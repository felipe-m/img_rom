--- Autcmatically generated VHDL ROM from a NES memory file----


---  Original memory dump file name: nespalette.pal --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_COLORS is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(6-1 downto 0);  --64 memory positions
    dout : out std_logic_vector(12-1 downto 0) -- memory data width
  );
end ROM_COLORS;

architecture BEHAVIORAL of ROM_COLORS is
  signal addr_int  : natural range 0 to 2**6-1;
  type memostruct is array (natural range<>) of std_logic_vector(12-1 downto 0);
  constant table_mem : memostruct := (
                    --    address   :    value 
                    --  dec -  hex  :  dec - hex(RGB)
    "010001000100", --    0 -  0x0  :  1092 - 0x444
    "000000000101", --    1 -  0x1  :     5 - 0x005
    "000000000111", --    2 -  0x2  :     7 - 0x007
    "000000000111", --    3 -  0x3  :     7 - 0x007
    "001100000100", --    4 -  0x4  :   772 - 0x304
    "010100000000", --    5 -  0x5  :  1280 - 0x500
    "010100000000", --    6 -  0x6  :  1280 - 0x500
    "010000000000", --    7 -  0x7  :  1024 - 0x400
    "000100000000", --    8 -  0x8  :   256 - 0x100
    "000000010000", --    9 -  0x9  :    16 - 0x010
    "000000010000", --   10 -  0xa  :    16 - 0x010
    "000000010000", --   11 -  0xb  :    16 - 0x010
    "000000010010", --   12 -  0xc  :    18 - 0x012
    "000000000000", --   13 -  0xd  :     0 - 0x000
    "000000000000", --   14 -  0xe  :     0 - 0x000
    "000000000000", --   15 -  0xf  :     0 - 0x000
    "100110011001", --   16 - 0x10  :  2457 - 0x999
    "000001001011", --   17 - 0x11  :    75 - 0x04B
    "000000111110", --   18 - 0x12  :    62 - 0x03E
    "010100011101", --   19 - 0x13  :  1309 - 0x51D
    "100100001010", --   20 - 0x14  :  2314 - 0x90A
    "110000000101", --   21 - 0x15  :  3077 - 0xC05
    "110000000000", --   22 - 0x16  :  3072 - 0xC00
    "101000100000", --   23 - 0x17  :  2592 - 0xA20
    "010100110000", --   24 - 0x18  :  1328 - 0x530
    "000001010000", --   25 - 0x19  :    80 - 0x050
    "000001100000", --   26 - 0x1a  :    96 - 0x060
    "000001100001", --   27 - 0x1b  :    97 - 0x061
    "000001010110", --   28 - 0x1c  :    86 - 0x056
    "000000000000", --   29 - 0x1d  :     0 - 0x000
    "000000000000", --   30 - 0x1e  :     0 - 0x000
    "000000000000", --   31 - 0x1f  :     0 - 0x000
    "111111111111", --   32 - 0x20  :  4095 - 0xFFF
    "000110011111", --   33 - 0x21  :   415 - 0x19F
    "010101111111", --   34 - 0x22  :  1407 - 0x57F
    "100101101111", --   35 - 0x23  :  2415 - 0x96F
    "111101101111", --   36 - 0x24  :  3951 - 0xF6F
    "111101101011", --   37 - 0x25  :  3947 - 0xF6B
    "111101110110", --   38 - 0x26  :  3958 - 0xF76
    "111110000001", --   39 - 0x27  :  3969 - 0xF81
    "110010010000", --   40 - 0x28  :  3216 - 0xC90
    "011110110000", --   41 - 0x29  :  1968 - 0x7B0
    "001011000010", --   42 - 0x2a  :   706 - 0x2C2
    "000011000111", --   43 - 0x2b  :   199 - 0x0C7
    "000010111101", --   44 - 0x2c  :   189 - 0x0BD
    "001000100010", --   45 - 0x2d  :   546 - 0x222
    "000000000000", --   46 - 0x2e  :     0 - 0x000
    "000000000000", --   47 - 0x2f  :     0 - 0x000
    "111111111111", --   48 - 0x30  :  4095 - 0xFFF
    "100111011111", --   49 - 0x31  :  2527 - 0x9DF
    "101011001111", --   50 - 0x32  :  2767 - 0xACF
    "110110111111", --   51 - 0x33  :  3519 - 0xDBF
    "111110111111", --   52 - 0x34  :  4031 - 0xFBF
    "111111001110", --   53 - 0x35  :  4046 - 0xFCE
    "111111001011", --   54 - 0x36  :  4043 - 0xFCB
    "111111001001", --   55 - 0x37  :  4041 - 0xFC9
    "111011011000", --   56 - 0x38  :  3800 - 0xED8
    "110011011000", --   57 - 0x39  :  3288 - 0xCD8
    "101011101010", --   58 - 0x3a  :  2794 - 0xAEA
    "100111101100", --   59 - 0x3b  :  2540 - 0x9EC
    "100111101110", --   60 - 0x3c  :  2542 - 0x9EE
    "101010101010", --   61 - 0x3d  :  2730 - 0xAAA
    "000000000000", --   62 - 0x3e  :     0 - 0x000
    "000000000000"  --   63 - 0x3f  :     0 - 0x000
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
