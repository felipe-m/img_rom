--- Autcmatically generated VHDL ROM from a NES memory file----
---   PATTERN TABLE
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


---  Original memory dump file name: donkeykong_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory with clock ------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_DONKEYKONG is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(13-1 downto 0);  --8192 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_DONKEYKONG;

architecture BEHAVIORAL of ROM_PTABLE_DONKEYKONG is
  signal addr_int  : natural range 0 to 2**13-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Pattern Table 0---------
    "00000000", --    0 -  0x0  :    0 - 0x0 -- Sprite 0x0
    "00000011", --    1 -  0x1  :    3 - 0x3
    "00000111", --    2 -  0x2  :    7 - 0x7
    "00000111", --    3 -  0x3  :    7 - 0x7
    "00001001", --    4 -  0x4  :    9 - 0x9
    "00001001", --    5 -  0x5  :    9 - 0x9
    "00011100", --    6 -  0x6  :   28 - 0x1c
    "00000000", --    7 -  0x7  :    0 - 0x0
    "00000000", --    8 -  0x8  :    0 - 0x0
    "00000011", --    9 -  0x9  :    3 - 0x3
    "00000111", --   10 -  0xa  :    7 - 0x7
    "00000000", --   11 -  0xb  :    0 - 0x0
    "00000110", --   12 -  0xc  :    6 - 0x6
    "00000110", --   13 -  0xd  :    6 - 0x6
    "00000011", --   14 -  0xe  :    3 - 0x3
    "00000011", --   15 -  0xf  :    3 - 0x3
    "00001111", --   16 - 0x10  :   15 - 0xf -- Sprite 0x1
    "00001111", --   17 - 0x11  :   15 - 0xf
    "00001111", --   18 - 0x12  :   15 - 0xf
    "11111111", --   19 - 0x13  :  255 - 0xff
    "11111111", --   20 - 0x14  :  255 - 0xff
    "11111100", --   21 - 0x15  :  252 - 0xfc
    "10000001", --   22 - 0x16  :  129 - 0x81
    "00000001", --   23 - 0x17  :    1 - 0x1
    "00000000", --   24 - 0x18  :    0 - 0x0
    "00010000", --   25 - 0x19  :   16 - 0x10
    "00111100", --   26 - 0x1a  :   60 - 0x3c
    "00111111", --   27 - 0x1b  :   63 - 0x3f
    "00111111", --   28 - 0x1c  :   63 - 0x3f
    "00111100", --   29 - 0x1d  :   60 - 0x3c
    "00000000", --   30 - 0x1e  :    0 - 0x0
    "00000000", --   31 - 0x1f  :    0 - 0x0
    "00000000", --   32 - 0x20  :    0 - 0x0 -- Sprite 0x2
    "11000000", --   33 - 0x21  :  192 - 0xc0
    "11111000", --   34 - 0x22  :  248 - 0xf8
    "10000000", --   35 - 0x23  :  128 - 0x80
    "00100000", --   36 - 0x24  :   32 - 0x20
    "10010000", --   37 - 0x25  :  144 - 0x90
    "00111100", --   38 - 0x26  :   60 - 0x3c
    "00000000", --   39 - 0x27  :    0 - 0x0
    "00000000", --   40 - 0x28  :    0 - 0x0
    "11000000", --   41 - 0x29  :  192 - 0xc0
    "11111000", --   42 - 0x2a  :  248 - 0xf8
    "01100000", --   43 - 0x2b  :   96 - 0x60
    "11011100", --   44 - 0x2c  :  220 - 0xdc
    "01101110", --   45 - 0x2d  :  110 - 0x6e
    "11000000", --   46 - 0x2e  :  192 - 0xc0
    "11111000", --   47 - 0x2f  :  248 - 0xf8
    "11000000", --   48 - 0x30  :  192 - 0xc0 -- Sprite 0x3
    "11000000", --   49 - 0x31  :  192 - 0xc0
    "11000000", --   50 - 0x32  :  192 - 0xc0
    "11110000", --   51 - 0x33  :  240 - 0xf0
    "11110000", --   52 - 0x34  :  240 - 0xf0
    "11100000", --   53 - 0x35  :  224 - 0xe0
    "11000000", --   54 - 0x36  :  192 - 0xc0
    "11100000", --   55 - 0x37  :  224 - 0xe0
    "01010000", --   56 - 0x38  :   80 - 0x50
    "00111000", --   57 - 0x39  :   56 - 0x38
    "00110000", --   58 - 0x3a  :   48 - 0x30
    "11110000", --   59 - 0x3b  :  240 - 0xf0
    "11110000", --   60 - 0x3c  :  240 - 0xf0
    "11100000", --   61 - 0x3d  :  224 - 0xe0
    "00000000", --   62 - 0x3e  :    0 - 0x0
    "00000000", --   63 - 0x3f  :    0 - 0x0
    "00000111", --   64 - 0x40  :    7 - 0x7 -- Sprite 0x4
    "00001111", --   65 - 0x41  :   15 - 0xf
    "00001111", --   66 - 0x42  :   15 - 0xf
    "00010010", --   67 - 0x43  :   18 - 0x12
    "00010011", --   68 - 0x44  :   19 - 0x13
    "00111000", --   69 - 0x45  :   56 - 0x38
    "00000000", --   70 - 0x46  :    0 - 0x0
    "00001111", --   71 - 0x47  :   15 - 0xf
    "00000111", --   72 - 0x48  :    7 - 0x7
    "00001111", --   73 - 0x49  :   15 - 0xf
    "00000000", --   74 - 0x4a  :    0 - 0x0
    "00001101", --   75 - 0x4b  :   13 - 0xd
    "00001100", --   76 - 0x4c  :   12 - 0xc
    "00000111", --   77 - 0x4d  :    7 - 0x7
    "00000111", --   78 - 0x4e  :    7 - 0x7
    "00000000", --   79 - 0x4f  :    0 - 0x0
    "00011111", --   80 - 0x50  :   31 - 0x1f -- Sprite 0x5
    "00011111", --   81 - 0x51  :   31 - 0x1f
    "00011111", --   82 - 0x52  :   31 - 0x1f
    "00011000", --   83 - 0x53  :   24 - 0x18
    "00011001", --   84 - 0x54  :   25 - 0x19
    "00011110", --   85 - 0x55  :   30 - 0x1e
    "00011100", --   86 - 0x56  :   28 - 0x1c
    "00011110", --   87 - 0x57  :   30 - 0x1e
    "00000001", --   88 - 0x58  :    1 - 0x1
    "00000011", --   89 - 0x59  :    3 - 0x3
    "00000001", --   90 - 0x5a  :    1 - 0x1
    "00010111", --   91 - 0x5b  :   23 - 0x17
    "00011111", --   92 - 0x5c  :   31 - 0x1f
    "00011110", --   93 - 0x5d  :   30 - 0x1e
    "00000000", --   94 - 0x5e  :    0 - 0x0
    "00000000", --   95 - 0x5f  :    0 - 0x0
    "10000000", --   96 - 0x60  :  128 - 0x80 -- Sprite 0x6
    "11110000", --   97 - 0x61  :  240 - 0xf0
    "00000000", --   98 - 0x62  :    0 - 0x0
    "01000000", --   99 - 0x63  :   64 - 0x40
    "00100000", --  100 - 0x64  :   32 - 0x20
    "01111000", --  101 - 0x65  :  120 - 0x78
    "00000000", --  102 - 0x66  :    0 - 0x0
    "11000000", --  103 - 0x67  :  192 - 0xc0
    "10000000", --  104 - 0x68  :  128 - 0x80
    "11110000", --  105 - 0x69  :  240 - 0xf0
    "11000000", --  106 - 0x6a  :  192 - 0xc0
    "10111000", --  107 - 0x6b  :  184 - 0xb8
    "11011100", --  108 - 0x6c  :  220 - 0xdc
    "10000000", --  109 - 0x6d  :  128 - 0x80
    "11110000", --  110 - 0x6e  :  240 - 0xf0
    "00000000", --  111 - 0x6f  :    0 - 0x0
    "11100000", --  112 - 0x70  :  224 - 0xe0 -- Sprite 0x7
    "01100000", --  113 - 0x71  :   96 - 0x60
    "11110000", --  114 - 0x72  :  240 - 0xf0
    "11110000", --  115 - 0x73  :  240 - 0xf0
    "11110000", --  116 - 0x74  :  240 - 0xf0
    "11100000", --  117 - 0x75  :  224 - 0xe0
    "11100000", --  118 - 0x76  :  224 - 0xe0
    "11110000", --  119 - 0x77  :  240 - 0xf0
    "10000000", --  120 - 0x78  :  128 - 0x80
    "11100000", --  121 - 0x79  :  224 - 0xe0
    "11110000", --  122 - 0x7a  :  240 - 0xf0
    "11110000", --  123 - 0x7b  :  240 - 0xf0
    "11110000", --  124 - 0x7c  :  240 - 0xf0
    "11100000", --  125 - 0x7d  :  224 - 0xe0
    "00000000", --  126 - 0x7e  :    0 - 0x0
    "00000000", --  127 - 0x7f  :    0 - 0x0
    "00000111", --  128 - 0x80  :    7 - 0x7 -- Sprite 0x8
    "00001111", --  129 - 0x81  :   15 - 0xf
    "00001111", --  130 - 0x82  :   15 - 0xf
    "00010010", --  131 - 0x83  :   18 - 0x12
    "00010011", --  132 - 0x84  :   19 - 0x13
    "00111000", --  133 - 0x85  :   56 - 0x38
    "00000000", --  134 - 0x86  :    0 - 0x0
    "00111111", --  135 - 0x87  :   63 - 0x3f
    "00000111", --  136 - 0x88  :    7 - 0x7
    "00001111", --  137 - 0x89  :   15 - 0xf
    "00000000", --  138 - 0x8a  :    0 - 0x0
    "00001101", --  139 - 0x8b  :   13 - 0xd
    "00001100", --  140 - 0x8c  :   12 - 0xc
    "00000111", --  141 - 0x8d  :    7 - 0x7
    "00000111", --  142 - 0x8e  :    7 - 0x7
    "00000011", --  143 - 0x8f  :    3 - 0x3
    "00111111", --  144 - 0x90  :   63 - 0x3f -- Sprite 0x9
    "00001110", --  145 - 0x91  :   14 - 0xe
    "00001111", --  146 - 0x92  :   15 - 0xf
    "00011111", --  147 - 0x93  :   31 - 0x1f
    "00111111", --  148 - 0x94  :   63 - 0x3f
    "01111100", --  149 - 0x95  :  124 - 0x7c
    "01110000", --  150 - 0x96  :  112 - 0x70
    "00111000", --  151 - 0x97  :   56 - 0x38
    "11000011", --  152 - 0x98  :  195 - 0xc3
    "11100011", --  153 - 0x99  :  227 - 0xe3
    "11001111", --  154 - 0x9a  :  207 - 0xcf
    "00011111", --  155 - 0x9b  :   31 - 0x1f
    "00111111", --  156 - 0x9c  :   63 - 0x3f
    "00001100", --  157 - 0x9d  :   12 - 0xc
    "00000000", --  158 - 0x9e  :    0 - 0x0
    "00000000", --  159 - 0x9f  :    0 - 0x0
    "10000000", --  160 - 0xa0  :  128 - 0x80 -- Sprite 0xa
    "11110000", --  161 - 0xa1  :  240 - 0xf0
    "00000000", --  162 - 0xa2  :    0 - 0x0
    "01000000", --  163 - 0xa3  :   64 - 0x40
    "00100000", --  164 - 0xa4  :   32 - 0x20
    "01111000", --  165 - 0xa5  :  120 - 0x78
    "00000000", --  166 - 0xa6  :    0 - 0x0
    "11000000", --  167 - 0xa7  :  192 - 0xc0
    "10000000", --  168 - 0xa8  :  128 - 0x80
    "11110000", --  169 - 0xa9  :  240 - 0xf0
    "11000000", --  170 - 0xaa  :  192 - 0xc0
    "10111000", --  171 - 0xab  :  184 - 0xb8
    "11011100", --  172 - 0xac  :  220 - 0xdc
    "10000000", --  173 - 0xad  :  128 - 0x80
    "11110000", --  174 - 0xae  :  240 - 0xf0
    "00000110", --  175 - 0xaf  :    6 - 0x6
    "11110000", --  176 - 0xb0  :  240 - 0xf0 -- Sprite 0xb
    "11111000", --  177 - 0xb1  :  248 - 0xf8
    "11100100", --  178 - 0xb2  :  228 - 0xe4
    "11111100", --  179 - 0xb3  :  252 - 0xfc
    "11111100", --  180 - 0xb4  :  252 - 0xfc
    "01111100", --  181 - 0xb5  :  124 - 0x7c
    "00000000", --  182 - 0xb6  :    0 - 0x0
    "00000000", --  183 - 0xb7  :    0 - 0x0
    "10001110", --  184 - 0xb8  :  142 - 0x8e
    "11100110", --  185 - 0xb9  :  230 - 0xe6
    "11100000", --  186 - 0xba  :  224 - 0xe0
    "11110000", --  187 - 0xbb  :  240 - 0xf0
    "11110000", --  188 - 0xbc  :  240 - 0xf0
    "01110000", --  189 - 0xbd  :  112 - 0x70
    "00000000", --  190 - 0xbe  :    0 - 0x0
    "00000000", --  191 - 0xbf  :    0 - 0x0
    "00000000", --  192 - 0xc0  :    0 - 0x0 -- Sprite 0xc
    "00000010", --  193 - 0xc1  :    2 - 0x2
    "00000110", --  194 - 0xc2  :    6 - 0x6
    "00000111", --  195 - 0xc3  :    7 - 0x7
    "00001001", --  196 - 0xc4  :    9 - 0x9
    "00001001", --  197 - 0xc5  :    9 - 0x9
    "00011101", --  198 - 0xc6  :   29 - 0x1d
    "00000011", --  199 - 0xc7  :    3 - 0x3
    "00000001", --  200 - 0xc8  :    1 - 0x1
    "00000011", --  201 - 0xc9  :    3 - 0x3
    "00000111", --  202 - 0xca  :    7 - 0x7
    "00000000", --  203 - 0xcb  :    0 - 0x0
    "00000110", --  204 - 0xcc  :    6 - 0x6
    "00000110", --  205 - 0xcd  :    6 - 0x6
    "00000010", --  206 - 0xce  :    2 - 0x2
    "00000000", --  207 - 0xcf  :    0 - 0x0
    "00001111", --  208 - 0xd0  :   15 - 0xf -- Sprite 0xd
    "00001111", --  209 - 0xd1  :   15 - 0xf
    "00001111", --  210 - 0xd2  :   15 - 0xf
    "11111111", --  211 - 0xd3  :  255 - 0xff
    "11111111", --  212 - 0xd4  :  255 - 0xff
    "11111100", --  213 - 0xd5  :  252 - 0xfc
    "10000001", --  214 - 0xd6  :  129 - 0x81
    "00000001", --  215 - 0xd7  :    1 - 0x1
    "00000000", --  216 - 0xd8  :    0 - 0x0
    "00000000", --  217 - 0xd9  :    0 - 0x0
    "00001100", --  218 - 0xda  :   12 - 0xc
    "00111111", --  219 - 0xdb  :   63 - 0x3f
    "00111111", --  220 - 0xdc  :   63 - 0x3f
    "00111100", --  221 - 0xdd  :   60 - 0x3c
    "00000000", --  222 - 0xde  :    0 - 0x0
    "00000000", --  223 - 0xdf  :    0 - 0x0
    "00000000", --  224 - 0xe0  :    0 - 0x0 -- Sprite 0xe
    "00000000", --  225 - 0xe1  :    0 - 0x0
    "00111000", --  226 - 0xe2  :   56 - 0x38
    "11000000", --  227 - 0xe3  :  192 - 0xc0
    "11100000", --  228 - 0xe4  :  224 - 0xe0
    "11010000", --  229 - 0xe5  :  208 - 0xd0
    "11111100", --  230 - 0xe6  :  252 - 0xfc
    "11000000", --  231 - 0xe7  :  192 - 0xc0
    "11000000", --  232 - 0xe8  :  192 - 0xc0
    "11000000", --  233 - 0xe9  :  192 - 0xc0
    "11111000", --  234 - 0xea  :  248 - 0xf8
    "00100000", --  235 - 0xeb  :   32 - 0x20
    "00011100", --  236 - 0xec  :   28 - 0x1c
    "00101110", --  237 - 0xed  :   46 - 0x2e
    "00000000", --  238 - 0xee  :    0 - 0x0
    "00111000", --  239 - 0xef  :   56 - 0x38
    "11100000", --  240 - 0xf0  :  224 - 0xe0 -- Sprite 0xf
    "11100000", --  241 - 0xf1  :  224 - 0xe0
    "10110000", --  242 - 0xf2  :  176 - 0xb0
    "11110000", --  243 - 0xf3  :  240 - 0xf0
    "11110000", --  244 - 0xf4  :  240 - 0xf0
    "11100000", --  245 - 0xf5  :  224 - 0xe0
    "11000000", --  246 - 0xf6  :  192 - 0xc0
    "11100000", --  247 - 0xf7  :  224 - 0xe0
    "00000000", --  248 - 0xf8  :    0 - 0x0
    "01100000", --  249 - 0xf9  :   96 - 0x60
    "11110000", --  250 - 0xfa  :  240 - 0xf0
    "11110000", --  251 - 0xfb  :  240 - 0xf0
    "11110000", --  252 - 0xfc  :  240 - 0xf0
    "11100000", --  253 - 0xfd  :  224 - 0xe0
    "00000000", --  254 - 0xfe  :    0 - 0x0
    "00000000", --  255 - 0xff  :    0 - 0x0
    "00000000", --  256 - 0x100  :    0 - 0x0 -- Sprite 0x10
    "00000011", --  257 - 0x101  :    3 - 0x3
    "00000111", --  258 - 0x102  :    7 - 0x7
    "00000111", --  259 - 0x103  :    7 - 0x7
    "00001001", --  260 - 0x104  :    9 - 0x9
    "00001001", --  261 - 0x105  :    9 - 0x9
    "00011100", --  262 - 0x106  :   28 - 0x1c
    "00000000", --  263 - 0x107  :    0 - 0x0
    "00000000", --  264 - 0x108  :    0 - 0x0
    "00000011", --  265 - 0x109  :    3 - 0x3
    "00000111", --  266 - 0x10a  :    7 - 0x7
    "00000000", --  267 - 0x10b  :    0 - 0x0
    "00000110", --  268 - 0x10c  :    6 - 0x6
    "00000110", --  269 - 0x10d  :    6 - 0x6
    "00000011", --  270 - 0x10e  :    3 - 0x3
    "00000011", --  271 - 0x10f  :    3 - 0x3
    "00001111", --  272 - 0x110  :   15 - 0xf -- Sprite 0x11
    "00001111", --  273 - 0x111  :   15 - 0xf
    "00001111", --  274 - 0x112  :   15 - 0xf
    "11111111", --  275 - 0x113  :  255 - 0xff
    "11111111", --  276 - 0x114  :  255 - 0xff
    "11111100", --  277 - 0x115  :  252 - 0xfc
    "10000001", --  278 - 0x116  :  129 - 0x81
    "00000001", --  279 - 0x117  :    1 - 0x1
    "00000000", --  280 - 0x118  :    0 - 0x0
    "00000000", --  281 - 0x119  :    0 - 0x0
    "00001100", --  282 - 0x11a  :   12 - 0xc
    "00111111", --  283 - 0x11b  :   63 - 0x3f
    "00111111", --  284 - 0x11c  :   63 - 0x3f
    "00111100", --  285 - 0x11d  :   60 - 0x3c
    "00000000", --  286 - 0x11e  :    0 - 0x0
    "00000000", --  287 - 0x11f  :    0 - 0x0
    "00000000", --  288 - 0x120  :    0 - 0x0 -- Sprite 0x12
    "11000000", --  289 - 0x121  :  192 - 0xc0
    "11111000", --  290 - 0x122  :  248 - 0xf8
    "10000000", --  291 - 0x123  :  128 - 0x80
    "00100000", --  292 - 0x124  :   32 - 0x20
    "10010000", --  293 - 0x125  :  144 - 0x90
    "00111100", --  294 - 0x126  :   60 - 0x3c
    "00000000", --  295 - 0x127  :    0 - 0x0
    "00000000", --  296 - 0x128  :    0 - 0x0
    "11000000", --  297 - 0x129  :  192 - 0xc0
    "11111000", --  298 - 0x12a  :  248 - 0xf8
    "01100000", --  299 - 0x12b  :   96 - 0x60
    "11011100", --  300 - 0x12c  :  220 - 0xdc
    "01101110", --  301 - 0x12d  :  110 - 0x6e
    "11000000", --  302 - 0x12e  :  192 - 0xc0
    "11111000", --  303 - 0x12f  :  248 - 0xf8
    "11100000", --  304 - 0x130  :  224 - 0xe0 -- Sprite 0x13
    "11110000", --  305 - 0x131  :  240 - 0xf0
    "11110000", --  306 - 0x132  :  240 - 0xf0
    "11110000", --  307 - 0x133  :  240 - 0xf0
    "11110000", --  308 - 0x134  :  240 - 0xf0
    "11100000", --  309 - 0x135  :  224 - 0xe0
    "11000000", --  310 - 0x136  :  192 - 0xc0
    "11100000", --  311 - 0x137  :  224 - 0xe0
    "01000111", --  312 - 0x138  :   71 - 0x47
    "00001111", --  313 - 0x139  :   15 - 0xf
    "00001110", --  314 - 0x13a  :   14 - 0xe
    "11110000", --  315 - 0x13b  :  240 - 0xf0
    "11110000", --  316 - 0x13c  :  240 - 0xf0
    "11100000", --  317 - 0x13d  :  224 - 0xe0
    "00000000", --  318 - 0x13e  :    0 - 0x0
    "00000000", --  319 - 0x13f  :    0 - 0x0
    "00000100", --  320 - 0x140  :    4 - 0x4 -- Sprite 0x14
    "00001100", --  321 - 0x141  :   12 - 0xc
    "00001100", --  322 - 0x142  :   12 - 0xc
    "00010011", --  323 - 0x143  :   19 - 0x13
    "00010011", --  324 - 0x144  :   19 - 0x13
    "00111011", --  325 - 0x145  :   59 - 0x3b
    "00000111", --  326 - 0x146  :    7 - 0x7
    "00001111", --  327 - 0x147  :   15 - 0xf
    "00000111", --  328 - 0x148  :    7 - 0x7
    "00001111", --  329 - 0x149  :   15 - 0xf
    "00000011", --  330 - 0x14a  :    3 - 0x3
    "00001100", --  331 - 0x14b  :   12 - 0xc
    "00001100", --  332 - 0x14c  :   12 - 0xc
    "00000100", --  333 - 0x14d  :    4 - 0x4
    "00000000", --  334 - 0x14e  :    0 - 0x0
    "00000000", --  335 - 0x14f  :    0 - 0x0
    "00001111", --  336 - 0x150  :   15 - 0xf -- Sprite 0x15
    "00001111", --  337 - 0x151  :   15 - 0xf
    "00001111", --  338 - 0x152  :   15 - 0xf
    "00011111", --  339 - 0x153  :   31 - 0x1f
    "00011111", --  340 - 0x154  :   31 - 0x1f
    "00011110", --  341 - 0x155  :   30 - 0x1e
    "00011100", --  342 - 0x156  :   28 - 0x1c
    "00011110", --  343 - 0x157  :   30 - 0x1e
    "00000000", --  344 - 0x158  :    0 - 0x0
    "00000001", --  345 - 0x159  :    1 - 0x1
    "00001111", --  346 - 0x15a  :   15 - 0xf
    "00011111", --  347 - 0x15b  :   31 - 0x1f
    "00011111", --  348 - 0x15c  :   31 - 0x1f
    "00011110", --  349 - 0x15d  :   30 - 0x1e
    "00000000", --  350 - 0x15e  :    0 - 0x0
    "00000000", --  351 - 0x15f  :    0 - 0x0
    "00000000", --  352 - 0x160  :    0 - 0x0 -- Sprite 0x16
    "01110000", --  353 - 0x161  :  112 - 0x70
    "00000000", --  354 - 0x162  :    0 - 0x0
    "11000000", --  355 - 0x163  :  192 - 0xc0
    "10100000", --  356 - 0x164  :  160 - 0xa0
    "11111000", --  357 - 0x165  :  248 - 0xf8
    "10000000", --  358 - 0x166  :  128 - 0x80
    "11000000", --  359 - 0x167  :  192 - 0xc0
    "10000000", --  360 - 0x168  :  128 - 0x80
    "11110000", --  361 - 0x169  :  240 - 0xf0
    "11000000", --  362 - 0x16a  :  192 - 0xc0
    "00111000", --  363 - 0x16b  :   56 - 0x38
    "01011100", --  364 - 0x16c  :   92 - 0x5c
    "00000000", --  365 - 0x16d  :    0 - 0x0
    "01110000", --  366 - 0x16e  :  112 - 0x70
    "01000000", --  367 - 0x16f  :   64 - 0x40
    "11100000", --  368 - 0x170  :  224 - 0xe0 -- Sprite 0x17
    "01100000", --  369 - 0x171  :   96 - 0x60
    "11110000", --  370 - 0x172  :  240 - 0xf0
    "11110000", --  371 - 0x173  :  240 - 0xf0
    "11110000", --  372 - 0x174  :  240 - 0xf0
    "11100000", --  373 - 0x175  :  224 - 0xe0
    "11100000", --  374 - 0x176  :  224 - 0xe0
    "11110000", --  375 - 0x177  :  240 - 0xf0
    "11000000", --  376 - 0x178  :  192 - 0xc0
    "11100000", --  377 - 0x179  :  224 - 0xe0
    "11110000", --  378 - 0x17a  :  240 - 0xf0
    "11110000", --  379 - 0x17b  :  240 - 0xf0
    "11110000", --  380 - 0x17c  :  240 - 0xf0
    "11100000", --  381 - 0x17d  :  224 - 0xe0
    "00000000", --  382 - 0x17e  :    0 - 0x0
    "00000000", --  383 - 0x17f  :    0 - 0x0
    "00000111", --  384 - 0x180  :    7 - 0x7 -- Sprite 0x18
    "00001111", --  385 - 0x181  :   15 - 0xf
    "00001111", --  386 - 0x182  :   15 - 0xf
    "00010010", --  387 - 0x183  :   18 - 0x12
    "00010011", --  388 - 0x184  :   19 - 0x13
    "00111000", --  389 - 0x185  :   56 - 0x38
    "00000000", --  390 - 0x186  :    0 - 0x0
    "00001111", --  391 - 0x187  :   15 - 0xf
    "00000111", --  392 - 0x188  :    7 - 0x7
    "00001111", --  393 - 0x189  :   15 - 0xf
    "00000000", --  394 - 0x18a  :    0 - 0x0
    "00001101", --  395 - 0x18b  :   13 - 0xd
    "00001100", --  396 - 0x18c  :   12 - 0xc
    "00000111", --  397 - 0x18d  :    7 - 0x7
    "00000111", --  398 - 0x18e  :    7 - 0x7
    "00000001", --  399 - 0x18f  :    1 - 0x1
    "00011111", --  400 - 0x190  :   31 - 0x1f -- Sprite 0x19
    "00011111", --  401 - 0x191  :   31 - 0x1f
    "00011111", --  402 - 0x192  :   31 - 0x1f
    "00011111", --  403 - 0x193  :   31 - 0x1f
    "00011111", --  404 - 0x194  :   31 - 0x1f
    "00011110", --  405 - 0x195  :   30 - 0x1e
    "00011100", --  406 - 0x196  :   28 - 0x1c
    "00011110", --  407 - 0x197  :   30 - 0x1e
    "00000000", --  408 - 0x198  :    0 - 0x0
    "00000000", --  409 - 0x199  :    0 - 0x0
    "00010011", --  410 - 0x19a  :   19 - 0x13
    "00011111", --  411 - 0x19b  :   31 - 0x1f
    "00011111", --  412 - 0x19c  :   31 - 0x1f
    "00011110", --  413 - 0x19d  :   30 - 0x1e
    "00000000", --  414 - 0x19e  :    0 - 0x0
    "00000000", --  415 - 0x19f  :    0 - 0x0
    "10000000", --  416 - 0x1a0  :  128 - 0x80 -- Sprite 0x1a
    "11110000", --  417 - 0x1a1  :  240 - 0xf0
    "00000000", --  418 - 0x1a2  :    0 - 0x0
    "01000000", --  419 - 0x1a3  :   64 - 0x40
    "00100000", --  420 - 0x1a4  :   32 - 0x20
    "01111000", --  421 - 0x1a5  :  120 - 0x78
    "00000000", --  422 - 0x1a6  :    0 - 0x0
    "11000000", --  423 - 0x1a7  :  192 - 0xc0
    "10000000", --  424 - 0x1a8  :  128 - 0x80
    "11110000", --  425 - 0x1a9  :  240 - 0xf0
    "11000000", --  426 - 0x1aa  :  192 - 0xc0
    "10111000", --  427 - 0x1ab  :  184 - 0xb8
    "11011100", --  428 - 0x1ac  :  220 - 0xdc
    "10000000", --  429 - 0x1ad  :  128 - 0x80
    "11110000", --  430 - 0x1ae  :  240 - 0xf0
    "10000000", --  431 - 0x1af  :  128 - 0x80
    "11111000", --  432 - 0x1b0  :  248 - 0xf8 -- Sprite 0x1b
    "11111000", --  433 - 0x1b1  :  248 - 0xf8
    "11110000", --  434 - 0x1b2  :  240 - 0xf0
    "11110000", --  435 - 0x1b3  :  240 - 0xf0
    "11110000", --  436 - 0x1b4  :  240 - 0xf0
    "11100000", --  437 - 0x1b5  :  224 - 0xe0
    "11100000", --  438 - 0x1b6  :  224 - 0xe0
    "11110000", --  439 - 0x1b7  :  240 - 0xf0
    "00000111", --  440 - 0x1b8  :    7 - 0x7
    "00000111", --  441 - 0x1b9  :    7 - 0x7
    "11111110", --  442 - 0x1ba  :  254 - 0xfe
    "11110000", --  443 - 0x1bb  :  240 - 0xf0
    "11110000", --  444 - 0x1bc  :  240 - 0xf0
    "11100000", --  445 - 0x1bd  :  224 - 0xe0
    "00000000", --  446 - 0x1be  :    0 - 0x0
    "00000000", --  447 - 0x1bf  :    0 - 0x0
    "00000100", --  448 - 0x1c0  :    4 - 0x4 -- Sprite 0x1c
    "00001100", --  449 - 0x1c1  :   12 - 0xc
    "00001100", --  450 - 0x1c2  :   12 - 0xc
    "00010011", --  451 - 0x1c3  :   19 - 0x13
    "00010011", --  452 - 0x1c4  :   19 - 0x13
    "00111111", --  453 - 0x1c5  :   63 - 0x3f
    "00000111", --  454 - 0x1c6  :    7 - 0x7
    "00001111", --  455 - 0x1c7  :   15 - 0xf
    "00000111", --  456 - 0x1c8  :    7 - 0x7
    "00001111", --  457 - 0x1c9  :   15 - 0xf
    "00000011", --  458 - 0x1ca  :    3 - 0x3
    "00001100", --  459 - 0x1cb  :   12 - 0xc
    "00001100", --  460 - 0x1cc  :   12 - 0xc
    "00000000", --  461 - 0x1cd  :    0 - 0x0
    "00000000", --  462 - 0x1ce  :    0 - 0x0
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "00001111", --  464 - 0x1d0  :   15 - 0xf -- Sprite 0x1d
    "00001111", --  465 - 0x1d1  :   15 - 0xf
    "00001111", --  466 - 0x1d2  :   15 - 0xf
    "00011111", --  467 - 0x1d3  :   31 - 0x1f
    "00111111", --  468 - 0x1d4  :   63 - 0x3f
    "01111100", --  469 - 0x1d5  :  124 - 0x7c
    "01110000", --  470 - 0x1d6  :  112 - 0x70
    "00111000", --  471 - 0x1d7  :   56 - 0x38
    "00000001", --  472 - 0x1d8  :    1 - 0x1
    "00000001", --  473 - 0x1d9  :    1 - 0x1
    "00001111", --  474 - 0x1da  :   15 - 0xf
    "00011111", --  475 - 0x1db  :   31 - 0x1f
    "00111111", --  476 - 0x1dc  :   63 - 0x3f
    "00011100", --  477 - 0x1dd  :   28 - 0x1c
    "00000000", --  478 - 0x1de  :    0 - 0x0
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "00000000", --  480 - 0x1e0  :    0 - 0x0 -- Sprite 0x1e
    "01110000", --  481 - 0x1e1  :  112 - 0x70
    "00000000", --  482 - 0x1e2  :    0 - 0x0
    "11000000", --  483 - 0x1e3  :  192 - 0xc0
    "10100000", --  484 - 0x1e4  :  160 - 0xa0
    "11111000", --  485 - 0x1e5  :  248 - 0xf8
    "10000000", --  486 - 0x1e6  :  128 - 0x80
    "11000000", --  487 - 0x1e7  :  192 - 0xc0
    "10000000", --  488 - 0x1e8  :  128 - 0x80
    "11110000", --  489 - 0x1e9  :  240 - 0xf0
    "11000000", --  490 - 0x1ea  :  192 - 0xc0
    "00111000", --  491 - 0x1eb  :   56 - 0x38
    "01011100", --  492 - 0x1ec  :   92 - 0x5c
    "00000000", --  493 - 0x1ed  :    0 - 0x0
    "01110000", --  494 - 0x1ee  :  112 - 0x70
    "01000000", --  495 - 0x1ef  :   64 - 0x40
    "11000000", --  496 - 0x1f0  :  192 - 0xc0 -- Sprite 0x1f
    "01100000", --  497 - 0x1f1  :   96 - 0x60
    "11100100", --  498 - 0x1f2  :  228 - 0xe4
    "11111100", --  499 - 0x1f3  :  252 - 0xfc
    "11111100", --  500 - 0x1f4  :  252 - 0xfc
    "01111100", --  501 - 0x1f5  :  124 - 0x7c
    "00000000", --  502 - 0x1f6  :    0 - 0x0
    "00000000", --  503 - 0x1f7  :    0 - 0x0
    "11000000", --  504 - 0x1f8  :  192 - 0xc0
    "11100000", --  505 - 0x1f9  :  224 - 0xe0
    "11100000", --  506 - 0x1fa  :  224 - 0xe0
    "11110000", --  507 - 0x1fb  :  240 - 0xf0
    "11110000", --  508 - 0x1fc  :  240 - 0xf0
    "01110000", --  509 - 0x1fd  :  112 - 0x70
    "00000000", --  510 - 0x1fe  :    0 - 0x0
    "00000000", --  511 - 0x1ff  :    0 - 0x0
    "00000111", --  512 - 0x200  :    7 - 0x7 -- Sprite 0x20
    "00001111", --  513 - 0x201  :   15 - 0xf
    "00001111", --  514 - 0x202  :   15 - 0xf
    "00010010", --  515 - 0x203  :   18 - 0x12
    "00010011", --  516 - 0x204  :   19 - 0x13
    "00111000", --  517 - 0x205  :   56 - 0x38
    "00000000", --  518 - 0x206  :    0 - 0x0
    "00000111", --  519 - 0x207  :    7 - 0x7
    "00000111", --  520 - 0x208  :    7 - 0x7
    "00001111", --  521 - 0x209  :   15 - 0xf
    "00000000", --  522 - 0x20a  :    0 - 0x0
    "00001101", --  523 - 0x20b  :   13 - 0xd
    "00001100", --  524 - 0x20c  :   12 - 0xc
    "00000111", --  525 - 0x20d  :    7 - 0x7
    "00000111", --  526 - 0x20e  :    7 - 0x7
    "00000001", --  527 - 0x20f  :    1 - 0x1
    "00001111", --  528 - 0x210  :   15 - 0xf -- Sprite 0x21
    "00001111", --  529 - 0x211  :   15 - 0xf
    "00001111", --  530 - 0x212  :   15 - 0xf
    "00011111", --  531 - 0x213  :   31 - 0x1f
    "00111111", --  532 - 0x214  :   63 - 0x3f
    "01111100", --  533 - 0x215  :  124 - 0x7c
    "01110000", --  534 - 0x216  :  112 - 0x70
    "00111000", --  535 - 0x217  :   56 - 0x38
    "00000000", --  536 - 0x218  :    0 - 0x0
    "00000000", --  537 - 0x219  :    0 - 0x0
    "00001001", --  538 - 0x21a  :    9 - 0x9
    "00011111", --  539 - 0x21b  :   31 - 0x1f
    "00111111", --  540 - 0x21c  :   63 - 0x3f
    "00011100", --  541 - 0x21d  :   28 - 0x1c
    "00000000", --  542 - 0x21e  :    0 - 0x0
    "00000000", --  543 - 0x21f  :    0 - 0x0
    "10000000", --  544 - 0x220  :  128 - 0x80 -- Sprite 0x22
    "11110000", --  545 - 0x221  :  240 - 0xf0
    "00000000", --  546 - 0x222  :    0 - 0x0
    "01000000", --  547 - 0x223  :   64 - 0x40
    "00100000", --  548 - 0x224  :   32 - 0x20
    "01111000", --  549 - 0x225  :  120 - 0x78
    "00000000", --  550 - 0x226  :    0 - 0x0
    "11000000", --  551 - 0x227  :  192 - 0xc0
    "10000000", --  552 - 0x228  :  128 - 0x80
    "11110000", --  553 - 0x229  :  240 - 0xf0
    "11000000", --  554 - 0x22a  :  192 - 0xc0
    "10111000", --  555 - 0x22b  :  184 - 0xb8
    "11011100", --  556 - 0x22c  :  220 - 0xdc
    "10000000", --  557 - 0x22d  :  128 - 0x80
    "11110000", --  558 - 0x22e  :  240 - 0xf0
    "10000000", --  559 - 0x22f  :  128 - 0x80
    "11111000", --  560 - 0x230  :  248 - 0xf8 -- Sprite 0x23
    "11111000", --  561 - 0x231  :  248 - 0xf8
    "11100000", --  562 - 0x232  :  224 - 0xe0
    "11111100", --  563 - 0x233  :  252 - 0xfc
    "11111100", --  564 - 0x234  :  252 - 0xfc
    "01111100", --  565 - 0x235  :  124 - 0x7c
    "00000000", --  566 - 0x236  :    0 - 0x0
    "00000000", --  567 - 0x237  :    0 - 0x0
    "00000111", --  568 - 0x238  :    7 - 0x7
    "00000111", --  569 - 0x239  :    7 - 0x7
    "11101110", --  570 - 0x23a  :  238 - 0xee
    "11110000", --  571 - 0x23b  :  240 - 0xf0
    "11110000", --  572 - 0x23c  :  240 - 0xf0
    "01110000", --  573 - 0x23d  :  112 - 0x70
    "00000000", --  574 - 0x23e  :    0 - 0x0
    "00000000", --  575 - 0x23f  :    0 - 0x0
    "00000000", --  576 - 0x240  :    0 - 0x0 -- Sprite 0x24
    "00000111", --  577 - 0x241  :    7 - 0x7
    "00000111", --  578 - 0x242  :    7 - 0x7
    "00001111", --  579 - 0x243  :   15 - 0xf
    "00001111", --  580 - 0x244  :   15 - 0xf
    "00111000", --  581 - 0x245  :   56 - 0x38
    "01111111", --  582 - 0x246  :  127 - 0x7f
    "01111111", --  583 - 0x247  :  127 - 0x7f
    "00000000", --  584 - 0x248  :    0 - 0x0
    "00000111", --  585 - 0x249  :    7 - 0x7
    "00000011", --  586 - 0x24a  :    3 - 0x3
    "00000000", --  587 - 0x24b  :    0 - 0x0
    "00000000", --  588 - 0x24c  :    0 - 0x0
    "00000111", --  589 - 0x24d  :    7 - 0x7
    "00000100", --  590 - 0x24e  :    4 - 0x4
    "00000100", --  591 - 0x24f  :    4 - 0x4
    "00011111", --  592 - 0x250  :   31 - 0x1f -- Sprite 0x25
    "00011111", --  593 - 0x251  :   31 - 0x1f
    "00011111", --  594 - 0x252  :   31 - 0x1f
    "00011111", --  595 - 0x253  :   31 - 0x1f
    "00001111", --  596 - 0x254  :   15 - 0xf
    "00001111", --  597 - 0x255  :   15 - 0xf
    "00001111", --  598 - 0x256  :   15 - 0xf
    "00000111", --  599 - 0x257  :    7 - 0x7
    "00011110", --  600 - 0x258  :   30 - 0x1e
    "00011111", --  601 - 0x259  :   31 - 0x1f
    "00011111", --  602 - 0x25a  :   31 - 0x1f
    "00011111", --  603 - 0x25b  :   31 - 0x1f
    "00001111", --  604 - 0x25c  :   15 - 0xf
    "00001000", --  605 - 0x25d  :    8 - 0x8
    "00000000", --  606 - 0x25e  :    0 - 0x0
    "00000000", --  607 - 0x25f  :    0 - 0x0
    "00000000", --  608 - 0x260  :    0 - 0x0 -- Sprite 0x26
    "11100000", --  609 - 0x261  :  224 - 0xe0
    "11111000", --  610 - 0x262  :  248 - 0xf8
    "11111100", --  611 - 0x263  :  252 - 0xfc
    "11111100", --  612 - 0x264  :  252 - 0xfc
    "00011100", --  613 - 0x265  :   28 - 0x1c
    "11111000", --  614 - 0x266  :  248 - 0xf8
    "11111000", --  615 - 0x267  :  248 - 0xf8
    "00111000", --  616 - 0x268  :   56 - 0x38
    "11111000", --  617 - 0x269  :  248 - 0xf8
    "11000000", --  618 - 0x26a  :  192 - 0xc0
    "00000000", --  619 - 0x26b  :    0 - 0x0
    "00000000", --  620 - 0x26c  :    0 - 0x0
    "11100000", --  621 - 0x26d  :  224 - 0xe0
    "00100000", --  622 - 0x26e  :   32 - 0x20
    "00100000", --  623 - 0x26f  :   32 - 0x20
    "11111000", --  624 - 0x270  :  248 - 0xf8 -- Sprite 0x27
    "11111100", --  625 - 0x271  :  252 - 0xfc
    "11111100", --  626 - 0x272  :  252 - 0xfc
    "11111000", --  627 - 0x273  :  248 - 0xf8
    "01111000", --  628 - 0x274  :  120 - 0x78
    "10000000", --  629 - 0x275  :  128 - 0x80
    "11000000", --  630 - 0x276  :  192 - 0xc0
    "11000000", --  631 - 0x277  :  192 - 0xc0
    "01111000", --  632 - 0x278  :  120 - 0x78
    "11111100", --  633 - 0x279  :  252 - 0xfc
    "11111100", --  634 - 0x27a  :  252 - 0xfc
    "11111000", --  635 - 0x27b  :  248 - 0xf8
    "00000000", --  636 - 0x27c  :    0 - 0x0
    "10000000", --  637 - 0x27d  :  128 - 0x80
    "00000000", --  638 - 0x27e  :    0 - 0x0
    "00000000", --  639 - 0x27f  :    0 - 0x0
    "00000000", --  640 - 0x280  :    0 - 0x0 -- Sprite 0x28
    "00000011", --  641 - 0x281  :    3 - 0x3
    "00000111", --  642 - 0x282  :    7 - 0x7
    "00000111", --  643 - 0x283  :    7 - 0x7
    "00001001", --  644 - 0x284  :    9 - 0x9
    "00001001", --  645 - 0x285  :    9 - 0x9
    "00011100", --  646 - 0x286  :   28 - 0x1c
    "00000000", --  647 - 0x287  :    0 - 0x0
    "00000000", --  648 - 0x288  :    0 - 0x0
    "00000011", --  649 - 0x289  :    3 - 0x3
    "00000111", --  650 - 0x28a  :    7 - 0x7
    "00000000", --  651 - 0x28b  :    0 - 0x0
    "00000110", --  652 - 0x28c  :    6 - 0x6
    "00000110", --  653 - 0x28d  :    6 - 0x6
    "00000011", --  654 - 0x28e  :    3 - 0x3
    "01100011", --  655 - 0x28f  :   99 - 0x63
    "00011111", --  656 - 0x290  :   31 - 0x1f -- Sprite 0x29
    "00001111", --  657 - 0x291  :   15 - 0xf
    "00000111", --  658 - 0x292  :    7 - 0x7
    "00110111", --  659 - 0x293  :   55 - 0x37
    "01111111", --  660 - 0x294  :  127 - 0x7f
    "11011111", --  661 - 0x295  :  223 - 0xdf
    "00001111", --  662 - 0x296  :   15 - 0xf
    "00000110", --  663 - 0x297  :    6 - 0x6
    "11100000", --  664 - 0x298  :  224 - 0xe0
    "00100001", --  665 - 0x299  :   33 - 0x21
    "00000001", --  666 - 0x29a  :    1 - 0x1
    "00000111", --  667 - 0x29b  :    7 - 0x7
    "00000111", --  668 - 0x29c  :    7 - 0x7
    "00011111", --  669 - 0x29d  :   31 - 0x1f
    "00001111", --  670 - 0x29e  :   15 - 0xf
    "00000110", --  671 - 0x29f  :    6 - 0x6
    "00000000", --  672 - 0x2a0  :    0 - 0x0 -- Sprite 0x2a
    "11000000", --  673 - 0x2a1  :  192 - 0xc0
    "11111000", --  674 - 0x2a2  :  248 - 0xf8
    "10000000", --  675 - 0x2a3  :  128 - 0x80
    "00100000", --  676 - 0x2a4  :   32 - 0x20
    "10010000", --  677 - 0x2a5  :  144 - 0x90
    "00111100", --  678 - 0x2a6  :   60 - 0x3c
    "00000000", --  679 - 0x2a7  :    0 - 0x0
    "00000000", --  680 - 0x2a8  :    0 - 0x0
    "11000000", --  681 - 0x2a9  :  192 - 0xc0
    "11111000", --  682 - 0x2aa  :  248 - 0xf8
    "01100000", --  683 - 0x2ab  :   96 - 0x60
    "11011100", --  684 - 0x2ac  :  220 - 0xdc
    "01101110", --  685 - 0x2ad  :  110 - 0x6e
    "11000000", --  686 - 0x2ae  :  192 - 0xc0
    "11111011", --  687 - 0x2af  :  251 - 0xfb
    "11100100", --  688 - 0x2b0  :  228 - 0xe4 -- Sprite 0x2b
    "11111110", --  689 - 0x2b1  :  254 - 0xfe
    "01110000", --  690 - 0x2b2  :  112 - 0x70
    "11110001", --  691 - 0x2b3  :  241 - 0xf1
    "11111111", --  692 - 0x2b4  :  255 - 0xff
    "11111111", --  693 - 0x2b5  :  255 - 0xff
    "00000000", --  694 - 0x2b6  :    0 - 0x0
    "00000000", --  695 - 0x2b7  :    0 - 0x0
    "10000011", --  696 - 0x2b8  :  131 - 0x83
    "11000000", --  697 - 0x2b9  :  192 - 0xc0
    "11110000", --  698 - 0x2ba  :  240 - 0xf0
    "11110000", --  699 - 0x2bb  :  240 - 0xf0
    "11111100", --  700 - 0x2bc  :  252 - 0xfc
    "11111100", --  701 - 0x2bd  :  252 - 0xfc
    "00000000", --  702 - 0x2be  :    0 - 0x0
    "00000000", --  703 - 0x2bf  :    0 - 0x0
    "00000111", --  704 - 0x2c0  :    7 - 0x7 -- Sprite 0x2c
    "00001111", --  705 - 0x2c1  :   15 - 0xf
    "00001111", --  706 - 0x2c2  :   15 - 0xf
    "00010010", --  707 - 0x2c3  :   18 - 0x12
    "00010011", --  708 - 0x2c4  :   19 - 0x13
    "00111000", --  709 - 0x2c5  :   56 - 0x38
    "01110000", --  710 - 0x2c6  :  112 - 0x70
    "11111111", --  711 - 0x2c7  :  255 - 0xff
    "00000111", --  712 - 0x2c8  :    7 - 0x7
    "00001111", --  713 - 0x2c9  :   15 - 0xf
    "00000000", --  714 - 0x2ca  :    0 - 0x0
    "00001101", --  715 - 0x2cb  :   13 - 0xd
    "00001100", --  716 - 0x2cc  :   12 - 0xc
    "00000111", --  717 - 0x2cd  :    7 - 0x7
    "00001111", --  718 - 0x2ce  :   15 - 0xf
    "00000010", --  719 - 0x2cf  :    2 - 0x2
    "11011111", --  720 - 0x2d0  :  223 - 0xdf -- Sprite 0x2d
    "00011110", --  721 - 0x2d1  :   30 - 0x1e
    "00011111", --  722 - 0x2d2  :   31 - 0x1f
    "00011111", --  723 - 0x2d3  :   31 - 0x1f
    "00011111", --  724 - 0x2d4  :   31 - 0x1f
    "00001111", --  725 - 0x2d5  :   15 - 0xf
    "00000111", --  726 - 0x2d6  :    7 - 0x7
    "00000001", --  727 - 0x2d7  :    1 - 0x1
    "00000001", --  728 - 0x2d8  :    1 - 0x1
    "11110011", --  729 - 0x2d9  :  243 - 0xf3
    "01011111", --  730 - 0x2da  :   95 - 0x5f
    "00011111", --  731 - 0x2db  :   31 - 0x1f
    "00011111", --  732 - 0x2dc  :   31 - 0x1f
    "01001111", --  733 - 0x2dd  :   79 - 0x4f
    "00110111", --  734 - 0x2de  :   55 - 0x37
    "11000000", --  735 - 0x2df  :  192 - 0xc0
    "10000000", --  736 - 0x2e0  :  128 - 0x80 -- Sprite 0x2e
    "11110000", --  737 - 0x2e1  :  240 - 0xf0
    "00000000", --  738 - 0x2e2  :    0 - 0x0
    "01000000", --  739 - 0x2e3  :   64 - 0x40
    "00100000", --  740 - 0x2e4  :   32 - 0x20
    "01111000", --  741 - 0x2e5  :  120 - 0x78
    "00000000", --  742 - 0x2e6  :    0 - 0x0
    "11111100", --  743 - 0x2e7  :  252 - 0xfc
    "10000000", --  744 - 0x2e8  :  128 - 0x80
    "11110000", --  745 - 0x2e9  :  240 - 0xf0
    "11000000", --  746 - 0x2ea  :  192 - 0xc0
    "10111000", --  747 - 0x2eb  :  184 - 0xb8
    "11011100", --  748 - 0x2ec  :  220 - 0xdc
    "10000000", --  749 - 0x2ed  :  128 - 0x80
    "11110000", --  750 - 0x2ee  :  240 - 0xf0
    "00000000", --  751 - 0x2ef  :    0 - 0x0
    "11110000", --  752 - 0x2f0  :  240 - 0xf0 -- Sprite 0x2f
    "11100000", --  753 - 0x2f1  :  224 - 0xe0
    "11100000", --  754 - 0x2f2  :  224 - 0xe0
    "11110000", --  755 - 0x2f3  :  240 - 0xf0
    "11111010", --  756 - 0x2f4  :  250 - 0xfa
    "11111110", --  757 - 0x2f5  :  254 - 0xfe
    "11111100", --  758 - 0x2f6  :  252 - 0xfc
    "11011000", --  759 - 0x2f7  :  216 - 0xd8
    "10001111", --  760 - 0x2f8  :  143 - 0x8f
    "11100111", --  761 - 0x2f9  :  231 - 0xe7
    "11100000", --  762 - 0x2fa  :  224 - 0xe0
    "11110000", --  763 - 0x2fb  :  240 - 0xf0
    "11001000", --  764 - 0x2fc  :  200 - 0xc8
    "10001000", --  765 - 0x2fd  :  136 - 0x88
    "00010000", --  766 - 0x2fe  :   16 - 0x10
    "00000000", --  767 - 0x2ff  :    0 - 0x0
    "00000000", --  768 - 0x300  :    0 - 0x0 -- Sprite 0x30
    "00000000", --  769 - 0x301  :    0 - 0x0
    "00000111", --  770 - 0x302  :    7 - 0x7
    "00001000", --  771 - 0x303  :    8 - 0x8
    "00010000", --  772 - 0x304  :   16 - 0x10
    "00100000", --  773 - 0x305  :   32 - 0x20
    "01000000", --  774 - 0x306  :   64 - 0x40
    "01000000", --  775 - 0x307  :   64 - 0x40
    "00000000", --  776 - 0x308  :    0 - 0x0
    "00000000", --  777 - 0x309  :    0 - 0x0
    "00000000", --  778 - 0x30a  :    0 - 0x0
    "00000111", --  779 - 0x30b  :    7 - 0x7
    "00001000", --  780 - 0x30c  :    8 - 0x8
    "00010000", --  781 - 0x30d  :   16 - 0x10
    "00100000", --  782 - 0x30e  :   32 - 0x20
    "00100000", --  783 - 0x30f  :   32 - 0x20
    "01000000", --  784 - 0x310  :   64 - 0x40 -- Sprite 0x31
    "01000000", --  785 - 0x311  :   64 - 0x40
    "00100000", --  786 - 0x312  :   32 - 0x20
    "00010000", --  787 - 0x313  :   16 - 0x10
    "00001000", --  788 - 0x314  :    8 - 0x8
    "00000111", --  789 - 0x315  :    7 - 0x7
    "00000000", --  790 - 0x316  :    0 - 0x0
    "00000000", --  791 - 0x317  :    0 - 0x0
    "00100000", --  792 - 0x318  :   32 - 0x20
    "00100000", --  793 - 0x319  :   32 - 0x20
    "00010000", --  794 - 0x31a  :   16 - 0x10
    "00001000", --  795 - 0x31b  :    8 - 0x8
    "00000111", --  796 - 0x31c  :    7 - 0x7
    "00000000", --  797 - 0x31d  :    0 - 0x0
    "00000000", --  798 - 0x31e  :    0 - 0x0
    "00000000", --  799 - 0x31f  :    0 - 0x0
    "00000000", --  800 - 0x320  :    0 - 0x0 -- Sprite 0x32
    "00000000", --  801 - 0x321  :    0 - 0x0
    "11100000", --  802 - 0x322  :  224 - 0xe0
    "00010000", --  803 - 0x323  :   16 - 0x10
    "00001000", --  804 - 0x324  :    8 - 0x8
    "00000100", --  805 - 0x325  :    4 - 0x4
    "00000010", --  806 - 0x326  :    2 - 0x2
    "00000010", --  807 - 0x327  :    2 - 0x2
    "00000000", --  808 - 0x328  :    0 - 0x0
    "00000000", --  809 - 0x329  :    0 - 0x0
    "00000000", --  810 - 0x32a  :    0 - 0x0
    "11100000", --  811 - 0x32b  :  224 - 0xe0
    "00010000", --  812 - 0x32c  :   16 - 0x10
    "00001000", --  813 - 0x32d  :    8 - 0x8
    "00000100", --  814 - 0x32e  :    4 - 0x4
    "00000100", --  815 - 0x32f  :    4 - 0x4
    "00000010", --  816 - 0x330  :    2 - 0x2 -- Sprite 0x33
    "00000010", --  817 - 0x331  :    2 - 0x2
    "00000100", --  818 - 0x332  :    4 - 0x4
    "00001000", --  819 - 0x333  :    8 - 0x8
    "00010000", --  820 - 0x334  :   16 - 0x10
    "11100000", --  821 - 0x335  :  224 - 0xe0
    "00000000", --  822 - 0x336  :    0 - 0x0
    "00000000", --  823 - 0x337  :    0 - 0x0
    "00000100", --  824 - 0x338  :    4 - 0x4
    "00000100", --  825 - 0x339  :    4 - 0x4
    "00001000", --  826 - 0x33a  :    8 - 0x8
    "00010000", --  827 - 0x33b  :   16 - 0x10
    "11100000", --  828 - 0x33c  :  224 - 0xe0
    "00000000", --  829 - 0x33d  :    0 - 0x0
    "00000000", --  830 - 0x33e  :    0 - 0x0
    "00000000", --  831 - 0x33f  :    0 - 0x0
    "00000000", --  832 - 0x340  :    0 - 0x0 -- Sprite 0x34
    "00000000", --  833 - 0x341  :    0 - 0x0
    "00000000", --  834 - 0x342  :    0 - 0x0
    "00000000", --  835 - 0x343  :    0 - 0x0
    "00000011", --  836 - 0x344  :    3 - 0x3
    "00000100", --  837 - 0x345  :    4 - 0x4
    "00001000", --  838 - 0x346  :    8 - 0x8
    "00010000", --  839 - 0x347  :   16 - 0x10
    "00000000", --  840 - 0x348  :    0 - 0x0
    "00000000", --  841 - 0x349  :    0 - 0x0
    "00000000", --  842 - 0x34a  :    0 - 0x0
    "00000000", --  843 - 0x34b  :    0 - 0x0
    "00000000", --  844 - 0x34c  :    0 - 0x0
    "00000011", --  845 - 0x34d  :    3 - 0x3
    "00000100", --  846 - 0x34e  :    4 - 0x4
    "00001000", --  847 - 0x34f  :    8 - 0x8
    "00010000", --  848 - 0x350  :   16 - 0x10 -- Sprite 0x35
    "00001000", --  849 - 0x351  :    8 - 0x8
    "00000100", --  850 - 0x352  :    4 - 0x4
    "00000011", --  851 - 0x353  :    3 - 0x3
    "00000000", --  852 - 0x354  :    0 - 0x0
    "00000000", --  853 - 0x355  :    0 - 0x0
    "00000000", --  854 - 0x356  :    0 - 0x0
    "00000000", --  855 - 0x357  :    0 - 0x0
    "00001000", --  856 - 0x358  :    8 - 0x8
    "00000100", --  857 - 0x359  :    4 - 0x4
    "00000011", --  858 - 0x35a  :    3 - 0x3
    "00000000", --  859 - 0x35b  :    0 - 0x0
    "00000000", --  860 - 0x35c  :    0 - 0x0
    "00000000", --  861 - 0x35d  :    0 - 0x0
    "00000000", --  862 - 0x35e  :    0 - 0x0
    "00000000", --  863 - 0x35f  :    0 - 0x0
    "00000000", --  864 - 0x360  :    0 - 0x0 -- Sprite 0x36
    "00000000", --  865 - 0x361  :    0 - 0x0
    "00000000", --  866 - 0x362  :    0 - 0x0
    "00000000", --  867 - 0x363  :    0 - 0x0
    "11000000", --  868 - 0x364  :  192 - 0xc0
    "00100000", --  869 - 0x365  :   32 - 0x20
    "00010000", --  870 - 0x366  :   16 - 0x10
    "00001000", --  871 - 0x367  :    8 - 0x8
    "00000000", --  872 - 0x368  :    0 - 0x0
    "00000000", --  873 - 0x369  :    0 - 0x0
    "00000000", --  874 - 0x36a  :    0 - 0x0
    "00000000", --  875 - 0x36b  :    0 - 0x0
    "00000000", --  876 - 0x36c  :    0 - 0x0
    "11000000", --  877 - 0x36d  :  192 - 0xc0
    "00100000", --  878 - 0x36e  :   32 - 0x20
    "00010000", --  879 - 0x36f  :   16 - 0x10
    "00001000", --  880 - 0x370  :    8 - 0x8 -- Sprite 0x37
    "00010000", --  881 - 0x371  :   16 - 0x10
    "00100000", --  882 - 0x372  :   32 - 0x20
    "11000000", --  883 - 0x373  :  192 - 0xc0
    "00000000", --  884 - 0x374  :    0 - 0x0
    "00000000", --  885 - 0x375  :    0 - 0x0
    "00000000", --  886 - 0x376  :    0 - 0x0
    "00000000", --  887 - 0x377  :    0 - 0x0
    "00010000", --  888 - 0x378  :   16 - 0x10
    "00100000", --  889 - 0x379  :   32 - 0x20
    "11000000", --  890 - 0x37a  :  192 - 0xc0
    "00000000", --  891 - 0x37b  :    0 - 0x0
    "00000000", --  892 - 0x37c  :    0 - 0x0
    "00000000", --  893 - 0x37d  :    0 - 0x0
    "00000000", --  894 - 0x37e  :    0 - 0x0
    "00000000", --  895 - 0x37f  :    0 - 0x0
    "00000000", --  896 - 0x380  :    0 - 0x0 -- Sprite 0x38
    "00000000", --  897 - 0x381  :    0 - 0x0
    "00000000", --  898 - 0x382  :    0 - 0x0
    "00000000", --  899 - 0x383  :    0 - 0x0
    "00000000", --  900 - 0x384  :    0 - 0x0
    "00000000", --  901 - 0x385  :    0 - 0x0
    "00000000", --  902 - 0x386  :    0 - 0x0
    "00000001", --  903 - 0x387  :    1 - 0x1
    "00000000", --  904 - 0x388  :    0 - 0x0
    "00000000", --  905 - 0x389  :    0 - 0x0
    "00000000", --  906 - 0x38a  :    0 - 0x0
    "00000000", --  907 - 0x38b  :    0 - 0x0
    "00000000", --  908 - 0x38c  :    0 - 0x0
    "00000000", --  909 - 0x38d  :    0 - 0x0
    "00000000", --  910 - 0x38e  :    0 - 0x0
    "00000000", --  911 - 0x38f  :    0 - 0x0
    "00000010", --  912 - 0x390  :    2 - 0x2 -- Sprite 0x39
    "00000001", --  913 - 0x391  :    1 - 0x1
    "00000000", --  914 - 0x392  :    0 - 0x0
    "00000000", --  915 - 0x393  :    0 - 0x0
    "00000000", --  916 - 0x394  :    0 - 0x0
    "00000000", --  917 - 0x395  :    0 - 0x0
    "00000000", --  918 - 0x396  :    0 - 0x0
    "00000000", --  919 - 0x397  :    0 - 0x0
    "00000001", --  920 - 0x398  :    1 - 0x1
    "00000000", --  921 - 0x399  :    0 - 0x0
    "00000000", --  922 - 0x39a  :    0 - 0x0
    "00000000", --  923 - 0x39b  :    0 - 0x0
    "00000000", --  924 - 0x39c  :    0 - 0x0
    "00000000", --  925 - 0x39d  :    0 - 0x0
    "00000000", --  926 - 0x39e  :    0 - 0x0
    "00000000", --  927 - 0x39f  :    0 - 0x0
    "00000000", --  928 - 0x3a0  :    0 - 0x0 -- Sprite 0x3a
    "00000000", --  929 - 0x3a1  :    0 - 0x0
    "00000000", --  930 - 0x3a2  :    0 - 0x0
    "00000000", --  931 - 0x3a3  :    0 - 0x0
    "00000000", --  932 - 0x3a4  :    0 - 0x0
    "00000000", --  933 - 0x3a5  :    0 - 0x0
    "00000000", --  934 - 0x3a6  :    0 - 0x0
    "00000000", --  935 - 0x3a7  :    0 - 0x0
    "00000000", --  936 - 0x3a8  :    0 - 0x0
    "00000000", --  937 - 0x3a9  :    0 - 0x0
    "00000000", --  938 - 0x3aa  :    0 - 0x0
    "00000000", --  939 - 0x3ab  :    0 - 0x0
    "00000000", --  940 - 0x3ac  :    0 - 0x0
    "00000000", --  941 - 0x3ad  :    0 - 0x0
    "00000000", --  942 - 0x3ae  :    0 - 0x0
    "00000000", --  943 - 0x3af  :    0 - 0x0
    "10000000", --  944 - 0x3b0  :  128 - 0x80 -- Sprite 0x3b
    "00000000", --  945 - 0x3b1  :    0 - 0x0
    "00000000", --  946 - 0x3b2  :    0 - 0x0
    "00000000", --  947 - 0x3b3  :    0 - 0x0
    "00000000", --  948 - 0x3b4  :    0 - 0x0
    "00000000", --  949 - 0x3b5  :    0 - 0x0
    "00000000", --  950 - 0x3b6  :    0 - 0x0
    "00000000", --  951 - 0x3b7  :    0 - 0x0
    "00000000", --  952 - 0x3b8  :    0 - 0x0
    "00000000", --  953 - 0x3b9  :    0 - 0x0
    "00000000", --  954 - 0x3ba  :    0 - 0x0
    "00000000", --  955 - 0x3bb  :    0 - 0x0
    "00000000", --  956 - 0x3bc  :    0 - 0x0
    "00000000", --  957 - 0x3bd  :    0 - 0x0
    "00000000", --  958 - 0x3be  :    0 - 0x0
    "00000000", --  959 - 0x3bf  :    0 - 0x0
    "00000000", --  960 - 0x3c0  :    0 - 0x0 -- Sprite 0x3c
    "00000000", --  961 - 0x3c1  :    0 - 0x0
    "00000000", --  962 - 0x3c2  :    0 - 0x0
    "00000001", --  963 - 0x3c3  :    1 - 0x1
    "00100001", --  964 - 0x3c4  :   33 - 0x21
    "00010000", --  965 - 0x3c5  :   16 - 0x10
    "00000000", --  966 - 0x3c6  :    0 - 0x0
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "00000000", --  968 - 0x3c8  :    0 - 0x0
    "00000001", --  969 - 0x3c9  :    1 - 0x1
    "00000001", --  970 - 0x3ca  :    1 - 0x1
    "01000000", --  971 - 0x3cb  :   64 - 0x40
    "00000000", --  972 - 0x3cc  :    0 - 0x0
    "00000000", --  973 - 0x3cd  :    0 - 0x0
    "00000000", --  974 - 0x3ce  :    0 - 0x0
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "01100000", --  976 - 0x3d0  :   96 - 0x60 -- Sprite 0x3d
    "00000000", --  977 - 0x3d1  :    0 - 0x0
    "00000000", --  978 - 0x3d2  :    0 - 0x0
    "00010000", --  979 - 0x3d3  :   16 - 0x10
    "00100001", --  980 - 0x3d4  :   33 - 0x21
    "00000001", --  981 - 0x3d5  :    1 - 0x1
    "00000000", --  982 - 0x3d6  :    0 - 0x0
    "00000000", --  983 - 0x3d7  :    0 - 0x0
    "10000000", --  984 - 0x3d8  :  128 - 0x80
    "00000000", --  985 - 0x3d9  :    0 - 0x0
    "00000000", --  986 - 0x3da  :    0 - 0x0
    "00000000", --  987 - 0x3db  :    0 - 0x0
    "00000000", --  988 - 0x3dc  :    0 - 0x0
    "01000000", --  989 - 0x3dd  :   64 - 0x40
    "00000001", --  990 - 0x3de  :    1 - 0x1
    "00000001", --  991 - 0x3df  :    1 - 0x1
    "00000000", --  992 - 0x3e0  :    0 - 0x0 -- Sprite 0x3e
    "00000000", --  993 - 0x3e1  :    0 - 0x0
    "00000000", --  994 - 0x3e2  :    0 - 0x0
    "00000000", --  995 - 0x3e3  :    0 - 0x0
    "00001000", --  996 - 0x3e4  :    8 - 0x8
    "00010000", --  997 - 0x3e5  :   16 - 0x10
    "00000000", --  998 - 0x3e6  :    0 - 0x0
    "00000000", --  999 - 0x3e7  :    0 - 0x0
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0
    "00000000", -- 1001 - 0x3e9  :    0 - 0x0
    "00000000", -- 1002 - 0x3ea  :    0 - 0x0
    "00000100", -- 1003 - 0x3eb  :    4 - 0x4
    "00000000", -- 1004 - 0x3ec  :    0 - 0x0
    "00000000", -- 1005 - 0x3ed  :    0 - 0x0
    "00000000", -- 1006 - 0x3ee  :    0 - 0x0
    "00000000", -- 1007 - 0x3ef  :    0 - 0x0
    "00001100", -- 1008 - 0x3f0  :   12 - 0xc -- Sprite 0x3f
    "00000000", -- 1009 - 0x3f1  :    0 - 0x0
    "00000000", -- 1010 - 0x3f2  :    0 - 0x0
    "00010000", -- 1011 - 0x3f3  :   16 - 0x10
    "00001000", -- 1012 - 0x3f4  :    8 - 0x8
    "00000000", -- 1013 - 0x3f5  :    0 - 0x0
    "00000000", -- 1014 - 0x3f6  :    0 - 0x0
    "00000000", -- 1015 - 0x3f7  :    0 - 0x0
    "00000010", -- 1016 - 0x3f8  :    2 - 0x2
    "00000000", -- 1017 - 0x3f9  :    0 - 0x0
    "00000000", -- 1018 - 0x3fa  :    0 - 0x0
    "00000000", -- 1019 - 0x3fb  :    0 - 0x0
    "00000000", -- 1020 - 0x3fc  :    0 - 0x0
    "00000100", -- 1021 - 0x3fd  :    4 - 0x4
    "00000000", -- 1022 - 0x3fe  :    0 - 0x0
    "00000000", -- 1023 - 0x3ff  :    0 - 0x0
    "00000100", -- 1024 - 0x400  :    4 - 0x4 -- Sprite 0x40
    "00000010", -- 1025 - 0x401  :    2 - 0x2
    "00000001", -- 1026 - 0x402  :    1 - 0x1
    "00000000", -- 1027 - 0x403  :    0 - 0x0
    "00000000", -- 1028 - 0x404  :    0 - 0x0
    "00000000", -- 1029 - 0x405  :    0 - 0x0
    "00000000", -- 1030 - 0x406  :    0 - 0x0
    "00000000", -- 1031 - 0x407  :    0 - 0x0
    "00001111", -- 1032 - 0x408  :   15 - 0xf
    "00000111", -- 1033 - 0x409  :    7 - 0x7
    "00000011", -- 1034 - 0x40a  :    3 - 0x3
    "00000000", -- 1035 - 0x40b  :    0 - 0x0
    "00000000", -- 1036 - 0x40c  :    0 - 0x0
    "00000001", -- 1037 - 0x40d  :    1 - 0x1
    "00000001", -- 1038 - 0x40e  :    1 - 0x1
    "00000001", -- 1039 - 0x40f  :    1 - 0x1
    "00000000", -- 1040 - 0x410  :    0 - 0x0 -- Sprite 0x41
    "00000000", -- 1041 - 0x411  :    0 - 0x0
    "00000000", -- 1042 - 0x412  :    0 - 0x0
    "00000000", -- 1043 - 0x413  :    0 - 0x0
    "00000000", -- 1044 - 0x414  :    0 - 0x0
    "00000000", -- 1045 - 0x415  :    0 - 0x0
    "00000001", -- 1046 - 0x416  :    1 - 0x1
    "00000011", -- 1047 - 0x417  :    3 - 0x3
    "00000000", -- 1048 - 0x418  :    0 - 0x0
    "00000000", -- 1049 - 0x419  :    0 - 0x0
    "00000000", -- 1050 - 0x41a  :    0 - 0x0
    "00000000", -- 1051 - 0x41b  :    0 - 0x0
    "00000000", -- 1052 - 0x41c  :    0 - 0x0
    "00000000", -- 1053 - 0x41d  :    0 - 0x0
    "00000001", -- 1054 - 0x41e  :    1 - 0x1
    "00000011", -- 1055 - 0x41f  :    3 - 0x3
    "00000111", -- 1056 - 0x420  :    7 - 0x7 -- Sprite 0x42
    "00000111", -- 1057 - 0x421  :    7 - 0x7
    "00000111", -- 1058 - 0x422  :    7 - 0x7
    "00000011", -- 1059 - 0x423  :    3 - 0x3
    "00000001", -- 1060 - 0x424  :    1 - 0x1
    "00000000", -- 1061 - 0x425  :    0 - 0x0
    "00000000", -- 1062 - 0x426  :    0 - 0x0
    "00000000", -- 1063 - 0x427  :    0 - 0x0
    "00000111", -- 1064 - 0x428  :    7 - 0x7
    "00000111", -- 1065 - 0x429  :    7 - 0x7
    "00000111", -- 1066 - 0x42a  :    7 - 0x7
    "00000111", -- 1067 - 0x42b  :    7 - 0x7
    "00000011", -- 1068 - 0x42c  :    3 - 0x3
    "00000001", -- 1069 - 0x42d  :    1 - 0x1
    "00000000", -- 1070 - 0x42e  :    0 - 0x0
    "00000000", -- 1071 - 0x42f  :    0 - 0x0
    "00000000", -- 1072 - 0x430  :    0 - 0x0 -- Sprite 0x43
    "00000000", -- 1073 - 0x431  :    0 - 0x0
    "00000000", -- 1074 - 0x432  :    0 - 0x0
    "00000000", -- 1075 - 0x433  :    0 - 0x0
    "00000000", -- 1076 - 0x434  :    0 - 0x0
    "00000000", -- 1077 - 0x435  :    0 - 0x0
    "00000000", -- 1078 - 0x436  :    0 - 0x0
    "00000000", -- 1079 - 0x437  :    0 - 0x0
    "00000000", -- 1080 - 0x438  :    0 - 0x0
    "00000000", -- 1081 - 0x439  :    0 - 0x0
    "00000000", -- 1082 - 0x43a  :    0 - 0x0
    "00000000", -- 1083 - 0x43b  :    0 - 0x0
    "00000000", -- 1084 - 0x43c  :    0 - 0x0
    "00000000", -- 1085 - 0x43d  :    0 - 0x0
    "00000000", -- 1086 - 0x43e  :    0 - 0x0
    "00000000", -- 1087 - 0x43f  :    0 - 0x0
    "00000000", -- 1088 - 0x440  :    0 - 0x0 -- Sprite 0x44
    "01000010", -- 1089 - 0x441  :   66 - 0x42
    "00111001", -- 1090 - 0x442  :   57 - 0x39
    "11111111", -- 1091 - 0x443  :  255 - 0xff
    "11111111", -- 1092 - 0x444  :  255 - 0xff
    "11111111", -- 1093 - 0x445  :  255 - 0xff
    "11111111", -- 1094 - 0x446  :  255 - 0xff
    "11111111", -- 1095 - 0x447  :  255 - 0xff
    "11111111", -- 1096 - 0x448  :  255 - 0xff
    "11111111", -- 1097 - 0x449  :  255 - 0xff
    "11111111", -- 1098 - 0x44a  :  255 - 0xff
    "11111111", -- 1099 - 0x44b  :  255 - 0xff
    "11111111", -- 1100 - 0x44c  :  255 - 0xff
    "11111111", -- 1101 - 0x44d  :  255 - 0xff
    "11111111", -- 1102 - 0x44e  :  255 - 0xff
    "11111111", -- 1103 - 0x44f  :  255 - 0xff
    "01111111", -- 1104 - 0x450  :  127 - 0x7f -- Sprite 0x45
    "00111111", -- 1105 - 0x451  :   63 - 0x3f
    "00011111", -- 1106 - 0x452  :   31 - 0x1f
    "00001111", -- 1107 - 0x453  :   15 - 0xf
    "00011111", -- 1108 - 0x454  :   31 - 0x1f
    "11111111", -- 1109 - 0x455  :  255 - 0xff
    "11111111", -- 1110 - 0x456  :  255 - 0xff
    "11111111", -- 1111 - 0x457  :  255 - 0xff
    "11111111", -- 1112 - 0x458  :  255 - 0xff
    "01111111", -- 1113 - 0x459  :  127 - 0x7f
    "00111111", -- 1114 - 0x45a  :   63 - 0x3f
    "00011111", -- 1115 - 0x45b  :   31 - 0x1f
    "00011111", -- 1116 - 0x45c  :   31 - 0x1f
    "11111111", -- 1117 - 0x45d  :  255 - 0xff
    "11111111", -- 1118 - 0x45e  :  255 - 0xff
    "11111111", -- 1119 - 0x45f  :  255 - 0xff
    "11111000", -- 1120 - 0x460  :  248 - 0xf8 -- Sprite 0x46
    "11110111", -- 1121 - 0x461  :  247 - 0xf7
    "11101111", -- 1122 - 0x462  :  239 - 0xef
    "11111111", -- 1123 - 0x463  :  255 - 0xff
    "11111111", -- 1124 - 0x464  :  255 - 0xff
    "11111110", -- 1125 - 0x465  :  254 - 0xfe
    "01111110", -- 1126 - 0x466  :  126 - 0x7e
    "00111110", -- 1127 - 0x467  :   62 - 0x3e
    "11111111", -- 1128 - 0x468  :  255 - 0xff
    "11111111", -- 1129 - 0x469  :  255 - 0xff
    "11111111", -- 1130 - 0x46a  :  255 - 0xff
    "11111111", -- 1131 - 0x46b  :  255 - 0xff
    "11111111", -- 1132 - 0x46c  :  255 - 0xff
    "11111111", -- 1133 - 0x46d  :  255 - 0xff
    "11111111", -- 1134 - 0x46e  :  255 - 0xff
    "01111111", -- 1135 - 0x46f  :  127 - 0x7f
    "00000111", -- 1136 - 0x470  :    7 - 0x7 -- Sprite 0x47
    "00000000", -- 1137 - 0x471  :    0 - 0x0
    "00000000", -- 1138 - 0x472  :    0 - 0x0
    "00000000", -- 1139 - 0x473  :    0 - 0x0
    "00000000", -- 1140 - 0x474  :    0 - 0x0
    "00000000", -- 1141 - 0x475  :    0 - 0x0
    "00000000", -- 1142 - 0x476  :    0 - 0x0
    "00000000", -- 1143 - 0x477  :    0 - 0x0
    "00000111", -- 1144 - 0x478  :    7 - 0x7
    "00000011", -- 1145 - 0x479  :    3 - 0x3
    "00000011", -- 1146 - 0x47a  :    3 - 0x3
    "00000001", -- 1147 - 0x47b  :    1 - 0x1
    "00000000", -- 1148 - 0x47c  :    0 - 0x0
    "00000000", -- 1149 - 0x47d  :    0 - 0x0
    "00000000", -- 1150 - 0x47e  :    0 - 0x0
    "00000000", -- 1151 - 0x47f  :    0 - 0x0
    "00000000", -- 1152 - 0x480  :    0 - 0x0 -- Sprite 0x48
    "00000000", -- 1153 - 0x481  :    0 - 0x0
    "00000000", -- 1154 - 0x482  :    0 - 0x0
    "11000000", -- 1155 - 0x483  :  192 - 0xc0
    "11100000", -- 1156 - 0x484  :  224 - 0xe0
    "11110000", -- 1157 - 0x485  :  240 - 0xf0
    "11011011", -- 1158 - 0x486  :  219 - 0xdb
    "11110110", -- 1159 - 0x487  :  246 - 0xf6
    "00000000", -- 1160 - 0x488  :    0 - 0x0
    "10000000", -- 1161 - 0x489  :  128 - 0x80
    "10000000", -- 1162 - 0x48a  :  128 - 0x80
    "11000000", -- 1163 - 0x48b  :  192 - 0xc0
    "11100000", -- 1164 - 0x48c  :  224 - 0xe0
    "11110000", -- 1165 - 0x48d  :  240 - 0xf0
    "11111111", -- 1166 - 0x48e  :  255 - 0xff
    "11111111", -- 1167 - 0x48f  :  255 - 0xff
    "11001011", -- 1168 - 0x490  :  203 - 0xcb -- Sprite 0x49
    "11100000", -- 1169 - 0x491  :  224 - 0xe0
    "11000100", -- 1170 - 0x492  :  196 - 0xc4
    "00000010", -- 1171 - 0x493  :    2 - 0x2
    "11010001", -- 1172 - 0x494  :  209 - 0xd1
    "11100001", -- 1173 - 0x495  :  225 - 0xe1
    "11010001", -- 1174 - 0x496  :  209 - 0xd1
    "10000011", -- 1175 - 0x497  :  131 - 0x83
    "11111111", -- 1176 - 0x498  :  255 - 0xff
    "11111111", -- 1177 - 0x499  :  255 - 0xff
    "11111111", -- 1178 - 0x49a  :  255 - 0xff
    "11111111", -- 1179 - 0x49b  :  255 - 0xff
    "11111111", -- 1180 - 0x49c  :  255 - 0xff
    "11111111", -- 1181 - 0x49d  :  255 - 0xff
    "11111111", -- 1182 - 0x49e  :  255 - 0xff
    "11111111", -- 1183 - 0x49f  :  255 - 0xff
    "00001111", -- 1184 - 0x4a0  :   15 - 0xf -- Sprite 0x4a
    "11111111", -- 1185 - 0x4a1  :  255 - 0xff
    "11100000", -- 1186 - 0x4a2  :  224 - 0xe0
    "10001111", -- 1187 - 0x4a3  :  143 - 0x8f
    "01101110", -- 1188 - 0x4a4  :  110 - 0x6e
    "01000100", -- 1189 - 0x4a5  :   68 - 0x44
    "11101110", -- 1190 - 0x4a6  :  238 - 0xee
    "01100000", -- 1191 - 0x4a7  :   96 - 0x60
    "11111111", -- 1192 - 0x4a8  :  255 - 0xff
    "11111111", -- 1193 - 0x4a9  :  255 - 0xff
    "11111111", -- 1194 - 0x4aa  :  255 - 0xff
    "11110000", -- 1195 - 0x4ab  :  240 - 0xf0
    "10000000", -- 1196 - 0x4ac  :  128 - 0x80
    "00000000", -- 1197 - 0x4ad  :    0 - 0x0
    "00000000", -- 1198 - 0x4ae  :    0 - 0x0
    "10011111", -- 1199 - 0x4af  :  159 - 0x9f
    "10000011", -- 1200 - 0x4b0  :  131 - 0x83 -- Sprite 0x4b
    "11100000", -- 1201 - 0x4b1  :  224 - 0xe0
    "11100100", -- 1202 - 0x4b2  :  228 - 0xe4
    "11000110", -- 1203 - 0x4b3  :  198 - 0xc6
    "01100001", -- 1204 - 0x4b4  :   97 - 0x61
    "00110011", -- 1205 - 0x4b5  :   51 - 0x33
    "00011111", -- 1206 - 0x4b6  :   31 - 0x1f
    "00001111", -- 1207 - 0x4b7  :   15 - 0xf
    "11111111", -- 1208 - 0x4b8  :  255 - 0xff
    "11111111", -- 1209 - 0x4b9  :  255 - 0xff
    "11111001", -- 1210 - 0x4ba  :  249 - 0xf9
    "11111001", -- 1211 - 0x4bb  :  249 - 0xf9
    "01111111", -- 1212 - 0x4bc  :  127 - 0x7f
    "00111111", -- 1213 - 0x4bd  :   63 - 0x3f
    "00011111", -- 1214 - 0x4be  :   31 - 0x1f
    "00001111", -- 1215 - 0x4bf  :   15 - 0xf
    "00000000", -- 1216 - 0x4c0  :    0 - 0x0 -- Sprite 0x4c
    "00000000", -- 1217 - 0x4c1  :    0 - 0x0
    "00000000", -- 1218 - 0x4c2  :    0 - 0x0
    "00000011", -- 1219 - 0x4c3  :    3 - 0x3
    "00000111", -- 1220 - 0x4c4  :    7 - 0x7
    "00001111", -- 1221 - 0x4c5  :   15 - 0xf
    "01011011", -- 1222 - 0x4c6  :   91 - 0x5b
    "10100111", -- 1223 - 0x4c7  :  167 - 0xa7
    "00000000", -- 1224 - 0x4c8  :    0 - 0x0
    "00000001", -- 1225 - 0x4c9  :    1 - 0x1
    "00000001", -- 1226 - 0x4ca  :    1 - 0x1
    "00000011", -- 1227 - 0x4cb  :    3 - 0x3
    "00000111", -- 1228 - 0x4cc  :    7 - 0x7
    "00001111", -- 1229 - 0x4cd  :   15 - 0xf
    "11111111", -- 1230 - 0x4ce  :  255 - 0xff
    "11111111", -- 1231 - 0x4cf  :  255 - 0xff
    "01110011", -- 1232 - 0x4d0  :  115 - 0x73 -- Sprite 0x4d
    "00000111", -- 1233 - 0x4d1  :    7 - 0x7
    "00100111", -- 1234 - 0x4d2  :   39 - 0x27
    "01000000", -- 1235 - 0x4d3  :   64 - 0x40
    "10001011", -- 1236 - 0x4d4  :  139 - 0x8b
    "10000111", -- 1237 - 0x4d5  :  135 - 0x87
    "10001011", -- 1238 - 0x4d6  :  139 - 0x8b
    "11000001", -- 1239 - 0x4d7  :  193 - 0xc1
    "11111111", -- 1240 - 0x4d8  :  255 - 0xff
    "11111111", -- 1241 - 0x4d9  :  255 - 0xff
    "11111111", -- 1242 - 0x4da  :  255 - 0xff
    "11111111", -- 1243 - 0x4db  :  255 - 0xff
    "11111111", -- 1244 - 0x4dc  :  255 - 0xff
    "11111111", -- 1245 - 0x4dd  :  255 - 0xff
    "11111111", -- 1246 - 0x4de  :  255 - 0xff
    "11111111", -- 1247 - 0x4df  :  255 - 0xff
    "11110000", -- 1248 - 0x4e0  :  240 - 0xf0 -- Sprite 0x4e
    "11111111", -- 1249 - 0x4e1  :  255 - 0xff
    "00001111", -- 1250 - 0x4e2  :   15 - 0xf
    "11100001", -- 1251 - 0x4e3  :  225 - 0xe1
    "11101100", -- 1252 - 0x4e4  :  236 - 0xec
    "01000100", -- 1253 - 0x4e5  :   68 - 0x44
    "11101110", -- 1254 - 0x4e6  :  238 - 0xee
    "00001100", -- 1255 - 0x4e7  :   12 - 0xc
    "11111111", -- 1256 - 0x4e8  :  255 - 0xff
    "11111111", -- 1257 - 0x4e9  :  255 - 0xff
    "11111111", -- 1258 - 0x4ea  :  255 - 0xff
    "00011111", -- 1259 - 0x4eb  :   31 - 0x1f
    "00000011", -- 1260 - 0x4ec  :    3 - 0x3
    "00000001", -- 1261 - 0x4ed  :    1 - 0x1
    "00000001", -- 1262 - 0x4ee  :    1 - 0x1
    "11110011", -- 1263 - 0x4ef  :  243 - 0xf3
    "10000000", -- 1264 - 0x4f0  :  128 - 0x80 -- Sprite 0x4f
    "00001110", -- 1265 - 0x4f1  :   14 - 0xe
    "01001110", -- 1266 - 0x4f2  :   78 - 0x4e
    "11000110", -- 1267 - 0x4f3  :  198 - 0xc6
    "00001100", -- 1268 - 0x4f4  :   12 - 0xc
    "10011000", -- 1269 - 0x4f5  :  152 - 0x98
    "11110000", -- 1270 - 0x4f6  :  240 - 0xf0
    "11100000", -- 1271 - 0x4f7  :  224 - 0xe0
    "11111111", -- 1272 - 0x4f8  :  255 - 0xff
    "11111111", -- 1273 - 0x4f9  :  255 - 0xff
    "00111111", -- 1274 - 0x4fa  :   63 - 0x3f
    "00111111", -- 1275 - 0x4fb  :   63 - 0x3f
    "11111100", -- 1276 - 0x4fc  :  252 - 0xfc
    "11111000", -- 1277 - 0x4fd  :  248 - 0xf8
    "11110000", -- 1278 - 0x4fe  :  240 - 0xf0
    "11100000", -- 1279 - 0x4ff  :  224 - 0xe0
    "00000000", -- 1280 - 0x500  :    0 - 0x0 -- Sprite 0x50
    "01000010", -- 1281 - 0x501  :   66 - 0x42
    "10011100", -- 1282 - 0x502  :  156 - 0x9c
    "11111111", -- 1283 - 0x503  :  255 - 0xff
    "11111111", -- 1284 - 0x504  :  255 - 0xff
    "11111111", -- 1285 - 0x505  :  255 - 0xff
    "11111111", -- 1286 - 0x506  :  255 - 0xff
    "11111111", -- 1287 - 0x507  :  255 - 0xff
    "11111111", -- 1288 - 0x508  :  255 - 0xff
    "11111111", -- 1289 - 0x509  :  255 - 0xff
    "11111111", -- 1290 - 0x50a  :  255 - 0xff
    "11111111", -- 1291 - 0x50b  :  255 - 0xff
    "11111111", -- 1292 - 0x50c  :  255 - 0xff
    "11111111", -- 1293 - 0x50d  :  255 - 0xff
    "11111111", -- 1294 - 0x50e  :  255 - 0xff
    "11111111", -- 1295 - 0x50f  :  255 - 0xff
    "11111110", -- 1296 - 0x510  :  254 - 0xfe -- Sprite 0x51
    "11111100", -- 1297 - 0x511  :  252 - 0xfc
    "11111000", -- 1298 - 0x512  :  248 - 0xf8
    "11110000", -- 1299 - 0x513  :  240 - 0xf0
    "11111000", -- 1300 - 0x514  :  248 - 0xf8
    "11111111", -- 1301 - 0x515  :  255 - 0xff
    "11111111", -- 1302 - 0x516  :  255 - 0xff
    "11111111", -- 1303 - 0x517  :  255 - 0xff
    "11111111", -- 1304 - 0x518  :  255 - 0xff
    "11111110", -- 1305 - 0x519  :  254 - 0xfe
    "11111100", -- 1306 - 0x51a  :  252 - 0xfc
    "11111000", -- 1307 - 0x51b  :  248 - 0xf8
    "11111000", -- 1308 - 0x51c  :  248 - 0xf8
    "11111111", -- 1309 - 0x51d  :  255 - 0xff
    "11111111", -- 1310 - 0x51e  :  255 - 0xff
    "11111111", -- 1311 - 0x51f  :  255 - 0xff
    "00011111", -- 1312 - 0x520  :   31 - 0x1f -- Sprite 0x52
    "11101111", -- 1313 - 0x521  :  239 - 0xef
    "11110111", -- 1314 - 0x522  :  247 - 0xf7
    "11111111", -- 1315 - 0x523  :  255 - 0xff
    "11111111", -- 1316 - 0x524  :  255 - 0xff
    "11111110", -- 1317 - 0x525  :  254 - 0xfe
    "01111100", -- 1318 - 0x526  :  124 - 0x7c
    "01110000", -- 1319 - 0x527  :  112 - 0x70
    "11111111", -- 1320 - 0x528  :  255 - 0xff
    "11111111", -- 1321 - 0x529  :  255 - 0xff
    "11111111", -- 1322 - 0x52a  :  255 - 0xff
    "11111111", -- 1323 - 0x52b  :  255 - 0xff
    "11111111", -- 1324 - 0x52c  :  255 - 0xff
    "11111111", -- 1325 - 0x52d  :  255 - 0xff
    "11111110", -- 1326 - 0x52e  :  254 - 0xfe
    "11111100", -- 1327 - 0x52f  :  252 - 0xfc
    "11100000", -- 1328 - 0x530  :  224 - 0xe0 -- Sprite 0x53
    "00000000", -- 1329 - 0x531  :    0 - 0x0
    "00000000", -- 1330 - 0x532  :    0 - 0x0
    "00000000", -- 1331 - 0x533  :    0 - 0x0
    "00000000", -- 1332 - 0x534  :    0 - 0x0
    "00000000", -- 1333 - 0x535  :    0 - 0x0
    "00000000", -- 1334 - 0x536  :    0 - 0x0
    "00000000", -- 1335 - 0x537  :    0 - 0x0
    "11100000", -- 1336 - 0x538  :  224 - 0xe0
    "10000000", -- 1337 - 0x539  :  128 - 0x80
    "10000000", -- 1338 - 0x53a  :  128 - 0x80
    "00000000", -- 1339 - 0x53b  :    0 - 0x0
    "00000000", -- 1340 - 0x53c  :    0 - 0x0
    "00000000", -- 1341 - 0x53d  :    0 - 0x0
    "00000000", -- 1342 - 0x53e  :    0 - 0x0
    "00000000", -- 1343 - 0x53f  :    0 - 0x0
    "00100000", -- 1344 - 0x540  :   32 - 0x20 -- Sprite 0x54
    "01000000", -- 1345 - 0x541  :   64 - 0x40
    "10000000", -- 1346 - 0x542  :  128 - 0x80
    "00000000", -- 1347 - 0x543  :    0 - 0x0
    "00000000", -- 1348 - 0x544  :    0 - 0x0
    "00000000", -- 1349 - 0x545  :    0 - 0x0
    "00000000", -- 1350 - 0x546  :    0 - 0x0
    "00000000", -- 1351 - 0x547  :    0 - 0x0
    "11110000", -- 1352 - 0x548  :  240 - 0xf0
    "11100000", -- 1353 - 0x549  :  224 - 0xe0
    "11000000", -- 1354 - 0x54a  :  192 - 0xc0
    "00000000", -- 1355 - 0x54b  :    0 - 0x0
    "00000000", -- 1356 - 0x54c  :    0 - 0x0
    "10000000", -- 1357 - 0x54d  :  128 - 0x80
    "10000000", -- 1358 - 0x54e  :  128 - 0x80
    "10000000", -- 1359 - 0x54f  :  128 - 0x80
    "00000000", -- 1360 - 0x550  :    0 - 0x0 -- Sprite 0x55
    "00000000", -- 1361 - 0x551  :    0 - 0x0
    "00000000", -- 1362 - 0x552  :    0 - 0x0
    "00000000", -- 1363 - 0x553  :    0 - 0x0
    "00000000", -- 1364 - 0x554  :    0 - 0x0
    "00000000", -- 1365 - 0x555  :    0 - 0x0
    "10000000", -- 1366 - 0x556  :  128 - 0x80
    "11000000", -- 1367 - 0x557  :  192 - 0xc0
    "00000000", -- 1368 - 0x558  :    0 - 0x0
    "00000000", -- 1369 - 0x559  :    0 - 0x0
    "00000000", -- 1370 - 0x55a  :    0 - 0x0
    "00000000", -- 1371 - 0x55b  :    0 - 0x0
    "00000000", -- 1372 - 0x55c  :    0 - 0x0
    "00000000", -- 1373 - 0x55d  :    0 - 0x0
    "10000000", -- 1374 - 0x55e  :  128 - 0x80
    "11000000", -- 1375 - 0x55f  :  192 - 0xc0
    "11100000", -- 1376 - 0x560  :  224 - 0xe0 -- Sprite 0x56
    "11100000", -- 1377 - 0x561  :  224 - 0xe0
    "11100000", -- 1378 - 0x562  :  224 - 0xe0
    "11000000", -- 1379 - 0x563  :  192 - 0xc0
    "10000000", -- 1380 - 0x564  :  128 - 0x80
    "00000000", -- 1381 - 0x565  :    0 - 0x0
    "00000000", -- 1382 - 0x566  :    0 - 0x0
    "00000000", -- 1383 - 0x567  :    0 - 0x0
    "11100000", -- 1384 - 0x568  :  224 - 0xe0
    "11100000", -- 1385 - 0x569  :  224 - 0xe0
    "11100000", -- 1386 - 0x56a  :  224 - 0xe0
    "11100000", -- 1387 - 0x56b  :  224 - 0xe0
    "11000000", -- 1388 - 0x56c  :  192 - 0xc0
    "10000000", -- 1389 - 0x56d  :  128 - 0x80
    "00000000", -- 1390 - 0x56e  :    0 - 0x0
    "00000000", -- 1391 - 0x56f  :    0 - 0x0
    "00000000", -- 1392 - 0x570  :    0 - 0x0 -- Sprite 0x57
    "00000000", -- 1393 - 0x571  :    0 - 0x0
    "00000000", -- 1394 - 0x572  :    0 - 0x0
    "00000000", -- 1395 - 0x573  :    0 - 0x0
    "00000000", -- 1396 - 0x574  :    0 - 0x0
    "00000000", -- 1397 - 0x575  :    0 - 0x0
    "00000000", -- 1398 - 0x576  :    0 - 0x0
    "00000000", -- 1399 - 0x577  :    0 - 0x0
    "00000000", -- 1400 - 0x578  :    0 - 0x0
    "00000000", -- 1401 - 0x579  :    0 - 0x0
    "00000000", -- 1402 - 0x57a  :    0 - 0x0
    "00000000", -- 1403 - 0x57b  :    0 - 0x0
    "00000000", -- 1404 - 0x57c  :    0 - 0x0
    "00000000", -- 1405 - 0x57d  :    0 - 0x0
    "00000000", -- 1406 - 0x57e  :    0 - 0x0
    "00000000", -- 1407 - 0x57f  :    0 - 0x0
    "11111111", -- 1408 - 0x580  :  255 - 0xff -- Sprite 0x58
    "11111111", -- 1409 - 0x581  :  255 - 0xff
    "11111111", -- 1410 - 0x582  :  255 - 0xff
    "11111111", -- 1411 - 0x583  :  255 - 0xff
    "11111111", -- 1412 - 0x584  :  255 - 0xff
    "11111111", -- 1413 - 0x585  :  255 - 0xff
    "11111111", -- 1414 - 0x586  :  255 - 0xff
    "11111111", -- 1415 - 0x587  :  255 - 0xff
    "11111111", -- 1416 - 0x588  :  255 - 0xff
    "11111111", -- 1417 - 0x589  :  255 - 0xff
    "11111111", -- 1418 - 0x58a  :  255 - 0xff
    "11111111", -- 1419 - 0x58b  :  255 - 0xff
    "11111111", -- 1420 - 0x58c  :  255 - 0xff
    "11111111", -- 1421 - 0x58d  :  255 - 0xff
    "11111111", -- 1422 - 0x58e  :  255 - 0xff
    "11111111", -- 1423 - 0x58f  :  255 - 0xff
    "11111111", -- 1424 - 0x590  :  255 - 0xff -- Sprite 0x59
    "11111111", -- 1425 - 0x591  :  255 - 0xff
    "11111111", -- 1426 - 0x592  :  255 - 0xff
    "11111111", -- 1427 - 0x593  :  255 - 0xff
    "11111111", -- 1428 - 0x594  :  255 - 0xff
    "11111111", -- 1429 - 0x595  :  255 - 0xff
    "11111111", -- 1430 - 0x596  :  255 - 0xff
    "11111111", -- 1431 - 0x597  :  255 - 0xff
    "11111111", -- 1432 - 0x598  :  255 - 0xff
    "11111111", -- 1433 - 0x599  :  255 - 0xff
    "11111111", -- 1434 - 0x59a  :  255 - 0xff
    "11111111", -- 1435 - 0x59b  :  255 - 0xff
    "11111111", -- 1436 - 0x59c  :  255 - 0xff
    "11111111", -- 1437 - 0x59d  :  255 - 0xff
    "11111111", -- 1438 - 0x59e  :  255 - 0xff
    "11111111", -- 1439 - 0x59f  :  255 - 0xff
    "11111111", -- 1440 - 0x5a0  :  255 - 0xff -- Sprite 0x5a
    "11111111", -- 1441 - 0x5a1  :  255 - 0xff
    "11111111", -- 1442 - 0x5a2  :  255 - 0xff
    "11111111", -- 1443 - 0x5a3  :  255 - 0xff
    "11111111", -- 1444 - 0x5a4  :  255 - 0xff
    "11111111", -- 1445 - 0x5a5  :  255 - 0xff
    "11111111", -- 1446 - 0x5a6  :  255 - 0xff
    "11111111", -- 1447 - 0x5a7  :  255 - 0xff
    "11111111", -- 1448 - 0x5a8  :  255 - 0xff
    "11111111", -- 1449 - 0x5a9  :  255 - 0xff
    "11111111", -- 1450 - 0x5aa  :  255 - 0xff
    "11111111", -- 1451 - 0x5ab  :  255 - 0xff
    "11111111", -- 1452 - 0x5ac  :  255 - 0xff
    "11111111", -- 1453 - 0x5ad  :  255 - 0xff
    "11111111", -- 1454 - 0x5ae  :  255 - 0xff
    "11111111", -- 1455 - 0x5af  :  255 - 0xff
    "11111111", -- 1456 - 0x5b0  :  255 - 0xff -- Sprite 0x5b
    "11111111", -- 1457 - 0x5b1  :  255 - 0xff
    "11111111", -- 1458 - 0x5b2  :  255 - 0xff
    "11111111", -- 1459 - 0x5b3  :  255 - 0xff
    "11111111", -- 1460 - 0x5b4  :  255 - 0xff
    "11111111", -- 1461 - 0x5b5  :  255 - 0xff
    "11111111", -- 1462 - 0x5b6  :  255 - 0xff
    "11111111", -- 1463 - 0x5b7  :  255 - 0xff
    "11111111", -- 1464 - 0x5b8  :  255 - 0xff
    "11111111", -- 1465 - 0x5b9  :  255 - 0xff
    "11111111", -- 1466 - 0x5ba  :  255 - 0xff
    "11111111", -- 1467 - 0x5bb  :  255 - 0xff
    "11111111", -- 1468 - 0x5bc  :  255 - 0xff
    "11111111", -- 1469 - 0x5bd  :  255 - 0xff
    "11111111", -- 1470 - 0x5be  :  255 - 0xff
    "11111111", -- 1471 - 0x5bf  :  255 - 0xff
    "11111111", -- 1472 - 0x5c0  :  255 - 0xff -- Sprite 0x5c
    "11111111", -- 1473 - 0x5c1  :  255 - 0xff
    "11111111", -- 1474 - 0x5c2  :  255 - 0xff
    "11111111", -- 1475 - 0x5c3  :  255 - 0xff
    "11111111", -- 1476 - 0x5c4  :  255 - 0xff
    "11111111", -- 1477 - 0x5c5  :  255 - 0xff
    "11111111", -- 1478 - 0x5c6  :  255 - 0xff
    "11111111", -- 1479 - 0x5c7  :  255 - 0xff
    "11111111", -- 1480 - 0x5c8  :  255 - 0xff
    "11111111", -- 1481 - 0x5c9  :  255 - 0xff
    "11111111", -- 1482 - 0x5ca  :  255 - 0xff
    "11111111", -- 1483 - 0x5cb  :  255 - 0xff
    "11111111", -- 1484 - 0x5cc  :  255 - 0xff
    "11111111", -- 1485 - 0x5cd  :  255 - 0xff
    "11111111", -- 1486 - 0x5ce  :  255 - 0xff
    "11111111", -- 1487 - 0x5cf  :  255 - 0xff
    "11111111", -- 1488 - 0x5d0  :  255 - 0xff -- Sprite 0x5d
    "11111111", -- 1489 - 0x5d1  :  255 - 0xff
    "11111111", -- 1490 - 0x5d2  :  255 - 0xff
    "11111111", -- 1491 - 0x5d3  :  255 - 0xff
    "11111111", -- 1492 - 0x5d4  :  255 - 0xff
    "11111111", -- 1493 - 0x5d5  :  255 - 0xff
    "11111111", -- 1494 - 0x5d6  :  255 - 0xff
    "11111111", -- 1495 - 0x5d7  :  255 - 0xff
    "11111111", -- 1496 - 0x5d8  :  255 - 0xff
    "11111111", -- 1497 - 0x5d9  :  255 - 0xff
    "11111111", -- 1498 - 0x5da  :  255 - 0xff
    "11111111", -- 1499 - 0x5db  :  255 - 0xff
    "11111111", -- 1500 - 0x5dc  :  255 - 0xff
    "11111111", -- 1501 - 0x5dd  :  255 - 0xff
    "11111111", -- 1502 - 0x5de  :  255 - 0xff
    "11111111", -- 1503 - 0x5df  :  255 - 0xff
    "11111111", -- 1504 - 0x5e0  :  255 - 0xff -- Sprite 0x5e
    "11111111", -- 1505 - 0x5e1  :  255 - 0xff
    "11111111", -- 1506 - 0x5e2  :  255 - 0xff
    "11111111", -- 1507 - 0x5e3  :  255 - 0xff
    "11111111", -- 1508 - 0x5e4  :  255 - 0xff
    "11111111", -- 1509 - 0x5e5  :  255 - 0xff
    "11111111", -- 1510 - 0x5e6  :  255 - 0xff
    "11111111", -- 1511 - 0x5e7  :  255 - 0xff
    "11111111", -- 1512 - 0x5e8  :  255 - 0xff
    "11111111", -- 1513 - 0x5e9  :  255 - 0xff
    "11111111", -- 1514 - 0x5ea  :  255 - 0xff
    "11111111", -- 1515 - 0x5eb  :  255 - 0xff
    "11111111", -- 1516 - 0x5ec  :  255 - 0xff
    "11111111", -- 1517 - 0x5ed  :  255 - 0xff
    "11111111", -- 1518 - 0x5ee  :  255 - 0xff
    "11111111", -- 1519 - 0x5ef  :  255 - 0xff
    "11111111", -- 1520 - 0x5f0  :  255 - 0xff -- Sprite 0x5f
    "11111111", -- 1521 - 0x5f1  :  255 - 0xff
    "11111111", -- 1522 - 0x5f2  :  255 - 0xff
    "11111111", -- 1523 - 0x5f3  :  255 - 0xff
    "11111111", -- 1524 - 0x5f4  :  255 - 0xff
    "11111111", -- 1525 - 0x5f5  :  255 - 0xff
    "11111111", -- 1526 - 0x5f6  :  255 - 0xff
    "11111111", -- 1527 - 0x5f7  :  255 - 0xff
    "11111111", -- 1528 - 0x5f8  :  255 - 0xff
    "11111111", -- 1529 - 0x5f9  :  255 - 0xff
    "11111111", -- 1530 - 0x5fa  :  255 - 0xff
    "11111111", -- 1531 - 0x5fb  :  255 - 0xff
    "11111111", -- 1532 - 0x5fc  :  255 - 0xff
    "11111111", -- 1533 - 0x5fd  :  255 - 0xff
    "11111111", -- 1534 - 0x5fe  :  255 - 0xff
    "11111111", -- 1535 - 0x5ff  :  255 - 0xff
    "00000000", -- 1536 - 0x600  :    0 - 0x0 -- Sprite 0x60
    "00000000", -- 1537 - 0x601  :    0 - 0x0
    "00011111", -- 1538 - 0x602  :   31 - 0x1f
    "00111111", -- 1539 - 0x603  :   63 - 0x3f
    "00111111", -- 1540 - 0x604  :   63 - 0x3f
    "01111111", -- 1541 - 0x605  :  127 - 0x7f
    "01111111", -- 1542 - 0x606  :  127 - 0x7f
    "01111111", -- 1543 - 0x607  :  127 - 0x7f
    "00000000", -- 1544 - 0x608  :    0 - 0x0
    "00001111", -- 1545 - 0x609  :   15 - 0xf
    "00101000", -- 1546 - 0x60a  :   40 - 0x28
    "01011100", -- 1547 - 0x60b  :   92 - 0x5c
    "00111111", -- 1548 - 0x60c  :   63 - 0x3f
    "01111111", -- 1549 - 0x60d  :  127 - 0x7f
    "01111111", -- 1550 - 0x60e  :  127 - 0x7f
    "01111111", -- 1551 - 0x60f  :  127 - 0x7f
    "01111111", -- 1552 - 0x610  :  127 - 0x7f -- Sprite 0x61
    "00111110", -- 1553 - 0x611  :   62 - 0x3e
    "00011111", -- 1554 - 0x612  :   31 - 0x1f
    "00011111", -- 1555 - 0x613  :   31 - 0x1f
    "00001111", -- 1556 - 0x614  :   15 - 0xf
    "00001111", -- 1557 - 0x615  :   15 - 0xf
    "00001111", -- 1558 - 0x616  :   15 - 0xf
    "00000111", -- 1559 - 0x617  :    7 - 0x7
    "01111111", -- 1560 - 0x618  :  127 - 0x7f
    "00111110", -- 1561 - 0x619  :   62 - 0x3e
    "00011111", -- 1562 - 0x61a  :   31 - 0x1f
    "00011111", -- 1563 - 0x61b  :   31 - 0x1f
    "00001000", -- 1564 - 0x61c  :    8 - 0x8
    "00000000", -- 1565 - 0x61d  :    0 - 0x0
    "00000000", -- 1566 - 0x61e  :    0 - 0x0
    "00000000", -- 1567 - 0x61f  :    0 - 0x0
    "00000000", -- 1568 - 0x620  :    0 - 0x0 -- Sprite 0x62
    "01100000", -- 1569 - 0x621  :   96 - 0x60
    "11110000", -- 1570 - 0x622  :  240 - 0xf0
    "11111000", -- 1571 - 0x623  :  248 - 0xf8
    "11111000", -- 1572 - 0x624  :  248 - 0xf8
    "11111000", -- 1573 - 0x625  :  248 - 0xf8
    "11111100", -- 1574 - 0x626  :  252 - 0xfc
    "11111100", -- 1575 - 0x627  :  252 - 0xfc
    "00000000", -- 1576 - 0x628  :    0 - 0x0
    "10000000", -- 1577 - 0x629  :  128 - 0x80
    "01000000", -- 1578 - 0x62a  :   64 - 0x40
    "11000100", -- 1579 - 0x62b  :  196 - 0xc4
    "11110110", -- 1580 - 0x62c  :  246 - 0xf6
    "11111110", -- 1581 - 0x62d  :  254 - 0xfe
    "11111100", -- 1582 - 0x62e  :  252 - 0xfc
    "11111100", -- 1583 - 0x62f  :  252 - 0xfc
    "11111000", -- 1584 - 0x630  :  248 - 0xf8 -- Sprite 0x63
    "11110000", -- 1585 - 0x631  :  240 - 0xf0
    "11110000", -- 1586 - 0x632  :  240 - 0xf0
    "11100000", -- 1587 - 0x633  :  224 - 0xe0
    "10000000", -- 1588 - 0x634  :  128 - 0x80
    "10000000", -- 1589 - 0x635  :  128 - 0x80
    "11000000", -- 1590 - 0x636  :  192 - 0xc0
    "11000000", -- 1591 - 0x637  :  192 - 0xc0
    "11111000", -- 1592 - 0x638  :  248 - 0xf8
    "11110000", -- 1593 - 0x639  :  240 - 0xf0
    "00000000", -- 1594 - 0x63a  :    0 - 0x0
    "00000000", -- 1595 - 0x63b  :    0 - 0x0
    "10000000", -- 1596 - 0x63c  :  128 - 0x80
    "00000000", -- 1597 - 0x63d  :    0 - 0x0
    "00000000", -- 1598 - 0x63e  :    0 - 0x0
    "00000000", -- 1599 - 0x63f  :    0 - 0x0
    "00000000", -- 1600 - 0x640  :    0 - 0x0 -- Sprite 0x64
    "00011111", -- 1601 - 0x641  :   31 - 0x1f
    "00111111", -- 1602 - 0x642  :   63 - 0x3f
    "01111111", -- 1603 - 0x643  :  127 - 0x7f
    "11111111", -- 1604 - 0x644  :  255 - 0xff
    "11111111", -- 1605 - 0x645  :  255 - 0xff
    "00111110", -- 1606 - 0x646  :   62 - 0x3e
    "00001111", -- 1607 - 0x647  :   15 - 0xf
    "00000000", -- 1608 - 0x648  :    0 - 0x0
    "00011100", -- 1609 - 0x649  :   28 - 0x1c
    "00111111", -- 1610 - 0x64a  :   63 - 0x3f
    "01111111", -- 1611 - 0x64b  :  127 - 0x7f
    "11111111", -- 1612 - 0x64c  :  255 - 0xff
    "11111111", -- 1613 - 0x64d  :  255 - 0xff
    "00111110", -- 1614 - 0x64e  :   62 - 0x3e
    "01110000", -- 1615 - 0x64f  :  112 - 0x70
    "00000000", -- 1616 - 0x650  :    0 - 0x0 -- Sprite 0x65
    "00000000", -- 1617 - 0x651  :    0 - 0x0
    "00000000", -- 1618 - 0x652  :    0 - 0x0
    "00000001", -- 1619 - 0x653  :    1 - 0x1
    "00000000", -- 1620 - 0x654  :    0 - 0x0
    "00000000", -- 1621 - 0x655  :    0 - 0x0
    "00000000", -- 1622 - 0x656  :    0 - 0x0
    "00000000", -- 1623 - 0x657  :    0 - 0x0
    "00000000", -- 1624 - 0x658  :    0 - 0x0
    "00000000", -- 1625 - 0x659  :    0 - 0x0
    "00000000", -- 1626 - 0x65a  :    0 - 0x0
    "00000000", -- 1627 - 0x65b  :    0 - 0x0
    "00000000", -- 1628 - 0x65c  :    0 - 0x0
    "00000000", -- 1629 - 0x65d  :    0 - 0x0
    "00000000", -- 1630 - 0x65e  :    0 - 0x0
    "00000000", -- 1631 - 0x65f  :    0 - 0x0
    "00000000", -- 1632 - 0x660  :    0 - 0x0 -- Sprite 0x66
    "11100000", -- 1633 - 0x661  :  224 - 0xe0
    "11110000", -- 1634 - 0x662  :  240 - 0xf0
    "11111100", -- 1635 - 0x663  :  252 - 0xfc
    "11111110", -- 1636 - 0x664  :  254 - 0xfe
    "11111110", -- 1637 - 0x665  :  254 - 0xfe
    "11111111", -- 1638 - 0x666  :  255 - 0xff
    "11111100", -- 1639 - 0x667  :  252 - 0xfc
    "00000000", -- 1640 - 0x668  :    0 - 0x0
    "01100000", -- 1641 - 0x669  :   96 - 0x60
    "11110000", -- 1642 - 0x66a  :  240 - 0xf0
    "11111000", -- 1643 - 0x66b  :  248 - 0xf8
    "11111100", -- 1644 - 0x66c  :  252 - 0xfc
    "11111100", -- 1645 - 0x66d  :  252 - 0xfc
    "11111100", -- 1646 - 0x66e  :  252 - 0xfc
    "11111111", -- 1647 - 0x66f  :  255 - 0xff
    "01111100", -- 1648 - 0x670  :  124 - 0x7c -- Sprite 0x67
    "11111100", -- 1649 - 0x671  :  252 - 0xfc
    "11111000", -- 1650 - 0x672  :  248 - 0xf8
    "11110000", -- 1651 - 0x673  :  240 - 0xf0
    "11100000", -- 1652 - 0x674  :  224 - 0xe0
    "00000000", -- 1653 - 0x675  :    0 - 0x0
    "00000000", -- 1654 - 0x676  :    0 - 0x0
    "00000000", -- 1655 - 0x677  :    0 - 0x0
    "01111100", -- 1656 - 0x678  :  124 - 0x7c
    "11111100", -- 1657 - 0x679  :  252 - 0xfc
    "10001000", -- 1658 - 0x67a  :  136 - 0x88
    "00000000", -- 1659 - 0x67b  :    0 - 0x0
    "00000000", -- 1660 - 0x67c  :    0 - 0x0
    "00000000", -- 1661 - 0x67d  :    0 - 0x0
    "00000000", -- 1662 - 0x67e  :    0 - 0x0
    "00000000", -- 1663 - 0x67f  :    0 - 0x0
    "00000000", -- 1664 - 0x680  :    0 - 0x0 -- Sprite 0x68
    "00000111", -- 1665 - 0x681  :    7 - 0x7
    "00000111", -- 1666 - 0x682  :    7 - 0x7
    "00001111", -- 1667 - 0x683  :   15 - 0xf
    "00001111", -- 1668 - 0x684  :   15 - 0xf
    "00000000", -- 1669 - 0x685  :    0 - 0x0
    "00011111", -- 1670 - 0x686  :   31 - 0x1f
    "00111111", -- 1671 - 0x687  :   63 - 0x3f
    "00000000", -- 1672 - 0x688  :    0 - 0x0
    "00000111", -- 1673 - 0x689  :    7 - 0x7
    "00000011", -- 1674 - 0x68a  :    3 - 0x3
    "00000000", -- 1675 - 0x68b  :    0 - 0x0
    "00000000", -- 1676 - 0x68c  :    0 - 0x0
    "00000111", -- 1677 - 0x68d  :    7 - 0x7
    "00000100", -- 1678 - 0x68e  :    4 - 0x4
    "00000100", -- 1679 - 0x68f  :    4 - 0x4
    "01111111", -- 1680 - 0x690  :  127 - 0x7f -- Sprite 0x69
    "01111111", -- 1681 - 0x691  :  127 - 0x7f
    "00011111", -- 1682 - 0x692  :   31 - 0x1f
    "00011111", -- 1683 - 0x693  :   31 - 0x1f
    "00011111", -- 1684 - 0x694  :   31 - 0x1f
    "00011110", -- 1685 - 0x695  :   30 - 0x1e
    "00001111", -- 1686 - 0x696  :   15 - 0xf
    "00011111", -- 1687 - 0x697  :   31 - 0x1f
    "00001100", -- 1688 - 0x698  :   12 - 0xc
    "10011110", -- 1689 - 0x699  :  158 - 0x9e
    "11111111", -- 1690 - 0x69a  :  255 - 0xff
    "00011111", -- 1691 - 0x69b  :   31 - 0x1f
    "00011111", -- 1692 - 0x69c  :   31 - 0x1f
    "00011110", -- 1693 - 0x69d  :   30 - 0x1e
    "00001111", -- 1694 - 0x69e  :   15 - 0xf
    "00000000", -- 1695 - 0x69f  :    0 - 0x0
    "00000000", -- 1696 - 0x6a0  :    0 - 0x0 -- Sprite 0x6a
    "11100000", -- 1697 - 0x6a1  :  224 - 0xe0
    "11100000", -- 1698 - 0x6a2  :  224 - 0xe0
    "11110000", -- 1699 - 0x6a3  :  240 - 0xf0
    "11110000", -- 1700 - 0x6a4  :  240 - 0xf0
    "00000000", -- 1701 - 0x6a5  :    0 - 0x0
    "11111000", -- 1702 - 0x6a6  :  248 - 0xf8
    "11111100", -- 1703 - 0x6a7  :  252 - 0xfc
    "00000000", -- 1704 - 0x6a8  :    0 - 0x0
    "11100000", -- 1705 - 0x6a9  :  224 - 0xe0
    "11000000", -- 1706 - 0x6aa  :  192 - 0xc0
    "00000000", -- 1707 - 0x6ab  :    0 - 0x0
    "00000000", -- 1708 - 0x6ac  :    0 - 0x0
    "11100000", -- 1709 - 0x6ad  :  224 - 0xe0
    "00100000", -- 1710 - 0x6ae  :   32 - 0x20
    "00100000", -- 1711 - 0x6af  :   32 - 0x20
    "11111110", -- 1712 - 0x6b0  :  254 - 0xfe -- Sprite 0x6b
    "11111110", -- 1713 - 0x6b1  :  254 - 0xfe
    "11111000", -- 1714 - 0x6b2  :  248 - 0xf8
    "11111000", -- 1715 - 0x6b3  :  248 - 0xf8
    "11111000", -- 1716 - 0x6b4  :  248 - 0xf8
    "01111000", -- 1717 - 0x6b5  :  120 - 0x78
    "11110000", -- 1718 - 0x6b6  :  240 - 0xf0
    "11111000", -- 1719 - 0x6b7  :  248 - 0xf8
    "00110000", -- 1720 - 0x6b8  :   48 - 0x30
    "01111001", -- 1721 - 0x6b9  :  121 - 0x79
    "11111111", -- 1722 - 0x6ba  :  255 - 0xff
    "11111000", -- 1723 - 0x6bb  :  248 - 0xf8
    "11111000", -- 1724 - 0x6bc  :  248 - 0xf8
    "01111000", -- 1725 - 0x6bd  :  120 - 0x78
    "11110000", -- 1726 - 0x6be  :  240 - 0xf0
    "00000000", -- 1727 - 0x6bf  :    0 - 0x0
    "00000011", -- 1728 - 0x6c0  :    3 - 0x3 -- Sprite 0x6c
    "00000111", -- 1729 - 0x6c1  :    7 - 0x7
    "00000101", -- 1730 - 0x6c2  :    5 - 0x5
    "00001000", -- 1731 - 0x6c3  :    8 - 0x8
    "00011011", -- 1732 - 0x6c4  :   27 - 0x1b
    "00011001", -- 1733 - 0x6c5  :   25 - 0x19
    "00000101", -- 1734 - 0x6c6  :    5 - 0x5
    "00111111", -- 1735 - 0x6c7  :   63 - 0x3f
    "00000011", -- 1736 - 0x6c8  :    3 - 0x3
    "00000111", -- 1737 - 0x6c9  :    7 - 0x7
    "00000010", -- 1738 - 0x6ca  :    2 - 0x2
    "00000111", -- 1739 - 0x6cb  :    7 - 0x7
    "00000100", -- 1740 - 0x6cc  :    4 - 0x4
    "01000110", -- 1741 - 0x6cd  :   70 - 0x46
    "11100011", -- 1742 - 0x6ce  :  227 - 0xe3
    "11000010", -- 1743 - 0x6cf  :  194 - 0xc2
    "00111111", -- 1744 - 0x6d0  :   63 - 0x3f -- Sprite 0x6d
    "00001111", -- 1745 - 0x6d1  :   15 - 0xf
    "00000101", -- 1746 - 0x6d2  :    5 - 0x5
    "00110111", -- 1747 - 0x6d3  :   55 - 0x37
    "00111111", -- 1748 - 0x6d4  :   63 - 0x3f
    "00111111", -- 1749 - 0x6d5  :   63 - 0x3f
    "00111110", -- 1750 - 0x6d6  :   62 - 0x3e
    "00011100", -- 1751 - 0x6d7  :   28 - 0x1c
    "01000010", -- 1752 - 0x6d8  :   66 - 0x42
    "00000111", -- 1753 - 0x6d9  :    7 - 0x7
    "00000111", -- 1754 - 0x6da  :    7 - 0x7
    "00000111", -- 1755 - 0x6db  :    7 - 0x7
    "00000111", -- 1756 - 0x6dc  :    7 - 0x7
    "00000011", -- 1757 - 0x6dd  :    3 - 0x3
    "00000010", -- 1758 - 0x6de  :    2 - 0x2
    "00000000", -- 1759 - 0x6df  :    0 - 0x0
    "11100000", -- 1760 - 0x6e0  :  224 - 0xe0 -- Sprite 0x6e
    "11110000", -- 1761 - 0x6e1  :  240 - 0xf0
    "01010000", -- 1762 - 0x6e2  :   80 - 0x50
    "00001000", -- 1763 - 0x6e3  :    8 - 0x8
    "01101100", -- 1764 - 0x6e4  :  108 - 0x6c
    "11001100", -- 1765 - 0x6e5  :  204 - 0xcc
    "11010000", -- 1766 - 0x6e6  :  208 - 0xd0
    "11111110", -- 1767 - 0x6e7  :  254 - 0xfe
    "11100000", -- 1768 - 0x6e8  :  224 - 0xe0
    "11110000", -- 1769 - 0x6e9  :  240 - 0xf0
    "10100000", -- 1770 - 0x6ea  :  160 - 0xa0
    "11110000", -- 1771 - 0x6eb  :  240 - 0xf0
    "10010000", -- 1772 - 0x6ec  :  144 - 0x90
    "00110010", -- 1773 - 0x6ed  :   50 - 0x32
    "11100011", -- 1774 - 0x6ee  :  227 - 0xe3
    "00100001", -- 1775 - 0x6ef  :   33 - 0x21
    "11111110", -- 1776 - 0x6f0  :  254 - 0xfe -- Sprite 0x6f
    "11111000", -- 1777 - 0x6f1  :  248 - 0xf8
    "11010000", -- 1778 - 0x6f2  :  208 - 0xd0
    "11111011", -- 1779 - 0x6f3  :  251 - 0xfb
    "11111111", -- 1780 - 0x6f4  :  255 - 0xff
    "11111111", -- 1781 - 0x6f5  :  255 - 0xff
    "00111110", -- 1782 - 0x6f6  :   62 - 0x3e
    "00001100", -- 1783 - 0x6f7  :   12 - 0xc
    "00100000", -- 1784 - 0x6f8  :   32 - 0x20
    "01110000", -- 1785 - 0x6f9  :  112 - 0x70
    "11110000", -- 1786 - 0x6fa  :  240 - 0xf0
    "11111000", -- 1787 - 0x6fb  :  248 - 0xf8
    "11111000", -- 1788 - 0x6fc  :  248 - 0xf8
    "11110000", -- 1789 - 0x6fd  :  240 - 0xf0
    "00110000", -- 1790 - 0x6fe  :   48 - 0x30
    "00000000", -- 1791 - 0x6ff  :    0 - 0x0
    "00000000", -- 1792 - 0x700  :    0 - 0x0 -- Sprite 0x70
    "00000000", -- 1793 - 0x701  :    0 - 0x0
    "01111001", -- 1794 - 0x702  :  121 - 0x79
    "11111001", -- 1795 - 0x703  :  249 - 0xf9
    "11110011", -- 1796 - 0x704  :  243 - 0xf3
    "11111111", -- 1797 - 0x705  :  255 - 0xff
    "01111011", -- 1798 - 0x706  :  123 - 0x7b
    "00111111", -- 1799 - 0x707  :   63 - 0x3f
    "00000000", -- 1800 - 0x708  :    0 - 0x0
    "00000001", -- 1801 - 0x709  :    1 - 0x1
    "00000000", -- 1802 - 0x70a  :    0 - 0x0
    "00000000", -- 1803 - 0x70b  :    0 - 0x0
    "00000000", -- 1804 - 0x70c  :    0 - 0x0
    "00011110", -- 1805 - 0x70d  :   30 - 0x1e
    "01111111", -- 1806 - 0x70e  :  127 - 0x7f
    "00111110", -- 1807 - 0x70f  :   62 - 0x3e
    "00111111", -- 1808 - 0x710  :   63 - 0x3f -- Sprite 0x71
    "00111111", -- 1809 - 0x711  :   63 - 0x3f
    "01111011", -- 1810 - 0x712  :  123 - 0x7b
    "01111111", -- 1811 - 0x713  :  127 - 0x7f
    "11111011", -- 1812 - 0x714  :  251 - 0xfb
    "11110001", -- 1813 - 0x715  :  241 - 0xf1
    "01111001", -- 1814 - 0x716  :  121 - 0x79
    "00111000", -- 1815 - 0x717  :   56 - 0x38
    "00111100", -- 1816 - 0x718  :   60 - 0x3c
    "00111110", -- 1817 - 0x719  :   62 - 0x3e
    "01111111", -- 1818 - 0x71a  :  127 - 0x7f
    "01111110", -- 1819 - 0x71b  :  126 - 0x7e
    "00011000", -- 1820 - 0x71c  :   24 - 0x18
    "00000000", -- 1821 - 0x71d  :    0 - 0x0
    "00000000", -- 1822 - 0x71e  :    0 - 0x0
    "00000000", -- 1823 - 0x71f  :    0 - 0x0
    "00000000", -- 1824 - 0x720  :    0 - 0x0 -- Sprite 0x72
    "00000000", -- 1825 - 0x721  :    0 - 0x0
    "10000000", -- 1826 - 0x722  :  128 - 0x80
    "10110000", -- 1827 - 0x723  :  176 - 0xb0
    "10111000", -- 1828 - 0x724  :  184 - 0xb8
    "11000110", -- 1829 - 0x725  :  198 - 0xc6
    "10010011", -- 1830 - 0x726  :  147 - 0x93
    "11110111", -- 1831 - 0x727  :  247 - 0xf7
    "11000000", -- 1832 - 0x728  :  192 - 0xc0
    "11100000", -- 1833 - 0x729  :  224 - 0xe0
    "01000000", -- 1834 - 0x72a  :   64 - 0x40
    "00000000", -- 1835 - 0x72b  :    0 - 0x0
    "00000000", -- 1836 - 0x72c  :    0 - 0x0
    "00111010", -- 1837 - 0x72d  :   58 - 0x3a
    "11101111", -- 1838 - 0x72e  :  239 - 0xef
    "01001011", -- 1839 - 0x72f  :   75 - 0x4b
    "11100011", -- 1840 - 0x730  :  227 - 0xe3 -- Sprite 0x73
    "11110111", -- 1841 - 0x731  :  247 - 0xf7
    "10010011", -- 1842 - 0x732  :  147 - 0x93
    "11000110", -- 1843 - 0x733  :  198 - 0xc6
    "10111000", -- 1844 - 0x734  :  184 - 0xb8
    "10110000", -- 1845 - 0x735  :  176 - 0xb0
    "10000000", -- 1846 - 0x736  :  128 - 0x80
    "00000000", -- 1847 - 0x737  :    0 - 0x0
    "01011111", -- 1848 - 0x738  :   95 - 0x5f
    "01001011", -- 1849 - 0x739  :   75 - 0x4b
    "11101111", -- 1850 - 0x73a  :  239 - 0xef
    "00111010", -- 1851 - 0x73b  :   58 - 0x3a
    "00000000", -- 1852 - 0x73c  :    0 - 0x0
    "00000000", -- 1853 - 0x73d  :    0 - 0x0
    "01100000", -- 1854 - 0x73e  :   96 - 0x60
    "11000000", -- 1855 - 0x73f  :  192 - 0xc0
    "00110000", -- 1856 - 0x740  :   48 - 0x30 -- Sprite 0x74
    "01111100", -- 1857 - 0x741  :  124 - 0x7c
    "11111111", -- 1858 - 0x742  :  255 - 0xff
    "11111111", -- 1859 - 0x743  :  255 - 0xff
    "11011111", -- 1860 - 0x744  :  223 - 0xdf
    "00001011", -- 1861 - 0x745  :   11 - 0xb
    "00011111", -- 1862 - 0x746  :   31 - 0x1f
    "01111111", -- 1863 - 0x747  :  127 - 0x7f
    "00000000", -- 1864 - 0x748  :    0 - 0x0
    "00001100", -- 1865 - 0x749  :   12 - 0xc
    "00001111", -- 1866 - 0x74a  :   15 - 0xf
    "00011111", -- 1867 - 0x74b  :   31 - 0x1f
    "00011111", -- 1868 - 0x74c  :   31 - 0x1f
    "00001111", -- 1869 - 0x74d  :   15 - 0xf
    "00001110", -- 1870 - 0x74e  :   14 - 0xe
    "00000100", -- 1871 - 0x74f  :    4 - 0x4
    "01111111", -- 1872 - 0x750  :  127 - 0x7f -- Sprite 0x75
    "00001011", -- 1873 - 0x751  :   11 - 0xb
    "00110011", -- 1874 - 0x752  :   51 - 0x33
    "00110110", -- 1875 - 0x753  :   54 - 0x36
    "00010000", -- 1876 - 0x754  :   16 - 0x10
    "00001010", -- 1877 - 0x755  :   10 - 0xa
    "00001111", -- 1878 - 0x756  :   15 - 0xf
    "00000111", -- 1879 - 0x757  :    7 - 0x7
    "10000100", -- 1880 - 0x758  :  132 - 0x84
    "11000111", -- 1881 - 0x759  :  199 - 0xc7
    "01001100", -- 1882 - 0x75a  :   76 - 0x4c
    "00001001", -- 1883 - 0x75b  :    9 - 0x9
    "00001111", -- 1884 - 0x75c  :   15 - 0xf
    "00000101", -- 1885 - 0x75d  :    5 - 0x5
    "00001111", -- 1886 - 0x75e  :   15 - 0xf
    "00000111", -- 1887 - 0x75f  :    7 - 0x7
    "00111000", -- 1888 - 0x760  :   56 - 0x38 -- Sprite 0x76
    "01111100", -- 1889 - 0x761  :  124 - 0x7c
    "11111100", -- 1890 - 0x762  :  252 - 0xfc
    "11111100", -- 1891 - 0x763  :  252 - 0xfc
    "11101100", -- 1892 - 0x764  :  236 - 0xec
    "10100000", -- 1893 - 0x765  :  160 - 0xa0
    "11110000", -- 1894 - 0x766  :  240 - 0xf0
    "11111100", -- 1895 - 0x767  :  252 - 0xfc
    "00000000", -- 1896 - 0x768  :    0 - 0x0
    "01000000", -- 1897 - 0x769  :   64 - 0x40
    "11000000", -- 1898 - 0x76a  :  192 - 0xc0
    "11100000", -- 1899 - 0x76b  :  224 - 0xe0
    "11100000", -- 1900 - 0x76c  :  224 - 0xe0
    "11100000", -- 1901 - 0x76d  :  224 - 0xe0
    "11100000", -- 1902 - 0x76e  :  224 - 0xe0
    "01000010", -- 1903 - 0x76f  :   66 - 0x42
    "11111100", -- 1904 - 0x770  :  252 - 0xfc -- Sprite 0x77
    "10100000", -- 1905 - 0x771  :  160 - 0xa0
    "10011000", -- 1906 - 0x772  :  152 - 0x98
    "11011000", -- 1907 - 0x773  :  216 - 0xd8
    "00010000", -- 1908 - 0x774  :   16 - 0x10
    "10100000", -- 1909 - 0x775  :  160 - 0xa0
    "11100000", -- 1910 - 0x776  :  224 - 0xe0
    "11000000", -- 1911 - 0x777  :  192 - 0xc0
    "01000011", -- 1912 - 0x778  :   67 - 0x43
    "11000111", -- 1913 - 0x779  :  199 - 0xc7
    "01100010", -- 1914 - 0x77a  :   98 - 0x62
    "00100000", -- 1915 - 0x77b  :   32 - 0x20
    "11100000", -- 1916 - 0x77c  :  224 - 0xe0
    "01000000", -- 1917 - 0x77d  :   64 - 0x40
    "11100000", -- 1918 - 0x77e  :  224 - 0xe0
    "11000000", -- 1919 - 0x77f  :  192 - 0xc0
    "00000000", -- 1920 - 0x780  :    0 - 0x0 -- Sprite 0x78
    "00000001", -- 1921 - 0x781  :    1 - 0x1
    "00001101", -- 1922 - 0x782  :   13 - 0xd
    "00011101", -- 1923 - 0x783  :   29 - 0x1d
    "01100011", -- 1924 - 0x784  :   99 - 0x63
    "11001001", -- 1925 - 0x785  :  201 - 0xc9
    "11101111", -- 1926 - 0x786  :  239 - 0xef
    "11000111", -- 1927 - 0x787  :  199 - 0xc7
    "00000011", -- 1928 - 0x788  :    3 - 0x3
    "00000100", -- 1929 - 0x789  :    4 - 0x4
    "00000000", -- 1930 - 0x78a  :    0 - 0x0
    "00000000", -- 1931 - 0x78b  :    0 - 0x0
    "01011100", -- 1932 - 0x78c  :   92 - 0x5c
    "11110111", -- 1933 - 0x78d  :  247 - 0xf7
    "11010010", -- 1934 - 0x78e  :  210 - 0xd2
    "11111010", -- 1935 - 0x78f  :  250 - 0xfa
    "11101111", -- 1936 - 0x790  :  239 - 0xef -- Sprite 0x79
    "11001001", -- 1937 - 0x791  :  201 - 0xc9
    "01100011", -- 1938 - 0x792  :   99 - 0x63
    "00011101", -- 1939 - 0x793  :   29 - 0x1d
    "00001101", -- 1940 - 0x794  :   13 - 0xd
    "00000001", -- 1941 - 0x795  :    1 - 0x1
    "00000000", -- 1942 - 0x796  :    0 - 0x0
    "00000000", -- 1943 - 0x797  :    0 - 0x0
    "11010010", -- 1944 - 0x798  :  210 - 0xd2
    "11110111", -- 1945 - 0x799  :  247 - 0xf7
    "01011100", -- 1946 - 0x79a  :   92 - 0x5c
    "00000000", -- 1947 - 0x79b  :    0 - 0x0
    "00000000", -- 1948 - 0x79c  :    0 - 0x0
    "00000010", -- 1949 - 0x79d  :    2 - 0x2
    "00000111", -- 1950 - 0x79e  :    7 - 0x7
    "00000011", -- 1951 - 0x79f  :    3 - 0x3
    "00011100", -- 1952 - 0x7a0  :   28 - 0x1c -- Sprite 0x7a
    "10011110", -- 1953 - 0x7a1  :  158 - 0x9e
    "10001111", -- 1954 - 0x7a2  :  143 - 0x8f
    "11011111", -- 1955 - 0x7a3  :  223 - 0xdf
    "11111110", -- 1956 - 0x7a4  :  254 - 0xfe
    "11011110", -- 1957 - 0x7a5  :  222 - 0xde
    "11111100", -- 1958 - 0x7a6  :  252 - 0xfc
    "11111100", -- 1959 - 0x7a7  :  252 - 0xfc
    "00000000", -- 1960 - 0x7a8  :    0 - 0x0
    "00000000", -- 1961 - 0x7a9  :    0 - 0x0
    "00000000", -- 1962 - 0x7aa  :    0 - 0x0
    "00011000", -- 1963 - 0x7ab  :   24 - 0x18
    "01111110", -- 1964 - 0x7ac  :  126 - 0x7e
    "11111110", -- 1965 - 0x7ad  :  254 - 0xfe
    "01111100", -- 1966 - 0x7ae  :  124 - 0x7c
    "00111100", -- 1967 - 0x7af  :   60 - 0x3c
    "11111100", -- 1968 - 0x7b0  :  252 - 0xfc -- Sprite 0x7b
    "11011110", -- 1969 - 0x7b1  :  222 - 0xde
    "11111111", -- 1970 - 0x7b2  :  255 - 0xff
    "11001111", -- 1971 - 0x7b3  :  207 - 0xcf
    "10011111", -- 1972 - 0x7b4  :  159 - 0x9f
    "10011110", -- 1973 - 0x7b5  :  158 - 0x9e
    "00000000", -- 1974 - 0x7b6  :    0 - 0x0
    "00000000", -- 1975 - 0x7b7  :    0 - 0x0
    "01111100", -- 1976 - 0x7b8  :  124 - 0x7c
    "11111110", -- 1977 - 0x7b9  :  254 - 0xfe
    "01111000", -- 1978 - 0x7ba  :  120 - 0x78
    "00000000", -- 1979 - 0x7bb  :    0 - 0x0
    "00000000", -- 1980 - 0x7bc  :    0 - 0x0
    "00000000", -- 1981 - 0x7bd  :    0 - 0x0
    "10000000", -- 1982 - 0x7be  :  128 - 0x80
    "00000000", -- 1983 - 0x7bf  :    0 - 0x0
    "00000000", -- 1984 - 0x7c0  :    0 - 0x0 -- Sprite 0x7c
    "00000000", -- 1985 - 0x7c1  :    0 - 0x0
    "00000000", -- 1986 - 0x7c2  :    0 - 0x0
    "00000000", -- 1987 - 0x7c3  :    0 - 0x0
    "00011110", -- 1988 - 0x7c4  :   30 - 0x1e
    "00111111", -- 1989 - 0x7c5  :   63 - 0x3f
    "01111101", -- 1990 - 0x7c6  :  125 - 0x7d
    "01111000", -- 1991 - 0x7c7  :  120 - 0x78
    "00000000", -- 1992 - 0x7c8  :    0 - 0x0
    "00000000", -- 1993 - 0x7c9  :    0 - 0x0
    "00000001", -- 1994 - 0x7ca  :    1 - 0x1
    "00000000", -- 1995 - 0x7cb  :    0 - 0x0
    "00000000", -- 1996 - 0x7cc  :    0 - 0x0
    "00100000", -- 1997 - 0x7cd  :   32 - 0x20
    "01111100", -- 1998 - 0x7ce  :  124 - 0x7c
    "01111000", -- 1999 - 0x7cf  :  120 - 0x78
    "01111100", -- 2000 - 0x7d0  :  124 - 0x7c -- Sprite 0x7d
    "11111011", -- 2001 - 0x7d1  :  251 - 0xfb
    "11111111", -- 2002 - 0x7d2  :  255 - 0xff
    "11111111", -- 2003 - 0x7d3  :  255 - 0xff
    "01011111", -- 2004 - 0x7d4  :   95 - 0x5f
    "00011111", -- 2005 - 0x7d5  :   31 - 0x1f
    "00011111", -- 2006 - 0x7d6  :   31 - 0x1f
    "00011111", -- 2007 - 0x7d7  :   31 - 0x1f
    "01111100", -- 2008 - 0x7d8  :  124 - 0x7c
    "11111110", -- 2009 - 0x7d9  :  254 - 0xfe
    "11111111", -- 2010 - 0x7da  :  255 - 0xff
    "11111110", -- 2011 - 0x7db  :  254 - 0xfe
    "01111100", -- 2012 - 0x7dc  :  124 - 0x7c
    "01100000", -- 2013 - 0x7dd  :   96 - 0x60
    "11100000", -- 2014 - 0x7de  :  224 - 0xe0
    "11100001", -- 2015 - 0x7df  :  225 - 0xe1
    "00000000", -- 2016 - 0x7e0  :    0 - 0x0 -- Sprite 0x7e
    "00000000", -- 2017 - 0x7e1  :    0 - 0x0
    "00000000", -- 2018 - 0x7e2  :    0 - 0x0
    "00000000", -- 2019 - 0x7e3  :    0 - 0x0
    "00000000", -- 2020 - 0x7e4  :    0 - 0x0
    "10000000", -- 2021 - 0x7e5  :  128 - 0x80
    "10000000", -- 2022 - 0x7e6  :  128 - 0x80
    "00000000", -- 2023 - 0x7e7  :    0 - 0x0
    "01111100", -- 2024 - 0x7e8  :  124 - 0x7c
    "10000010", -- 2025 - 0x7e9  :  130 - 0x82
    "00000001", -- 2026 - 0x7ea  :    1 - 0x1
    "10000010", -- 2027 - 0x7eb  :  130 - 0x82
    "01111100", -- 2028 - 0x7ec  :  124 - 0x7c
    "00000000", -- 2029 - 0x7ed  :    0 - 0x0
    "00000000", -- 2030 - 0x7ee  :    0 - 0x0
    "00000000", -- 2031 - 0x7ef  :    0 - 0x0
    "00000000", -- 2032 - 0x7f0  :    0 - 0x0 -- Sprite 0x7f
    "00100001", -- 2033 - 0x7f1  :   33 - 0x21
    "10100010", -- 2034 - 0x7f2  :  162 - 0xa2
    "10100011", -- 2035 - 0x7f3  :  163 - 0xa3
    "10110011", -- 2036 - 0x7f4  :  179 - 0xb3
    "10001111", -- 2037 - 0x7f5  :  143 - 0x8f
    "00100111", -- 2038 - 0x7f6  :   39 - 0x27
    "11111110", -- 2039 - 0x7f7  :  254 - 0xfe
    "00010000", -- 2040 - 0x7f8  :   16 - 0x10
    "00011001", -- 2041 - 0x7f9  :   25 - 0x19
    "01011010", -- 2042 - 0x7fa  :   90 - 0x5a
    "11011111", -- 2043 - 0x7fb  :  223 - 0xdf
    "01001111", -- 2044 - 0x7fc  :   79 - 0x4f
    "01110011", -- 2045 - 0x7fd  :  115 - 0x73
    "11011011", -- 2046 - 0x7fe  :  219 - 0xdb
    "00000010", -- 2047 - 0x7ff  :    2 - 0x2
    "00000000", -- 2048 - 0x800  :    0 - 0x0 -- Sprite 0x80
    "00000000", -- 2049 - 0x801  :    0 - 0x0
    "00000000", -- 2050 - 0x802  :    0 - 0x0
    "00000000", -- 2051 - 0x803  :    0 - 0x0
    "00000011", -- 2052 - 0x804  :    3 - 0x3
    "00001111", -- 2053 - 0x805  :   15 - 0xf
    "00011111", -- 2054 - 0x806  :   31 - 0x1f
    "00011111", -- 2055 - 0x807  :   31 - 0x1f
    "00000000", -- 2056 - 0x808  :    0 - 0x0
    "00000000", -- 2057 - 0x809  :    0 - 0x0
    "00000000", -- 2058 - 0x80a  :    0 - 0x0
    "00000011", -- 2059 - 0x80b  :    3 - 0x3
    "00001100", -- 2060 - 0x80c  :   12 - 0xc
    "00010000", -- 2061 - 0x80d  :   16 - 0x10
    "00100010", -- 2062 - 0x80e  :   34 - 0x22
    "00100000", -- 2063 - 0x80f  :   32 - 0x20
    "00011111", -- 2064 - 0x810  :   31 - 0x1f -- Sprite 0x81
    "00011111", -- 2065 - 0x811  :   31 - 0x1f
    "00001111", -- 2066 - 0x812  :   15 - 0xf
    "00000011", -- 2067 - 0x813  :    3 - 0x3
    "00000000", -- 2068 - 0x814  :    0 - 0x0
    "00000000", -- 2069 - 0x815  :    0 - 0x0
    "00000000", -- 2070 - 0x816  :    0 - 0x0
    "00000000", -- 2071 - 0x817  :    0 - 0x0
    "00100001", -- 2072 - 0x818  :   33 - 0x21
    "00100011", -- 2073 - 0x819  :   35 - 0x23
    "00010000", -- 2074 - 0x81a  :   16 - 0x10
    "00001100", -- 2075 - 0x81b  :   12 - 0xc
    "00000011", -- 2076 - 0x81c  :    3 - 0x3
    "00000000", -- 2077 - 0x81d  :    0 - 0x0
    "00000000", -- 2078 - 0x81e  :    0 - 0x0
    "00000000", -- 2079 - 0x81f  :    0 - 0x0
    "00000000", -- 2080 - 0x820  :    0 - 0x0 -- Sprite 0x82
    "00000000", -- 2081 - 0x821  :    0 - 0x0
    "00000000", -- 2082 - 0x822  :    0 - 0x0
    "00000000", -- 2083 - 0x823  :    0 - 0x0
    "11000000", -- 2084 - 0x824  :  192 - 0xc0
    "11110000", -- 2085 - 0x825  :  240 - 0xf0
    "11111000", -- 2086 - 0x826  :  248 - 0xf8
    "11111000", -- 2087 - 0x827  :  248 - 0xf8
    "00000000", -- 2088 - 0x828  :    0 - 0x0
    "00000000", -- 2089 - 0x829  :    0 - 0x0
    "00000000", -- 2090 - 0x82a  :    0 - 0x0
    "11000000", -- 2091 - 0x82b  :  192 - 0xc0
    "00110000", -- 2092 - 0x82c  :   48 - 0x30
    "00001000", -- 2093 - 0x82d  :    8 - 0x8
    "01100100", -- 2094 - 0x82e  :  100 - 0x64
    "11000100", -- 2095 - 0x82f  :  196 - 0xc4
    "11111000", -- 2096 - 0x830  :  248 - 0xf8 -- Sprite 0x83
    "11111000", -- 2097 - 0x831  :  248 - 0xf8
    "11110000", -- 2098 - 0x832  :  240 - 0xf0
    "11000000", -- 2099 - 0x833  :  192 - 0xc0
    "00000000", -- 2100 - 0x834  :    0 - 0x0
    "00000000", -- 2101 - 0x835  :    0 - 0x0
    "00000000", -- 2102 - 0x836  :    0 - 0x0
    "00000000", -- 2103 - 0x837  :    0 - 0x0
    "10000100", -- 2104 - 0x838  :  132 - 0x84
    "00000100", -- 2105 - 0x839  :    4 - 0x4
    "00001000", -- 2106 - 0x83a  :    8 - 0x8
    "00110000", -- 2107 - 0x83b  :   48 - 0x30
    "11000000", -- 2108 - 0x83c  :  192 - 0xc0
    "00000000", -- 2109 - 0x83d  :    0 - 0x0
    "00000000", -- 2110 - 0x83e  :    0 - 0x0
    "00000000", -- 2111 - 0x83f  :    0 - 0x0
    "00000000", -- 2112 - 0x840  :    0 - 0x0 -- Sprite 0x84
    "00000000", -- 2113 - 0x841  :    0 - 0x0
    "00000000", -- 2114 - 0x842  :    0 - 0x0
    "00000000", -- 2115 - 0x843  :    0 - 0x0
    "00000011", -- 2116 - 0x844  :    3 - 0x3
    "00001111", -- 2117 - 0x845  :   15 - 0xf
    "00011111", -- 2118 - 0x846  :   31 - 0x1f
    "00011111", -- 2119 - 0x847  :   31 - 0x1f
    "00000000", -- 2120 - 0x848  :    0 - 0x0
    "00000000", -- 2121 - 0x849  :    0 - 0x0
    "00000000", -- 2122 - 0x84a  :    0 - 0x0
    "00000011", -- 2123 - 0x84b  :    3 - 0x3
    "00001100", -- 2124 - 0x84c  :   12 - 0xc
    "00010000", -- 2125 - 0x84d  :   16 - 0x10
    "00100110", -- 2126 - 0x84e  :   38 - 0x26
    "00100011", -- 2127 - 0x84f  :   35 - 0x23
    "00011111", -- 2128 - 0x850  :   31 - 0x1f -- Sprite 0x85
    "00011111", -- 2129 - 0x851  :   31 - 0x1f
    "00001111", -- 2130 - 0x852  :   15 - 0xf
    "00000011", -- 2131 - 0x853  :    3 - 0x3
    "00000000", -- 2132 - 0x854  :    0 - 0x0
    "00000000", -- 2133 - 0x855  :    0 - 0x0
    "00000000", -- 2134 - 0x856  :    0 - 0x0
    "00000000", -- 2135 - 0x857  :    0 - 0x0
    "00100001", -- 2136 - 0x858  :   33 - 0x21
    "00100000", -- 2137 - 0x859  :   32 - 0x20
    "00010000", -- 2138 - 0x85a  :   16 - 0x10
    "00001100", -- 2139 - 0x85b  :   12 - 0xc
    "00000011", -- 2140 - 0x85c  :    3 - 0x3
    "00000000", -- 2141 - 0x85d  :    0 - 0x0
    "00000000", -- 2142 - 0x85e  :    0 - 0x0
    "00000000", -- 2143 - 0x85f  :    0 - 0x0
    "00000000", -- 2144 - 0x860  :    0 - 0x0 -- Sprite 0x86
    "00000000", -- 2145 - 0x861  :    0 - 0x0
    "00000000", -- 2146 - 0x862  :    0 - 0x0
    "00000000", -- 2147 - 0x863  :    0 - 0x0
    "11000000", -- 2148 - 0x864  :  192 - 0xc0
    "11110000", -- 2149 - 0x865  :  240 - 0xf0
    "11111000", -- 2150 - 0x866  :  248 - 0xf8
    "11111000", -- 2151 - 0x867  :  248 - 0xf8
    "00000000", -- 2152 - 0x868  :    0 - 0x0
    "00000000", -- 2153 - 0x869  :    0 - 0x0
    "00000000", -- 2154 - 0x86a  :    0 - 0x0
    "11000000", -- 2155 - 0x86b  :  192 - 0xc0
    "00110000", -- 2156 - 0x86c  :   48 - 0x30
    "00001000", -- 2157 - 0x86d  :    8 - 0x8
    "01000100", -- 2158 - 0x86e  :   68 - 0x44
    "00000100", -- 2159 - 0x86f  :    4 - 0x4
    "11111000", -- 2160 - 0x870  :  248 - 0xf8 -- Sprite 0x87
    "11111000", -- 2161 - 0x871  :  248 - 0xf8
    "11110000", -- 2162 - 0x872  :  240 - 0xf0
    "11000000", -- 2163 - 0x873  :  192 - 0xc0
    "00000000", -- 2164 - 0x874  :    0 - 0x0
    "00000000", -- 2165 - 0x875  :    0 - 0x0
    "00000000", -- 2166 - 0x876  :    0 - 0x0
    "00000000", -- 2167 - 0x877  :    0 - 0x0
    "10000100", -- 2168 - 0x878  :  132 - 0x84
    "11000100", -- 2169 - 0x879  :  196 - 0xc4
    "00001000", -- 2170 - 0x87a  :    8 - 0x8
    "00110000", -- 2171 - 0x87b  :   48 - 0x30
    "11000000", -- 2172 - 0x87c  :  192 - 0xc0
    "00000000", -- 2173 - 0x87d  :    0 - 0x0
    "00000000", -- 2174 - 0x87e  :    0 - 0x0
    "00000000", -- 2175 - 0x87f  :    0 - 0x0
    "00000000", -- 2176 - 0x880  :    0 - 0x0 -- Sprite 0x88
    "00000000", -- 2177 - 0x881  :    0 - 0x0
    "00000000", -- 2178 - 0x882  :    0 - 0x0
    "00000000", -- 2179 - 0x883  :    0 - 0x0
    "00000011", -- 2180 - 0x884  :    3 - 0x3
    "00001111", -- 2181 - 0x885  :   15 - 0xf
    "00011111", -- 2182 - 0x886  :   31 - 0x1f
    "00011111", -- 2183 - 0x887  :   31 - 0x1f
    "00000000", -- 2184 - 0x888  :    0 - 0x0
    "00000000", -- 2185 - 0x889  :    0 - 0x0
    "00000000", -- 2186 - 0x88a  :    0 - 0x0
    "00000011", -- 2187 - 0x88b  :    3 - 0x3
    "00001100", -- 2188 - 0x88c  :   12 - 0xc
    "00010000", -- 2189 - 0x88d  :   16 - 0x10
    "00100000", -- 2190 - 0x88e  :   32 - 0x20
    "00100001", -- 2191 - 0x88f  :   33 - 0x21
    "00011111", -- 2192 - 0x890  :   31 - 0x1f -- Sprite 0x89
    "00011111", -- 2193 - 0x891  :   31 - 0x1f
    "00001111", -- 2194 - 0x892  :   15 - 0xf
    "00000011", -- 2195 - 0x893  :    3 - 0x3
    "00000000", -- 2196 - 0x894  :    0 - 0x0
    "00000000", -- 2197 - 0x895  :    0 - 0x0
    "00000000", -- 2198 - 0x896  :    0 - 0x0
    "00000000", -- 2199 - 0x897  :    0 - 0x0
    "00100011", -- 2200 - 0x898  :   35 - 0x23
    "00100110", -- 2201 - 0x899  :   38 - 0x26
    "00010000", -- 2202 - 0x89a  :   16 - 0x10
    "00001100", -- 2203 - 0x89b  :   12 - 0xc
    "00000011", -- 2204 - 0x89c  :    3 - 0x3
    "00000000", -- 2205 - 0x89d  :    0 - 0x0
    "00000000", -- 2206 - 0x89e  :    0 - 0x0
    "00000000", -- 2207 - 0x89f  :    0 - 0x0
    "00000000", -- 2208 - 0x8a0  :    0 - 0x0 -- Sprite 0x8a
    "00000000", -- 2209 - 0x8a1  :    0 - 0x0
    "00000000", -- 2210 - 0x8a2  :    0 - 0x0
    "00000000", -- 2211 - 0x8a3  :    0 - 0x0
    "11000000", -- 2212 - 0x8a4  :  192 - 0xc0
    "11110000", -- 2213 - 0x8a5  :  240 - 0xf0
    "11111000", -- 2214 - 0x8a6  :  248 - 0xf8
    "11111000", -- 2215 - 0x8a7  :  248 - 0xf8
    "00000000", -- 2216 - 0x8a8  :    0 - 0x0
    "00000000", -- 2217 - 0x8a9  :    0 - 0x0
    "00000000", -- 2218 - 0x8aa  :    0 - 0x0
    "11000000", -- 2219 - 0x8ab  :  192 - 0xc0
    "00110000", -- 2220 - 0x8ac  :   48 - 0x30
    "00001000", -- 2221 - 0x8ad  :    8 - 0x8
    "11000100", -- 2222 - 0x8ae  :  196 - 0xc4
    "10000100", -- 2223 - 0x8af  :  132 - 0x84
    "11111000", -- 2224 - 0x8b0  :  248 - 0xf8 -- Sprite 0x8b
    "11111000", -- 2225 - 0x8b1  :  248 - 0xf8
    "11110000", -- 2226 - 0x8b2  :  240 - 0xf0
    "11000000", -- 2227 - 0x8b3  :  192 - 0xc0
    "00000000", -- 2228 - 0x8b4  :    0 - 0x0
    "00000000", -- 2229 - 0x8b5  :    0 - 0x0
    "00000000", -- 2230 - 0x8b6  :    0 - 0x0
    "00000000", -- 2231 - 0x8b7  :    0 - 0x0
    "00000100", -- 2232 - 0x8b8  :    4 - 0x4
    "01000100", -- 2233 - 0x8b9  :   68 - 0x44
    "00001000", -- 2234 - 0x8ba  :    8 - 0x8
    "00110000", -- 2235 - 0x8bb  :   48 - 0x30
    "11000000", -- 2236 - 0x8bc  :  192 - 0xc0
    "00000000", -- 2237 - 0x8bd  :    0 - 0x0
    "00000000", -- 2238 - 0x8be  :    0 - 0x0
    "00000000", -- 2239 - 0x8bf  :    0 - 0x0
    "00000000", -- 2240 - 0x8c0  :    0 - 0x0 -- Sprite 0x8c
    "00000000", -- 2241 - 0x8c1  :    0 - 0x0
    "00000000", -- 2242 - 0x8c2  :    0 - 0x0
    "00000000", -- 2243 - 0x8c3  :    0 - 0x0
    "00000011", -- 2244 - 0x8c4  :    3 - 0x3
    "00001111", -- 2245 - 0x8c5  :   15 - 0xf
    "00011111", -- 2246 - 0x8c6  :   31 - 0x1f
    "00011111", -- 2247 - 0x8c7  :   31 - 0x1f
    "00000000", -- 2248 - 0x8c8  :    0 - 0x0
    "00000000", -- 2249 - 0x8c9  :    0 - 0x0
    "00000000", -- 2250 - 0x8ca  :    0 - 0x0
    "00000011", -- 2251 - 0x8cb  :    3 - 0x3
    "00001100", -- 2252 - 0x8cc  :   12 - 0xc
    "00010000", -- 2253 - 0x8cd  :   16 - 0x10
    "00100011", -- 2254 - 0x8ce  :   35 - 0x23
    "00100001", -- 2255 - 0x8cf  :   33 - 0x21
    "00011111", -- 2256 - 0x8d0  :   31 - 0x1f -- Sprite 0x8d
    "00011111", -- 2257 - 0x8d1  :   31 - 0x1f
    "00001111", -- 2258 - 0x8d2  :   15 - 0xf
    "00000011", -- 2259 - 0x8d3  :    3 - 0x3
    "00000000", -- 2260 - 0x8d4  :    0 - 0x0
    "00000000", -- 2261 - 0x8d5  :    0 - 0x0
    "00000000", -- 2262 - 0x8d6  :    0 - 0x0
    "00000000", -- 2263 - 0x8d7  :    0 - 0x0
    "00100000", -- 2264 - 0x8d8  :   32 - 0x20
    "00100010", -- 2265 - 0x8d9  :   34 - 0x22
    "00010000", -- 2266 - 0x8da  :   16 - 0x10
    "00001100", -- 2267 - 0x8db  :   12 - 0xc
    "00000011", -- 2268 - 0x8dc  :    3 - 0x3
    "00000000", -- 2269 - 0x8dd  :    0 - 0x0
    "00000000", -- 2270 - 0x8de  :    0 - 0x0
    "00000000", -- 2271 - 0x8df  :    0 - 0x0
    "00000000", -- 2272 - 0x8e0  :    0 - 0x0 -- Sprite 0x8e
    "00000000", -- 2273 - 0x8e1  :    0 - 0x0
    "00000000", -- 2274 - 0x8e2  :    0 - 0x0
    "00000000", -- 2275 - 0x8e3  :    0 - 0x0
    "11000000", -- 2276 - 0x8e4  :  192 - 0xc0
    "11110000", -- 2277 - 0x8e5  :  240 - 0xf0
    "11111000", -- 2278 - 0x8e6  :  248 - 0xf8
    "11111000", -- 2279 - 0x8e7  :  248 - 0xf8
    "00000000", -- 2280 - 0x8e8  :    0 - 0x0
    "00000000", -- 2281 - 0x8e9  :    0 - 0x0
    "00000000", -- 2282 - 0x8ea  :    0 - 0x0
    "11000000", -- 2283 - 0x8eb  :  192 - 0xc0
    "00110000", -- 2284 - 0x8ec  :   48 - 0x30
    "00001000", -- 2285 - 0x8ed  :    8 - 0x8
    "00000100", -- 2286 - 0x8ee  :    4 - 0x4
    "10000100", -- 2287 - 0x8ef  :  132 - 0x84
    "11111000", -- 2288 - 0x8f0  :  248 - 0xf8 -- Sprite 0x8f
    "11111000", -- 2289 - 0x8f1  :  248 - 0xf8
    "11110000", -- 2290 - 0x8f2  :  240 - 0xf0
    "11000000", -- 2291 - 0x8f3  :  192 - 0xc0
    "00000000", -- 2292 - 0x8f4  :    0 - 0x0
    "00000000", -- 2293 - 0x8f5  :    0 - 0x0
    "00000000", -- 2294 - 0x8f6  :    0 - 0x0
    "00000000", -- 2295 - 0x8f7  :    0 - 0x0
    "11000100", -- 2296 - 0x8f8  :  196 - 0xc4
    "01100100", -- 2297 - 0x8f9  :  100 - 0x64
    "00001000", -- 2298 - 0x8fa  :    8 - 0x8
    "00110000", -- 2299 - 0x8fb  :   48 - 0x30
    "11000000", -- 2300 - 0x8fc  :  192 - 0xc0
    "00000000", -- 2301 - 0x8fd  :    0 - 0x0
    "00000000", -- 2302 - 0x8fe  :    0 - 0x0
    "00000000", -- 2303 - 0x8ff  :    0 - 0x0
    "00000000", -- 2304 - 0x900  :    0 - 0x0 -- Sprite 0x90
    "00000000", -- 2305 - 0x901  :    0 - 0x0
    "00000000", -- 2306 - 0x902  :    0 - 0x0
    "00001111", -- 2307 - 0x903  :   15 - 0xf
    "00110000", -- 2308 - 0x904  :   48 - 0x30
    "01100000", -- 2309 - 0x905  :   96 - 0x60
    "00111111", -- 2310 - 0x906  :   63 - 0x3f
    "01111111", -- 2311 - 0x907  :  127 - 0x7f
    "00000000", -- 2312 - 0x908  :    0 - 0x0
    "00000000", -- 2313 - 0x909  :    0 - 0x0
    "00000000", -- 2314 - 0x90a  :    0 - 0x0
    "00000000", -- 2315 - 0x90b  :    0 - 0x0
    "00101111", -- 2316 - 0x90c  :   47 - 0x2f
    "00111111", -- 2317 - 0x90d  :   63 - 0x3f
    "01100000", -- 2318 - 0x90e  :   96 - 0x60
    "00100000", -- 2319 - 0x90f  :   32 - 0x20
    "01111111", -- 2320 - 0x910  :  127 - 0x7f -- Sprite 0x91
    "00111111", -- 2321 - 0x911  :   63 - 0x3f
    "01100000", -- 2322 - 0x912  :   96 - 0x60
    "00110000", -- 2323 - 0x913  :   48 - 0x30
    "00001111", -- 2324 - 0x914  :   15 - 0xf
    "00000000", -- 2325 - 0x915  :    0 - 0x0
    "00000000", -- 2326 - 0x916  :    0 - 0x0
    "00000000", -- 2327 - 0x917  :    0 - 0x0
    "00100000", -- 2328 - 0x918  :   32 - 0x20
    "01100000", -- 2329 - 0x919  :   96 - 0x60
    "00111111", -- 2330 - 0x91a  :   63 - 0x3f
    "00101111", -- 2331 - 0x91b  :   47 - 0x2f
    "00000000", -- 2332 - 0x91c  :    0 - 0x0
    "00000000", -- 2333 - 0x91d  :    0 - 0x0
    "00000000", -- 2334 - 0x91e  :    0 - 0x0
    "00000000", -- 2335 - 0x91f  :    0 - 0x0
    "00000000", -- 2336 - 0x920  :    0 - 0x0 -- Sprite 0x92
    "00000000", -- 2337 - 0x921  :    0 - 0x0
    "00000000", -- 2338 - 0x922  :    0 - 0x0
    "11111000", -- 2339 - 0x923  :  248 - 0xf8
    "00000110", -- 2340 - 0x924  :    6 - 0x6
    "00000011", -- 2341 - 0x925  :    3 - 0x3
    "11111110", -- 2342 - 0x926  :  254 - 0xfe
    "11111111", -- 2343 - 0x927  :  255 - 0xff
    "00000000", -- 2344 - 0x928  :    0 - 0x0
    "00000000", -- 2345 - 0x929  :    0 - 0x0
    "00000000", -- 2346 - 0x92a  :    0 - 0x0
    "00000000", -- 2347 - 0x92b  :    0 - 0x0
    "11111010", -- 2348 - 0x92c  :  250 - 0xfa
    "11111110", -- 2349 - 0x92d  :  254 - 0xfe
    "00000011", -- 2350 - 0x92e  :    3 - 0x3
    "00000010", -- 2351 - 0x92f  :    2 - 0x2
    "11111111", -- 2352 - 0x930  :  255 - 0xff -- Sprite 0x93
    "11111110", -- 2353 - 0x931  :  254 - 0xfe
    "00000011", -- 2354 - 0x932  :    3 - 0x3
    "00000110", -- 2355 - 0x933  :    6 - 0x6
    "11111000", -- 2356 - 0x934  :  248 - 0xf8
    "00000000", -- 2357 - 0x935  :    0 - 0x0
    "00000000", -- 2358 - 0x936  :    0 - 0x0
    "00000000", -- 2359 - 0x937  :    0 - 0x0
    "00000010", -- 2360 - 0x938  :    2 - 0x2
    "00000011", -- 2361 - 0x939  :    3 - 0x3
    "11111110", -- 2362 - 0x93a  :  254 - 0xfe
    "11111010", -- 2363 - 0x93b  :  250 - 0xfa
    "00000000", -- 2364 - 0x93c  :    0 - 0x0
    "00000000", -- 2365 - 0x93d  :    0 - 0x0
    "00000000", -- 2366 - 0x93e  :    0 - 0x0
    "00000000", -- 2367 - 0x93f  :    0 - 0x0
    "00000000", -- 2368 - 0x940  :    0 - 0x0 -- Sprite 0x94
    "00000000", -- 2369 - 0x941  :    0 - 0x0
    "00000000", -- 2370 - 0x942  :    0 - 0x0
    "00000000", -- 2371 - 0x943  :    0 - 0x0
    "00101111", -- 2372 - 0x944  :   47 - 0x2f
    "00111111", -- 2373 - 0x945  :   63 - 0x3f
    "01100000", -- 2374 - 0x946  :   96 - 0x60
    "00100000", -- 2375 - 0x947  :   32 - 0x20
    "00000000", -- 2376 - 0x948  :    0 - 0x0
    "00000000", -- 2377 - 0x949  :    0 - 0x0
    "00000000", -- 2378 - 0x94a  :    0 - 0x0
    "00001111", -- 2379 - 0x94b  :   15 - 0xf
    "00110000", -- 2380 - 0x94c  :   48 - 0x30
    "01100000", -- 2381 - 0x94d  :   96 - 0x60
    "00111111", -- 2382 - 0x94e  :   63 - 0x3f
    "01111111", -- 2383 - 0x94f  :  127 - 0x7f
    "00100000", -- 2384 - 0x950  :   32 - 0x20 -- Sprite 0x95
    "01100000", -- 2385 - 0x951  :   96 - 0x60
    "00111111", -- 2386 - 0x952  :   63 - 0x3f
    "00101111", -- 2387 - 0x953  :   47 - 0x2f
    "00000000", -- 2388 - 0x954  :    0 - 0x0
    "00000000", -- 2389 - 0x955  :    0 - 0x0
    "00000000", -- 2390 - 0x956  :    0 - 0x0
    "00000000", -- 2391 - 0x957  :    0 - 0x0
    "01111111", -- 2392 - 0x958  :  127 - 0x7f
    "00111111", -- 2393 - 0x959  :   63 - 0x3f
    "01100000", -- 2394 - 0x95a  :   96 - 0x60
    "00110000", -- 2395 - 0x95b  :   48 - 0x30
    "00001111", -- 2396 - 0x95c  :   15 - 0xf
    "00000000", -- 2397 - 0x95d  :    0 - 0x0
    "00000000", -- 2398 - 0x95e  :    0 - 0x0
    "00000000", -- 2399 - 0x95f  :    0 - 0x0
    "00000000", -- 2400 - 0x960  :    0 - 0x0 -- Sprite 0x96
    "00000000", -- 2401 - 0x961  :    0 - 0x0
    "00000000", -- 2402 - 0x962  :    0 - 0x0
    "00000000", -- 2403 - 0x963  :    0 - 0x0
    "11111010", -- 2404 - 0x964  :  250 - 0xfa
    "11111110", -- 2405 - 0x965  :  254 - 0xfe
    "00000011", -- 2406 - 0x966  :    3 - 0x3
    "00000010", -- 2407 - 0x967  :    2 - 0x2
    "00000000", -- 2408 - 0x968  :    0 - 0x0
    "00000000", -- 2409 - 0x969  :    0 - 0x0
    "00000000", -- 2410 - 0x96a  :    0 - 0x0
    "11111000", -- 2411 - 0x96b  :  248 - 0xf8
    "00000110", -- 2412 - 0x96c  :    6 - 0x6
    "00000011", -- 2413 - 0x96d  :    3 - 0x3
    "11111110", -- 2414 - 0x96e  :  254 - 0xfe
    "11111111", -- 2415 - 0x96f  :  255 - 0xff
    "00000010", -- 2416 - 0x970  :    2 - 0x2 -- Sprite 0x97
    "00000011", -- 2417 - 0x971  :    3 - 0x3
    "11111110", -- 2418 - 0x972  :  254 - 0xfe
    "11111010", -- 2419 - 0x973  :  250 - 0xfa
    "00000000", -- 2420 - 0x974  :    0 - 0x0
    "00000000", -- 2421 - 0x975  :    0 - 0x0
    "00000000", -- 2422 - 0x976  :    0 - 0x0
    "00000000", -- 2423 - 0x977  :    0 - 0x0
    "11111111", -- 2424 - 0x978  :  255 - 0xff
    "11111110", -- 2425 - 0x979  :  254 - 0xfe
    "00000011", -- 2426 - 0x97a  :    3 - 0x3
    "00000110", -- 2427 - 0x97b  :    6 - 0x6
    "11111000", -- 2428 - 0x97c  :  248 - 0xf8
    "00000000", -- 2429 - 0x97d  :    0 - 0x0
    "00000000", -- 2430 - 0x97e  :    0 - 0x0
    "00000000", -- 2431 - 0x97f  :    0 - 0x0
    "00000000", -- 2432 - 0x980  :    0 - 0x0 -- Sprite 0x98
    "01000100", -- 2433 - 0x981  :   68 - 0x44
    "00000000", -- 2434 - 0x982  :    0 - 0x0
    "01000001", -- 2435 - 0x983  :   65 - 0x41
    "00100000", -- 2436 - 0x984  :   32 - 0x20
    "01001011", -- 2437 - 0x985  :   75 - 0x4b
    "00100111", -- 2438 - 0x986  :   39 - 0x27
    "00011111", -- 2439 - 0x987  :   31 - 0x1f
    "00000000", -- 2440 - 0x988  :    0 - 0x0
    "00000000", -- 2441 - 0x989  :    0 - 0x0
    "00000000", -- 2442 - 0x98a  :    0 - 0x0
    "01000000", -- 2443 - 0x98b  :   64 - 0x40
    "00100000", -- 2444 - 0x98c  :   32 - 0x20
    "00000000", -- 2445 - 0x98d  :    0 - 0x0
    "00000000", -- 2446 - 0x98e  :    0 - 0x0
    "00000001", -- 2447 - 0x98f  :    1 - 0x1
    "00001111", -- 2448 - 0x990  :   15 - 0xf -- Sprite 0x99
    "00011110", -- 2449 - 0x991  :   30 - 0x1e
    "00011111", -- 2450 - 0x992  :   31 - 0x1f
    "00011111", -- 2451 - 0x993  :   31 - 0x1f
    "00011111", -- 2452 - 0x994  :   31 - 0x1f
    "00001111", -- 2453 - 0x995  :   15 - 0xf
    "00001111", -- 2454 - 0x996  :   15 - 0xf
    "00000011", -- 2455 - 0x997  :    3 - 0x3
    "00000011", -- 2456 - 0x998  :    3 - 0x3
    "00000111", -- 2457 - 0x999  :    7 - 0x7
    "00000110", -- 2458 - 0x99a  :    6 - 0x6
    "00000110", -- 2459 - 0x99b  :    6 - 0x6
    "00000111", -- 2460 - 0x99c  :    7 - 0x7
    "00000011", -- 2461 - 0x99d  :    3 - 0x3
    "00000000", -- 2462 - 0x99e  :    0 - 0x0
    "00000000", -- 2463 - 0x99f  :    0 - 0x0
    "00000000", -- 2464 - 0x9a0  :    0 - 0x0 -- Sprite 0x9a
    "00100000", -- 2465 - 0x9a1  :   32 - 0x20
    "01010000", -- 2466 - 0x9a2  :   80 - 0x50
    "00100000", -- 2467 - 0x9a3  :   32 - 0x20
    "01100000", -- 2468 - 0x9a4  :   96 - 0x60
    "01001000", -- 2469 - 0x9a5  :   72 - 0x48
    "11100000", -- 2470 - 0x9a6  :  224 - 0xe0
    "11110000", -- 2471 - 0x9a7  :  240 - 0xf0
    "00000000", -- 2472 - 0x9a8  :    0 - 0x0
    "00000000", -- 2473 - 0x9a9  :    0 - 0x0
    "01000000", -- 2474 - 0x9aa  :   64 - 0x40
    "00000000", -- 2475 - 0x9ab  :    0 - 0x0
    "00000000", -- 2476 - 0x9ac  :    0 - 0x0
    "00001000", -- 2477 - 0x9ad  :    8 - 0x8
    "00000000", -- 2478 - 0x9ae  :    0 - 0x0
    "01000000", -- 2479 - 0x9af  :   64 - 0x40
    "11111000", -- 2480 - 0x9b0  :  248 - 0xf8 -- Sprite 0x9b
    "01111000", -- 2481 - 0x9b1  :  120 - 0x78
    "00111100", -- 2482 - 0x9b2  :   60 - 0x3c
    "00111100", -- 2483 - 0x9b3  :   60 - 0x3c
    "00111100", -- 2484 - 0x9b4  :   60 - 0x3c
    "11111100", -- 2485 - 0x9b5  :  252 - 0xfc
    "11111000", -- 2486 - 0x9b6  :  248 - 0xf8
    "11100000", -- 2487 - 0x9b7  :  224 - 0xe0
    "11100000", -- 2488 - 0x9b8  :  224 - 0xe0
    "11110000", -- 2489 - 0x9b9  :  240 - 0xf0
    "11010000", -- 2490 - 0x9ba  :  208 - 0xd0
    "11010000", -- 2491 - 0x9bb  :  208 - 0xd0
    "11110000", -- 2492 - 0x9bc  :  240 - 0xf0
    "11100000", -- 2493 - 0x9bd  :  224 - 0xe0
    "00000000", -- 2494 - 0x9be  :    0 - 0x0
    "00000000", -- 2495 - 0x9bf  :    0 - 0x0
    "00010000", -- 2496 - 0x9c0  :   16 - 0x10 -- Sprite 0x9c
    "00000001", -- 2497 - 0x9c1  :    1 - 0x1
    "00101010", -- 2498 - 0x9c2  :   42 - 0x2a
    "00001100", -- 2499 - 0x9c3  :   12 - 0xc
    "10100110", -- 2500 - 0x9c4  :  166 - 0xa6
    "00010111", -- 2501 - 0x9c5  :   23 - 0x17
    "00011111", -- 2502 - 0x9c6  :   31 - 0x1f
    "00011111", -- 2503 - 0x9c7  :   31 - 0x1f
    "00000000", -- 2504 - 0x9c8  :    0 - 0x0
    "00000000", -- 2505 - 0x9c9  :    0 - 0x0
    "00000010", -- 2506 - 0x9ca  :    2 - 0x2
    "00000000", -- 2507 - 0x9cb  :    0 - 0x0
    "10000000", -- 2508 - 0x9cc  :  128 - 0x80
    "00000000", -- 2509 - 0x9cd  :    0 - 0x0
    "00000011", -- 2510 - 0x9ce  :    3 - 0x3
    "00000111", -- 2511 - 0x9cf  :    7 - 0x7
    "01011110", -- 2512 - 0x9d0  :   94 - 0x5e -- Sprite 0x9d
    "00111100", -- 2513 - 0x9d1  :   60 - 0x3c
    "00111101", -- 2514 - 0x9d2  :   61 - 0x3d
    "00111101", -- 2515 - 0x9d3  :   61 - 0x3d
    "00111110", -- 2516 - 0x9d4  :   62 - 0x3e
    "00011111", -- 2517 - 0x9d5  :   31 - 0x1f
    "00001111", -- 2518 - 0x9d6  :   15 - 0xf
    "00000111", -- 2519 - 0x9d7  :    7 - 0x7
    "00000111", -- 2520 - 0x9d8  :    7 - 0x7
    "00001111", -- 2521 - 0x9d9  :   15 - 0xf
    "00001110", -- 2522 - 0x9da  :   14 - 0xe
    "00001110", -- 2523 - 0x9db  :   14 - 0xe
    "00001111", -- 2524 - 0x9dc  :   15 - 0xf
    "00000111", -- 2525 - 0x9dd  :    7 - 0x7
    "00000011", -- 2526 - 0x9de  :    3 - 0x3
    "00000000", -- 2527 - 0x9df  :    0 - 0x0
    "00000000", -- 2528 - 0x9e0  :    0 - 0x0 -- Sprite 0x9e
    "00000000", -- 2529 - 0x9e1  :    0 - 0x0
    "10000000", -- 2530 - 0x9e2  :  128 - 0x80
    "11001000", -- 2531 - 0x9e3  :  200 - 0xc8
    "01100000", -- 2532 - 0x9e4  :   96 - 0x60
    "11100000", -- 2533 - 0x9e5  :  224 - 0xe0
    "11110100", -- 2534 - 0x9e6  :  244 - 0xf4
    "11111000", -- 2535 - 0x9e7  :  248 - 0xf8
    "00000000", -- 2536 - 0x9e8  :    0 - 0x0
    "00000000", -- 2537 - 0x9e9  :    0 - 0x0
    "00000000", -- 2538 - 0x9ea  :    0 - 0x0
    "00001000", -- 2539 - 0x9eb  :    8 - 0x8
    "00000000", -- 2540 - 0x9ec  :    0 - 0x0
    "10000000", -- 2541 - 0x9ed  :  128 - 0x80
    "00100100", -- 2542 - 0x9ee  :   36 - 0x24
    "11000000", -- 2543 - 0x9ef  :  192 - 0xc0
    "01111100", -- 2544 - 0x9f0  :  124 - 0x7c -- Sprite 0x9f
    "00011100", -- 2545 - 0x9f1  :   28 - 0x1c
    "00101110", -- 2546 - 0x9f2  :   46 - 0x2e
    "00101110", -- 2547 - 0x9f3  :   46 - 0x2e
    "00011110", -- 2548 - 0x9f4  :   30 - 0x1e
    "11111100", -- 2549 - 0x9f5  :  252 - 0xfc
    "11111000", -- 2550 - 0x9f6  :  248 - 0xf8
    "11100000", -- 2551 - 0x9f7  :  224 - 0xe0
    "11110000", -- 2552 - 0x9f8  :  240 - 0xf0
    "11111000", -- 2553 - 0x9f9  :  248 - 0xf8
    "11011000", -- 2554 - 0x9fa  :  216 - 0xd8
    "11011000", -- 2555 - 0x9fb  :  216 - 0xd8
    "11111000", -- 2556 - 0x9fc  :  248 - 0xf8
    "11110000", -- 2557 - 0x9fd  :  240 - 0xf0
    "11000000", -- 2558 - 0x9fe  :  192 - 0xc0
    "00000000", -- 2559 - 0x9ff  :    0 - 0x0
    "11111111", -- 2560 - 0xa00  :  255 - 0xff -- Sprite 0xa0
    "11111111", -- 2561 - 0xa01  :  255 - 0xff
    "00111000", -- 2562 - 0xa02  :   56 - 0x38
    "01101100", -- 2563 - 0xa03  :  108 - 0x6c
    "11000110", -- 2564 - 0xa04  :  198 - 0xc6
    "10000011", -- 2565 - 0xa05  :  131 - 0x83
    "11111111", -- 2566 - 0xa06  :  255 - 0xff
    "11111111", -- 2567 - 0xa07  :  255 - 0xff
    "11111111", -- 2568 - 0xa08  :  255 - 0xff
    "11111111", -- 2569 - 0xa09  :  255 - 0xff
    "00111000", -- 2570 - 0xa0a  :   56 - 0x38
    "01101100", -- 2571 - 0xa0b  :  108 - 0x6c
    "11000110", -- 2572 - 0xa0c  :  198 - 0xc6
    "10000011", -- 2573 - 0xa0d  :  131 - 0x83
    "11111111", -- 2574 - 0xa0e  :  255 - 0xff
    "11111111", -- 2575 - 0xa0f  :  255 - 0xff
    "11111111", -- 2576 - 0xa10  :  255 - 0xff -- Sprite 0xa1
    "11111111", -- 2577 - 0xa11  :  255 - 0xff
    "00111000", -- 2578 - 0xa12  :   56 - 0x38
    "01101100", -- 2579 - 0xa13  :  108 - 0x6c
    "11000110", -- 2580 - 0xa14  :  198 - 0xc6
    "10000011", -- 2581 - 0xa15  :  131 - 0x83
    "11111111", -- 2582 - 0xa16  :  255 - 0xff
    "11111111", -- 2583 - 0xa17  :  255 - 0xff
    "11111111", -- 2584 - 0xa18  :  255 - 0xff
    "11111111", -- 2585 - 0xa19  :  255 - 0xff
    "00111000", -- 2586 - 0xa1a  :   56 - 0x38
    "01101100", -- 2587 - 0xa1b  :  108 - 0x6c
    "11000110", -- 2588 - 0xa1c  :  198 - 0xc6
    "10000011", -- 2589 - 0xa1d  :  131 - 0x83
    "11111111", -- 2590 - 0xa1e  :  255 - 0xff
    "11111111", -- 2591 - 0xa1f  :  255 - 0xff
    "10010010", -- 2592 - 0xa20  :  146 - 0x92 -- Sprite 0xa2
    "01010100", -- 2593 - 0xa21  :   84 - 0x54
    "00111000", -- 2594 - 0xa22  :   56 - 0x38
    "11111110", -- 2595 - 0xa23  :  254 - 0xfe
    "00111000", -- 2596 - 0xa24  :   56 - 0x38
    "01010100", -- 2597 - 0xa25  :   84 - 0x54
    "10010010", -- 2598 - 0xa26  :  146 - 0x92
    "00000000", -- 2599 - 0xa27  :    0 - 0x0
    "00000000", -- 2600 - 0xa28  :    0 - 0x0
    "00000000", -- 2601 - 0xa29  :    0 - 0x0
    "00000000", -- 2602 - 0xa2a  :    0 - 0x0
    "00000000", -- 2603 - 0xa2b  :    0 - 0x0
    "00000000", -- 2604 - 0xa2c  :    0 - 0x0
    "00000000", -- 2605 - 0xa2d  :    0 - 0x0
    "00000000", -- 2606 - 0xa2e  :    0 - 0x0
    "00000000", -- 2607 - 0xa2f  :    0 - 0x0
    "11111111", -- 2608 - 0xa30  :  255 - 0xff -- Sprite 0xa3
    "11111111", -- 2609 - 0xa31  :  255 - 0xff
    "11111111", -- 2610 - 0xa32  :  255 - 0xff
    "11111111", -- 2611 - 0xa33  :  255 - 0xff
    "11111111", -- 2612 - 0xa34  :  255 - 0xff
    "11111111", -- 2613 - 0xa35  :  255 - 0xff
    "11111111", -- 2614 - 0xa36  :  255 - 0xff
    "11111111", -- 2615 - 0xa37  :  255 - 0xff
    "11111111", -- 2616 - 0xa38  :  255 - 0xff
    "11111111", -- 2617 - 0xa39  :  255 - 0xff
    "11111111", -- 2618 - 0xa3a  :  255 - 0xff
    "11111111", -- 2619 - 0xa3b  :  255 - 0xff
    "11111111", -- 2620 - 0xa3c  :  255 - 0xff
    "11111111", -- 2621 - 0xa3d  :  255 - 0xff
    "11111111", -- 2622 - 0xa3e  :  255 - 0xff
    "11111111", -- 2623 - 0xa3f  :  255 - 0xff
    "11111111", -- 2624 - 0xa40  :  255 - 0xff -- Sprite 0xa4
    "11111111", -- 2625 - 0xa41  :  255 - 0xff
    "11111111", -- 2626 - 0xa42  :  255 - 0xff
    "11111111", -- 2627 - 0xa43  :  255 - 0xff
    "11111111", -- 2628 - 0xa44  :  255 - 0xff
    "11111111", -- 2629 - 0xa45  :  255 - 0xff
    "11111111", -- 2630 - 0xa46  :  255 - 0xff
    "11111111", -- 2631 - 0xa47  :  255 - 0xff
    "11111111", -- 2632 - 0xa48  :  255 - 0xff
    "11111111", -- 2633 - 0xa49  :  255 - 0xff
    "11111111", -- 2634 - 0xa4a  :  255 - 0xff
    "11111111", -- 2635 - 0xa4b  :  255 - 0xff
    "11111111", -- 2636 - 0xa4c  :  255 - 0xff
    "11111111", -- 2637 - 0xa4d  :  255 - 0xff
    "11111111", -- 2638 - 0xa4e  :  255 - 0xff
    "11111111", -- 2639 - 0xa4f  :  255 - 0xff
    "11111111", -- 2640 - 0xa50  :  255 - 0xff -- Sprite 0xa5
    "11111111", -- 2641 - 0xa51  :  255 - 0xff
    "11111111", -- 2642 - 0xa52  :  255 - 0xff
    "11111111", -- 2643 - 0xa53  :  255 - 0xff
    "11111111", -- 2644 - 0xa54  :  255 - 0xff
    "11111111", -- 2645 - 0xa55  :  255 - 0xff
    "11111111", -- 2646 - 0xa56  :  255 - 0xff
    "11111111", -- 2647 - 0xa57  :  255 - 0xff
    "11111111", -- 2648 - 0xa58  :  255 - 0xff
    "11111111", -- 2649 - 0xa59  :  255 - 0xff
    "11111111", -- 2650 - 0xa5a  :  255 - 0xff
    "11111111", -- 2651 - 0xa5b  :  255 - 0xff
    "11111111", -- 2652 - 0xa5c  :  255 - 0xff
    "11111111", -- 2653 - 0xa5d  :  255 - 0xff
    "11111111", -- 2654 - 0xa5e  :  255 - 0xff
    "11111111", -- 2655 - 0xa5f  :  255 - 0xff
    "11111111", -- 2656 - 0xa60  :  255 - 0xff -- Sprite 0xa6
    "11111111", -- 2657 - 0xa61  :  255 - 0xff
    "11111111", -- 2658 - 0xa62  :  255 - 0xff
    "11111111", -- 2659 - 0xa63  :  255 - 0xff
    "11111111", -- 2660 - 0xa64  :  255 - 0xff
    "11111111", -- 2661 - 0xa65  :  255 - 0xff
    "11111111", -- 2662 - 0xa66  :  255 - 0xff
    "11111111", -- 2663 - 0xa67  :  255 - 0xff
    "11111111", -- 2664 - 0xa68  :  255 - 0xff
    "11111111", -- 2665 - 0xa69  :  255 - 0xff
    "11111111", -- 2666 - 0xa6a  :  255 - 0xff
    "11111111", -- 2667 - 0xa6b  :  255 - 0xff
    "11111111", -- 2668 - 0xa6c  :  255 - 0xff
    "11111111", -- 2669 - 0xa6d  :  255 - 0xff
    "11111111", -- 2670 - 0xa6e  :  255 - 0xff
    "11111111", -- 2671 - 0xa6f  :  255 - 0xff
    "11111111", -- 2672 - 0xa70  :  255 - 0xff -- Sprite 0xa7
    "11111111", -- 2673 - 0xa71  :  255 - 0xff
    "11111111", -- 2674 - 0xa72  :  255 - 0xff
    "11111111", -- 2675 - 0xa73  :  255 - 0xff
    "11111111", -- 2676 - 0xa74  :  255 - 0xff
    "11111111", -- 2677 - 0xa75  :  255 - 0xff
    "11111111", -- 2678 - 0xa76  :  255 - 0xff
    "11111111", -- 2679 - 0xa77  :  255 - 0xff
    "11111111", -- 2680 - 0xa78  :  255 - 0xff
    "11111111", -- 2681 - 0xa79  :  255 - 0xff
    "11111111", -- 2682 - 0xa7a  :  255 - 0xff
    "11111111", -- 2683 - 0xa7b  :  255 - 0xff
    "11111111", -- 2684 - 0xa7c  :  255 - 0xff
    "11111111", -- 2685 - 0xa7d  :  255 - 0xff
    "11111111", -- 2686 - 0xa7e  :  255 - 0xff
    "11111111", -- 2687 - 0xa7f  :  255 - 0xff
    "00000000", -- 2688 - 0xa80  :    0 - 0x0 -- Sprite 0xa8
    "00000000", -- 2689 - 0xa81  :    0 - 0x0
    "00000000", -- 2690 - 0xa82  :    0 - 0x0
    "00000000", -- 2691 - 0xa83  :    0 - 0x0
    "00000000", -- 2692 - 0xa84  :    0 - 0x0
    "00100011", -- 2693 - 0xa85  :   35 - 0x23
    "10010111", -- 2694 - 0xa86  :  151 - 0x97
    "00101111", -- 2695 - 0xa87  :   47 - 0x2f
    "00000000", -- 2696 - 0xa88  :    0 - 0x0
    "00000000", -- 2697 - 0xa89  :    0 - 0x0
    "00000000", -- 2698 - 0xa8a  :    0 - 0x0
    "00000000", -- 2699 - 0xa8b  :    0 - 0x0
    "00000000", -- 2700 - 0xa8c  :    0 - 0x0
    "00000000", -- 2701 - 0xa8d  :    0 - 0x0
    "00000001", -- 2702 - 0xa8e  :    1 - 0x1
    "00000011", -- 2703 - 0xa8f  :    3 - 0x3
    "01101110", -- 2704 - 0xa90  :  110 - 0x6e -- Sprite 0xa9
    "11101111", -- 2705 - 0xa91  :  239 - 0xef
    "11110111", -- 2706 - 0xa92  :  247 - 0xf7
    "11111111", -- 2707 - 0xa93  :  255 - 0xff
    "01111111", -- 2708 - 0xa94  :  127 - 0x7f
    "00111111", -- 2709 - 0xa95  :   63 - 0x3f
    "01011111", -- 2710 - 0xa96  :   95 - 0x5f
    "00001111", -- 2711 - 0xa97  :   15 - 0xf
    "00000111", -- 2712 - 0xa98  :    7 - 0x7
    "00000111", -- 2713 - 0xa99  :    7 - 0x7
    "00000011", -- 2714 - 0xa9a  :    3 - 0x3
    "00100111", -- 2715 - 0xa9b  :   39 - 0x27
    "00011111", -- 2716 - 0xa9c  :   31 - 0x1f
    "00000111", -- 2717 - 0xa9d  :    7 - 0x7
    "00000000", -- 2718 - 0xa9e  :    0 - 0x0
    "00000000", -- 2719 - 0xa9f  :    0 - 0x0
    "00000000", -- 2720 - 0xaa0  :    0 - 0x0 -- Sprite 0xaa
    "00000000", -- 2721 - 0xaa1  :    0 - 0x0
    "00000000", -- 2722 - 0xaa2  :    0 - 0x0
    "00000000", -- 2723 - 0xaa3  :    0 - 0x0
    "11111000", -- 2724 - 0xaa4  :  248 - 0xf8
    "11111100", -- 2725 - 0xaa5  :  252 - 0xfc
    "11111110", -- 2726 - 0xaa6  :  254 - 0xfe
    "01011110", -- 2727 - 0xaa7  :   94 - 0x5e
    "00000000", -- 2728 - 0xaa8  :    0 - 0x0
    "00000000", -- 2729 - 0xaa9  :    0 - 0x0
    "00000000", -- 2730 - 0xaaa  :    0 - 0x0
    "00000000", -- 2731 - 0xaab  :    0 - 0x0
    "00000000", -- 2732 - 0xaac  :    0 - 0x0
    "11110000", -- 2733 - 0xaad  :  240 - 0xf0
    "11111000", -- 2734 - 0xaae  :  248 - 0xf8
    "10101100", -- 2735 - 0xaaf  :  172 - 0xac
    "01011110", -- 2736 - 0xab0  :   94 - 0x5e -- Sprite 0xab
    "00001100", -- 2737 - 0xab1  :   12 - 0xc
    "10011110", -- 2738 - 0xab2  :  158 - 0x9e
    "11111110", -- 2739 - 0xab3  :  254 - 0xfe
    "11111110", -- 2740 - 0xab4  :  254 - 0xfe
    "11111110", -- 2741 - 0xab5  :  254 - 0xfe
    "11111000", -- 2742 - 0xab6  :  248 - 0xf8
    "11000000", -- 2743 - 0xab7  :  192 - 0xc0
    "10101100", -- 2744 - 0xab8  :  172 - 0xac
    "11111000", -- 2745 - 0xab9  :  248 - 0xf8
    "11111000", -- 2746 - 0xaba  :  248 - 0xf8
    "11111000", -- 2747 - 0xabb  :  248 - 0xf8
    "11110000", -- 2748 - 0xabc  :  240 - 0xf0
    "11000000", -- 2749 - 0xabd  :  192 - 0xc0
    "00000000", -- 2750 - 0xabe  :    0 - 0x0
    "00000000", -- 2751 - 0xabf  :    0 - 0x0
    "00000000", -- 2752 - 0xac0  :    0 - 0x0 -- Sprite 0xac
    "00000000", -- 2753 - 0xac1  :    0 - 0x0
    "00000000", -- 2754 - 0xac2  :    0 - 0x0
    "00000000", -- 2755 - 0xac3  :    0 - 0x0
    "00000000", -- 2756 - 0xac4  :    0 - 0x0
    "00000011", -- 2757 - 0xac5  :    3 - 0x3
    "00000111", -- 2758 - 0xac6  :    7 - 0x7
    "00101111", -- 2759 - 0xac7  :   47 - 0x2f
    "00000000", -- 2760 - 0xac8  :    0 - 0x0
    "00000000", -- 2761 - 0xac9  :    0 - 0x0
    "00000000", -- 2762 - 0xaca  :    0 - 0x0
    "00000000", -- 2763 - 0xacb  :    0 - 0x0
    "00000000", -- 2764 - 0xacc  :    0 - 0x0
    "00000000", -- 2765 - 0xacd  :    0 - 0x0
    "00000001", -- 2766 - 0xace  :    1 - 0x1
    "00000011", -- 2767 - 0xacf  :    3 - 0x3
    "01001110", -- 2768 - 0xad0  :   78 - 0x4e -- Sprite 0xad
    "01101110", -- 2769 - 0xad1  :  110 - 0x6e
    "11111110", -- 2770 - 0xad2  :  254 - 0xfe
    "01111111", -- 2771 - 0xad3  :  127 - 0x7f
    "00111111", -- 2772 - 0xad4  :   63 - 0x3f
    "00011111", -- 2773 - 0xad5  :   31 - 0x1f
    "00001111", -- 2774 - 0xad6  :   15 - 0xf
    "00000011", -- 2775 - 0xad7  :    3 - 0x3
    "00000111", -- 2776 - 0xad8  :    7 - 0x7
    "00000111", -- 2777 - 0xad9  :    7 - 0x7
    "00000111", -- 2778 - 0xada  :    7 - 0x7
    "00100111", -- 2779 - 0xadb  :   39 - 0x27
    "00011111", -- 2780 - 0xadc  :   31 - 0x1f
    "00000111", -- 2781 - 0xadd  :    7 - 0x7
    "00000001", -- 2782 - 0xade  :    1 - 0x1
    "00000000", -- 2783 - 0xadf  :    0 - 0x0
    "00000000", -- 2784 - 0xae0  :    0 - 0x0 -- Sprite 0xae
    "00000000", -- 2785 - 0xae1  :    0 - 0x0
    "00000000", -- 2786 - 0xae2  :    0 - 0x0
    "00000000", -- 2787 - 0xae3  :    0 - 0x0
    "11111000", -- 2788 - 0xae4  :  248 - 0xf8
    "11111100", -- 2789 - 0xae5  :  252 - 0xfc
    "11111110", -- 2790 - 0xae6  :  254 - 0xfe
    "01010110", -- 2791 - 0xae7  :   86 - 0x56
    "00000000", -- 2792 - 0xae8  :    0 - 0x0
    "00000000", -- 2793 - 0xae9  :    0 - 0x0
    "00000000", -- 2794 - 0xaea  :    0 - 0x0
    "00000000", -- 2795 - 0xaeb  :    0 - 0x0
    "00000000", -- 2796 - 0xaec  :    0 - 0x0
    "11110000", -- 2797 - 0xaed  :  240 - 0xf0
    "11111000", -- 2798 - 0xaee  :  248 - 0xf8
    "10101100", -- 2799 - 0xaef  :  172 - 0xac
    "01010110", -- 2800 - 0xaf0  :   86 - 0x56 -- Sprite 0xaf
    "00001100", -- 2801 - 0xaf1  :   12 - 0xc
    "00001110", -- 2802 - 0xaf2  :   14 - 0xe
    "00011111", -- 2803 - 0xaf3  :   31 - 0x1f
    "11111111", -- 2804 - 0xaf4  :  255 - 0xff
    "11111111", -- 2805 - 0xaf5  :  255 - 0xff
    "11111110", -- 2806 - 0xaf6  :  254 - 0xfe
    "11111000", -- 2807 - 0xaf7  :  248 - 0xf8
    "10101100", -- 2808 - 0xaf8  :  172 - 0xac
    "11111000", -- 2809 - 0xaf9  :  248 - 0xf8
    "11111000", -- 2810 - 0xafa  :  248 - 0xf8
    "11111100", -- 2811 - 0xafb  :  252 - 0xfc
    "11111100", -- 2812 - 0xafc  :  252 - 0xfc
    "11111000", -- 2813 - 0xafd  :  248 - 0xf8
    "11110000", -- 2814 - 0xafe  :  240 - 0xf0
    "00000000", -- 2815 - 0xaff  :    0 - 0x0
    "11111111", -- 2816 - 0xb00  :  255 - 0xff -- Sprite 0xb0
    "11111111", -- 2817 - 0xb01  :  255 - 0xff
    "11111111", -- 2818 - 0xb02  :  255 - 0xff
    "11111111", -- 2819 - 0xb03  :  255 - 0xff
    "11111111", -- 2820 - 0xb04  :  255 - 0xff
    "11111111", -- 2821 - 0xb05  :  255 - 0xff
    "11111111", -- 2822 - 0xb06  :  255 - 0xff
    "11111111", -- 2823 - 0xb07  :  255 - 0xff
    "11111111", -- 2824 - 0xb08  :  255 - 0xff
    "11111111", -- 2825 - 0xb09  :  255 - 0xff
    "11111111", -- 2826 - 0xb0a  :  255 - 0xff
    "11111111", -- 2827 - 0xb0b  :  255 - 0xff
    "11111111", -- 2828 - 0xb0c  :  255 - 0xff
    "11111111", -- 2829 - 0xb0d  :  255 - 0xff
    "11111111", -- 2830 - 0xb0e  :  255 - 0xff
    "11111111", -- 2831 - 0xb0f  :  255 - 0xff
    "11111111", -- 2832 - 0xb10  :  255 - 0xff -- Sprite 0xb1
    "11111111", -- 2833 - 0xb11  :  255 - 0xff
    "11111111", -- 2834 - 0xb12  :  255 - 0xff
    "11111111", -- 2835 - 0xb13  :  255 - 0xff
    "11111111", -- 2836 - 0xb14  :  255 - 0xff
    "11111111", -- 2837 - 0xb15  :  255 - 0xff
    "11111111", -- 2838 - 0xb16  :  255 - 0xff
    "11111111", -- 2839 - 0xb17  :  255 - 0xff
    "11111111", -- 2840 - 0xb18  :  255 - 0xff
    "11111111", -- 2841 - 0xb19  :  255 - 0xff
    "11111111", -- 2842 - 0xb1a  :  255 - 0xff
    "11111111", -- 2843 - 0xb1b  :  255 - 0xff
    "11111111", -- 2844 - 0xb1c  :  255 - 0xff
    "11111111", -- 2845 - 0xb1d  :  255 - 0xff
    "11111111", -- 2846 - 0xb1e  :  255 - 0xff
    "11111111", -- 2847 - 0xb1f  :  255 - 0xff
    "11111111", -- 2848 - 0xb20  :  255 - 0xff -- Sprite 0xb2
    "11111111", -- 2849 - 0xb21  :  255 - 0xff
    "11111111", -- 2850 - 0xb22  :  255 - 0xff
    "11111111", -- 2851 - 0xb23  :  255 - 0xff
    "11111111", -- 2852 - 0xb24  :  255 - 0xff
    "11111111", -- 2853 - 0xb25  :  255 - 0xff
    "11111111", -- 2854 - 0xb26  :  255 - 0xff
    "11111111", -- 2855 - 0xb27  :  255 - 0xff
    "11111111", -- 2856 - 0xb28  :  255 - 0xff
    "11111111", -- 2857 - 0xb29  :  255 - 0xff
    "11111111", -- 2858 - 0xb2a  :  255 - 0xff
    "11111111", -- 2859 - 0xb2b  :  255 - 0xff
    "11111111", -- 2860 - 0xb2c  :  255 - 0xff
    "11111111", -- 2861 - 0xb2d  :  255 - 0xff
    "11111111", -- 2862 - 0xb2e  :  255 - 0xff
    "11111111", -- 2863 - 0xb2f  :  255 - 0xff
    "11111111", -- 2864 - 0xb30  :  255 - 0xff -- Sprite 0xb3
    "11111111", -- 2865 - 0xb31  :  255 - 0xff
    "11111111", -- 2866 - 0xb32  :  255 - 0xff
    "11111111", -- 2867 - 0xb33  :  255 - 0xff
    "11111111", -- 2868 - 0xb34  :  255 - 0xff
    "11111111", -- 2869 - 0xb35  :  255 - 0xff
    "11111111", -- 2870 - 0xb36  :  255 - 0xff
    "11111111", -- 2871 - 0xb37  :  255 - 0xff
    "11111111", -- 2872 - 0xb38  :  255 - 0xff
    "11111111", -- 2873 - 0xb39  :  255 - 0xff
    "11111111", -- 2874 - 0xb3a  :  255 - 0xff
    "11111111", -- 2875 - 0xb3b  :  255 - 0xff
    "11111111", -- 2876 - 0xb3c  :  255 - 0xff
    "11111111", -- 2877 - 0xb3d  :  255 - 0xff
    "11111111", -- 2878 - 0xb3e  :  255 - 0xff
    "11111111", -- 2879 - 0xb3f  :  255 - 0xff
    "11111111", -- 2880 - 0xb40  :  255 - 0xff -- Sprite 0xb4
    "11111111", -- 2881 - 0xb41  :  255 - 0xff
    "11111111", -- 2882 - 0xb42  :  255 - 0xff
    "11111111", -- 2883 - 0xb43  :  255 - 0xff
    "11111111", -- 2884 - 0xb44  :  255 - 0xff
    "11111111", -- 2885 - 0xb45  :  255 - 0xff
    "11111111", -- 2886 - 0xb46  :  255 - 0xff
    "11111111", -- 2887 - 0xb47  :  255 - 0xff
    "11111111", -- 2888 - 0xb48  :  255 - 0xff
    "11111111", -- 2889 - 0xb49  :  255 - 0xff
    "11111111", -- 2890 - 0xb4a  :  255 - 0xff
    "11111111", -- 2891 - 0xb4b  :  255 - 0xff
    "11111111", -- 2892 - 0xb4c  :  255 - 0xff
    "11111111", -- 2893 - 0xb4d  :  255 - 0xff
    "11111111", -- 2894 - 0xb4e  :  255 - 0xff
    "11111111", -- 2895 - 0xb4f  :  255 - 0xff
    "11111111", -- 2896 - 0xb50  :  255 - 0xff -- Sprite 0xb5
    "11111111", -- 2897 - 0xb51  :  255 - 0xff
    "11111111", -- 2898 - 0xb52  :  255 - 0xff
    "11111111", -- 2899 - 0xb53  :  255 - 0xff
    "11111111", -- 2900 - 0xb54  :  255 - 0xff
    "11111111", -- 2901 - 0xb55  :  255 - 0xff
    "11111111", -- 2902 - 0xb56  :  255 - 0xff
    "11111111", -- 2903 - 0xb57  :  255 - 0xff
    "11111111", -- 2904 - 0xb58  :  255 - 0xff
    "11111111", -- 2905 - 0xb59  :  255 - 0xff
    "11111111", -- 2906 - 0xb5a  :  255 - 0xff
    "11111111", -- 2907 - 0xb5b  :  255 - 0xff
    "11111111", -- 2908 - 0xb5c  :  255 - 0xff
    "11111111", -- 2909 - 0xb5d  :  255 - 0xff
    "11111111", -- 2910 - 0xb5e  :  255 - 0xff
    "11111111", -- 2911 - 0xb5f  :  255 - 0xff
    "11111111", -- 2912 - 0xb60  :  255 - 0xff -- Sprite 0xb6
    "11111111", -- 2913 - 0xb61  :  255 - 0xff
    "11111111", -- 2914 - 0xb62  :  255 - 0xff
    "11111111", -- 2915 - 0xb63  :  255 - 0xff
    "11111111", -- 2916 - 0xb64  :  255 - 0xff
    "11111111", -- 2917 - 0xb65  :  255 - 0xff
    "11111111", -- 2918 - 0xb66  :  255 - 0xff
    "11111111", -- 2919 - 0xb67  :  255 - 0xff
    "11111111", -- 2920 - 0xb68  :  255 - 0xff
    "11111111", -- 2921 - 0xb69  :  255 - 0xff
    "11111111", -- 2922 - 0xb6a  :  255 - 0xff
    "11111111", -- 2923 - 0xb6b  :  255 - 0xff
    "11111111", -- 2924 - 0xb6c  :  255 - 0xff
    "11111111", -- 2925 - 0xb6d  :  255 - 0xff
    "11111111", -- 2926 - 0xb6e  :  255 - 0xff
    "11111111", -- 2927 - 0xb6f  :  255 - 0xff
    "11111111", -- 2928 - 0xb70  :  255 - 0xff -- Sprite 0xb7
    "11111111", -- 2929 - 0xb71  :  255 - 0xff
    "11111111", -- 2930 - 0xb72  :  255 - 0xff
    "11111111", -- 2931 - 0xb73  :  255 - 0xff
    "11111111", -- 2932 - 0xb74  :  255 - 0xff
    "11111111", -- 2933 - 0xb75  :  255 - 0xff
    "11111111", -- 2934 - 0xb76  :  255 - 0xff
    "11111111", -- 2935 - 0xb77  :  255 - 0xff
    "11111111", -- 2936 - 0xb78  :  255 - 0xff
    "11111111", -- 2937 - 0xb79  :  255 - 0xff
    "11111111", -- 2938 - 0xb7a  :  255 - 0xff
    "11111111", -- 2939 - 0xb7b  :  255 - 0xff
    "11111111", -- 2940 - 0xb7c  :  255 - 0xff
    "11111111", -- 2941 - 0xb7d  :  255 - 0xff
    "11111111", -- 2942 - 0xb7e  :  255 - 0xff
    "11111111", -- 2943 - 0xb7f  :  255 - 0xff
    "00000000", -- 2944 - 0xb80  :    0 - 0x0 -- Sprite 0xb8
    "00000111", -- 2945 - 0xb81  :    7 - 0x7
    "00001000", -- 2946 - 0xb82  :    8 - 0x8
    "00010000", -- 2947 - 0xb83  :   16 - 0x10
    "00010000", -- 2948 - 0xb84  :   16 - 0x10
    "00100000", -- 2949 - 0xb85  :   32 - 0x20
    "00100000", -- 2950 - 0xb86  :   32 - 0x20
    "00100000", -- 2951 - 0xb87  :   32 - 0x20
    "00000000", -- 2952 - 0xb88  :    0 - 0x0
    "00000111", -- 2953 - 0xb89  :    7 - 0x7
    "00001000", -- 2954 - 0xb8a  :    8 - 0x8
    "00010000", -- 2955 - 0xb8b  :   16 - 0x10
    "00010000", -- 2956 - 0xb8c  :   16 - 0x10
    "00100000", -- 2957 - 0xb8d  :   32 - 0x20
    "00100000", -- 2958 - 0xb8e  :   32 - 0x20
    "00100000", -- 2959 - 0xb8f  :   32 - 0x20
    "00011111", -- 2960 - 0xb90  :   31 - 0x1f -- Sprite 0xb9
    "00101111", -- 2961 - 0xb91  :   47 - 0x2f
    "00110111", -- 2962 - 0xb92  :   55 - 0x37
    "00111010", -- 2963 - 0xb93  :   58 - 0x3a
    "00111101", -- 2964 - 0xb94  :   61 - 0x3d
    "00111110", -- 2965 - 0xb95  :   62 - 0x3e
    "00111111", -- 2966 - 0xb96  :   63 - 0x3f
    "00000000", -- 2967 - 0xb97  :    0 - 0x0
    "00011111", -- 2968 - 0xb98  :   31 - 0x1f
    "00111111", -- 2969 - 0xb99  :   63 - 0x3f
    "00111111", -- 2970 - 0xb9a  :   63 - 0x3f
    "00111111", -- 2971 - 0xb9b  :   63 - 0x3f
    "00111110", -- 2972 - 0xb9c  :   62 - 0x3e
    "00111111", -- 2973 - 0xb9d  :   63 - 0x3f
    "00111111", -- 2974 - 0xb9e  :   63 - 0x3f
    "00000000", -- 2975 - 0xb9f  :    0 - 0x0
    "00000000", -- 2976 - 0xba0  :    0 - 0x0 -- Sprite 0xba
    "00000101", -- 2977 - 0xba1  :    5 - 0x5
    "00011001", -- 2978 - 0xba2  :   25 - 0x19
    "00110011", -- 2979 - 0xba3  :   51 - 0x33
    "01100011", -- 2980 - 0xba4  :   99 - 0x63
    "11000111", -- 2981 - 0xba5  :  199 - 0xc7
    "11000111", -- 2982 - 0xba6  :  199 - 0xc7
    "11000100", -- 2983 - 0xba7  :  196 - 0xc4
    "00000000", -- 2984 - 0xba8  :    0 - 0x0
    "00000111", -- 2985 - 0xba9  :    7 - 0x7
    "00011111", -- 2986 - 0xbaa  :   31 - 0x1f
    "00111111", -- 2987 - 0xbab  :   63 - 0x3f
    "01111111", -- 2988 - 0xbac  :  127 - 0x7f
    "11111111", -- 2989 - 0xbad  :  255 - 0xff
    "11111111", -- 2990 - 0xbae  :  255 - 0xff
    "11011101", -- 2991 - 0xbaf  :  221 - 0xdd
    "10000000", -- 2992 - 0xbb0  :  128 - 0x80 -- Sprite 0xbb
    "00000000", -- 2993 - 0xbb1  :    0 - 0x0
    "00000000", -- 2994 - 0xbb2  :    0 - 0x0
    "00000000", -- 2995 - 0xbb3  :    0 - 0x0
    "00000000", -- 2996 - 0xbb4  :    0 - 0x0
    "00000011", -- 2997 - 0xbb5  :    3 - 0x3
    "00000011", -- 2998 - 0xbb6  :    3 - 0x3
    "00000000", -- 2999 - 0xbb7  :    0 - 0x0
    "10001001", -- 3000 - 0xbb8  :  137 - 0x89
    "00000001", -- 3001 - 0xbb9  :    1 - 0x1
    "00000001", -- 3002 - 0xbba  :    1 - 0x1
    "00000001", -- 3003 - 0xbbb  :    1 - 0x1
    "00000001", -- 3004 - 0xbbc  :    1 - 0x1
    "00000000", -- 3005 - 0xbbd  :    0 - 0x0
    "00000000", -- 3006 - 0xbbe  :    0 - 0x0
    "00000000", -- 3007 - 0xbbf  :    0 - 0x0
    "00000000", -- 3008 - 0xbc0  :    0 - 0x0 -- Sprite 0xbc
    "00000000", -- 3009 - 0xbc1  :    0 - 0x0
    "00000000", -- 3010 - 0xbc2  :    0 - 0x0
    "00000000", -- 3011 - 0xbc3  :    0 - 0x0
    "00000000", -- 3012 - 0xbc4  :    0 - 0x0
    "00000000", -- 3013 - 0xbc5  :    0 - 0x0
    "00000000", -- 3014 - 0xbc6  :    0 - 0x0
    "00000000", -- 3015 - 0xbc7  :    0 - 0x0
    "00000000", -- 3016 - 0xbc8  :    0 - 0x0
    "00000000", -- 3017 - 0xbc9  :    0 - 0x0
    "00000000", -- 3018 - 0xbca  :    0 - 0x0
    "00000000", -- 3019 - 0xbcb  :    0 - 0x0
    "00000000", -- 3020 - 0xbcc  :    0 - 0x0
    "00000000", -- 3021 - 0xbcd  :    0 - 0x0
    "00000011", -- 3022 - 0xbce  :    3 - 0x3
    "00000111", -- 3023 - 0xbcf  :    7 - 0x7
    "00000000", -- 3024 - 0xbd0  :    0 - 0x0 -- Sprite 0xbd
    "00000000", -- 3025 - 0xbd1  :    0 - 0x0
    "00001111", -- 3026 - 0xbd2  :   15 - 0xf
    "00000000", -- 3027 - 0xbd3  :    0 - 0x0
    "10000000", -- 3028 - 0xbd4  :  128 - 0x80
    "01100011", -- 3029 - 0xbd5  :   99 - 0x63
    "00011110", -- 3030 - 0xbd6  :   30 - 0x1e
    "00000000", -- 3031 - 0xbd7  :    0 - 0x0
    "00001111", -- 3032 - 0xbd8  :   15 - 0xf
    "00001111", -- 3033 - 0xbd9  :   15 - 0xf
    "00000000", -- 3034 - 0xbda  :    0 - 0x0
    "00011111", -- 3035 - 0xbdb  :   31 - 0x1f
    "01111111", -- 3036 - 0xbdc  :  127 - 0x7f
    "00011100", -- 3037 - 0xbdd  :   28 - 0x1c
    "00000000", -- 3038 - 0xbde  :    0 - 0x0
    "00000000", -- 3039 - 0xbdf  :    0 - 0x0
    "00000001", -- 3040 - 0xbe0  :    1 - 0x1 -- Sprite 0xbe
    "00000011", -- 3041 - 0xbe1  :    3 - 0x3
    "00011001", -- 3042 - 0xbe2  :   25 - 0x19
    "00111100", -- 3043 - 0xbe3  :   60 - 0x3c
    "00011001", -- 3044 - 0xbe4  :   25 - 0x19
    "00100011", -- 3045 - 0xbe5  :   35 - 0x23
    "01010001", -- 3046 - 0xbe6  :   81 - 0x51
    "00100000", -- 3047 - 0xbe7  :   32 - 0x20
    "00000001", -- 3048 - 0xbe8  :    1 - 0x1
    "00000010", -- 3049 - 0xbe9  :    2 - 0x2
    "00011001", -- 3050 - 0xbea  :   25 - 0x19
    "00100100", -- 3051 - 0xbeb  :   36 - 0x24
    "00011001", -- 3052 - 0xbec  :   25 - 0x19
    "00100010", -- 3053 - 0xbed  :   34 - 0x22
    "00010001", -- 3054 - 0xbee  :   17 - 0x11
    "00101100", -- 3055 - 0xbef  :   44 - 0x2c
    "00000000", -- 3056 - 0xbf0  :    0 - 0x0 -- Sprite 0xbf
    "00000000", -- 3057 - 0xbf1  :    0 - 0x0
    "00000000", -- 3058 - 0xbf2  :    0 - 0x0
    "00000000", -- 3059 - 0xbf3  :    0 - 0x0
    "00000000", -- 3060 - 0xbf4  :    0 - 0x0
    "00000000", -- 3061 - 0xbf5  :    0 - 0x0
    "00000000", -- 3062 - 0xbf6  :    0 - 0x0
    "00000000", -- 3063 - 0xbf7  :    0 - 0x0
    "00011111", -- 3064 - 0xbf8  :   31 - 0x1f
    "00000111", -- 3065 - 0xbf9  :    7 - 0x7
    "00000011", -- 3066 - 0xbfa  :    3 - 0x3
    "00000011", -- 3067 - 0xbfb  :    3 - 0x3
    "00000001", -- 3068 - 0xbfc  :    1 - 0x1
    "00000001", -- 3069 - 0xbfd  :    1 - 0x1
    "00000001", -- 3070 - 0xbfe  :    1 - 0x1
    "00000000", -- 3071 - 0xbff  :    0 - 0x0
    "00000000", -- 3072 - 0xc00  :    0 - 0x0 -- Sprite 0xc0
    "00111111", -- 3073 - 0xc01  :   63 - 0x3f
    "00011111", -- 3074 - 0xc02  :   31 - 0x1f
    "00000000", -- 3075 - 0xc03  :    0 - 0x0
    "00000001", -- 3076 - 0xc04  :    1 - 0x1
    "00000000", -- 3077 - 0xc05  :    0 - 0x0
    "00000001", -- 3078 - 0xc06  :    1 - 0x1
    "00000000", -- 3079 - 0xc07  :    0 - 0x0
    "00000000", -- 3080 - 0xc08  :    0 - 0x0
    "00000000", -- 3081 - 0xc09  :    0 - 0x0
    "00000000", -- 3082 - 0xc0a  :    0 - 0x0
    "00000001", -- 3083 - 0xc0b  :    1 - 0x1
    "00000011", -- 3084 - 0xc0c  :    3 - 0x3
    "00000111", -- 3085 - 0xc0d  :    7 - 0x7
    "00001101", -- 3086 - 0xc0e  :   13 - 0xd
    "00011001", -- 3087 - 0xc0f  :   25 - 0x19
    "00010001", -- 3088 - 0xc10  :   17 - 0x11 -- Sprite 0xc1
    "00000000", -- 3089 - 0xc11  :    0 - 0x0
    "00000001", -- 3090 - 0xc12  :    1 - 0x1
    "00000000", -- 3091 - 0xc13  :    0 - 0x0
    "00000001", -- 3092 - 0xc14  :    1 - 0x1
    "00000000", -- 3093 - 0xc15  :    0 - 0x0
    "00011111", -- 3094 - 0xc16  :   31 - 0x1f
    "00111111", -- 3095 - 0xc17  :   63 - 0x3f
    "00101001", -- 3096 - 0xc18  :   41 - 0x29
    "00011001", -- 3097 - 0xc19  :   25 - 0x19
    "00001101", -- 3098 - 0xc1a  :   13 - 0xd
    "00000111", -- 3099 - 0xc1b  :    7 - 0x7
    "00000011", -- 3100 - 0xc1c  :    3 - 0x3
    "00000001", -- 3101 - 0xc1d  :    1 - 0x1
    "00000000", -- 3102 - 0xc1e  :    0 - 0x0
    "00000000", -- 3103 - 0xc1f  :    0 - 0x0
    "00000000", -- 3104 - 0xc20  :    0 - 0x0 -- Sprite 0xc2
    "11111100", -- 3105 - 0xc21  :  252 - 0xfc
    "11111000", -- 3106 - 0xc22  :  248 - 0xf8
    "00000000", -- 3107 - 0xc23  :    0 - 0x0
    "10000000", -- 3108 - 0xc24  :  128 - 0x80
    "00000000", -- 3109 - 0xc25  :    0 - 0x0
    "10000000", -- 3110 - 0xc26  :  128 - 0x80
    "00000000", -- 3111 - 0xc27  :    0 - 0x0
    "00000000", -- 3112 - 0xc28  :    0 - 0x0
    "00000000", -- 3113 - 0xc29  :    0 - 0x0
    "00000000", -- 3114 - 0xc2a  :    0 - 0x0
    "10000000", -- 3115 - 0xc2b  :  128 - 0x80
    "11000000", -- 3116 - 0xc2c  :  192 - 0xc0
    "11100000", -- 3117 - 0xc2d  :  224 - 0xe0
    "10110000", -- 3118 - 0xc2e  :  176 - 0xb0
    "10011000", -- 3119 - 0xc2f  :  152 - 0x98
    "10001000", -- 3120 - 0xc30  :  136 - 0x88 -- Sprite 0xc3
    "00000000", -- 3121 - 0xc31  :    0 - 0x0
    "10000000", -- 3122 - 0xc32  :  128 - 0x80
    "00000000", -- 3123 - 0xc33  :    0 - 0x0
    "10000000", -- 3124 - 0xc34  :  128 - 0x80
    "00000000", -- 3125 - 0xc35  :    0 - 0x0
    "11111000", -- 3126 - 0xc36  :  248 - 0xf8
    "11111100", -- 3127 - 0xc37  :  252 - 0xfc
    "10010100", -- 3128 - 0xc38  :  148 - 0x94
    "10011000", -- 3129 - 0xc39  :  152 - 0x98
    "10110000", -- 3130 - 0xc3a  :  176 - 0xb0
    "11100000", -- 3131 - 0xc3b  :  224 - 0xe0
    "11000000", -- 3132 - 0xc3c  :  192 - 0xc0
    "10000000", -- 3133 - 0xc3d  :  128 - 0x80
    "00000000", -- 3134 - 0xc3e  :    0 - 0x0
    "00000000", -- 3135 - 0xc3f  :    0 - 0x0
    "00000000", -- 3136 - 0xc40  :    0 - 0x0 -- Sprite 0xc4
    "00000000", -- 3137 - 0xc41  :    0 - 0x0
    "00000000", -- 3138 - 0xc42  :    0 - 0x0
    "00000000", -- 3139 - 0xc43  :    0 - 0x0
    "00000000", -- 3140 - 0xc44  :    0 - 0x0
    "00111111", -- 3141 - 0xc45  :   63 - 0x3f
    "00011111", -- 3142 - 0xc46  :   31 - 0x1f
    "00000000", -- 3143 - 0xc47  :    0 - 0x0
    "00000000", -- 3144 - 0xc48  :    0 - 0x0
    "00000000", -- 3145 - 0xc49  :    0 - 0x0
    "00000000", -- 3146 - 0xc4a  :    0 - 0x0
    "00000000", -- 3147 - 0xc4b  :    0 - 0x0
    "00000000", -- 3148 - 0xc4c  :    0 - 0x0
    "00000000", -- 3149 - 0xc4d  :    0 - 0x0
    "00000000", -- 3150 - 0xc4e  :    0 - 0x0
    "00000001", -- 3151 - 0xc4f  :    1 - 0x1
    "00000001", -- 3152 - 0xc50  :    1 - 0x1 -- Sprite 0xc5
    "00000001", -- 3153 - 0xc51  :    1 - 0x1
    "01000001", -- 3154 - 0xc52  :   65 - 0x41
    "00000001", -- 3155 - 0xc53  :    1 - 0x1
    "00000001", -- 3156 - 0xc54  :    1 - 0x1
    "00000000", -- 3157 - 0xc55  :    0 - 0x0
    "00011111", -- 3158 - 0xc56  :   31 - 0x1f
    "00111111", -- 3159 - 0xc57  :   63 - 0x3f
    "00001111", -- 3160 - 0xc58  :   15 - 0xf
    "01111001", -- 3161 - 0xc59  :  121 - 0x79
    "10100001", -- 3162 - 0xc5a  :  161 - 0xa1
    "01111001", -- 3163 - 0xc5b  :  121 - 0x79
    "00001111", -- 3164 - 0xc5c  :   15 - 0xf
    "00000001", -- 3165 - 0xc5d  :    1 - 0x1
    "00000000", -- 3166 - 0xc5e  :    0 - 0x0
    "00000000", -- 3167 - 0xc5f  :    0 - 0x0
    "00000000", -- 3168 - 0xc60  :    0 - 0x0 -- Sprite 0xc6
    "00000000", -- 3169 - 0xc61  :    0 - 0x0
    "00000000", -- 3170 - 0xc62  :    0 - 0x0
    "00000000", -- 3171 - 0xc63  :    0 - 0x0
    "00000000", -- 3172 - 0xc64  :    0 - 0x0
    "11111100", -- 3173 - 0xc65  :  252 - 0xfc
    "11111000", -- 3174 - 0xc66  :  248 - 0xf8
    "00000000", -- 3175 - 0xc67  :    0 - 0x0
    "00000000", -- 3176 - 0xc68  :    0 - 0x0
    "00000000", -- 3177 - 0xc69  :    0 - 0x0
    "00000000", -- 3178 - 0xc6a  :    0 - 0x0
    "00000000", -- 3179 - 0xc6b  :    0 - 0x0
    "00000000", -- 3180 - 0xc6c  :    0 - 0x0
    "00000000", -- 3181 - 0xc6d  :    0 - 0x0
    "00000000", -- 3182 - 0xc6e  :    0 - 0x0
    "10000000", -- 3183 - 0xc6f  :  128 - 0x80
    "10000000", -- 3184 - 0xc70  :  128 - 0x80 -- Sprite 0xc7
    "10000000", -- 3185 - 0xc71  :  128 - 0x80
    "10000010", -- 3186 - 0xc72  :  130 - 0x82
    "10000000", -- 3187 - 0xc73  :  128 - 0x80
    "10000000", -- 3188 - 0xc74  :  128 - 0x80
    "00000000", -- 3189 - 0xc75  :    0 - 0x0
    "11111000", -- 3190 - 0xc76  :  248 - 0xf8
    "11111100", -- 3191 - 0xc77  :  252 - 0xfc
    "11110000", -- 3192 - 0xc78  :  240 - 0xf0
    "10011110", -- 3193 - 0xc79  :  158 - 0x9e
    "10000101", -- 3194 - 0xc7a  :  133 - 0x85
    "10011110", -- 3195 - 0xc7b  :  158 - 0x9e
    "11110000", -- 3196 - 0xc7c  :  240 - 0xf0
    "10000000", -- 3197 - 0xc7d  :  128 - 0x80
    "00000000", -- 3198 - 0xc7e  :    0 - 0x0
    "00000000", -- 3199 - 0xc7f  :    0 - 0x0
    "00000000", -- 3200 - 0xc80  :    0 - 0x0 -- Sprite 0xc8
    "00000000", -- 3201 - 0xc81  :    0 - 0x0
    "00000000", -- 3202 - 0xc82  :    0 - 0x0
    "00011110", -- 3203 - 0xc83  :   30 - 0x1e
    "00111111", -- 3204 - 0xc84  :   63 - 0x3f
    "00111111", -- 3205 - 0xc85  :   63 - 0x3f
    "00111111", -- 3206 - 0xc86  :   63 - 0x3f
    "00111111", -- 3207 - 0xc87  :   63 - 0x3f
    "00000000", -- 3208 - 0xc88  :    0 - 0x0
    "00000000", -- 3209 - 0xc89  :    0 - 0x0
    "00000000", -- 3210 - 0xc8a  :    0 - 0x0
    "00011110", -- 3211 - 0xc8b  :   30 - 0x1e
    "00111111", -- 3212 - 0xc8c  :   63 - 0x3f
    "00111111", -- 3213 - 0xc8d  :   63 - 0x3f
    "00111111", -- 3214 - 0xc8e  :   63 - 0x3f
    "00111111", -- 3215 - 0xc8f  :   63 - 0x3f
    "00011111", -- 3216 - 0xc90  :   31 - 0x1f -- Sprite 0xc9
    "00001111", -- 3217 - 0xc91  :   15 - 0xf
    "00000111", -- 3218 - 0xc92  :    7 - 0x7
    "00000011", -- 3219 - 0xc93  :    3 - 0x3
    "00000001", -- 3220 - 0xc94  :    1 - 0x1
    "00000000", -- 3221 - 0xc95  :    0 - 0x0
    "00000000", -- 3222 - 0xc96  :    0 - 0x0
    "00000000", -- 3223 - 0xc97  :    0 - 0x0
    "00011111", -- 3224 - 0xc98  :   31 - 0x1f
    "00001111", -- 3225 - 0xc99  :   15 - 0xf
    "00000111", -- 3226 - 0xc9a  :    7 - 0x7
    "00000011", -- 3227 - 0xc9b  :    3 - 0x3
    "00000001", -- 3228 - 0xc9c  :    1 - 0x1
    "00000000", -- 3229 - 0xc9d  :    0 - 0x0
    "00000000", -- 3230 - 0xc9e  :    0 - 0x0
    "00000000", -- 3231 - 0xc9f  :    0 - 0x0
    "00000000", -- 3232 - 0xca0  :    0 - 0x0 -- Sprite 0xca
    "00000000", -- 3233 - 0xca1  :    0 - 0x0
    "00000000", -- 3234 - 0xca2  :    0 - 0x0
    "00111100", -- 3235 - 0xca3  :   60 - 0x3c
    "01111110", -- 3236 - 0xca4  :  126 - 0x7e
    "11111110", -- 3237 - 0xca5  :  254 - 0xfe
    "11111110", -- 3238 - 0xca6  :  254 - 0xfe
    "11111110", -- 3239 - 0xca7  :  254 - 0xfe
    "00000000", -- 3240 - 0xca8  :    0 - 0x0
    "00000000", -- 3241 - 0xca9  :    0 - 0x0
    "00000000", -- 3242 - 0xcaa  :    0 - 0x0
    "00111100", -- 3243 - 0xcab  :   60 - 0x3c
    "01111110", -- 3244 - 0xcac  :  126 - 0x7e
    "11111110", -- 3245 - 0xcad  :  254 - 0xfe
    "11111110", -- 3246 - 0xcae  :  254 - 0xfe
    "11111110", -- 3247 - 0xcaf  :  254 - 0xfe
    "11111100", -- 3248 - 0xcb0  :  252 - 0xfc -- Sprite 0xcb
    "11111000", -- 3249 - 0xcb1  :  248 - 0xf8
    "11110000", -- 3250 - 0xcb2  :  240 - 0xf0
    "11100000", -- 3251 - 0xcb3  :  224 - 0xe0
    "11000000", -- 3252 - 0xcb4  :  192 - 0xc0
    "10000000", -- 3253 - 0xcb5  :  128 - 0x80
    "00000000", -- 3254 - 0xcb6  :    0 - 0x0
    "00000000", -- 3255 - 0xcb7  :    0 - 0x0
    "11111100", -- 3256 - 0xcb8  :  252 - 0xfc
    "11111000", -- 3257 - 0xcb9  :  248 - 0xf8
    "11110000", -- 3258 - 0xcba  :  240 - 0xf0
    "11100000", -- 3259 - 0xcbb  :  224 - 0xe0
    "11000000", -- 3260 - 0xcbc  :  192 - 0xc0
    "10000000", -- 3261 - 0xcbd  :  128 - 0x80
    "00000000", -- 3262 - 0xcbe  :    0 - 0x0
    "00000000", -- 3263 - 0xcbf  :    0 - 0x0
    "11111111", -- 3264 - 0xcc0  :  255 - 0xff -- Sprite 0xcc
    "11111111", -- 3265 - 0xcc1  :  255 - 0xff
    "11111111", -- 3266 - 0xcc2  :  255 - 0xff
    "11111111", -- 3267 - 0xcc3  :  255 - 0xff
    "11111111", -- 3268 - 0xcc4  :  255 - 0xff
    "11111111", -- 3269 - 0xcc5  :  255 - 0xff
    "11111111", -- 3270 - 0xcc6  :  255 - 0xff
    "11111111", -- 3271 - 0xcc7  :  255 - 0xff
    "11111111", -- 3272 - 0xcc8  :  255 - 0xff
    "11111111", -- 3273 - 0xcc9  :  255 - 0xff
    "11111111", -- 3274 - 0xcca  :  255 - 0xff
    "11111111", -- 3275 - 0xccb  :  255 - 0xff
    "11111111", -- 3276 - 0xccc  :  255 - 0xff
    "11111111", -- 3277 - 0xccd  :  255 - 0xff
    "11111111", -- 3278 - 0xcce  :  255 - 0xff
    "11111111", -- 3279 - 0xccf  :  255 - 0xff
    "11111111", -- 3280 - 0xcd0  :  255 - 0xff -- Sprite 0xcd
    "11111111", -- 3281 - 0xcd1  :  255 - 0xff
    "11111111", -- 3282 - 0xcd2  :  255 - 0xff
    "11111111", -- 3283 - 0xcd3  :  255 - 0xff
    "11111111", -- 3284 - 0xcd4  :  255 - 0xff
    "11111111", -- 3285 - 0xcd5  :  255 - 0xff
    "11111111", -- 3286 - 0xcd6  :  255 - 0xff
    "11111111", -- 3287 - 0xcd7  :  255 - 0xff
    "11111111", -- 3288 - 0xcd8  :  255 - 0xff
    "11111111", -- 3289 - 0xcd9  :  255 - 0xff
    "11111111", -- 3290 - 0xcda  :  255 - 0xff
    "11111111", -- 3291 - 0xcdb  :  255 - 0xff
    "11111111", -- 3292 - 0xcdc  :  255 - 0xff
    "11111111", -- 3293 - 0xcdd  :  255 - 0xff
    "11111111", -- 3294 - 0xcde  :  255 - 0xff
    "11111111", -- 3295 - 0xcdf  :  255 - 0xff
    "11111111", -- 3296 - 0xce0  :  255 - 0xff -- Sprite 0xce
    "11111111", -- 3297 - 0xce1  :  255 - 0xff
    "11111111", -- 3298 - 0xce2  :  255 - 0xff
    "11111111", -- 3299 - 0xce3  :  255 - 0xff
    "11111111", -- 3300 - 0xce4  :  255 - 0xff
    "11111111", -- 3301 - 0xce5  :  255 - 0xff
    "11111111", -- 3302 - 0xce6  :  255 - 0xff
    "11111111", -- 3303 - 0xce7  :  255 - 0xff
    "11111111", -- 3304 - 0xce8  :  255 - 0xff
    "11111111", -- 3305 - 0xce9  :  255 - 0xff
    "11111111", -- 3306 - 0xcea  :  255 - 0xff
    "11111111", -- 3307 - 0xceb  :  255 - 0xff
    "11111111", -- 3308 - 0xcec  :  255 - 0xff
    "11111111", -- 3309 - 0xced  :  255 - 0xff
    "11111111", -- 3310 - 0xcee  :  255 - 0xff
    "11111111", -- 3311 - 0xcef  :  255 - 0xff
    "11111111", -- 3312 - 0xcf0  :  255 - 0xff -- Sprite 0xcf
    "11111111", -- 3313 - 0xcf1  :  255 - 0xff
    "11111111", -- 3314 - 0xcf2  :  255 - 0xff
    "11111111", -- 3315 - 0xcf3  :  255 - 0xff
    "11111111", -- 3316 - 0xcf4  :  255 - 0xff
    "11111111", -- 3317 - 0xcf5  :  255 - 0xff
    "11111111", -- 3318 - 0xcf6  :  255 - 0xff
    "11111111", -- 3319 - 0xcf7  :  255 - 0xff
    "11111111", -- 3320 - 0xcf8  :  255 - 0xff
    "11111111", -- 3321 - 0xcf9  :  255 - 0xff
    "11111111", -- 3322 - 0xcfa  :  255 - 0xff
    "11111111", -- 3323 - 0xcfb  :  255 - 0xff
    "11111111", -- 3324 - 0xcfc  :  255 - 0xff
    "11111111", -- 3325 - 0xcfd  :  255 - 0xff
    "11111111", -- 3326 - 0xcfe  :  255 - 0xff
    "11111111", -- 3327 - 0xcff  :  255 - 0xff
    "00001000", -- 3328 - 0xd00  :    8 - 0x8 -- Sprite 0xd0
    "00011001", -- 3329 - 0xd01  :   25 - 0x19
    "00001001", -- 3330 - 0xd02  :    9 - 0x9
    "00001001", -- 3331 - 0xd03  :    9 - 0x9
    "00001001", -- 3332 - 0xd04  :    9 - 0x9
    "00001001", -- 3333 - 0xd05  :    9 - 0x9
    "00011100", -- 3334 - 0xd06  :   28 - 0x1c
    "00000000", -- 3335 - 0xd07  :    0 - 0x0
    "00000000", -- 3336 - 0xd08  :    0 - 0x0
    "00000000", -- 3337 - 0xd09  :    0 - 0x0
    "00000000", -- 3338 - 0xd0a  :    0 - 0x0
    "00000000", -- 3339 - 0xd0b  :    0 - 0x0
    "00000000", -- 3340 - 0xd0c  :    0 - 0x0
    "00000000", -- 3341 - 0xd0d  :    0 - 0x0
    "00000000", -- 3342 - 0xd0e  :    0 - 0x0
    "00000000", -- 3343 - 0xd0f  :    0 - 0x0
    "00111000", -- 3344 - 0xd10  :   56 - 0x38 -- Sprite 0xd1
    "00000101", -- 3345 - 0xd11  :    5 - 0x5
    "00000101", -- 3346 - 0xd12  :    5 - 0x5
    "00011001", -- 3347 - 0xd13  :   25 - 0x19
    "00000101", -- 3348 - 0xd14  :    5 - 0x5
    "00000101", -- 3349 - 0xd15  :    5 - 0x5
    "00111000", -- 3350 - 0xd16  :   56 - 0x38
    "00000000", -- 3351 - 0xd17  :    0 - 0x0
    "00000000", -- 3352 - 0xd18  :    0 - 0x0
    "00000000", -- 3353 - 0xd19  :    0 - 0x0
    "00000000", -- 3354 - 0xd1a  :    0 - 0x0
    "00000000", -- 3355 - 0xd1b  :    0 - 0x0
    "00000000", -- 3356 - 0xd1c  :    0 - 0x0
    "00000000", -- 3357 - 0xd1d  :    0 - 0x0
    "00000000", -- 3358 - 0xd1e  :    0 - 0x0
    "00000000", -- 3359 - 0xd1f  :    0 - 0x0
    "00111100", -- 3360 - 0xd20  :   60 - 0x3c -- Sprite 0xd2
    "00100001", -- 3361 - 0xd21  :   33 - 0x21
    "00100001", -- 3362 - 0xd22  :   33 - 0x21
    "00111101", -- 3363 - 0xd23  :   61 - 0x3d
    "00000101", -- 3364 - 0xd24  :    5 - 0x5
    "00000101", -- 3365 - 0xd25  :    5 - 0x5
    "00111000", -- 3366 - 0xd26  :   56 - 0x38
    "00000000", -- 3367 - 0xd27  :    0 - 0x0
    "00000000", -- 3368 - 0xd28  :    0 - 0x0
    "00000000", -- 3369 - 0xd29  :    0 - 0x0
    "00000000", -- 3370 - 0xd2a  :    0 - 0x0
    "00000000", -- 3371 - 0xd2b  :    0 - 0x0
    "00000000", -- 3372 - 0xd2c  :    0 - 0x0
    "00000000", -- 3373 - 0xd2d  :    0 - 0x0
    "00000000", -- 3374 - 0xd2e  :    0 - 0x0
    "00000000", -- 3375 - 0xd2f  :    0 - 0x0
    "00011000", -- 3376 - 0xd30  :   24 - 0x18 -- Sprite 0xd3
    "00100101", -- 3377 - 0xd31  :   37 - 0x25
    "00100101", -- 3378 - 0xd32  :   37 - 0x25
    "00011001", -- 3379 - 0xd33  :   25 - 0x19
    "00100101", -- 3380 - 0xd34  :   37 - 0x25
    "00100101", -- 3381 - 0xd35  :   37 - 0x25
    "00011000", -- 3382 - 0xd36  :   24 - 0x18
    "00000000", -- 3383 - 0xd37  :    0 - 0x0
    "00000000", -- 3384 - 0xd38  :    0 - 0x0
    "00000000", -- 3385 - 0xd39  :    0 - 0x0
    "00000000", -- 3386 - 0xd3a  :    0 - 0x0
    "00000000", -- 3387 - 0xd3b  :    0 - 0x0
    "00000000", -- 3388 - 0xd3c  :    0 - 0x0
    "00000000", -- 3389 - 0xd3d  :    0 - 0x0
    "00000000", -- 3390 - 0xd3e  :    0 - 0x0
    "00000000", -- 3391 - 0xd3f  :    0 - 0x0
    "11000110", -- 3392 - 0xd40  :  198 - 0xc6 -- Sprite 0xd4
    "00101001", -- 3393 - 0xd41  :   41 - 0x29
    "00101001", -- 3394 - 0xd42  :   41 - 0x29
    "00101001", -- 3395 - 0xd43  :   41 - 0x29
    "00101001", -- 3396 - 0xd44  :   41 - 0x29
    "00101001", -- 3397 - 0xd45  :   41 - 0x29
    "11000110", -- 3398 - 0xd46  :  198 - 0xc6
    "00000000", -- 3399 - 0xd47  :    0 - 0x0
    "00000000", -- 3400 - 0xd48  :    0 - 0x0
    "00000000", -- 3401 - 0xd49  :    0 - 0x0
    "00000000", -- 3402 - 0xd4a  :    0 - 0x0
    "00000000", -- 3403 - 0xd4b  :    0 - 0x0
    "00000000", -- 3404 - 0xd4c  :    0 - 0x0
    "00000000", -- 3405 - 0xd4d  :    0 - 0x0
    "00000000", -- 3406 - 0xd4e  :    0 - 0x0
    "00000000", -- 3407 - 0xd4f  :    0 - 0x0
    "00000000", -- 3408 - 0xd50  :    0 - 0x0 -- Sprite 0xd5
    "00000000", -- 3409 - 0xd51  :    0 - 0x0
    "00000000", -- 3410 - 0xd52  :    0 - 0x0
    "00000000", -- 3411 - 0xd53  :    0 - 0x0
    "00000000", -- 3412 - 0xd54  :    0 - 0x0
    "00000000", -- 3413 - 0xd55  :    0 - 0x0
    "00000000", -- 3414 - 0xd56  :    0 - 0x0
    "00000000", -- 3415 - 0xd57  :    0 - 0x0
    "00000000", -- 3416 - 0xd58  :    0 - 0x0
    "00000000", -- 3417 - 0xd59  :    0 - 0x0
    "00000000", -- 3418 - 0xd5a  :    0 - 0x0
    "00000001", -- 3419 - 0xd5b  :    1 - 0x1
    "00000011", -- 3420 - 0xd5c  :    3 - 0x3
    "01100011", -- 3421 - 0xd5d  :   99 - 0x63
    "00110001", -- 3422 - 0xd5e  :   49 - 0x31
    "00011111", -- 3423 - 0xd5f  :   31 - 0x1f
    "00000000", -- 3424 - 0xd60  :    0 - 0x0 -- Sprite 0xd6
    "00000000", -- 3425 - 0xd61  :    0 - 0x0
    "00000000", -- 3426 - 0xd62  :    0 - 0x0
    "00000000", -- 3427 - 0xd63  :    0 - 0x0
    "00111100", -- 3428 - 0xd64  :   60 - 0x3c
    "10110110", -- 3429 - 0xd65  :  182 - 0xb6
    "01111100", -- 3430 - 0xd66  :  124 - 0x7c
    "11111000", -- 3431 - 0xd67  :  248 - 0xf8
    "00000000", -- 3432 - 0xd68  :    0 - 0x0
    "00000000", -- 3433 - 0xd69  :    0 - 0x0
    "11111100", -- 3434 - 0xd6a  :  252 - 0xfc
    "11111110", -- 3435 - 0xd6b  :  254 - 0xfe
    "11000000", -- 3436 - 0xd6c  :  192 - 0xc0
    "01000000", -- 3437 - 0xd6d  :   64 - 0x40
    "10000000", -- 3438 - 0xd6e  :  128 - 0x80
    "00000000", -- 3439 - 0xd6f  :    0 - 0x0
    "00000011", -- 3440 - 0xd70  :    3 - 0x3 -- Sprite 0xd7
    "00000011", -- 3441 - 0xd71  :    3 - 0x3
    "00000011", -- 3442 - 0xd72  :    3 - 0x3
    "00000111", -- 3443 - 0xd73  :    7 - 0x7
    "00001100", -- 3444 - 0xd74  :   12 - 0xc
    "00011011", -- 3445 - 0xd75  :   27 - 0x1b
    "01110111", -- 3446 - 0xd76  :  119 - 0x77
    "00000111", -- 3447 - 0xd77  :    7 - 0x7
    "01111111", -- 3448 - 0xd78  :  127 - 0x7f
    "00111111", -- 3449 - 0xd79  :   63 - 0x3f
    "01010011", -- 3450 - 0xd7a  :   83 - 0x53
    "00000111", -- 3451 - 0xd7b  :    7 - 0x7
    "00001100", -- 3452 - 0xd7c  :   12 - 0xc
    "00011011", -- 3453 - 0xd7d  :   27 - 0x1b
    "00000111", -- 3454 - 0xd7e  :    7 - 0x7
    "00000111", -- 3455 - 0xd7f  :    7 - 0x7
    "00001111", -- 3456 - 0xd80  :   15 - 0xf -- Sprite 0xd8
    "00001111", -- 3457 - 0xd81  :   15 - 0xf
    "00011111", -- 3458 - 0xd82  :   31 - 0x1f
    "00111111", -- 3459 - 0xd83  :   63 - 0x3f
    "01111111", -- 3460 - 0xd84  :  127 - 0x7f
    "00111111", -- 3461 - 0xd85  :   63 - 0x3f
    "00000000", -- 3462 - 0xd86  :    0 - 0x0
    "00000000", -- 3463 - 0xd87  :    0 - 0x0
    "00001111", -- 3464 - 0xd88  :   15 - 0xf
    "00001111", -- 3465 - 0xd89  :   15 - 0xf
    "00000011", -- 3466 - 0xd8a  :    3 - 0x3
    "00111000", -- 3467 - 0xd8b  :   56 - 0x38
    "00111111", -- 3468 - 0xd8c  :   63 - 0x3f
    "00001110", -- 3469 - 0xd8d  :   14 - 0xe
    "00011100", -- 3470 - 0xd8e  :   28 - 0x1c
    "00001110", -- 3471 - 0xd8f  :   14 - 0xe
    "11100000", -- 3472 - 0xd90  :  224 - 0xe0 -- Sprite 0xd9
    "11110000", -- 3473 - 0xd91  :  240 - 0xf0
    "11110000", -- 3474 - 0xd92  :  240 - 0xf0
    "11110000", -- 3475 - 0xd93  :  240 - 0xf0
    "00011000", -- 3476 - 0xd94  :   24 - 0x18
    "11111100", -- 3477 - 0xd95  :  252 - 0xfc
    "11111100", -- 3478 - 0xd96  :  252 - 0xfc
    "11111100", -- 3479 - 0xd97  :  252 - 0xfc
    "00000000", -- 3480 - 0xd98  :    0 - 0x0
    "10010000", -- 3481 - 0xd99  :  144 - 0x90
    "11110000", -- 3482 - 0xd9a  :  240 - 0xf0
    "11110000", -- 3483 - 0xd9b  :  240 - 0xf0
    "00011000", -- 3484 - 0xd9c  :   24 - 0x18
    "11111100", -- 3485 - 0xd9d  :  252 - 0xfc
    "11110000", -- 3486 - 0xd9e  :  240 - 0xf0
    "11111000", -- 3487 - 0xd9f  :  248 - 0xf8
    "11111000", -- 3488 - 0xda0  :  248 - 0xf8 -- Sprite 0xda
    "11111100", -- 3489 - 0xda1  :  252 - 0xfc
    "11111111", -- 3490 - 0xda2  :  255 - 0xff
    "11111111", -- 3491 - 0xda3  :  255 - 0xff
    "11111110", -- 3492 - 0xda4  :  254 - 0xfe
    "11110000", -- 3493 - 0xda5  :  240 - 0xf0
    "00000000", -- 3494 - 0xda6  :    0 - 0x0
    "00000000", -- 3495 - 0xda7  :    0 - 0x0
    "11111000", -- 3496 - 0xda8  :  248 - 0xf8
    "11110000", -- 3497 - 0xda9  :  240 - 0xf0
    "10000111", -- 3498 - 0xdaa  :  135 - 0x87
    "00111101", -- 3499 - 0xdab  :   61 - 0x3d
    "11111110", -- 3500 - 0xdac  :  254 - 0xfe
    "00011100", -- 3501 - 0xdad  :   28 - 0x1c
    "00001000", -- 3502 - 0xdae  :    8 - 0x8
    "00000000", -- 3503 - 0xdaf  :    0 - 0x0
    "00000011", -- 3504 - 0xdb0  :    3 - 0x3 -- Sprite 0xdb
    "00000011", -- 3505 - 0xdb1  :    3 - 0x3
    "00000011", -- 3506 - 0xdb2  :    3 - 0x3
    "00000011", -- 3507 - 0xdb3  :    3 - 0x3
    "00000001", -- 3508 - 0xdb4  :    1 - 0x1
    "00000000", -- 3509 - 0xdb5  :    0 - 0x0
    "00000111", -- 3510 - 0xdb6  :    7 - 0x7
    "00011111", -- 3511 - 0xdb7  :   31 - 0x1f
    "01111111", -- 3512 - 0xdb8  :  127 - 0x7f
    "00111111", -- 3513 - 0xdb9  :   63 - 0x3f
    "01010011", -- 3514 - 0xdba  :   83 - 0x53
    "00000011", -- 3515 - 0xdbb  :    3 - 0x3
    "00000001", -- 3516 - 0xdbc  :    1 - 0x1
    "00000000", -- 3517 - 0xdbd  :    0 - 0x0
    "00000111", -- 3518 - 0xdbe  :    7 - 0x7
    "00011111", -- 3519 - 0xdbf  :   31 - 0x1f
    "11111111", -- 3520 - 0xdc0  :  255 - 0xff -- Sprite 0xdc
    "11111111", -- 3521 - 0xdc1  :  255 - 0xff
    "01111111", -- 3522 - 0xdc2  :  127 - 0x7f
    "00111111", -- 3523 - 0xdc3  :   63 - 0x3f
    "00001111", -- 3524 - 0xdc4  :   15 - 0xf
    "00000011", -- 3525 - 0xdc5  :    3 - 0x3
    "00000000", -- 3526 - 0xdc6  :    0 - 0x0
    "00000000", -- 3527 - 0xdc7  :    0 - 0x0
    "11001111", -- 3528 - 0xdc8  :  207 - 0xcf
    "01100011", -- 3529 - 0xdc9  :   99 - 0x63
    "00111000", -- 3530 - 0xdca  :   56 - 0x38
    "00111110", -- 3531 - 0xdcb  :   62 - 0x3e
    "01111011", -- 3532 - 0xdcc  :  123 - 0x7b
    "00110000", -- 3533 - 0xdcd  :   48 - 0x30
    "00011000", -- 3534 - 0xdce  :   24 - 0x18
    "00000000", -- 3535 - 0xdcf  :    0 - 0x0
    "11100000", -- 3536 - 0xdd0  :  224 - 0xe0 -- Sprite 0xdd
    "11110000", -- 3537 - 0xdd1  :  240 - 0xf0
    "11110000", -- 3538 - 0xdd2  :  240 - 0xf0
    "11100000", -- 3539 - 0xdd3  :  224 - 0xe0
    "11111110", -- 3540 - 0xdd4  :  254 - 0xfe
    "00111100", -- 3541 - 0xdd5  :   60 - 0x3c
    "11110000", -- 3542 - 0xdd6  :  240 - 0xf0
    "11111100", -- 3543 - 0xdd7  :  252 - 0xfc
    "00000000", -- 3544 - 0xdd8  :    0 - 0x0
    "10010000", -- 3545 - 0xdd9  :  144 - 0x90
    "11110000", -- 3546 - 0xdda  :  240 - 0xf0
    "11100000", -- 3547 - 0xddb  :  224 - 0xe0
    "11111000", -- 3548 - 0xddc  :  248 - 0xf8
    "00111000", -- 3549 - 0xddd  :   56 - 0x38
    "11110000", -- 3550 - 0xdde  :  240 - 0xf0
    "11110000", -- 3551 - 0xddf  :  240 - 0xf0
    "11111100", -- 3552 - 0xde0  :  252 - 0xfc -- Sprite 0xde
    "11111000", -- 3553 - 0xde1  :  248 - 0xf8
    "11111000", -- 3554 - 0xde2  :  248 - 0xf8
    "11111000", -- 3555 - 0xde3  :  248 - 0xf8
    "11111000", -- 3556 - 0xde4  :  248 - 0xf8
    "11111000", -- 3557 - 0xde5  :  248 - 0xf8
    "11111000", -- 3558 - 0xde6  :  248 - 0xf8
    "00000000", -- 3559 - 0xde7  :    0 - 0x0
    "11111000", -- 3560 - 0xde8  :  248 - 0xf8
    "11111000", -- 3561 - 0xde9  :  248 - 0xf8
    "11111000", -- 3562 - 0xdea  :  248 - 0xf8
    "00111000", -- 3563 - 0xdeb  :   56 - 0x38
    "10000000", -- 3564 - 0xdec  :  128 - 0x80
    "11111000", -- 3565 - 0xded  :  248 - 0xf8
    "00000000", -- 3566 - 0xdee  :    0 - 0x0
    "01011100", -- 3567 - 0xdef  :   92 - 0x5c
    "11111111", -- 3568 - 0xdf0  :  255 - 0xff -- Sprite 0xdf
    "11111111", -- 3569 - 0xdf1  :  255 - 0xff
    "11111111", -- 3570 - 0xdf2  :  255 - 0xff
    "11111111", -- 3571 - 0xdf3  :  255 - 0xff
    "11111111", -- 3572 - 0xdf4  :  255 - 0xff
    "11111111", -- 3573 - 0xdf5  :  255 - 0xff
    "11111111", -- 3574 - 0xdf6  :  255 - 0xff
    "11111111", -- 3575 - 0xdf7  :  255 - 0xff
    "11111111", -- 3576 - 0xdf8  :  255 - 0xff
    "11111111", -- 3577 - 0xdf9  :  255 - 0xff
    "11111111", -- 3578 - 0xdfa  :  255 - 0xff
    "11111111", -- 3579 - 0xdfb  :  255 - 0xff
    "11111111", -- 3580 - 0xdfc  :  255 - 0xff
    "11111111", -- 3581 - 0xdfd  :  255 - 0xff
    "11111111", -- 3582 - 0xdfe  :  255 - 0xff
    "11111111", -- 3583 - 0xdff  :  255 - 0xff
    "11111111", -- 3584 - 0xe00  :  255 - 0xff -- Sprite 0xe0
    "11111111", -- 3585 - 0xe01  :  255 - 0xff
    "11111111", -- 3586 - 0xe02  :  255 - 0xff
    "11111111", -- 3587 - 0xe03  :  255 - 0xff
    "11111111", -- 3588 - 0xe04  :  255 - 0xff
    "11111111", -- 3589 - 0xe05  :  255 - 0xff
    "11111111", -- 3590 - 0xe06  :  255 - 0xff
    "11111111", -- 3591 - 0xe07  :  255 - 0xff
    "11111111", -- 3592 - 0xe08  :  255 - 0xff
    "11111111", -- 3593 - 0xe09  :  255 - 0xff
    "11111111", -- 3594 - 0xe0a  :  255 - 0xff
    "11111111", -- 3595 - 0xe0b  :  255 - 0xff
    "11111111", -- 3596 - 0xe0c  :  255 - 0xff
    "11111111", -- 3597 - 0xe0d  :  255 - 0xff
    "11111111", -- 3598 - 0xe0e  :  255 - 0xff
    "11111111", -- 3599 - 0xe0f  :  255 - 0xff
    "11111111", -- 3600 - 0xe10  :  255 - 0xff -- Sprite 0xe1
    "11111111", -- 3601 - 0xe11  :  255 - 0xff
    "11111111", -- 3602 - 0xe12  :  255 - 0xff
    "11111111", -- 3603 - 0xe13  :  255 - 0xff
    "11111111", -- 3604 - 0xe14  :  255 - 0xff
    "11111111", -- 3605 - 0xe15  :  255 - 0xff
    "11111111", -- 3606 - 0xe16  :  255 - 0xff
    "11111111", -- 3607 - 0xe17  :  255 - 0xff
    "11111111", -- 3608 - 0xe18  :  255 - 0xff
    "11111111", -- 3609 - 0xe19  :  255 - 0xff
    "11111111", -- 3610 - 0xe1a  :  255 - 0xff
    "11111111", -- 3611 - 0xe1b  :  255 - 0xff
    "11111111", -- 3612 - 0xe1c  :  255 - 0xff
    "11111111", -- 3613 - 0xe1d  :  255 - 0xff
    "11111111", -- 3614 - 0xe1e  :  255 - 0xff
    "11111111", -- 3615 - 0xe1f  :  255 - 0xff
    "11111111", -- 3616 - 0xe20  :  255 - 0xff -- Sprite 0xe2
    "11111111", -- 3617 - 0xe21  :  255 - 0xff
    "11111111", -- 3618 - 0xe22  :  255 - 0xff
    "11111111", -- 3619 - 0xe23  :  255 - 0xff
    "11111111", -- 3620 - 0xe24  :  255 - 0xff
    "11111111", -- 3621 - 0xe25  :  255 - 0xff
    "11111111", -- 3622 - 0xe26  :  255 - 0xff
    "11111111", -- 3623 - 0xe27  :  255 - 0xff
    "11111111", -- 3624 - 0xe28  :  255 - 0xff
    "11111111", -- 3625 - 0xe29  :  255 - 0xff
    "11111111", -- 3626 - 0xe2a  :  255 - 0xff
    "11111111", -- 3627 - 0xe2b  :  255 - 0xff
    "11111111", -- 3628 - 0xe2c  :  255 - 0xff
    "11111111", -- 3629 - 0xe2d  :  255 - 0xff
    "11111111", -- 3630 - 0xe2e  :  255 - 0xff
    "11111111", -- 3631 - 0xe2f  :  255 - 0xff
    "11111111", -- 3632 - 0xe30  :  255 - 0xff -- Sprite 0xe3
    "11111111", -- 3633 - 0xe31  :  255 - 0xff
    "11111111", -- 3634 - 0xe32  :  255 - 0xff
    "11111111", -- 3635 - 0xe33  :  255 - 0xff
    "11111111", -- 3636 - 0xe34  :  255 - 0xff
    "11111111", -- 3637 - 0xe35  :  255 - 0xff
    "11111111", -- 3638 - 0xe36  :  255 - 0xff
    "11111111", -- 3639 - 0xe37  :  255 - 0xff
    "11111111", -- 3640 - 0xe38  :  255 - 0xff
    "11111111", -- 3641 - 0xe39  :  255 - 0xff
    "11111111", -- 3642 - 0xe3a  :  255 - 0xff
    "11111111", -- 3643 - 0xe3b  :  255 - 0xff
    "11111111", -- 3644 - 0xe3c  :  255 - 0xff
    "11111111", -- 3645 - 0xe3d  :  255 - 0xff
    "11111111", -- 3646 - 0xe3e  :  255 - 0xff
    "11111111", -- 3647 - 0xe3f  :  255 - 0xff
    "11111111", -- 3648 - 0xe40  :  255 - 0xff -- Sprite 0xe4
    "11111111", -- 3649 - 0xe41  :  255 - 0xff
    "11111111", -- 3650 - 0xe42  :  255 - 0xff
    "11111111", -- 3651 - 0xe43  :  255 - 0xff
    "11111111", -- 3652 - 0xe44  :  255 - 0xff
    "11111111", -- 3653 - 0xe45  :  255 - 0xff
    "11111111", -- 3654 - 0xe46  :  255 - 0xff
    "11111111", -- 3655 - 0xe47  :  255 - 0xff
    "11111111", -- 3656 - 0xe48  :  255 - 0xff
    "11111111", -- 3657 - 0xe49  :  255 - 0xff
    "11111111", -- 3658 - 0xe4a  :  255 - 0xff
    "11111111", -- 3659 - 0xe4b  :  255 - 0xff
    "11111111", -- 3660 - 0xe4c  :  255 - 0xff
    "11111111", -- 3661 - 0xe4d  :  255 - 0xff
    "11111111", -- 3662 - 0xe4e  :  255 - 0xff
    "11111111", -- 3663 - 0xe4f  :  255 - 0xff
    "11111111", -- 3664 - 0xe50  :  255 - 0xff -- Sprite 0xe5
    "11111111", -- 3665 - 0xe51  :  255 - 0xff
    "11111111", -- 3666 - 0xe52  :  255 - 0xff
    "11111111", -- 3667 - 0xe53  :  255 - 0xff
    "11111111", -- 3668 - 0xe54  :  255 - 0xff
    "11111111", -- 3669 - 0xe55  :  255 - 0xff
    "11111111", -- 3670 - 0xe56  :  255 - 0xff
    "11111111", -- 3671 - 0xe57  :  255 - 0xff
    "11111111", -- 3672 - 0xe58  :  255 - 0xff
    "11111111", -- 3673 - 0xe59  :  255 - 0xff
    "11111111", -- 3674 - 0xe5a  :  255 - 0xff
    "11111111", -- 3675 - 0xe5b  :  255 - 0xff
    "11111111", -- 3676 - 0xe5c  :  255 - 0xff
    "11111111", -- 3677 - 0xe5d  :  255 - 0xff
    "11111111", -- 3678 - 0xe5e  :  255 - 0xff
    "11111111", -- 3679 - 0xe5f  :  255 - 0xff
    "11111111", -- 3680 - 0xe60  :  255 - 0xff -- Sprite 0xe6
    "11111111", -- 3681 - 0xe61  :  255 - 0xff
    "11111111", -- 3682 - 0xe62  :  255 - 0xff
    "11111111", -- 3683 - 0xe63  :  255 - 0xff
    "11111111", -- 3684 - 0xe64  :  255 - 0xff
    "11111111", -- 3685 - 0xe65  :  255 - 0xff
    "11111111", -- 3686 - 0xe66  :  255 - 0xff
    "11111111", -- 3687 - 0xe67  :  255 - 0xff
    "11111111", -- 3688 - 0xe68  :  255 - 0xff
    "11111111", -- 3689 - 0xe69  :  255 - 0xff
    "11111111", -- 3690 - 0xe6a  :  255 - 0xff
    "11111111", -- 3691 - 0xe6b  :  255 - 0xff
    "11111111", -- 3692 - 0xe6c  :  255 - 0xff
    "11111111", -- 3693 - 0xe6d  :  255 - 0xff
    "11111111", -- 3694 - 0xe6e  :  255 - 0xff
    "11111111", -- 3695 - 0xe6f  :  255 - 0xff
    "11111111", -- 3696 - 0xe70  :  255 - 0xff -- Sprite 0xe7
    "11111111", -- 3697 - 0xe71  :  255 - 0xff
    "11111111", -- 3698 - 0xe72  :  255 - 0xff
    "11111111", -- 3699 - 0xe73  :  255 - 0xff
    "11111111", -- 3700 - 0xe74  :  255 - 0xff
    "11111111", -- 3701 - 0xe75  :  255 - 0xff
    "11111111", -- 3702 - 0xe76  :  255 - 0xff
    "11111111", -- 3703 - 0xe77  :  255 - 0xff
    "11111111", -- 3704 - 0xe78  :  255 - 0xff
    "11111111", -- 3705 - 0xe79  :  255 - 0xff
    "11111111", -- 3706 - 0xe7a  :  255 - 0xff
    "11111111", -- 3707 - 0xe7b  :  255 - 0xff
    "11111111", -- 3708 - 0xe7c  :  255 - 0xff
    "11111111", -- 3709 - 0xe7d  :  255 - 0xff
    "11111111", -- 3710 - 0xe7e  :  255 - 0xff
    "11111111", -- 3711 - 0xe7f  :  255 - 0xff
    "11111111", -- 3712 - 0xe80  :  255 - 0xff -- Sprite 0xe8
    "11111111", -- 3713 - 0xe81  :  255 - 0xff
    "11111111", -- 3714 - 0xe82  :  255 - 0xff
    "11111111", -- 3715 - 0xe83  :  255 - 0xff
    "11111111", -- 3716 - 0xe84  :  255 - 0xff
    "11111111", -- 3717 - 0xe85  :  255 - 0xff
    "11111111", -- 3718 - 0xe86  :  255 - 0xff
    "11111111", -- 3719 - 0xe87  :  255 - 0xff
    "11111111", -- 3720 - 0xe88  :  255 - 0xff
    "11111111", -- 3721 - 0xe89  :  255 - 0xff
    "11111111", -- 3722 - 0xe8a  :  255 - 0xff
    "11111111", -- 3723 - 0xe8b  :  255 - 0xff
    "11111111", -- 3724 - 0xe8c  :  255 - 0xff
    "11111111", -- 3725 - 0xe8d  :  255 - 0xff
    "11111111", -- 3726 - 0xe8e  :  255 - 0xff
    "11111111", -- 3727 - 0xe8f  :  255 - 0xff
    "11111111", -- 3728 - 0xe90  :  255 - 0xff -- Sprite 0xe9
    "11111111", -- 3729 - 0xe91  :  255 - 0xff
    "11111111", -- 3730 - 0xe92  :  255 - 0xff
    "11111111", -- 3731 - 0xe93  :  255 - 0xff
    "11111111", -- 3732 - 0xe94  :  255 - 0xff
    "11111111", -- 3733 - 0xe95  :  255 - 0xff
    "11111111", -- 3734 - 0xe96  :  255 - 0xff
    "11111111", -- 3735 - 0xe97  :  255 - 0xff
    "11111111", -- 3736 - 0xe98  :  255 - 0xff
    "11111111", -- 3737 - 0xe99  :  255 - 0xff
    "11111111", -- 3738 - 0xe9a  :  255 - 0xff
    "11111111", -- 3739 - 0xe9b  :  255 - 0xff
    "11111111", -- 3740 - 0xe9c  :  255 - 0xff
    "11111111", -- 3741 - 0xe9d  :  255 - 0xff
    "11111111", -- 3742 - 0xe9e  :  255 - 0xff
    "11111111", -- 3743 - 0xe9f  :  255 - 0xff
    "11111111", -- 3744 - 0xea0  :  255 - 0xff -- Sprite 0xea
    "11111111", -- 3745 - 0xea1  :  255 - 0xff
    "11111111", -- 3746 - 0xea2  :  255 - 0xff
    "11111111", -- 3747 - 0xea3  :  255 - 0xff
    "11111111", -- 3748 - 0xea4  :  255 - 0xff
    "11111111", -- 3749 - 0xea5  :  255 - 0xff
    "11111111", -- 3750 - 0xea6  :  255 - 0xff
    "11111111", -- 3751 - 0xea7  :  255 - 0xff
    "11111111", -- 3752 - 0xea8  :  255 - 0xff
    "11111111", -- 3753 - 0xea9  :  255 - 0xff
    "11111111", -- 3754 - 0xeaa  :  255 - 0xff
    "11111111", -- 3755 - 0xeab  :  255 - 0xff
    "11111111", -- 3756 - 0xeac  :  255 - 0xff
    "11111111", -- 3757 - 0xead  :  255 - 0xff
    "11111111", -- 3758 - 0xeae  :  255 - 0xff
    "11111111", -- 3759 - 0xeaf  :  255 - 0xff
    "11111111", -- 3760 - 0xeb0  :  255 - 0xff -- Sprite 0xeb
    "11111111", -- 3761 - 0xeb1  :  255 - 0xff
    "11111111", -- 3762 - 0xeb2  :  255 - 0xff
    "11111111", -- 3763 - 0xeb3  :  255 - 0xff
    "11111111", -- 3764 - 0xeb4  :  255 - 0xff
    "11111111", -- 3765 - 0xeb5  :  255 - 0xff
    "11111111", -- 3766 - 0xeb6  :  255 - 0xff
    "11111111", -- 3767 - 0xeb7  :  255 - 0xff
    "11111111", -- 3768 - 0xeb8  :  255 - 0xff
    "11111111", -- 3769 - 0xeb9  :  255 - 0xff
    "11111111", -- 3770 - 0xeba  :  255 - 0xff
    "11111111", -- 3771 - 0xebb  :  255 - 0xff
    "11111111", -- 3772 - 0xebc  :  255 - 0xff
    "11111111", -- 3773 - 0xebd  :  255 - 0xff
    "11111111", -- 3774 - 0xebe  :  255 - 0xff
    "11111111", -- 3775 - 0xebf  :  255 - 0xff
    "00000000", -- 3776 - 0xec0  :    0 - 0x0 -- Sprite 0xec
    "00000001", -- 3777 - 0xec1  :    1 - 0x1
    "00000011", -- 3778 - 0xec2  :    3 - 0x3
    "00110011", -- 3779 - 0xec3  :   51 - 0x33
    "00011001", -- 3780 - 0xec4  :   25 - 0x19
    "00001111", -- 3781 - 0xec5  :   15 - 0xf
    "00111111", -- 3782 - 0xec6  :   63 - 0x3f
    "00011111", -- 3783 - 0xec7  :   31 - 0x1f
    "00000000", -- 3784 - 0xec8  :    0 - 0x0
    "00000001", -- 3785 - 0xec9  :    1 - 0x1
    "00000011", -- 3786 - 0xeca  :    3 - 0x3
    "00110011", -- 3787 - 0xecb  :   51 - 0x33
    "00011001", -- 3788 - 0xecc  :   25 - 0x19
    "00001111", -- 3789 - 0xecd  :   15 - 0xf
    "00111111", -- 3790 - 0xece  :   63 - 0x3f
    "00011111", -- 3791 - 0xecf  :   31 - 0x1f
    "00101011", -- 3792 - 0xed0  :   43 - 0x2b -- Sprite 0xed
    "00000111", -- 3793 - 0xed1  :    7 - 0x7
    "00000101", -- 3794 - 0xed2  :    5 - 0x5
    "00001101", -- 3795 - 0xed3  :   13 - 0xd
    "00001011", -- 3796 - 0xed4  :   11 - 0xb
    "00011011", -- 3797 - 0xed5  :   27 - 0x1b
    "00011011", -- 3798 - 0xed6  :   27 - 0x1b
    "00111011", -- 3799 - 0xed7  :   59 - 0x3b
    "00101011", -- 3800 - 0xed8  :   43 - 0x2b
    "00000111", -- 3801 - 0xed9  :    7 - 0x7
    "00000101", -- 3802 - 0xeda  :    5 - 0x5
    "00001101", -- 3803 - 0xedb  :   13 - 0xd
    "00001011", -- 3804 - 0xedc  :   11 - 0xb
    "00011011", -- 3805 - 0xedd  :   27 - 0x1b
    "00011011", -- 3806 - 0xede  :   27 - 0x1b
    "00000011", -- 3807 - 0xedf  :    3 - 0x3
    "00001001", -- 3808 - 0xee0  :    9 - 0x9 -- Sprite 0xee
    "00000000", -- 3809 - 0xee1  :    0 - 0x0
    "00000111", -- 3810 - 0xee2  :    7 - 0x7
    "00000111", -- 3811 - 0xee3  :    7 - 0x7
    "00001111", -- 3812 - 0xee4  :   15 - 0xf
    "00001101", -- 3813 - 0xee5  :   13 - 0xd
    "00000001", -- 3814 - 0xee6  :    1 - 0x1
    "00000000", -- 3815 - 0xee7  :    0 - 0x0
    "00000001", -- 3816 - 0xee8  :    1 - 0x1
    "00000000", -- 3817 - 0xee9  :    0 - 0x0
    "00000011", -- 3818 - 0xeea  :    3 - 0x3
    "00000101", -- 3819 - 0xeeb  :    5 - 0x5
    "00001110", -- 3820 - 0xeec  :   14 - 0xe
    "00001101", -- 3821 - 0xeed  :   13 - 0xd
    "00000001", -- 3822 - 0xeee  :    1 - 0x1
    "00000000", -- 3823 - 0xeef  :    0 - 0x0
    "11111000", -- 3824 - 0xef0  :  248 - 0xf8 -- Sprite 0xef
    "11111100", -- 3825 - 0xef1  :  252 - 0xfc
    "11111000", -- 3826 - 0xef2  :  248 - 0xf8
    "11101100", -- 3827 - 0xef3  :  236 - 0xec
    "11111000", -- 3828 - 0xef4  :  248 - 0xf8
    "11110000", -- 3829 - 0xef5  :  240 - 0xf0
    "11000000", -- 3830 - 0xef6  :  192 - 0xc0
    "11000000", -- 3831 - 0xef7  :  192 - 0xc0
    "11111000", -- 3832 - 0xef8  :  248 - 0xf8
    "11111100", -- 3833 - 0xef9  :  252 - 0xfc
    "11000000", -- 3834 - 0xefa  :  192 - 0xc0
    "01000000", -- 3835 - 0xefb  :   64 - 0x40
    "10000000", -- 3836 - 0xefc  :  128 - 0x80
    "10000000", -- 3837 - 0xefd  :  128 - 0x80
    "00000000", -- 3838 - 0xefe  :    0 - 0x0
    "10000000", -- 3839 - 0xeff  :  128 - 0x80
    "11110000", -- 3840 - 0xf00  :  240 - 0xf0 -- Sprite 0xf0
    "11111000", -- 3841 - 0xf01  :  248 - 0xf8
    "11111000", -- 3842 - 0xf02  :  248 - 0xf8
    "11101000", -- 3843 - 0xf03  :  232 - 0xe8
    "11001100", -- 3844 - 0xf04  :  204 - 0xcc
    "11100110", -- 3845 - 0xf05  :  230 - 0xe6
    "11111011", -- 3846 - 0xf06  :  251 - 0xfb
    "11111111", -- 3847 - 0xf07  :  255 - 0xff
    "11010000", -- 3848 - 0xf08  :  208 - 0xd0
    "11111000", -- 3849 - 0xf09  :  248 - 0xf8
    "11111000", -- 3850 - 0xf0a  :  248 - 0xf8
    "11101000", -- 3851 - 0xf0b  :  232 - 0xe8
    "11001100", -- 3852 - 0xf0c  :  204 - 0xcc
    "11100110", -- 3853 - 0xf0d  :  230 - 0xe6
    "11111000", -- 3854 - 0xf0e  :  248 - 0xf8
    "11111110", -- 3855 - 0xf0f  :  254 - 0xfe
    "11111111", -- 3856 - 0xf10  :  255 - 0xff -- Sprite 0xf1
    "11111110", -- 3857 - 0xf11  :  254 - 0xfe
    "11111110", -- 3858 - 0xf12  :  254 - 0xfe
    "11111110", -- 3859 - 0xf13  :  254 - 0xfe
    "11111110", -- 3860 - 0xf14  :  254 - 0xfe
    "10001111", -- 3861 - 0xf15  :  143 - 0x8f
    "00000000", -- 3862 - 0xf16  :    0 - 0x0
    "00000000", -- 3863 - 0xf17  :    0 - 0x0
    "11111110", -- 3864 - 0xf18  :  254 - 0xfe
    "11111110", -- 3865 - 0xf19  :  254 - 0xfe
    "00000110", -- 3866 - 0xf1a  :    6 - 0x6
    "11111000", -- 3867 - 0xf1b  :  248 - 0xf8
    "00001110", -- 3868 - 0xf1c  :   14 - 0xe
    "10000000", -- 3869 - 0xf1d  :  128 - 0x80
    "00000000", -- 3870 - 0xf1e  :    0 - 0x0
    "00000000", -- 3871 - 0xf1f  :    0 - 0x0
    "00000001", -- 3872 - 0xf20  :    1 - 0x1 -- Sprite 0xf2
    "00001111", -- 3873 - 0xf21  :   15 - 0xf
    "00000000", -- 3874 - 0xf22  :    0 - 0x0
    "00000000", -- 3875 - 0xf23  :    0 - 0x0
    "00000100", -- 3876 - 0xf24  :    4 - 0x4
    "00011110", -- 3877 - 0xf25  :   30 - 0x1e
    "00000000", -- 3878 - 0xf26  :    0 - 0x0
    "00000011", -- 3879 - 0xf27  :    3 - 0x3
    "00000001", -- 3880 - 0xf28  :    1 - 0x1
    "00001111", -- 3881 - 0xf29  :   15 - 0xf
    "00000111", -- 3882 - 0xf2a  :    7 - 0x7
    "00011101", -- 3883 - 0xf2b  :   29 - 0x1d
    "00111011", -- 3884 - 0xf2c  :   59 - 0x3b
    "00000001", -- 3885 - 0xf2d  :    1 - 0x1
    "00001111", -- 3886 - 0xf2e  :   15 - 0xf
    "00000010", -- 3887 - 0xf2f  :    2 - 0x2
    "00000111", -- 3888 - 0xf30  :    7 - 0x7 -- Sprite 0xf3
    "00001111", -- 3889 - 0xf31  :   15 - 0xf
    "00011111", -- 3890 - 0xf32  :   31 - 0x1f
    "00001111", -- 3891 - 0xf33  :   15 - 0xf
    "00000111", -- 3892 - 0xf34  :    7 - 0x7
    "00001111", -- 3893 - 0xf35  :   15 - 0xf
    "00001111", -- 3894 - 0xf36  :   15 - 0xf
    "00000011", -- 3895 - 0xf37  :    3 - 0x3
    "00000010", -- 3896 - 0xf38  :    2 - 0x2
    "00000011", -- 3897 - 0xf39  :    3 - 0x3
    "00000010", -- 3898 - 0xf3a  :    2 - 0x2
    "01110111", -- 3899 - 0xf3b  :  119 - 0x77
    "00010111", -- 3900 - 0xf3c  :   23 - 0x17
    "00000001", -- 3901 - 0xf3d  :    1 - 0x1
    "00000000", -- 3902 - 0xf3e  :    0 - 0x0
    "00000000", -- 3903 - 0xf3f  :    0 - 0x0
    "11100000", -- 3904 - 0xf40  :  224 - 0xe0 -- Sprite 0xf4
    "11110000", -- 3905 - 0xf41  :  240 - 0xf0
    "11110000", -- 3906 - 0xf42  :  240 - 0xf0
    "01001000", -- 3907 - 0xf43  :   72 - 0x48
    "11001000", -- 3908 - 0xf44  :  200 - 0xc8
    "10011100", -- 3909 - 0xf45  :  156 - 0x9c
    "00000000", -- 3910 - 0xf46  :    0 - 0x0
    "11110000", -- 3911 - 0xf47  :  240 - 0xf0
    "11100000", -- 3912 - 0xf48  :  224 - 0xe0
    "11110000", -- 3913 - 0xf49  :  240 - 0xf0
    "00000000", -- 3914 - 0xf4a  :    0 - 0x0
    "10110000", -- 3915 - 0xf4b  :  176 - 0xb0
    "00110000", -- 3916 - 0xf4c  :   48 - 0x30
    "01100000", -- 3917 - 0xf4d  :   96 - 0x60
    "11110000", -- 3918 - 0xf4e  :  240 - 0xf0
    "00010000", -- 3919 - 0xf4f  :   16 - 0x10
    "11111000", -- 3920 - 0xf50  :  248 - 0xf8 -- Sprite 0xf5
    "11111100", -- 3921 - 0xf51  :  252 - 0xfc
    "11111100", -- 3922 - 0xf52  :  252 - 0xfc
    "11111000", -- 3923 - 0xf53  :  248 - 0xf8
    "11111000", -- 3924 - 0xf54  :  248 - 0xf8
    "01111000", -- 3925 - 0xf55  :  120 - 0x78
    "01110000", -- 3926 - 0xf56  :  112 - 0x70
    "01100000", -- 3927 - 0xf57  :   96 - 0x60
    "00110000", -- 3928 - 0xf58  :   48 - 0x30
    "11110000", -- 3929 - 0xf59  :  240 - 0xf0
    "11010000", -- 3930 - 0xf5a  :  208 - 0xd0
    "11111100", -- 3931 - 0xf5b  :  252 - 0xfc
    "11111110", -- 3932 - 0xf5c  :  254 - 0xfe
    "00001000", -- 3933 - 0xf5d  :    8 - 0x8
    "00000000", -- 3934 - 0xf5e  :    0 - 0x0
    "00000000", -- 3935 - 0xf5f  :    0 - 0x0
    "00000000", -- 3936 - 0xf60  :    0 - 0x0 -- Sprite 0xf6
    "00000000", -- 3937 - 0xf61  :    0 - 0x0
    "01111100", -- 3938 - 0xf62  :  124 - 0x7c
    "10001010", -- 3939 - 0xf63  :  138 - 0x8a
    "11111110", -- 3940 - 0xf64  :  254 - 0xfe
    "11111110", -- 3941 - 0xf65  :  254 - 0xfe
    "11111110", -- 3942 - 0xf66  :  254 - 0xfe
    "11111110", -- 3943 - 0xf67  :  254 - 0xfe
    "00000000", -- 3944 - 0xf68  :    0 - 0x0
    "00010000", -- 3945 - 0xf69  :   16 - 0x10
    "00000000", -- 3946 - 0xf6a  :    0 - 0x0
    "01110100", -- 3947 - 0xf6b  :  116 - 0x74
    "00000000", -- 3948 - 0xf6c  :    0 - 0x0
    "00000000", -- 3949 - 0xf6d  :    0 - 0x0
    "00000000", -- 3950 - 0xf6e  :    0 - 0x0
    "00000000", -- 3951 - 0xf6f  :    0 - 0x0
    "11111110", -- 3952 - 0xf70  :  254 - 0xfe -- Sprite 0xf7
    "01111100", -- 3953 - 0xf71  :  124 - 0x7c
    "00000000", -- 3954 - 0xf72  :    0 - 0x0
    "00000000", -- 3955 - 0xf73  :    0 - 0x0
    "00000000", -- 3956 - 0xf74  :    0 - 0x0
    "00000000", -- 3957 - 0xf75  :    0 - 0x0
    "00000000", -- 3958 - 0xf76  :    0 - 0x0
    "00000000", -- 3959 - 0xf77  :    0 - 0x0
    "00000000", -- 3960 - 0xf78  :    0 - 0x0
    "00000000", -- 3961 - 0xf79  :    0 - 0x0
    "00010000", -- 3962 - 0xf7a  :   16 - 0x10
    "00010000", -- 3963 - 0xf7b  :   16 - 0x10
    "00010000", -- 3964 - 0xf7c  :   16 - 0x10
    "00010000", -- 3965 - 0xf7d  :   16 - 0x10
    "00010000", -- 3966 - 0xf7e  :   16 - 0x10
    "00010000", -- 3967 - 0xf7f  :   16 - 0x10
    "00000111", -- 3968 - 0xf80  :    7 - 0x7 -- Sprite 0xf8
    "00001011", -- 3969 - 0xf81  :   11 - 0xb
    "00001111", -- 3970 - 0xf82  :   15 - 0xf
    "00001011", -- 3971 - 0xf83  :   11 - 0xb
    "00001011", -- 3972 - 0xf84  :   11 - 0xb
    "00001011", -- 3973 - 0xf85  :   11 - 0xb
    "00001011", -- 3974 - 0xf86  :   11 - 0xb
    "00000111", -- 3975 - 0xf87  :    7 - 0x7
    "00000000", -- 3976 - 0xf88  :    0 - 0x0
    "00000100", -- 3977 - 0xf89  :    4 - 0x4
    "00000000", -- 3978 - 0xf8a  :    0 - 0x0
    "00010100", -- 3979 - 0xf8b  :   20 - 0x14
    "00000100", -- 3980 - 0xf8c  :    4 - 0x4
    "00000100", -- 3981 - 0xf8d  :    4 - 0x4
    "00000100", -- 3982 - 0xf8e  :    4 - 0x4
    "00000000", -- 3983 - 0xf8f  :    0 - 0x0
    "11000000", -- 3984 - 0xf90  :  192 - 0xc0 -- Sprite 0xf9
    "11100000", -- 3985 - 0xf91  :  224 - 0xe0
    "11100000", -- 3986 - 0xf92  :  224 - 0xe0
    "11100000", -- 3987 - 0xf93  :  224 - 0xe0
    "11100000", -- 3988 - 0xf94  :  224 - 0xe0
    "11100000", -- 3989 - 0xf95  :  224 - 0xe0
    "11100000", -- 3990 - 0xf96  :  224 - 0xe0
    "11000000", -- 3991 - 0xf97  :  192 - 0xc0
    "00000000", -- 3992 - 0xf98  :    0 - 0x0
    "00000000", -- 3993 - 0xf99  :    0 - 0x0
    "00000000", -- 3994 - 0xf9a  :    0 - 0x0
    "00011111", -- 3995 - 0xf9b  :   31 - 0x1f
    "00000000", -- 3996 - 0xf9c  :    0 - 0x0
    "00000000", -- 3997 - 0xf9d  :    0 - 0x0
    "00000000", -- 3998 - 0xf9e  :    0 - 0x0
    "00000000", -- 3999 - 0xf9f  :    0 - 0x0
    "00000011", -- 4000 - 0xfa0  :    3 - 0x3 -- Sprite 0xfa
    "00000111", -- 4001 - 0xfa1  :    7 - 0x7
    "00000111", -- 4002 - 0xfa2  :    7 - 0x7
    "00000111", -- 4003 - 0xfa3  :    7 - 0x7
    "00000111", -- 4004 - 0xfa4  :    7 - 0x7
    "00000111", -- 4005 - 0xfa5  :    7 - 0x7
    "00000111", -- 4006 - 0xfa6  :    7 - 0x7
    "00000011", -- 4007 - 0xfa7  :    3 - 0x3
    "00000000", -- 4008 - 0xfa8  :    0 - 0x0
    "00000000", -- 4009 - 0xfa9  :    0 - 0x0
    "00000000", -- 4010 - 0xfaa  :    0 - 0x0
    "11111000", -- 4011 - 0xfab  :  248 - 0xf8
    "00000000", -- 4012 - 0xfac  :    0 - 0x0
    "00000000", -- 4013 - 0xfad  :    0 - 0x0
    "00000000", -- 4014 - 0xfae  :    0 - 0x0
    "00000000", -- 4015 - 0xfaf  :    0 - 0x0
    "11100000", -- 4016 - 0xfb0  :  224 - 0xe0 -- Sprite 0xfb
    "11010000", -- 4017 - 0xfb1  :  208 - 0xd0
    "11010000", -- 4018 - 0xfb2  :  208 - 0xd0
    "11010000", -- 4019 - 0xfb3  :  208 - 0xd0
    "11010000", -- 4020 - 0xfb4  :  208 - 0xd0
    "11110000", -- 4021 - 0xfb5  :  240 - 0xf0
    "11010000", -- 4022 - 0xfb6  :  208 - 0xd0
    "11100000", -- 4023 - 0xfb7  :  224 - 0xe0
    "00000000", -- 4024 - 0xfb8  :    0 - 0x0
    "00100000", -- 4025 - 0xfb9  :   32 - 0x20
    "00100000", -- 4026 - 0xfba  :   32 - 0x20
    "00101000", -- 4027 - 0xfbb  :   40 - 0x28
    "00100000", -- 4028 - 0xfbc  :   32 - 0x20
    "00000000", -- 4029 - 0xfbd  :    0 - 0x0
    "00100000", -- 4030 - 0xfbe  :   32 - 0x20
    "00000000", -- 4031 - 0xfbf  :    0 - 0x0
    "00000000", -- 4032 - 0xfc0  :    0 - 0x0 -- Sprite 0xfc
    "00000001", -- 4033 - 0xfc1  :    1 - 0x1
    "00010011", -- 4034 - 0xfc2  :   19 - 0x13
    "00110111", -- 4035 - 0xfc3  :   55 - 0x37
    "00111011", -- 4036 - 0xfc4  :   59 - 0x3b
    "01110100", -- 4037 - 0xfc5  :  116 - 0x74
    "01111010", -- 4038 - 0xfc6  :  122 - 0x7a
    "00111110", -- 4039 - 0xfc7  :   62 - 0x3e
    "00000000", -- 4040 - 0xfc8  :    0 - 0x0
    "00000000", -- 4041 - 0xfc9  :    0 - 0x0
    "00001000", -- 4042 - 0xfca  :    8 - 0x8
    "00100101", -- 4043 - 0xfcb  :   37 - 0x25
    "00010010", -- 4044 - 0xfcc  :   18 - 0x12
    "01010011", -- 4045 - 0xfcd  :   83 - 0x53
    "00110011", -- 4046 - 0xfce  :   51 - 0x33
    "00111001", -- 4047 - 0xfcf  :   57 - 0x39
    "11011000", -- 4048 - 0xfd0  :  216 - 0xd8 -- Sprite 0xfd
    "10011000", -- 4049 - 0xfd1  :  152 - 0x98
    "10101000", -- 4050 - 0xfd2  :  168 - 0xa8
    "11011000", -- 4051 - 0xfd3  :  216 - 0xd8
    "11011010", -- 4052 - 0xfd4  :  218 - 0xda
    "01110100", -- 4053 - 0xfd5  :  116 - 0x74
    "00101000", -- 4054 - 0xfd6  :   40 - 0x28
    "11001000", -- 4055 - 0xfd7  :  200 - 0xc8
    "00001000", -- 4056 - 0xfd8  :    8 - 0x8
    "10000000", -- 4057 - 0xfd9  :  128 - 0x80
    "00110000", -- 4058 - 0xfda  :   48 - 0x30
    "10011100", -- 4059 - 0xfdb  :  156 - 0x9c
    "11001010", -- 4060 - 0xfdc  :  202 - 0xca
    "10111000", -- 4061 - 0xfdd  :  184 - 0xb8
    "10011000", -- 4062 - 0xfde  :  152 - 0x98
    "01111000", -- 4063 - 0xfdf  :  120 - 0x78
    "00001000", -- 4064 - 0xfe0  :    8 - 0x8 -- Sprite 0xfe
    "01011001", -- 4065 - 0xfe1  :   89 - 0x59
    "00110000", -- 4066 - 0xfe2  :   48 - 0x30
    "01110001", -- 4067 - 0xfe3  :  113 - 0x71
    "01111001", -- 4068 - 0xfe4  :  121 - 0x79
    "00101011", -- 4069 - 0xfe5  :   43 - 0x2b
    "00110110", -- 4070 - 0xfe6  :   54 - 0x36
    "00010110", -- 4071 - 0xfe7  :   22 - 0x16
    "00000000", -- 4072 - 0xfe8  :    0 - 0x0
    "00001000", -- 4073 - 0xfe9  :    8 - 0x8
    "00000000", -- 4074 - 0xfea  :    0 - 0x0
    "01000000", -- 4075 - 0xfeb  :   64 - 0x40
    "00000000", -- 4076 - 0xfec  :    0 - 0x0
    "00110001", -- 4077 - 0xfed  :   49 - 0x31
    "00111101", -- 4078 - 0xfee  :   61 - 0x3d
    "00011001", -- 4079 - 0xfef  :   25 - 0x19
    "11000110", -- 4080 - 0xff0  :  198 - 0xc6 -- Sprite 0xff
    "11000100", -- 4081 - 0xff1  :  196 - 0xc4
    "11001100", -- 4082 - 0xff2  :  204 - 0xcc
    "11001100", -- 4083 - 0xff3  :  204 - 0xcc
    "10111000", -- 4084 - 0xff4  :  184 - 0xb8
    "01111100", -- 4085 - 0xff5  :  124 - 0x7c
    "11101100", -- 4086 - 0xff6  :  236 - 0xec
    "11001000", -- 4087 - 0xff7  :  200 - 0xc8
    "00000000", -- 4088 - 0xff8  :    0 - 0x0
    "10000000", -- 4089 - 0xff9  :  128 - 0x80
    "11000000", -- 4090 - 0xffa  :  192 - 0xc0
    "11000000", -- 4091 - 0xffb  :  192 - 0xc0
    "11000000", -- 4092 - 0xffc  :  192 - 0xc0
    "10001000", -- 4093 - 0xffd  :  136 - 0x88
    "10111000", -- 4094 - 0xffe  :  184 - 0xb8
    "10111000", -- 4095 - 0xfff  :  184 - 0xb8
          -- Pattern Table 1---------
    "00111000", -- 4096 - 0x1000  :   56 - 0x38 -- Background 0x0
    "01001100", -- 4097 - 0x1001  :   76 - 0x4c
    "11000110", -- 4098 - 0x1002  :  198 - 0xc6
    "11000110", -- 4099 - 0x1003  :  198 - 0xc6
    "11000110", -- 4100 - 0x1004  :  198 - 0xc6
    "01100100", -- 4101 - 0x1005  :  100 - 0x64
    "00111000", -- 4102 - 0x1006  :   56 - 0x38
    "00000000", -- 4103 - 0x1007  :    0 - 0x0
    "00000000", -- 4104 - 0x1008  :    0 - 0x0
    "00000000", -- 4105 - 0x1009  :    0 - 0x0
    "00000000", -- 4106 - 0x100a  :    0 - 0x0
    "00000000", -- 4107 - 0x100b  :    0 - 0x0
    "00000000", -- 4108 - 0x100c  :    0 - 0x0
    "00000000", -- 4109 - 0x100d  :    0 - 0x0
    "00000000", -- 4110 - 0x100e  :    0 - 0x0
    "00000000", -- 4111 - 0x100f  :    0 - 0x0
    "00011000", -- 4112 - 0x1010  :   24 - 0x18 -- Background 0x1
    "00111000", -- 4113 - 0x1011  :   56 - 0x38
    "00011000", -- 4114 - 0x1012  :   24 - 0x18
    "00011000", -- 4115 - 0x1013  :   24 - 0x18
    "00011000", -- 4116 - 0x1014  :   24 - 0x18
    "00011000", -- 4117 - 0x1015  :   24 - 0x18
    "01111110", -- 4118 - 0x1016  :  126 - 0x7e
    "00000000", -- 4119 - 0x1017  :    0 - 0x0
    "00000000", -- 4120 - 0x1018  :    0 - 0x0
    "00000000", -- 4121 - 0x1019  :    0 - 0x0
    "00000000", -- 4122 - 0x101a  :    0 - 0x0
    "00000000", -- 4123 - 0x101b  :    0 - 0x0
    "00000000", -- 4124 - 0x101c  :    0 - 0x0
    "00000000", -- 4125 - 0x101d  :    0 - 0x0
    "00000000", -- 4126 - 0x101e  :    0 - 0x0
    "00000000", -- 4127 - 0x101f  :    0 - 0x0
    "01111100", -- 4128 - 0x1020  :  124 - 0x7c -- Background 0x2
    "11000110", -- 4129 - 0x1021  :  198 - 0xc6
    "00001110", -- 4130 - 0x1022  :   14 - 0xe
    "00111100", -- 4131 - 0x1023  :   60 - 0x3c
    "01111000", -- 4132 - 0x1024  :  120 - 0x78
    "11100000", -- 4133 - 0x1025  :  224 - 0xe0
    "11111110", -- 4134 - 0x1026  :  254 - 0xfe
    "00000000", -- 4135 - 0x1027  :    0 - 0x0
    "00000000", -- 4136 - 0x1028  :    0 - 0x0
    "00000000", -- 4137 - 0x1029  :    0 - 0x0
    "00000000", -- 4138 - 0x102a  :    0 - 0x0
    "00000000", -- 4139 - 0x102b  :    0 - 0x0
    "00000000", -- 4140 - 0x102c  :    0 - 0x0
    "00000000", -- 4141 - 0x102d  :    0 - 0x0
    "00000000", -- 4142 - 0x102e  :    0 - 0x0
    "00000000", -- 4143 - 0x102f  :    0 - 0x0
    "01111110", -- 4144 - 0x1030  :  126 - 0x7e -- Background 0x3
    "00001100", -- 4145 - 0x1031  :   12 - 0xc
    "00011000", -- 4146 - 0x1032  :   24 - 0x18
    "00111100", -- 4147 - 0x1033  :   60 - 0x3c
    "00000110", -- 4148 - 0x1034  :    6 - 0x6
    "11000110", -- 4149 - 0x1035  :  198 - 0xc6
    "01111100", -- 4150 - 0x1036  :  124 - 0x7c
    "00000000", -- 4151 - 0x1037  :    0 - 0x0
    "00000000", -- 4152 - 0x1038  :    0 - 0x0
    "00000000", -- 4153 - 0x1039  :    0 - 0x0
    "00000000", -- 4154 - 0x103a  :    0 - 0x0
    "00000000", -- 4155 - 0x103b  :    0 - 0x0
    "00000000", -- 4156 - 0x103c  :    0 - 0x0
    "00000000", -- 4157 - 0x103d  :    0 - 0x0
    "00000000", -- 4158 - 0x103e  :    0 - 0x0
    "00000000", -- 4159 - 0x103f  :    0 - 0x0
    "00011100", -- 4160 - 0x1040  :   28 - 0x1c -- Background 0x4
    "00111100", -- 4161 - 0x1041  :   60 - 0x3c
    "01101100", -- 4162 - 0x1042  :  108 - 0x6c
    "11001100", -- 4163 - 0x1043  :  204 - 0xcc
    "11111110", -- 4164 - 0x1044  :  254 - 0xfe
    "00001100", -- 4165 - 0x1045  :   12 - 0xc
    "00001100", -- 4166 - 0x1046  :   12 - 0xc
    "00000000", -- 4167 - 0x1047  :    0 - 0x0
    "00000000", -- 4168 - 0x1048  :    0 - 0x0
    "00000000", -- 4169 - 0x1049  :    0 - 0x0
    "00000000", -- 4170 - 0x104a  :    0 - 0x0
    "00000000", -- 4171 - 0x104b  :    0 - 0x0
    "00000000", -- 4172 - 0x104c  :    0 - 0x0
    "00000000", -- 4173 - 0x104d  :    0 - 0x0
    "00000000", -- 4174 - 0x104e  :    0 - 0x0
    "00000000", -- 4175 - 0x104f  :    0 - 0x0
    "11111100", -- 4176 - 0x1050  :  252 - 0xfc -- Background 0x5
    "11000000", -- 4177 - 0x1051  :  192 - 0xc0
    "11111100", -- 4178 - 0x1052  :  252 - 0xfc
    "00000110", -- 4179 - 0x1053  :    6 - 0x6
    "00000110", -- 4180 - 0x1054  :    6 - 0x6
    "11000110", -- 4181 - 0x1055  :  198 - 0xc6
    "01111100", -- 4182 - 0x1056  :  124 - 0x7c
    "00000000", -- 4183 - 0x1057  :    0 - 0x0
    "00000000", -- 4184 - 0x1058  :    0 - 0x0
    "00000000", -- 4185 - 0x1059  :    0 - 0x0
    "00000000", -- 4186 - 0x105a  :    0 - 0x0
    "00000000", -- 4187 - 0x105b  :    0 - 0x0
    "00000000", -- 4188 - 0x105c  :    0 - 0x0
    "00000000", -- 4189 - 0x105d  :    0 - 0x0
    "00000000", -- 4190 - 0x105e  :    0 - 0x0
    "00000000", -- 4191 - 0x105f  :    0 - 0x0
    "00111100", -- 4192 - 0x1060  :   60 - 0x3c -- Background 0x6
    "01100000", -- 4193 - 0x1061  :   96 - 0x60
    "11000000", -- 4194 - 0x1062  :  192 - 0xc0
    "11111100", -- 4195 - 0x1063  :  252 - 0xfc
    "11000110", -- 4196 - 0x1064  :  198 - 0xc6
    "11000110", -- 4197 - 0x1065  :  198 - 0xc6
    "01111100", -- 4198 - 0x1066  :  124 - 0x7c
    "00000000", -- 4199 - 0x1067  :    0 - 0x0
    "00000000", -- 4200 - 0x1068  :    0 - 0x0
    "00000000", -- 4201 - 0x1069  :    0 - 0x0
    "00000000", -- 4202 - 0x106a  :    0 - 0x0
    "00000000", -- 4203 - 0x106b  :    0 - 0x0
    "00000000", -- 4204 - 0x106c  :    0 - 0x0
    "00000000", -- 4205 - 0x106d  :    0 - 0x0
    "00000000", -- 4206 - 0x106e  :    0 - 0x0
    "00000000", -- 4207 - 0x106f  :    0 - 0x0
    "11111110", -- 4208 - 0x1070  :  254 - 0xfe -- Background 0x7
    "11000110", -- 4209 - 0x1071  :  198 - 0xc6
    "00001100", -- 4210 - 0x1072  :   12 - 0xc
    "00011000", -- 4211 - 0x1073  :   24 - 0x18
    "00110000", -- 4212 - 0x1074  :   48 - 0x30
    "00110000", -- 4213 - 0x1075  :   48 - 0x30
    "00110000", -- 4214 - 0x1076  :   48 - 0x30
    "00000000", -- 4215 - 0x1077  :    0 - 0x0
    "00000000", -- 4216 - 0x1078  :    0 - 0x0
    "00000000", -- 4217 - 0x1079  :    0 - 0x0
    "00000000", -- 4218 - 0x107a  :    0 - 0x0
    "00000000", -- 4219 - 0x107b  :    0 - 0x0
    "00000000", -- 4220 - 0x107c  :    0 - 0x0
    "00000000", -- 4221 - 0x107d  :    0 - 0x0
    "00000000", -- 4222 - 0x107e  :    0 - 0x0
    "00000000", -- 4223 - 0x107f  :    0 - 0x0
    "01111000", -- 4224 - 0x1080  :  120 - 0x78 -- Background 0x8
    "11000100", -- 4225 - 0x1081  :  196 - 0xc4
    "11100100", -- 4226 - 0x1082  :  228 - 0xe4
    "01111000", -- 4227 - 0x1083  :  120 - 0x78
    "10000110", -- 4228 - 0x1084  :  134 - 0x86
    "10000110", -- 4229 - 0x1085  :  134 - 0x86
    "01111100", -- 4230 - 0x1086  :  124 - 0x7c
    "00000000", -- 4231 - 0x1087  :    0 - 0x0
    "00000000", -- 4232 - 0x1088  :    0 - 0x0
    "00000000", -- 4233 - 0x1089  :    0 - 0x0
    "00000000", -- 4234 - 0x108a  :    0 - 0x0
    "00000000", -- 4235 - 0x108b  :    0 - 0x0
    "00000000", -- 4236 - 0x108c  :    0 - 0x0
    "00000000", -- 4237 - 0x108d  :    0 - 0x0
    "00000000", -- 4238 - 0x108e  :    0 - 0x0
    "00000000", -- 4239 - 0x108f  :    0 - 0x0
    "01111100", -- 4240 - 0x1090  :  124 - 0x7c -- Background 0x9
    "11000110", -- 4241 - 0x1091  :  198 - 0xc6
    "11000110", -- 4242 - 0x1092  :  198 - 0xc6
    "01111110", -- 4243 - 0x1093  :  126 - 0x7e
    "00000110", -- 4244 - 0x1094  :    6 - 0x6
    "00001100", -- 4245 - 0x1095  :   12 - 0xc
    "01111000", -- 4246 - 0x1096  :  120 - 0x78
    "00000000", -- 4247 - 0x1097  :    0 - 0x0
    "00000000", -- 4248 - 0x1098  :    0 - 0x0
    "00000000", -- 4249 - 0x1099  :    0 - 0x0
    "00000000", -- 4250 - 0x109a  :    0 - 0x0
    "00000000", -- 4251 - 0x109b  :    0 - 0x0
    "00000000", -- 4252 - 0x109c  :    0 - 0x0
    "00000000", -- 4253 - 0x109d  :    0 - 0x0
    "00000000", -- 4254 - 0x109e  :    0 - 0x0
    "00000000", -- 4255 - 0x109f  :    0 - 0x0
    "00111000", -- 4256 - 0x10a0  :   56 - 0x38 -- Background 0xa
    "01101100", -- 4257 - 0x10a1  :  108 - 0x6c
    "11000110", -- 4258 - 0x10a2  :  198 - 0xc6
    "11000110", -- 4259 - 0x10a3  :  198 - 0xc6
    "11111110", -- 4260 - 0x10a4  :  254 - 0xfe
    "11000110", -- 4261 - 0x10a5  :  198 - 0xc6
    "11000110", -- 4262 - 0x10a6  :  198 - 0xc6
    "00000000", -- 4263 - 0x10a7  :    0 - 0x0
    "00000000", -- 4264 - 0x10a8  :    0 - 0x0
    "00000000", -- 4265 - 0x10a9  :    0 - 0x0
    "00000000", -- 4266 - 0x10aa  :    0 - 0x0
    "00000000", -- 4267 - 0x10ab  :    0 - 0x0
    "00000000", -- 4268 - 0x10ac  :    0 - 0x0
    "00000000", -- 4269 - 0x10ad  :    0 - 0x0
    "00000000", -- 4270 - 0x10ae  :    0 - 0x0
    "00000000", -- 4271 - 0x10af  :    0 - 0x0
    "11111100", -- 4272 - 0x10b0  :  252 - 0xfc -- Background 0xb
    "11000110", -- 4273 - 0x10b1  :  198 - 0xc6
    "11000110", -- 4274 - 0x10b2  :  198 - 0xc6
    "11111100", -- 4275 - 0x10b3  :  252 - 0xfc
    "11000110", -- 4276 - 0x10b4  :  198 - 0xc6
    "11000110", -- 4277 - 0x10b5  :  198 - 0xc6
    "11111100", -- 4278 - 0x10b6  :  252 - 0xfc
    "00000000", -- 4279 - 0x10b7  :    0 - 0x0
    "00000000", -- 4280 - 0x10b8  :    0 - 0x0
    "00000000", -- 4281 - 0x10b9  :    0 - 0x0
    "00000000", -- 4282 - 0x10ba  :    0 - 0x0
    "00000000", -- 4283 - 0x10bb  :    0 - 0x0
    "00000000", -- 4284 - 0x10bc  :    0 - 0x0
    "00000000", -- 4285 - 0x10bd  :    0 - 0x0
    "00000000", -- 4286 - 0x10be  :    0 - 0x0
    "00000000", -- 4287 - 0x10bf  :    0 - 0x0
    "00111100", -- 4288 - 0x10c0  :   60 - 0x3c -- Background 0xc
    "01100110", -- 4289 - 0x10c1  :  102 - 0x66
    "11000000", -- 4290 - 0x10c2  :  192 - 0xc0
    "11000000", -- 4291 - 0x10c3  :  192 - 0xc0
    "11000000", -- 4292 - 0x10c4  :  192 - 0xc0
    "01100110", -- 4293 - 0x10c5  :  102 - 0x66
    "00111100", -- 4294 - 0x10c6  :   60 - 0x3c
    "00000000", -- 4295 - 0x10c7  :    0 - 0x0
    "00000000", -- 4296 - 0x10c8  :    0 - 0x0
    "00000000", -- 4297 - 0x10c9  :    0 - 0x0
    "00000000", -- 4298 - 0x10ca  :    0 - 0x0
    "00000000", -- 4299 - 0x10cb  :    0 - 0x0
    "00000000", -- 4300 - 0x10cc  :    0 - 0x0
    "00000000", -- 4301 - 0x10cd  :    0 - 0x0
    "00000000", -- 4302 - 0x10ce  :    0 - 0x0
    "00000000", -- 4303 - 0x10cf  :    0 - 0x0
    "11111000", -- 4304 - 0x10d0  :  248 - 0xf8 -- Background 0xd
    "11001100", -- 4305 - 0x10d1  :  204 - 0xcc
    "11000110", -- 4306 - 0x10d2  :  198 - 0xc6
    "11000110", -- 4307 - 0x10d3  :  198 - 0xc6
    "11000110", -- 4308 - 0x10d4  :  198 - 0xc6
    "11001100", -- 4309 - 0x10d5  :  204 - 0xcc
    "11111000", -- 4310 - 0x10d6  :  248 - 0xf8
    "00000000", -- 4311 - 0x10d7  :    0 - 0x0
    "00000000", -- 4312 - 0x10d8  :    0 - 0x0
    "00000000", -- 4313 - 0x10d9  :    0 - 0x0
    "00000000", -- 4314 - 0x10da  :    0 - 0x0
    "00000000", -- 4315 - 0x10db  :    0 - 0x0
    "00000000", -- 4316 - 0x10dc  :    0 - 0x0
    "00000000", -- 4317 - 0x10dd  :    0 - 0x0
    "00000000", -- 4318 - 0x10de  :    0 - 0x0
    "00000000", -- 4319 - 0x10df  :    0 - 0x0
    "11111110", -- 4320 - 0x10e0  :  254 - 0xfe -- Background 0xe
    "11000000", -- 4321 - 0x10e1  :  192 - 0xc0
    "11000000", -- 4322 - 0x10e2  :  192 - 0xc0
    "11111100", -- 4323 - 0x10e3  :  252 - 0xfc
    "11000000", -- 4324 - 0x10e4  :  192 - 0xc0
    "11000000", -- 4325 - 0x10e5  :  192 - 0xc0
    "11111110", -- 4326 - 0x10e6  :  254 - 0xfe
    "00000000", -- 4327 - 0x10e7  :    0 - 0x0
    "00000000", -- 4328 - 0x10e8  :    0 - 0x0
    "00000000", -- 4329 - 0x10e9  :    0 - 0x0
    "00000000", -- 4330 - 0x10ea  :    0 - 0x0
    "00000000", -- 4331 - 0x10eb  :    0 - 0x0
    "00000000", -- 4332 - 0x10ec  :    0 - 0x0
    "00000000", -- 4333 - 0x10ed  :    0 - 0x0
    "00000000", -- 4334 - 0x10ee  :    0 - 0x0
    "00000000", -- 4335 - 0x10ef  :    0 - 0x0
    "11111110", -- 4336 - 0x10f0  :  254 - 0xfe -- Background 0xf
    "11000000", -- 4337 - 0x10f1  :  192 - 0xc0
    "11000000", -- 4338 - 0x10f2  :  192 - 0xc0
    "11111100", -- 4339 - 0x10f3  :  252 - 0xfc
    "11000000", -- 4340 - 0x10f4  :  192 - 0xc0
    "11000000", -- 4341 - 0x10f5  :  192 - 0xc0
    "11000000", -- 4342 - 0x10f6  :  192 - 0xc0
    "00000000", -- 4343 - 0x10f7  :    0 - 0x0
    "00000000", -- 4344 - 0x10f8  :    0 - 0x0
    "00000000", -- 4345 - 0x10f9  :    0 - 0x0
    "00000000", -- 4346 - 0x10fa  :    0 - 0x0
    "00000000", -- 4347 - 0x10fb  :    0 - 0x0
    "00000000", -- 4348 - 0x10fc  :    0 - 0x0
    "00000000", -- 4349 - 0x10fd  :    0 - 0x0
    "00000000", -- 4350 - 0x10fe  :    0 - 0x0
    "00000000", -- 4351 - 0x10ff  :    0 - 0x0
    "00111110", -- 4352 - 0x1100  :   62 - 0x3e -- Background 0x10
    "01100000", -- 4353 - 0x1101  :   96 - 0x60
    "11000000", -- 4354 - 0x1102  :  192 - 0xc0
    "11011110", -- 4355 - 0x1103  :  222 - 0xde
    "11000110", -- 4356 - 0x1104  :  198 - 0xc6
    "01100110", -- 4357 - 0x1105  :  102 - 0x66
    "01111110", -- 4358 - 0x1106  :  126 - 0x7e
    "00000000", -- 4359 - 0x1107  :    0 - 0x0
    "00000000", -- 4360 - 0x1108  :    0 - 0x0
    "00000000", -- 4361 - 0x1109  :    0 - 0x0
    "00000000", -- 4362 - 0x110a  :    0 - 0x0
    "00000000", -- 4363 - 0x110b  :    0 - 0x0
    "00000000", -- 4364 - 0x110c  :    0 - 0x0
    "00000000", -- 4365 - 0x110d  :    0 - 0x0
    "00000000", -- 4366 - 0x110e  :    0 - 0x0
    "00000000", -- 4367 - 0x110f  :    0 - 0x0
    "11000110", -- 4368 - 0x1110  :  198 - 0xc6 -- Background 0x11
    "11000110", -- 4369 - 0x1111  :  198 - 0xc6
    "11000110", -- 4370 - 0x1112  :  198 - 0xc6
    "11111110", -- 4371 - 0x1113  :  254 - 0xfe
    "11000110", -- 4372 - 0x1114  :  198 - 0xc6
    "11000110", -- 4373 - 0x1115  :  198 - 0xc6
    "11000110", -- 4374 - 0x1116  :  198 - 0xc6
    "00000000", -- 4375 - 0x1117  :    0 - 0x0
    "00000000", -- 4376 - 0x1118  :    0 - 0x0
    "00000000", -- 4377 - 0x1119  :    0 - 0x0
    "00000000", -- 4378 - 0x111a  :    0 - 0x0
    "00000000", -- 4379 - 0x111b  :    0 - 0x0
    "00000000", -- 4380 - 0x111c  :    0 - 0x0
    "00000000", -- 4381 - 0x111d  :    0 - 0x0
    "00000000", -- 4382 - 0x111e  :    0 - 0x0
    "00000000", -- 4383 - 0x111f  :    0 - 0x0
    "01111110", -- 4384 - 0x1120  :  126 - 0x7e -- Background 0x12
    "00011000", -- 4385 - 0x1121  :   24 - 0x18
    "00011000", -- 4386 - 0x1122  :   24 - 0x18
    "00011000", -- 4387 - 0x1123  :   24 - 0x18
    "00011000", -- 4388 - 0x1124  :   24 - 0x18
    "00011000", -- 4389 - 0x1125  :   24 - 0x18
    "01111110", -- 4390 - 0x1126  :  126 - 0x7e
    "00000000", -- 4391 - 0x1127  :    0 - 0x0
    "00000000", -- 4392 - 0x1128  :    0 - 0x0
    "00000000", -- 4393 - 0x1129  :    0 - 0x0
    "00000000", -- 4394 - 0x112a  :    0 - 0x0
    "00000000", -- 4395 - 0x112b  :    0 - 0x0
    "00000000", -- 4396 - 0x112c  :    0 - 0x0
    "00000000", -- 4397 - 0x112d  :    0 - 0x0
    "00000000", -- 4398 - 0x112e  :    0 - 0x0
    "00000000", -- 4399 - 0x112f  :    0 - 0x0
    "00011110", -- 4400 - 0x1130  :   30 - 0x1e -- Background 0x13
    "00000110", -- 4401 - 0x1131  :    6 - 0x6
    "00000110", -- 4402 - 0x1132  :    6 - 0x6
    "00000110", -- 4403 - 0x1133  :    6 - 0x6
    "11000110", -- 4404 - 0x1134  :  198 - 0xc6
    "11000110", -- 4405 - 0x1135  :  198 - 0xc6
    "01111100", -- 4406 - 0x1136  :  124 - 0x7c
    "00000000", -- 4407 - 0x1137  :    0 - 0x0
    "00000000", -- 4408 - 0x1138  :    0 - 0x0
    "00000000", -- 4409 - 0x1139  :    0 - 0x0
    "00000000", -- 4410 - 0x113a  :    0 - 0x0
    "00000000", -- 4411 - 0x113b  :    0 - 0x0
    "00000000", -- 4412 - 0x113c  :    0 - 0x0
    "00000000", -- 4413 - 0x113d  :    0 - 0x0
    "00000000", -- 4414 - 0x113e  :    0 - 0x0
    "00000000", -- 4415 - 0x113f  :    0 - 0x0
    "11000110", -- 4416 - 0x1140  :  198 - 0xc6 -- Background 0x14
    "11001100", -- 4417 - 0x1141  :  204 - 0xcc
    "11011000", -- 4418 - 0x1142  :  216 - 0xd8
    "11110000", -- 4419 - 0x1143  :  240 - 0xf0
    "11111000", -- 4420 - 0x1144  :  248 - 0xf8
    "11011100", -- 4421 - 0x1145  :  220 - 0xdc
    "11001110", -- 4422 - 0x1146  :  206 - 0xce
    "00000000", -- 4423 - 0x1147  :    0 - 0x0
    "00000000", -- 4424 - 0x1148  :    0 - 0x0
    "00000000", -- 4425 - 0x1149  :    0 - 0x0
    "00000000", -- 4426 - 0x114a  :    0 - 0x0
    "00000000", -- 4427 - 0x114b  :    0 - 0x0
    "00000000", -- 4428 - 0x114c  :    0 - 0x0
    "00000000", -- 4429 - 0x114d  :    0 - 0x0
    "00000000", -- 4430 - 0x114e  :    0 - 0x0
    "00000000", -- 4431 - 0x114f  :    0 - 0x0
    "01100000", -- 4432 - 0x1150  :   96 - 0x60 -- Background 0x15
    "01100000", -- 4433 - 0x1151  :   96 - 0x60
    "01100000", -- 4434 - 0x1152  :   96 - 0x60
    "01100000", -- 4435 - 0x1153  :   96 - 0x60
    "01100000", -- 4436 - 0x1154  :   96 - 0x60
    "01100000", -- 4437 - 0x1155  :   96 - 0x60
    "01111110", -- 4438 - 0x1156  :  126 - 0x7e
    "00000000", -- 4439 - 0x1157  :    0 - 0x0
    "00000000", -- 4440 - 0x1158  :    0 - 0x0
    "00000000", -- 4441 - 0x1159  :    0 - 0x0
    "00000000", -- 4442 - 0x115a  :    0 - 0x0
    "00000000", -- 4443 - 0x115b  :    0 - 0x0
    "00000000", -- 4444 - 0x115c  :    0 - 0x0
    "00000000", -- 4445 - 0x115d  :    0 - 0x0
    "00000000", -- 4446 - 0x115e  :    0 - 0x0
    "00000000", -- 4447 - 0x115f  :    0 - 0x0
    "11000110", -- 4448 - 0x1160  :  198 - 0xc6 -- Background 0x16
    "11101110", -- 4449 - 0x1161  :  238 - 0xee
    "11111110", -- 4450 - 0x1162  :  254 - 0xfe
    "11111110", -- 4451 - 0x1163  :  254 - 0xfe
    "11010110", -- 4452 - 0x1164  :  214 - 0xd6
    "11000110", -- 4453 - 0x1165  :  198 - 0xc6
    "11000110", -- 4454 - 0x1166  :  198 - 0xc6
    "00000000", -- 4455 - 0x1167  :    0 - 0x0
    "00000000", -- 4456 - 0x1168  :    0 - 0x0
    "00000000", -- 4457 - 0x1169  :    0 - 0x0
    "00000000", -- 4458 - 0x116a  :    0 - 0x0
    "00000000", -- 4459 - 0x116b  :    0 - 0x0
    "00000000", -- 4460 - 0x116c  :    0 - 0x0
    "00000000", -- 4461 - 0x116d  :    0 - 0x0
    "00000000", -- 4462 - 0x116e  :    0 - 0x0
    "00000000", -- 4463 - 0x116f  :    0 - 0x0
    "11000110", -- 4464 - 0x1170  :  198 - 0xc6 -- Background 0x17
    "11100110", -- 4465 - 0x1171  :  230 - 0xe6
    "11110110", -- 4466 - 0x1172  :  246 - 0xf6
    "11111110", -- 4467 - 0x1173  :  254 - 0xfe
    "11011110", -- 4468 - 0x1174  :  222 - 0xde
    "11001110", -- 4469 - 0x1175  :  206 - 0xce
    "11000110", -- 4470 - 0x1176  :  198 - 0xc6
    "00000000", -- 4471 - 0x1177  :    0 - 0x0
    "00000000", -- 4472 - 0x1178  :    0 - 0x0
    "00000000", -- 4473 - 0x1179  :    0 - 0x0
    "00000000", -- 4474 - 0x117a  :    0 - 0x0
    "00000000", -- 4475 - 0x117b  :    0 - 0x0
    "00000000", -- 4476 - 0x117c  :    0 - 0x0
    "00000000", -- 4477 - 0x117d  :    0 - 0x0
    "00000000", -- 4478 - 0x117e  :    0 - 0x0
    "00000000", -- 4479 - 0x117f  :    0 - 0x0
    "01111100", -- 4480 - 0x1180  :  124 - 0x7c -- Background 0x18
    "11000110", -- 4481 - 0x1181  :  198 - 0xc6
    "11000110", -- 4482 - 0x1182  :  198 - 0xc6
    "11000110", -- 4483 - 0x1183  :  198 - 0xc6
    "11000110", -- 4484 - 0x1184  :  198 - 0xc6
    "11000110", -- 4485 - 0x1185  :  198 - 0xc6
    "01111100", -- 4486 - 0x1186  :  124 - 0x7c
    "00000000", -- 4487 - 0x1187  :    0 - 0x0
    "00000000", -- 4488 - 0x1188  :    0 - 0x0
    "00000000", -- 4489 - 0x1189  :    0 - 0x0
    "00000000", -- 4490 - 0x118a  :    0 - 0x0
    "00000000", -- 4491 - 0x118b  :    0 - 0x0
    "00000000", -- 4492 - 0x118c  :    0 - 0x0
    "00000000", -- 4493 - 0x118d  :    0 - 0x0
    "00000000", -- 4494 - 0x118e  :    0 - 0x0
    "00000000", -- 4495 - 0x118f  :    0 - 0x0
    "11111100", -- 4496 - 0x1190  :  252 - 0xfc -- Background 0x19
    "11000110", -- 4497 - 0x1191  :  198 - 0xc6
    "11000110", -- 4498 - 0x1192  :  198 - 0xc6
    "11000110", -- 4499 - 0x1193  :  198 - 0xc6
    "11111100", -- 4500 - 0x1194  :  252 - 0xfc
    "11000000", -- 4501 - 0x1195  :  192 - 0xc0
    "11000000", -- 4502 - 0x1196  :  192 - 0xc0
    "00000000", -- 4503 - 0x1197  :    0 - 0x0
    "00000000", -- 4504 - 0x1198  :    0 - 0x0
    "00000000", -- 4505 - 0x1199  :    0 - 0x0
    "00000000", -- 4506 - 0x119a  :    0 - 0x0
    "00000000", -- 4507 - 0x119b  :    0 - 0x0
    "00000000", -- 4508 - 0x119c  :    0 - 0x0
    "00000000", -- 4509 - 0x119d  :    0 - 0x0
    "00000000", -- 4510 - 0x119e  :    0 - 0x0
    "00000000", -- 4511 - 0x119f  :    0 - 0x0
    "01111100", -- 4512 - 0x11a0  :  124 - 0x7c -- Background 0x1a
    "11000110", -- 4513 - 0x11a1  :  198 - 0xc6
    "11000110", -- 4514 - 0x11a2  :  198 - 0xc6
    "11000110", -- 4515 - 0x11a3  :  198 - 0xc6
    "11011110", -- 4516 - 0x11a4  :  222 - 0xde
    "11001100", -- 4517 - 0x11a5  :  204 - 0xcc
    "01111010", -- 4518 - 0x11a6  :  122 - 0x7a
    "00000000", -- 4519 - 0x11a7  :    0 - 0x0
    "00000000", -- 4520 - 0x11a8  :    0 - 0x0
    "00000000", -- 4521 - 0x11a9  :    0 - 0x0
    "00000000", -- 4522 - 0x11aa  :    0 - 0x0
    "00000000", -- 4523 - 0x11ab  :    0 - 0x0
    "00000000", -- 4524 - 0x11ac  :    0 - 0x0
    "00000000", -- 4525 - 0x11ad  :    0 - 0x0
    "00000000", -- 4526 - 0x11ae  :    0 - 0x0
    "00000000", -- 4527 - 0x11af  :    0 - 0x0
    "11111100", -- 4528 - 0x11b0  :  252 - 0xfc -- Background 0x1b
    "11000110", -- 4529 - 0x11b1  :  198 - 0xc6
    "11000110", -- 4530 - 0x11b2  :  198 - 0xc6
    "11001110", -- 4531 - 0x11b3  :  206 - 0xce
    "11111000", -- 4532 - 0x11b4  :  248 - 0xf8
    "11011100", -- 4533 - 0x11b5  :  220 - 0xdc
    "11001110", -- 4534 - 0x11b6  :  206 - 0xce
    "00000000", -- 4535 - 0x11b7  :    0 - 0x0
    "00000000", -- 4536 - 0x11b8  :    0 - 0x0
    "00000000", -- 4537 - 0x11b9  :    0 - 0x0
    "00000000", -- 4538 - 0x11ba  :    0 - 0x0
    "00000000", -- 4539 - 0x11bb  :    0 - 0x0
    "00000000", -- 4540 - 0x11bc  :    0 - 0x0
    "00000000", -- 4541 - 0x11bd  :    0 - 0x0
    "00000000", -- 4542 - 0x11be  :    0 - 0x0
    "00000000", -- 4543 - 0x11bf  :    0 - 0x0
    "01111000", -- 4544 - 0x11c0  :  120 - 0x78 -- Background 0x1c
    "11001100", -- 4545 - 0x11c1  :  204 - 0xcc
    "11000000", -- 4546 - 0x11c2  :  192 - 0xc0
    "01111100", -- 4547 - 0x11c3  :  124 - 0x7c
    "00000110", -- 4548 - 0x11c4  :    6 - 0x6
    "11000110", -- 4549 - 0x11c5  :  198 - 0xc6
    "01111100", -- 4550 - 0x11c6  :  124 - 0x7c
    "00000000", -- 4551 - 0x11c7  :    0 - 0x0
    "00000000", -- 4552 - 0x11c8  :    0 - 0x0
    "00000000", -- 4553 - 0x11c9  :    0 - 0x0
    "00000000", -- 4554 - 0x11ca  :    0 - 0x0
    "00000000", -- 4555 - 0x11cb  :    0 - 0x0
    "00000000", -- 4556 - 0x11cc  :    0 - 0x0
    "00000000", -- 4557 - 0x11cd  :    0 - 0x0
    "00000000", -- 4558 - 0x11ce  :    0 - 0x0
    "00000000", -- 4559 - 0x11cf  :    0 - 0x0
    "01111110", -- 4560 - 0x11d0  :  126 - 0x7e -- Background 0x1d
    "00011000", -- 4561 - 0x11d1  :   24 - 0x18
    "00011000", -- 4562 - 0x11d2  :   24 - 0x18
    "00011000", -- 4563 - 0x11d3  :   24 - 0x18
    "00011000", -- 4564 - 0x11d4  :   24 - 0x18
    "00011000", -- 4565 - 0x11d5  :   24 - 0x18
    "00011000", -- 4566 - 0x11d6  :   24 - 0x18
    "00000000", -- 4567 - 0x11d7  :    0 - 0x0
    "00000000", -- 4568 - 0x11d8  :    0 - 0x0
    "00000000", -- 4569 - 0x11d9  :    0 - 0x0
    "00000000", -- 4570 - 0x11da  :    0 - 0x0
    "00000000", -- 4571 - 0x11db  :    0 - 0x0
    "00000000", -- 4572 - 0x11dc  :    0 - 0x0
    "00000000", -- 4573 - 0x11dd  :    0 - 0x0
    "00000000", -- 4574 - 0x11de  :    0 - 0x0
    "00000000", -- 4575 - 0x11df  :    0 - 0x0
    "11000110", -- 4576 - 0x11e0  :  198 - 0xc6 -- Background 0x1e
    "11000110", -- 4577 - 0x11e1  :  198 - 0xc6
    "11000110", -- 4578 - 0x11e2  :  198 - 0xc6
    "11000110", -- 4579 - 0x11e3  :  198 - 0xc6
    "11000110", -- 4580 - 0x11e4  :  198 - 0xc6
    "11000110", -- 4581 - 0x11e5  :  198 - 0xc6
    "01111100", -- 4582 - 0x11e6  :  124 - 0x7c
    "00000000", -- 4583 - 0x11e7  :    0 - 0x0
    "00000000", -- 4584 - 0x11e8  :    0 - 0x0
    "00000000", -- 4585 - 0x11e9  :    0 - 0x0
    "00000000", -- 4586 - 0x11ea  :    0 - 0x0
    "00000000", -- 4587 - 0x11eb  :    0 - 0x0
    "00000000", -- 4588 - 0x11ec  :    0 - 0x0
    "00000000", -- 4589 - 0x11ed  :    0 - 0x0
    "00000000", -- 4590 - 0x11ee  :    0 - 0x0
    "00000000", -- 4591 - 0x11ef  :    0 - 0x0
    "11000110", -- 4592 - 0x11f0  :  198 - 0xc6 -- Background 0x1f
    "11000110", -- 4593 - 0x11f1  :  198 - 0xc6
    "11000110", -- 4594 - 0x11f2  :  198 - 0xc6
    "11101110", -- 4595 - 0x11f3  :  238 - 0xee
    "01111100", -- 4596 - 0x11f4  :  124 - 0x7c
    "00111000", -- 4597 - 0x11f5  :   56 - 0x38
    "00010000", -- 4598 - 0x11f6  :   16 - 0x10
    "00000000", -- 4599 - 0x11f7  :    0 - 0x0
    "00000000", -- 4600 - 0x11f8  :    0 - 0x0
    "00000000", -- 4601 - 0x11f9  :    0 - 0x0
    "00000000", -- 4602 - 0x11fa  :    0 - 0x0
    "00000000", -- 4603 - 0x11fb  :    0 - 0x0
    "00000000", -- 4604 - 0x11fc  :    0 - 0x0
    "00000000", -- 4605 - 0x11fd  :    0 - 0x0
    "00000000", -- 4606 - 0x11fe  :    0 - 0x0
    "00000000", -- 4607 - 0x11ff  :    0 - 0x0
    "11000110", -- 4608 - 0x1200  :  198 - 0xc6 -- Background 0x20
    "11000110", -- 4609 - 0x1201  :  198 - 0xc6
    "11010110", -- 4610 - 0x1202  :  214 - 0xd6
    "11111110", -- 4611 - 0x1203  :  254 - 0xfe
    "11111110", -- 4612 - 0x1204  :  254 - 0xfe
    "11101110", -- 4613 - 0x1205  :  238 - 0xee
    "11000110", -- 4614 - 0x1206  :  198 - 0xc6
    "00000000", -- 4615 - 0x1207  :    0 - 0x0
    "00000000", -- 4616 - 0x1208  :    0 - 0x0
    "00000000", -- 4617 - 0x1209  :    0 - 0x0
    "00000000", -- 4618 - 0x120a  :    0 - 0x0
    "00000000", -- 4619 - 0x120b  :    0 - 0x0
    "00000000", -- 4620 - 0x120c  :    0 - 0x0
    "00000000", -- 4621 - 0x120d  :    0 - 0x0
    "00000000", -- 4622 - 0x120e  :    0 - 0x0
    "00000000", -- 4623 - 0x120f  :    0 - 0x0
    "11000110", -- 4624 - 0x1210  :  198 - 0xc6 -- Background 0x21
    "11101110", -- 4625 - 0x1211  :  238 - 0xee
    "01111100", -- 4626 - 0x1212  :  124 - 0x7c
    "00111000", -- 4627 - 0x1213  :   56 - 0x38
    "01111100", -- 4628 - 0x1214  :  124 - 0x7c
    "11101110", -- 4629 - 0x1215  :  238 - 0xee
    "11000110", -- 4630 - 0x1216  :  198 - 0xc6
    "00000000", -- 4631 - 0x1217  :    0 - 0x0
    "00000000", -- 4632 - 0x1218  :    0 - 0x0
    "00000000", -- 4633 - 0x1219  :    0 - 0x0
    "00000000", -- 4634 - 0x121a  :    0 - 0x0
    "00000000", -- 4635 - 0x121b  :    0 - 0x0
    "00000000", -- 4636 - 0x121c  :    0 - 0x0
    "00000000", -- 4637 - 0x121d  :    0 - 0x0
    "00000000", -- 4638 - 0x121e  :    0 - 0x0
    "00000000", -- 4639 - 0x121f  :    0 - 0x0
    "01100110", -- 4640 - 0x1220  :  102 - 0x66 -- Background 0x22
    "01100110", -- 4641 - 0x1221  :  102 - 0x66
    "01100110", -- 4642 - 0x1222  :  102 - 0x66
    "00111100", -- 4643 - 0x1223  :   60 - 0x3c
    "00011000", -- 4644 - 0x1224  :   24 - 0x18
    "00011000", -- 4645 - 0x1225  :   24 - 0x18
    "00011000", -- 4646 - 0x1226  :   24 - 0x18
    "00000000", -- 4647 - 0x1227  :    0 - 0x0
    "00000000", -- 4648 - 0x1228  :    0 - 0x0
    "00000000", -- 4649 - 0x1229  :    0 - 0x0
    "00000000", -- 4650 - 0x122a  :    0 - 0x0
    "00000000", -- 4651 - 0x122b  :    0 - 0x0
    "00000000", -- 4652 - 0x122c  :    0 - 0x0
    "00000000", -- 4653 - 0x122d  :    0 - 0x0
    "00000000", -- 4654 - 0x122e  :    0 - 0x0
    "00000000", -- 4655 - 0x122f  :    0 - 0x0
    "11111110", -- 4656 - 0x1230  :  254 - 0xfe -- Background 0x23
    "00001110", -- 4657 - 0x1231  :   14 - 0xe
    "00011100", -- 4658 - 0x1232  :   28 - 0x1c
    "00111000", -- 4659 - 0x1233  :   56 - 0x38
    "01110000", -- 4660 - 0x1234  :  112 - 0x70
    "11100000", -- 4661 - 0x1235  :  224 - 0xe0
    "11111110", -- 4662 - 0x1236  :  254 - 0xfe
    "00000000", -- 4663 - 0x1237  :    0 - 0x0
    "00000000", -- 4664 - 0x1238  :    0 - 0x0
    "00000000", -- 4665 - 0x1239  :    0 - 0x0
    "00000000", -- 4666 - 0x123a  :    0 - 0x0
    "00000000", -- 4667 - 0x123b  :    0 - 0x0
    "00000000", -- 4668 - 0x123c  :    0 - 0x0
    "00000000", -- 4669 - 0x123d  :    0 - 0x0
    "00000000", -- 4670 - 0x123e  :    0 - 0x0
    "00000000", -- 4671 - 0x123f  :    0 - 0x0
    "00000000", -- 4672 - 0x1240  :    0 - 0x0 -- Background 0x24
    "00000000", -- 4673 - 0x1241  :    0 - 0x0
    "00000000", -- 4674 - 0x1242  :    0 - 0x0
    "00000000", -- 4675 - 0x1243  :    0 - 0x0
    "00000000", -- 4676 - 0x1244  :    0 - 0x0
    "00000000", -- 4677 - 0x1245  :    0 - 0x0
    "00000000", -- 4678 - 0x1246  :    0 - 0x0
    "00000000", -- 4679 - 0x1247  :    0 - 0x0
    "00000000", -- 4680 - 0x1248  :    0 - 0x0
    "00000000", -- 4681 - 0x1249  :    0 - 0x0
    "00000000", -- 4682 - 0x124a  :    0 - 0x0
    "00000000", -- 4683 - 0x124b  :    0 - 0x0
    "00000000", -- 4684 - 0x124c  :    0 - 0x0
    "00000000", -- 4685 - 0x124d  :    0 - 0x0
    "00000000", -- 4686 - 0x124e  :    0 - 0x0
    "00000000", -- 4687 - 0x124f  :    0 - 0x0
    "00000000", -- 4688 - 0x1250  :    0 - 0x0 -- Background 0x25
    "00000000", -- 4689 - 0x1251  :    0 - 0x0
    "00000110", -- 4690 - 0x1252  :    6 - 0x6
    "00001110", -- 4691 - 0x1253  :   14 - 0xe
    "00001000", -- 4692 - 0x1254  :    8 - 0x8
    "00001000", -- 4693 - 0x1255  :    8 - 0x8
    "00001000", -- 4694 - 0x1256  :    8 - 0x8
    "00001000", -- 4695 - 0x1257  :    8 - 0x8
    "00000000", -- 4696 - 0x1258  :    0 - 0x0
    "00000000", -- 4697 - 0x1259  :    0 - 0x0
    "00000000", -- 4698 - 0x125a  :    0 - 0x0
    "00000000", -- 4699 - 0x125b  :    0 - 0x0
    "00000000", -- 4700 - 0x125c  :    0 - 0x0
    "00000000", -- 4701 - 0x125d  :    0 - 0x0
    "00000000", -- 4702 - 0x125e  :    0 - 0x0
    "00000000", -- 4703 - 0x125f  :    0 - 0x0
    "00000000", -- 4704 - 0x1260  :    0 - 0x0 -- Background 0x26
    "01111000", -- 4705 - 0x1261  :  120 - 0x78
    "01100101", -- 4706 - 0x1262  :  101 - 0x65
    "01111001", -- 4707 - 0x1263  :  121 - 0x79
    "01100101", -- 4708 - 0x1264  :  101 - 0x65
    "01100101", -- 4709 - 0x1265  :  101 - 0x65
    "01111000", -- 4710 - 0x1266  :  120 - 0x78
    "00000000", -- 4711 - 0x1267  :    0 - 0x0
    "00000000", -- 4712 - 0x1268  :    0 - 0x0
    "00000000", -- 4713 - 0x1269  :    0 - 0x0
    "00000000", -- 4714 - 0x126a  :    0 - 0x0
    "00000000", -- 4715 - 0x126b  :    0 - 0x0
    "00000000", -- 4716 - 0x126c  :    0 - 0x0
    "00000000", -- 4717 - 0x126d  :    0 - 0x0
    "00000000", -- 4718 - 0x126e  :    0 - 0x0
    "00000000", -- 4719 - 0x126f  :    0 - 0x0
    "00000000", -- 4720 - 0x1270  :    0 - 0x0 -- Background 0x27
    "11100100", -- 4721 - 0x1271  :  228 - 0xe4
    "10010110", -- 4722 - 0x1272  :  150 - 0x96
    "10010110", -- 4723 - 0x1273  :  150 - 0x96
    "10010111", -- 4724 - 0x1274  :  151 - 0x97
    "10010110", -- 4725 - 0x1275  :  150 - 0x96
    "11100110", -- 4726 - 0x1276  :  230 - 0xe6
    "00000000", -- 4727 - 0x1277  :    0 - 0x0
    "00000000", -- 4728 - 0x1278  :    0 - 0x0
    "00000000", -- 4729 - 0x1279  :    0 - 0x0
    "00000000", -- 4730 - 0x127a  :    0 - 0x0
    "00000000", -- 4731 - 0x127b  :    0 - 0x0
    "00000000", -- 4732 - 0x127c  :    0 - 0x0
    "00000000", -- 4733 - 0x127d  :    0 - 0x0
    "00000000", -- 4734 - 0x127e  :    0 - 0x0
    "00000000", -- 4735 - 0x127f  :    0 - 0x0
    "00000000", -- 4736 - 0x1280  :    0 - 0x0 -- Background 0x28
    "01011001", -- 4737 - 0x1281  :   89 - 0x59
    "01011001", -- 4738 - 0x1282  :   89 - 0x59
    "01011001", -- 4739 - 0x1283  :   89 - 0x59
    "01011001", -- 4740 - 0x1284  :   89 - 0x59
    "11011001", -- 4741 - 0x1285  :  217 - 0xd9
    "01001110", -- 4742 - 0x1286  :   78 - 0x4e
    "00000000", -- 4743 - 0x1287  :    0 - 0x0
    "00000000", -- 4744 - 0x1288  :    0 - 0x0
    "00000000", -- 4745 - 0x1289  :    0 - 0x0
    "00000000", -- 4746 - 0x128a  :    0 - 0x0
    "00000000", -- 4747 - 0x128b  :    0 - 0x0
    "00000000", -- 4748 - 0x128c  :    0 - 0x0
    "00000000", -- 4749 - 0x128d  :    0 - 0x0
    "00000000", -- 4750 - 0x128e  :    0 - 0x0
    "00000000", -- 4751 - 0x128f  :    0 - 0x0
    "00000000", -- 4752 - 0x1290  :    0 - 0x0 -- Background 0x29
    "00111100", -- 4753 - 0x1291  :   60 - 0x3c
    "01110000", -- 4754 - 0x1292  :  112 - 0x70
    "01110000", -- 4755 - 0x1293  :  112 - 0x70
    "00111100", -- 4756 - 0x1294  :   60 - 0x3c
    "00001100", -- 4757 - 0x1295  :   12 - 0xc
    "01111000", -- 4758 - 0x1296  :  120 - 0x78
    "00000000", -- 4759 - 0x1297  :    0 - 0x0
    "00000000", -- 4760 - 0x1298  :    0 - 0x0
    "00000000", -- 4761 - 0x1299  :    0 - 0x0
    "00000000", -- 4762 - 0x129a  :    0 - 0x0
    "00000000", -- 4763 - 0x129b  :    0 - 0x0
    "00000000", -- 4764 - 0x129c  :    0 - 0x0
    "00000000", -- 4765 - 0x129d  :    0 - 0x0
    "00000000", -- 4766 - 0x129e  :    0 - 0x0
    "00000000", -- 4767 - 0x129f  :    0 - 0x0
    "00000000", -- 4768 - 0x12a0  :    0 - 0x0 -- Background 0x2a
    "00000000", -- 4769 - 0x12a1  :    0 - 0x0
    "11000110", -- 4770 - 0x12a2  :  198 - 0xc6
    "11101110", -- 4771 - 0x12a3  :  238 - 0xee
    "00101000", -- 4772 - 0x12a4  :   40 - 0x28
    "00101000", -- 4773 - 0x12a5  :   40 - 0x28
    "00101000", -- 4774 - 0x12a6  :   40 - 0x28
    "00101000", -- 4775 - 0x12a7  :   40 - 0x28
    "00000000", -- 4776 - 0x12a8  :    0 - 0x0
    "00000000", -- 4777 - 0x12a9  :    0 - 0x0
    "00000000", -- 4778 - 0x12aa  :    0 - 0x0
    "00000000", -- 4779 - 0x12ab  :    0 - 0x0
    "00000000", -- 4780 - 0x12ac  :    0 - 0x0
    "00000000", -- 4781 - 0x12ad  :    0 - 0x0
    "00000000", -- 4782 - 0x12ae  :    0 - 0x0
    "00000000", -- 4783 - 0x12af  :    0 - 0x0
    "00001000", -- 4784 - 0x12b0  :    8 - 0x8 -- Background 0x2b
    "00001000", -- 4785 - 0x12b1  :    8 - 0x8
    "00001000", -- 4786 - 0x12b2  :    8 - 0x8
    "00001000", -- 4787 - 0x12b3  :    8 - 0x8
    "00001110", -- 4788 - 0x12b4  :   14 - 0xe
    "00000110", -- 4789 - 0x12b5  :    6 - 0x6
    "00000000", -- 4790 - 0x12b6  :    0 - 0x0
    "00000000", -- 4791 - 0x12b7  :    0 - 0x0
    "00000000", -- 4792 - 0x12b8  :    0 - 0x0
    "00000000", -- 4793 - 0x12b9  :    0 - 0x0
    "00000000", -- 4794 - 0x12ba  :    0 - 0x0
    "00000000", -- 4795 - 0x12bb  :    0 - 0x0
    "00000000", -- 4796 - 0x12bc  :    0 - 0x0
    "00000000", -- 4797 - 0x12bd  :    0 - 0x0
    "00000000", -- 4798 - 0x12be  :    0 - 0x0
    "00000000", -- 4799 - 0x12bf  :    0 - 0x0
    "00101000", -- 4800 - 0x12c0  :   40 - 0x28 -- Background 0x2c
    "00101000", -- 4801 - 0x12c1  :   40 - 0x28
    "00101000", -- 4802 - 0x12c2  :   40 - 0x28
    "00101000", -- 4803 - 0x12c3  :   40 - 0x28
    "11101110", -- 4804 - 0x12c4  :  238 - 0xee
    "11000110", -- 4805 - 0x12c5  :  198 - 0xc6
    "00000000", -- 4806 - 0x12c6  :    0 - 0x0
    "00000000", -- 4807 - 0x12c7  :    0 - 0x0
    "00000000", -- 4808 - 0x12c8  :    0 - 0x0
    "00000000", -- 4809 - 0x12c9  :    0 - 0x0
    "00000000", -- 4810 - 0x12ca  :    0 - 0x0
    "00000000", -- 4811 - 0x12cb  :    0 - 0x0
    "00000000", -- 4812 - 0x12cc  :    0 - 0x0
    "00000000", -- 4813 - 0x12cd  :    0 - 0x0
    "00000000", -- 4814 - 0x12ce  :    0 - 0x0
    "00000000", -- 4815 - 0x12cf  :    0 - 0x0
    "00000000", -- 4816 - 0x12d0  :    0 - 0x0 -- Background 0x2d
    "00000000", -- 4817 - 0x12d1  :    0 - 0x0
    "01100000", -- 4818 - 0x12d2  :   96 - 0x60
    "01110000", -- 4819 - 0x12d3  :  112 - 0x70
    "00010000", -- 4820 - 0x12d4  :   16 - 0x10
    "00010000", -- 4821 - 0x12d5  :   16 - 0x10
    "00010000", -- 4822 - 0x12d6  :   16 - 0x10
    "00010000", -- 4823 - 0x12d7  :   16 - 0x10
    "00000000", -- 4824 - 0x12d8  :    0 - 0x0
    "00000000", -- 4825 - 0x12d9  :    0 - 0x0
    "00000000", -- 4826 - 0x12da  :    0 - 0x0
    "00000000", -- 4827 - 0x12db  :    0 - 0x0
    "00000000", -- 4828 - 0x12dc  :    0 - 0x0
    "00000000", -- 4829 - 0x12dd  :    0 - 0x0
    "00000000", -- 4830 - 0x12de  :    0 - 0x0
    "00000000", -- 4831 - 0x12df  :    0 - 0x0
    "00011100", -- 4832 - 0x12e0  :   28 - 0x1c -- Background 0x2e
    "00111110", -- 4833 - 0x12e1  :   62 - 0x3e
    "00111100", -- 4834 - 0x12e2  :   60 - 0x3c
    "00111000", -- 4835 - 0x12e3  :   56 - 0x38
    "00110000", -- 4836 - 0x12e4  :   48 - 0x30
    "00000000", -- 4837 - 0x12e5  :    0 - 0x0
    "01100000", -- 4838 - 0x12e6  :   96 - 0x60
    "00000000", -- 4839 - 0x12e7  :    0 - 0x0
    "00000000", -- 4840 - 0x12e8  :    0 - 0x0
    "00000000", -- 4841 - 0x12e9  :    0 - 0x0
    "00000000", -- 4842 - 0x12ea  :    0 - 0x0
    "00000000", -- 4843 - 0x12eb  :    0 - 0x0
    "00000000", -- 4844 - 0x12ec  :    0 - 0x0
    "00000000", -- 4845 - 0x12ed  :    0 - 0x0
    "00000000", -- 4846 - 0x12ee  :    0 - 0x0
    "00000000", -- 4847 - 0x12ef  :    0 - 0x0
    "00010000", -- 4848 - 0x12f0  :   16 - 0x10 -- Background 0x2f
    "00010000", -- 4849 - 0x12f1  :   16 - 0x10
    "00010000", -- 4850 - 0x12f2  :   16 - 0x10
    "00010000", -- 4851 - 0x12f3  :   16 - 0x10
    "01110000", -- 4852 - 0x12f4  :  112 - 0x70
    "01100000", -- 4853 - 0x12f5  :   96 - 0x60
    "00000000", -- 4854 - 0x12f6  :    0 - 0x0
    "00000000", -- 4855 - 0x12f7  :    0 - 0x0
    "00000000", -- 4856 - 0x12f8  :    0 - 0x0
    "00000000", -- 4857 - 0x12f9  :    0 - 0x0
    "00000000", -- 4858 - 0x12fa  :    0 - 0x0
    "00000000", -- 4859 - 0x12fb  :    0 - 0x0
    "00000000", -- 4860 - 0x12fc  :    0 - 0x0
    "00000000", -- 4861 - 0x12fd  :    0 - 0x0
    "00000000", -- 4862 - 0x12fe  :    0 - 0x0
    "00000000", -- 4863 - 0x12ff  :    0 - 0x0
    "11111111", -- 4864 - 0x1300  :  255 - 0xff -- Background 0x30
    "11111111", -- 4865 - 0x1301  :  255 - 0xff
    "00111000", -- 4866 - 0x1302  :   56 - 0x38
    "01101100", -- 4867 - 0x1303  :  108 - 0x6c
    "11000110", -- 4868 - 0x1304  :  198 - 0xc6
    "10000011", -- 4869 - 0x1305  :  131 - 0x83
    "11111111", -- 4870 - 0x1306  :  255 - 0xff
    "11111111", -- 4871 - 0x1307  :  255 - 0xff
    "00000000", -- 4872 - 0x1308  :    0 - 0x0
    "00000000", -- 4873 - 0x1309  :    0 - 0x0
    "00000000", -- 4874 - 0x130a  :    0 - 0x0
    "00000000", -- 4875 - 0x130b  :    0 - 0x0
    "00000000", -- 4876 - 0x130c  :    0 - 0x0
    "00000000", -- 4877 - 0x130d  :    0 - 0x0
    "00000000", -- 4878 - 0x130e  :    0 - 0x0
    "00000000", -- 4879 - 0x130f  :    0 - 0x0
    "11111111", -- 4880 - 0x1310  :  255 - 0xff -- Background 0x31
    "00111000", -- 4881 - 0x1311  :   56 - 0x38
    "01101100", -- 4882 - 0x1312  :  108 - 0x6c
    "11000110", -- 4883 - 0x1313  :  198 - 0xc6
    "10000011", -- 4884 - 0x1314  :  131 - 0x83
    "11111111", -- 4885 - 0x1315  :  255 - 0xff
    "11111111", -- 4886 - 0x1316  :  255 - 0xff
    "00000000", -- 4887 - 0x1317  :    0 - 0x0
    "00000000", -- 4888 - 0x1318  :    0 - 0x0
    "00000000", -- 4889 - 0x1319  :    0 - 0x0
    "00000000", -- 4890 - 0x131a  :    0 - 0x0
    "00000000", -- 4891 - 0x131b  :    0 - 0x0
    "00000000", -- 4892 - 0x131c  :    0 - 0x0
    "00000000", -- 4893 - 0x131d  :    0 - 0x0
    "00000000", -- 4894 - 0x131e  :    0 - 0x0
    "00000000", -- 4895 - 0x131f  :    0 - 0x0
    "00111000", -- 4896 - 0x1320  :   56 - 0x38 -- Background 0x32
    "01101100", -- 4897 - 0x1321  :  108 - 0x6c
    "11000110", -- 4898 - 0x1322  :  198 - 0xc6
    "10000011", -- 4899 - 0x1323  :  131 - 0x83
    "11111111", -- 4900 - 0x1324  :  255 - 0xff
    "11111111", -- 4901 - 0x1325  :  255 - 0xff
    "00000000", -- 4902 - 0x1326  :    0 - 0x0
    "00000000", -- 4903 - 0x1327  :    0 - 0x0
    "00000000", -- 4904 - 0x1328  :    0 - 0x0
    "00000000", -- 4905 - 0x1329  :    0 - 0x0
    "00000000", -- 4906 - 0x132a  :    0 - 0x0
    "00000000", -- 4907 - 0x132b  :    0 - 0x0
    "00000000", -- 4908 - 0x132c  :    0 - 0x0
    "00000000", -- 4909 - 0x132d  :    0 - 0x0
    "00000000", -- 4910 - 0x132e  :    0 - 0x0
    "00000000", -- 4911 - 0x132f  :    0 - 0x0
    "01101100", -- 4912 - 0x1330  :  108 - 0x6c -- Background 0x33
    "11000110", -- 4913 - 0x1331  :  198 - 0xc6
    "10000011", -- 4914 - 0x1332  :  131 - 0x83
    "11111111", -- 4915 - 0x1333  :  255 - 0xff
    "11111111", -- 4916 - 0x1334  :  255 - 0xff
    "00000000", -- 4917 - 0x1335  :    0 - 0x0
    "00000000", -- 4918 - 0x1336  :    0 - 0x0
    "00000000", -- 4919 - 0x1337  :    0 - 0x0
    "00000000", -- 4920 - 0x1338  :    0 - 0x0
    "00000000", -- 4921 - 0x1339  :    0 - 0x0
    "00000000", -- 4922 - 0x133a  :    0 - 0x0
    "00000000", -- 4923 - 0x133b  :    0 - 0x0
    "00000000", -- 4924 - 0x133c  :    0 - 0x0
    "00000000", -- 4925 - 0x133d  :    0 - 0x0
    "00000000", -- 4926 - 0x133e  :    0 - 0x0
    "00000000", -- 4927 - 0x133f  :    0 - 0x0
    "11000110", -- 4928 - 0x1340  :  198 - 0xc6 -- Background 0x34
    "10000011", -- 4929 - 0x1341  :  131 - 0x83
    "11111111", -- 4930 - 0x1342  :  255 - 0xff
    "11111111", -- 4931 - 0x1343  :  255 - 0xff
    "00000000", -- 4932 - 0x1344  :    0 - 0x0
    "00000000", -- 4933 - 0x1345  :    0 - 0x0
    "00000000", -- 4934 - 0x1346  :    0 - 0x0
    "00000000", -- 4935 - 0x1347  :    0 - 0x0
    "00000000", -- 4936 - 0x1348  :    0 - 0x0
    "00000000", -- 4937 - 0x1349  :    0 - 0x0
    "00000000", -- 4938 - 0x134a  :    0 - 0x0
    "00000000", -- 4939 - 0x134b  :    0 - 0x0
    "00000000", -- 4940 - 0x134c  :    0 - 0x0
    "00000000", -- 4941 - 0x134d  :    0 - 0x0
    "00000000", -- 4942 - 0x134e  :    0 - 0x0
    "00000000", -- 4943 - 0x134f  :    0 - 0x0
    "10000011", -- 4944 - 0x1350  :  131 - 0x83 -- Background 0x35
    "11111111", -- 4945 - 0x1351  :  255 - 0xff
    "11111111", -- 4946 - 0x1352  :  255 - 0xff
    "00000000", -- 4947 - 0x1353  :    0 - 0x0
    "00000000", -- 4948 - 0x1354  :    0 - 0x0
    "00000000", -- 4949 - 0x1355  :    0 - 0x0
    "00000000", -- 4950 - 0x1356  :    0 - 0x0
    "00000000", -- 4951 - 0x1357  :    0 - 0x0
    "00000000", -- 4952 - 0x1358  :    0 - 0x0
    "00000000", -- 4953 - 0x1359  :    0 - 0x0
    "00000000", -- 4954 - 0x135a  :    0 - 0x0
    "00000000", -- 4955 - 0x135b  :    0 - 0x0
    "00000000", -- 4956 - 0x135c  :    0 - 0x0
    "00000000", -- 4957 - 0x135d  :    0 - 0x0
    "00000000", -- 4958 - 0x135e  :    0 - 0x0
    "00000000", -- 4959 - 0x135f  :    0 - 0x0
    "11111111", -- 4960 - 0x1360  :  255 - 0xff -- Background 0x36
    "11111111", -- 4961 - 0x1361  :  255 - 0xff
    "00000000", -- 4962 - 0x1362  :    0 - 0x0
    "00000000", -- 4963 - 0x1363  :    0 - 0x0
    "00000000", -- 4964 - 0x1364  :    0 - 0x0
    "00000000", -- 4965 - 0x1365  :    0 - 0x0
    "00000000", -- 4966 - 0x1366  :    0 - 0x0
    "00000000", -- 4967 - 0x1367  :    0 - 0x0
    "00000000", -- 4968 - 0x1368  :    0 - 0x0
    "00000000", -- 4969 - 0x1369  :    0 - 0x0
    "00000000", -- 4970 - 0x136a  :    0 - 0x0
    "00000000", -- 4971 - 0x136b  :    0 - 0x0
    "00000000", -- 4972 - 0x136c  :    0 - 0x0
    "00000000", -- 4973 - 0x136d  :    0 - 0x0
    "00000000", -- 4974 - 0x136e  :    0 - 0x0
    "00000000", -- 4975 - 0x136f  :    0 - 0x0
    "11111111", -- 4976 - 0x1370  :  255 - 0xff -- Background 0x37
    "00000000", -- 4977 - 0x1371  :    0 - 0x0
    "00000000", -- 4978 - 0x1372  :    0 - 0x0
    "00000000", -- 4979 - 0x1373  :    0 - 0x0
    "00000000", -- 4980 - 0x1374  :    0 - 0x0
    "00000000", -- 4981 - 0x1375  :    0 - 0x0
    "00000000", -- 4982 - 0x1376  :    0 - 0x0
    "00000000", -- 4983 - 0x1377  :    0 - 0x0
    "00000000", -- 4984 - 0x1378  :    0 - 0x0
    "00000000", -- 4985 - 0x1379  :    0 - 0x0
    "00000000", -- 4986 - 0x137a  :    0 - 0x0
    "00000000", -- 4987 - 0x137b  :    0 - 0x0
    "00000000", -- 4988 - 0x137c  :    0 - 0x0
    "00000000", -- 4989 - 0x137d  :    0 - 0x0
    "00000000", -- 4990 - 0x137e  :    0 - 0x0
    "00000000", -- 4991 - 0x137f  :    0 - 0x0
    "00000000", -- 4992 - 0x1380  :    0 - 0x0 -- Background 0x38
    "00000000", -- 4993 - 0x1381  :    0 - 0x0
    "00000000", -- 4994 - 0x1382  :    0 - 0x0
    "00000000", -- 4995 - 0x1383  :    0 - 0x0
    "00000000", -- 4996 - 0x1384  :    0 - 0x0
    "00000000", -- 4997 - 0x1385  :    0 - 0x0
    "00000000", -- 4998 - 0x1386  :    0 - 0x0
    "11111111", -- 4999 - 0x1387  :  255 - 0xff
    "00000000", -- 5000 - 0x1388  :    0 - 0x0
    "00000000", -- 5001 - 0x1389  :    0 - 0x0
    "00000000", -- 5002 - 0x138a  :    0 - 0x0
    "00000000", -- 5003 - 0x138b  :    0 - 0x0
    "00000000", -- 5004 - 0x138c  :    0 - 0x0
    "00000000", -- 5005 - 0x138d  :    0 - 0x0
    "00000000", -- 5006 - 0x138e  :    0 - 0x0
    "00000000", -- 5007 - 0x138f  :    0 - 0x0
    "00000000", -- 5008 - 0x1390  :    0 - 0x0 -- Background 0x39
    "00000000", -- 5009 - 0x1391  :    0 - 0x0
    "00000000", -- 5010 - 0x1392  :    0 - 0x0
    "00000000", -- 5011 - 0x1393  :    0 - 0x0
    "00000000", -- 5012 - 0x1394  :    0 - 0x0
    "00000000", -- 5013 - 0x1395  :    0 - 0x0
    "11111111", -- 5014 - 0x1396  :  255 - 0xff
    "11111111", -- 5015 - 0x1397  :  255 - 0xff
    "00000000", -- 5016 - 0x1398  :    0 - 0x0
    "00000000", -- 5017 - 0x1399  :    0 - 0x0
    "00000000", -- 5018 - 0x139a  :    0 - 0x0
    "00000000", -- 5019 - 0x139b  :    0 - 0x0
    "00000000", -- 5020 - 0x139c  :    0 - 0x0
    "00000000", -- 5021 - 0x139d  :    0 - 0x0
    "00000000", -- 5022 - 0x139e  :    0 - 0x0
    "00000000", -- 5023 - 0x139f  :    0 - 0x0
    "00000000", -- 5024 - 0x13a0  :    0 - 0x0 -- Background 0x3a
    "00000000", -- 5025 - 0x13a1  :    0 - 0x0
    "00000000", -- 5026 - 0x13a2  :    0 - 0x0
    "00000000", -- 5027 - 0x13a3  :    0 - 0x0
    "00000000", -- 5028 - 0x13a4  :    0 - 0x0
    "11111111", -- 5029 - 0x13a5  :  255 - 0xff
    "11111111", -- 5030 - 0x13a6  :  255 - 0xff
    "00111000", -- 5031 - 0x13a7  :   56 - 0x38
    "00000000", -- 5032 - 0x13a8  :    0 - 0x0
    "00000000", -- 5033 - 0x13a9  :    0 - 0x0
    "00000000", -- 5034 - 0x13aa  :    0 - 0x0
    "00000000", -- 5035 - 0x13ab  :    0 - 0x0
    "00000000", -- 5036 - 0x13ac  :    0 - 0x0
    "00000000", -- 5037 - 0x13ad  :    0 - 0x0
    "00000000", -- 5038 - 0x13ae  :    0 - 0x0
    "00000000", -- 5039 - 0x13af  :    0 - 0x0
    "00000000", -- 5040 - 0x13b0  :    0 - 0x0 -- Background 0x3b
    "00000000", -- 5041 - 0x13b1  :    0 - 0x0
    "00000000", -- 5042 - 0x13b2  :    0 - 0x0
    "00000000", -- 5043 - 0x13b3  :    0 - 0x0
    "11111111", -- 5044 - 0x13b4  :  255 - 0xff
    "11111111", -- 5045 - 0x13b5  :  255 - 0xff
    "00111000", -- 5046 - 0x13b6  :   56 - 0x38
    "01101100", -- 5047 - 0x13b7  :  108 - 0x6c
    "00000000", -- 5048 - 0x13b8  :    0 - 0x0
    "00000000", -- 5049 - 0x13b9  :    0 - 0x0
    "00000000", -- 5050 - 0x13ba  :    0 - 0x0
    "00000000", -- 5051 - 0x13bb  :    0 - 0x0
    "00000000", -- 5052 - 0x13bc  :    0 - 0x0
    "00000000", -- 5053 - 0x13bd  :    0 - 0x0
    "00000000", -- 5054 - 0x13be  :    0 - 0x0
    "00000000", -- 5055 - 0x13bf  :    0 - 0x0
    "00000000", -- 5056 - 0x13c0  :    0 - 0x0 -- Background 0x3c
    "00000000", -- 5057 - 0x13c1  :    0 - 0x0
    "00000000", -- 5058 - 0x13c2  :    0 - 0x0
    "11111111", -- 5059 - 0x13c3  :  255 - 0xff
    "11111111", -- 5060 - 0x13c4  :  255 - 0xff
    "00111000", -- 5061 - 0x13c5  :   56 - 0x38
    "01101100", -- 5062 - 0x13c6  :  108 - 0x6c
    "11000110", -- 5063 - 0x13c7  :  198 - 0xc6
    "00000000", -- 5064 - 0x13c8  :    0 - 0x0
    "00000000", -- 5065 - 0x13c9  :    0 - 0x0
    "00000000", -- 5066 - 0x13ca  :    0 - 0x0
    "00000000", -- 5067 - 0x13cb  :    0 - 0x0
    "00000000", -- 5068 - 0x13cc  :    0 - 0x0
    "00000000", -- 5069 - 0x13cd  :    0 - 0x0
    "00000000", -- 5070 - 0x13ce  :    0 - 0x0
    "00000000", -- 5071 - 0x13cf  :    0 - 0x0
    "00000000", -- 5072 - 0x13d0  :    0 - 0x0 -- Background 0x3d
    "00000000", -- 5073 - 0x13d1  :    0 - 0x0
    "11111111", -- 5074 - 0x13d2  :  255 - 0xff
    "11111111", -- 5075 - 0x13d3  :  255 - 0xff
    "00111000", -- 5076 - 0x13d4  :   56 - 0x38
    "01101100", -- 5077 - 0x13d5  :  108 - 0x6c
    "11000110", -- 5078 - 0x13d6  :  198 - 0xc6
    "10000011", -- 5079 - 0x13d7  :  131 - 0x83
    "00000000", -- 5080 - 0x13d8  :    0 - 0x0
    "00000000", -- 5081 - 0x13d9  :    0 - 0x0
    "00000000", -- 5082 - 0x13da  :    0 - 0x0
    "00000000", -- 5083 - 0x13db  :    0 - 0x0
    "00000000", -- 5084 - 0x13dc  :    0 - 0x0
    "00000000", -- 5085 - 0x13dd  :    0 - 0x0
    "00000000", -- 5086 - 0x13de  :    0 - 0x0
    "00000000", -- 5087 - 0x13df  :    0 - 0x0
    "00000000", -- 5088 - 0x13e0  :    0 - 0x0 -- Background 0x3e
    "11111111", -- 5089 - 0x13e1  :  255 - 0xff
    "11111111", -- 5090 - 0x13e2  :  255 - 0xff
    "00111000", -- 5091 - 0x13e3  :   56 - 0x38
    "01101100", -- 5092 - 0x13e4  :  108 - 0x6c
    "11000110", -- 5093 - 0x13e5  :  198 - 0xc6
    "10000011", -- 5094 - 0x13e6  :  131 - 0x83
    "11111111", -- 5095 - 0x13e7  :  255 - 0xff
    "00000000", -- 5096 - 0x13e8  :    0 - 0x0
    "00000000", -- 5097 - 0x13e9  :    0 - 0x0
    "00000000", -- 5098 - 0x13ea  :    0 - 0x0
    "00000000", -- 5099 - 0x13eb  :    0 - 0x0
    "00000000", -- 5100 - 0x13ec  :    0 - 0x0
    "00000000", -- 5101 - 0x13ed  :    0 - 0x0
    "00000000", -- 5102 - 0x13ee  :    0 - 0x0
    "00000000", -- 5103 - 0x13ef  :    0 - 0x0
    "00000000", -- 5104 - 0x13f0  :    0 - 0x0 -- Background 0x3f
    "00000000", -- 5105 - 0x13f1  :    0 - 0x0
    "00000000", -- 5106 - 0x13f2  :    0 - 0x0
    "00000000", -- 5107 - 0x13f3  :    0 - 0x0
    "00000000", -- 5108 - 0x13f4  :    0 - 0x0
    "00000000", -- 5109 - 0x13f5  :    0 - 0x0
    "00000000", -- 5110 - 0x13f6  :    0 - 0x0
    "00000000", -- 5111 - 0x13f7  :    0 - 0x0
    "10000001", -- 5112 - 0x13f8  :  129 - 0x81
    "11111111", -- 5113 - 0x13f9  :  255 - 0xff
    "10000001", -- 5114 - 0x13fa  :  129 - 0x81
    "10000001", -- 5115 - 0x13fb  :  129 - 0x81
    "10000001", -- 5116 - 0x13fc  :  129 - 0x81
    "11111111", -- 5117 - 0x13fd  :  255 - 0xff
    "10000001", -- 5118 - 0x13fe  :  129 - 0x81
    "10000001", -- 5119 - 0x13ff  :  129 - 0x81
    "00000000", -- 5120 - 0x1400  :    0 - 0x0 -- Background 0x40
    "00000000", -- 5121 - 0x1401  :    0 - 0x0
    "00000000", -- 5122 - 0x1402  :    0 - 0x0
    "00000000", -- 5123 - 0x1403  :    0 - 0x0
    "00000000", -- 5124 - 0x1404  :    0 - 0x0
    "00000000", -- 5125 - 0x1405  :    0 - 0x0
    "00000000", -- 5126 - 0x1406  :    0 - 0x0
    "11111111", -- 5127 - 0x1407  :  255 - 0xff
    "10000001", -- 5128 - 0x1408  :  129 - 0x81
    "11111111", -- 5129 - 0x1409  :  255 - 0xff
    "10000001", -- 5130 - 0x140a  :  129 - 0x81
    "10000001", -- 5131 - 0x140b  :  129 - 0x81
    "10000001", -- 5132 - 0x140c  :  129 - 0x81
    "11111111", -- 5133 - 0x140d  :  255 - 0xff
    "10000001", -- 5134 - 0x140e  :  129 - 0x81
    "00000000", -- 5135 - 0x140f  :    0 - 0x0
    "00000000", -- 5136 - 0x1410  :    0 - 0x0 -- Background 0x41
    "00000000", -- 5137 - 0x1411  :    0 - 0x0
    "00000000", -- 5138 - 0x1412  :    0 - 0x0
    "00000000", -- 5139 - 0x1413  :    0 - 0x0
    "00000000", -- 5140 - 0x1414  :    0 - 0x0
    "11111111", -- 5141 - 0x1415  :  255 - 0xff
    "11111111", -- 5142 - 0x1416  :  255 - 0xff
    "00111000", -- 5143 - 0x1417  :   56 - 0x38
    "10000001", -- 5144 - 0x1418  :  129 - 0x81
    "11111111", -- 5145 - 0x1419  :  255 - 0xff
    "10000001", -- 5146 - 0x141a  :  129 - 0x81
    "10000001", -- 5147 - 0x141b  :  129 - 0x81
    "10000001", -- 5148 - 0x141c  :  129 - 0x81
    "00000000", -- 5149 - 0x141d  :    0 - 0x0
    "00000000", -- 5150 - 0x141e  :    0 - 0x0
    "00000000", -- 5151 - 0x141f  :    0 - 0x0
    "00000000", -- 5152 - 0x1420  :    0 - 0x0 -- Background 0x42
    "00000000", -- 5153 - 0x1421  :    0 - 0x0
    "00000000", -- 5154 - 0x1422  :    0 - 0x0
    "00000000", -- 5155 - 0x1423  :    0 - 0x0
    "11111111", -- 5156 - 0x1424  :  255 - 0xff
    "11111111", -- 5157 - 0x1425  :  255 - 0xff
    "00111000", -- 5158 - 0x1426  :   56 - 0x38
    "01101100", -- 5159 - 0x1427  :  108 - 0x6c
    "10000001", -- 5160 - 0x1428  :  129 - 0x81
    "11111111", -- 5161 - 0x1429  :  255 - 0xff
    "10000001", -- 5162 - 0x142a  :  129 - 0x81
    "10000001", -- 5163 - 0x142b  :  129 - 0x81
    "00000000", -- 5164 - 0x142c  :    0 - 0x0
    "00000000", -- 5165 - 0x142d  :    0 - 0x0
    "00000000", -- 5166 - 0x142e  :    0 - 0x0
    "00000000", -- 5167 - 0x142f  :    0 - 0x0
    "00000000", -- 5168 - 0x1430  :    0 - 0x0 -- Background 0x43
    "00000000", -- 5169 - 0x1431  :    0 - 0x0
    "00000000", -- 5170 - 0x1432  :    0 - 0x0
    "11111111", -- 5171 - 0x1433  :  255 - 0xff
    "11111111", -- 5172 - 0x1434  :  255 - 0xff
    "00111000", -- 5173 - 0x1435  :   56 - 0x38
    "01101100", -- 5174 - 0x1436  :  108 - 0x6c
    "11000110", -- 5175 - 0x1437  :  198 - 0xc6
    "10000001", -- 5176 - 0x1438  :  129 - 0x81
    "11111111", -- 5177 - 0x1439  :  255 - 0xff
    "10000001", -- 5178 - 0x143a  :  129 - 0x81
    "00000000", -- 5179 - 0x143b  :    0 - 0x0
    "00000000", -- 5180 - 0x143c  :    0 - 0x0
    "00000000", -- 5181 - 0x143d  :    0 - 0x0
    "00000000", -- 5182 - 0x143e  :    0 - 0x0
    "00000000", -- 5183 - 0x143f  :    0 - 0x0
    "00000000", -- 5184 - 0x1440  :    0 - 0x0 -- Background 0x44
    "00000000", -- 5185 - 0x1441  :    0 - 0x0
    "11111111", -- 5186 - 0x1442  :  255 - 0xff
    "11111111", -- 5187 - 0x1443  :  255 - 0xff
    "00111000", -- 5188 - 0x1444  :   56 - 0x38
    "01101100", -- 5189 - 0x1445  :  108 - 0x6c
    "11000110", -- 5190 - 0x1446  :  198 - 0xc6
    "10000011", -- 5191 - 0x1447  :  131 - 0x83
    "10000001", -- 5192 - 0x1448  :  129 - 0x81
    "11111111", -- 5193 - 0x1449  :  255 - 0xff
    "00000000", -- 5194 - 0x144a  :    0 - 0x0
    "00000000", -- 5195 - 0x144b  :    0 - 0x0
    "00000000", -- 5196 - 0x144c  :    0 - 0x0
    "00000000", -- 5197 - 0x144d  :    0 - 0x0
    "00000000", -- 5198 - 0x144e  :    0 - 0x0
    "00000000", -- 5199 - 0x144f  :    0 - 0x0
    "00000000", -- 5200 - 0x1450  :    0 - 0x0 -- Background 0x45
    "11111111", -- 5201 - 0x1451  :  255 - 0xff
    "11111111", -- 5202 - 0x1452  :  255 - 0xff
    "00111000", -- 5203 - 0x1453  :   56 - 0x38
    "01101100", -- 5204 - 0x1454  :  108 - 0x6c
    "11000110", -- 5205 - 0x1455  :  198 - 0xc6
    "10000011", -- 5206 - 0x1456  :  131 - 0x83
    "11111111", -- 5207 - 0x1457  :  255 - 0xff
    "10000001", -- 5208 - 0x1458  :  129 - 0x81
    "00000000", -- 5209 - 0x1459  :    0 - 0x0
    "00000000", -- 5210 - 0x145a  :    0 - 0x0
    "00000000", -- 5211 - 0x145b  :    0 - 0x0
    "00000000", -- 5212 - 0x145c  :    0 - 0x0
    "00000000", -- 5213 - 0x145d  :    0 - 0x0
    "00000000", -- 5214 - 0x145e  :    0 - 0x0
    "00000000", -- 5215 - 0x145f  :    0 - 0x0
    "11111111", -- 5216 - 0x1460  :  255 - 0xff -- Background 0x46
    "00111000", -- 5217 - 0x1461  :   56 - 0x38
    "01101100", -- 5218 - 0x1462  :  108 - 0x6c
    "11000110", -- 5219 - 0x1463  :  198 - 0xc6
    "10000011", -- 5220 - 0x1464  :  131 - 0x83
    "11111111", -- 5221 - 0x1465  :  255 - 0xff
    "11111111", -- 5222 - 0x1466  :  255 - 0xff
    "00000000", -- 5223 - 0x1467  :    0 - 0x0
    "00000000", -- 5224 - 0x1468  :    0 - 0x0
    "00000000", -- 5225 - 0x1469  :    0 - 0x0
    "00000000", -- 5226 - 0x146a  :    0 - 0x0
    "00000000", -- 5227 - 0x146b  :    0 - 0x0
    "00000000", -- 5228 - 0x146c  :    0 - 0x0
    "00000000", -- 5229 - 0x146d  :    0 - 0x0
    "00000000", -- 5230 - 0x146e  :    0 - 0x0
    "10000001", -- 5231 - 0x146f  :  129 - 0x81
    "00111000", -- 5232 - 0x1470  :   56 - 0x38 -- Background 0x47
    "01101100", -- 5233 - 0x1471  :  108 - 0x6c
    "11000110", -- 5234 - 0x1472  :  198 - 0xc6
    "10000011", -- 5235 - 0x1473  :  131 - 0x83
    "11111111", -- 5236 - 0x1474  :  255 - 0xff
    "11111111", -- 5237 - 0x1475  :  255 - 0xff
    "00000000", -- 5238 - 0x1476  :    0 - 0x0
    "00000000", -- 5239 - 0x1477  :    0 - 0x0
    "00000000", -- 5240 - 0x1478  :    0 - 0x0
    "00000000", -- 5241 - 0x1479  :    0 - 0x0
    "00000000", -- 5242 - 0x147a  :    0 - 0x0
    "00000000", -- 5243 - 0x147b  :    0 - 0x0
    "00000000", -- 5244 - 0x147c  :    0 - 0x0
    "00000000", -- 5245 - 0x147d  :    0 - 0x0
    "10000001", -- 5246 - 0x147e  :  129 - 0x81
    "10000001", -- 5247 - 0x147f  :  129 - 0x81
    "01101100", -- 5248 - 0x1480  :  108 - 0x6c -- Background 0x48
    "11000110", -- 5249 - 0x1481  :  198 - 0xc6
    "10000011", -- 5250 - 0x1482  :  131 - 0x83
    "11111111", -- 5251 - 0x1483  :  255 - 0xff
    "11111111", -- 5252 - 0x1484  :  255 - 0xff
    "00000000", -- 5253 - 0x1485  :    0 - 0x0
    "00000000", -- 5254 - 0x1486  :    0 - 0x0
    "00000000", -- 5255 - 0x1487  :    0 - 0x0
    "00000000", -- 5256 - 0x1488  :    0 - 0x0
    "00000000", -- 5257 - 0x1489  :    0 - 0x0
    "00000000", -- 5258 - 0x148a  :    0 - 0x0
    "00000000", -- 5259 - 0x148b  :    0 - 0x0
    "00000000", -- 5260 - 0x148c  :    0 - 0x0
    "11111111", -- 5261 - 0x148d  :  255 - 0xff
    "10000001", -- 5262 - 0x148e  :  129 - 0x81
    "10000001", -- 5263 - 0x148f  :  129 - 0x81
    "11000110", -- 5264 - 0x1490  :  198 - 0xc6 -- Background 0x49
    "10000011", -- 5265 - 0x1491  :  131 - 0x83
    "11111111", -- 5266 - 0x1492  :  255 - 0xff
    "11111111", -- 5267 - 0x1493  :  255 - 0xff
    "00000000", -- 5268 - 0x1494  :    0 - 0x0
    "00000000", -- 5269 - 0x1495  :    0 - 0x0
    "00000000", -- 5270 - 0x1496  :    0 - 0x0
    "00000000", -- 5271 - 0x1497  :    0 - 0x0
    "00000000", -- 5272 - 0x1498  :    0 - 0x0
    "00000000", -- 5273 - 0x1499  :    0 - 0x0
    "00000000", -- 5274 - 0x149a  :    0 - 0x0
    "00000000", -- 5275 - 0x149b  :    0 - 0x0
    "10000001", -- 5276 - 0x149c  :  129 - 0x81
    "11111111", -- 5277 - 0x149d  :  255 - 0xff
    "10000001", -- 5278 - 0x149e  :  129 - 0x81
    "10000001", -- 5279 - 0x149f  :  129 - 0x81
    "10000011", -- 5280 - 0x14a0  :  131 - 0x83 -- Background 0x4a
    "11111111", -- 5281 - 0x14a1  :  255 - 0xff
    "11111111", -- 5282 - 0x14a2  :  255 - 0xff
    "00000000", -- 5283 - 0x14a3  :    0 - 0x0
    "00000000", -- 5284 - 0x14a4  :    0 - 0x0
    "00000000", -- 5285 - 0x14a5  :    0 - 0x0
    "00000000", -- 5286 - 0x14a6  :    0 - 0x0
    "00000000", -- 5287 - 0x14a7  :    0 - 0x0
    "00000000", -- 5288 - 0x14a8  :    0 - 0x0
    "00000000", -- 5289 - 0x14a9  :    0 - 0x0
    "00000000", -- 5290 - 0x14aa  :    0 - 0x0
    "10000001", -- 5291 - 0x14ab  :  129 - 0x81
    "10000001", -- 5292 - 0x14ac  :  129 - 0x81
    "11111111", -- 5293 - 0x14ad  :  255 - 0xff
    "10000001", -- 5294 - 0x14ae  :  129 - 0x81
    "10000001", -- 5295 - 0x14af  :  129 - 0x81
    "11111111", -- 5296 - 0x14b0  :  255 - 0xff -- Background 0x4b
    "11111111", -- 5297 - 0x14b1  :  255 - 0xff
    "00000000", -- 5298 - 0x14b2  :    0 - 0x0
    "00000000", -- 5299 - 0x14b3  :    0 - 0x0
    "00000000", -- 5300 - 0x14b4  :    0 - 0x0
    "00000000", -- 5301 - 0x14b5  :    0 - 0x0
    "00000000", -- 5302 - 0x14b6  :    0 - 0x0
    "00000000", -- 5303 - 0x14b7  :    0 - 0x0
    "00000000", -- 5304 - 0x14b8  :    0 - 0x0
    "00000000", -- 5305 - 0x14b9  :    0 - 0x0
    "10000001", -- 5306 - 0x14ba  :  129 - 0x81
    "10000001", -- 5307 - 0x14bb  :  129 - 0x81
    "10000001", -- 5308 - 0x14bc  :  129 - 0x81
    "11111111", -- 5309 - 0x14bd  :  255 - 0xff
    "10000001", -- 5310 - 0x14be  :  129 - 0x81
    "10000001", -- 5311 - 0x14bf  :  129 - 0x81
    "10111111", -- 5312 - 0x14c0  :  191 - 0xbf -- Background 0x4c
    "01011111", -- 5313 - 0x14c1  :   95 - 0x5f
    "01011111", -- 5314 - 0x14c2  :   95 - 0x5f
    "01011111", -- 5315 - 0x14c3  :   95 - 0x5f
    "00000000", -- 5316 - 0x14c4  :    0 - 0x0
    "01011111", -- 5317 - 0x14c5  :   95 - 0x5f
    "01010001", -- 5318 - 0x14c6  :   81 - 0x51
    "01010101", -- 5319 - 0x14c7  :   85 - 0x55
    "11111111", -- 5320 - 0x14c8  :  255 - 0xff
    "01111111", -- 5321 - 0x14c9  :  127 - 0x7f
    "01111111", -- 5322 - 0x14ca  :  127 - 0x7f
    "01111111", -- 5323 - 0x14cb  :  127 - 0x7f
    "01111111", -- 5324 - 0x14cc  :  127 - 0x7f
    "01111111", -- 5325 - 0x14cd  :  127 - 0x7f
    "01111111", -- 5326 - 0x14ce  :  127 - 0x7f
    "01111111", -- 5327 - 0x14cf  :  127 - 0x7f
    "01010001", -- 5328 - 0x14d0  :   81 - 0x51 -- Background 0x4d
    "01011111", -- 5329 - 0x14d1  :   95 - 0x5f
    "00000000", -- 5330 - 0x14d2  :    0 - 0x0
    "01011111", -- 5331 - 0x14d3  :   95 - 0x5f
    "01011111", -- 5332 - 0x14d4  :   95 - 0x5f
    "01011111", -- 5333 - 0x14d5  :   95 - 0x5f
    "01011111", -- 5334 - 0x14d6  :   95 - 0x5f
    "10111111", -- 5335 - 0x14d7  :  191 - 0xbf
    "01111111", -- 5336 - 0x14d8  :  127 - 0x7f
    "01111111", -- 5337 - 0x14d9  :  127 - 0x7f
    "01111111", -- 5338 - 0x14da  :  127 - 0x7f
    "01111111", -- 5339 - 0x14db  :  127 - 0x7f
    "01110010", -- 5340 - 0x14dc  :  114 - 0x72
    "01111111", -- 5341 - 0x14dd  :  127 - 0x7f
    "01111111", -- 5342 - 0x14de  :  127 - 0x7f
    "11111111", -- 5343 - 0x14df  :  255 - 0xff
    "11111111", -- 5344 - 0x14e0  :  255 - 0xff -- Background 0x4e
    "11111110", -- 5345 - 0x14e1  :  254 - 0xfe
    "11111110", -- 5346 - 0x14e2  :  254 - 0xfe
    "11111110", -- 5347 - 0x14e3  :  254 - 0xfe
    "00000000", -- 5348 - 0x14e4  :    0 - 0x0
    "11111110", -- 5349 - 0x14e5  :  254 - 0xfe
    "00100110", -- 5350 - 0x14e6  :   38 - 0x26
    "00100110", -- 5351 - 0x14e7  :   38 - 0x26
    "11111111", -- 5352 - 0x14e8  :  255 - 0xff
    "11111110", -- 5353 - 0x14e9  :  254 - 0xfe
    "11111110", -- 5354 - 0x14ea  :  254 - 0xfe
    "11111110", -- 5355 - 0x14eb  :  254 - 0xfe
    "11111110", -- 5356 - 0x14ec  :  254 - 0xfe
    "11111110", -- 5357 - 0x14ed  :  254 - 0xfe
    "11111110", -- 5358 - 0x14ee  :  254 - 0xfe
    "11111110", -- 5359 - 0x14ef  :  254 - 0xfe
    "00100010", -- 5360 - 0x14f0  :   34 - 0x22 -- Background 0x4f
    "11111110", -- 5361 - 0x14f1  :  254 - 0xfe
    "00000000", -- 5362 - 0x14f2  :    0 - 0x0
    "11111110", -- 5363 - 0x14f3  :  254 - 0xfe
    "11111110", -- 5364 - 0x14f4  :  254 - 0xfe
    "11111110", -- 5365 - 0x14f5  :  254 - 0xfe
    "11111110", -- 5366 - 0x14f6  :  254 - 0xfe
    "11111111", -- 5367 - 0x14f7  :  255 - 0xff
    "11111110", -- 5368 - 0x14f8  :  254 - 0xfe
    "11111110", -- 5369 - 0x14f9  :  254 - 0xfe
    "11111110", -- 5370 - 0x14fa  :  254 - 0xfe
    "11111110", -- 5371 - 0x14fb  :  254 - 0xfe
    "01001010", -- 5372 - 0x14fc  :   74 - 0x4a
    "11111110", -- 5373 - 0x14fd  :  254 - 0xfe
    "11111110", -- 5374 - 0x14fe  :  254 - 0xfe
    "11111111", -- 5375 - 0x14ff  :  255 - 0xff
    "00000111", -- 5376 - 0x1500  :    7 - 0x7 -- Background 0x50
    "00000000", -- 5377 - 0x1501  :    0 - 0x0
    "00001111", -- 5378 - 0x1502  :   15 - 0xf
    "00011111", -- 5379 - 0x1503  :   31 - 0x1f
    "00011111", -- 5380 - 0x1504  :   31 - 0x1f
    "00011111", -- 5381 - 0x1505  :   31 - 0x1f
    "00011111", -- 5382 - 0x1506  :   31 - 0x1f
    "00011111", -- 5383 - 0x1507  :   31 - 0x1f
    "00000101", -- 5384 - 0x1508  :    5 - 0x5
    "00001111", -- 5385 - 0x1509  :   15 - 0xf
    "00001011", -- 5386 - 0x150a  :   11 - 0xb
    "00011011", -- 5387 - 0x150b  :   27 - 0x1b
    "00010011", -- 5388 - 0x150c  :   19 - 0x13
    "00010011", -- 5389 - 0x150d  :   19 - 0x13
    "00010011", -- 5390 - 0x150e  :   19 - 0x13
    "00010011", -- 5391 - 0x150f  :   19 - 0x13
    "00011111", -- 5392 - 0x1510  :   31 - 0x1f -- Background 0x51
    "00011111", -- 5393 - 0x1511  :   31 - 0x1f
    "00011111", -- 5394 - 0x1512  :   31 - 0x1f
    "00011111", -- 5395 - 0x1513  :   31 - 0x1f
    "00011111", -- 5396 - 0x1514  :   31 - 0x1f
    "00001111", -- 5397 - 0x1515  :   15 - 0xf
    "00000000", -- 5398 - 0x1516  :    0 - 0x0
    "00000111", -- 5399 - 0x1517  :    7 - 0x7
    "00010011", -- 5400 - 0x1518  :   19 - 0x13
    "00010011", -- 5401 - 0x1519  :   19 - 0x13
    "00010011", -- 5402 - 0x151a  :   19 - 0x13
    "00010011", -- 5403 - 0x151b  :   19 - 0x13
    "00011011", -- 5404 - 0x151c  :   27 - 0x1b
    "00001011", -- 5405 - 0x151d  :   11 - 0xb
    "00001111", -- 5406 - 0x151e  :   15 - 0xf
    "00000101", -- 5407 - 0x151f  :    5 - 0x5
    "00000111", -- 5408 - 0x1520  :    7 - 0x7 -- Background 0x52
    "00000000", -- 5409 - 0x1521  :    0 - 0x0
    "00001111", -- 5410 - 0x1522  :   15 - 0xf
    "00011111", -- 5411 - 0x1523  :   31 - 0x1f
    "00011111", -- 5412 - 0x1524  :   31 - 0x1f
    "00011111", -- 5413 - 0x1525  :   31 - 0x1f
    "00011111", -- 5414 - 0x1526  :   31 - 0x1f
    "00011111", -- 5415 - 0x1527  :   31 - 0x1f
    "00000101", -- 5416 - 0x1528  :    5 - 0x5
    "00001111", -- 5417 - 0x1529  :   15 - 0xf
    "00001011", -- 5418 - 0x152a  :   11 - 0xb
    "00011011", -- 5419 - 0x152b  :   27 - 0x1b
    "00010011", -- 5420 - 0x152c  :   19 - 0x13
    "00010011", -- 5421 - 0x152d  :   19 - 0x13
    "00010011", -- 5422 - 0x152e  :   19 - 0x13
    "00010011", -- 5423 - 0x152f  :   19 - 0x13
    "00011111", -- 5424 - 0x1530  :   31 - 0x1f -- Background 0x53
    "00011111", -- 5425 - 0x1531  :   31 - 0x1f
    "00011111", -- 5426 - 0x1532  :   31 - 0x1f
    "00011111", -- 5427 - 0x1533  :   31 - 0x1f
    "00011111", -- 5428 - 0x1534  :   31 - 0x1f
    "00001111", -- 5429 - 0x1535  :   15 - 0xf
    "00000000", -- 5430 - 0x1536  :    0 - 0x0
    "00000111", -- 5431 - 0x1537  :    7 - 0x7
    "00010011", -- 5432 - 0x1538  :   19 - 0x13
    "00010011", -- 5433 - 0x1539  :   19 - 0x13
    "00010011", -- 5434 - 0x153a  :   19 - 0x13
    "00010011", -- 5435 - 0x153b  :   19 - 0x13
    "00011011", -- 5436 - 0x153c  :   27 - 0x1b
    "00001011", -- 5437 - 0x153d  :   11 - 0xb
    "00001111", -- 5438 - 0x153e  :   15 - 0xf
    "00000101", -- 5439 - 0x153f  :    5 - 0x5
    "11100000", -- 5440 - 0x1540  :  224 - 0xe0 -- Background 0x54
    "00000000", -- 5441 - 0x1541  :    0 - 0x0
    "11110001", -- 5442 - 0x1542  :  241 - 0xf1
    "11111011", -- 5443 - 0x1543  :  251 - 0xfb
    "11111011", -- 5444 - 0x1544  :  251 - 0xfb
    "11111011", -- 5445 - 0x1545  :  251 - 0xfb
    "11111011", -- 5446 - 0x1546  :  251 - 0xfb
    "11111011", -- 5447 - 0x1547  :  251 - 0xfb
    "10100000", -- 5448 - 0x1548  :  160 - 0xa0
    "11110001", -- 5449 - 0x1549  :  241 - 0xf1
    "11010001", -- 5450 - 0x154a  :  209 - 0xd1
    "11011011", -- 5451 - 0x154b  :  219 - 0xdb
    "11001010", -- 5452 - 0x154c  :  202 - 0xca
    "11001010", -- 5453 - 0x154d  :  202 - 0xca
    "11001010", -- 5454 - 0x154e  :  202 - 0xca
    "11001010", -- 5455 - 0x154f  :  202 - 0xca
    "11111011", -- 5456 - 0x1550  :  251 - 0xfb -- Background 0x55
    "11111011", -- 5457 - 0x1551  :  251 - 0xfb
    "11111011", -- 5458 - 0x1552  :  251 - 0xfb
    "11111011", -- 5459 - 0x1553  :  251 - 0xfb
    "11111011", -- 5460 - 0x1554  :  251 - 0xfb
    "11110001", -- 5461 - 0x1555  :  241 - 0xf1
    "00000000", -- 5462 - 0x1556  :    0 - 0x0
    "11100000", -- 5463 - 0x1557  :  224 - 0xe0
    "11001010", -- 5464 - 0x1558  :  202 - 0xca
    "11001010", -- 5465 - 0x1559  :  202 - 0xca
    "11001010", -- 5466 - 0x155a  :  202 - 0xca
    "11001010", -- 5467 - 0x155b  :  202 - 0xca
    "11011011", -- 5468 - 0x155c  :  219 - 0xdb
    "11010001", -- 5469 - 0x155d  :  209 - 0xd1
    "11110001", -- 5470 - 0x155e  :  241 - 0xf1
    "10100000", -- 5471 - 0x155f  :  160 - 0xa0
    "11100000", -- 5472 - 0x1560  :  224 - 0xe0 -- Background 0x56
    "00000000", -- 5473 - 0x1561  :    0 - 0x0
    "11110001", -- 5474 - 0x1562  :  241 - 0xf1
    "11111011", -- 5475 - 0x1563  :  251 - 0xfb
    "11111011", -- 5476 - 0x1564  :  251 - 0xfb
    "11111011", -- 5477 - 0x1565  :  251 - 0xfb
    "11111011", -- 5478 - 0x1566  :  251 - 0xfb
    "11111011", -- 5479 - 0x1567  :  251 - 0xfb
    "10100000", -- 5480 - 0x1568  :  160 - 0xa0
    "11110001", -- 5481 - 0x1569  :  241 - 0xf1
    "11010001", -- 5482 - 0x156a  :  209 - 0xd1
    "11011011", -- 5483 - 0x156b  :  219 - 0xdb
    "11001010", -- 5484 - 0x156c  :  202 - 0xca
    "11001010", -- 5485 - 0x156d  :  202 - 0xca
    "11001010", -- 5486 - 0x156e  :  202 - 0xca
    "11001010", -- 5487 - 0x156f  :  202 - 0xca
    "11111011", -- 5488 - 0x1570  :  251 - 0xfb -- Background 0x57
    "11111011", -- 5489 - 0x1571  :  251 - 0xfb
    "11111011", -- 5490 - 0x1572  :  251 - 0xfb
    "11111011", -- 5491 - 0x1573  :  251 - 0xfb
    "11111011", -- 5492 - 0x1574  :  251 - 0xfb
    "11110001", -- 5493 - 0x1575  :  241 - 0xf1
    "00000000", -- 5494 - 0x1576  :    0 - 0x0
    "11100000", -- 5495 - 0x1577  :  224 - 0xe0
    "11001010", -- 5496 - 0x1578  :  202 - 0xca
    "11001010", -- 5497 - 0x1579  :  202 - 0xca
    "11001010", -- 5498 - 0x157a  :  202 - 0xca
    "11001010", -- 5499 - 0x157b  :  202 - 0xca
    "11011011", -- 5500 - 0x157c  :  219 - 0xdb
    "11010001", -- 5501 - 0x157d  :  209 - 0xd1
    "11110000", -- 5502 - 0x157e  :  240 - 0xf0
    "10100000", -- 5503 - 0x157f  :  160 - 0xa0
    "11111100", -- 5504 - 0x1580  :  252 - 0xfc -- Background 0x58
    "00000000", -- 5505 - 0x1581  :    0 - 0x0
    "11111110", -- 5506 - 0x1582  :  254 - 0xfe
    "11111111", -- 5507 - 0x1583  :  255 - 0xff
    "11111111", -- 5508 - 0x1584  :  255 - 0xff
    "11111111", -- 5509 - 0x1585  :  255 - 0xff
    "11111111", -- 5510 - 0x1586  :  255 - 0xff
    "11111111", -- 5511 - 0x1587  :  255 - 0xff
    "10110100", -- 5512 - 0x1588  :  180 - 0xb4
    "11111110", -- 5513 - 0x1589  :  254 - 0xfe
    "01111010", -- 5514 - 0x158a  :  122 - 0x7a
    "01111011", -- 5515 - 0x158b  :  123 - 0x7b
    "01111001", -- 5516 - 0x158c  :  121 - 0x79
    "01111001", -- 5517 - 0x158d  :  121 - 0x79
    "01111001", -- 5518 - 0x158e  :  121 - 0x79
    "01111001", -- 5519 - 0x158f  :  121 - 0x79
    "11111111", -- 5520 - 0x1590  :  255 - 0xff -- Background 0x59
    "11111111", -- 5521 - 0x1591  :  255 - 0xff
    "11111111", -- 5522 - 0x1592  :  255 - 0xff
    "11111111", -- 5523 - 0x1593  :  255 - 0xff
    "11111111", -- 5524 - 0x1594  :  255 - 0xff
    "11111110", -- 5525 - 0x1595  :  254 - 0xfe
    "00000000", -- 5526 - 0x1596  :    0 - 0x0
    "11111100", -- 5527 - 0x1597  :  252 - 0xfc
    "01111001", -- 5528 - 0x1598  :  121 - 0x79
    "01111001", -- 5529 - 0x1599  :  121 - 0x79
    "01111001", -- 5530 - 0x159a  :  121 - 0x79
    "01111001", -- 5531 - 0x159b  :  121 - 0x79
    "01111011", -- 5532 - 0x159c  :  123 - 0x7b
    "01111010", -- 5533 - 0x159d  :  122 - 0x7a
    "11111110", -- 5534 - 0x159e  :  254 - 0xfe
    "10110100", -- 5535 - 0x159f  :  180 - 0xb4
    "11111100", -- 5536 - 0x15a0  :  252 - 0xfc -- Background 0x5a
    "00000000", -- 5537 - 0x15a1  :    0 - 0x0
    "11111110", -- 5538 - 0x15a2  :  254 - 0xfe
    "11111111", -- 5539 - 0x15a3  :  255 - 0xff
    "11111111", -- 5540 - 0x15a4  :  255 - 0xff
    "11111111", -- 5541 - 0x15a5  :  255 - 0xff
    "11111111", -- 5542 - 0x15a6  :  255 - 0xff
    "11111111", -- 5543 - 0x15a7  :  255 - 0xff
    "10110100", -- 5544 - 0x15a8  :  180 - 0xb4
    "11111110", -- 5545 - 0x15a9  :  254 - 0xfe
    "01111010", -- 5546 - 0x15aa  :  122 - 0x7a
    "01111011", -- 5547 - 0x15ab  :  123 - 0x7b
    "01111001", -- 5548 - 0x15ac  :  121 - 0x79
    "01111001", -- 5549 - 0x15ad  :  121 - 0x79
    "01111001", -- 5550 - 0x15ae  :  121 - 0x79
    "01111001", -- 5551 - 0x15af  :  121 - 0x79
    "11111111", -- 5552 - 0x15b0  :  255 - 0xff -- Background 0x5b
    "11111111", -- 5553 - 0x15b1  :  255 - 0xff
    "11111111", -- 5554 - 0x15b2  :  255 - 0xff
    "11111111", -- 5555 - 0x15b3  :  255 - 0xff
    "11111111", -- 5556 - 0x15b4  :  255 - 0xff
    "11111110", -- 5557 - 0x15b5  :  254 - 0xfe
    "00000000", -- 5558 - 0x15b6  :    0 - 0x0
    "11111100", -- 5559 - 0x15b7  :  252 - 0xfc
    "01111001", -- 5560 - 0x15b8  :  121 - 0x79
    "01111001", -- 5561 - 0x15b9  :  121 - 0x79
    "01111001", -- 5562 - 0x15ba  :  121 - 0x79
    "01111001", -- 5563 - 0x15bb  :  121 - 0x79
    "01111011", -- 5564 - 0x15bc  :  123 - 0x7b
    "01111010", -- 5565 - 0x15bd  :  122 - 0x7a
    "11111110", -- 5566 - 0x15be  :  254 - 0xfe
    "10110100", -- 5567 - 0x15bf  :  180 - 0xb4
    "00000000", -- 5568 - 0x15c0  :    0 - 0x0 -- Background 0x5c
    "00000000", -- 5569 - 0x15c1  :    0 - 0x0
    "00011111", -- 5570 - 0x15c2  :   31 - 0x1f
    "00010000", -- 5571 - 0x15c3  :   16 - 0x10
    "00010000", -- 5572 - 0x15c4  :   16 - 0x10
    "00011111", -- 5573 - 0x15c5  :   31 - 0x1f
    "00000000", -- 5574 - 0x15c6  :    0 - 0x0
    "00000000", -- 5575 - 0x15c7  :    0 - 0x0
    "01111111", -- 5576 - 0x15c8  :  127 - 0x7f
    "10111111", -- 5577 - 0x15c9  :  191 - 0xbf
    "11111111", -- 5578 - 0x15ca  :  255 - 0xff
    "10110010", -- 5579 - 0x15cb  :  178 - 0xb2
    "10110001", -- 5580 - 0x15cc  :  177 - 0xb1
    "11111111", -- 5581 - 0x15cd  :  255 - 0xff
    "10111111", -- 5582 - 0x15ce  :  191 - 0xbf
    "01111111", -- 5583 - 0x15cf  :  127 - 0x7f
    "00000000", -- 5584 - 0x15d0  :    0 - 0x0 -- Background 0x5d
    "00000000", -- 5585 - 0x15d1  :    0 - 0x0
    "11111000", -- 5586 - 0x15d2  :  248 - 0xf8
    "00001000", -- 5587 - 0x15d3  :    8 - 0x8
    "00001000", -- 5588 - 0x15d4  :    8 - 0x8
    "11111000", -- 5589 - 0x15d5  :  248 - 0xf8
    "00000000", -- 5590 - 0x15d6  :    0 - 0x0
    "00000000", -- 5591 - 0x15d7  :    0 - 0x0
    "11111110", -- 5592 - 0x15d8  :  254 - 0xfe
    "11111101", -- 5593 - 0x15d9  :  253 - 0xfd
    "11111111", -- 5594 - 0x15da  :  255 - 0xff
    "11001101", -- 5595 - 0x15db  :  205 - 0xcd
    "01101101", -- 5596 - 0x15dc  :  109 - 0x6d
    "11111111", -- 5597 - 0x15dd  :  255 - 0xff
    "11111101", -- 5598 - 0x15de  :  253 - 0xfd
    "11111110", -- 5599 - 0x15df  :  254 - 0xfe
    "00000000", -- 5600 - 0x15e0  :    0 - 0x0 -- Background 0x5e
    "00000001", -- 5601 - 0x15e1  :    1 - 0x1
    "00000010", -- 5602 - 0x15e2  :    2 - 0x2
    "00000010", -- 5603 - 0x15e3  :    2 - 0x2
    "11110001", -- 5604 - 0x15e4  :  241 - 0xf1
    "00001000", -- 5605 - 0x15e5  :    8 - 0x8
    "00000100", -- 5606 - 0x15e6  :    4 - 0x4
    "00000011", -- 5607 - 0x15e7  :    3 - 0x3
    "11111111", -- 5608 - 0x15e8  :  255 - 0xff
    "11111111", -- 5609 - 0x15e9  :  255 - 0xff
    "10101110", -- 5610 - 0x15ea  :  174 - 0xae
    "11111110", -- 5611 - 0x15eb  :  254 - 0xfe
    "11111111", -- 5612 - 0x15ec  :  255 - 0xff
    "00001111", -- 5613 - 0x15ed  :   15 - 0xf
    "00000111", -- 5614 - 0x15ee  :    7 - 0x7
    "00000011", -- 5615 - 0x15ef  :    3 - 0x3
    "00000000", -- 5616 - 0x15f0  :    0 - 0x0 -- Background 0x5f
    "10000000", -- 5617 - 0x15f1  :  128 - 0x80
    "01000000", -- 5618 - 0x15f2  :   64 - 0x40
    "01000000", -- 5619 - 0x15f3  :   64 - 0x40
    "10001111", -- 5620 - 0x15f4  :  143 - 0x8f
    "00010000", -- 5621 - 0x15f5  :   16 - 0x10
    "00100000", -- 5622 - 0x15f6  :   32 - 0x20
    "11000000", -- 5623 - 0x15f7  :  192 - 0xc0
    "11111111", -- 5624 - 0x15f8  :  255 - 0xff
    "11111111", -- 5625 - 0x15f9  :  255 - 0xff
    "01110101", -- 5626 - 0x15fa  :  117 - 0x75
    "01111111", -- 5627 - 0x15fb  :  127 - 0x7f
    "11111111", -- 5628 - 0x15fc  :  255 - 0xff
    "11110000", -- 5629 - 0x15fd  :  240 - 0xf0
    "11100000", -- 5630 - 0x15fe  :  224 - 0xe0
    "11000000", -- 5631 - 0x15ff  :  192 - 0xc0
    "00000011", -- 5632 - 0x1600  :    3 - 0x3 -- Background 0x60
    "00000100", -- 5633 - 0x1601  :    4 - 0x4
    "00001000", -- 5634 - 0x1602  :    8 - 0x8
    "11110001", -- 5635 - 0x1603  :  241 - 0xf1
    "00000010", -- 5636 - 0x1604  :    2 - 0x2
    "00000010", -- 5637 - 0x1605  :    2 - 0x2
    "00000001", -- 5638 - 0x1606  :    1 - 0x1
    "00000000", -- 5639 - 0x1607  :    0 - 0x0
    "00000011", -- 5640 - 0x1608  :    3 - 0x3
    "00000111", -- 5641 - 0x1609  :    7 - 0x7
    "00001111", -- 5642 - 0x160a  :   15 - 0xf
    "11111111", -- 5643 - 0x160b  :  255 - 0xff
    "11111110", -- 5644 - 0x160c  :  254 - 0xfe
    "10101110", -- 5645 - 0x160d  :  174 - 0xae
    "11111111", -- 5646 - 0x160e  :  255 - 0xff
    "11111111", -- 5647 - 0x160f  :  255 - 0xff
    "11000000", -- 5648 - 0x1610  :  192 - 0xc0 -- Background 0x61
    "00100000", -- 5649 - 0x1611  :   32 - 0x20
    "00010000", -- 5650 - 0x1612  :   16 - 0x10
    "10001111", -- 5651 - 0x1613  :  143 - 0x8f
    "01000000", -- 5652 - 0x1614  :   64 - 0x40
    "01000000", -- 5653 - 0x1615  :   64 - 0x40
    "10000000", -- 5654 - 0x1616  :  128 - 0x80
    "00000000", -- 5655 - 0x1617  :    0 - 0x0
    "11000000", -- 5656 - 0x1618  :  192 - 0xc0
    "11100000", -- 5657 - 0x1619  :  224 - 0xe0
    "11110000", -- 5658 - 0x161a  :  240 - 0xf0
    "11111111", -- 5659 - 0x161b  :  255 - 0xff
    "01111111", -- 5660 - 0x161c  :  127 - 0x7f
    "01110101", -- 5661 - 0x161d  :  117 - 0x75
    "11111111", -- 5662 - 0x161e  :  255 - 0xff
    "11111111", -- 5663 - 0x161f  :  255 - 0xff
    "11111111", -- 5664 - 0x1620  :  255 - 0xff -- Background 0x62
    "11111111", -- 5665 - 0x1621  :  255 - 0xff
    "11000011", -- 5666 - 0x1622  :  195 - 0xc3
    "10000001", -- 5667 - 0x1623  :  129 - 0x81
    "10000001", -- 5668 - 0x1624  :  129 - 0x81
    "11000011", -- 5669 - 0x1625  :  195 - 0xc3
    "11111111", -- 5670 - 0x1626  :  255 - 0xff
    "11111111", -- 5671 - 0x1627  :  255 - 0xff
    "11111111", -- 5672 - 0x1628  :  255 - 0xff
    "00000000", -- 5673 - 0x1629  :    0 - 0x0
    "11000011", -- 5674 - 0x162a  :  195 - 0xc3
    "10000001", -- 5675 - 0x162b  :  129 - 0x81
    "10000001", -- 5676 - 0x162c  :  129 - 0x81
    "11000011", -- 5677 - 0x162d  :  195 - 0xc3
    "11111111", -- 5678 - 0x162e  :  255 - 0xff
    "00000000", -- 5679 - 0x162f  :    0 - 0x0
    "11111111", -- 5680 - 0x1630  :  255 - 0xff -- Background 0x63
    "10011001", -- 5681 - 0x1631  :  153 - 0x99
    "00000000", -- 5682 - 0x1632  :    0 - 0x0
    "00000000", -- 5683 - 0x1633  :    0 - 0x0
    "00000000", -- 5684 - 0x1634  :    0 - 0x0
    "10000001", -- 5685 - 0x1635  :  129 - 0x81
    "10000001", -- 5686 - 0x1636  :  129 - 0x81
    "10000001", -- 5687 - 0x1637  :  129 - 0x81
    "10000001", -- 5688 - 0x1638  :  129 - 0x81
    "01100110", -- 5689 - 0x1639  :  102 - 0x66
    "01111110", -- 5690 - 0x163a  :  126 - 0x7e
    "01111110", -- 5691 - 0x163b  :  126 - 0x7e
    "01111110", -- 5692 - 0x163c  :  126 - 0x7e
    "11111111", -- 5693 - 0x163d  :  255 - 0xff
    "11111111", -- 5694 - 0x163e  :  255 - 0xff
    "01111110", -- 5695 - 0x163f  :  126 - 0x7e
    "00000000", -- 5696 - 0x1640  :    0 - 0x0 -- Background 0x64
    "00000000", -- 5697 - 0x1641  :    0 - 0x0
    "00000000", -- 5698 - 0x1642  :    0 - 0x0
    "00000000", -- 5699 - 0x1643  :    0 - 0x0
    "01100000", -- 5700 - 0x1644  :   96 - 0x60
    "01100000", -- 5701 - 0x1645  :   96 - 0x60
    "00000000", -- 5702 - 0x1646  :    0 - 0x0
    "00000000", -- 5703 - 0x1647  :    0 - 0x0
    "00000000", -- 5704 - 0x1648  :    0 - 0x0
    "00000000", -- 5705 - 0x1649  :    0 - 0x0
    "00000000", -- 5706 - 0x164a  :    0 - 0x0
    "00000000", -- 5707 - 0x164b  :    0 - 0x0
    "00000000", -- 5708 - 0x164c  :    0 - 0x0
    "00000000", -- 5709 - 0x164d  :    0 - 0x0
    "00000000", -- 5710 - 0x164e  :    0 - 0x0
    "00000000", -- 5711 - 0x164f  :    0 - 0x0
    "00000000", -- 5712 - 0x1650  :    0 - 0x0 -- Background 0x65
    "00000000", -- 5713 - 0x1651  :    0 - 0x0
    "00000000", -- 5714 - 0x1652  :    0 - 0x0
    "00000000", -- 5715 - 0x1653  :    0 - 0x0
    "01101100", -- 5716 - 0x1654  :  108 - 0x6c
    "01101100", -- 5717 - 0x1655  :  108 - 0x6c
    "00001000", -- 5718 - 0x1656  :    8 - 0x8
    "00000000", -- 5719 - 0x1657  :    0 - 0x0
    "00000000", -- 5720 - 0x1658  :    0 - 0x0
    "00000000", -- 5721 - 0x1659  :    0 - 0x0
    "00000000", -- 5722 - 0x165a  :    0 - 0x0
    "00000000", -- 5723 - 0x165b  :    0 - 0x0
    "00000000", -- 5724 - 0x165c  :    0 - 0x0
    "00000000", -- 5725 - 0x165d  :    0 - 0x0
    "00000000", -- 5726 - 0x165e  :    0 - 0x0
    "00000000", -- 5727 - 0x165f  :    0 - 0x0
    "00111100", -- 5728 - 0x1660  :   60 - 0x3c -- Background 0x66
    "00011000", -- 5729 - 0x1661  :   24 - 0x18
    "00011000", -- 5730 - 0x1662  :   24 - 0x18
    "00011000", -- 5731 - 0x1663  :   24 - 0x18
    "00011000", -- 5732 - 0x1664  :   24 - 0x18
    "00011000", -- 5733 - 0x1665  :   24 - 0x18
    "00111100", -- 5734 - 0x1666  :   60 - 0x3c
    "00000000", -- 5735 - 0x1667  :    0 - 0x0
    "00000000", -- 5736 - 0x1668  :    0 - 0x0
    "00000000", -- 5737 - 0x1669  :    0 - 0x0
    "00000000", -- 5738 - 0x166a  :    0 - 0x0
    "00000000", -- 5739 - 0x166b  :    0 - 0x0
    "00000000", -- 5740 - 0x166c  :    0 - 0x0
    "00000000", -- 5741 - 0x166d  :    0 - 0x0
    "00000000", -- 5742 - 0x166e  :    0 - 0x0
    "00000000", -- 5743 - 0x166f  :    0 - 0x0
    "11111111", -- 5744 - 0x1670  :  255 - 0xff -- Background 0x67
    "01100110", -- 5745 - 0x1671  :  102 - 0x66
    "01100110", -- 5746 - 0x1672  :  102 - 0x66
    "01100110", -- 5747 - 0x1673  :  102 - 0x66
    "01100110", -- 5748 - 0x1674  :  102 - 0x66
    "01100110", -- 5749 - 0x1675  :  102 - 0x66
    "01100110", -- 5750 - 0x1676  :  102 - 0x66
    "11111111", -- 5751 - 0x1677  :  255 - 0xff
    "00000000", -- 5752 - 0x1678  :    0 - 0x0
    "00000000", -- 5753 - 0x1679  :    0 - 0x0
    "00000000", -- 5754 - 0x167a  :    0 - 0x0
    "00000000", -- 5755 - 0x167b  :    0 - 0x0
    "00000000", -- 5756 - 0x167c  :    0 - 0x0
    "00000000", -- 5757 - 0x167d  :    0 - 0x0
    "00000000", -- 5758 - 0x167e  :    0 - 0x0
    "00000000", -- 5759 - 0x167f  :    0 - 0x0
    "00000011", -- 5760 - 0x1680  :    3 - 0x3 -- Background 0x68
    "00000001", -- 5761 - 0x1681  :    1 - 0x1
    "00000000", -- 5762 - 0x1682  :    0 - 0x0
    "00000000", -- 5763 - 0x1683  :    0 - 0x0
    "00000000", -- 5764 - 0x1684  :    0 - 0x0
    "00000000", -- 5765 - 0x1685  :    0 - 0x0
    "00000000", -- 5766 - 0x1686  :    0 - 0x0
    "00000000", -- 5767 - 0x1687  :    0 - 0x0
    "00000011", -- 5768 - 0x1688  :    3 - 0x3
    "00000001", -- 5769 - 0x1689  :    1 - 0x1
    "00000000", -- 5770 - 0x168a  :    0 - 0x0
    "00000000", -- 5771 - 0x168b  :    0 - 0x0
    "00000000", -- 5772 - 0x168c  :    0 - 0x0
    "00000000", -- 5773 - 0x168d  :    0 - 0x0
    "00000000", -- 5774 - 0x168e  :    0 - 0x0
    "00000000", -- 5775 - 0x168f  :    0 - 0x0
    "10000011", -- 5776 - 0x1690  :  131 - 0x83 -- Background 0x69
    "11010001", -- 5777 - 0x1691  :  209 - 0xd1
    "11100001", -- 5778 - 0x1692  :  225 - 0xe1
    "11010001", -- 5779 - 0x1693  :  209 - 0xd1
    "00000010", -- 5780 - 0x1694  :    2 - 0x2
    "10000100", -- 5781 - 0x1695  :  132 - 0x84
    "11110000", -- 5782 - 0x1696  :  240 - 0xf0
    "11001110", -- 5783 - 0x1697  :  206 - 0xce
    "11111111", -- 5784 - 0x1698  :  255 - 0xff
    "11111111", -- 5785 - 0x1699  :  255 - 0xff
    "11111111", -- 5786 - 0x169a  :  255 - 0xff
    "11111111", -- 5787 - 0x169b  :  255 - 0xff
    "11111111", -- 5788 - 0x169c  :  255 - 0xff
    "11111111", -- 5789 - 0x169d  :  255 - 0xff
    "11111111", -- 5790 - 0x169e  :  255 - 0xff
    "11111111", -- 5791 - 0x169f  :  255 - 0xff
    "11000000", -- 5792 - 0x16a0  :  192 - 0xc0 -- Background 0x6a
    "10000000", -- 5793 - 0x16a1  :  128 - 0x80
    "00000000", -- 5794 - 0x16a2  :    0 - 0x0
    "00000000", -- 5795 - 0x16a3  :    0 - 0x0
    "00000000", -- 5796 - 0x16a4  :    0 - 0x0
    "00000000", -- 5797 - 0x16a5  :    0 - 0x0
    "00000000", -- 5798 - 0x16a6  :    0 - 0x0
    "00000000", -- 5799 - 0x16a7  :    0 - 0x0
    "11000000", -- 5800 - 0x16a8  :  192 - 0xc0
    "10000000", -- 5801 - 0x16a9  :  128 - 0x80
    "00000000", -- 5802 - 0x16aa  :    0 - 0x0
    "00000000", -- 5803 - 0x16ab  :    0 - 0x0
    "00000000", -- 5804 - 0x16ac  :    0 - 0x0
    "00000000", -- 5805 - 0x16ad  :    0 - 0x0
    "00000000", -- 5806 - 0x16ae  :    0 - 0x0
    "00000000", -- 5807 - 0x16af  :    0 - 0x0
    "11000001", -- 5808 - 0x16b0  :  193 - 0xc1 -- Background 0x6b
    "10001011", -- 5809 - 0x16b1  :  139 - 0x8b
    "10000111", -- 5810 - 0x16b2  :  135 - 0x87
    "10001011", -- 5811 - 0x16b3  :  139 - 0x8b
    "01000000", -- 5812 - 0x16b4  :   64 - 0x40
    "00100001", -- 5813 - 0x16b5  :   33 - 0x21
    "00001111", -- 5814 - 0x16b6  :   15 - 0xf
    "11010011", -- 5815 - 0x16b7  :  211 - 0xd3
    "11111111", -- 5816 - 0x16b8  :  255 - 0xff
    "11111111", -- 5817 - 0x16b9  :  255 - 0xff
    "11111111", -- 5818 - 0x16ba  :  255 - 0xff
    "11111111", -- 5819 - 0x16bb  :  255 - 0xff
    "11111111", -- 5820 - 0x16bc  :  255 - 0xff
    "11111111", -- 5821 - 0x16bd  :  255 - 0xff
    "11111111", -- 5822 - 0x16be  :  255 - 0xff
    "11111111", -- 5823 - 0x16bf  :  255 - 0xff
    "11111111", -- 5824 - 0x16c0  :  255 - 0xff -- Background 0x6c
    "11111111", -- 5825 - 0x16c1  :  255 - 0xff
    "11111111", -- 5826 - 0x16c2  :  255 - 0xff
    "00011111", -- 5827 - 0x16c3  :   31 - 0x1f
    "00001111", -- 5828 - 0x16c4  :   15 - 0xf
    "00011110", -- 5829 - 0x16c5  :   30 - 0x1e
    "00111111", -- 5830 - 0x16c6  :   63 - 0x3f
    "01111111", -- 5831 - 0x16c7  :  127 - 0x7f
    "11111111", -- 5832 - 0x16c8  :  255 - 0xff
    "11111111", -- 5833 - 0x16c9  :  255 - 0xff
    "11111111", -- 5834 - 0x16ca  :  255 - 0xff
    "00011111", -- 5835 - 0x16cb  :   31 - 0x1f
    "00011111", -- 5836 - 0x16cc  :   31 - 0x1f
    "00111111", -- 5837 - 0x16cd  :   63 - 0x3f
    "01111111", -- 5838 - 0x16ce  :  127 - 0x7f
    "11111111", -- 5839 - 0x16cf  :  255 - 0xff
    "11111111", -- 5840 - 0x16d0  :  255 - 0xff -- Background 0x6d
    "11111111", -- 5841 - 0x16d1  :  255 - 0xff
    "11111111", -- 5842 - 0x16d2  :  255 - 0xff
    "11111000", -- 5843 - 0x16d3  :  248 - 0xf8
    "11110000", -- 5844 - 0x16d4  :  240 - 0xf0
    "01111000", -- 5845 - 0x16d5  :  120 - 0x78
    "11111100", -- 5846 - 0x16d6  :  252 - 0xfc
    "11111110", -- 5847 - 0x16d7  :  254 - 0xfe
    "11111111", -- 5848 - 0x16d8  :  255 - 0xff
    "11111111", -- 5849 - 0x16d9  :  255 - 0xff
    "11111111", -- 5850 - 0x16da  :  255 - 0xff
    "11111000", -- 5851 - 0x16db  :  248 - 0xf8
    "11111000", -- 5852 - 0x16dc  :  248 - 0xf8
    "11111100", -- 5853 - 0x16dd  :  252 - 0xfc
    "11111110", -- 5854 - 0x16de  :  254 - 0xfe
    "11111111", -- 5855 - 0x16df  :  255 - 0xff
    "00000000", -- 5856 - 0x16e0  :    0 - 0x0 -- Background 0x6e
    "00000000", -- 5857 - 0x16e1  :    0 - 0x0
    "00000000", -- 5858 - 0x16e2  :    0 - 0x0
    "00000000", -- 5859 - 0x16e3  :    0 - 0x0
    "00000000", -- 5860 - 0x16e4  :    0 - 0x0
    "00111100", -- 5861 - 0x16e5  :   60 - 0x3c
    "01000010", -- 5862 - 0x16e6  :   66 - 0x42
    "10000001", -- 5863 - 0x16e7  :  129 - 0x81
    "00000000", -- 5864 - 0x16e8  :    0 - 0x0
    "00000000", -- 5865 - 0x16e9  :    0 - 0x0
    "00000000", -- 5866 - 0x16ea  :    0 - 0x0
    "00000000", -- 5867 - 0x16eb  :    0 - 0x0
    "00000000", -- 5868 - 0x16ec  :    0 - 0x0
    "00111100", -- 5869 - 0x16ed  :   60 - 0x3c
    "01000010", -- 5870 - 0x16ee  :   66 - 0x42
    "10000001", -- 5871 - 0x16ef  :  129 - 0x81
    "10000001", -- 5872 - 0x16f0  :  129 - 0x81 -- Background 0x6f
    "10111101", -- 5873 - 0x16f1  :  189 - 0xbd
    "01111110", -- 5874 - 0x16f2  :  126 - 0x7e
    "11111111", -- 5875 - 0x16f3  :  255 - 0xff
    "11100111", -- 5876 - 0x16f4  :  231 - 0xe7
    "11111111", -- 5877 - 0x16f5  :  255 - 0xff
    "11111111", -- 5878 - 0x16f6  :  255 - 0xff
    "11111111", -- 5879 - 0x16f7  :  255 - 0xff
    "10000001", -- 5880 - 0x16f8  :  129 - 0x81
    "10111101", -- 5881 - 0x16f9  :  189 - 0xbd
    "01111110", -- 5882 - 0x16fa  :  126 - 0x7e
    "10100101", -- 5883 - 0x16fb  :  165 - 0xa5
    "11011011", -- 5884 - 0x16fc  :  219 - 0xdb
    "11100111", -- 5885 - 0x16fd  :  231 - 0xe7
    "11111111", -- 5886 - 0x16fe  :  255 - 0xff
    "11111111", -- 5887 - 0x16ff  :  255 - 0xff
    "00000001", -- 5888 - 0x1700  :    1 - 0x1 -- Background 0x70
    "00000111", -- 5889 - 0x1701  :    7 - 0x7
    "00011111", -- 5890 - 0x1702  :   31 - 0x1f
    "00111111", -- 5891 - 0x1703  :   63 - 0x3f
    "01111111", -- 5892 - 0x1704  :  127 - 0x7f
    "11111111", -- 5893 - 0x1705  :  255 - 0xff
    "11111111", -- 5894 - 0x1706  :  255 - 0xff
    "11011101", -- 5895 - 0x1707  :  221 - 0xdd
    "00000000", -- 5896 - 0x1708  :    0 - 0x0
    "00000101", -- 5897 - 0x1709  :    5 - 0x5
    "00011001", -- 5898 - 0x170a  :   25 - 0x19
    "00110011", -- 5899 - 0x170b  :   51 - 0x33
    "01100011", -- 5900 - 0x170c  :   99 - 0x63
    "11000111", -- 5901 - 0x170d  :  199 - 0xc7
    "11000111", -- 5902 - 0x170e  :  199 - 0xc7
    "11000100", -- 5903 - 0x170f  :  196 - 0xc4
    "10001001", -- 5904 - 0x1710  :  137 - 0x89 -- Background 0x71
    "00000001", -- 5905 - 0x1711  :    1 - 0x1
    "00000001", -- 5906 - 0x1712  :    1 - 0x1
    "00000001", -- 5907 - 0x1713  :    1 - 0x1
    "00000001", -- 5908 - 0x1714  :    1 - 0x1
    "00000001", -- 5909 - 0x1715  :    1 - 0x1
    "00000000", -- 5910 - 0x1716  :    0 - 0x0
    "00000000", -- 5911 - 0x1717  :    0 - 0x0
    "10000000", -- 5912 - 0x1718  :  128 - 0x80
    "00000000", -- 5913 - 0x1719  :    0 - 0x0
    "00000000", -- 5914 - 0x171a  :    0 - 0x0
    "00000001", -- 5915 - 0x171b  :    1 - 0x1
    "00000001", -- 5916 - 0x171c  :    1 - 0x1
    "00000001", -- 5917 - 0x171d  :    1 - 0x1
    "00000000", -- 5918 - 0x171e  :    0 - 0x0
    "00000000", -- 5919 - 0x171f  :    0 - 0x0
    "10000000", -- 5920 - 0x1720  :  128 - 0x80 -- Background 0x72
    "11100000", -- 5921 - 0x1721  :  224 - 0xe0
    "11111000", -- 5922 - 0x1722  :  248 - 0xf8
    "11111100", -- 5923 - 0x1723  :  252 - 0xfc
    "11111110", -- 5924 - 0x1724  :  254 - 0xfe
    "11111111", -- 5925 - 0x1725  :  255 - 0xff
    "11111111", -- 5926 - 0x1726  :  255 - 0xff
    "00111011", -- 5927 - 0x1727  :   59 - 0x3b
    "00000000", -- 5928 - 0x1728  :    0 - 0x0
    "10100000", -- 5929 - 0x1729  :  160 - 0xa0
    "10011000", -- 5930 - 0x172a  :  152 - 0x98
    "11001100", -- 5931 - 0x172b  :  204 - 0xcc
    "11000110", -- 5932 - 0x172c  :  198 - 0xc6
    "11100011", -- 5933 - 0x172d  :  227 - 0xe3
    "11100011", -- 5934 - 0x172e  :  227 - 0xe3
    "00100011", -- 5935 - 0x172f  :   35 - 0x23
    "00010001", -- 5936 - 0x1730  :   17 - 0x11 -- Background 0x73
    "00000000", -- 5937 - 0x1731  :    0 - 0x0
    "00000000", -- 5938 - 0x1732  :    0 - 0x0
    "00000000", -- 5939 - 0x1733  :    0 - 0x0
    "00000000", -- 5940 - 0x1734  :    0 - 0x0
    "01000000", -- 5941 - 0x1735  :   64 - 0x40
    "10000000", -- 5942 - 0x1736  :  128 - 0x80
    "00000000", -- 5943 - 0x1737  :    0 - 0x0
    "00000001", -- 5944 - 0x1738  :    1 - 0x1
    "00000000", -- 5945 - 0x1739  :    0 - 0x0
    "00000000", -- 5946 - 0x173a  :    0 - 0x0
    "00000000", -- 5947 - 0x173b  :    0 - 0x0
    "00000000", -- 5948 - 0x173c  :    0 - 0x0
    "01000000", -- 5949 - 0x173d  :   64 - 0x40
    "10000000", -- 5950 - 0x173e  :  128 - 0x80
    "00000000", -- 5951 - 0x173f  :    0 - 0x0
    "00000001", -- 5952 - 0x1740  :    1 - 0x1 -- Background 0x74
    "00000001", -- 5953 - 0x1741  :    1 - 0x1
    "00000001", -- 5954 - 0x1742  :    1 - 0x1
    "00000001", -- 5955 - 0x1743  :    1 - 0x1
    "00000001", -- 5956 - 0x1744  :    1 - 0x1
    "00000001", -- 5957 - 0x1745  :    1 - 0x1
    "00000001", -- 5958 - 0x1746  :    1 - 0x1
    "00000001", -- 5959 - 0x1747  :    1 - 0x1
    "00000001", -- 5960 - 0x1748  :    1 - 0x1
    "00000001", -- 5961 - 0x1749  :    1 - 0x1
    "00000001", -- 5962 - 0x174a  :    1 - 0x1
    "00000001", -- 5963 - 0x174b  :    1 - 0x1
    "00000001", -- 5964 - 0x174c  :    1 - 0x1
    "00000001", -- 5965 - 0x174d  :    1 - 0x1
    "00000001", -- 5966 - 0x174e  :    1 - 0x1
    "00000001", -- 5967 - 0x174f  :    1 - 0x1
    "10000000", -- 5968 - 0x1750  :  128 - 0x80 -- Background 0x75
    "10000000", -- 5969 - 0x1751  :  128 - 0x80
    "10000000", -- 5970 - 0x1752  :  128 - 0x80
    "10000000", -- 5971 - 0x1753  :  128 - 0x80
    "10000000", -- 5972 - 0x1754  :  128 - 0x80
    "10000000", -- 5973 - 0x1755  :  128 - 0x80
    "10000000", -- 5974 - 0x1756  :  128 - 0x80
    "10000000", -- 5975 - 0x1757  :  128 - 0x80
    "10000000", -- 5976 - 0x1758  :  128 - 0x80
    "10000000", -- 5977 - 0x1759  :  128 - 0x80
    "10000000", -- 5978 - 0x175a  :  128 - 0x80
    "10000000", -- 5979 - 0x175b  :  128 - 0x80
    "10000000", -- 5980 - 0x175c  :  128 - 0x80
    "10000000", -- 5981 - 0x175d  :  128 - 0x80
    "10000000", -- 5982 - 0x175e  :  128 - 0x80
    "10000000", -- 5983 - 0x175f  :  128 - 0x80
    "00000001", -- 5984 - 0x1760  :    1 - 0x1 -- Background 0x76
    "00000011", -- 5985 - 0x1761  :    3 - 0x3
    "00000000", -- 5986 - 0x1762  :    0 - 0x0
    "00000000", -- 5987 - 0x1763  :    0 - 0x0
    "00000011", -- 5988 - 0x1764  :    3 - 0x3
    "00011001", -- 5989 - 0x1765  :   25 - 0x19
    "00000000", -- 5990 - 0x1766  :    0 - 0x0
    "00000000", -- 5991 - 0x1767  :    0 - 0x0
    "00000001", -- 5992 - 0x1768  :    1 - 0x1
    "00000011", -- 5993 - 0x1769  :    3 - 0x3
    "00000011", -- 5994 - 0x176a  :    3 - 0x3
    "00000111", -- 5995 - 0x176b  :    7 - 0x7
    "00000100", -- 5996 - 0x176c  :    4 - 0x4
    "00011100", -- 5997 - 0x176d  :   28 - 0x1c
    "00111111", -- 5998 - 0x176e  :   63 - 0x3f
    "01111111", -- 5999 - 0x176f  :  127 - 0x7f
    "00000000", -- 6000 - 0x1770  :    0 - 0x0 -- Background 0x77
    "00000000", -- 6001 - 0x1771  :    0 - 0x0
    "01111100", -- 6002 - 0x1772  :  124 - 0x7c
    "00000010", -- 6003 - 0x1773  :    2 - 0x2
    "00000001", -- 6004 - 0x1774  :    1 - 0x1
    "00000000", -- 6005 - 0x1775  :    0 - 0x0
    "00000000", -- 6006 - 0x1776  :    0 - 0x0
    "00000000", -- 6007 - 0x1777  :    0 - 0x0
    "01111111", -- 6008 - 0x1778  :  127 - 0x7f
    "11111111", -- 6009 - 0x1779  :  255 - 0xff
    "11111111", -- 6010 - 0x177a  :  255 - 0xff
    "01111111", -- 6011 - 0x177b  :  127 - 0x7f
    "01111111", -- 6012 - 0x177c  :  127 - 0x7f
    "00011111", -- 6013 - 0x177d  :   31 - 0x1f
    "00000011", -- 6014 - 0x177e  :    3 - 0x3
    "00000000", -- 6015 - 0x177f  :    0 - 0x0
    "00000000", -- 6016 - 0x1780  :    0 - 0x0 -- Background 0x78
    "00000000", -- 6017 - 0x1781  :    0 - 0x0
    "00000001", -- 6018 - 0x1782  :    1 - 0x1
    "00000001", -- 6019 - 0x1783  :    1 - 0x1
    "00000011", -- 6020 - 0x1784  :    3 - 0x3
    "00000111", -- 6021 - 0x1785  :    7 - 0x7
    "00000111", -- 6022 - 0x1786  :    7 - 0x7
    "00001111", -- 6023 - 0x1787  :   15 - 0xf
    "00000000", -- 6024 - 0x1788  :    0 - 0x0
    "00000000", -- 6025 - 0x1789  :    0 - 0x0
    "00000001", -- 6026 - 0x178a  :    1 - 0x1
    "00000001", -- 6027 - 0x178b  :    1 - 0x1
    "00000011", -- 6028 - 0x178c  :    3 - 0x3
    "00000111", -- 6029 - 0x178d  :    7 - 0x7
    "00000111", -- 6030 - 0x178e  :    7 - 0x7
    "00001111", -- 6031 - 0x178f  :   15 - 0xf
    "00001111", -- 6032 - 0x1790  :   15 - 0xf -- Background 0x79
    "00000111", -- 6033 - 0x1791  :    7 - 0x7
    "00001111", -- 6034 - 0x1792  :   15 - 0xf
    "00000111", -- 6035 - 0x1793  :    7 - 0x7
    "00000001", -- 6036 - 0x1794  :    1 - 0x1
    "00010000", -- 6037 - 0x1795  :   16 - 0x10
    "00100000", -- 6038 - 0x1796  :   32 - 0x20
    "00000000", -- 6039 - 0x1797  :    0 - 0x0
    "11111111", -- 6040 - 0x1798  :  255 - 0xff
    "11111111", -- 6041 - 0x1799  :  255 - 0xff
    "00111111", -- 6042 - 0x179a  :   63 - 0x3f
    "00111111", -- 6043 - 0x179b  :   63 - 0x3f
    "01111111", -- 6044 - 0x179c  :  127 - 0x7f
    "11111110", -- 6045 - 0x179d  :  254 - 0xfe
    "11111100", -- 6046 - 0x179e  :  252 - 0xfc
    "00110000", -- 6047 - 0x179f  :   48 - 0x30
    "11111000", -- 6048 - 0x17a0  :  248 - 0xf8 -- Background 0x7a
    "11111110", -- 6049 - 0x17a1  :  254 - 0xfe
    "01111111", -- 6050 - 0x17a2  :  127 - 0x7f
    "00011111", -- 6051 - 0x17a3  :   31 - 0x1f
    "00001111", -- 6052 - 0x17a4  :   15 - 0xf
    "00011001", -- 6053 - 0x17a5  :   25 - 0x19
    "00110000", -- 6054 - 0x17a6  :   48 - 0x30
    "01110000", -- 6055 - 0x17a7  :  112 - 0x70
    "11111000", -- 6056 - 0x17a8  :  248 - 0xf8
    "11111110", -- 6057 - 0x17a9  :  254 - 0xfe
    "11111111", -- 6058 - 0x17aa  :  255 - 0xff
    "11111111", -- 6059 - 0x17ab  :  255 - 0xff
    "11111111", -- 6060 - 0x17ac  :  255 - 0xff
    "11111111", -- 6061 - 0x17ad  :  255 - 0xff
    "11111111", -- 6062 - 0x17ae  :  255 - 0xff
    "11111111", -- 6063 - 0x17af  :  255 - 0xff
    "11111011", -- 6064 - 0x17b0  :  251 - 0xfb -- Background 0x7b
    "01110011", -- 6065 - 0x17b1  :  115 - 0x73
    "00100111", -- 6066 - 0x17b2  :   39 - 0x27
    "00001111", -- 6067 - 0x17b3  :   15 - 0xf
    "00011111", -- 6068 - 0x17b4  :   31 - 0x1f
    "00011111", -- 6069 - 0x17b5  :   31 - 0x1f
    "00111111", -- 6070 - 0x17b6  :   63 - 0x3f
    "01111111", -- 6071 - 0x17b7  :  127 - 0x7f
    "11111111", -- 6072 - 0x17b8  :  255 - 0xff
    "11111111", -- 6073 - 0x17b9  :  255 - 0xff
    "11111111", -- 6074 - 0x17ba  :  255 - 0xff
    "11111111", -- 6075 - 0x17bb  :  255 - 0xff
    "11111111", -- 6076 - 0x17bc  :  255 - 0xff
    "11111111", -- 6077 - 0x17bd  :  255 - 0xff
    "11111111", -- 6078 - 0x17be  :  255 - 0xff
    "01111111", -- 6079 - 0x17bf  :  127 - 0x7f
    "11111111", -- 6080 - 0x17c0  :  255 - 0xff -- Background 0x7c
    "11111111", -- 6081 - 0x17c1  :  255 - 0xff
    "11111111", -- 6082 - 0x17c2  :  255 - 0xff
    "11111111", -- 6083 - 0x17c3  :  255 - 0xff
    "11111110", -- 6084 - 0x17c4  :  254 - 0xfe
    "11111101", -- 6085 - 0x17c5  :  253 - 0xfd
    "11111000", -- 6086 - 0x17c6  :  248 - 0xf8
    "11110110", -- 6087 - 0x17c7  :  246 - 0xf6
    "11111111", -- 6088 - 0x17c8  :  255 - 0xff
    "11111111", -- 6089 - 0x17c9  :  255 - 0xff
    "11111111", -- 6090 - 0x17ca  :  255 - 0xff
    "11111111", -- 6091 - 0x17cb  :  255 - 0xff
    "11111111", -- 6092 - 0x17cc  :  255 - 0xff
    "11111111", -- 6093 - 0x17cd  :  255 - 0xff
    "11111111", -- 6094 - 0x17ce  :  255 - 0xff
    "11111111", -- 6095 - 0x17cf  :  255 - 0xff
    "11101111", -- 6096 - 0x17d0  :  239 - 0xef -- Background 0x7d
    "11001111", -- 6097 - 0x17d1  :  207 - 0xcf
    "10011111", -- 6098 - 0x17d2  :  159 - 0x9f
    "00011111", -- 6099 - 0x17d3  :   31 - 0x1f
    "00001111", -- 6100 - 0x17d4  :   15 - 0xf
    "00101101", -- 6101 - 0x17d5  :   45 - 0x2d
    "01010000", -- 6102 - 0x17d6  :   80 - 0x50
    "01000000", -- 6103 - 0x17d7  :   64 - 0x40
    "11101111", -- 6104 - 0x17d8  :  239 - 0xef
    "11001111", -- 6105 - 0x17d9  :  207 - 0xcf
    "10011111", -- 6106 - 0x17da  :  159 - 0x9f
    "00011111", -- 6107 - 0x17db  :   31 - 0x1f
    "00001111", -- 6108 - 0x17dc  :   15 - 0xf
    "01111111", -- 6109 - 0x17dd  :  127 - 0x7f
    "11111111", -- 6110 - 0x17de  :  255 - 0xff
    "11111111", -- 6111 - 0x17df  :  255 - 0xff
    "00000000", -- 6112 - 0x17e0  :    0 - 0x0 -- Background 0x7e
    "00000000", -- 6113 - 0x17e1  :    0 - 0x0
    "00000000", -- 6114 - 0x17e2  :    0 - 0x0
    "00000000", -- 6115 - 0x17e3  :    0 - 0x0
    "11100000", -- 6116 - 0x17e4  :  224 - 0xe0
    "11111110", -- 6117 - 0x17e5  :  254 - 0xfe
    "11111111", -- 6118 - 0x17e6  :  255 - 0xff
    "11110011", -- 6119 - 0x17e7  :  243 - 0xf3
    "00000000", -- 6120 - 0x17e8  :    0 - 0x0
    "00000000", -- 6121 - 0x17e9  :    0 - 0x0
    "00000000", -- 6122 - 0x17ea  :    0 - 0x0
    "11110000", -- 6123 - 0x17eb  :  240 - 0xf0
    "11111110", -- 6124 - 0x17ec  :  254 - 0xfe
    "11111111", -- 6125 - 0x17ed  :  255 - 0xff
    "11111111", -- 6126 - 0x17ee  :  255 - 0xff
    "11111111", -- 6127 - 0x17ef  :  255 - 0xff
    "11111011", -- 6128 - 0x17f0  :  251 - 0xfb -- Background 0x7f
    "11111011", -- 6129 - 0x17f1  :  251 - 0xfb
    "11111011", -- 6130 - 0x17f2  :  251 - 0xfb
    "11111011", -- 6131 - 0x17f3  :  251 - 0xfb
    "11111011", -- 6132 - 0x17f4  :  251 - 0xfb
    "11110011", -- 6133 - 0x17f5  :  243 - 0xf3
    "11110111", -- 6134 - 0x17f6  :  247 - 0xf7
    "11100111", -- 6135 - 0x17f7  :  231 - 0xe7
    "11111111", -- 6136 - 0x17f8  :  255 - 0xff
    "11111111", -- 6137 - 0x17f9  :  255 - 0xff
    "11111111", -- 6138 - 0x17fa  :  255 - 0xff
    "11111111", -- 6139 - 0x17fb  :  255 - 0xff
    "11111111", -- 6140 - 0x17fc  :  255 - 0xff
    "11111111", -- 6141 - 0x17fd  :  255 - 0xff
    "11111111", -- 6142 - 0x17fe  :  255 - 0xff
    "11111111", -- 6143 - 0x17ff  :  255 - 0xff
    "11001111", -- 6144 - 0x1800  :  207 - 0xcf -- Background 0x80
    "10011111", -- 6145 - 0x1801  :  159 - 0x9f
    "00111111", -- 6146 - 0x1802  :   63 - 0x3f
    "00111111", -- 6147 - 0x1803  :   63 - 0x3f
    "00111111", -- 6148 - 0x1804  :   63 - 0x3f
    "00001111", -- 6149 - 0x1805  :   15 - 0xf
    "00000011", -- 6150 - 0x1806  :    3 - 0x3
    "00000000", -- 6151 - 0x1807  :    0 - 0x0
    "11111111", -- 6152 - 0x1808  :  255 - 0xff
    "11111111", -- 6153 - 0x1809  :  255 - 0xff
    "11111111", -- 6154 - 0x180a  :  255 - 0xff
    "11111111", -- 6155 - 0x180b  :  255 - 0xff
    "11111111", -- 6156 - 0x180c  :  255 - 0xff
    "11111111", -- 6157 - 0x180d  :  255 - 0xff
    "11111111", -- 6158 - 0x180e  :  255 - 0xff
    "11111111", -- 6159 - 0x180f  :  255 - 0xff
    "11000000", -- 6160 - 0x1810  :  192 - 0xc0 -- Background 0x81
    "11110000", -- 6161 - 0x1811  :  240 - 0xf0
    "11111100", -- 6162 - 0x1812  :  252 - 0xfc
    "11110000", -- 6163 - 0x1813  :  240 - 0xf0
    "11110000", -- 6164 - 0x1814  :  240 - 0xf0
    "10011000", -- 6165 - 0x1815  :  152 - 0x98
    "00001000", -- 6166 - 0x1816  :    8 - 0x8
    "00000000", -- 6167 - 0x1817  :    0 - 0x0
    "11111111", -- 6168 - 0x1818  :  255 - 0xff
    "11111111", -- 6169 - 0x1819  :  255 - 0xff
    "11111111", -- 6170 - 0x181a  :  255 - 0xff
    "11110000", -- 6171 - 0x181b  :  240 - 0xf0
    "11110000", -- 6172 - 0x181c  :  240 - 0xf0
    "11111000", -- 6173 - 0x181d  :  248 - 0xf8
    "11111000", -- 6174 - 0x181e  :  248 - 0xf8
    "11111000", -- 6175 - 0x181f  :  248 - 0xf8
    "00000000", -- 6176 - 0x1820  :    0 - 0x0 -- Background 0x82
    "00000000", -- 6177 - 0x1821  :    0 - 0x0
    "00000000", -- 6178 - 0x1822  :    0 - 0x0
    "00000000", -- 6179 - 0x1823  :    0 - 0x0
    "00000000", -- 6180 - 0x1824  :    0 - 0x0
    "00000000", -- 6181 - 0x1825  :    0 - 0x0
    "10000000", -- 6182 - 0x1826  :  128 - 0x80
    "11000000", -- 6183 - 0x1827  :  192 - 0xc0
    "00000000", -- 6184 - 0x1828  :    0 - 0x0
    "00000000", -- 6185 - 0x1829  :    0 - 0x0
    "00000000", -- 6186 - 0x182a  :    0 - 0x0
    "00000000", -- 6187 - 0x182b  :    0 - 0x0
    "00000000", -- 6188 - 0x182c  :    0 - 0x0
    "10000000", -- 6189 - 0x182d  :  128 - 0x80
    "11000000", -- 6190 - 0x182e  :  192 - 0xc0
    "11100000", -- 6191 - 0x182f  :  224 - 0xe0
    "11100000", -- 6192 - 0x1830  :  224 - 0xe0 -- Background 0x83
    "11100000", -- 6193 - 0x1831  :  224 - 0xe0
    "11110000", -- 6194 - 0x1832  :  240 - 0xf0
    "11110000", -- 6195 - 0x1833  :  240 - 0xf0
    "11110000", -- 6196 - 0x1834  :  240 - 0xf0
    "11110000", -- 6197 - 0x1835  :  240 - 0xf0
    "11111000", -- 6198 - 0x1836  :  248 - 0xf8
    "11111000", -- 6199 - 0x1837  :  248 - 0xf8
    "11110000", -- 6200 - 0x1838  :  240 - 0xf0
    "11110000", -- 6201 - 0x1839  :  240 - 0xf0
    "11111000", -- 6202 - 0x183a  :  248 - 0xf8
    "11111000", -- 6203 - 0x183b  :  248 - 0xf8
    "11111000", -- 6204 - 0x183c  :  248 - 0xf8
    "11111100", -- 6205 - 0x183d  :  252 - 0xfc
    "11111100", -- 6206 - 0x183e  :  252 - 0xfc
    "11111110", -- 6207 - 0x183f  :  254 - 0xfe
    "11111110", -- 6208 - 0x1840  :  254 - 0xfe -- Background 0x84
    "11111111", -- 6209 - 0x1841  :  255 - 0xff
    "11111111", -- 6210 - 0x1842  :  255 - 0xff
    "11111111", -- 6211 - 0x1843  :  255 - 0xff
    "11111111", -- 6212 - 0x1844  :  255 - 0xff
    "11111111", -- 6213 - 0x1845  :  255 - 0xff
    "11111111", -- 6214 - 0x1846  :  255 - 0xff
    "11111111", -- 6215 - 0x1847  :  255 - 0xff
    "11111111", -- 6216 - 0x1848  :  255 - 0xff
    "11111111", -- 6217 - 0x1849  :  255 - 0xff
    "11111111", -- 6218 - 0x184a  :  255 - 0xff
    "11111111", -- 6219 - 0x184b  :  255 - 0xff
    "11111111", -- 6220 - 0x184c  :  255 - 0xff
    "11111111", -- 6221 - 0x184d  :  255 - 0xff
    "11111111", -- 6222 - 0x184e  :  255 - 0xff
    "11111111", -- 6223 - 0x184f  :  255 - 0xff
    "00111111", -- 6224 - 0x1850  :   63 - 0x3f -- Background 0x85
    "00011111", -- 6225 - 0x1851  :   31 - 0x1f
    "00011111", -- 6226 - 0x1852  :   31 - 0x1f
    "00001111", -- 6227 - 0x1853  :   15 - 0xf
    "00000111", -- 6228 - 0x1854  :    7 - 0x7
    "00000000", -- 6229 - 0x1855  :    0 - 0x0
    "00000000", -- 6230 - 0x1856  :    0 - 0x0
    "00000000", -- 6231 - 0x1857  :    0 - 0x0
    "11111111", -- 6232 - 0x1858  :  255 - 0xff
    "11111111", -- 6233 - 0x1859  :  255 - 0xff
    "11111111", -- 6234 - 0x185a  :  255 - 0xff
    "00001111", -- 6235 - 0x185b  :   15 - 0xf
    "00000111", -- 6236 - 0x185c  :    7 - 0x7
    "00000000", -- 6237 - 0x185d  :    0 - 0x0
    "00000000", -- 6238 - 0x185e  :    0 - 0x0
    "00000000", -- 6239 - 0x185f  :    0 - 0x0
    "00000000", -- 6240 - 0x1860  :    0 - 0x0 -- Background 0x86
    "00000000", -- 6241 - 0x1861  :    0 - 0x0
    "11000000", -- 6242 - 0x1862  :  192 - 0xc0
    "11100000", -- 6243 - 0x1863  :  224 - 0xe0
    "11110000", -- 6244 - 0x1864  :  240 - 0xf0
    "11110000", -- 6245 - 0x1865  :  240 - 0xf0
    "11110000", -- 6246 - 0x1866  :  240 - 0xf0
    "11111000", -- 6247 - 0x1867  :  248 - 0xf8
    "00000000", -- 6248 - 0x1868  :    0 - 0x0
    "10000000", -- 6249 - 0x1869  :  128 - 0x80
    "11000000", -- 6250 - 0x186a  :  192 - 0xc0
    "11100000", -- 6251 - 0x186b  :  224 - 0xe0
    "11110000", -- 6252 - 0x186c  :  240 - 0xf0
    "11110000", -- 6253 - 0x186d  :  240 - 0xf0
    "11110000", -- 6254 - 0x186e  :  240 - 0xf0
    "11111100", -- 6255 - 0x186f  :  252 - 0xfc
    "11111001", -- 6256 - 0x1870  :  249 - 0xf9 -- Background 0x87
    "11111111", -- 6257 - 0x1871  :  255 - 0xff
    "11111111", -- 6258 - 0x1872  :  255 - 0xff
    "11111111", -- 6259 - 0x1873  :  255 - 0xff
    "11111111", -- 6260 - 0x1874  :  255 - 0xff
    "00001110", -- 6261 - 0x1875  :   14 - 0xe
    "00000010", -- 6262 - 0x1876  :    2 - 0x2
    "00010100", -- 6263 - 0x1877  :   20 - 0x14
    "11111111", -- 6264 - 0x1878  :  255 - 0xff
    "11111111", -- 6265 - 0x1879  :  255 - 0xff
    "11111111", -- 6266 - 0x187a  :  255 - 0xff
    "11111111", -- 6267 - 0x187b  :  255 - 0xff
    "11111111", -- 6268 - 0x187c  :  255 - 0xff
    "00001111", -- 6269 - 0x187d  :   15 - 0xf
    "00011111", -- 6270 - 0x187e  :   31 - 0x1f
    "00111111", -- 6271 - 0x187f  :   63 - 0x3f
    "10000000", -- 6272 - 0x1880  :  128 - 0x80 -- Background 0x88
    "10100000", -- 6273 - 0x1881  :  160 - 0xa0
    "00100000", -- 6274 - 0x1882  :   32 - 0x20
    "00100000", -- 6275 - 0x1883  :   32 - 0x20
    "10100000", -- 6276 - 0x1884  :  160 - 0xa0
    "10000000", -- 6277 - 0x1885  :  128 - 0x80
    "00000000", -- 6278 - 0x1886  :    0 - 0x0
    "00000000", -- 6279 - 0x1887  :    0 - 0x0
    "11000000", -- 6280 - 0x1888  :  192 - 0xc0
    "11100000", -- 6281 - 0x1889  :  224 - 0xe0
    "11100000", -- 6282 - 0x188a  :  224 - 0xe0
    "11100000", -- 6283 - 0x188b  :  224 - 0xe0
    "11100000", -- 6284 - 0x188c  :  224 - 0xe0
    "11000000", -- 6285 - 0x188d  :  192 - 0xc0
    "11000000", -- 6286 - 0x188e  :  192 - 0xc0
    "10000000", -- 6287 - 0x188f  :  128 - 0x80
    "00000001", -- 6288 - 0x1890  :    1 - 0x1 -- Background 0x89
    "00000101", -- 6289 - 0x1891  :    5 - 0x5
    "00000100", -- 6290 - 0x1892  :    4 - 0x4
    "00000100", -- 6291 - 0x1893  :    4 - 0x4
    "00000101", -- 6292 - 0x1894  :    5 - 0x5
    "00000001", -- 6293 - 0x1895  :    1 - 0x1
    "00000000", -- 6294 - 0x1896  :    0 - 0x0
    "00000000", -- 6295 - 0x1897  :    0 - 0x0
    "00000011", -- 6296 - 0x1898  :    3 - 0x3
    "00000111", -- 6297 - 0x1899  :    7 - 0x7
    "00000111", -- 6298 - 0x189a  :    7 - 0x7
    "00000111", -- 6299 - 0x189b  :    7 - 0x7
    "00000111", -- 6300 - 0x189c  :    7 - 0x7
    "00000011", -- 6301 - 0x189d  :    3 - 0x3
    "00000011", -- 6302 - 0x189e  :    3 - 0x3
    "00000001", -- 6303 - 0x189f  :    1 - 0x1
    "00000000", -- 6304 - 0x18a0  :    0 - 0x0 -- Background 0x8a
    "00000000", -- 6305 - 0x18a1  :    0 - 0x0
    "00000011", -- 6306 - 0x18a2  :    3 - 0x3
    "00000111", -- 6307 - 0x18a3  :    7 - 0x7
    "00001111", -- 6308 - 0x18a4  :   15 - 0xf
    "00001111", -- 6309 - 0x18a5  :   15 - 0xf
    "00001111", -- 6310 - 0x18a6  :   15 - 0xf
    "00001111", -- 6311 - 0x18a7  :   15 - 0xf
    "00000000", -- 6312 - 0x18a8  :    0 - 0x0
    "00000001", -- 6313 - 0x18a9  :    1 - 0x1
    "00000011", -- 6314 - 0x18aa  :    3 - 0x3
    "00000111", -- 6315 - 0x18ab  :    7 - 0x7
    "00001111", -- 6316 - 0x18ac  :   15 - 0xf
    "00001111", -- 6317 - 0x18ad  :   15 - 0xf
    "00001111", -- 6318 - 0x18ae  :   15 - 0xf
    "00111111", -- 6319 - 0x18af  :   63 - 0x3f
    "10011111", -- 6320 - 0x18b0  :  159 - 0x9f -- Background 0x8b
    "11111111", -- 6321 - 0x18b1  :  255 - 0xff
    "11111111", -- 6322 - 0x18b2  :  255 - 0xff
    "11111111", -- 6323 - 0x18b3  :  255 - 0xff
    "11111111", -- 6324 - 0x18b4  :  255 - 0xff
    "01110000", -- 6325 - 0x18b5  :  112 - 0x70
    "01000000", -- 6326 - 0x18b6  :   64 - 0x40
    "00101000", -- 6327 - 0x18b7  :   40 - 0x28
    "11111111", -- 6328 - 0x18b8  :  255 - 0xff
    "11111111", -- 6329 - 0x18b9  :  255 - 0xff
    "11111111", -- 6330 - 0x18ba  :  255 - 0xff
    "11111111", -- 6331 - 0x18bb  :  255 - 0xff
    "11111111", -- 6332 - 0x18bc  :  255 - 0xff
    "11110000", -- 6333 - 0x18bd  :  240 - 0xf0
    "11111000", -- 6334 - 0x18be  :  248 - 0xf8
    "11111100", -- 6335 - 0x18bf  :  252 - 0xfc
    "00000000", -- 6336 - 0x18c0  :    0 - 0x0 -- Background 0x8c
    "00000000", -- 6337 - 0x18c1  :    0 - 0x0
    "00000000", -- 6338 - 0x18c2  :    0 - 0x0
    "00000000", -- 6339 - 0x18c3  :    0 - 0x0
    "00000000", -- 6340 - 0x18c4  :    0 - 0x0
    "00000000", -- 6341 - 0x18c5  :    0 - 0x0
    "00000001", -- 6342 - 0x18c6  :    1 - 0x1
    "00000011", -- 6343 - 0x18c7  :    3 - 0x3
    "00000000", -- 6344 - 0x18c8  :    0 - 0x0
    "00000000", -- 6345 - 0x18c9  :    0 - 0x0
    "00000000", -- 6346 - 0x18ca  :    0 - 0x0
    "00000000", -- 6347 - 0x18cb  :    0 - 0x0
    "00000000", -- 6348 - 0x18cc  :    0 - 0x0
    "00000001", -- 6349 - 0x18cd  :    1 - 0x1
    "00000011", -- 6350 - 0x18ce  :    3 - 0x3
    "00000111", -- 6351 - 0x18cf  :    7 - 0x7
    "00000111", -- 6352 - 0x18d0  :    7 - 0x7 -- Background 0x8d
    "00000111", -- 6353 - 0x18d1  :    7 - 0x7
    "00001111", -- 6354 - 0x18d2  :   15 - 0xf
    "00001111", -- 6355 - 0x18d3  :   15 - 0xf
    "00001111", -- 6356 - 0x18d4  :   15 - 0xf
    "00001111", -- 6357 - 0x18d5  :   15 - 0xf
    "00011111", -- 6358 - 0x18d6  :   31 - 0x1f
    "00011111", -- 6359 - 0x18d7  :   31 - 0x1f
    "00001111", -- 6360 - 0x18d8  :   15 - 0xf
    "00001111", -- 6361 - 0x18d9  :   15 - 0xf
    "00011111", -- 6362 - 0x18da  :   31 - 0x1f
    "00011111", -- 6363 - 0x18db  :   31 - 0x1f
    "00011111", -- 6364 - 0x18dc  :   31 - 0x1f
    "00111111", -- 6365 - 0x18dd  :   63 - 0x3f
    "00111111", -- 6366 - 0x18de  :   63 - 0x3f
    "01111111", -- 6367 - 0x18df  :  127 - 0x7f
    "01111111", -- 6368 - 0x18e0  :  127 - 0x7f -- Background 0x8e
    "11111111", -- 6369 - 0x18e1  :  255 - 0xff
    "11111111", -- 6370 - 0x18e2  :  255 - 0xff
    "11111111", -- 6371 - 0x18e3  :  255 - 0xff
    "11111111", -- 6372 - 0x18e4  :  255 - 0xff
    "11111111", -- 6373 - 0x18e5  :  255 - 0xff
    "11111111", -- 6374 - 0x18e6  :  255 - 0xff
    "11111111", -- 6375 - 0x18e7  :  255 - 0xff
    "11111111", -- 6376 - 0x18e8  :  255 - 0xff
    "11111111", -- 6377 - 0x18e9  :  255 - 0xff
    "11111111", -- 6378 - 0x18ea  :  255 - 0xff
    "11111111", -- 6379 - 0x18eb  :  255 - 0xff
    "11111111", -- 6380 - 0x18ec  :  255 - 0xff
    "11111111", -- 6381 - 0x18ed  :  255 - 0xff
    "11111111", -- 6382 - 0x18ee  :  255 - 0xff
    "11111111", -- 6383 - 0x18ef  :  255 - 0xff
    "11111100", -- 6384 - 0x18f0  :  252 - 0xfc -- Background 0x8f
    "11111000", -- 6385 - 0x18f1  :  248 - 0xf8
    "11111000", -- 6386 - 0x18f2  :  248 - 0xf8
    "11110000", -- 6387 - 0x18f3  :  240 - 0xf0
    "11100000", -- 6388 - 0x18f4  :  224 - 0xe0
    "00000000", -- 6389 - 0x18f5  :    0 - 0x0
    "00000000", -- 6390 - 0x18f6  :    0 - 0x0
    "00000000", -- 6391 - 0x18f7  :    0 - 0x0
    "11111111", -- 6392 - 0x18f8  :  255 - 0xff
    "11111111", -- 6393 - 0x18f9  :  255 - 0xff
    "11111111", -- 6394 - 0x18fa  :  255 - 0xff
    "11110000", -- 6395 - 0x18fb  :  240 - 0xf0
    "11100000", -- 6396 - 0x18fc  :  224 - 0xe0
    "00000000", -- 6397 - 0x18fd  :    0 - 0x0
    "00000000", -- 6398 - 0x18fe  :    0 - 0x0
    "00000000", -- 6399 - 0x18ff  :    0 - 0x0
    "00000000", -- 6400 - 0x1900  :    0 - 0x0 -- Background 0x90
    "00000000", -- 6401 - 0x1901  :    0 - 0x0
    "00000000", -- 6402 - 0x1902  :    0 - 0x0
    "00000000", -- 6403 - 0x1903  :    0 - 0x0
    "00000111", -- 6404 - 0x1904  :    7 - 0x7
    "01111111", -- 6405 - 0x1905  :  127 - 0x7f
    "11111111", -- 6406 - 0x1906  :  255 - 0xff
    "11001111", -- 6407 - 0x1907  :  207 - 0xcf
    "00000000", -- 6408 - 0x1908  :    0 - 0x0
    "00000000", -- 6409 - 0x1909  :    0 - 0x0
    "00000000", -- 6410 - 0x190a  :    0 - 0x0
    "00001111", -- 6411 - 0x190b  :   15 - 0xf
    "01111111", -- 6412 - 0x190c  :  127 - 0x7f
    "11111111", -- 6413 - 0x190d  :  255 - 0xff
    "11111111", -- 6414 - 0x190e  :  255 - 0xff
    "11111111", -- 6415 - 0x190f  :  255 - 0xff
    "11011111", -- 6416 - 0x1910  :  223 - 0xdf -- Background 0x91
    "11011111", -- 6417 - 0x1911  :  223 - 0xdf
    "11011111", -- 6418 - 0x1912  :  223 - 0xdf
    "11011111", -- 6419 - 0x1913  :  223 - 0xdf
    "11011111", -- 6420 - 0x1914  :  223 - 0xdf
    "11001111", -- 6421 - 0x1915  :  207 - 0xcf
    "11101111", -- 6422 - 0x1916  :  239 - 0xef
    "11100111", -- 6423 - 0x1917  :  231 - 0xe7
    "11111111", -- 6424 - 0x1918  :  255 - 0xff
    "11111111", -- 6425 - 0x1919  :  255 - 0xff
    "11111111", -- 6426 - 0x191a  :  255 - 0xff
    "11111111", -- 6427 - 0x191b  :  255 - 0xff
    "11111111", -- 6428 - 0x191c  :  255 - 0xff
    "11111111", -- 6429 - 0x191d  :  255 - 0xff
    "11111111", -- 6430 - 0x191e  :  255 - 0xff
    "11111111", -- 6431 - 0x191f  :  255 - 0xff
    "11110011", -- 6432 - 0x1920  :  243 - 0xf3 -- Background 0x92
    "11111001", -- 6433 - 0x1921  :  249 - 0xf9
    "11111100", -- 6434 - 0x1922  :  252 - 0xfc
    "11111100", -- 6435 - 0x1923  :  252 - 0xfc
    "11111100", -- 6436 - 0x1924  :  252 - 0xfc
    "11110000", -- 6437 - 0x1925  :  240 - 0xf0
    "11000000", -- 6438 - 0x1926  :  192 - 0xc0
    "00000000", -- 6439 - 0x1927  :    0 - 0x0
    "11111111", -- 6440 - 0x1928  :  255 - 0xff
    "11111111", -- 6441 - 0x1929  :  255 - 0xff
    "11111111", -- 6442 - 0x192a  :  255 - 0xff
    "11111111", -- 6443 - 0x192b  :  255 - 0xff
    "11111111", -- 6444 - 0x192c  :  255 - 0xff
    "11111111", -- 6445 - 0x192d  :  255 - 0xff
    "11111111", -- 6446 - 0x192e  :  255 - 0xff
    "11111111", -- 6447 - 0x192f  :  255 - 0xff
    "00000011", -- 6448 - 0x1930  :    3 - 0x3 -- Background 0x93
    "00001111", -- 6449 - 0x1931  :   15 - 0xf
    "00111111", -- 6450 - 0x1932  :   63 - 0x3f
    "00001111", -- 6451 - 0x1933  :   15 - 0xf
    "00001111", -- 6452 - 0x1934  :   15 - 0xf
    "00011001", -- 6453 - 0x1935  :   25 - 0x19
    "00010000", -- 6454 - 0x1936  :   16 - 0x10
    "00000000", -- 6455 - 0x1937  :    0 - 0x0
    "11111111", -- 6456 - 0x1938  :  255 - 0xff
    "11111111", -- 6457 - 0x1939  :  255 - 0xff
    "11111111", -- 6458 - 0x193a  :  255 - 0xff
    "00001111", -- 6459 - 0x193b  :   15 - 0xf
    "00001111", -- 6460 - 0x193c  :   15 - 0xf
    "00011111", -- 6461 - 0x193d  :   31 - 0x1f
    "00011111", -- 6462 - 0x193e  :   31 - 0x1f
    "00011111", -- 6463 - 0x193f  :   31 - 0x1f
    "00011111", -- 6464 - 0x1940  :   31 - 0x1f -- Background 0x94
    "01111111", -- 6465 - 0x1941  :  127 - 0x7f
    "11111110", -- 6466 - 0x1942  :  254 - 0xfe
    "11111000", -- 6467 - 0x1943  :  248 - 0xf8
    "11110000", -- 6468 - 0x1944  :  240 - 0xf0
    "10011000", -- 6469 - 0x1945  :  152 - 0x98
    "00001100", -- 6470 - 0x1946  :   12 - 0xc
    "00001110", -- 6471 - 0x1947  :   14 - 0xe
    "00011111", -- 6472 - 0x1948  :   31 - 0x1f
    "01111111", -- 6473 - 0x1949  :  127 - 0x7f
    "11111111", -- 6474 - 0x194a  :  255 - 0xff
    "11111111", -- 6475 - 0x194b  :  255 - 0xff
    "11111111", -- 6476 - 0x194c  :  255 - 0xff
    "11111111", -- 6477 - 0x194d  :  255 - 0xff
    "11111111", -- 6478 - 0x194e  :  255 - 0xff
    "11111111", -- 6479 - 0x194f  :  255 - 0xff
    "11011111", -- 6480 - 0x1950  :  223 - 0xdf -- Background 0x95
    "11001110", -- 6481 - 0x1951  :  206 - 0xce
    "11100100", -- 6482 - 0x1952  :  228 - 0xe4
    "11110000", -- 6483 - 0x1953  :  240 - 0xf0
    "11111000", -- 6484 - 0x1954  :  248 - 0xf8
    "11111000", -- 6485 - 0x1955  :  248 - 0xf8
    "11111100", -- 6486 - 0x1956  :  252 - 0xfc
    "11111110", -- 6487 - 0x1957  :  254 - 0xfe
    "11111111", -- 6488 - 0x1958  :  255 - 0xff
    "11111111", -- 6489 - 0x1959  :  255 - 0xff
    "11111111", -- 6490 - 0x195a  :  255 - 0xff
    "11111111", -- 6491 - 0x195b  :  255 - 0xff
    "11111111", -- 6492 - 0x195c  :  255 - 0xff
    "11111111", -- 6493 - 0x195d  :  255 - 0xff
    "11111111", -- 6494 - 0x195e  :  255 - 0xff
    "11111110", -- 6495 - 0x195f  :  254 - 0xfe
    "11111111", -- 6496 - 0x1960  :  255 - 0xff -- Background 0x96
    "11111111", -- 6497 - 0x1961  :  255 - 0xff
    "11111111", -- 6498 - 0x1962  :  255 - 0xff
    "11111111", -- 6499 - 0x1963  :  255 - 0xff
    "01111111", -- 6500 - 0x1964  :  127 - 0x7f
    "10111111", -- 6501 - 0x1965  :  191 - 0xbf
    "00011111", -- 6502 - 0x1966  :   31 - 0x1f
    "01101111", -- 6503 - 0x1967  :  111 - 0x6f
    "11111111", -- 6504 - 0x1968  :  255 - 0xff
    "11111111", -- 6505 - 0x1969  :  255 - 0xff
    "11111111", -- 6506 - 0x196a  :  255 - 0xff
    "11111111", -- 6507 - 0x196b  :  255 - 0xff
    "11111111", -- 6508 - 0x196c  :  255 - 0xff
    "11111111", -- 6509 - 0x196d  :  255 - 0xff
    "11111111", -- 6510 - 0x196e  :  255 - 0xff
    "11111111", -- 6511 - 0x196f  :  255 - 0xff
    "11110111", -- 6512 - 0x1970  :  247 - 0xf7 -- Background 0x97
    "11110011", -- 6513 - 0x1971  :  243 - 0xf3
    "11111001", -- 6514 - 0x1972  :  249 - 0xf9
    "11111000", -- 6515 - 0x1973  :  248 - 0xf8
    "11110000", -- 6516 - 0x1974  :  240 - 0xf0
    "10110100", -- 6517 - 0x1975  :  180 - 0xb4
    "00001010", -- 6518 - 0x1976  :   10 - 0xa
    "00000010", -- 6519 - 0x1977  :    2 - 0x2
    "11110111", -- 6520 - 0x1978  :  247 - 0xf7
    "11110011", -- 6521 - 0x1979  :  243 - 0xf3
    "11111001", -- 6522 - 0x197a  :  249 - 0xf9
    "11111000", -- 6523 - 0x197b  :  248 - 0xf8
    "11110000", -- 6524 - 0x197c  :  240 - 0xf0
    "11111110", -- 6525 - 0x197d  :  254 - 0xfe
    "11111111", -- 6526 - 0x197e  :  255 - 0xff
    "11111111", -- 6527 - 0x197f  :  255 - 0xff
    "10000000", -- 6528 - 0x1980  :  128 - 0x80 -- Background 0x98
    "11000000", -- 6529 - 0x1981  :  192 - 0xc0
    "00000000", -- 6530 - 0x1982  :    0 - 0x0
    "00000000", -- 6531 - 0x1983  :    0 - 0x0
    "11000000", -- 6532 - 0x1984  :  192 - 0xc0
    "10011000", -- 6533 - 0x1985  :  152 - 0x98
    "00000000", -- 6534 - 0x1986  :    0 - 0x0
    "00000000", -- 6535 - 0x1987  :    0 - 0x0
    "10000000", -- 6536 - 0x1988  :  128 - 0x80
    "11000000", -- 6537 - 0x1989  :  192 - 0xc0
    "11000000", -- 6538 - 0x198a  :  192 - 0xc0
    "11100000", -- 6539 - 0x198b  :  224 - 0xe0
    "00100000", -- 6540 - 0x198c  :   32 - 0x20
    "00111000", -- 6541 - 0x198d  :   56 - 0x38
    "11111100", -- 6542 - 0x198e  :  252 - 0xfc
    "11111110", -- 6543 - 0x198f  :  254 - 0xfe
    "00000000", -- 6544 - 0x1990  :    0 - 0x0 -- Background 0x99
    "00000000", -- 6545 - 0x1991  :    0 - 0x0
    "00111110", -- 6546 - 0x1992  :   62 - 0x3e
    "01000000", -- 6547 - 0x1993  :   64 - 0x40
    "10000000", -- 6548 - 0x1994  :  128 - 0x80
    "00000000", -- 6549 - 0x1995  :    0 - 0x0
    "00000000", -- 6550 - 0x1996  :    0 - 0x0
    "00000000", -- 6551 - 0x1997  :    0 - 0x0
    "11111110", -- 6552 - 0x1998  :  254 - 0xfe
    "11111111", -- 6553 - 0x1999  :  255 - 0xff
    "11111111", -- 6554 - 0x199a  :  255 - 0xff
    "11111110", -- 6555 - 0x199b  :  254 - 0xfe
    "11111100", -- 6556 - 0x199c  :  252 - 0xfc
    "11111000", -- 6557 - 0x199d  :  248 - 0xf8
    "11000000", -- 6558 - 0x199e  :  192 - 0xc0
    "00000000", -- 6559 - 0x199f  :    0 - 0x0
    "00000000", -- 6560 - 0x19a0  :    0 - 0x0 -- Background 0x9a
    "00000000", -- 6561 - 0x19a1  :    0 - 0x0
    "10000000", -- 6562 - 0x19a2  :  128 - 0x80
    "10000000", -- 6563 - 0x19a3  :  128 - 0x80
    "11000000", -- 6564 - 0x19a4  :  192 - 0xc0
    "11100000", -- 6565 - 0x19a5  :  224 - 0xe0
    "11100000", -- 6566 - 0x19a6  :  224 - 0xe0
    "11110000", -- 6567 - 0x19a7  :  240 - 0xf0
    "00000000", -- 6568 - 0x19a8  :    0 - 0x0
    "00000000", -- 6569 - 0x19a9  :    0 - 0x0
    "10000000", -- 6570 - 0x19aa  :  128 - 0x80
    "10000000", -- 6571 - 0x19ab  :  128 - 0x80
    "11000000", -- 6572 - 0x19ac  :  192 - 0xc0
    "11100000", -- 6573 - 0x19ad  :  224 - 0xe0
    "11100000", -- 6574 - 0x19ae  :  224 - 0xe0
    "11110000", -- 6575 - 0x19af  :  240 - 0xf0
    "11110000", -- 6576 - 0x19b0  :  240 - 0xf0 -- Background 0x9b
    "11100000", -- 6577 - 0x19b1  :  224 - 0xe0
    "11110000", -- 6578 - 0x19b2  :  240 - 0xf0
    "11100000", -- 6579 - 0x19b3  :  224 - 0xe0
    "10000000", -- 6580 - 0x19b4  :  128 - 0x80
    "00001000", -- 6581 - 0x19b5  :    8 - 0x8
    "00000100", -- 6582 - 0x19b6  :    4 - 0x4
    "00000000", -- 6583 - 0x19b7  :    0 - 0x0
    "11111111", -- 6584 - 0x19b8  :  255 - 0xff
    "11111111", -- 6585 - 0x19b9  :  255 - 0xff
    "11111100", -- 6586 - 0x19ba  :  252 - 0xfc
    "11111100", -- 6587 - 0x19bb  :  252 - 0xfc
    "11111110", -- 6588 - 0x19bc  :  254 - 0xfe
    "01111110", -- 6589 - 0x19bd  :  126 - 0x7e
    "00111111", -- 6590 - 0x19be  :   63 - 0x3f
    "00001100", -- 6591 - 0x19bf  :   12 - 0xc
    "00000000", -- 6592 - 0x19c0  :    0 - 0x0 -- Background 0x9c
    "00000000", -- 6593 - 0x19c1  :    0 - 0x0
    "00000001", -- 6594 - 0x19c2  :    1 - 0x1
    "00000011", -- 6595 - 0x19c3  :    3 - 0x3
    "00000011", -- 6596 - 0x19c4  :    3 - 0x3
    "00000011", -- 6597 - 0x19c5  :    3 - 0x3
    "00000111", -- 6598 - 0x19c6  :    7 - 0x7
    "00000111", -- 6599 - 0x19c7  :    7 - 0x7
    "00000000", -- 6600 - 0x19c8  :    0 - 0x0
    "00000001", -- 6601 - 0x19c9  :    1 - 0x1
    "00000011", -- 6602 - 0x19ca  :    3 - 0x3
    "00000111", -- 6603 - 0x19cb  :    7 - 0x7
    "00000111", -- 6604 - 0x19cc  :    7 - 0x7
    "00000111", -- 6605 - 0x19cd  :    7 - 0x7
    "00001111", -- 6606 - 0x19ce  :   15 - 0xf
    "00001111", -- 6607 - 0x19cf  :   15 - 0xf
    "00000111", -- 6608 - 0x19d0  :    7 - 0x7 -- Background 0x9d
    "00000011", -- 6609 - 0x19d1  :    3 - 0x3
    "00000011", -- 6610 - 0x19d2  :    3 - 0x3
    "00000011", -- 6611 - 0x19d3  :    3 - 0x3
    "00000011", -- 6612 - 0x19d4  :    3 - 0x3
    "00000011", -- 6613 - 0x19d5  :    3 - 0x3
    "00000011", -- 6614 - 0x19d6  :    3 - 0x3
    "00000001", -- 6615 - 0x19d7  :    1 - 0x1
    "00001111", -- 6616 - 0x19d8  :   15 - 0xf
    "00001111", -- 6617 - 0x19d9  :   15 - 0xf
    "00000111", -- 6618 - 0x19da  :    7 - 0x7
    "00000111", -- 6619 - 0x19db  :    7 - 0x7
    "00000111", -- 6620 - 0x19dc  :    7 - 0x7
    "00000011", -- 6621 - 0x19dd  :    3 - 0x3
    "00000011", -- 6622 - 0x19de  :    3 - 0x3
    "00000001", -- 6623 - 0x19df  :    1 - 0x1
    "00000000", -- 6624 - 0x19e0  :    0 - 0x0 -- Background 0x9e
    "00000000", -- 6625 - 0x19e1  :    0 - 0x0
    "00000000", -- 6626 - 0x19e2  :    0 - 0x0
    "00000000", -- 6627 - 0x19e3  :    0 - 0x0
    "00000000", -- 6628 - 0x19e4  :    0 - 0x0
    "00000001", -- 6629 - 0x19e5  :    1 - 0x1
    "00000010", -- 6630 - 0x19e6  :    2 - 0x2
    "00000100", -- 6631 - 0x19e7  :    4 - 0x4
    "00000001", -- 6632 - 0x19e8  :    1 - 0x1
    "00000001", -- 6633 - 0x19e9  :    1 - 0x1
    "00000001", -- 6634 - 0x19ea  :    1 - 0x1
    "00000000", -- 6635 - 0x19eb  :    0 - 0x0
    "00000000", -- 6636 - 0x19ec  :    0 - 0x0
    "00000011", -- 6637 - 0x19ed  :    3 - 0x3
    "00000111", -- 6638 - 0x19ee  :    7 - 0x7
    "00001111", -- 6639 - 0x19ef  :   15 - 0xf
    "00000000", -- 6640 - 0x19f0  :    0 - 0x0 -- Background 0x9f
    "00000000", -- 6641 - 0x19f1  :    0 - 0x0
    "00000000", -- 6642 - 0x19f2  :    0 - 0x0
    "00000000", -- 6643 - 0x19f3  :    0 - 0x0
    "00000000", -- 6644 - 0x19f4  :    0 - 0x0
    "00000000", -- 6645 - 0x19f5  :    0 - 0x0
    "00011100", -- 6646 - 0x19f6  :   28 - 0x1c
    "00111011", -- 6647 - 0x19f7  :   59 - 0x3b
    "00000000", -- 6648 - 0x19f8  :    0 - 0x0
    "00000000", -- 6649 - 0x19f9  :    0 - 0x0
    "00000000", -- 6650 - 0x19fa  :    0 - 0x0
    "00000000", -- 6651 - 0x19fb  :    0 - 0x0
    "00000001", -- 6652 - 0x19fc  :    1 - 0x1
    "00000011", -- 6653 - 0x19fd  :    3 - 0x3
    "00111111", -- 6654 - 0x19fe  :   63 - 0x3f
    "01111111", -- 6655 - 0x19ff  :  127 - 0x7f
    "01111110", -- 6656 - 0x1a00  :  126 - 0x7e -- Background 0xa0
    "11111110", -- 6657 - 0x1a01  :  254 - 0xfe
    "11111111", -- 6658 - 0x1a02  :  255 - 0xff
    "11111111", -- 6659 - 0x1a03  :  255 - 0xff
    "11111111", -- 6660 - 0x1a04  :  255 - 0xff
    "11111111", -- 6661 - 0x1a05  :  255 - 0xff
    "11111101", -- 6662 - 0x1a06  :  253 - 0xfd
    "11111001", -- 6663 - 0x1a07  :  249 - 0xf9
    "11111111", -- 6664 - 0x1a08  :  255 - 0xff
    "11111111", -- 6665 - 0x1a09  :  255 - 0xff
    "11111111", -- 6666 - 0x1a0a  :  255 - 0xff
    "11111111", -- 6667 - 0x1a0b  :  255 - 0xff
    "11111111", -- 6668 - 0x1a0c  :  255 - 0xff
    "11111111", -- 6669 - 0x1a0d  :  255 - 0xff
    "11111101", -- 6670 - 0x1a0e  :  253 - 0xfd
    "11111001", -- 6671 - 0x1a0f  :  249 - 0xf9
    "11110011", -- 6672 - 0x1a10  :  243 - 0xf3 -- Background 0xa1
    "11110111", -- 6673 - 0x1a11  :  247 - 0xf7
    "11110110", -- 6674 - 0x1a12  :  246 - 0xf6
    "11101110", -- 6675 - 0x1a13  :  238 - 0xee
    "11111101", -- 6676 - 0x1a14  :  253 - 0xfd
    "11111100", -- 6677 - 0x1a15  :  252 - 0xfc
    "11111000", -- 6678 - 0x1a16  :  248 - 0xf8
    "11100001", -- 6679 - 0x1a17  :  225 - 0xe1
    "11110011", -- 6680 - 0x1a18  :  243 - 0xf3
    "11111111", -- 6681 - 0x1a19  :  255 - 0xff
    "11111111", -- 6682 - 0x1a1a  :  255 - 0xff
    "11111111", -- 6683 - 0x1a1b  :  255 - 0xff
    "11111111", -- 6684 - 0x1a1c  :  255 - 0xff
    "11111111", -- 6685 - 0x1a1d  :  255 - 0xff
    "11111111", -- 6686 - 0x1a1e  :  255 - 0xff
    "11111111", -- 6687 - 0x1a1f  :  255 - 0xff
    "11010011", -- 6688 - 0x1a20  :  211 - 0xd3 -- Background 0xa2
    "11001011", -- 6689 - 0x1a21  :  203 - 0xcb
    "11000011", -- 6690 - 0x1a22  :  195 - 0xc3
    "11100001", -- 6691 - 0x1a23  :  225 - 0xe1
    "11111001", -- 6692 - 0x1a24  :  249 - 0xf9
    "00111001", -- 6693 - 0x1a25  :   57 - 0x39
    "01000010", -- 6694 - 0x1a26  :   66 - 0x42
    "00000000", -- 6695 - 0x1a27  :    0 - 0x0
    "11111111", -- 6696 - 0x1a28  :  255 - 0xff
    "11111111", -- 6697 - 0x1a29  :  255 - 0xff
    "11111111", -- 6698 - 0x1a2a  :  255 - 0xff
    "11111111", -- 6699 - 0x1a2b  :  255 - 0xff
    "11111111", -- 6700 - 0x1a2c  :  255 - 0xff
    "11111111", -- 6701 - 0x1a2d  :  255 - 0xff
    "11111111", -- 6702 - 0x1a2e  :  255 - 0xff
    "11111111", -- 6703 - 0x1a2f  :  255 - 0xff
    "00000111", -- 6704 - 0x1a30  :    7 - 0x7 -- Background 0xa3
    "00001111", -- 6705 - 0x1a31  :   15 - 0xf
    "00011001", -- 6706 - 0x1a32  :   25 - 0x19
    "00110000", -- 6707 - 0x1a33  :   48 - 0x30
    "01100011", -- 6708 - 0x1a34  :   99 - 0x63
    "01110010", -- 6709 - 0x1a35  :  114 - 0x72
    "01110000", -- 6710 - 0x1a36  :  112 - 0x70
    "00000001", -- 6711 - 0x1a37  :    1 - 0x1
    "00000111", -- 6712 - 0x1a38  :    7 - 0x7
    "00001111", -- 6713 - 0x1a39  :   15 - 0xf
    "00011111", -- 6714 - 0x1a3a  :   31 - 0x1f
    "00111111", -- 6715 - 0x1a3b  :   63 - 0x3f
    "11111100", -- 6716 - 0x1a3c  :  252 - 0xfc
    "11111100", -- 6717 - 0x1a3d  :  252 - 0xfc
    "11111111", -- 6718 - 0x1a3e  :  255 - 0xff
    "11111111", -- 6719 - 0x1a3f  :  255 - 0xff
    "00000000", -- 6720 - 0x1a40  :    0 - 0x0 -- Background 0xa4
    "00011111", -- 6721 - 0x1a41  :   31 - 0x1f
    "00100000", -- 6722 - 0x1a42  :   32 - 0x20
    "11000000", -- 6723 - 0x1a43  :  192 - 0xc0
    "11000000", -- 6724 - 0x1a44  :  192 - 0xc0
    "11110000", -- 6725 - 0x1a45  :  240 - 0xf0
    "11111111", -- 6726 - 0x1a46  :  255 - 0xff
    "11111111", -- 6727 - 0x1a47  :  255 - 0xff
    "11111111", -- 6728 - 0x1a48  :  255 - 0xff
    "11111111", -- 6729 - 0x1a49  :  255 - 0xff
    "11111111", -- 6730 - 0x1a4a  :  255 - 0xff
    "11111111", -- 6731 - 0x1a4b  :  255 - 0xff
    "11111111", -- 6732 - 0x1a4c  :  255 - 0xff
    "11111111", -- 6733 - 0x1a4d  :  255 - 0xff
    "11111111", -- 6734 - 0x1a4e  :  255 - 0xff
    "11111111", -- 6735 - 0x1a4f  :  255 - 0xff
    "10101011", -- 6736 - 0x1a50  :  171 - 0xab -- Background 0xa5
    "11000001", -- 6737 - 0x1a51  :  193 - 0xc1
    "10000001", -- 6738 - 0x1a52  :  129 - 0x81
    "10010001", -- 6739 - 0x1a53  :  145 - 0x91
    "10000010", -- 6740 - 0x1a54  :  130 - 0x82
    "11111100", -- 6741 - 0x1a55  :  252 - 0xfc
    "11100000", -- 6742 - 0x1a56  :  224 - 0xe0
    "11001110", -- 6743 - 0x1a57  :  206 - 0xce
    "11111111", -- 6744 - 0x1a58  :  255 - 0xff
    "11111111", -- 6745 - 0x1a59  :  255 - 0xff
    "11111111", -- 6746 - 0x1a5a  :  255 - 0xff
    "11111111", -- 6747 - 0x1a5b  :  255 - 0xff
    "11111111", -- 6748 - 0x1a5c  :  255 - 0xff
    "11111111", -- 6749 - 0x1a5d  :  255 - 0xff
    "11111111", -- 6750 - 0x1a5e  :  255 - 0xff
    "11111111", -- 6751 - 0x1a5f  :  255 - 0xff
    "11100101", -- 6752 - 0x1a60  :  229 - 0xe5 -- Background 0xa6
    "11011010", -- 6753 - 0x1a61  :  218 - 0xda
    "11110000", -- 6754 - 0x1a62  :  240 - 0xf0
    "11100000", -- 6755 - 0x1a63  :  224 - 0xe0
    "11000000", -- 6756 - 0x1a64  :  192 - 0xc0
    "00000000", -- 6757 - 0x1a65  :    0 - 0x0
    "00000000", -- 6758 - 0x1a66  :    0 - 0x0
    "00000000", -- 6759 - 0x1a67  :    0 - 0x0
    "11111111", -- 6760 - 0x1a68  :  255 - 0xff
    "11111111", -- 6761 - 0x1a69  :  255 - 0xff
    "11110000", -- 6762 - 0x1a6a  :  240 - 0xf0
    "11100000", -- 6763 - 0x1a6b  :  224 - 0xe0
    "11000000", -- 6764 - 0x1a6c  :  192 - 0xc0
    "10000000", -- 6765 - 0x1a6d  :  128 - 0x80
    "10000000", -- 6766 - 0x1a6e  :  128 - 0x80
    "00000000", -- 6767 - 0x1a6f  :    0 - 0x0
    "11110000", -- 6768 - 0x1a70  :  240 - 0xf0 -- Background 0xa7
    "11111000", -- 6769 - 0x1a71  :  248 - 0xf8
    "11001100", -- 6770 - 0x1a72  :  204 - 0xcc
    "10000110", -- 6771 - 0x1a73  :  134 - 0x86
    "01100010", -- 6772 - 0x1a74  :   98 - 0x62
    "00100110", -- 6773 - 0x1a75  :   38 - 0x26
    "00000110", -- 6774 - 0x1a76  :    6 - 0x6
    "11000000", -- 6775 - 0x1a77  :  192 - 0xc0
    "11110000", -- 6776 - 0x1a78  :  240 - 0xf0
    "11111000", -- 6777 - 0x1a79  :  248 - 0xf8
    "11111100", -- 6778 - 0x1a7a  :  252 - 0xfc
    "11111110", -- 6779 - 0x1a7b  :  254 - 0xfe
    "10011111", -- 6780 - 0x1a7c  :  159 - 0x9f
    "10011111", -- 6781 - 0x1a7d  :  159 - 0x9f
    "11111111", -- 6782 - 0x1a7e  :  255 - 0xff
    "11111111", -- 6783 - 0x1a7f  :  255 - 0xff
    "00000000", -- 6784 - 0x1a80  :    0 - 0x0 -- Background 0xa8
    "11111100", -- 6785 - 0x1a81  :  252 - 0xfc
    "00000110", -- 6786 - 0x1a82  :    6 - 0x6
    "00000011", -- 6787 - 0x1a83  :    3 - 0x3
    "00000001", -- 6788 - 0x1a84  :    1 - 0x1
    "00000111", -- 6789 - 0x1a85  :    7 - 0x7
    "11111111", -- 6790 - 0x1a86  :  255 - 0xff
    "11111111", -- 6791 - 0x1a87  :  255 - 0xff
    "11111111", -- 6792 - 0x1a88  :  255 - 0xff
    "11111111", -- 6793 - 0x1a89  :  255 - 0xff
    "11111111", -- 6794 - 0x1a8a  :  255 - 0xff
    "11111111", -- 6795 - 0x1a8b  :  255 - 0xff
    "11111111", -- 6796 - 0x1a8c  :  255 - 0xff
    "11111111", -- 6797 - 0x1a8d  :  255 - 0xff
    "11111111", -- 6798 - 0x1a8e  :  255 - 0xff
    "11111111", -- 6799 - 0x1a8f  :  255 - 0xff
    "11010101", -- 6800 - 0x1a90  :  213 - 0xd5 -- Background 0xa9
    "10000011", -- 6801 - 0x1a91  :  131 - 0x83
    "10000001", -- 6802 - 0x1a92  :  129 - 0x81
    "10001001", -- 6803 - 0x1a93  :  137 - 0x89
    "01000001", -- 6804 - 0x1a94  :   65 - 0x41
    "00111111", -- 6805 - 0x1a95  :   63 - 0x3f
    "00000111", -- 6806 - 0x1a96  :    7 - 0x7
    "11010011", -- 6807 - 0x1a97  :  211 - 0xd3
    "11111111", -- 6808 - 0x1a98  :  255 - 0xff
    "11111111", -- 6809 - 0x1a99  :  255 - 0xff
    "11111111", -- 6810 - 0x1a9a  :  255 - 0xff
    "11111111", -- 6811 - 0x1a9b  :  255 - 0xff
    "11111111", -- 6812 - 0x1a9c  :  255 - 0xff
    "11111111", -- 6813 - 0x1a9d  :  255 - 0xff
    "11111111", -- 6814 - 0x1a9e  :  255 - 0xff
    "11111111", -- 6815 - 0x1a9f  :  255 - 0xff
    "01101111", -- 6816 - 0x1aa0  :  111 - 0x6f -- Background 0xaa
    "11011011", -- 6817 - 0x1aa1  :  219 - 0xdb
    "00001111", -- 6818 - 0x1aa2  :   15 - 0xf
    "00000111", -- 6819 - 0x1aa3  :    7 - 0x7
    "00000011", -- 6820 - 0x1aa4  :    3 - 0x3
    "00000000", -- 6821 - 0x1aa5  :    0 - 0x0
    "00000000", -- 6822 - 0x1aa6  :    0 - 0x0
    "00000000", -- 6823 - 0x1aa7  :    0 - 0x0
    "11111111", -- 6824 - 0x1aa8  :  255 - 0xff
    "11111111", -- 6825 - 0x1aa9  :  255 - 0xff
    "00001111", -- 6826 - 0x1aaa  :   15 - 0xf
    "00000111", -- 6827 - 0x1aab  :    7 - 0x7
    "00000011", -- 6828 - 0x1aac  :    3 - 0x3
    "00000001", -- 6829 - 0x1aad  :    1 - 0x1
    "00000001", -- 6830 - 0x1aae  :    1 - 0x1
    "00000000", -- 6831 - 0x1aaf  :    0 - 0x0
    "00000000", -- 6832 - 0x1ab0  :    0 - 0x0 -- Background 0xab
    "00000000", -- 6833 - 0x1ab1  :    0 - 0x0
    "00000000", -- 6834 - 0x1ab2  :    0 - 0x0
    "00000000", -- 6835 - 0x1ab3  :    0 - 0x0
    "00000000", -- 6836 - 0x1ab4  :    0 - 0x0
    "00000000", -- 6837 - 0x1ab5  :    0 - 0x0
    "00111000", -- 6838 - 0x1ab6  :   56 - 0x38
    "11011100", -- 6839 - 0x1ab7  :  220 - 0xdc
    "00000000", -- 6840 - 0x1ab8  :    0 - 0x0
    "00000000", -- 6841 - 0x1ab9  :    0 - 0x0
    "00000000", -- 6842 - 0x1aba  :    0 - 0x0
    "00000000", -- 6843 - 0x1abb  :    0 - 0x0
    "10000000", -- 6844 - 0x1abc  :  128 - 0x80
    "11000000", -- 6845 - 0x1abd  :  192 - 0xc0
    "11111100", -- 6846 - 0x1abe  :  252 - 0xfc
    "11111110", -- 6847 - 0x1abf  :  254 - 0xfe
    "01111110", -- 6848 - 0x1ac0  :  126 - 0x7e -- Background 0xac
    "01111111", -- 6849 - 0x1ac1  :  127 - 0x7f
    "01111111", -- 6850 - 0x1ac2  :  127 - 0x7f
    "11111111", -- 6851 - 0x1ac3  :  255 - 0xff
    "11111111", -- 6852 - 0x1ac4  :  255 - 0xff
    "11111111", -- 6853 - 0x1ac5  :  255 - 0xff
    "10111111", -- 6854 - 0x1ac6  :  191 - 0xbf
    "10011111", -- 6855 - 0x1ac7  :  159 - 0x9f
    "11111111", -- 6856 - 0x1ac8  :  255 - 0xff
    "11111111", -- 6857 - 0x1ac9  :  255 - 0xff
    "11111111", -- 6858 - 0x1aca  :  255 - 0xff
    "11111111", -- 6859 - 0x1acb  :  255 - 0xff
    "11111111", -- 6860 - 0x1acc  :  255 - 0xff
    "11111111", -- 6861 - 0x1acd  :  255 - 0xff
    "10111111", -- 6862 - 0x1ace  :  191 - 0xbf
    "10011111", -- 6863 - 0x1acf  :  159 - 0x9f
    "11001111", -- 6864 - 0x1ad0  :  207 - 0xcf -- Background 0xad
    "11101111", -- 6865 - 0x1ad1  :  239 - 0xef
    "01101111", -- 6866 - 0x1ad2  :  111 - 0x6f
    "01110111", -- 6867 - 0x1ad3  :  119 - 0x77
    "10111111", -- 6868 - 0x1ad4  :  191 - 0xbf
    "00111111", -- 6869 - 0x1ad5  :   63 - 0x3f
    "00011111", -- 6870 - 0x1ad6  :   31 - 0x1f
    "10000111", -- 6871 - 0x1ad7  :  135 - 0x87
    "11001111", -- 6872 - 0x1ad8  :  207 - 0xcf
    "11111111", -- 6873 - 0x1ad9  :  255 - 0xff
    "11111111", -- 6874 - 0x1ada  :  255 - 0xff
    "11111111", -- 6875 - 0x1adb  :  255 - 0xff
    "11111111", -- 6876 - 0x1adc  :  255 - 0xff
    "11111111", -- 6877 - 0x1add  :  255 - 0xff
    "11111111", -- 6878 - 0x1ade  :  255 - 0xff
    "11111111", -- 6879 - 0x1adf  :  255 - 0xff
    "11001011", -- 6880 - 0x1ae0  :  203 - 0xcb -- Background 0xae
    "11010011", -- 6881 - 0x1ae1  :  211 - 0xd3
    "11000011", -- 6882 - 0x1ae2  :  195 - 0xc3
    "10000111", -- 6883 - 0x1ae3  :  135 - 0x87
    "10011111", -- 6884 - 0x1ae4  :  159 - 0x9f
    "10011100", -- 6885 - 0x1ae5  :  156 - 0x9c
    "01000010", -- 6886 - 0x1ae6  :   66 - 0x42
    "00000000", -- 6887 - 0x1ae7  :    0 - 0x0
    "11111111", -- 6888 - 0x1ae8  :  255 - 0xff
    "11111111", -- 6889 - 0x1ae9  :  255 - 0xff
    "11111111", -- 6890 - 0x1aea  :  255 - 0xff
    "11111111", -- 6891 - 0x1aeb  :  255 - 0xff
    "11111111", -- 6892 - 0x1aec  :  255 - 0xff
    "11111111", -- 6893 - 0x1aed  :  255 - 0xff
    "11111111", -- 6894 - 0x1aee  :  255 - 0xff
    "11111111", -- 6895 - 0x1aef  :  255 - 0xff
    "00000000", -- 6896 - 0x1af0  :    0 - 0x0 -- Background 0xaf
    "00000000", -- 6897 - 0x1af1  :    0 - 0x0
    "10000000", -- 6898 - 0x1af2  :  128 - 0x80
    "11000000", -- 6899 - 0x1af3  :  192 - 0xc0
    "11000000", -- 6900 - 0x1af4  :  192 - 0xc0
    "11000000", -- 6901 - 0x1af5  :  192 - 0xc0
    "11100000", -- 6902 - 0x1af6  :  224 - 0xe0
    "11100000", -- 6903 - 0x1af7  :  224 - 0xe0
    "00000000", -- 6904 - 0x1af8  :    0 - 0x0
    "10000000", -- 6905 - 0x1af9  :  128 - 0x80
    "11000000", -- 6906 - 0x1afa  :  192 - 0xc0
    "11100000", -- 6907 - 0x1afb  :  224 - 0xe0
    "11100000", -- 6908 - 0x1afc  :  224 - 0xe0
    "11100000", -- 6909 - 0x1afd  :  224 - 0xe0
    "11110000", -- 6910 - 0x1afe  :  240 - 0xf0
    "11110000", -- 6911 - 0x1aff  :  240 - 0xf0
    "11100000", -- 6912 - 0x1b00  :  224 - 0xe0 -- Background 0xb0
    "11000000", -- 6913 - 0x1b01  :  192 - 0xc0
    "11000000", -- 6914 - 0x1b02  :  192 - 0xc0
    "11000000", -- 6915 - 0x1b03  :  192 - 0xc0
    "11000000", -- 6916 - 0x1b04  :  192 - 0xc0
    "11000000", -- 6917 - 0x1b05  :  192 - 0xc0
    "11000000", -- 6918 - 0x1b06  :  192 - 0xc0
    "10000000", -- 6919 - 0x1b07  :  128 - 0x80
    "11110000", -- 6920 - 0x1b08  :  240 - 0xf0
    "11110000", -- 6921 - 0x1b09  :  240 - 0xf0
    "11100000", -- 6922 - 0x1b0a  :  224 - 0xe0
    "11100000", -- 6923 - 0x1b0b  :  224 - 0xe0
    "11100000", -- 6924 - 0x1b0c  :  224 - 0xe0
    "11000000", -- 6925 - 0x1b0d  :  192 - 0xc0
    "11000000", -- 6926 - 0x1b0e  :  192 - 0xc0
    "10000000", -- 6927 - 0x1b0f  :  128 - 0x80
    "00000000", -- 6928 - 0x1b10  :    0 - 0x0 -- Background 0xb1
    "00000000", -- 6929 - 0x1b11  :    0 - 0x0
    "00000000", -- 6930 - 0x1b12  :    0 - 0x0
    "00000000", -- 6931 - 0x1b13  :    0 - 0x0
    "00000000", -- 6932 - 0x1b14  :    0 - 0x0
    "10000000", -- 6933 - 0x1b15  :  128 - 0x80
    "01000000", -- 6934 - 0x1b16  :   64 - 0x40
    "00100000", -- 6935 - 0x1b17  :   32 - 0x20
    "10000000", -- 6936 - 0x1b18  :  128 - 0x80
    "10000000", -- 6937 - 0x1b19  :  128 - 0x80
    "10000000", -- 6938 - 0x1b1a  :  128 - 0x80
    "00000000", -- 6939 - 0x1b1b  :    0 - 0x0
    "00000000", -- 6940 - 0x1b1c  :    0 - 0x0
    "11000000", -- 6941 - 0x1b1d  :  192 - 0xc0
    "11100000", -- 6942 - 0x1b1e  :  224 - 0xe0
    "11110000", -- 6943 - 0x1b1f  :  240 - 0xf0
    "00000000", -- 6944 - 0x1b20  :    0 - 0x0 -- Background 0xb2
    "00000000", -- 6945 - 0x1b21  :    0 - 0x0
    "00000000", -- 6946 - 0x1b22  :    0 - 0x0
    "00000001", -- 6947 - 0x1b23  :    1 - 0x1
    "00000011", -- 6948 - 0x1b24  :    3 - 0x3
    "00000111", -- 6949 - 0x1b25  :    7 - 0x7
    "00000111", -- 6950 - 0x1b26  :    7 - 0x7
    "00000111", -- 6951 - 0x1b27  :    7 - 0x7
    "00000000", -- 6952 - 0x1b28  :    0 - 0x0
    "00000000", -- 6953 - 0x1b29  :    0 - 0x0
    "00000001", -- 6954 - 0x1b2a  :    1 - 0x1
    "00000011", -- 6955 - 0x1b2b  :    3 - 0x3
    "00000111", -- 6956 - 0x1b2c  :    7 - 0x7
    "00000111", -- 6957 - 0x1b2d  :    7 - 0x7
    "00000111", -- 6958 - 0x1b2e  :    7 - 0x7
    "00000111", -- 6959 - 0x1b2f  :    7 - 0x7
    "00000011", -- 6960 - 0x1b30  :    3 - 0x3 -- Background 0xb3
    "00000001", -- 6961 - 0x1b31  :    1 - 0x1
    "00000000", -- 6962 - 0x1b32  :    0 - 0x0
    "00000000", -- 6963 - 0x1b33  :    0 - 0x0
    "00000000", -- 6964 - 0x1b34  :    0 - 0x0
    "00000000", -- 6965 - 0x1b35  :    0 - 0x0
    "00000001", -- 6966 - 0x1b36  :    1 - 0x1
    "00000001", -- 6967 - 0x1b37  :    1 - 0x1
    "00000011", -- 6968 - 0x1b38  :    3 - 0x3
    "00000001", -- 6969 - 0x1b39  :    1 - 0x1
    "00000000", -- 6970 - 0x1b3a  :    0 - 0x0
    "00000000", -- 6971 - 0x1b3b  :    0 - 0x0
    "00000000", -- 6972 - 0x1b3c  :    0 - 0x0
    "00000001", -- 6973 - 0x1b3d  :    1 - 0x1
    "00000011", -- 6974 - 0x1b3e  :    3 - 0x3
    "00000011", -- 6975 - 0x1b3f  :    3 - 0x3
    "00000001", -- 6976 - 0x1b40  :    1 - 0x1 -- Background 0xb4
    "00000001", -- 6977 - 0x1b41  :    1 - 0x1
    "00000111", -- 6978 - 0x1b42  :    7 - 0x7
    "00000011", -- 6979 - 0x1b43  :    3 - 0x3
    "00000100", -- 6980 - 0x1b44  :    4 - 0x4
    "00000000", -- 6981 - 0x1b45  :    0 - 0x0
    "00000000", -- 6982 - 0x1b46  :    0 - 0x0
    "00000000", -- 6983 - 0x1b47  :    0 - 0x0
    "00000011", -- 6984 - 0x1b48  :    3 - 0x3
    "00000011", -- 6985 - 0x1b49  :    3 - 0x3
    "00000111", -- 6986 - 0x1b4a  :    7 - 0x7
    "00011111", -- 6987 - 0x1b4b  :   31 - 0x1f
    "00111111", -- 6988 - 0x1b4c  :   63 - 0x3f
    "00111111", -- 6989 - 0x1b4d  :   63 - 0x3f
    "00000000", -- 6990 - 0x1b4e  :    0 - 0x0
    "00000000", -- 6991 - 0x1b4f  :    0 - 0x0
    "00000000", -- 6992 - 0x1b50  :    0 - 0x0 -- Background 0xb5
    "00000000", -- 6993 - 0x1b51  :    0 - 0x0
    "00000000", -- 6994 - 0x1b52  :    0 - 0x0
    "00000000", -- 6995 - 0x1b53  :    0 - 0x0
    "00000000", -- 6996 - 0x1b54  :    0 - 0x0
    "00000000", -- 6997 - 0x1b55  :    0 - 0x0
    "00000000", -- 6998 - 0x1b56  :    0 - 0x0
    "00000111", -- 6999 - 0x1b57  :    7 - 0x7
    "00000000", -- 7000 - 0x1b58  :    0 - 0x0
    "00000000", -- 7001 - 0x1b59  :    0 - 0x0
    "00000000", -- 7002 - 0x1b5a  :    0 - 0x0
    "00000000", -- 7003 - 0x1b5b  :    0 - 0x0
    "00000001", -- 7004 - 0x1b5c  :    1 - 0x1
    "00000011", -- 7005 - 0x1b5d  :    3 - 0x3
    "00000011", -- 7006 - 0x1b5e  :    3 - 0x3
    "00001111", -- 7007 - 0x1b5f  :   15 - 0xf
    "00001110", -- 7008 - 0x1b60  :   14 - 0xe -- Background 0xb6
    "00111110", -- 7009 - 0x1b61  :   62 - 0x3e
    "01111111", -- 7010 - 0x1b62  :  127 - 0x7f
    "11111111", -- 7011 - 0x1b63  :  255 - 0xff
    "11111111", -- 7012 - 0x1b64  :  255 - 0xff
    "11101111", -- 7013 - 0x1b65  :  239 - 0xef
    "11110111", -- 7014 - 0x1b66  :  247 - 0xf7
    "11111000", -- 7015 - 0x1b67  :  248 - 0xf8
    "00111111", -- 7016 - 0x1b68  :   63 - 0x3f
    "01111111", -- 7017 - 0x1b69  :  127 - 0x7f
    "11111111", -- 7018 - 0x1b6a  :  255 - 0xff
    "11111111", -- 7019 - 0x1b6b  :  255 - 0xff
    "11111111", -- 7020 - 0x1b6c  :  255 - 0xff
    "11111111", -- 7021 - 0x1b6d  :  255 - 0xff
    "11111111", -- 7022 - 0x1b6e  :  255 - 0xff
    "11111111", -- 7023 - 0x1b6f  :  255 - 0xff
    "11111111", -- 7024 - 0x1b70  :  255 - 0xff -- Background 0xb7
    "11111111", -- 7025 - 0x1b71  :  255 - 0xff
    "11111111", -- 7026 - 0x1b72  :  255 - 0xff
    "00011111", -- 7027 - 0x1b73  :   31 - 0x1f
    "00011111", -- 7028 - 0x1b74  :   31 - 0x1f
    "01111111", -- 7029 - 0x1b75  :  127 - 0x7f
    "11111111", -- 7030 - 0x1b76  :  255 - 0xff
    "11111110", -- 7031 - 0x1b77  :  254 - 0xfe
    "11111111", -- 7032 - 0x1b78  :  255 - 0xff
    "11111111", -- 7033 - 0x1b79  :  255 - 0xff
    "11111111", -- 7034 - 0x1b7a  :  255 - 0xff
    "00011111", -- 7035 - 0x1b7b  :   31 - 0x1f
    "01111111", -- 7036 - 0x1b7c  :  127 - 0x7f
    "11111111", -- 7037 - 0x1b7d  :  255 - 0xff
    "11111111", -- 7038 - 0x1b7e  :  255 - 0xff
    "11111111", -- 7039 - 0x1b7f  :  255 - 0xff
    "11111111", -- 7040 - 0x1b80  :  255 - 0xff -- Background 0xb8
    "11111111", -- 7041 - 0x1b81  :  255 - 0xff
    "11111111", -- 7042 - 0x1b82  :  255 - 0xff
    "11111100", -- 7043 - 0x1b83  :  252 - 0xfc
    "11111000", -- 7044 - 0x1b84  :  248 - 0xf8
    "10000000", -- 7045 - 0x1b85  :  128 - 0x80
    "00000000", -- 7046 - 0x1b86  :    0 - 0x0
    "00000000", -- 7047 - 0x1b87  :    0 - 0x0
    "11111111", -- 7048 - 0x1b88  :  255 - 0xff
    "11111111", -- 7049 - 0x1b89  :  255 - 0xff
    "11111111", -- 7050 - 0x1b8a  :  255 - 0xff
    "11111100", -- 7051 - 0x1b8b  :  252 - 0xfc
    "11111000", -- 7052 - 0x1b8c  :  248 - 0xf8
    "11111000", -- 7053 - 0x1b8d  :  248 - 0xf8
    "00000000", -- 7054 - 0x1b8e  :    0 - 0x0
    "00000000", -- 7055 - 0x1b8f  :    0 - 0x0
    "00110000", -- 7056 - 0x1b90  :   48 - 0x30 -- Background 0xb9
    "01111111", -- 7057 - 0x1b91  :  127 - 0x7f
    "01111111", -- 7058 - 0x1b92  :  127 - 0x7f
    "00111111", -- 7059 - 0x1b93  :   63 - 0x3f
    "10000111", -- 7060 - 0x1b94  :  135 - 0x87
    "11110000", -- 7061 - 0x1b95  :  240 - 0xf0
    "11111111", -- 7062 - 0x1b96  :  255 - 0xff
    "11111111", -- 7063 - 0x1b97  :  255 - 0xff
    "11001111", -- 7064 - 0x1b98  :  207 - 0xcf
    "10001000", -- 7065 - 0x1b99  :  136 - 0x88
    "11011101", -- 7066 - 0x1b9a  :  221 - 0xdd
    "11001000", -- 7067 - 0x1b9b  :  200 - 0xc8
    "11111000", -- 7068 - 0x1b9c  :  248 - 0xf8
    "11111111", -- 7069 - 0x1b9d  :  255 - 0xff
    "11111111", -- 7070 - 0x1b9e  :  255 - 0xff
    "11111111", -- 7071 - 0x1b9f  :  255 - 0xff
    "11100101", -- 7072 - 0x1ba0  :  229 - 0xe5 -- Background 0xba
    "11011010", -- 7073 - 0x1ba1  :  218 - 0xda
    "11000000", -- 7074 - 0x1ba2  :  192 - 0xc0
    "00000000", -- 7075 - 0x1ba3  :    0 - 0x0
    "00000000", -- 7076 - 0x1ba4  :    0 - 0x0
    "00000000", -- 7077 - 0x1ba5  :    0 - 0x0
    "00000000", -- 7078 - 0x1ba6  :    0 - 0x0
    "00000000", -- 7079 - 0x1ba7  :    0 - 0x0
    "11111111", -- 7080 - 0x1ba8  :  255 - 0xff
    "11111111", -- 7081 - 0x1ba9  :  255 - 0xff
    "11000000", -- 7082 - 0x1baa  :  192 - 0xc0
    "00000000", -- 7083 - 0x1bab  :    0 - 0x0
    "00000000", -- 7084 - 0x1bac  :    0 - 0x0
    "00000000", -- 7085 - 0x1bad  :    0 - 0x0
    "00000000", -- 7086 - 0x1bae  :    0 - 0x0
    "00000000", -- 7087 - 0x1baf  :    0 - 0x0
    "00000110", -- 7088 - 0x1bb0  :    6 - 0x6 -- Background 0xbb
    "11111111", -- 7089 - 0x1bb1  :  255 - 0xff
    "11111111", -- 7090 - 0x1bb2  :  255 - 0xff
    "11111110", -- 7091 - 0x1bb3  :  254 - 0xfe
    "11110001", -- 7092 - 0x1bb4  :  241 - 0xf1
    "00000111", -- 7093 - 0x1bb5  :    7 - 0x7
    "11111111", -- 7094 - 0x1bb6  :  255 - 0xff
    "11111111", -- 7095 - 0x1bb7  :  255 - 0xff
    "11111001", -- 7096 - 0x1bb8  :  249 - 0xf9
    "10001000", -- 7097 - 0x1bb9  :  136 - 0x88
    "11011101", -- 7098 - 0x1bba  :  221 - 0xdd
    "10001001", -- 7099 - 0x1bbb  :  137 - 0x89
    "00001111", -- 7100 - 0x1bbc  :   15 - 0xf
    "11111111", -- 7101 - 0x1bbd  :  255 - 0xff
    "11111111", -- 7102 - 0x1bbe  :  255 - 0xff
    "11111111", -- 7103 - 0x1bbf  :  255 - 0xff
    "00000000", -- 7104 - 0x1bc0  :    0 - 0x0 -- Background 0xbc
    "00000001", -- 7105 - 0x1bc1  :    1 - 0x1
    "00000010", -- 7106 - 0x1bc2  :    2 - 0x2
    "00000111", -- 7107 - 0x1bc3  :    7 - 0x7
    "00000000", -- 7108 - 0x1bc4  :    0 - 0x0
    "00000000", -- 7109 - 0x1bc5  :    0 - 0x0
    "00100000", -- 7110 - 0x1bc6  :   32 - 0x20
    "11111111", -- 7111 - 0x1bc7  :  255 - 0xff
    "00000011", -- 7112 - 0x1bc8  :    3 - 0x3
    "00000111", -- 7113 - 0x1bc9  :    7 - 0x7
    "00001111", -- 7114 - 0x1bca  :   15 - 0xf
    "00000111", -- 7115 - 0x1bcb  :    7 - 0x7
    "10000111", -- 7116 - 0x1bcc  :  135 - 0x87
    "11000011", -- 7117 - 0x1bcd  :  195 - 0xc3
    "11100000", -- 7118 - 0x1bce  :  224 - 0xe0
    "11111111", -- 7119 - 0x1bcf  :  255 - 0xff
    "01111111", -- 7120 - 0x1bd0  :  127 - 0x7f -- Background 0xbd
    "01111111", -- 7121 - 0x1bd1  :  127 - 0x7f
    "01111111", -- 7122 - 0x1bd2  :  127 - 0x7f
    "11111111", -- 7123 - 0x1bd3  :  255 - 0xff
    "11111111", -- 7124 - 0x1bd4  :  255 - 0xff
    "11111111", -- 7125 - 0x1bd5  :  255 - 0xff
    "11111111", -- 7126 - 0x1bd6  :  255 - 0xff
    "11111110", -- 7127 - 0x1bd7  :  254 - 0xfe
    "11111111", -- 7128 - 0x1bd8  :  255 - 0xff
    "11111111", -- 7129 - 0x1bd9  :  255 - 0xff
    "11111111", -- 7130 - 0x1bda  :  255 - 0xff
    "11111111", -- 7131 - 0x1bdb  :  255 - 0xff
    "11111111", -- 7132 - 0x1bdc  :  255 - 0xff
    "11111111", -- 7133 - 0x1bdd  :  255 - 0xff
    "11111111", -- 7134 - 0x1bde  :  255 - 0xff
    "11111110", -- 7135 - 0x1bdf  :  254 - 0xfe
    "11111100", -- 7136 - 0x1be0  :  252 - 0xfc -- Background 0xbe
    "10111000", -- 7137 - 0x1be1  :  184 - 0xb8
    "01111000", -- 7138 - 0x1be2  :  120 - 0x78
    "01111000", -- 7139 - 0x1be3  :  120 - 0x78
    "10110000", -- 7140 - 0x1be4  :  176 - 0xb0
    "01111000", -- 7141 - 0x1be5  :  120 - 0x78
    "11111100", -- 7142 - 0x1be6  :  252 - 0xfc
    "11111110", -- 7143 - 0x1be7  :  254 - 0xfe
    "11111100", -- 7144 - 0x1be8  :  252 - 0xfc
    "11111000", -- 7145 - 0x1be9  :  248 - 0xf8
    "11111000", -- 7146 - 0x1bea  :  248 - 0xf8
    "11111000", -- 7147 - 0x1beb  :  248 - 0xf8
    "11111000", -- 7148 - 0x1bec  :  248 - 0xf8
    "11111100", -- 7149 - 0x1bed  :  252 - 0xfc
    "11111110", -- 7150 - 0x1bee  :  254 - 0xfe
    "11111111", -- 7151 - 0x1bef  :  255 - 0xff
    "11111111", -- 7152 - 0x1bf0  :  255 - 0xff -- Background 0xbf
    "11111111", -- 7153 - 0x1bf1  :  255 - 0xff
    "11111111", -- 7154 - 0x1bf2  :  255 - 0xff
    "11111111", -- 7155 - 0x1bf3  :  255 - 0xff
    "11111111", -- 7156 - 0x1bf4  :  255 - 0xff
    "10011100", -- 7157 - 0x1bf5  :  156 - 0x9c
    "01000010", -- 7158 - 0x1bf6  :   66 - 0x42
    "00000000", -- 7159 - 0x1bf7  :    0 - 0x0
    "11111111", -- 7160 - 0x1bf8  :  255 - 0xff
    "11111111", -- 7161 - 0x1bf9  :  255 - 0xff
    "11111111", -- 7162 - 0x1bfa  :  255 - 0xff
    "11111111", -- 7163 - 0x1bfb  :  255 - 0xff
    "11111111", -- 7164 - 0x1bfc  :  255 - 0xff
    "11111111", -- 7165 - 0x1bfd  :  255 - 0xff
    "11111111", -- 7166 - 0x1bfe  :  255 - 0xff
    "11111111", -- 7167 - 0x1bff  :  255 - 0xff
    "00000000", -- 7168 - 0x1c00  :    0 - 0x0 -- Background 0xc0
    "00000000", -- 7169 - 0x1c01  :    0 - 0x0
    "00100000", -- 7170 - 0x1c02  :   32 - 0x20
    "01000000", -- 7171 - 0x1c03  :   64 - 0x40
    "10001010", -- 7172 - 0x1c04  :  138 - 0x8a
    "00011110", -- 7173 - 0x1c05  :   30 - 0x1e
    "01111110", -- 7174 - 0x1c06  :  126 - 0x7e
    "10111110", -- 7175 - 0x1c07  :  190 - 0xbe
    "11000000", -- 7176 - 0x1c08  :  192 - 0xc0
    "11110000", -- 7177 - 0x1c09  :  240 - 0xf0
    "11111100", -- 7178 - 0x1c0a  :  252 - 0xfc
    "11111100", -- 7179 - 0x1c0b  :  252 - 0xfc
    "11111110", -- 7180 - 0x1c0c  :  254 - 0xfe
    "11111110", -- 7181 - 0x1c0d  :  254 - 0xfe
    "11111110", -- 7182 - 0x1c0e  :  254 - 0xfe
    "11111110", -- 7183 - 0x1c0f  :  254 - 0xfe
    "11011111", -- 7184 - 0x1c10  :  223 - 0xdf -- Background 0xc1
    "11111111", -- 7185 - 0x1c11  :  255 - 0xff
    "11111110", -- 7186 - 0x1c12  :  254 - 0xfe
    "11111100", -- 7187 - 0x1c13  :  252 - 0xfc
    "11110000", -- 7188 - 0x1c14  :  240 - 0xf0
    "11100000", -- 7189 - 0x1c15  :  224 - 0xe0
    "10000000", -- 7190 - 0x1c16  :  128 - 0x80
    "00000000", -- 7191 - 0x1c17  :    0 - 0x0
    "11111111", -- 7192 - 0x1c18  :  255 - 0xff
    "11111111", -- 7193 - 0x1c19  :  255 - 0xff
    "11111110", -- 7194 - 0x1c1a  :  254 - 0xfe
    "11111100", -- 7195 - 0x1c1b  :  252 - 0xfc
    "11110000", -- 7196 - 0x1c1c  :  240 - 0xf0
    "11100000", -- 7197 - 0x1c1d  :  224 - 0xe0
    "10000000", -- 7198 - 0x1c1e  :  128 - 0x80
    "00000000", -- 7199 - 0x1c1f  :    0 - 0x0
    "00000000", -- 7200 - 0x1c20  :    0 - 0x0 -- Background 0xc2
    "00000000", -- 7201 - 0x1c21  :    0 - 0x0
    "00000100", -- 7202 - 0x1c22  :    4 - 0x4
    "00000010", -- 7203 - 0x1c23  :    2 - 0x2
    "01010001", -- 7204 - 0x1c24  :   81 - 0x51
    "01111000", -- 7205 - 0x1c25  :  120 - 0x78
    "01111110", -- 7206 - 0x1c26  :  126 - 0x7e
    "11111101", -- 7207 - 0x1c27  :  253 - 0xfd
    "00000011", -- 7208 - 0x1c28  :    3 - 0x3
    "00001111", -- 7209 - 0x1c29  :   15 - 0xf
    "00111111", -- 7210 - 0x1c2a  :   63 - 0x3f
    "00111111", -- 7211 - 0x1c2b  :   63 - 0x3f
    "01111111", -- 7212 - 0x1c2c  :  127 - 0x7f
    "01111111", -- 7213 - 0x1c2d  :  127 - 0x7f
    "01111110", -- 7214 - 0x1c2e  :  126 - 0x7e
    "11111111", -- 7215 - 0x1c2f  :  255 - 0xff
    "11111011", -- 7216 - 0x1c30  :  251 - 0xfb -- Background 0xc3
    "11111111", -- 7217 - 0x1c31  :  255 - 0xff
    "01111111", -- 7218 - 0x1c32  :  127 - 0x7f
    "00111111", -- 7219 - 0x1c33  :   63 - 0x3f
    "00001111", -- 7220 - 0x1c34  :   15 - 0xf
    "00000111", -- 7221 - 0x1c35  :    7 - 0x7
    "00000001", -- 7222 - 0x1c36  :    1 - 0x1
    "00000000", -- 7223 - 0x1c37  :    0 - 0x0
    "11111111", -- 7224 - 0x1c38  :  255 - 0xff
    "11111111", -- 7225 - 0x1c39  :  255 - 0xff
    "01111111", -- 7226 - 0x1c3a  :  127 - 0x7f
    "00111111", -- 7227 - 0x1c3b  :   63 - 0x3f
    "00001111", -- 7228 - 0x1c3c  :   15 - 0xf
    "00000111", -- 7229 - 0x1c3d  :    7 - 0x7
    "00000001", -- 7230 - 0x1c3e  :    1 - 0x1
    "00000000", -- 7231 - 0x1c3f  :    0 - 0x0
    "00000000", -- 7232 - 0x1c40  :    0 - 0x0 -- Background 0xc4
    "10000000", -- 7233 - 0x1c41  :  128 - 0x80
    "01000000", -- 7234 - 0x1c42  :   64 - 0x40
    "11100000", -- 7235 - 0x1c43  :  224 - 0xe0
    "00000000", -- 7236 - 0x1c44  :    0 - 0x0
    "00000000", -- 7237 - 0x1c45  :    0 - 0x0
    "00000100", -- 7238 - 0x1c46  :    4 - 0x4
    "11111111", -- 7239 - 0x1c47  :  255 - 0xff
    "11000000", -- 7240 - 0x1c48  :  192 - 0xc0
    "11100000", -- 7241 - 0x1c49  :  224 - 0xe0
    "11110000", -- 7242 - 0x1c4a  :  240 - 0xf0
    "11100000", -- 7243 - 0x1c4b  :  224 - 0xe0
    "11100001", -- 7244 - 0x1c4c  :  225 - 0xe1
    "11000011", -- 7245 - 0x1c4d  :  195 - 0xc3
    "00000111", -- 7246 - 0x1c4e  :    7 - 0x7
    "11111111", -- 7247 - 0x1c4f  :  255 - 0xff
    "11111110", -- 7248 - 0x1c50  :  254 - 0xfe -- Background 0xc5
    "11111110", -- 7249 - 0x1c51  :  254 - 0xfe
    "11111110", -- 7250 - 0x1c52  :  254 - 0xfe
    "11111111", -- 7251 - 0x1c53  :  255 - 0xff
    "11111111", -- 7252 - 0x1c54  :  255 - 0xff
    "11111111", -- 7253 - 0x1c55  :  255 - 0xff
    "11111111", -- 7254 - 0x1c56  :  255 - 0xff
    "01111111", -- 7255 - 0x1c57  :  127 - 0x7f
    "11111111", -- 7256 - 0x1c58  :  255 - 0xff
    "11111111", -- 7257 - 0x1c59  :  255 - 0xff
    "11111111", -- 7258 - 0x1c5a  :  255 - 0xff
    "11111111", -- 7259 - 0x1c5b  :  255 - 0xff
    "11111111", -- 7260 - 0x1c5c  :  255 - 0xff
    "11111111", -- 7261 - 0x1c5d  :  255 - 0xff
    "11111111", -- 7262 - 0x1c5e  :  255 - 0xff
    "01111111", -- 7263 - 0x1c5f  :  127 - 0x7f
    "00111111", -- 7264 - 0x1c60  :   63 - 0x3f -- Background 0xc6
    "00011101", -- 7265 - 0x1c61  :   29 - 0x1d
    "00011110", -- 7266 - 0x1c62  :   30 - 0x1e
    "00011110", -- 7267 - 0x1c63  :   30 - 0x1e
    "00001101", -- 7268 - 0x1c64  :   13 - 0xd
    "00011110", -- 7269 - 0x1c65  :   30 - 0x1e
    "00111111", -- 7270 - 0x1c66  :   63 - 0x3f
    "01111111", -- 7271 - 0x1c67  :  127 - 0x7f
    "00111111", -- 7272 - 0x1c68  :   63 - 0x3f
    "00011111", -- 7273 - 0x1c69  :   31 - 0x1f
    "00011111", -- 7274 - 0x1c6a  :   31 - 0x1f
    "00011111", -- 7275 - 0x1c6b  :   31 - 0x1f
    "00011111", -- 7276 - 0x1c6c  :   31 - 0x1f
    "00111111", -- 7277 - 0x1c6d  :   63 - 0x3f
    "01111111", -- 7278 - 0x1c6e  :  127 - 0x7f
    "11111111", -- 7279 - 0x1c6f  :  255 - 0xff
    "11111111", -- 7280 - 0x1c70  :  255 - 0xff -- Background 0xc7
    "11111111", -- 7281 - 0x1c71  :  255 - 0xff
    "11111111", -- 7282 - 0x1c72  :  255 - 0xff
    "11111111", -- 7283 - 0x1c73  :  255 - 0xff
    "11111111", -- 7284 - 0x1c74  :  255 - 0xff
    "00111001", -- 7285 - 0x1c75  :   57 - 0x39
    "01000010", -- 7286 - 0x1c76  :   66 - 0x42
    "00000000", -- 7287 - 0x1c77  :    0 - 0x0
    "11111111", -- 7288 - 0x1c78  :  255 - 0xff
    "11111111", -- 7289 - 0x1c79  :  255 - 0xff
    "11111111", -- 7290 - 0x1c7a  :  255 - 0xff
    "11111111", -- 7291 - 0x1c7b  :  255 - 0xff
    "11111111", -- 7292 - 0x1c7c  :  255 - 0xff
    "11111111", -- 7293 - 0x1c7d  :  255 - 0xff
    "11111111", -- 7294 - 0x1c7e  :  255 - 0xff
    "11111111", -- 7295 - 0x1c7f  :  255 - 0xff
    "01101111", -- 7296 - 0x1c80  :  111 - 0x6f -- Background 0xc8
    "11011011", -- 7297 - 0x1c81  :  219 - 0xdb
    "00000011", -- 7298 - 0x1c82  :    3 - 0x3
    "00000000", -- 7299 - 0x1c83  :    0 - 0x0
    "00000000", -- 7300 - 0x1c84  :    0 - 0x0
    "00000000", -- 7301 - 0x1c85  :    0 - 0x0
    "00000000", -- 7302 - 0x1c86  :    0 - 0x0
    "00000000", -- 7303 - 0x1c87  :    0 - 0x0
    "11111111", -- 7304 - 0x1c88  :  255 - 0xff
    "11111111", -- 7305 - 0x1c89  :  255 - 0xff
    "00000011", -- 7306 - 0x1c8a  :    3 - 0x3
    "00000000", -- 7307 - 0x1c8b  :    0 - 0x0
    "00000000", -- 7308 - 0x1c8c  :    0 - 0x0
    "00000000", -- 7309 - 0x1c8d  :    0 - 0x0
    "00000000", -- 7310 - 0x1c8e  :    0 - 0x0
    "00000000", -- 7311 - 0x1c8f  :    0 - 0x0
    "00000000", -- 7312 - 0x1c90  :    0 - 0x0 -- Background 0xc9
    "00000000", -- 7313 - 0x1c91  :    0 - 0x0
    "00000000", -- 7314 - 0x1c92  :    0 - 0x0
    "00000000", -- 7315 - 0x1c93  :    0 - 0x0
    "00000000", -- 7316 - 0x1c94  :    0 - 0x0
    "00000000", -- 7317 - 0x1c95  :    0 - 0x0
    "00000000", -- 7318 - 0x1c96  :    0 - 0x0
    "11100000", -- 7319 - 0x1c97  :  224 - 0xe0
    "00000000", -- 7320 - 0x1c98  :    0 - 0x0
    "00000000", -- 7321 - 0x1c99  :    0 - 0x0
    "00000000", -- 7322 - 0x1c9a  :    0 - 0x0
    "00000000", -- 7323 - 0x1c9b  :    0 - 0x0
    "10000000", -- 7324 - 0x1c9c  :  128 - 0x80
    "11000000", -- 7325 - 0x1c9d  :  192 - 0xc0
    "11000000", -- 7326 - 0x1c9e  :  192 - 0xc0
    "11110000", -- 7327 - 0x1c9f  :  240 - 0xf0
    "01110000", -- 7328 - 0x1ca0  :  112 - 0x70 -- Background 0xca
    "01111100", -- 7329 - 0x1ca1  :  124 - 0x7c
    "01111110", -- 7330 - 0x1ca2  :  126 - 0x7e
    "11111111", -- 7331 - 0x1ca3  :  255 - 0xff
    "11111111", -- 7332 - 0x1ca4  :  255 - 0xff
    "11110111", -- 7333 - 0x1ca5  :  247 - 0xf7
    "11101111", -- 7334 - 0x1ca6  :  239 - 0xef
    "00011111", -- 7335 - 0x1ca7  :   31 - 0x1f
    "11111100", -- 7336 - 0x1ca8  :  252 - 0xfc
    "11111110", -- 7337 - 0x1ca9  :  254 - 0xfe
    "11111111", -- 7338 - 0x1caa  :  255 - 0xff
    "11111111", -- 7339 - 0x1cab  :  255 - 0xff
    "11111111", -- 7340 - 0x1cac  :  255 - 0xff
    "11111111", -- 7341 - 0x1cad  :  255 - 0xff
    "11111111", -- 7342 - 0x1cae  :  255 - 0xff
    "11111111", -- 7343 - 0x1caf  :  255 - 0xff
    "11111111", -- 7344 - 0x1cb0  :  255 - 0xff -- Background 0xcb
    "11111111", -- 7345 - 0x1cb1  :  255 - 0xff
    "11111111", -- 7346 - 0x1cb2  :  255 - 0xff
    "11111000", -- 7347 - 0x1cb3  :  248 - 0xf8
    "11111000", -- 7348 - 0x1cb4  :  248 - 0xf8
    "11111110", -- 7349 - 0x1cb5  :  254 - 0xfe
    "11111111", -- 7350 - 0x1cb6  :  255 - 0xff
    "11111111", -- 7351 - 0x1cb7  :  255 - 0xff
    "11111111", -- 7352 - 0x1cb8  :  255 - 0xff
    "11111111", -- 7353 - 0x1cb9  :  255 - 0xff
    "11111111", -- 7354 - 0x1cba  :  255 - 0xff
    "11111000", -- 7355 - 0x1cbb  :  248 - 0xf8
    "11111110", -- 7356 - 0x1cbc  :  254 - 0xfe
    "11111111", -- 7357 - 0x1cbd  :  255 - 0xff
    "11111111", -- 7358 - 0x1cbe  :  255 - 0xff
    "11111111", -- 7359 - 0x1cbf  :  255 - 0xff
    "11111111", -- 7360 - 0x1cc0  :  255 - 0xff -- Background 0xcc
    "11111111", -- 7361 - 0x1cc1  :  255 - 0xff
    "11111111", -- 7362 - 0x1cc2  :  255 - 0xff
    "00111111", -- 7363 - 0x1cc3  :   63 - 0x3f
    "00011110", -- 7364 - 0x1cc4  :   30 - 0x1e
    "00000001", -- 7365 - 0x1cc5  :    1 - 0x1
    "00000000", -- 7366 - 0x1cc6  :    0 - 0x0
    "00000000", -- 7367 - 0x1cc7  :    0 - 0x0
    "11111111", -- 7368 - 0x1cc8  :  255 - 0xff
    "11111111", -- 7369 - 0x1cc9  :  255 - 0xff
    "11111111", -- 7370 - 0x1cca  :  255 - 0xff
    "00111111", -- 7371 - 0x1ccb  :   63 - 0x3f
    "00011111", -- 7372 - 0x1ccc  :   31 - 0x1f
    "00011111", -- 7373 - 0x1ccd  :   31 - 0x1f
    "00000000", -- 7374 - 0x1cce  :    0 - 0x0
    "00000000", -- 7375 - 0x1ccf  :    0 - 0x0
    "00000000", -- 7376 - 0x1cd0  :    0 - 0x0 -- Background 0xcd
    "00000000", -- 7377 - 0x1cd1  :    0 - 0x0
    "00000000", -- 7378 - 0x1cd2  :    0 - 0x0
    "10000000", -- 7379 - 0x1cd3  :  128 - 0x80
    "11000000", -- 7380 - 0x1cd4  :  192 - 0xc0
    "11100000", -- 7381 - 0x1cd5  :  224 - 0xe0
    "11100000", -- 7382 - 0x1cd6  :  224 - 0xe0
    "11100000", -- 7383 - 0x1cd7  :  224 - 0xe0
    "00000000", -- 7384 - 0x1cd8  :    0 - 0x0
    "00000000", -- 7385 - 0x1cd9  :    0 - 0x0
    "10000000", -- 7386 - 0x1cda  :  128 - 0x80
    "11000000", -- 7387 - 0x1cdb  :  192 - 0xc0
    "11100000", -- 7388 - 0x1cdc  :  224 - 0xe0
    "11100000", -- 7389 - 0x1cdd  :  224 - 0xe0
    "11100000", -- 7390 - 0x1cde  :  224 - 0xe0
    "11100000", -- 7391 - 0x1cdf  :  224 - 0xe0
    "11000000", -- 7392 - 0x1ce0  :  192 - 0xc0 -- Background 0xce
    "10000000", -- 7393 - 0x1ce1  :  128 - 0x80
    "00000000", -- 7394 - 0x1ce2  :    0 - 0x0
    "00000000", -- 7395 - 0x1ce3  :    0 - 0x0
    "00000000", -- 7396 - 0x1ce4  :    0 - 0x0
    "00000000", -- 7397 - 0x1ce5  :    0 - 0x0
    "10000000", -- 7398 - 0x1ce6  :  128 - 0x80
    "10000000", -- 7399 - 0x1ce7  :  128 - 0x80
    "11000000", -- 7400 - 0x1ce8  :  192 - 0xc0
    "10000000", -- 7401 - 0x1ce9  :  128 - 0x80
    "00000000", -- 7402 - 0x1cea  :    0 - 0x0
    "00000000", -- 7403 - 0x1ceb  :    0 - 0x0
    "00000000", -- 7404 - 0x1cec  :    0 - 0x0
    "10000000", -- 7405 - 0x1ced  :  128 - 0x80
    "11000000", -- 7406 - 0x1cee  :  192 - 0xc0
    "11000000", -- 7407 - 0x1cef  :  192 - 0xc0
    "10000000", -- 7408 - 0x1cf0  :  128 - 0x80 -- Background 0xcf
    "10000000", -- 7409 - 0x1cf1  :  128 - 0x80
    "11100000", -- 7410 - 0x1cf2  :  224 - 0xe0
    "11000000", -- 7411 - 0x1cf3  :  192 - 0xc0
    "00100000", -- 7412 - 0x1cf4  :   32 - 0x20
    "00000000", -- 7413 - 0x1cf5  :    0 - 0x0
    "00000000", -- 7414 - 0x1cf6  :    0 - 0x0
    "00000000", -- 7415 - 0x1cf7  :    0 - 0x0
    "11000000", -- 7416 - 0x1cf8  :  192 - 0xc0
    "11000000", -- 7417 - 0x1cf9  :  192 - 0xc0
    "11100000", -- 7418 - 0x1cfa  :  224 - 0xe0
    "11111000", -- 7419 - 0x1cfb  :  248 - 0xf8
    "11111100", -- 7420 - 0x1cfc  :  252 - 0xfc
    "11111100", -- 7421 - 0x1cfd  :  252 - 0xfc
    "00000000", -- 7422 - 0x1cfe  :    0 - 0x0
    "00000000", -- 7423 - 0x1cff  :    0 - 0x0
    "00011111", -- 7424 - 0x1d00  :   31 - 0x1f -- Background 0xd0
    "00000110", -- 7425 - 0x1d01  :    6 - 0x6
    "00000110", -- 7426 - 0x1d02  :    6 - 0x6
    "00000110", -- 7427 - 0x1d03  :    6 - 0x6
    "00000110", -- 7428 - 0x1d04  :    6 - 0x6
    "00000110", -- 7429 - 0x1d05  :    6 - 0x6
    "00000110", -- 7430 - 0x1d06  :    6 - 0x6
    "00000000", -- 7431 - 0x1d07  :    0 - 0x0
    "00000000", -- 7432 - 0x1d08  :    0 - 0x0
    "00000000", -- 7433 - 0x1d09  :    0 - 0x0
    "00000000", -- 7434 - 0x1d0a  :    0 - 0x0
    "00000000", -- 7435 - 0x1d0b  :    0 - 0x0
    "00000000", -- 7436 - 0x1d0c  :    0 - 0x0
    "00000000", -- 7437 - 0x1d0d  :    0 - 0x0
    "00000000", -- 7438 - 0x1d0e  :    0 - 0x0
    "00000000", -- 7439 - 0x1d0f  :    0 - 0x0
    "00111001", -- 7440 - 0x1d10  :   57 - 0x39 -- Background 0xd1
    "01100101", -- 7441 - 0x1d11  :  101 - 0x65
    "01100101", -- 7442 - 0x1d12  :  101 - 0x65
    "01100101", -- 7443 - 0x1d13  :  101 - 0x65
    "01100101", -- 7444 - 0x1d14  :  101 - 0x65
    "01100101", -- 7445 - 0x1d15  :  101 - 0x65
    "00111001", -- 7446 - 0x1d16  :   57 - 0x39
    "00000000", -- 7447 - 0x1d17  :    0 - 0x0
    "00000000", -- 7448 - 0x1d18  :    0 - 0x0
    "00000000", -- 7449 - 0x1d19  :    0 - 0x0
    "00000000", -- 7450 - 0x1d1a  :    0 - 0x0
    "00000000", -- 7451 - 0x1d1b  :    0 - 0x0
    "00000000", -- 7452 - 0x1d1c  :    0 - 0x0
    "00000000", -- 7453 - 0x1d1d  :    0 - 0x0
    "00000000", -- 7454 - 0x1d1e  :    0 - 0x0
    "00000000", -- 7455 - 0x1d1f  :    0 - 0x0
    "11100000", -- 7456 - 0x1d20  :  224 - 0xe0 -- Background 0xd2
    "10110000", -- 7457 - 0x1d21  :  176 - 0xb0
    "10110000", -- 7458 - 0x1d22  :  176 - 0xb0
    "10110110", -- 7459 - 0x1d23  :  182 - 0xb6
    "11100110", -- 7460 - 0x1d24  :  230 - 0xe6
    "10000000", -- 7461 - 0x1d25  :  128 - 0x80
    "10000000", -- 7462 - 0x1d26  :  128 - 0x80
    "00000000", -- 7463 - 0x1d27  :    0 - 0x0
    "00000000", -- 7464 - 0x1d28  :    0 - 0x0
    "00000000", -- 7465 - 0x1d29  :    0 - 0x0
    "00000000", -- 7466 - 0x1d2a  :    0 - 0x0
    "00000000", -- 7467 - 0x1d2b  :    0 - 0x0
    "00000000", -- 7468 - 0x1d2c  :    0 - 0x0
    "00000000", -- 7469 - 0x1d2d  :    0 - 0x0
    "00000000", -- 7470 - 0x1d2e  :    0 - 0x0
    "00000000", -- 7471 - 0x1d2f  :    0 - 0x0
    "00111100", -- 7472 - 0x1d30  :   60 - 0x3c -- Background 0xd3
    "01000010", -- 7473 - 0x1d31  :   66 - 0x42
    "10011001", -- 7474 - 0x1d32  :  153 - 0x99
    "10100001", -- 7475 - 0x1d33  :  161 - 0xa1
    "10100001", -- 7476 - 0x1d34  :  161 - 0xa1
    "10011001", -- 7477 - 0x1d35  :  153 - 0x99
    "01000010", -- 7478 - 0x1d36  :   66 - 0x42
    "00111100", -- 7479 - 0x1d37  :   60 - 0x3c
    "00000000", -- 7480 - 0x1d38  :    0 - 0x0
    "00000000", -- 7481 - 0x1d39  :    0 - 0x0
    "00000000", -- 7482 - 0x1d3a  :    0 - 0x0
    "00000000", -- 7483 - 0x1d3b  :    0 - 0x0
    "00000000", -- 7484 - 0x1d3c  :    0 - 0x0
    "00000000", -- 7485 - 0x1d3d  :    0 - 0x0
    "00000000", -- 7486 - 0x1d3e  :    0 - 0x0
    "00000000", -- 7487 - 0x1d3f  :    0 - 0x0
    "00000000", -- 7488 - 0x1d40  :    0 - 0x0 -- Background 0xd4
    "00000000", -- 7489 - 0x1d41  :    0 - 0x0
    "00000000", -- 7490 - 0x1d42  :    0 - 0x0
    "00000011", -- 7491 - 0x1d43  :    3 - 0x3
    "00000110", -- 7492 - 0x1d44  :    6 - 0x6
    "00000000", -- 7493 - 0x1d45  :    0 - 0x0
    "00000001", -- 7494 - 0x1d46  :    1 - 0x1
    "00000111", -- 7495 - 0x1d47  :    7 - 0x7
    "00000000", -- 7496 - 0x1d48  :    0 - 0x0
    "00000000", -- 7497 - 0x1d49  :    0 - 0x0
    "00000000", -- 7498 - 0x1d4a  :    0 - 0x0
    "00000000", -- 7499 - 0x1d4b  :    0 - 0x0
    "00000011", -- 7500 - 0x1d4c  :    3 - 0x3
    "00000111", -- 7501 - 0x1d4d  :    7 - 0x7
    "00000011", -- 7502 - 0x1d4e  :    3 - 0x3
    "00000111", -- 7503 - 0x1d4f  :    7 - 0x7
    "00001111", -- 7504 - 0x1d50  :   15 - 0xf -- Background 0xd5
    "00011111", -- 7505 - 0x1d51  :   31 - 0x1f
    "00111111", -- 7506 - 0x1d52  :   63 - 0x3f
    "01111111", -- 7507 - 0x1d53  :  127 - 0x7f
    "01111111", -- 7508 - 0x1d54  :  127 - 0x7f
    "01111111", -- 7509 - 0x1d55  :  127 - 0x7f
    "11111111", -- 7510 - 0x1d56  :  255 - 0xff
    "01111111", -- 7511 - 0x1d57  :  127 - 0x7f
    "00011111", -- 7512 - 0x1d58  :   31 - 0x1f
    "00111111", -- 7513 - 0x1d59  :   63 - 0x3f
    "01111111", -- 7514 - 0x1d5a  :  127 - 0x7f
    "11111111", -- 7515 - 0x1d5b  :  255 - 0xff
    "11111111", -- 7516 - 0x1d5c  :  255 - 0xff
    "11111111", -- 7517 - 0x1d5d  :  255 - 0xff
    "11111111", -- 7518 - 0x1d5e  :  255 - 0xff
    "01111111", -- 7519 - 0x1d5f  :  127 - 0x7f
    "00000000", -- 7520 - 0x1d60  :    0 - 0x0 -- Background 0xd6
    "00000000", -- 7521 - 0x1d61  :    0 - 0x0
    "00000000", -- 7522 - 0x1d62  :    0 - 0x0
    "10000000", -- 7523 - 0x1d63  :  128 - 0x80
    "00000000", -- 7524 - 0x1d64  :    0 - 0x0
    "00000000", -- 7525 - 0x1d65  :    0 - 0x0
    "00000000", -- 7526 - 0x1d66  :    0 - 0x0
    "10100000", -- 7527 - 0x1d67  :  160 - 0xa0
    "00000000", -- 7528 - 0x1d68  :    0 - 0x0
    "00000000", -- 7529 - 0x1d69  :    0 - 0x0
    "00000000", -- 7530 - 0x1d6a  :    0 - 0x0
    "11000000", -- 7531 - 0x1d6b  :  192 - 0xc0
    "11100000", -- 7532 - 0x1d6c  :  224 - 0xe0
    "11110000", -- 7533 - 0x1d6d  :  240 - 0xf0
    "11110000", -- 7534 - 0x1d6e  :  240 - 0xf0
    "11111000", -- 7535 - 0x1d6f  :  248 - 0xf8
    "11100000", -- 7536 - 0x1d70  :  224 - 0xe0 -- Background 0xd7
    "11110000", -- 7537 - 0x1d71  :  240 - 0xf0
    "11100000", -- 7538 - 0x1d72  :  224 - 0xe0
    "11011101", -- 7539 - 0x1d73  :  221 - 0xdd
    "11111010", -- 7540 - 0x1d74  :  250 - 0xfa
    "11101011", -- 7541 - 0x1d75  :  235 - 0xeb
    "10000000", -- 7542 - 0x1d76  :  128 - 0x80
    "00000000", -- 7543 - 0x1d77  :    0 - 0x0
    "11111100", -- 7544 - 0x1d78  :  252 - 0xfc
    "11111000", -- 7545 - 0x1d79  :  248 - 0xf8
    "11110000", -- 7546 - 0x1d7a  :  240 - 0xf0
    "11111111", -- 7547 - 0x1d7b  :  255 - 0xff
    "11111111", -- 7548 - 0x1d7c  :  255 - 0xff
    "11111111", -- 7549 - 0x1d7d  :  255 - 0xff
    "11111111", -- 7550 - 0x1d7e  :  255 - 0xff
    "11111111", -- 7551 - 0x1d7f  :  255 - 0xff
    "00000000", -- 7552 - 0x1d80  :    0 - 0x0 -- Background 0xd8
    "00000000", -- 7553 - 0x1d81  :    0 - 0x0
    "00000000", -- 7554 - 0x1d82  :    0 - 0x0
    "00000011", -- 7555 - 0x1d83  :    3 - 0x3
    "00000110", -- 7556 - 0x1d84  :    6 - 0x6
    "00000000", -- 7557 - 0x1d85  :    0 - 0x0
    "00000001", -- 7558 - 0x1d86  :    1 - 0x1
    "00000001", -- 7559 - 0x1d87  :    1 - 0x1
    "00000000", -- 7560 - 0x1d88  :    0 - 0x0
    "00000000", -- 7561 - 0x1d89  :    0 - 0x0
    "00000000", -- 7562 - 0x1d8a  :    0 - 0x0
    "00000000", -- 7563 - 0x1d8b  :    0 - 0x0
    "00000011", -- 7564 - 0x1d8c  :    3 - 0x3
    "00000111", -- 7565 - 0x1d8d  :    7 - 0x7
    "00001111", -- 7566 - 0x1d8e  :   15 - 0xf
    "00011111", -- 7567 - 0x1d8f  :   31 - 0x1f
    "00001011", -- 7568 - 0x1d90  :   11 - 0xb -- Background 0xd9
    "00000111", -- 7569 - 0x1d91  :    7 - 0x7
    "00000011", -- 7570 - 0x1d92  :    3 - 0x3
    "01011101", -- 7571 - 0x1d93  :   93 - 0x5d
    "10101111", -- 7572 - 0x1d94  :  175 - 0xaf
    "01010011", -- 7573 - 0x1d95  :   83 - 0x53
    "00000000", -- 7574 - 0x1d96  :    0 - 0x0
    "00000000", -- 7575 - 0x1d97  :    0 - 0x0
    "00111111", -- 7576 - 0x1d98  :   63 - 0x3f
    "00011111", -- 7577 - 0x1d99  :   31 - 0x1f
    "00000111", -- 7578 - 0x1d9a  :    7 - 0x7
    "11111111", -- 7579 - 0x1d9b  :  255 - 0xff
    "11111111", -- 7580 - 0x1d9c  :  255 - 0xff
    "11111111", -- 7581 - 0x1d9d  :  255 - 0xff
    "11111111", -- 7582 - 0x1d9e  :  255 - 0xff
    "11111111", -- 7583 - 0x1d9f  :  255 - 0xff
    "00000000", -- 7584 - 0x1da0  :    0 - 0x0 -- Background 0xda
    "00000000", -- 7585 - 0x1da1  :    0 - 0x0
    "00000000", -- 7586 - 0x1da2  :    0 - 0x0
    "10000000", -- 7587 - 0x1da3  :  128 - 0x80
    "00000000", -- 7588 - 0x1da4  :    0 - 0x0
    "00000000", -- 7589 - 0x1da5  :    0 - 0x0
    "01100000", -- 7590 - 0x1da6  :   96 - 0x60
    "11110000", -- 7591 - 0x1da7  :  240 - 0xf0
    "00000000", -- 7592 - 0x1da8  :    0 - 0x0
    "00000000", -- 7593 - 0x1da9  :    0 - 0x0
    "00000000", -- 7594 - 0x1daa  :    0 - 0x0
    "11000000", -- 7595 - 0x1dab  :  192 - 0xc0
    "11000000", -- 7596 - 0x1dac  :  192 - 0xc0
    "11000000", -- 7597 - 0x1dad  :  192 - 0xc0
    "11100000", -- 7598 - 0x1dae  :  224 - 0xe0
    "11111000", -- 7599 - 0x1daf  :  248 - 0xf8
    "11111000", -- 7600 - 0x1db0  :  248 - 0xf8 -- Background 0xdb
    "11111100", -- 7601 - 0x1db1  :  252 - 0xfc
    "11111100", -- 7602 - 0x1db2  :  252 - 0xfc
    "11111110", -- 7603 - 0x1db3  :  254 - 0xfe
    "11111110", -- 7604 - 0x1db4  :  254 - 0xfe
    "11111111", -- 7605 - 0x1db5  :  255 - 0xff
    "11111111", -- 7606 - 0x1db6  :  255 - 0xff
    "01111110", -- 7607 - 0x1db7  :  126 - 0x7e
    "11111100", -- 7608 - 0x1db8  :  252 - 0xfc
    "11111110", -- 7609 - 0x1db9  :  254 - 0xfe
    "11111110", -- 7610 - 0x1dba  :  254 - 0xfe
    "11111111", -- 7611 - 0x1dbb  :  255 - 0xff
    "11111111", -- 7612 - 0x1dbc  :  255 - 0xff
    "11111111", -- 7613 - 0x1dbd  :  255 - 0xff
    "11111111", -- 7614 - 0x1dbe  :  255 - 0xff
    "11111110", -- 7615 - 0x1dbf  :  254 - 0xfe
    "00000000", -- 7616 - 0x1dc0  :    0 - 0x0 -- Background 0xdc
    "00000000", -- 7617 - 0x1dc1  :    0 - 0x0
    "00000000", -- 7618 - 0x1dc2  :    0 - 0x0
    "00000000", -- 7619 - 0x1dc3  :    0 - 0x0
    "00000000", -- 7620 - 0x1dc4  :    0 - 0x0
    "00000000", -- 7621 - 0x1dc5  :    0 - 0x0
    "00100001", -- 7622 - 0x1dc6  :   33 - 0x21
    "00111111", -- 7623 - 0x1dc7  :   63 - 0x3f
    "00110110", -- 7624 - 0x1dc8  :   54 - 0x36
    "00110110", -- 7625 - 0x1dc9  :   54 - 0x36
    "01111110", -- 7626 - 0x1dca  :  126 - 0x7e
    "01111111", -- 7627 - 0x1dcb  :  127 - 0x7f
    "01111111", -- 7628 - 0x1dcc  :  127 - 0x7f
    "01111111", -- 7629 - 0x1dcd  :  127 - 0x7f
    "00111111", -- 7630 - 0x1dce  :   63 - 0x3f
    "00111111", -- 7631 - 0x1dcf  :   63 - 0x3f
    "00111111", -- 7632 - 0x1dd0  :   63 - 0x3f -- Background 0xdd
    "00011111", -- 7633 - 0x1dd1  :   31 - 0x1f
    "00011111", -- 7634 - 0x1dd2  :   31 - 0x1f
    "00001111", -- 7635 - 0x1dd3  :   15 - 0xf
    "00000111", -- 7636 - 0x1dd4  :    7 - 0x7
    "00000011", -- 7637 - 0x1dd5  :    3 - 0x3
    "00000000", -- 7638 - 0x1dd6  :    0 - 0x0
    "00000000", -- 7639 - 0x1dd7  :    0 - 0x0
    "00111111", -- 7640 - 0x1dd8  :   63 - 0x3f
    "00011111", -- 7641 - 0x1dd9  :   31 - 0x1f
    "00011111", -- 7642 - 0x1dda  :   31 - 0x1f
    "00001111", -- 7643 - 0x1ddb  :   15 - 0xf
    "00000111", -- 7644 - 0x1ddc  :    7 - 0x7
    "00000011", -- 7645 - 0x1ddd  :    3 - 0x3
    "00000000", -- 7646 - 0x1dde  :    0 - 0x0
    "00000000", -- 7647 - 0x1ddf  :    0 - 0x0
    "00111110", -- 7648 - 0x1de0  :   62 - 0x3e -- Background 0xde
    "00011110", -- 7649 - 0x1de1  :   30 - 0x1e
    "00011110", -- 7650 - 0x1de2  :   30 - 0x1e
    "00001110", -- 7651 - 0x1de3  :   14 - 0xe
    "00001111", -- 7652 - 0x1de4  :   15 - 0xf
    "00011111", -- 7653 - 0x1de5  :   31 - 0x1f
    "10011111", -- 7654 - 0x1de6  :  159 - 0x9f
    "10011111", -- 7655 - 0x1de7  :  159 - 0x9f
    "00111111", -- 7656 - 0x1de8  :   63 - 0x3f
    "00011111", -- 7657 - 0x1de9  :   31 - 0x1f
    "11011111", -- 7658 - 0x1dea  :  223 - 0xdf
    "11001111", -- 7659 - 0x1deb  :  207 - 0xcf
    "11001111", -- 7660 - 0x1dec  :  207 - 0xcf
    "10011111", -- 7661 - 0x1ded  :  159 - 0x9f
    "11011111", -- 7662 - 0x1dee  :  223 - 0xdf
    "11111111", -- 7663 - 0x1def  :  255 - 0xff
    "11011111", -- 7664 - 0x1df0  :  223 - 0xdf -- Background 0xdf
    "11111111", -- 7665 - 0x1df1  :  255 - 0xff
    "11111111", -- 7666 - 0x1df2  :  255 - 0xff
    "11111111", -- 7667 - 0x1df3  :  255 - 0xff
    "11111111", -- 7668 - 0x1df4  :  255 - 0xff
    "11011111", -- 7669 - 0x1df5  :  223 - 0xdf
    "11100111", -- 7670 - 0x1df6  :  231 - 0xe7
    "00000000", -- 7671 - 0x1df7  :    0 - 0x0
    "11111111", -- 7672 - 0x1df8  :  255 - 0xff
    "11111111", -- 7673 - 0x1df9  :  255 - 0xff
    "11111111", -- 7674 - 0x1dfa  :  255 - 0xff
    "11111111", -- 7675 - 0x1dfb  :  255 - 0xff
    "11111111", -- 7676 - 0x1dfc  :  255 - 0xff
    "11111111", -- 7677 - 0x1dfd  :  255 - 0xff
    "11111111", -- 7678 - 0x1dfe  :  255 - 0xff
    "00001111", -- 7679 - 0x1dff  :   15 - 0xf
    "00100000", -- 7680 - 0x1e00  :   32 - 0x20 -- Background 0xe0
    "00001111", -- 7681 - 0x1e01  :   15 - 0xf
    "00110000", -- 7682 - 0x1e02  :   48 - 0x30
    "01000000", -- 7683 - 0x1e03  :   64 - 0x40
    "10011000", -- 7684 - 0x1e04  :  152 - 0x98
    "00111110", -- 7685 - 0x1e05  :   62 - 0x3e
    "00011111", -- 7686 - 0x1e06  :   31 - 0x1f
    "00000000", -- 7687 - 0x1e07  :    0 - 0x0
    "11111111", -- 7688 - 0x1e08  :  255 - 0xff
    "11111111", -- 7689 - 0x1e09  :  255 - 0xff
    "11111111", -- 7690 - 0x1e0a  :  255 - 0xff
    "11111111", -- 7691 - 0x1e0b  :  255 - 0xff
    "11111111", -- 7692 - 0x1e0c  :  255 - 0xff
    "11111111", -- 7693 - 0x1e0d  :  255 - 0xff
    "11111111", -- 7694 - 0x1e0e  :  255 - 0xff
    "11111111", -- 7695 - 0x1e0f  :  255 - 0xff
    "10000001", -- 7696 - 0x1e10  :  129 - 0x81 -- Background 0xe1
    "00110110", -- 7697 - 0x1e11  :   54 - 0x36
    "00101110", -- 7698 - 0x1e12  :   46 - 0x2e
    "10101111", -- 7699 - 0x1e13  :  175 - 0xaf
    "10101110", -- 7700 - 0x1e14  :  174 - 0xae
    "11010001", -- 7701 - 0x1e15  :  209 - 0xd1
    "11101111", -- 7702 - 0x1e16  :  239 - 0xef
    "10000111", -- 7703 - 0x1e17  :  135 - 0x87
    "11111111", -- 7704 - 0x1e18  :  255 - 0xff
    "11111001", -- 7705 - 0x1e19  :  249 - 0xf9
    "11110000", -- 7706 - 0x1e1a  :  240 - 0xf0
    "11110000", -- 7707 - 0x1e1b  :  240 - 0xf0
    "10110001", -- 7708 - 0x1e1c  :  177 - 0xb1
    "11011111", -- 7709 - 0x1e1d  :  223 - 0xdf
    "11101111", -- 7710 - 0x1e1e  :  239 - 0xef
    "10000111", -- 7711 - 0x1e1f  :  135 - 0x87
    "00000010", -- 7712 - 0x1e20  :    2 - 0x2 -- Background 0xe2
    "11111000", -- 7713 - 0x1e21  :  248 - 0xf8
    "00000110", -- 7714 - 0x1e22  :    6 - 0x6
    "00000001", -- 7715 - 0x1e23  :    1 - 0x1
    "00001100", -- 7716 - 0x1e24  :   12 - 0xc
    "00111110", -- 7717 - 0x1e25  :   62 - 0x3e
    "11111100", -- 7718 - 0x1e26  :  252 - 0xfc
    "00000000", -- 7719 - 0x1e27  :    0 - 0x0
    "11111111", -- 7720 - 0x1e28  :  255 - 0xff
    "11111111", -- 7721 - 0x1e29  :  255 - 0xff
    "11111111", -- 7722 - 0x1e2a  :  255 - 0xff
    "11111111", -- 7723 - 0x1e2b  :  255 - 0xff
    "11111111", -- 7724 - 0x1e2c  :  255 - 0xff
    "11111111", -- 7725 - 0x1e2d  :  255 - 0xff
    "11111111", -- 7726 - 0x1e2e  :  255 - 0xff
    "11111111", -- 7727 - 0x1e2f  :  255 - 0xff
    "11000000", -- 7728 - 0x1e30  :  192 - 0xc0 -- Background 0xe3
    "00110110", -- 7729 - 0x1e31  :   54 - 0x36
    "00111110", -- 7730 - 0x1e32  :   62 - 0x3e
    "01111010", -- 7731 - 0x1e33  :  122 - 0x7a
    "10110110", -- 7732 - 0x1e34  :  182 - 0xb6
    "11001101", -- 7733 - 0x1e35  :  205 - 0xcd
    "11111011", -- 7734 - 0x1e36  :  251 - 0xfb
    "11110000", -- 7735 - 0x1e37  :  240 - 0xf0
    "11111111", -- 7736 - 0x1e38  :  255 - 0xff
    "11001111", -- 7737 - 0x1e39  :  207 - 0xcf
    "10000111", -- 7738 - 0x1e3a  :  135 - 0x87
    "10000111", -- 7739 - 0x1e3b  :  135 - 0x87
    "11001110", -- 7740 - 0x1e3c  :  206 - 0xce
    "11111101", -- 7741 - 0x1e3d  :  253 - 0xfd
    "11111011", -- 7742 - 0x1e3e  :  251 - 0xfb
    "11110000", -- 7743 - 0x1e3f  :  240 - 0xf0
    "00111110", -- 7744 - 0x1e40  :   62 - 0x3e -- Background 0xe4
    "00111100", -- 7745 - 0x1e41  :   60 - 0x3c
    "00111100", -- 7746 - 0x1e42  :   60 - 0x3c
    "00111000", -- 7747 - 0x1e43  :   56 - 0x38
    "11111000", -- 7748 - 0x1e44  :  248 - 0xf8
    "01111100", -- 7749 - 0x1e45  :  124 - 0x7c
    "01111110", -- 7750 - 0x1e46  :  126 - 0x7e
    "01111000", -- 7751 - 0x1e47  :  120 - 0x78
    "11111110", -- 7752 - 0x1e48  :  254 - 0xfe
    "11111100", -- 7753 - 0x1e49  :  252 - 0xfc
    "11111100", -- 7754 - 0x1e4a  :  252 - 0xfc
    "11111000", -- 7755 - 0x1e4b  :  248 - 0xf8
    "11111011", -- 7756 - 0x1e4c  :  251 - 0xfb
    "11111101", -- 7757 - 0x1e4d  :  253 - 0xfd
    "11111110", -- 7758 - 0x1e4e  :  254 - 0xfe
    "11111111", -- 7759 - 0x1e4f  :  255 - 0xff
    "11111000", -- 7760 - 0x1e50  :  248 - 0xf8 -- Background 0xe5
    "01111111", -- 7761 - 0x1e51  :  127 - 0x7f
    "01111111", -- 7762 - 0x1e52  :  127 - 0x7f
    "11111110", -- 7763 - 0x1e53  :  254 - 0xfe
    "11111111", -- 7764 - 0x1e54  :  255 - 0xff
    "11111111", -- 7765 - 0x1e55  :  255 - 0xff
    "11110011", -- 7766 - 0x1e56  :  243 - 0xf3
    "10000001", -- 7767 - 0x1e57  :  129 - 0x81
    "11111111", -- 7768 - 0x1e58  :  255 - 0xff
    "11111111", -- 7769 - 0x1e59  :  255 - 0xff
    "11111111", -- 7770 - 0x1e5a  :  255 - 0xff
    "11111111", -- 7771 - 0x1e5b  :  255 - 0xff
    "11111111", -- 7772 - 0x1e5c  :  255 - 0xff
    "11111111", -- 7773 - 0x1e5d  :  255 - 0xff
    "11111111", -- 7774 - 0x1e5e  :  255 - 0xff
    "11111001", -- 7775 - 0x1e5f  :  249 - 0xf9
    "00000000", -- 7776 - 0x1e60  :    0 - 0x0 -- Background 0xe6
    "00000000", -- 7777 - 0x1e61  :    0 - 0x0
    "00000000", -- 7778 - 0x1e62  :    0 - 0x0
    "00010000", -- 7779 - 0x1e63  :   16 - 0x10
    "01000000", -- 7780 - 0x1e64  :   64 - 0x40
    "00100000", -- 7781 - 0x1e65  :   32 - 0x20
    "00000000", -- 7782 - 0x1e66  :    0 - 0x0
    "00000000", -- 7783 - 0x1e67  :    0 - 0x0
    "00000000", -- 7784 - 0x1e68  :    0 - 0x0
    "00000000", -- 7785 - 0x1e69  :    0 - 0x0
    "00000000", -- 7786 - 0x1e6a  :    0 - 0x0
    "01111000", -- 7787 - 0x1e6b  :  120 - 0x78
    "11111100", -- 7788 - 0x1e6c  :  252 - 0xfc
    "11111100", -- 7789 - 0x1e6d  :  252 - 0xfc
    "11111100", -- 7790 - 0x1e6e  :  252 - 0xfc
    "11111100", -- 7791 - 0x1e6f  :  252 - 0xfc
    "00000110", -- 7792 - 0x1e70  :    6 - 0x6 -- Background 0xe7
    "00001110", -- 7793 - 0x1e71  :   14 - 0xe
    "01111110", -- 7794 - 0x1e72  :  126 - 0x7e
    "11111110", -- 7795 - 0x1e73  :  254 - 0xfe
    "11111110", -- 7796 - 0x1e74  :  254 - 0xfe
    "11111100", -- 7797 - 0x1e75  :  252 - 0xfc
    "11111000", -- 7798 - 0x1e76  :  248 - 0xf8
    "11110000", -- 7799 - 0x1e77  :  240 - 0xf0
    "11111110", -- 7800 - 0x1e78  :  254 - 0xfe
    "11111110", -- 7801 - 0x1e79  :  254 - 0xfe
    "11111110", -- 7802 - 0x1e7a  :  254 - 0xfe
    "11111110", -- 7803 - 0x1e7b  :  254 - 0xfe
    "11111110", -- 7804 - 0x1e7c  :  254 - 0xfe
    "11111100", -- 7805 - 0x1e7d  :  252 - 0xfc
    "11111000", -- 7806 - 0x1e7e  :  248 - 0xf8
    "11110000", -- 7807 - 0x1e7f  :  240 - 0xf0
    "00000000", -- 7808 - 0x1e80  :    0 - 0x0 -- Background 0xe8
    "00000000", -- 7809 - 0x1e81  :    0 - 0x0
    "00000000", -- 7810 - 0x1e82  :    0 - 0x0
    "00000000", -- 7811 - 0x1e83  :    0 - 0x0
    "00000000", -- 7812 - 0x1e84  :    0 - 0x0
    "00000000", -- 7813 - 0x1e85  :    0 - 0x0
    "00000000", -- 7814 - 0x1e86  :    0 - 0x0
    "00000001", -- 7815 - 0x1e87  :    1 - 0x1
    "00000000", -- 7816 - 0x1e88  :    0 - 0x0
    "00000000", -- 7817 - 0x1e89  :    0 - 0x0
    "00000000", -- 7818 - 0x1e8a  :    0 - 0x0
    "00000000", -- 7819 - 0x1e8b  :    0 - 0x0
    "00000000", -- 7820 - 0x1e8c  :    0 - 0x0
    "00000000", -- 7821 - 0x1e8d  :    0 - 0x0
    "00000000", -- 7822 - 0x1e8e  :    0 - 0x0
    "00000000", -- 7823 - 0x1e8f  :    0 - 0x0
    "00000010", -- 7824 - 0x1e90  :    2 - 0x2 -- Background 0xe9
    "00000000", -- 7825 - 0x1e91  :    0 - 0x0
    "00001000", -- 7826 - 0x1e92  :    8 - 0x8
    "00000001", -- 7827 - 0x1e93  :    1 - 0x1
    "00010011", -- 7828 - 0x1e94  :   19 - 0x13
    "00000001", -- 7829 - 0x1e95  :    1 - 0x1
    "00000000", -- 7830 - 0x1e96  :    0 - 0x0
    "00000000", -- 7831 - 0x1e97  :    0 - 0x0
    "00000001", -- 7832 - 0x1e98  :    1 - 0x1
    "00001111", -- 7833 - 0x1e99  :   15 - 0xf
    "00011111", -- 7834 - 0x1e9a  :   31 - 0x1f
    "00011111", -- 7835 - 0x1e9b  :   31 - 0x1f
    "00111011", -- 7836 - 0x1e9c  :   59 - 0x3b
    "00110011", -- 7837 - 0x1e9d  :   51 - 0x33
    "00000001", -- 7838 - 0x1e9e  :    1 - 0x1
    "00000001", -- 7839 - 0x1e9f  :    1 - 0x1
    "00000000", -- 7840 - 0x1ea0  :    0 - 0x0 -- Background 0xea
    "00000000", -- 7841 - 0x1ea1  :    0 - 0x0
    "00000000", -- 7842 - 0x1ea2  :    0 - 0x0
    "00000000", -- 7843 - 0x1ea3  :    0 - 0x0
    "00000000", -- 7844 - 0x1ea4  :    0 - 0x0
    "00000000", -- 7845 - 0x1ea5  :    0 - 0x0
    "00000000", -- 7846 - 0x1ea6  :    0 - 0x0
    "00000000", -- 7847 - 0x1ea7  :    0 - 0x0
    "00000000", -- 7848 - 0x1ea8  :    0 - 0x0
    "00000000", -- 7849 - 0x1ea9  :    0 - 0x0
    "00000000", -- 7850 - 0x1eaa  :    0 - 0x0
    "00110110", -- 7851 - 0x1eab  :   54 - 0x36
    "01101100", -- 7852 - 0x1eac  :  108 - 0x6c
    "11111101", -- 7853 - 0x1ead  :  253 - 0xfd
    "11111111", -- 7854 - 0x1eae  :  255 - 0xff
    "11111111", -- 7855 - 0x1eaf  :  255 - 0xff
    "00000000", -- 7856 - 0x1eb0  :    0 - 0x0 -- Background 0xeb
    "01000011", -- 7857 - 0x1eb1  :   67 - 0x43
    "01111111", -- 7858 - 0x1eb2  :  127 - 0x7f
    "01111111", -- 7859 - 0x1eb3  :  127 - 0x7f
    "01111111", -- 7860 - 0x1eb4  :  127 - 0x7f
    "00111111", -- 7861 - 0x1eb5  :   63 - 0x3f
    "00011111", -- 7862 - 0x1eb6  :   31 - 0x1f
    "00000111", -- 7863 - 0x1eb7  :    7 - 0x7
    "11111111", -- 7864 - 0x1eb8  :  255 - 0xff
    "01111111", -- 7865 - 0x1eb9  :  127 - 0x7f
    "01111111", -- 7866 - 0x1eba  :  127 - 0x7f
    "01111111", -- 7867 - 0x1ebb  :  127 - 0x7f
    "01111111", -- 7868 - 0x1ebc  :  127 - 0x7f
    "00111111", -- 7869 - 0x1ebd  :   63 - 0x3f
    "00011111", -- 7870 - 0x1ebe  :   31 - 0x1f
    "00000111", -- 7871 - 0x1ebf  :    7 - 0x7
    "00000000", -- 7872 - 0x1ec0  :    0 - 0x0 -- Background 0xec
    "00000000", -- 7873 - 0x1ec1  :    0 - 0x0
    "00000000", -- 7874 - 0x1ec2  :    0 - 0x0
    "00000000", -- 7875 - 0x1ec3  :    0 - 0x0
    "00000000", -- 7876 - 0x1ec4  :    0 - 0x0
    "00000000", -- 7877 - 0x1ec5  :    0 - 0x0
    "11000000", -- 7878 - 0x1ec6  :  192 - 0xc0
    "00000000", -- 7879 - 0x1ec7  :    0 - 0x0
    "00000000", -- 7880 - 0x1ec8  :    0 - 0x0
    "00000000", -- 7881 - 0x1ec9  :    0 - 0x0
    "00000000", -- 7882 - 0x1eca  :    0 - 0x0
    "00000000", -- 7883 - 0x1ecb  :    0 - 0x0
    "00000000", -- 7884 - 0x1ecc  :    0 - 0x0
    "00000000", -- 7885 - 0x1ecd  :    0 - 0x0
    "00000000", -- 7886 - 0x1ece  :    0 - 0x0
    "11100000", -- 7887 - 0x1ecf  :  224 - 0xe0
    "00010000", -- 7888 - 0x1ed0  :   16 - 0x10 -- Background 0xed
    "00111000", -- 7889 - 0x1ed1  :   56 - 0x38
    "10111111", -- 7890 - 0x1ed2  :  191 - 0xbf
    "11111111", -- 7891 - 0x1ed3  :  255 - 0xff
    "11111111", -- 7892 - 0x1ed4  :  255 - 0xff
    "11111111", -- 7893 - 0x1ed5  :  255 - 0xff
    "11111111", -- 7894 - 0x1ed6  :  255 - 0xff
    "11111111", -- 7895 - 0x1ed7  :  255 - 0xff
    "11111000", -- 7896 - 0x1ed8  :  248 - 0xf8
    "11111111", -- 7897 - 0x1ed9  :  255 - 0xff
    "11111111", -- 7898 - 0x1eda  :  255 - 0xff
    "11111111", -- 7899 - 0x1edb  :  255 - 0xff
    "11111111", -- 7900 - 0x1edc  :  255 - 0xff
    "11111111", -- 7901 - 0x1edd  :  255 - 0xff
    "11111111", -- 7902 - 0x1ede  :  255 - 0xff
    "11111111", -- 7903 - 0x1edf  :  255 - 0xff
    "01111110", -- 7904 - 0x1ee0  :  126 - 0x7e -- Background 0xee
    "00011110", -- 7905 - 0x1ee1  :   30 - 0x1e
    "00011110", -- 7906 - 0x1ee2  :   30 - 0x1e
    "00001110", -- 7907 - 0x1ee3  :   14 - 0xe
    "00001111", -- 7908 - 0x1ee4  :   15 - 0xf
    "00011110", -- 7909 - 0x1ee5  :   30 - 0x1e
    "00011110", -- 7910 - 0x1ee6  :   30 - 0x1e
    "00111110", -- 7911 - 0x1ee7  :   62 - 0x3e
    "11111111", -- 7912 - 0x1ee8  :  255 - 0xff
    "01111111", -- 7913 - 0x1ee9  :  127 - 0x7f
    "00011111", -- 7914 - 0x1eea  :   31 - 0x1f
    "00001111", -- 7915 - 0x1eeb  :   15 - 0xf
    "00001111", -- 7916 - 0x1eec  :   15 - 0xf
    "10011111", -- 7917 - 0x1eed  :  159 - 0x9f
    "10011111", -- 7918 - 0x1eee  :  159 - 0x9f
    "10111111", -- 7919 - 0x1eef  :  191 - 0xbf
    "01111111", -- 7920 - 0x1ef0  :  127 - 0x7f -- Background 0xef
    "01111111", -- 7921 - 0x1ef1  :  127 - 0x7f
    "10111111", -- 7922 - 0x1ef2  :  191 - 0xbf
    "11111111", -- 7923 - 0x1ef3  :  255 - 0xff
    "11111111", -- 7924 - 0x1ef4  :  255 - 0xff
    "11111111", -- 7925 - 0x1ef5  :  255 - 0xff
    "11100111", -- 7926 - 0x1ef6  :  231 - 0xe7
    "11000000", -- 7927 - 0x1ef7  :  192 - 0xc0
    "01111111", -- 7928 - 0x1ef8  :  127 - 0x7f
    "11111111", -- 7929 - 0x1ef9  :  255 - 0xff
    "11111111", -- 7930 - 0x1efa  :  255 - 0xff
    "11111111", -- 7931 - 0x1efb  :  255 - 0xff
    "11111111", -- 7932 - 0x1efc  :  255 - 0xff
    "11111111", -- 7933 - 0x1efd  :  255 - 0xff
    "11111111", -- 7934 - 0x1efe  :  255 - 0xff
    "11001111", -- 7935 - 0x1eff  :  207 - 0xcf
    "00000000", -- 7936 - 0x1f00  :    0 - 0x0 -- Background 0xf0
    "00000000", -- 7937 - 0x1f01  :    0 - 0x0
    "00010000", -- 7938 - 0x1f02  :   16 - 0x10
    "11111101", -- 7939 - 0x1f03  :  253 - 0xfd
    "11111010", -- 7940 - 0x1f04  :  250 - 0xfa
    "11101011", -- 7941 - 0x1f05  :  235 - 0xeb
    "10000000", -- 7942 - 0x1f06  :  128 - 0x80
    "00000000", -- 7943 - 0x1f07  :    0 - 0x0
    "00000000", -- 7944 - 0x1f08  :    0 - 0x0
    "00000000", -- 7945 - 0x1f09  :    0 - 0x0
    "11110000", -- 7946 - 0x1f0a  :  240 - 0xf0
    "11111111", -- 7947 - 0x1f0b  :  255 - 0xff
    "11111111", -- 7948 - 0x1f0c  :  255 - 0xff
    "11111111", -- 7949 - 0x1f0d  :  255 - 0xff
    "11111111", -- 7950 - 0x1f0e  :  255 - 0xff
    "11111111", -- 7951 - 0x1f0f  :  255 - 0xff
    "00100000", -- 7952 - 0x1f10  :   32 - 0x20 -- Background 0xf1
    "00011111", -- 7953 - 0x1f11  :   31 - 0x1f
    "01100000", -- 7954 - 0x1f12  :   96 - 0x60
    "10001110", -- 7955 - 0x1f13  :  142 - 0x8e
    "00111111", -- 7956 - 0x1f14  :   63 - 0x3f
    "01111111", -- 7957 - 0x1f15  :  127 - 0x7f
    "01111111", -- 7958 - 0x1f16  :  127 - 0x7f
    "01111100", -- 7959 - 0x1f17  :  124 - 0x7c
    "11111111", -- 7960 - 0x1f18  :  255 - 0xff
    "11111111", -- 7961 - 0x1f19  :  255 - 0xff
    "11111111", -- 7962 - 0x1f1a  :  255 - 0xff
    "11110001", -- 7963 - 0x1f1b  :  241 - 0xf1
    "11000100", -- 7964 - 0x1f1c  :  196 - 0xc4
    "11101110", -- 7965 - 0x1f1d  :  238 - 0xee
    "11000100", -- 7966 - 0x1f1e  :  196 - 0xc4
    "10000011", -- 7967 - 0x1f1f  :  131 - 0x83
    "00111001", -- 7968 - 0x1f20  :   57 - 0x39 -- Background 0xf2
    "00110110", -- 7969 - 0x1f21  :   54 - 0x36
    "00101110", -- 7970 - 0x1f22  :   46 - 0x2e
    "10101111", -- 7971 - 0x1f23  :  175 - 0xaf
    "10101110", -- 7972 - 0x1f24  :  174 - 0xae
    "11010001", -- 7973 - 0x1f25  :  209 - 0xd1
    "11101111", -- 7974 - 0x1f26  :  239 - 0xef
    "10000111", -- 7975 - 0x1f27  :  135 - 0x87
    "11000111", -- 7976 - 0x1f28  :  199 - 0xc7
    "11111001", -- 7977 - 0x1f29  :  249 - 0xf9
    "11110000", -- 7978 - 0x1f2a  :  240 - 0xf0
    "11110000", -- 7979 - 0x1f2b  :  240 - 0xf0
    "10110001", -- 7980 - 0x1f2c  :  177 - 0xb1
    "11011111", -- 7981 - 0x1f2d  :  223 - 0xdf
    "11101111", -- 7982 - 0x1f2e  :  239 - 0xef
    "10000111", -- 7983 - 0x1f2f  :  135 - 0x87
    "00000000", -- 7984 - 0x1f30  :    0 - 0x0 -- Background 0xf3
    "00000000", -- 7985 - 0x1f31  :    0 - 0x0
    "00000100", -- 7986 - 0x1f32  :    4 - 0x4
    "01011111", -- 7987 - 0x1f33  :   95 - 0x5f
    "10101111", -- 7988 - 0x1f34  :  175 - 0xaf
    "01010011", -- 7989 - 0x1f35  :   83 - 0x53
    "00000000", -- 7990 - 0x1f36  :    0 - 0x0
    "00000000", -- 7991 - 0x1f37  :    0 - 0x0
    "00000000", -- 7992 - 0x1f38  :    0 - 0x0
    "00000000", -- 7993 - 0x1f39  :    0 - 0x0
    "00000111", -- 7994 - 0x1f3a  :    7 - 0x7
    "11111111", -- 7995 - 0x1f3b  :  255 - 0xff
    "11111111", -- 7996 - 0x1f3c  :  255 - 0xff
    "11111111", -- 7997 - 0x1f3d  :  255 - 0xff
    "11111111", -- 7998 - 0x1f3e  :  255 - 0xff
    "11111111", -- 7999 - 0x1f3f  :  255 - 0xff
    "00000010", -- 8000 - 0x1f40  :    2 - 0x2 -- Background 0xf4
    "11111100", -- 8001 - 0x1f41  :  252 - 0xfc
    "00000011", -- 8002 - 0x1f42  :    3 - 0x3
    "00111000", -- 8003 - 0x1f43  :   56 - 0x38
    "11111110", -- 8004 - 0x1f44  :  254 - 0xfe
    "11111111", -- 8005 - 0x1f45  :  255 - 0xff
    "11111111", -- 8006 - 0x1f46  :  255 - 0xff
    "00011110", -- 8007 - 0x1f47  :   30 - 0x1e
    "11111111", -- 8008 - 0x1f48  :  255 - 0xff
    "11111111", -- 8009 - 0x1f49  :  255 - 0xff
    "11111111", -- 8010 - 0x1f4a  :  255 - 0xff
    "11000111", -- 8011 - 0x1f4b  :  199 - 0xc7
    "01000101", -- 8012 - 0x1f4c  :   69 - 0x45
    "11101110", -- 8013 - 0x1f4d  :  238 - 0xee
    "01000100", -- 8014 - 0x1f4e  :   68 - 0x44
    "11100001", -- 8015 - 0x1f4f  :  225 - 0xe1
    "11000000", -- 8016 - 0x1f50  :  192 - 0xc0 -- Background 0xf5
    "00110110", -- 8017 - 0x1f51  :   54 - 0x36
    "00111110", -- 8018 - 0x1f52  :   62 - 0x3e
    "01111010", -- 8019 - 0x1f53  :  122 - 0x7a
    "10110110", -- 8020 - 0x1f54  :  182 - 0xb6
    "11001101", -- 8021 - 0x1f55  :  205 - 0xcd
    "11111011", -- 8022 - 0x1f56  :  251 - 0xfb
    "11110000", -- 8023 - 0x1f57  :  240 - 0xf0
    "11111111", -- 8024 - 0x1f58  :  255 - 0xff
    "11001111", -- 8025 - 0x1f59  :  207 - 0xcf
    "10000111", -- 8026 - 0x1f5a  :  135 - 0x87
    "10000111", -- 8027 - 0x1f5b  :  135 - 0x87
    "11001110", -- 8028 - 0x1f5c  :  206 - 0xce
    "11111101", -- 8029 - 0x1f5d  :  253 - 0xfd
    "11111011", -- 8030 - 0x1f5e  :  251 - 0xfb
    "11110000", -- 8031 - 0x1f5f  :  240 - 0xf0
    "00000000", -- 8032 - 0x1f60  :    0 - 0x0 -- Background 0xf6
    "00000000", -- 8033 - 0x1f61  :    0 - 0x0
    "00000000", -- 8034 - 0x1f62  :    0 - 0x0
    "00000000", -- 8035 - 0x1f63  :    0 - 0x0
    "00000000", -- 8036 - 0x1f64  :    0 - 0x0
    "00001110", -- 8037 - 0x1f65  :   14 - 0xe
    "00001000", -- 8038 - 0x1f66  :    8 - 0x8
    "00001000", -- 8039 - 0x1f67  :    8 - 0x8
    "00000000", -- 8040 - 0x1f68  :    0 - 0x0
    "00000000", -- 8041 - 0x1f69  :    0 - 0x0
    "00000000", -- 8042 - 0x1f6a  :    0 - 0x0
    "00000000", -- 8043 - 0x1f6b  :    0 - 0x0
    "00000000", -- 8044 - 0x1f6c  :    0 - 0x0
    "00000001", -- 8045 - 0x1f6d  :    1 - 0x1
    "00000111", -- 8046 - 0x1f6e  :    7 - 0x7
    "00001111", -- 8047 - 0x1f6f  :   15 - 0xf
    "00011111", -- 8048 - 0x1f70  :   31 - 0x1f -- Background 0xf7
    "00111111", -- 8049 - 0x1f71  :   63 - 0x3f
    "11111111", -- 8050 - 0x1f72  :  255 - 0xff
    "11111111", -- 8051 - 0x1f73  :  255 - 0xff
    "11111111", -- 8052 - 0x1f74  :  255 - 0xff
    "11111111", -- 8053 - 0x1f75  :  255 - 0xff
    "11111111", -- 8054 - 0x1f76  :  255 - 0xff
    "01111111", -- 8055 - 0x1f77  :  127 - 0x7f
    "00111111", -- 8056 - 0x1f78  :   63 - 0x3f
    "11111111", -- 8057 - 0x1f79  :  255 - 0xff
    "11111111", -- 8058 - 0x1f7a  :  255 - 0xff
    "11111111", -- 8059 - 0x1f7b  :  255 - 0xff
    "11111111", -- 8060 - 0x1f7c  :  255 - 0xff
    "11111111", -- 8061 - 0x1f7d  :  255 - 0xff
    "11111111", -- 8062 - 0x1f7e  :  255 - 0xff
    "11111111", -- 8063 - 0x1f7f  :  255 - 0xff
    "00111111", -- 8064 - 0x1f80  :   63 - 0x3f -- Background 0xf8
    "00111110", -- 8065 - 0x1f81  :   62 - 0x3e
    "00111100", -- 8066 - 0x1f82  :   60 - 0x3c
    "10111000", -- 8067 - 0x1f83  :  184 - 0xb8
    "01111000", -- 8068 - 0x1f84  :  120 - 0x78
    "01111000", -- 8069 - 0x1f85  :  120 - 0x78
    "01111110", -- 8070 - 0x1f86  :  126 - 0x7e
    "01111110", -- 8071 - 0x1f87  :  126 - 0x7e
    "11111111", -- 8072 - 0x1f88  :  255 - 0xff
    "11111111", -- 8073 - 0x1f89  :  255 - 0xff
    "11111101", -- 8074 - 0x1f8a  :  253 - 0xfd
    "11111000", -- 8075 - 0x1f8b  :  248 - 0xf8
    "11111111", -- 8076 - 0x1f8c  :  255 - 0xff
    "11111111", -- 8077 - 0x1f8d  :  255 - 0xff
    "11111110", -- 8078 - 0x1f8e  :  254 - 0xfe
    "11111111", -- 8079 - 0x1f8f  :  255 - 0xff
    "11111101", -- 8080 - 0x1f90  :  253 - 0xfd -- Background 0xf9
    "01111001", -- 8081 - 0x1f91  :  121 - 0x79
    "01111011", -- 8082 - 0x1f92  :  123 - 0x7b
    "11111111", -- 8083 - 0x1f93  :  255 - 0xff
    "11111111", -- 8084 - 0x1f94  :  255 - 0xff
    "11111111", -- 8085 - 0x1f95  :  255 - 0xff
    "11110011", -- 8086 - 0x1f96  :  243 - 0xf3
    "10000000", -- 8087 - 0x1f97  :  128 - 0x80
    "11111111", -- 8088 - 0x1f98  :  255 - 0xff
    "11111111", -- 8089 - 0x1f99  :  255 - 0xff
    "11111111", -- 8090 - 0x1f9a  :  255 - 0xff
    "11111111", -- 8091 - 0x1f9b  :  255 - 0xff
    "11111111", -- 8092 - 0x1f9c  :  255 - 0xff
    "11111111", -- 8093 - 0x1f9d  :  255 - 0xff
    "11111111", -- 8094 - 0x1f9e  :  255 - 0xff
    "11111000", -- 8095 - 0x1f9f  :  248 - 0xf8
    "00000000", -- 8096 - 0x1fa0  :    0 - 0x0 -- Background 0xfa
    "00000000", -- 8097 - 0x1fa1  :    0 - 0x0
    "00000000", -- 8098 - 0x1fa2  :    0 - 0x0
    "00000000", -- 8099 - 0x1fa3  :    0 - 0x0
    "00000000", -- 8100 - 0x1fa4  :    0 - 0x0
    "00000000", -- 8101 - 0x1fa5  :    0 - 0x0
    "00000000", -- 8102 - 0x1fa6  :    0 - 0x0
    "00000000", -- 8103 - 0x1fa7  :    0 - 0x0
    "00000000", -- 8104 - 0x1fa8  :    0 - 0x0
    "00000000", -- 8105 - 0x1fa9  :    0 - 0x0
    "00000000", -- 8106 - 0x1faa  :    0 - 0x0
    "00000000", -- 8107 - 0x1fab  :    0 - 0x0
    "00000000", -- 8108 - 0x1fac  :    0 - 0x0
    "00000000", -- 8109 - 0x1fad  :    0 - 0x0
    "11000000", -- 8110 - 0x1fae  :  192 - 0xc0
    "11110000", -- 8111 - 0x1faf  :  240 - 0xf0
    "00010000", -- 8112 - 0x1fb0  :   16 - 0x10 -- Background 0xfb
    "10000100", -- 8113 - 0x1fb1  :  132 - 0x84
    "11100000", -- 8114 - 0x1fb2  :  224 - 0xe0
    "11000000", -- 8115 - 0x1fb3  :  192 - 0xc0
    "10000000", -- 8116 - 0x1fb4  :  128 - 0x80
    "10000000", -- 8117 - 0x1fb5  :  128 - 0x80
    "00000000", -- 8118 - 0x1fb6  :    0 - 0x0
    "00000000", -- 8119 - 0x1fb7  :    0 - 0x0
    "11111100", -- 8120 - 0x1fb8  :  252 - 0xfc
    "11111110", -- 8121 - 0x1fb9  :  254 - 0xfe
    "11101100", -- 8122 - 0x1fba  :  236 - 0xec
    "11100000", -- 8123 - 0x1fbb  :  224 - 0xe0
    "11000000", -- 8124 - 0x1fbc  :  192 - 0xc0
    "11000000", -- 8125 - 0x1fbd  :  192 - 0xc0
    "10000000", -- 8126 - 0x1fbe  :  128 - 0x80
    "10000000", -- 8127 - 0x1fbf  :  128 - 0x80
    "00000000", -- 8128 - 0x1fc0  :    0 - 0x0 -- Background 0xfc
    "01001000", -- 8129 - 0x1fc1  :   72 - 0x48
    "00100000", -- 8130 - 0x1fc2  :   32 - 0x20
    "00000000", -- 8131 - 0x1fc3  :    0 - 0x0
    "00000000", -- 8132 - 0x1fc4  :    0 - 0x0
    "00000100", -- 8133 - 0x1fc5  :    4 - 0x4
    "00001110", -- 8134 - 0x1fc6  :   14 - 0xe
    "11111110", -- 8135 - 0x1fc7  :  254 - 0xfe
    "01110000", -- 8136 - 0x1fc8  :  112 - 0x70
    "11111100", -- 8137 - 0x1fc9  :  252 - 0xfc
    "11111100", -- 8138 - 0x1fca  :  252 - 0xfc
    "11111100", -- 8139 - 0x1fcb  :  252 - 0xfc
    "11111100", -- 8140 - 0x1fcc  :  252 - 0xfc
    "11111100", -- 8141 - 0x1fcd  :  252 - 0xfc
    "11111110", -- 8142 - 0x1fce  :  254 - 0xfe
    "11111110", -- 8143 - 0x1fcf  :  254 - 0xfe
    "11111110", -- 8144 - 0x1fd0  :  254 - 0xfe -- Background 0xfd
    "11111100", -- 8145 - 0x1fd1  :  252 - 0xfc
    "11111100", -- 8146 - 0x1fd2  :  252 - 0xfc
    "11111000", -- 8147 - 0x1fd3  :  248 - 0xf8
    "11110000", -- 8148 - 0x1fd4  :  240 - 0xf0
    "11100000", -- 8149 - 0x1fd5  :  224 - 0xe0
    "10000000", -- 8150 - 0x1fd6  :  128 - 0x80
    "00000000", -- 8151 - 0x1fd7  :    0 - 0x0
    "11111110", -- 8152 - 0x1fd8  :  254 - 0xfe
    "11111100", -- 8153 - 0x1fd9  :  252 - 0xfc
    "11111100", -- 8154 - 0x1fda  :  252 - 0xfc
    "11111000", -- 8155 - 0x1fdb  :  248 - 0xf8
    "11110000", -- 8156 - 0x1fdc  :  240 - 0xf0
    "11100000", -- 8157 - 0x1fdd  :  224 - 0xe0
    "10000000", -- 8158 - 0x1fde  :  128 - 0x80
    "00000000", -- 8159 - 0x1fdf  :    0 - 0x0
    "00001111", -- 8160 - 0x1fe0  :   15 - 0xf -- Background 0xfe
    "00000110", -- 8161 - 0x1fe1  :    6 - 0x6
    "00000110", -- 8162 - 0x1fe2  :    6 - 0x6
    "00000110", -- 8163 - 0x1fe3  :    6 - 0x6
    "00000110", -- 8164 - 0x1fe4  :    6 - 0x6
    "00000110", -- 8165 - 0x1fe5  :    6 - 0x6
    "00001111", -- 8166 - 0x1fe6  :   15 - 0xf
    "00000000", -- 8167 - 0x1fe7  :    0 - 0x0
    "00000000", -- 8168 - 0x1fe8  :    0 - 0x0
    "00000000", -- 8169 - 0x1fe9  :    0 - 0x0
    "00000000", -- 8170 - 0x1fea  :    0 - 0x0
    "00000000", -- 8171 - 0x1feb  :    0 - 0x0
    "00000000", -- 8172 - 0x1fec  :    0 - 0x0
    "00000000", -- 8173 - 0x1fed  :    0 - 0x0
    "00000000", -- 8174 - 0x1fee  :    0 - 0x0
    "00000000", -- 8175 - 0x1fef  :    0 - 0x0
    "11110000", -- 8176 - 0x1ff0  :  240 - 0xf0 -- Background 0xff
    "01100000", -- 8177 - 0x1ff1  :   96 - 0x60
    "01100000", -- 8178 - 0x1ff2  :   96 - 0x60
    "01100110", -- 8179 - 0x1ff3  :  102 - 0x66
    "01100110", -- 8180 - 0x1ff4  :  102 - 0x66
    "01100000", -- 8181 - 0x1ff5  :   96 - 0x60
    "11110000", -- 8182 - 0x1ff6  :  240 - 0xf0
    "00000000", -- 8183 - 0x1ff7  :    0 - 0x0
    "00000000", -- 8184 - 0x1ff8  :    0 - 0x0
    "00000000", -- 8185 - 0x1ff9  :    0 - 0x0
    "00000000", -- 8186 - 0x1ffa  :    0 - 0x0
    "00000000", -- 8187 - 0x1ffb  :    0 - 0x0
    "00000000", -- 8188 - 0x1ffc  :    0 - 0x0
    "00000000", -- 8189 - 0x1ffd  :    0 - 0x0
    "00000000", -- 8190 - 0x1ffe  :    0 - 0x0
    "00000000"  -- 8191 - 0x1fff  :    0 - 0x0
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
