---   Sprites Pattern table COLOR PLANE 1
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
--- Autcmatically generated VHDL ROM from a NES memory file----


---  Original memory dump file name: lawnmower_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_LAWN_SPR_PLN1 is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(11-1 downto 0);  --2048 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_LAWN_SPR_PLN1;

architecture BEHAVIORAL of ROM_PTABLE_LAWN_SPR_PLN1 is
  signal addr_int  : natural range 0 to 2**11-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Sprite pattern Table COLOR PLANE 1
    "00000000", --    0 -  0x0  :    0 - 0x0 -- Sprite 0x0
    "00000000", --    1 -  0x1  :    0 - 0x0
    "00000000", --    2 -  0x2  :    0 - 0x0
    "00000000", --    3 -  0x3  :    0 - 0x0
    "00000000", --    4 -  0x4  :    0 - 0x0
    "00000000", --    5 -  0x5  :    0 - 0x0
    "00000000", --    6 -  0x6  :    0 - 0x0
    "00000000", --    7 -  0x7  :    0 - 0x0
    "00000000", --    8 -  0x8  :    0 - 0x0 -- Sprite 0x1
    "00000000", --    9 -  0x9  :    0 - 0x0
    "00000000", --   10 -  0xa  :    0 - 0x0
    "00000000", --   11 -  0xb  :    0 - 0x0
    "00000000", --   12 -  0xc  :    0 - 0x0
    "00000111", --   13 -  0xd  :    7 - 0x7
    "00000111", --   14 -  0xe  :    7 - 0x7
    "00000110", --   15 -  0xf  :    6 - 0x6
    "00000000", --   16 - 0x10  :    0 - 0x0 -- Sprite 0x2
    "00000000", --   17 - 0x11  :    0 - 0x0
    "00000000", --   18 - 0x12  :    0 - 0x0
    "00000000", --   19 - 0x13  :    0 - 0x0
    "00000000", --   20 - 0x14  :    0 - 0x0
    "11111111", --   21 - 0x15  :  255 - 0xff
    "11111111", --   22 - 0x16  :  255 - 0xff
    "00000000", --   23 - 0x17  :    0 - 0x0
    "00000000", --   24 - 0x18  :    0 - 0x0 -- Sprite 0x3
    "00000000", --   25 - 0x19  :    0 - 0x0
    "00000000", --   26 - 0x1a  :    0 - 0x0
    "00000000", --   27 - 0x1b  :    0 - 0x0
    "00000000", --   28 - 0x1c  :    0 - 0x0
    "11100000", --   29 - 0x1d  :  224 - 0xe0
    "11100000", --   30 - 0x1e  :  224 - 0xe0
    "01100000", --   31 - 0x1f  :   96 - 0x60
    "00000000", --   32 - 0x20  :    0 - 0x0 -- Sprite 0x4
    "00000000", --   33 - 0x21  :    0 - 0x0
    "00000000", --   34 - 0x22  :    0 - 0x0
    "00000000", --   35 - 0x23  :    0 - 0x0
    "00000000", --   36 - 0x24  :    0 - 0x0
    "00011111", --   37 - 0x25  :   31 - 0x1f
    "01111111", --   38 - 0x26  :  127 - 0x7f
    "11110000", --   39 - 0x27  :  240 - 0xf0
    "00000000", --   40 - 0x28  :    0 - 0x0 -- Sprite 0x5
    "00000000", --   41 - 0x29  :    0 - 0x0
    "00000000", --   42 - 0x2a  :    0 - 0x0
    "00000000", --   43 - 0x2b  :    0 - 0x0
    "00000000", --   44 - 0x2c  :    0 - 0x0
    "11111000", --   45 - 0x2d  :  248 - 0xf8
    "11111110", --   46 - 0x2e  :  254 - 0xfe
    "00001111", --   47 - 0x2f  :   15 - 0xf
    "00000000", --   48 - 0x30  :    0 - 0x0 -- Sprite 0x6
    "00000000", --   49 - 0x31  :    0 - 0x0
    "00000000", --   50 - 0x32  :    0 - 0x0
    "00000000", --   51 - 0x33  :    0 - 0x0
    "00000000", --   52 - 0x34  :    0 - 0x0
    "11100111", --   53 - 0x35  :  231 - 0xe7
    "11100111", --   54 - 0x36  :  231 - 0xe7
    "01100110", --   55 - 0x37  :  102 - 0x66
    "00000000", --   56 - 0x38  :    0 - 0x0 -- Sprite 0x7
    "00000000", --   57 - 0x39  :    0 - 0x0
    "00000000", --   58 - 0x3a  :    0 - 0x0
    "00000000", --   59 - 0x3b  :    0 - 0x0
    "00000000", --   60 - 0x3c  :    0 - 0x0
    "11000111", --   61 - 0x3d  :  199 - 0xc7
    "11000111", --   62 - 0x3e  :  199 - 0xc7
    "01100110", --   63 - 0x3f  :  102 - 0x66
    "00000110", --   64 - 0x40  :    6 - 0x6 -- Sprite 0x8
    "00000110", --   65 - 0x41  :    6 - 0x6
    "00000110", --   66 - 0x42  :    6 - 0x6
    "00000110", --   67 - 0x43  :    6 - 0x6
    "00000110", --   68 - 0x44  :    6 - 0x6
    "00000110", --   69 - 0x45  :    6 - 0x6
    "00000110", --   70 - 0x46  :    6 - 0x6
    "00000110", --   71 - 0x47  :    6 - 0x6
    "11111111", --   72 - 0x48  :  255 - 0xff -- Sprite 0x9
    "11111111", --   73 - 0x49  :  255 - 0xff
    "11111111", --   74 - 0x4a  :  255 - 0xff
    "11111111", --   75 - 0x4b  :  255 - 0xff
    "11111111", --   76 - 0x4c  :  255 - 0xff
    "11111111", --   77 - 0x4d  :  255 - 0xff
    "11111111", --   78 - 0x4e  :  255 - 0xff
    "11111111", --   79 - 0x4f  :  255 - 0xff
    "01100000", --   80 - 0x50  :   96 - 0x60 -- Sprite 0xa
    "01100000", --   81 - 0x51  :   96 - 0x60
    "01100000", --   82 - 0x52  :   96 - 0x60
    "01100000", --   83 - 0x53  :   96 - 0x60
    "01100000", --   84 - 0x54  :   96 - 0x60
    "01100000", --   85 - 0x55  :   96 - 0x60
    "01100000", --   86 - 0x56  :   96 - 0x60
    "01100000", --   87 - 0x57  :   96 - 0x60
    "00000001", --   88 - 0x58  :    1 - 0x1 -- Sprite 0xb
    "00000011", --   89 - 0x59  :    3 - 0x3
    "00000011", --   90 - 0x5a  :    3 - 0x3
    "00000111", --   91 - 0x5b  :    7 - 0x7
    "00000110", --   92 - 0x5c  :    6 - 0x6
    "00000110", --   93 - 0x5d  :    6 - 0x6
    "00000110", --   94 - 0x5e  :    6 - 0x6
    "00000110", --   95 - 0x5f  :    6 - 0x6
    "11000111", --   96 - 0x60  :  199 - 0xc7 -- Sprite 0xc
    "10011111", --   97 - 0x61  :  159 - 0x9f
    "00111111", --   98 - 0x62  :   63 - 0x3f
    "01111111", --   99 - 0x63  :  127 - 0x7f
    "01111111", --  100 - 0x64  :  127 - 0x7f
    "11111111", --  101 - 0x65  :  255 - 0xff
    "11111111", --  102 - 0x66  :  255 - 0xff
    "11111111", --  103 - 0x67  :  255 - 0xff
    "11100011", --  104 - 0x68  :  227 - 0xe3 -- Sprite 0xd
    "11111001", --  105 - 0x69  :  249 - 0xf9
    "11111100", --  106 - 0x6a  :  252 - 0xfc
    "11111110", --  107 - 0x6b  :  254 - 0xfe
    "11111110", --  108 - 0x6c  :  254 - 0xfe
    "11111111", --  109 - 0x6d  :  255 - 0xff
    "11111111", --  110 - 0x6e  :  255 - 0xff
    "11111111", --  111 - 0x6f  :  255 - 0xff
    "10000110", --  112 - 0x70  :  134 - 0x86 -- Sprite 0xe
    "11000110", --  113 - 0x71  :  198 - 0xc6
    "11000110", --  114 - 0x72  :  198 - 0xc6
    "11100110", --  115 - 0x73  :  230 - 0xe6
    "01100110", --  116 - 0x74  :  102 - 0x66
    "01100110", --  117 - 0x75  :  102 - 0x66
    "01100110", --  118 - 0x76  :  102 - 0x66
    "01100110", --  119 - 0x77  :  102 - 0x66
    "01100110", --  120 - 0x78  :  102 - 0x66 -- Sprite 0xf
    "01100110", --  121 - 0x79  :  102 - 0x66
    "01100110", --  122 - 0x7a  :  102 - 0x66
    "01100110", --  123 - 0x7b  :  102 - 0x66
    "01100110", --  124 - 0x7c  :  102 - 0x66
    "01100110", --  125 - 0x7d  :  102 - 0x66
    "01100110", --  126 - 0x7e  :  102 - 0x66
    "01100110", --  127 - 0x7f  :  102 - 0x66
    "01100110", --  128 - 0x80  :  102 - 0x66 -- Sprite 0x10
    "00110110", --  129 - 0x81  :   54 - 0x36
    "10110110", --  130 - 0x82  :  182 - 0xb6
    "10011110", --  131 - 0x83  :  158 - 0x9e
    "11011110", --  132 - 0x84  :  222 - 0xde
    "11001110", --  133 - 0x85  :  206 - 0xce
    "11101110", --  134 - 0x86  :  238 - 0xee
    "11100110", --  135 - 0x87  :  230 - 0xe6
    "10000001", --  136 - 0x88  :  129 - 0x81 -- Sprite 0x11
    "00111100", --  137 - 0x89  :   60 - 0x3c
    "01111110", --  138 - 0x8a  :  126 - 0x7e
    "01100110", --  139 - 0x8b  :  102 - 0x66
    "01100110", --  140 - 0x8c  :  102 - 0x66
    "01100110", --  141 - 0x8d  :  102 - 0x66
    "01100110", --  142 - 0x8e  :  102 - 0x66
    "01100110", --  143 - 0x8f  :  102 - 0x66
    "11110110", --  144 - 0x90  :  246 - 0xf6 -- Sprite 0x12
    "11110010", --  145 - 0x91  :  242 - 0xf2
    "11111010", --  146 - 0x92  :  250 - 0xfa
    "11111000", --  147 - 0x93  :  248 - 0xf8
    "11111100", --  148 - 0x94  :  252 - 0xfc
    "11111100", --  149 - 0x95  :  252 - 0xfc
    "11111110", --  150 - 0x96  :  254 - 0xfe
    "11111110", --  151 - 0x97  :  254 - 0xfe
    "01100110", --  152 - 0x98  :  102 - 0x66 -- Sprite 0x13
    "01100110", --  153 - 0x99  :  102 - 0x66
    "01100110", --  154 - 0x9a  :  102 - 0x66
    "01100110", --  155 - 0x9b  :  102 - 0x66
    "01100110", --  156 - 0x9c  :  102 - 0x66
    "01100110", --  157 - 0x9d  :  102 - 0x66
    "01100110", --  158 - 0x9e  :  102 - 0x66
    "01111110", --  159 - 0x9f  :  126 - 0x7e
    "11111111", --  160 - 0xa0  :  255 - 0xff -- Sprite 0x14
    "01111111", --  161 - 0xa1  :  127 - 0x7f
    "01111111", --  162 - 0xa2  :  127 - 0x7f
    "00111111", --  163 - 0xa3  :   63 - 0x3f
    "00111111", --  164 - 0xa4  :   63 - 0x3f
    "00011111", --  165 - 0xa5  :   31 - 0x1f
    "01011111", --  166 - 0xa6  :   95 - 0x5f
    "01001111", --  167 - 0xa7  :   79 - 0x4f
    "01100110", --  168 - 0xa8  :  102 - 0x66 -- Sprite 0x15
    "01100110", --  169 - 0xa9  :  102 - 0x66
    "01100110", --  170 - 0xaa  :  102 - 0x66
    "01100110", --  171 - 0xab  :  102 - 0x66
    "01100110", --  172 - 0xac  :  102 - 0x66
    "01111110", --  173 - 0xad  :  126 - 0x7e
    "01111110", --  174 - 0xae  :  126 - 0x7e
    "00000000", --  175 - 0xaf  :    0 - 0x0
    "01111110", --  176 - 0xb0  :  126 - 0x7e -- Sprite 0x16
    "01100110", --  177 - 0xb1  :  102 - 0x66
    "01000010", --  178 - 0xb2  :   66 - 0x42
    "00011000", --  179 - 0xb3  :   24 - 0x18
    "00111100", --  180 - 0xb4  :   60 - 0x3c
    "01111110", --  181 - 0xb5  :  126 - 0x7e
    "11111111", --  182 - 0xb6  :  255 - 0xff
    "11111111", --  183 - 0xb7  :  255 - 0xff
    "01101111", --  184 - 0xb8  :  111 - 0x6f -- Sprite 0x17
    "01100111", --  185 - 0xb9  :  103 - 0x67
    "01110111", --  186 - 0xba  :  119 - 0x77
    "01110011", --  187 - 0xbb  :  115 - 0x73
    "01111011", --  188 - 0xbc  :  123 - 0x7b
    "01111001", --  189 - 0xbd  :  121 - 0x79
    "01101101", --  190 - 0xbe  :  109 - 0x6d
    "01101100", --  191 - 0xbf  :  108 - 0x6c
    "01100000", --  192 - 0xc0  :   96 - 0x60 -- Sprite 0x18
    "01100000", --  193 - 0xc1  :   96 - 0x60
    "01100000", --  194 - 0xc2  :   96 - 0x60
    "01100000", --  195 - 0xc3  :   96 - 0x60
    "01100000", --  196 - 0xc4  :   96 - 0x60
    "01111111", --  197 - 0xc5  :  127 - 0x7f
    "01111111", --  198 - 0xc6  :  127 - 0x7f
    "00000000", --  199 - 0xc7  :    0 - 0x0
    "00000110", --  200 - 0xc8  :    6 - 0x6 -- Sprite 0x19
    "00000110", --  201 - 0xc9  :    6 - 0x6
    "00000110", --  202 - 0xca  :    6 - 0x6
    "00000110", --  203 - 0xcb  :    6 - 0x6
    "00000110", --  204 - 0xcc  :    6 - 0x6
    "11100110", --  205 - 0xcd  :  230 - 0xe6
    "11100110", --  206 - 0xce  :  230 - 0xe6
    "01100110", --  207 - 0xcf  :  102 - 0x66
    "11111111", --  208 - 0xd0  :  255 - 0xff -- Sprite 0x1a
    "11111111", --  209 - 0xd1  :  255 - 0xff
    "11111111", --  210 - 0xd2  :  255 - 0xff
    "11111111", --  211 - 0xd3  :  255 - 0xff
    "11100111", --  212 - 0xd4  :  231 - 0xe7
    "11000011", --  213 - 0xd5  :  195 - 0xc3
    "10011001", --  214 - 0xd6  :  153 - 0x99
    "00111100", --  215 - 0xd7  :   60 - 0x3c
    "00000000", --  216 - 0xd8  :    0 - 0x0 -- Sprite 0x1b
    "01111110", --  217 - 0xd9  :  126 - 0x7e
    "01111110", --  218 - 0xda  :  126 - 0x7e
    "01100110", --  219 - 0xdb  :  102 - 0x66
    "01100110", --  220 - 0xdc  :  102 - 0x66
    "01100110", --  221 - 0xdd  :  102 - 0x66
    "01100110", --  222 - 0xde  :  102 - 0x66
    "01100110", --  223 - 0xdf  :  102 - 0x66
    "11111110", --  224 - 0xe0  :  254 - 0xfe -- Sprite 0x1c
    "11111100", --  225 - 0xe1  :  252 - 0xfc
    "11111001", --  226 - 0xe2  :  249 - 0xf9
    "11110011", --  227 - 0xe3  :  243 - 0xf3
    "11100111", --  228 - 0xe4  :  231 - 0xe7
    "11001110", --  229 - 0xe5  :  206 - 0xce
    "10011100", --  230 - 0xe6  :  156 - 0x9c
    "00111000", --  231 - 0xe7  :   56 - 0x38
    "01111110", --  232 - 0xe8  :  126 - 0x7e -- Sprite 0x1d
    "11100111", --  233 - 0xe9  :  231 - 0xe7
    "11000011", --  234 - 0xea  :  195 - 0xc3
    "10000001", --  235 - 0xeb  :  129 - 0x81
    "00000000", --  236 - 0xec  :    0 - 0x0
    "00000000", --  237 - 0xed  :    0 - 0x0
    "00000000", --  238 - 0xee  :    0 - 0x0
    "00000000", --  239 - 0xef  :    0 - 0x0
    "01111111", --  240 - 0xf0  :  127 - 0x7f -- Sprite 0x1e
    "00111111", --  241 - 0xf1  :   63 - 0x3f
    "10011111", --  242 - 0xf2  :  159 - 0x9f
    "11001111", --  243 - 0xf3  :  207 - 0xcf
    "11100111", --  244 - 0xf4  :  231 - 0xe7
    "01110011", --  245 - 0xf5  :  115 - 0x73
    "00111001", --  246 - 0xf6  :   57 - 0x39
    "00011100", --  247 - 0xf7  :   28 - 0x1c
    "00000110", --  248 - 0xf8  :    6 - 0x6 -- Sprite 0x1f
    "00000111", --  249 - 0xf9  :    7 - 0x7
    "00000111", --  250 - 0xfa  :    7 - 0x7
    "00000000", --  251 - 0xfb  :    0 - 0x0
    "00000000", --  252 - 0xfc  :    0 - 0x0
    "00000000", --  253 - 0xfd  :    0 - 0x0
    "00000000", --  254 - 0xfe  :    0 - 0x0
    "00000000", --  255 - 0xff  :    0 - 0x0
    "00000000", --  256 - 0x100  :    0 - 0x0 -- Sprite 0x20
    "11111111", --  257 - 0x101  :  255 - 0xff
    "11111111", --  258 - 0x102  :  255 - 0xff
    "00000000", --  259 - 0x103  :    0 - 0x0
    "00000000", --  260 - 0x104  :    0 - 0x0
    "00000000", --  261 - 0x105  :    0 - 0x0
    "00000000", --  262 - 0x106  :    0 - 0x0
    "00000000", --  263 - 0x107  :    0 - 0x0
    "01100110", --  264 - 0x108  :  102 - 0x66 -- Sprite 0x21
    "11100111", --  265 - 0x109  :  231 - 0xe7
    "11100111", --  266 - 0x10a  :  231 - 0xe7
    "00000000", --  267 - 0x10b  :    0 - 0x0
    "00000000", --  268 - 0x10c  :    0 - 0x0
    "00000000", --  269 - 0x10d  :    0 - 0x0
    "00000000", --  270 - 0x10e  :    0 - 0x0
    "00000000", --  271 - 0x10f  :    0 - 0x0
    "01110000", --  272 - 0x110  :  112 - 0x70 -- Sprite 0x22
    "11100000", --  273 - 0x111  :  224 - 0xe0
    "11000000", --  274 - 0x112  :  192 - 0xc0
    "00000000", --  275 - 0x113  :    0 - 0x0
    "00000000", --  276 - 0x114  :    0 - 0x0
    "00000000", --  277 - 0x115  :    0 - 0x0
    "00000000", --  278 - 0x116  :    0 - 0x0
    "00000000", --  279 - 0x117  :    0 - 0x0
    "00001110", --  280 - 0x118  :   14 - 0xe -- Sprite 0x23
    "00000111", --  281 - 0x119  :    7 - 0x7
    "00000011", --  282 - 0x11a  :    3 - 0x3
    "00000000", --  283 - 0x11b  :    0 - 0x0
    "00000000", --  284 - 0x11c  :    0 - 0x0
    "00000000", --  285 - 0x11d  :    0 - 0x0
    "00000000", --  286 - 0x11e  :    0 - 0x0
    "00000000", --  287 - 0x11f  :    0 - 0x0
    "01100000", --  288 - 0x120  :   96 - 0x60 -- Sprite 0x24
    "11100000", --  289 - 0x121  :  224 - 0xe0
    "11100000", --  290 - 0x122  :  224 - 0xe0
    "00000000", --  291 - 0x123  :    0 - 0x0
    "00000000", --  292 - 0x124  :    0 - 0x0
    "00000000", --  293 - 0x125  :    0 - 0x0
    "00000000", --  294 - 0x126  :    0 - 0x0
    "00000000", --  295 - 0x127  :    0 - 0x0
    "00000000", --  296 - 0x128  :    0 - 0x0 -- Sprite 0x25
    "00000000", --  297 - 0x129  :    0 - 0x0
    "00000000", --  298 - 0x12a  :    0 - 0x0
    "00000000", --  299 - 0x12b  :    0 - 0x0
    "00000000", --  300 - 0x12c  :    0 - 0x0
    "11000000", --  301 - 0x12d  :  192 - 0xc0
    "11100000", --  302 - 0x12e  :  224 - 0xe0
    "01110000", --  303 - 0x12f  :  112 - 0x70
    "00000000", --  304 - 0x130  :    0 - 0x0 -- Sprite 0x26
    "00000000", --  305 - 0x131  :    0 - 0x0
    "00000000", --  306 - 0x132  :    0 - 0x0
    "00000000", --  307 - 0x133  :    0 - 0x0
    "00000000", --  308 - 0x134  :    0 - 0x0
    "00000011", --  309 - 0x135  :    3 - 0x3
    "00000111", --  310 - 0x136  :    7 - 0x7
    "00001110", --  311 - 0x137  :   14 - 0xe
    "00111000", --  312 - 0x138  :   56 - 0x38 -- Sprite 0x27
    "10011100", --  313 - 0x139  :  156 - 0x9c
    "11001110", --  314 - 0x13a  :  206 - 0xce
    "11100111", --  315 - 0x13b  :  231 - 0xe7
    "11110011", --  316 - 0x13c  :  243 - 0xf3
    "11111001", --  317 - 0x13d  :  249 - 0xf9
    "11111100", --  318 - 0x13e  :  252 - 0xfc
    "11111110", --  319 - 0x13f  :  254 - 0xfe
    "00000000", --  320 - 0x140  :    0 - 0x0 -- Sprite 0x28
    "00000000", --  321 - 0x141  :    0 - 0x0
    "00000000", --  322 - 0x142  :    0 - 0x0
    "00000000", --  323 - 0x143  :    0 - 0x0
    "10000001", --  324 - 0x144  :  129 - 0x81
    "11000011", --  325 - 0x145  :  195 - 0xc3
    "11100111", --  326 - 0x146  :  231 - 0xe7
    "01111110", --  327 - 0x147  :  126 - 0x7e
    "00011100", --  328 - 0x148  :   28 - 0x1c -- Sprite 0x29
    "00111001", --  329 - 0x149  :   57 - 0x39
    "01110011", --  330 - 0x14a  :  115 - 0x73
    "11100111", --  331 - 0x14b  :  231 - 0xe7
    "11001111", --  332 - 0x14c  :  207 - 0xcf
    "10011111", --  333 - 0x14d  :  159 - 0x9f
    "00111111", --  334 - 0x14e  :   63 - 0x3f
    "01111111", --  335 - 0x14f  :  127 - 0x7f
    "01100001", --  336 - 0x150  :   97 - 0x61 -- Sprite 0x2a
    "01100011", --  337 - 0x151  :   99 - 0x63
    "01100011", --  338 - 0x152  :   99 - 0x63
    "01100111", --  339 - 0x153  :  103 - 0x67
    "01100110", --  340 - 0x154  :  102 - 0x66
    "01100110", --  341 - 0x155  :  102 - 0x66
    "01100110", --  342 - 0x156  :  102 - 0x66
    "01100110", --  343 - 0x157  :  102 - 0x66
    "10000000", --  344 - 0x158  :  128 - 0x80 -- Sprite 0x2b
    "11000000", --  345 - 0x159  :  192 - 0xc0
    "11000000", --  346 - 0x15a  :  192 - 0xc0
    "11100000", --  347 - 0x15b  :  224 - 0xe0
    "01100000", --  348 - 0x15c  :   96 - 0x60
    "01100000", --  349 - 0x15d  :   96 - 0x60
    "01100000", --  350 - 0x15e  :   96 - 0x60
    "01100000", --  351 - 0x15f  :   96 - 0x60
    "00111100", --  352 - 0x160  :   60 - 0x3c -- Sprite 0x2c
    "10011001", --  353 - 0x161  :  153 - 0x99
    "11000011", --  354 - 0x162  :  195 - 0xc3
    "11100111", --  355 - 0x163  :  231 - 0xe7
    "11111111", --  356 - 0x164  :  255 - 0xff
    "11111111", --  357 - 0x165  :  255 - 0xff
    "11111111", --  358 - 0x166  :  255 - 0xff
    "11111111", --  359 - 0x167  :  255 - 0xff
    "00000000", --  360 - 0x168  :    0 - 0x0 -- Sprite 0x2d
    "01111111", --  361 - 0x169  :  127 - 0x7f
    "01111111", --  362 - 0x16a  :  127 - 0x7f
    "01100000", --  363 - 0x16b  :   96 - 0x60
    "01100000", --  364 - 0x16c  :   96 - 0x60
    "01100000", --  365 - 0x16d  :   96 - 0x60
    "01100000", --  366 - 0x16e  :   96 - 0x60
    "01100000", --  367 - 0x16f  :   96 - 0x60
    "01100110", --  368 - 0x170  :  102 - 0x66 -- Sprite 0x2e
    "11100110", --  369 - 0x171  :  230 - 0xe6
    "11100110", --  370 - 0x172  :  230 - 0xe6
    "00000110", --  371 - 0x173  :    6 - 0x6
    "00000110", --  372 - 0x174  :    6 - 0x6
    "00000110", --  373 - 0x175  :    6 - 0x6
    "00000110", --  374 - 0x176  :    6 - 0x6
    "00000110", --  375 - 0x177  :    6 - 0x6
    "00000001", --  376 - 0x178  :    1 - 0x1 -- Sprite 0x2f
    "01111100", --  377 - 0x179  :  124 - 0x7c
    "01111110", --  378 - 0x17a  :  126 - 0x7e
    "01100110", --  379 - 0x17b  :  102 - 0x66
    "01100110", --  380 - 0x17c  :  102 - 0x66
    "01100110", --  381 - 0x17d  :  102 - 0x66
    "01100110", --  382 - 0x17e  :  102 - 0x66
    "01100110", --  383 - 0x17f  :  102 - 0x66
    "11111111", --  384 - 0x180  :  255 - 0xff -- Sprite 0x30
    "11111111", --  385 - 0x181  :  255 - 0xff
    "01111110", --  386 - 0x182  :  126 - 0x7e
    "00111100", --  387 - 0x183  :   60 - 0x3c
    "00011000", --  388 - 0x184  :   24 - 0x18
    "01000010", --  389 - 0x185  :   66 - 0x42
    "01100110", --  390 - 0x186  :  102 - 0x66
    "01111110", --  391 - 0x187  :  126 - 0x7e
    "01100000", --  392 - 0x188  :   96 - 0x60 -- Sprite 0x31
    "01111111", --  393 - 0x189  :  127 - 0x7f
    "01111111", --  394 - 0x18a  :  127 - 0x7f
    "00000000", --  395 - 0x18b  :    0 - 0x0
    "11111111", --  396 - 0x18c  :  255 - 0xff
    "11111111", --  397 - 0x18d  :  255 - 0xff
    "11111111", --  398 - 0x18e  :  255 - 0xff
    "11111111", --  399 - 0x18f  :  255 - 0xff
    "00000000", --  400 - 0x190  :    0 - 0x0 -- Sprite 0x32
    "11111111", --  401 - 0x191  :  255 - 0xff
    "11111111", --  402 - 0x192  :  255 - 0xff
    "00000000", --  403 - 0x193  :    0 - 0x0
    "11111111", --  404 - 0x194  :  255 - 0xff
    "11111111", --  405 - 0x195  :  255 - 0xff
    "11111111", --  406 - 0x196  :  255 - 0xff
    "11111111", --  407 - 0x197  :  255 - 0xff
    "00000000", --  408 - 0x198  :    0 - 0x0 -- Sprite 0x33
    "11100000", --  409 - 0x199  :  224 - 0xe0
    "11100000", --  410 - 0x19a  :  224 - 0xe0
    "01100000", --  411 - 0x19b  :   96 - 0x60
    "01100000", --  412 - 0x19c  :   96 - 0x60
    "01100000", --  413 - 0x19d  :   96 - 0x60
    "01100000", --  414 - 0x19e  :   96 - 0x60
    "01100000", --  415 - 0x19f  :   96 - 0x60
    "01111110", --  416 - 0x1a0  :  126 - 0x7e -- Sprite 0x34
    "01100110", --  417 - 0x1a1  :  102 - 0x66
    "01100110", --  418 - 0x1a2  :  102 - 0x66
    "01100110", --  419 - 0x1a3  :  102 - 0x66
    "01100110", --  420 - 0x1a4  :  102 - 0x66
    "01100110", --  421 - 0x1a5  :  102 - 0x66
    "01100110", --  422 - 0x1a6  :  102 - 0x66
    "01100110", --  423 - 0x1a7  :  102 - 0x66
    "11111111", --  424 - 0x1a8  :  255 - 0xff -- Sprite 0x35
    "11111111", --  425 - 0x1a9  :  255 - 0xff
    "11111111", --  426 - 0x1aa  :  255 - 0xff
    "11111111", --  427 - 0x1ab  :  255 - 0xff
    "00000000", --  428 - 0x1ac  :    0 - 0x0
    "01111111", --  429 - 0x1ad  :  127 - 0x7f
    "01111111", --  430 - 0x1ae  :  127 - 0x7f
    "01100000", --  431 - 0x1af  :   96 - 0x60
    "11111111", --  432 - 0x1b0  :  255 - 0xff -- Sprite 0x36
    "11111111", --  433 - 0x1b1  :  255 - 0xff
    "11111111", --  434 - 0x1b2  :  255 - 0xff
    "11111111", --  435 - 0x1b3  :  255 - 0xff
    "00000000", --  436 - 0x1b4  :    0 - 0x0
    "11111111", --  437 - 0x1b5  :  255 - 0xff
    "11111111", --  438 - 0x1b6  :  255 - 0xff
    "00000000", --  439 - 0x1b7  :    0 - 0x0
    "01100000", --  440 - 0x1b8  :   96 - 0x60 -- Sprite 0x37
    "01100000", --  441 - 0x1b9  :   96 - 0x60
    "01100000", --  442 - 0x1ba  :   96 - 0x60
    "01100000", --  443 - 0x1bb  :   96 - 0x60
    "01100000", --  444 - 0x1bc  :   96 - 0x60
    "11100000", --  445 - 0x1bd  :  224 - 0xe0
    "11100000", --  446 - 0x1be  :  224 - 0xe0
    "00000000", --  447 - 0x1bf  :    0 - 0x0
    "01100110", --  448 - 0x1c0  :  102 - 0x66 -- Sprite 0x38
    "01100110", --  449 - 0x1c1  :  102 - 0x66
    "01100110", --  450 - 0x1c2  :  102 - 0x66
    "01100110", --  451 - 0x1c3  :  102 - 0x66
    "01100110", --  452 - 0x1c4  :  102 - 0x66
    "01111110", --  453 - 0x1c5  :  126 - 0x7e
    "01111100", --  454 - 0x1c6  :  124 - 0x7c
    "00000001", --  455 - 0x1c7  :    1 - 0x1
    "11111111", --  456 - 0x1c8  :  255 - 0xff -- Sprite 0x39
    "11111111", --  457 - 0x1c9  :  255 - 0xff
    "11111111", --  458 - 0x1ca  :  255 - 0xff
    "11111111", --  459 - 0x1cb  :  255 - 0xff
    "11111111", --  460 - 0x1cc  :  255 - 0xff
    "11111111", --  461 - 0x1cd  :  255 - 0xff
    "11111111", --  462 - 0x1ce  :  255 - 0xff
    "11111110", --  463 - 0x1cf  :  254 - 0xfe
    "01100110", --  464 - 0x1d0  :  102 - 0x66 -- Sprite 0x3a
    "01100110", --  465 - 0x1d1  :  102 - 0x66
    "01100110", --  466 - 0x1d2  :  102 - 0x66
    "01100110", --  467 - 0x1d3  :  102 - 0x66
    "01100110", --  468 - 0x1d4  :  102 - 0x66
    "01111110", --  469 - 0x1d5  :  126 - 0x7e
    "00111100", --  470 - 0x1d6  :   60 - 0x3c
    "10000001", --  471 - 0x1d7  :  129 - 0x81
    "01100000", --  472 - 0x1d8  :   96 - 0x60 -- Sprite 0x3b
    "01100000", --  473 - 0x1d9  :   96 - 0x60
    "01100000", --  474 - 0x1da  :   96 - 0x60
    "01100000", --  475 - 0x1db  :   96 - 0x60
    "01100000", --  476 - 0x1dc  :   96 - 0x60
    "01111111", --  477 - 0x1dd  :  127 - 0x7f
    "01111111", --  478 - 0x1de  :  127 - 0x7f
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "00000000", --  480 - 0x1e0  :    0 - 0x0 -- Sprite 0x3c
    "00000000", --  481 - 0x1e1  :    0 - 0x0
    "00000000", --  482 - 0x1e2  :    0 - 0x0
    "00000000", --  483 - 0x1e3  :    0 - 0x0
    "00000000", --  484 - 0x1e4  :    0 - 0x0
    "11111111", --  485 - 0x1e5  :  255 - 0xff
    "11111111", --  486 - 0x1e6  :  255 - 0xff
    "00000000", --  487 - 0x1e7  :    0 - 0x0
    "00000000", --  488 - 0x1e8  :    0 - 0x0 -- Sprite 0x3d
    "00000000", --  489 - 0x1e9  :    0 - 0x0
    "00000000", --  490 - 0x1ea  :    0 - 0x0
    "00000000", --  491 - 0x1eb  :    0 - 0x0
    "00000000", --  492 - 0x1ec  :    0 - 0x0
    "11111111", --  493 - 0x1ed  :  255 - 0xff
    "11111111", --  494 - 0x1ee  :  255 - 0xff
    "00000000", --  495 - 0x1ef  :    0 - 0x0
    "11111110", --  496 - 0x1f0  :  254 - 0xfe -- Sprite 0x3e
    "11111100", --  497 - 0x1f1  :  252 - 0xfc
    "11111001", --  498 - 0x1f2  :  249 - 0xf9
    "11110011", --  499 - 0x1f3  :  243 - 0xf3
    "11110011", --  500 - 0x1f4  :  243 - 0xf3
    "11111001", --  501 - 0x1f5  :  249 - 0xf9
    "11111100", --  502 - 0x1f6  :  252 - 0xfc
    "11111110", --  503 - 0x1f7  :  254 - 0xfe
    "11100000", --  504 - 0x1f8  :  224 - 0xe0 -- Sprite 0x3f
    "11000000", --  505 - 0x1f9  :  192 - 0xc0
    "11000000", --  506 - 0x1fa  :  192 - 0xc0
    "10000000", --  507 - 0x1fb  :  128 - 0x80
    "10000000", --  508 - 0x1fc  :  128 - 0x80
    "11000000", --  509 - 0x1fd  :  192 - 0xc0
    "11000000", --  510 - 0x1fe  :  192 - 0xc0
    "11100000", --  511 - 0x1ff  :  224 - 0xe0
    "01100110", --  512 - 0x200  :  102 - 0x66 -- Sprite 0x40
    "01100110", --  513 - 0x201  :  102 - 0x66
    "01100110", --  514 - 0x202  :  102 - 0x66
    "01100110", --  515 - 0x203  :  102 - 0x66
    "01100111", --  516 - 0x204  :  103 - 0x67
    "01100011", --  517 - 0x205  :   99 - 0x63
    "01100011", --  518 - 0x206  :   99 - 0x63
    "01100001", --  519 - 0x207  :   97 - 0x61
    "11111111", --  520 - 0x208  :  255 - 0xff -- Sprite 0x41
    "11111111", --  521 - 0x209  :  255 - 0xff
    "11111111", --  522 - 0x20a  :  255 - 0xff
    "01111111", --  523 - 0x20b  :  127 - 0x7f
    "01111111", --  524 - 0x20c  :  127 - 0x7f
    "00111111", --  525 - 0x20d  :   63 - 0x3f
    "10011111", --  526 - 0x20e  :  159 - 0x9f
    "11000111", --  527 - 0x20f  :  199 - 0xc7
    "11111111", --  528 - 0x210  :  255 - 0xff -- Sprite 0x42
    "11111111", --  529 - 0x211  :  255 - 0xff
    "11111111", --  530 - 0x212  :  255 - 0xff
    "11111110", --  531 - 0x213  :  254 - 0xfe
    "11111110", --  532 - 0x214  :  254 - 0xfe
    "11111100", --  533 - 0x215  :  252 - 0xfc
    "11111001", --  534 - 0x216  :  249 - 0xf9
    "11100011", --  535 - 0x217  :  227 - 0xe3
    "01100110", --  536 - 0x218  :  102 - 0x66 -- Sprite 0x43
    "01100110", --  537 - 0x219  :  102 - 0x66
    "01100110", --  538 - 0x21a  :  102 - 0x66
    "01100110", --  539 - 0x21b  :  102 - 0x66
    "11100110", --  540 - 0x21c  :  230 - 0xe6
    "11000110", --  541 - 0x21d  :  198 - 0xc6
    "11000110", --  542 - 0x21e  :  198 - 0xc6
    "10000110", --  543 - 0x21f  :  134 - 0x86
    "11111110", --  544 - 0x220  :  254 - 0xfe -- Sprite 0x44
    "11111111", --  545 - 0x221  :  255 - 0xff
    "11111111", --  546 - 0x222  :  255 - 0xff
    "11111111", --  547 - 0x223  :  255 - 0xff
    "11111111", --  548 - 0x224  :  255 - 0xff
    "11111111", --  549 - 0x225  :  255 - 0xff
    "11111111", --  550 - 0x226  :  255 - 0xff
    "11111111", --  551 - 0x227  :  255 - 0xff
    "01100000", --  552 - 0x228  :   96 - 0x60 -- Sprite 0x45
    "01100000", --  553 - 0x229  :   96 - 0x60
    "01100000", --  554 - 0x22a  :   96 - 0x60
    "01100000", --  555 - 0x22b  :   96 - 0x60
    "01100000", --  556 - 0x22c  :   96 - 0x60
    "01100000", --  557 - 0x22d  :   96 - 0x60
    "01100000", --  558 - 0x22e  :   96 - 0x60
    "01100000", --  559 - 0x22f  :   96 - 0x60
    "11110000", --  560 - 0x230  :  240 - 0xf0 -- Sprite 0x46
    "01111111", --  561 - 0x231  :  127 - 0x7f
    "00011111", --  562 - 0x232  :   31 - 0x1f
    "00000000", --  563 - 0x233  :    0 - 0x0
    "00000000", --  564 - 0x234  :    0 - 0x0
    "00000000", --  565 - 0x235  :    0 - 0x0
    "00000000", --  566 - 0x236  :    0 - 0x0
    "00000000", --  567 - 0x237  :    0 - 0x0
    "00001111", --  568 - 0x238  :   15 - 0xf -- Sprite 0x47
    "11111110", --  569 - 0x239  :  254 - 0xfe
    "11111000", --  570 - 0x23a  :  248 - 0xf8
    "00000000", --  571 - 0x23b  :    0 - 0x0
    "00000000", --  572 - 0x23c  :    0 - 0x0
    "00000000", --  573 - 0x23d  :    0 - 0x0
    "00000000", --  574 - 0x23e  :    0 - 0x0
    "00000000", --  575 - 0x23f  :    0 - 0x0
    "00000110", --  576 - 0x240  :    6 - 0x6 -- Sprite 0x48
    "00000111", --  577 - 0x241  :    7 - 0x7
    "00000111", --  578 - 0x242  :    7 - 0x7
    "00000000", --  579 - 0x243  :    0 - 0x0
    "00000000", --  580 - 0x244  :    0 - 0x0
    "00000000", --  581 - 0x245  :    0 - 0x0
    "00000000", --  582 - 0x246  :    0 - 0x0
    "00000000", --  583 - 0x247  :    0 - 0x0
    "00000000", --  584 - 0x248  :    0 - 0x0 -- Sprite 0x49
    "00000000", --  585 - 0x249  :    0 - 0x0
    "00000000", --  586 - 0x24a  :    0 - 0x0
    "00000000", --  587 - 0x24b  :    0 - 0x0
    "00000000", --  588 - 0x24c  :    0 - 0x0
    "00000000", --  589 - 0x24d  :    0 - 0x0
    "00000000", --  590 - 0x24e  :    0 - 0x0
    "00000000", --  591 - 0x24f  :    0 - 0x0
    "00000000", --  592 - 0x250  :    0 - 0x0 -- Sprite 0x4a
    "01110110", --  593 - 0x251  :  118 - 0x76
    "01010111", --  594 - 0x252  :   87 - 0x57
    "01010101", --  595 - 0x253  :   85 - 0x55
    "01010101", --  596 - 0x254  :   85 - 0x55
    "01110101", --  597 - 0x255  :  117 - 0x75
    "01000111", --  598 - 0x256  :   71 - 0x47
    "00000000", --  599 - 0x257  :    0 - 0x0
    "00000000", --  600 - 0x258  :    0 - 0x0 -- Sprite 0x4b
    "01110111", --  601 - 0x259  :  119 - 0x77
    "00010101", --  602 - 0x25a  :   21 - 0x15
    "01110101", --  603 - 0x25b  :  117 - 0x75
    "01000101", --  604 - 0x25c  :   69 - 0x45
    "01000101", --  605 - 0x25d  :   69 - 0x45
    "01110111", --  606 - 0x25e  :  119 - 0x77
    "00000000", --  607 - 0x25f  :    0 - 0x0
    "00000000", --  608 - 0x260  :    0 - 0x0 -- Sprite 0x4c
    "00100100", --  609 - 0x261  :   36 - 0x24
    "01101100", --  610 - 0x262  :  108 - 0x6c
    "00100100", --  611 - 0x263  :   36 - 0x24
    "00100100", --  612 - 0x264  :   36 - 0x24
    "00100100", --  613 - 0x265  :   36 - 0x24
    "00100101", --  614 - 0x266  :   37 - 0x25
    "00000000", --  615 - 0x267  :    0 - 0x0
    "00000000", --  616 - 0x268  :    0 - 0x0 -- Sprite 0x4d
    "01110100", --  617 - 0x269  :  116 - 0x74
    "01000111", --  618 - 0x26a  :   71 - 0x47
    "01110101", --  619 - 0x26b  :  117 - 0x75
    "00010101", --  620 - 0x26c  :   21 - 0x15
    "00010101", --  621 - 0x26d  :   21 - 0x15
    "01110101", --  622 - 0x26e  :  117 - 0x75
    "00000000", --  623 - 0x26f  :    0 - 0x0
    "00000000", --  624 - 0x270  :    0 - 0x0 -- Sprite 0x4e
    "01000000", --  625 - 0x271  :   64 - 0x40
    "00011101", --  626 - 0x272  :   29 - 0x1d
    "01010101", --  627 - 0x273  :   85 - 0x55
    "01010001", --  628 - 0x274  :   81 - 0x51
    "01010001", --  629 - 0x275  :   81 - 0x51
    "01010001", --  630 - 0x276  :   81 - 0x51
    "00000000", --  631 - 0x277  :    0 - 0x0
    "00000000", --  632 - 0x278  :    0 - 0x0 -- Sprite 0x4f
    "00000000", --  633 - 0x279  :    0 - 0x0
    "01001000", --  634 - 0x27a  :   72 - 0x48
    "01000001", --  635 - 0x27b  :   65 - 0x41
    "01000100", --  636 - 0x27c  :   68 - 0x44
    "01000000", --  637 - 0x27d  :   64 - 0x40
    "11010000", --  638 - 0x27e  :  208 - 0xd0
    "00000010", --  639 - 0x27f  :    2 - 0x2
    "00000000", --  640 - 0x280  :    0 - 0x0 -- Sprite 0x50
    "00000000", --  641 - 0x281  :    0 - 0x0
    "11111100", --  642 - 0x282  :  252 - 0xfc
    "11111110", --  643 - 0x283  :  254 - 0xfe
    "11101110", --  644 - 0x284  :  238 - 0xee
    "11101110", --  645 - 0x285  :  238 - 0xee
    "11101110", --  646 - 0x286  :  238 - 0xee
    "11101110", --  647 - 0x287  :  238 - 0xee
    "00000000", --  648 - 0x288  :    0 - 0x0 -- Sprite 0x51
    "00000000", --  649 - 0x289  :    0 - 0x0
    "11111100", --  650 - 0x28a  :  252 - 0xfc
    "11111110", --  651 - 0x28b  :  254 - 0xfe
    "11101110", --  652 - 0x28c  :  238 - 0xee
    "11101110", --  653 - 0x28d  :  238 - 0xee
    "11101110", --  654 - 0x28e  :  238 - 0xee
    "11101110", --  655 - 0x28f  :  238 - 0xee
    "00000000", --  656 - 0x290  :    0 - 0x0 -- Sprite 0x52
    "00000000", --  657 - 0x291  :    0 - 0x0
    "11111110", --  658 - 0x292  :  254 - 0xfe
    "11111110", --  659 - 0x293  :  254 - 0xfe
    "11100000", --  660 - 0x294  :  224 - 0xe0
    "11100000", --  661 - 0x295  :  224 - 0xe0
    "11111000", --  662 - 0x296  :  248 - 0xf8
    "11111000", --  663 - 0x297  :  248 - 0xf8
    "00000000", --  664 - 0x298  :    0 - 0x0 -- Sprite 0x53
    "00000000", --  665 - 0x299  :    0 - 0x0
    "01111100", --  666 - 0x29a  :  124 - 0x7c
    "11111110", --  667 - 0x29b  :  254 - 0xfe
    "11101110", --  668 - 0x29c  :  238 - 0xee
    "11100000", --  669 - 0x29d  :  224 - 0xe0
    "11111100", --  670 - 0x29e  :  252 - 0xfc
    "01111110", --  671 - 0x29f  :  126 - 0x7e
    "00000000", --  672 - 0x2a0  :    0 - 0x0 -- Sprite 0x54
    "00000000", --  673 - 0x2a1  :    0 - 0x0
    "11111110", --  674 - 0x2a2  :  254 - 0xfe
    "11111110", --  675 - 0x2a3  :  254 - 0xfe
    "00111000", --  676 - 0x2a4  :   56 - 0x38
    "00111000", --  677 - 0x2a5  :   56 - 0x38
    "00111000", --  678 - 0x2a6  :   56 - 0x38
    "00111000", --  679 - 0x2a7  :   56 - 0x38
    "00000000", --  680 - 0x2a8  :    0 - 0x0 -- Sprite 0x55
    "00000000", --  681 - 0x2a9  :    0 - 0x0
    "01111100", --  682 - 0x2aa  :  124 - 0x7c
    "11111110", --  683 - 0x2ab  :  254 - 0xfe
    "11101110", --  684 - 0x2ac  :  238 - 0xee
    "11101110", --  685 - 0x2ad  :  238 - 0xee
    "11101110", --  686 - 0x2ae  :  238 - 0xee
    "11101110", --  687 - 0x2af  :  238 - 0xee
    "00000000", --  688 - 0x2b0  :    0 - 0x0 -- Sprite 0x56
    "00000000", --  689 - 0x2b1  :    0 - 0x0
    "11100000", --  690 - 0x2b2  :  224 - 0xe0
    "11100000", --  691 - 0x2b3  :  224 - 0xe0
    "11100000", --  692 - 0x2b4  :  224 - 0xe0
    "11100000", --  693 - 0x2b5  :  224 - 0xe0
    "11100000", --  694 - 0x2b6  :  224 - 0xe0
    "11100000", --  695 - 0x2b7  :  224 - 0xe0
    "00000000", --  696 - 0x2b8  :    0 - 0x0 -- Sprite 0x57
    "00000000", --  697 - 0x2b9  :    0 - 0x0
    "11101110", --  698 - 0x2ba  :  238 - 0xee
    "11101110", --  699 - 0x2bb  :  238 - 0xee
    "11101110", --  700 - 0x2bc  :  238 - 0xee
    "11101110", --  701 - 0x2bd  :  238 - 0xee
    "11101110", --  702 - 0x2be  :  238 - 0xee
    "11101110", --  703 - 0x2bf  :  238 - 0xee
    "00000000", --  704 - 0x2c0  :    0 - 0x0 -- Sprite 0x58
    "00000000", --  705 - 0x2c1  :    0 - 0x0
    "10001110", --  706 - 0x2c2  :  142 - 0x8e
    "11001110", --  707 - 0x2c3  :  206 - 0xce
    "11101110", --  708 - 0x2c4  :  238 - 0xee
    "11111110", --  709 - 0x2c5  :  254 - 0xfe
    "11111110", --  710 - 0x2c6  :  254 - 0xfe
    "11101110", --  711 - 0x2c7  :  238 - 0xee
    "00000000", --  712 - 0x2c8  :    0 - 0x0 -- Sprite 0x59
    "00000000", --  713 - 0x2c9  :    0 - 0x0
    "11111100", --  714 - 0x2ca  :  252 - 0xfc
    "11111110", --  715 - 0x2cb  :  254 - 0xfe
    "11101110", --  716 - 0x2cc  :  238 - 0xee
    "11101110", --  717 - 0x2cd  :  238 - 0xee
    "11101110", --  718 - 0x2ce  :  238 - 0xee
    "11101110", --  719 - 0x2cf  :  238 - 0xee
    "00000000", --  720 - 0x2d0  :    0 - 0x0 -- Sprite 0x5a
    "00000000", --  721 - 0x2d1  :    0 - 0x0
    "01111100", --  722 - 0x2d2  :  124 - 0x7c
    "11111110", --  723 - 0x2d3  :  254 - 0xfe
    "11101110", --  724 - 0x2d4  :  238 - 0xee
    "11101110", --  725 - 0x2d5  :  238 - 0xee
    "11101110", --  726 - 0x2d6  :  238 - 0xee
    "11101110", --  727 - 0x2d7  :  238 - 0xee
    "00000000", --  728 - 0x2d8  :    0 - 0x0 -- Sprite 0x5b
    "00000000", --  729 - 0x2d9  :    0 - 0x0
    "11111110", --  730 - 0x2da  :  254 - 0xfe
    "11111110", --  731 - 0x2db  :  254 - 0xfe
    "11100000", --  732 - 0x2dc  :  224 - 0xe0
    "11100000", --  733 - 0x2dd  :  224 - 0xe0
    "11111000", --  734 - 0x2de  :  248 - 0xf8
    "11111000", --  735 - 0x2df  :  248 - 0xf8
    "00000000", --  736 - 0x2e0  :    0 - 0x0 -- Sprite 0x5c
    "00000000", --  737 - 0x2e1  :    0 - 0x0
    "00000000", --  738 - 0x2e2  :    0 - 0x0
    "00000000", --  739 - 0x2e3  :    0 - 0x0
    "00000000", --  740 - 0x2e4  :    0 - 0x0
    "00000000", --  741 - 0x2e5  :    0 - 0x0
    "11001100", --  742 - 0x2e6  :  204 - 0xcc
    "11001100", --  743 - 0x2e7  :  204 - 0xcc
    "00000000", --  744 - 0x2e8  :    0 - 0x0 -- Sprite 0x5d
    "00000000", --  745 - 0x2e9  :    0 - 0x0
    "11111110", --  746 - 0x2ea  :  254 - 0xfe
    "11111110", --  747 - 0x2eb  :  254 - 0xfe
    "11100000", --  748 - 0x2ec  :  224 - 0xe0
    "11100000", --  749 - 0x2ed  :  224 - 0xe0
    "11111000", --  750 - 0x2ee  :  248 - 0xf8
    "11111000", --  751 - 0x2ef  :  248 - 0xf8
    "00000000", --  752 - 0x2f0  :    0 - 0x0 -- Sprite 0x5e
    "00000000", --  753 - 0x2f1  :    0 - 0x0
    "11101110", --  754 - 0x2f2  :  238 - 0xee
    "11101110", --  755 - 0x2f3  :  238 - 0xee
    "11101110", --  756 - 0x2f4  :  238 - 0xee
    "11101110", --  757 - 0x2f5  :  238 - 0xee
    "11101110", --  758 - 0x2f6  :  238 - 0xee
    "11101110", --  759 - 0x2f7  :  238 - 0xee
    "01111110", --  760 - 0x2f8  :  126 - 0x7e -- Sprite 0x5f
    "01111110", --  761 - 0x2f9  :  126 - 0x7e
    "01111110", --  762 - 0x2fa  :  126 - 0x7e
    "01111110", --  763 - 0x2fb  :  126 - 0x7e
    "01111110", --  764 - 0x2fc  :  126 - 0x7e
    "01111110", --  765 - 0x2fd  :  126 - 0x7e
    "01111110", --  766 - 0x2fe  :  126 - 0x7e
    "01111110", --  767 - 0x2ff  :  126 - 0x7e
    "11101110", --  768 - 0x300  :  238 - 0xee -- Sprite 0x60
    "11101110", --  769 - 0x301  :  238 - 0xee
    "11111110", --  770 - 0x302  :  254 - 0xfe
    "11111100", --  771 - 0x303  :  252 - 0xfc
    "11100000", --  772 - 0x304  :  224 - 0xe0
    "11100000", --  773 - 0x305  :  224 - 0xe0
    "00000000", --  774 - 0x306  :    0 - 0x0
    "00000000", --  775 - 0x307  :    0 - 0x0
    "11101110", --  776 - 0x308  :  238 - 0xee -- Sprite 0x61
    "11101110", --  777 - 0x309  :  238 - 0xee
    "11111100", --  778 - 0x30a  :  252 - 0xfc
    "11111100", --  779 - 0x30b  :  252 - 0xfc
    "11101110", --  780 - 0x30c  :  238 - 0xee
    "11101110", --  781 - 0x30d  :  238 - 0xee
    "00000000", --  782 - 0x30e  :    0 - 0x0
    "00000000", --  783 - 0x30f  :    0 - 0x0
    "11100000", --  784 - 0x310  :  224 - 0xe0 -- Sprite 0x62
    "11100000", --  785 - 0x311  :  224 - 0xe0
    "11100000", --  786 - 0x312  :  224 - 0xe0
    "11100000", --  787 - 0x313  :  224 - 0xe0
    "11111110", --  788 - 0x314  :  254 - 0xfe
    "11111110", --  789 - 0x315  :  254 - 0xfe
    "00000000", --  790 - 0x316  :    0 - 0x0
    "00000000", --  791 - 0x317  :    0 - 0x0
    "00001110", --  792 - 0x318  :   14 - 0xe -- Sprite 0x63
    "00001110", --  793 - 0x319  :   14 - 0xe
    "00001110", --  794 - 0x31a  :   14 - 0xe
    "11101110", --  795 - 0x31b  :  238 - 0xee
    "11111110", --  796 - 0x31c  :  254 - 0xfe
    "01111100", --  797 - 0x31d  :  124 - 0x7c
    "00000000", --  798 - 0x31e  :    0 - 0x0
    "00000000", --  799 - 0x31f  :    0 - 0x0
    "00111000", --  800 - 0x320  :   56 - 0x38 -- Sprite 0x64
    "00111000", --  801 - 0x321  :   56 - 0x38
    "00111000", --  802 - 0x322  :   56 - 0x38
    "00111000", --  803 - 0x323  :   56 - 0x38
    "00111000", --  804 - 0x324  :   56 - 0x38
    "00111000", --  805 - 0x325  :   56 - 0x38
    "00000000", --  806 - 0x326  :    0 - 0x0
    "00000000", --  807 - 0x327  :    0 - 0x0
    "11101110", --  808 - 0x328  :  238 - 0xee -- Sprite 0x65
    "11101110", --  809 - 0x329  :  238 - 0xee
    "11111110", --  810 - 0x32a  :  254 - 0xfe
    "11111110", --  811 - 0x32b  :  254 - 0xfe
    "11101110", --  812 - 0x32c  :  238 - 0xee
    "11101110", --  813 - 0x32d  :  238 - 0xee
    "00000000", --  814 - 0x32e  :    0 - 0x0
    "00000000", --  815 - 0x32f  :    0 - 0x0
    "11100000", --  816 - 0x330  :  224 - 0xe0 -- Sprite 0x66
    "11100000", --  817 - 0x331  :  224 - 0xe0
    "11100000", --  818 - 0x332  :  224 - 0xe0
    "11101110", --  819 - 0x333  :  238 - 0xee
    "11111110", --  820 - 0x334  :  254 - 0xfe
    "11111110", --  821 - 0x335  :  254 - 0xfe
    "00000000", --  822 - 0x336  :    0 - 0x0
    "00000000", --  823 - 0x337  :    0 - 0x0
    "11101110", --  824 - 0x338  :  238 - 0xee -- Sprite 0x67
    "11101110", --  825 - 0x339  :  238 - 0xee
    "11111110", --  826 - 0x33a  :  254 - 0xfe
    "11111110", --  827 - 0x33b  :  254 - 0xfe
    "11101110", --  828 - 0x33c  :  238 - 0xee
    "11000110", --  829 - 0x33d  :  198 - 0xc6
    "00000000", --  830 - 0x33e  :    0 - 0x0
    "00000000", --  831 - 0x33f  :    0 - 0x0
    "11101110", --  832 - 0x340  :  238 - 0xee -- Sprite 0x68
    "11101110", --  833 - 0x341  :  238 - 0xee
    "11101110", --  834 - 0x342  :  238 - 0xee
    "11101110", --  835 - 0x343  :  238 - 0xee
    "11101110", --  836 - 0x344  :  238 - 0xee
    "11101110", --  837 - 0x345  :  238 - 0xee
    "00000000", --  838 - 0x346  :    0 - 0x0
    "00000000", --  839 - 0x347  :    0 - 0x0
    "11101110", --  840 - 0x348  :  238 - 0xee -- Sprite 0x69
    "11101110", --  841 - 0x349  :  238 - 0xee
    "11101110", --  842 - 0x34a  :  238 - 0xee
    "11101110", --  843 - 0x34b  :  238 - 0xee
    "11111110", --  844 - 0x34c  :  254 - 0xfe
    "11111100", --  845 - 0x34d  :  252 - 0xfc
    "00000000", --  846 - 0x34e  :    0 - 0x0
    "00000000", --  847 - 0x34f  :    0 - 0x0
    "11101110", --  848 - 0x350  :  238 - 0xee -- Sprite 0x6a
    "11101110", --  849 - 0x351  :  238 - 0xee
    "11101110", --  850 - 0x352  :  238 - 0xee
    "11101110", --  851 - 0x353  :  238 - 0xee
    "11111110", --  852 - 0x354  :  254 - 0xfe
    "01111100", --  853 - 0x355  :  124 - 0x7c
    "00000000", --  854 - 0x356  :    0 - 0x0
    "00000000", --  855 - 0x357  :    0 - 0x0
    "11100000", --  856 - 0x358  :  224 - 0xe0 -- Sprite 0x6b
    "11100000", --  857 - 0x359  :  224 - 0xe0
    "11100000", --  858 - 0x35a  :  224 - 0xe0
    "11100000", --  859 - 0x35b  :  224 - 0xe0
    "11111110", --  860 - 0x35c  :  254 - 0xfe
    "11111110", --  861 - 0x35d  :  254 - 0xfe
    "00000000", --  862 - 0x35e  :    0 - 0x0
    "00000000", --  863 - 0x35f  :    0 - 0x0
    "00011000", --  864 - 0x360  :   24 - 0x18 -- Sprite 0x6c
    "00011000", --  865 - 0x361  :   24 - 0x18
    "00110000", --  866 - 0x362  :   48 - 0x30
    "00110000", --  867 - 0x363  :   48 - 0x30
    "01100110", --  868 - 0x364  :  102 - 0x66
    "01100110", --  869 - 0x365  :  102 - 0x66
    "00000000", --  870 - 0x366  :    0 - 0x0
    "00000000", --  871 - 0x367  :    0 - 0x0
    "11100000", --  872 - 0x368  :  224 - 0xe0 -- Sprite 0x6d
    "11100000", --  873 - 0x369  :  224 - 0xe0
    "11100000", --  874 - 0x36a  :  224 - 0xe0
    "11100000", --  875 - 0x36b  :  224 - 0xe0
    "11100000", --  876 - 0x36c  :  224 - 0xe0
    "11100000", --  877 - 0x36d  :  224 - 0xe0
    "00000000", --  878 - 0x36e  :    0 - 0x0
    "00000000", --  879 - 0x36f  :    0 - 0x0
    "11101110", --  880 - 0x370  :  238 - 0xee -- Sprite 0x6e
    "11101110", --  881 - 0x371  :  238 - 0xee
    "11101110", --  882 - 0x372  :  238 - 0xee
    "11101110", --  883 - 0x373  :  238 - 0xee
    "11111110", --  884 - 0x374  :  254 - 0xfe
    "01111100", --  885 - 0x375  :  124 - 0x7c
    "00000000", --  886 - 0x376  :    0 - 0x0
    "00000000", --  887 - 0x377  :    0 - 0x0
    "01111110", --  888 - 0x378  :  126 - 0x7e -- Sprite 0x6f
    "01111110", --  889 - 0x379  :  126 - 0x7e
    "01111110", --  890 - 0x37a  :  126 - 0x7e
    "01111110", --  891 - 0x37b  :  126 - 0x7e
    "00111100", --  892 - 0x37c  :   60 - 0x3c
    "00111100", --  893 - 0x37d  :   60 - 0x3c
    "00000000", --  894 - 0x37e  :    0 - 0x0
    "00000000", --  895 - 0x37f  :    0 - 0x0
    "00000111", --  896 - 0x380  :    7 - 0x7 -- Sprite 0x70
    "00011111", --  897 - 0x381  :   31 - 0x1f
    "00111111", --  898 - 0x382  :   63 - 0x3f
    "00111111", --  899 - 0x383  :   63 - 0x3f
    "01111111", --  900 - 0x384  :  127 - 0x7f
    "01111111", --  901 - 0x385  :  127 - 0x7f
    "01111111", --  902 - 0x386  :  127 - 0x7f
    "01111110", --  903 - 0x387  :  126 - 0x7e
    "11100000", --  904 - 0x388  :  224 - 0xe0 -- Sprite 0x71
    "11111000", --  905 - 0x389  :  248 - 0xf8
    "11111100", --  906 - 0x38a  :  252 - 0xfc
    "11111100", --  907 - 0x38b  :  252 - 0xfc
    "11111110", --  908 - 0x38c  :  254 - 0xfe
    "11111110", --  909 - 0x38d  :  254 - 0xfe
    "11111110", --  910 - 0x38e  :  254 - 0xfe
    "01111110", --  911 - 0x38f  :  126 - 0x7e
    "01111110", --  912 - 0x390  :  126 - 0x7e -- Sprite 0x72
    "01111110", --  913 - 0x391  :  126 - 0x7e
    "01111110", --  914 - 0x392  :  126 - 0x7e
    "01111110", --  915 - 0x393  :  126 - 0x7e
    "01111110", --  916 - 0x394  :  126 - 0x7e
    "01111110", --  917 - 0x395  :  126 - 0x7e
    "01111110", --  918 - 0x396  :  126 - 0x7e
    "01111110", --  919 - 0x397  :  126 - 0x7e
    "01111110", --  920 - 0x398  :  126 - 0x7e -- Sprite 0x73
    "01111111", --  921 - 0x399  :  127 - 0x7f
    "01111111", --  922 - 0x39a  :  127 - 0x7f
    "01111111", --  923 - 0x39b  :  127 - 0x7f
    "00111111", --  924 - 0x39c  :   63 - 0x3f
    "00111111", --  925 - 0x39d  :   63 - 0x3f
    "00011111", --  926 - 0x39e  :   31 - 0x1f
    "00000111", --  927 - 0x39f  :    7 - 0x7
    "01111110", --  928 - 0x3a0  :  126 - 0x7e -- Sprite 0x74
    "11111110", --  929 - 0x3a1  :  254 - 0xfe
    "11111110", --  930 - 0x3a2  :  254 - 0xfe
    "11111110", --  931 - 0x3a3  :  254 - 0xfe
    "11111100", --  932 - 0x3a4  :  252 - 0xfc
    "11111100", --  933 - 0x3a5  :  252 - 0xfc
    "11111000", --  934 - 0x3a6  :  248 - 0xf8
    "11100000", --  935 - 0x3a7  :  224 - 0xe0
    "01111111", --  936 - 0x3a8  :  127 - 0x7f -- Sprite 0x75
    "01111111", --  937 - 0x3a9  :  127 - 0x7f
    "01111111", --  938 - 0x3aa  :  127 - 0x7f
    "01111111", --  939 - 0x3ab  :  127 - 0x7f
    "01111111", --  940 - 0x3ac  :  127 - 0x7f
    "01111111", --  941 - 0x3ad  :  127 - 0x7f
    "00000111", --  942 - 0x3ae  :    7 - 0x7
    "00000111", --  943 - 0x3af  :    7 - 0x7
    "11111110", --  944 - 0x3b0  :  254 - 0xfe -- Sprite 0x76
    "11111110", --  945 - 0x3b1  :  254 - 0xfe
    "11111110", --  946 - 0x3b2  :  254 - 0xfe
    "11111110", --  947 - 0x3b3  :  254 - 0xfe
    "11111110", --  948 - 0x3b4  :  254 - 0xfe
    "11111110", --  949 - 0x3b5  :  254 - 0xfe
    "11100000", --  950 - 0x3b6  :  224 - 0xe0
    "11100000", --  951 - 0x3b7  :  224 - 0xe0
    "00000111", --  952 - 0x3b8  :    7 - 0x7 -- Sprite 0x77
    "00000111", --  953 - 0x3b9  :    7 - 0x7
    "00000111", --  954 - 0x3ba  :    7 - 0x7
    "00000111", --  955 - 0x3bb  :    7 - 0x7
    "00000111", --  956 - 0x3bc  :    7 - 0x7
    "00000111", --  957 - 0x3bd  :    7 - 0x7
    "00000111", --  958 - 0x3be  :    7 - 0x7
    "00000111", --  959 - 0x3bf  :    7 - 0x7
    "11100000", --  960 - 0x3c0  :  224 - 0xe0 -- Sprite 0x78
    "11100000", --  961 - 0x3c1  :  224 - 0xe0
    "11100000", --  962 - 0x3c2  :  224 - 0xe0
    "11100000", --  963 - 0x3c3  :  224 - 0xe0
    "11100000", --  964 - 0x3c4  :  224 - 0xe0
    "11100000", --  965 - 0x3c5  :  224 - 0xe0
    "11100000", --  966 - 0x3c6  :  224 - 0xe0
    "11100000", --  967 - 0x3c7  :  224 - 0xe0
    "01111111", --  968 - 0x3c8  :  127 - 0x7f -- Sprite 0x79
    "01111111", --  969 - 0x3c9  :  127 - 0x7f
    "01111111", --  970 - 0x3ca  :  127 - 0x7f
    "01111111", --  971 - 0x3cb  :  127 - 0x7f
    "01111111", --  972 - 0x3cc  :  127 - 0x7f
    "01111111", --  973 - 0x3cd  :  127 - 0x7f
    "01111110", --  974 - 0x3ce  :  126 - 0x7e
    "01111110", --  975 - 0x3cf  :  126 - 0x7e
    "11111110", --  976 - 0x3d0  :  254 - 0xfe -- Sprite 0x7a
    "11111110", --  977 - 0x3d1  :  254 - 0xfe
    "11111110", --  978 - 0x3d2  :  254 - 0xfe
    "11111110", --  979 - 0x3d3  :  254 - 0xfe
    "11111110", --  980 - 0x3d4  :  254 - 0xfe
    "11111110", --  981 - 0x3d5  :  254 - 0xfe
    "00000000", --  982 - 0x3d6  :    0 - 0x0
    "00000000", --  983 - 0x3d7  :    0 - 0x0
    "01111110", --  984 - 0x3d8  :  126 - 0x7e -- Sprite 0x7b
    "01111111", --  985 - 0x3d9  :  127 - 0x7f
    "01111111", --  986 - 0x3da  :  127 - 0x7f
    "01111111", --  987 - 0x3db  :  127 - 0x7f
    "01111111", --  988 - 0x3dc  :  127 - 0x7f
    "01111111", --  989 - 0x3dd  :  127 - 0x7f
    "01111111", --  990 - 0x3de  :  127 - 0x7f
    "01111110", --  991 - 0x3df  :  126 - 0x7e
    "00000000", --  992 - 0x3e0  :    0 - 0x0 -- Sprite 0x7c
    "11110000", --  993 - 0x3e1  :  240 - 0xf0
    "11110000", --  994 - 0x3e2  :  240 - 0xf0
    "11110000", --  995 - 0x3e3  :  240 - 0xf0
    "11110000", --  996 - 0x3e4  :  240 - 0xf0
    "11110000", --  997 - 0x3e5  :  240 - 0xf0
    "11110000", --  998 - 0x3e6  :  240 - 0xf0
    "00000000", --  999 - 0x3e7  :    0 - 0x0
    "01111110", -- 1000 - 0x3e8  :  126 - 0x7e -- Sprite 0x7d
    "01111110", -- 1001 - 0x3e9  :  126 - 0x7e
    "01111111", -- 1002 - 0x3ea  :  127 - 0x7f
    "01111111", -- 1003 - 0x3eb  :  127 - 0x7f
    "01111111", -- 1004 - 0x3ec  :  127 - 0x7f
    "01111111", -- 1005 - 0x3ed  :  127 - 0x7f
    "01111111", -- 1006 - 0x3ee  :  127 - 0x7f
    "01111111", -- 1007 - 0x3ef  :  127 - 0x7f
    "00000000", -- 1008 - 0x3f0  :    0 - 0x0 -- Sprite 0x7e
    "00000000", -- 1009 - 0x3f1  :    0 - 0x0
    "11111110", -- 1010 - 0x3f2  :  254 - 0xfe
    "11111110", -- 1011 - 0x3f3  :  254 - 0xfe
    "11111110", -- 1012 - 0x3f4  :  254 - 0xfe
    "11111110", -- 1013 - 0x3f5  :  254 - 0xfe
    "11111110", -- 1014 - 0x3f6  :  254 - 0xfe
    "11111110", -- 1015 - 0x3f7  :  254 - 0xfe
    "01111110", -- 1016 - 0x3f8  :  126 - 0x7e -- Sprite 0x7f
    "11111110", -- 1017 - 0x3f9  :  254 - 0xfe
    "11111110", -- 1018 - 0x3fa  :  254 - 0xfe
    "11111110", -- 1019 - 0x3fb  :  254 - 0xfe
    "11111110", -- 1020 - 0x3fc  :  254 - 0xfe
    "11111110", -- 1021 - 0x3fd  :  254 - 0xfe
    "11111110", -- 1022 - 0x3fe  :  254 - 0xfe
    "01111110", -- 1023 - 0x3ff  :  126 - 0x7e
    "01000000", -- 1024 - 0x400  :   64 - 0x40 -- Sprite 0x80
    "00001000", -- 1025 - 0x401  :    8 - 0x8
    "00000010", -- 1026 - 0x402  :    2 - 0x2
    "00100000", -- 1027 - 0x403  :   32 - 0x20
    "00000100", -- 1028 - 0x404  :    4 - 0x4
    "01000000", -- 1029 - 0x405  :   64 - 0x40
    "00000001", -- 1030 - 0x406  :    1 - 0x1
    "00010000", -- 1031 - 0x407  :   16 - 0x10
    "00000000", -- 1032 - 0x408  :    0 - 0x0 -- Sprite 0x81
    "00010001", -- 1033 - 0x409  :   17 - 0x11
    "00000000", -- 1034 - 0x40a  :    0 - 0x0
    "00100000", -- 1035 - 0x40b  :   32 - 0x20
    "10001000", -- 1036 - 0x40c  :  136 - 0x88
    "00000010", -- 1037 - 0x40d  :    2 - 0x2
    "00100000", -- 1038 - 0x40e  :   32 - 0x20
    "01000000", -- 1039 - 0x40f  :   64 - 0x40
    "00000001", -- 1040 - 0x410  :    1 - 0x1 -- Sprite 0x82
    "00010000", -- 1041 - 0x411  :   16 - 0x10
    "01000000", -- 1042 - 0x412  :   64 - 0x40
    "00001000", -- 1043 - 0x413  :    8 - 0x8
    "00000010", -- 1044 - 0x414  :    2 - 0x2
    "00100000", -- 1045 - 0x415  :   32 - 0x20
    "00000100", -- 1046 - 0x416  :    4 - 0x4
    "01000000", -- 1047 - 0x417  :   64 - 0x40
    "00010000", -- 1048 - 0x418  :   16 - 0x10 -- Sprite 0x83
    "00000000", -- 1049 - 0x419  :    0 - 0x0
    "01000100", -- 1050 - 0x41a  :   68 - 0x44
    "00000000", -- 1051 - 0x41b  :    0 - 0x0
    "00001000", -- 1052 - 0x41c  :    8 - 0x8
    "00100010", -- 1053 - 0x41d  :   34 - 0x22
    "10000000", -- 1054 - 0x41e  :  128 - 0x80
    "00001000", -- 1055 - 0x41f  :    8 - 0x8
    "00010100", -- 1056 - 0x420  :   20 - 0x14 -- Sprite 0x84
    "10110101", -- 1057 - 0x421  :  181 - 0xb5
    "01000100", -- 1058 - 0x422  :   68 - 0x44
    "01001010", -- 1059 - 0x423  :   74 - 0x4a
    "10010010", -- 1060 - 0x424  :  146 - 0x92
    "10010010", -- 1061 - 0x425  :  146 - 0x92
    "01000100", -- 1062 - 0x426  :   68 - 0x44
    "01001001", -- 1063 - 0x427  :   73 - 0x49
    "01000010", -- 1064 - 0x428  :   66 - 0x42 -- Sprite 0x85
    "01001010", -- 1065 - 0x429  :   74 - 0x4a
    "11001010", -- 1066 - 0x42a  :  202 - 0xca
    "00101001", -- 1067 - 0x42b  :   41 - 0x29
    "10100110", -- 1068 - 0x42c  :  166 - 0xa6
    "10010010", -- 1069 - 0x42d  :  146 - 0x92
    "10001001", -- 1070 - 0x42e  :  137 - 0x89
    "00101101", -- 1071 - 0x42f  :   45 - 0x2d
    "10001000", -- 1072 - 0x430  :  136 - 0x88 -- Sprite 0x86
    "00101001", -- 1073 - 0x431  :   41 - 0x29
    "10000010", -- 1074 - 0x432  :  130 - 0x82
    "10110110", -- 1075 - 0x433  :  182 - 0xb6
    "10001000", -- 1076 - 0x434  :  136 - 0x88
    "01001001", -- 1077 - 0x435  :   73 - 0x49
    "01010010", -- 1078 - 0x436  :   82 - 0x52
    "01010010", -- 1079 - 0x437  :   82 - 0x52
    "10110010", -- 1080 - 0x438  :  178 - 0xb2 -- Sprite 0x87
    "01001010", -- 1081 - 0x439  :   74 - 0x4a
    "10101001", -- 1082 - 0x43a  :  169 - 0xa9
    "10100100", -- 1083 - 0x43b  :  164 - 0xa4
    "01100010", -- 1084 - 0x43c  :   98 - 0x62
    "01001011", -- 1085 - 0x43d  :   75 - 0x4b
    "10010000", -- 1086 - 0x43e  :  144 - 0x90
    "10010010", -- 1087 - 0x43f  :  146 - 0x92
    "00000000", -- 1088 - 0x440  :    0 - 0x0 -- Sprite 0x88
    "01100000", -- 1089 - 0x441  :   96 - 0x60
    "11111110", -- 1090 - 0x442  :  254 - 0xfe
    "11111111", -- 1091 - 0x443  :  255 - 0xff
    "01111111", -- 1092 - 0x444  :  127 - 0x7f
    "00011111", -- 1093 - 0x445  :   31 - 0x1f
    "00001110", -- 1094 - 0x446  :   14 - 0xe
    "00000000", -- 1095 - 0x447  :    0 - 0x0
    "00110000", -- 1096 - 0x448  :   48 - 0x30 -- Sprite 0x89
    "01111000", -- 1097 - 0x449  :  120 - 0x78
    "01111000", -- 1098 - 0x44a  :  120 - 0x78
    "00111110", -- 1099 - 0x44b  :   62 - 0x3e
    "00011111", -- 1100 - 0x44c  :   31 - 0x1f
    "00011111", -- 1101 - 0x44d  :   31 - 0x1f
    "00011111", -- 1102 - 0x44e  :   31 - 0x1f
    "00001110", -- 1103 - 0x44f  :   14 - 0xe
    "01000000", -- 1104 - 0x450  :   64 - 0x40 -- Sprite 0x8a
    "00001000", -- 1105 - 0x451  :    8 - 0x8
    "00000010", -- 1106 - 0x452  :    2 - 0x2
    "00101000", -- 1107 - 0x453  :   40 - 0x28
    "00010100", -- 1108 - 0x454  :   20 - 0x14
    "01010100", -- 1109 - 0x455  :   84 - 0x54
    "00000001", -- 1110 - 0x456  :    1 - 0x1
    "00010000", -- 1111 - 0x457  :   16 - 0x10
    "01000000", -- 1112 - 0x458  :   64 - 0x40 -- Sprite 0x8b
    "00000000", -- 1113 - 0x459  :    0 - 0x0
    "10010001", -- 1114 - 0x45a  :  145 - 0x91
    "00010100", -- 1115 - 0x45b  :   20 - 0x14
    "00101000", -- 1116 - 0x45c  :   40 - 0x28
    "10001010", -- 1117 - 0x45d  :  138 - 0x8a
    "01000000", -- 1118 - 0x45e  :   64 - 0x40
    "00100000", -- 1119 - 0x45f  :   32 - 0x20
    "00000000", -- 1120 - 0x460  :    0 - 0x0 -- Sprite 0x8c
    "00000111", -- 1121 - 0x461  :    7 - 0x7
    "00011111", -- 1122 - 0x462  :   31 - 0x1f
    "00111111", -- 1123 - 0x463  :   63 - 0x3f
    "00111111", -- 1124 - 0x464  :   63 - 0x3f
    "01111111", -- 1125 - 0x465  :  127 - 0x7f
    "01111111", -- 1126 - 0x466  :  127 - 0x7f
    "01111111", -- 1127 - 0x467  :  127 - 0x7f
    "00000000", -- 1128 - 0x468  :    0 - 0x0 -- Sprite 0x8d
    "11100000", -- 1129 - 0x469  :  224 - 0xe0
    "11111000", -- 1130 - 0x46a  :  248 - 0xf8
    "11111000", -- 1131 - 0x46b  :  248 - 0xf8
    "11110000", -- 1132 - 0x46c  :  240 - 0xf0
    "11111000", -- 1133 - 0x46d  :  248 - 0xf8
    "11110100", -- 1134 - 0x46e  :  244 - 0xf4
    "11111000", -- 1135 - 0x46f  :  248 - 0xf8
    "01111111", -- 1136 - 0x470  :  127 - 0x7f -- Sprite 0x8e
    "00111111", -- 1137 - 0x471  :   63 - 0x3f
    "00111111", -- 1138 - 0x472  :   63 - 0x3f
    "00011111", -- 1139 - 0x473  :   31 - 0x1f
    "00011111", -- 1140 - 0x474  :   31 - 0x1f
    "00001111", -- 1141 - 0x475  :   15 - 0xf
    "00001111", -- 1142 - 0x476  :   15 - 0xf
    "00000111", -- 1143 - 0x477  :    7 - 0x7
    "11111110", -- 1144 - 0x478  :  254 - 0xfe -- Sprite 0x8f
    "11111100", -- 1145 - 0x479  :  252 - 0xfc
    "11111100", -- 1146 - 0x47a  :  252 - 0xfc
    "11111000", -- 1147 - 0x47b  :  248 - 0xf8
    "11111000", -- 1148 - 0x47c  :  248 - 0xf8
    "11110000", -- 1149 - 0x47d  :  240 - 0xf0
    "11110000", -- 1150 - 0x47e  :  240 - 0xf0
    "11100000", -- 1151 - 0x47f  :  224 - 0xe0
    "01000001", -- 1152 - 0x480  :   65 - 0x41 -- Sprite 0x90
    "00001000", -- 1153 - 0x481  :    8 - 0x8
    "00000000", -- 1154 - 0x482  :    0 - 0x0
    "00100000", -- 1155 - 0x483  :   32 - 0x20
    "00000100", -- 1156 - 0x484  :    4 - 0x4
    "00000001", -- 1157 - 0x485  :    1 - 0x1
    "01000000", -- 1158 - 0x486  :   64 - 0x40
    "00001000", -- 1159 - 0x487  :    8 - 0x8
    "00010001", -- 1160 - 0x488  :   17 - 0x11 -- Sprite 0x91
    "00000000", -- 1161 - 0x489  :    0 - 0x0
    "10000100", -- 1162 - 0x48a  :  132 - 0x84
    "00000010", -- 1163 - 0x48b  :    2 - 0x2
    "00010000", -- 1164 - 0x48c  :   16 - 0x10
    "00000000", -- 1165 - 0x48d  :    0 - 0x0
    "01000010", -- 1166 - 0x48e  :   66 - 0x42
    "00000000", -- 1167 - 0x48f  :    0 - 0x0
    "00000100", -- 1168 - 0x490  :    4 - 0x4 -- Sprite 0x92
    "01000000", -- 1169 - 0x491  :   64 - 0x40
    "00010000", -- 1170 - 0x492  :   16 - 0x10
    "00000010", -- 1171 - 0x493  :    2 - 0x2
    "00000000", -- 1172 - 0x494  :    0 - 0x0
    "01000000", -- 1173 - 0x495  :   64 - 0x40
    "00000100", -- 1174 - 0x496  :    4 - 0x4
    "00100000", -- 1175 - 0x497  :   32 - 0x20
    "01000010", -- 1176 - 0x498  :   66 - 0x42 -- Sprite 0x93
    "00000000", -- 1177 - 0x499  :    0 - 0x0
    "10001000", -- 1178 - 0x49a  :  136 - 0x88
    "00000001", -- 1179 - 0x49b  :    1 - 0x1
    "00100000", -- 1180 - 0x49c  :   32 - 0x20
    "00000100", -- 1181 - 0x49d  :    4 - 0x4
    "00010000", -- 1182 - 0x49e  :   16 - 0x10
    "10000000", -- 1183 - 0x49f  :  128 - 0x80
    "11001000", -- 1184 - 0x4a0  :  200 - 0xc8 -- Sprite 0x94
    "00101010", -- 1185 - 0x4a1  :   42 - 0x2a
    "10100010", -- 1186 - 0x4a2  :  162 - 0xa2
    "10010100", -- 1187 - 0x4a3  :  148 - 0x94
    "10010001", -- 1188 - 0x4a4  :  145 - 0x91
    "01010101", -- 1189 - 0x4a5  :   85 - 0x55
    "01000100", -- 1190 - 0x4a6  :   68 - 0x44
    "00010010", -- 1191 - 0x4a7  :   18 - 0x12
    "10101010", -- 1192 - 0x4a8  :  170 - 0xaa -- Sprite 0x95
    "10100010", -- 1193 - 0x4a9  :  162 - 0xa2
    "00010010", -- 1194 - 0x4aa  :   18 - 0x12
    "01010011", -- 1195 - 0x4ab  :   83 - 0x53
    "01001100", -- 1196 - 0x4ac  :   76 - 0x4c
    "01010101", -- 1197 - 0x4ad  :   85 - 0x55
    "10010001", -- 1198 - 0x4ae  :  145 - 0x91
    "01001000", -- 1199 - 0x4af  :   72 - 0x48
    "01010001", -- 1200 - 0x4b0  :   81 - 0x51 -- Sprite 0x96
    "00010101", -- 1201 - 0x4b1  :   21 - 0x15
    "10100100", -- 1202 - 0x4b2  :  164 - 0xa4
    "10001100", -- 1203 - 0x4b3  :  140 - 0x8c
    "10101010", -- 1204 - 0x4b4  :  170 - 0xaa
    "00100010", -- 1205 - 0x4b5  :   34 - 0x22
    "10010000", -- 1206 - 0x4b6  :  144 - 0x90
    "01000110", -- 1207 - 0x4b7  :   70 - 0x46
    "00010011", -- 1208 - 0x4b8  :   19 - 0x13 -- Sprite 0x97
    "01010101", -- 1209 - 0x4b9  :   85 - 0x55
    "01100100", -- 1210 - 0x4ba  :  100 - 0x64
    "00010010", -- 1211 - 0x4bb  :   18 - 0x12
    "10101010", -- 1212 - 0x4bc  :  170 - 0xaa
    "10101000", -- 1213 - 0x4bd  :  168 - 0xa8
    "10000100", -- 1214 - 0x4be  :  132 - 0x84
    "11010100", -- 1215 - 0x4bf  :  212 - 0xd4
    "00110000", -- 1216 - 0x4c0  :   48 - 0x30 -- Sprite 0x98
    "01111000", -- 1217 - 0x4c1  :  120 - 0x78
    "01111000", -- 1218 - 0x4c2  :  120 - 0x78
    "00111110", -- 1219 - 0x4c3  :   62 - 0x3e
    "00011111", -- 1220 - 0x4c4  :   31 - 0x1f
    "00011111", -- 1221 - 0x4c5  :   31 - 0x1f
    "00011111", -- 1222 - 0x4c6  :   31 - 0x1f
    "00001110", -- 1223 - 0x4c7  :   14 - 0xe
    "00000000", -- 1224 - 0x4c8  :    0 - 0x0 -- Sprite 0x99
    "01100000", -- 1225 - 0x4c9  :   96 - 0x60
    "11111110", -- 1226 - 0x4ca  :  254 - 0xfe
    "11111111", -- 1227 - 0x4cb  :  255 - 0xff
    "01111111", -- 1228 - 0x4cc  :  127 - 0x7f
    "00011111", -- 1229 - 0x4cd  :   31 - 0x1f
    "00001110", -- 1230 - 0x4ce  :   14 - 0xe
    "00000000", -- 1231 - 0x4cf  :    0 - 0x0
    "01000000", -- 1232 - 0x4d0  :   64 - 0x40 -- Sprite 0x9a
    "00001100", -- 1233 - 0x4d1  :   12 - 0xc
    "00000000", -- 1234 - 0x4d2  :    0 - 0x0
    "00101000", -- 1235 - 0x4d3  :   40 - 0x28
    "00101100", -- 1236 - 0x4d4  :   44 - 0x2c
    "00010001", -- 1237 - 0x4d5  :   17 - 0x11
    "01000000", -- 1238 - 0x4d6  :   64 - 0x40
    "00001000", -- 1239 - 0x4d7  :    8 - 0x8
    "00100000", -- 1240 - 0x4d8  :   32 - 0x20 -- Sprite 0x9b
    "00000000", -- 1241 - 0x4d9  :    0 - 0x0
    "10010100", -- 1242 - 0x4da  :  148 - 0x94
    "01001000", -- 1243 - 0x4db  :   72 - 0x48
    "00011000", -- 1244 - 0x4dc  :   24 - 0x18
    "00000110", -- 1245 - 0x4dd  :    6 - 0x6
    "01000000", -- 1246 - 0x4de  :   64 - 0x40
    "00000000", -- 1247 - 0x4df  :    0 - 0x0
    "01111111", -- 1248 - 0x4e0  :  127 - 0x7f -- Sprite 0x9c
    "01111111", -- 1249 - 0x4e1  :  127 - 0x7f
    "01111111", -- 1250 - 0x4e2  :  127 - 0x7f
    "00111111", -- 1251 - 0x4e3  :   63 - 0x3f
    "00110101", -- 1252 - 0x4e4  :   53 - 0x35
    "00000010", -- 1253 - 0x4e5  :    2 - 0x2
    "00000000", -- 1254 - 0x4e6  :    0 - 0x0
    "00000000", -- 1255 - 0x4e7  :    0 - 0x0
    "11110100", -- 1256 - 0x4e8  :  244 - 0xf4 -- Sprite 0x9d
    "11111000", -- 1257 - 0x4e9  :  248 - 0xf8
    "11110000", -- 1258 - 0x4ea  :  240 - 0xf0
    "11101000", -- 1259 - 0x4eb  :  232 - 0xe8
    "01010000", -- 1260 - 0x4ec  :   80 - 0x50
    "10000000", -- 1261 - 0x4ed  :  128 - 0x80
    "00000000", -- 1262 - 0x4ee  :    0 - 0x0
    "00000000", -- 1263 - 0x4ef  :    0 - 0x0
    "11111110", -- 1264 - 0x4f0  :  254 - 0xfe -- Sprite 0x9e
    "11111100", -- 1265 - 0x4f1  :  252 - 0xfc
    "11111100", -- 1266 - 0x4f2  :  252 - 0xfc
    "11111000", -- 1267 - 0x4f3  :  248 - 0xf8
    "11111000", -- 1268 - 0x4f4  :  248 - 0xf8
    "11111100", -- 1269 - 0x4f5  :  252 - 0xfc
    "11111100", -- 1270 - 0x4f6  :  252 - 0xfc
    "11111110", -- 1271 - 0x4f7  :  254 - 0xfe
    "00000000", -- 1272 - 0x4f8  :    0 - 0x0 -- Sprite 0x9f
    "00000000", -- 1273 - 0x4f9  :    0 - 0x0
    "01111110", -- 1274 - 0x4fa  :  126 - 0x7e
    "01111110", -- 1275 - 0x4fb  :  126 - 0x7e
    "01111110", -- 1276 - 0x4fc  :  126 - 0x7e
    "01111110", -- 1277 - 0x4fd  :  126 - 0x7e
    "01111110", -- 1278 - 0x4fe  :  126 - 0x7e
    "01111110", -- 1279 - 0x4ff  :  126 - 0x7e
    "00010000", -- 1280 - 0x500  :   16 - 0x10 -- Sprite 0xa0
    "00111000", -- 1281 - 0x501  :   56 - 0x38
    "01111100", -- 1282 - 0x502  :  124 - 0x7c
    "11111000", -- 1283 - 0x503  :  248 - 0xf8
    "01110000", -- 1284 - 0x504  :  112 - 0x70
    "00100010", -- 1285 - 0x505  :   34 - 0x22
    "00000101", -- 1286 - 0x506  :    5 - 0x5
    "00000010", -- 1287 - 0x507  :    2 - 0x2
    "00010000", -- 1288 - 0x508  :   16 - 0x10 -- Sprite 0xa1
    "00111000", -- 1289 - 0x509  :   56 - 0x38
    "01111100", -- 1290 - 0x50a  :  124 - 0x7c
    "11100000", -- 1291 - 0x50b  :  224 - 0xe0
    "01100000", -- 1292 - 0x50c  :   96 - 0x60
    "00100000", -- 1293 - 0x50d  :   32 - 0x20
    "00000000", -- 1294 - 0x50e  :    0 - 0x0
    "00000000", -- 1295 - 0x50f  :    0 - 0x0
    "00010000", -- 1296 - 0x510  :   16 - 0x10 -- Sprite 0xa2
    "00111000", -- 1297 - 0x511  :   56 - 0x38
    "01111100", -- 1298 - 0x512  :  124 - 0x7c
    "00000000", -- 1299 - 0x513  :    0 - 0x0
    "00000000", -- 1300 - 0x514  :    0 - 0x0
    "00000000", -- 1301 - 0x515  :    0 - 0x0
    "00000000", -- 1302 - 0x516  :    0 - 0x0
    "00000000", -- 1303 - 0x517  :    0 - 0x0
    "00000000", -- 1304 - 0x518  :    0 - 0x0 -- Sprite 0xa3
    "00100000", -- 1305 - 0x519  :   32 - 0x20
    "01100000", -- 1306 - 0x51a  :   96 - 0x60
    "11100000", -- 1307 - 0x51b  :  224 - 0xe0
    "01100000", -- 1308 - 0x51c  :   96 - 0x60
    "00100000", -- 1309 - 0x51d  :   32 - 0x20
    "00000000", -- 1310 - 0x51e  :    0 - 0x0
    "00000000", -- 1311 - 0x51f  :    0 - 0x0
    "00000000", -- 1312 - 0x520  :    0 - 0x0 -- Sprite 0xa4
    "00100000", -- 1313 - 0x521  :   32 - 0x20
    "01100011", -- 1314 - 0x522  :   99 - 0x63
    "11100111", -- 1315 - 0x523  :  231 - 0xe7
    "01100000", -- 1316 - 0x524  :   96 - 0x60
    "00100010", -- 1317 - 0x525  :   34 - 0x22
    "00000101", -- 1318 - 0x526  :    5 - 0x5
    "00000010", -- 1319 - 0x527  :    2 - 0x2
    "00000000", -- 1320 - 0x528  :    0 - 0x0 -- Sprite 0xa5
    "00000000", -- 1321 - 0x529  :    0 - 0x0
    "11111111", -- 1322 - 0x52a  :  255 - 0xff
    "11111111", -- 1323 - 0x52b  :  255 - 0xff
    "00000000", -- 1324 - 0x52c  :    0 - 0x0
    "00100010", -- 1325 - 0x52d  :   34 - 0x22
    "00000101", -- 1326 - 0x52e  :    5 - 0x5
    "00000010", -- 1327 - 0x52f  :    2 - 0x2
    "00010000", -- 1328 - 0x530  :   16 - 0x10 -- Sprite 0xa6
    "00111000", -- 1329 - 0x531  :   56 - 0x38
    "01111100", -- 1330 - 0x532  :  124 - 0x7c
    "00000000", -- 1331 - 0x533  :    0 - 0x0
    "00000000", -- 1332 - 0x534  :    0 - 0x0
    "00010010", -- 1333 - 0x535  :   18 - 0x12
    "00110101", -- 1334 - 0x536  :   53 - 0x35
    "00110010", -- 1335 - 0x537  :   50 - 0x32
    "00110000", -- 1336 - 0x538  :   48 - 0x30 -- Sprite 0xa7
    "00110000", -- 1337 - 0x539  :   48 - 0x30
    "00110100", -- 1338 - 0x53a  :   52 - 0x34
    "00110000", -- 1339 - 0x53b  :   48 - 0x30
    "00110000", -- 1340 - 0x53c  :   48 - 0x30
    "00110010", -- 1341 - 0x53d  :   50 - 0x32
    "00110101", -- 1342 - 0x53e  :   53 - 0x35
    "00110010", -- 1343 - 0x53f  :   50 - 0x32
    "00110000", -- 1344 - 0x540  :   48 - 0x30 -- Sprite 0xa8
    "00110000", -- 1345 - 0x541  :   48 - 0x30
    "11110100", -- 1346 - 0x542  :  244 - 0xf4
    "11110000", -- 1347 - 0x543  :  240 - 0xf0
    "00000000", -- 1348 - 0x544  :    0 - 0x0
    "00100010", -- 1349 - 0x545  :   34 - 0x22
    "00000101", -- 1350 - 0x546  :    5 - 0x5
    "00000010", -- 1351 - 0x547  :    2 - 0x2
    "00000000", -- 1352 - 0x548  :    0 - 0x0 -- Sprite 0xa9
    "00000000", -- 1353 - 0x549  :    0 - 0x0
    "00000000", -- 1354 - 0x54a  :    0 - 0x0
    "00000000", -- 1355 - 0x54b  :    0 - 0x0
    "00000000", -- 1356 - 0x54c  :    0 - 0x0
    "00000000", -- 1357 - 0x54d  :    0 - 0x0
    "00000000", -- 1358 - 0x54e  :    0 - 0x0
    "00000000", -- 1359 - 0x54f  :    0 - 0x0
    "00000000", -- 1360 - 0x550  :    0 - 0x0 -- Sprite 0xaa
    "00000000", -- 1361 - 0x551  :    0 - 0x0
    "01010000", -- 1362 - 0x552  :   80 - 0x50
    "10101000", -- 1363 - 0x553  :  168 - 0xa8
    "01110000", -- 1364 - 0x554  :  112 - 0x70
    "00100010", -- 1365 - 0x555  :   34 - 0x22
    "00000101", -- 1366 - 0x556  :    5 - 0x5
    "00000010", -- 1367 - 0x557  :    2 - 0x2
    "00000000", -- 1368 - 0x558  :    0 - 0x0 -- Sprite 0xab
    "00000000", -- 1369 - 0x559  :    0 - 0x0
    "00000000", -- 1370 - 0x55a  :    0 - 0x0
    "00000000", -- 1371 - 0x55b  :    0 - 0x0
    "00000000", -- 1372 - 0x55c  :    0 - 0x0
    "00000000", -- 1373 - 0x55d  :    0 - 0x0
    "00000000", -- 1374 - 0x55e  :    0 - 0x0
    "00000000", -- 1375 - 0x55f  :    0 - 0x0
    "00000000", -- 1376 - 0x560  :    0 - 0x0 -- Sprite 0xac
    "00000000", -- 1377 - 0x561  :    0 - 0x0
    "00000000", -- 1378 - 0x562  :    0 - 0x0
    "00000000", -- 1379 - 0x563  :    0 - 0x0
    "00000000", -- 1380 - 0x564  :    0 - 0x0
    "00000000", -- 1381 - 0x565  :    0 - 0x0
    "00000000", -- 1382 - 0x566  :    0 - 0x0
    "00000000", -- 1383 - 0x567  :    0 - 0x0
    "00000000", -- 1384 - 0x568  :    0 - 0x0 -- Sprite 0xad
    "00000000", -- 1385 - 0x569  :    0 - 0x0
    "11111111", -- 1386 - 0x56a  :  255 - 0xff
    "00000000", -- 1387 - 0x56b  :    0 - 0x0
    "00000000", -- 1388 - 0x56c  :    0 - 0x0
    "00000000", -- 1389 - 0x56d  :    0 - 0x0
    "00000000", -- 1390 - 0x56e  :    0 - 0x0
    "00000000", -- 1391 - 0x56f  :    0 - 0x0
    "00000000", -- 1392 - 0x570  :    0 - 0x0 -- Sprite 0xae
    "00000000", -- 1393 - 0x571  :    0 - 0x0
    "00000000", -- 1394 - 0x572  :    0 - 0x0
    "00000000", -- 1395 - 0x573  :    0 - 0x0
    "00000000", -- 1396 - 0x574  :    0 - 0x0
    "11111111", -- 1397 - 0x575  :  255 - 0xff
    "00000000", -- 1398 - 0x576  :    0 - 0x0
    "00000000", -- 1399 - 0x577  :    0 - 0x0
    "00000000", -- 1400 - 0x578  :    0 - 0x0 -- Sprite 0xaf
    "00000000", -- 1401 - 0x579  :    0 - 0x0
    "00000000", -- 1402 - 0x57a  :    0 - 0x0
    "00000000", -- 1403 - 0x57b  :    0 - 0x0
    "00000000", -- 1404 - 0x57c  :    0 - 0x0
    "00000000", -- 1405 - 0x57d  :    0 - 0x0
    "00000000", -- 1406 - 0x57e  :    0 - 0x0
    "00000000", -- 1407 - 0x57f  :    0 - 0x0
    "00000000", -- 1408 - 0x580  :    0 - 0x0 -- Sprite 0xb0
    "00011111", -- 1409 - 0x581  :   31 - 0x1f
    "00011111", -- 1410 - 0x582  :   31 - 0x1f
    "00011111", -- 1411 - 0x583  :   31 - 0x1f
    "00011111", -- 1412 - 0x584  :   31 - 0x1f
    "00011111", -- 1413 - 0x585  :   31 - 0x1f
    "00011111", -- 1414 - 0x586  :   31 - 0x1f
    "00011111", -- 1415 - 0x587  :   31 - 0x1f
    "00000000", -- 1416 - 0x588  :    0 - 0x0 -- Sprite 0xb1
    "11110000", -- 1417 - 0x589  :  240 - 0xf0
    "11110000", -- 1418 - 0x58a  :  240 - 0xf0
    "11110000", -- 1419 - 0x58b  :  240 - 0xf0
    "11110000", -- 1420 - 0x58c  :  240 - 0xf0
    "11110000", -- 1421 - 0x58d  :  240 - 0xf0
    "11110000", -- 1422 - 0x58e  :  240 - 0xf0
    "11110000", -- 1423 - 0x58f  :  240 - 0xf0
    "00011111", -- 1424 - 0x590  :   31 - 0x1f -- Sprite 0xb2
    "00011111", -- 1425 - 0x591  :   31 - 0x1f
    "00011111", -- 1426 - 0x592  :   31 - 0x1f
    "00011111", -- 1427 - 0x593  :   31 - 0x1f
    "00000000", -- 1428 - 0x594  :    0 - 0x0
    "00000000", -- 1429 - 0x595  :    0 - 0x0
    "00000000", -- 1430 - 0x596  :    0 - 0x0
    "00000000", -- 1431 - 0x597  :    0 - 0x0
    "11110000", -- 1432 - 0x598  :  240 - 0xf0 -- Sprite 0xb3
    "11110000", -- 1433 - 0x599  :  240 - 0xf0
    "11110000", -- 1434 - 0x59a  :  240 - 0xf0
    "11110000", -- 1435 - 0x59b  :  240 - 0xf0
    "00000000", -- 1436 - 0x59c  :    0 - 0x0
    "00000000", -- 1437 - 0x59d  :    0 - 0x0
    "00000000", -- 1438 - 0x59e  :    0 - 0x0
    "00000000", -- 1439 - 0x59f  :    0 - 0x0
    "00000000", -- 1440 - 0x5a0  :    0 - 0x0 -- Sprite 0xb4
    "00000000", -- 1441 - 0x5a1  :    0 - 0x0
    "00111111", -- 1442 - 0x5a2  :   63 - 0x3f
    "01111111", -- 1443 - 0x5a3  :  127 - 0x7f
    "01111111", -- 1444 - 0x5a4  :  127 - 0x7f
    "01111111", -- 1445 - 0x5a5  :  127 - 0x7f
    "01111111", -- 1446 - 0x5a6  :  127 - 0x7f
    "01111111", -- 1447 - 0x5a7  :  127 - 0x7f
    "00000000", -- 1448 - 0x5a8  :    0 - 0x0 -- Sprite 0xb5
    "00000000", -- 1449 - 0x5a9  :    0 - 0x0
    "11111000", -- 1450 - 0x5aa  :  248 - 0xf8
    "11111000", -- 1451 - 0x5ab  :  248 - 0xf8
    "11111000", -- 1452 - 0x5ac  :  248 - 0xf8
    "11111000", -- 1453 - 0x5ad  :  248 - 0xf8
    "11111000", -- 1454 - 0x5ae  :  248 - 0xf8
    "11111000", -- 1455 - 0x5af  :  248 - 0xf8
    "01111111", -- 1456 - 0x5b0  :  127 - 0x7f -- Sprite 0xb6
    "01111111", -- 1457 - 0x5b1  :  127 - 0x7f
    "01111111", -- 1458 - 0x5b2  :  127 - 0x7f
    "01000000", -- 1459 - 0x5b3  :   64 - 0x40
    "00000000", -- 1460 - 0x5b4  :    0 - 0x0
    "00000000", -- 1461 - 0x5b5  :    0 - 0x0
    "00000000", -- 1462 - 0x5b6  :    0 - 0x0
    "00000000", -- 1463 - 0x5b7  :    0 - 0x0
    "11111000", -- 1464 - 0x5b8  :  248 - 0xf8 -- Sprite 0xb7
    "11111000", -- 1465 - 0x5b9  :  248 - 0xf8
    "11111000", -- 1466 - 0x5ba  :  248 - 0xf8
    "00000000", -- 1467 - 0x5bb  :    0 - 0x0
    "00000000", -- 1468 - 0x5bc  :    0 - 0x0
    "00000000", -- 1469 - 0x5bd  :    0 - 0x0
    "00000000", -- 1470 - 0x5be  :    0 - 0x0
    "00000000", -- 1471 - 0x5bf  :    0 - 0x0
    "00000000", -- 1472 - 0x5c0  :    0 - 0x0 -- Sprite 0xb8
    "00000011", -- 1473 - 0x5c1  :    3 - 0x3
    "00000111", -- 1474 - 0x5c2  :    7 - 0x7
    "00000111", -- 1475 - 0x5c3  :    7 - 0x7
    "00000111", -- 1476 - 0x5c4  :    7 - 0x7
    "00000011", -- 1477 - 0x5c5  :    3 - 0x3
    "00000000", -- 1478 - 0x5c6  :    0 - 0x0
    "00000000", -- 1479 - 0x5c7  :    0 - 0x0
    "00000000", -- 1480 - 0x5c8  :    0 - 0x0 -- Sprite 0xb9
    "11000001", -- 1481 - 0x5c9  :  193 - 0xc1
    "11100010", -- 1482 - 0x5ca  :  226 - 0xe2
    "11001100", -- 1483 - 0x5cb  :  204 - 0xcc
    "11000000", -- 1484 - 0x5cc  :  192 - 0xc0
    "10000000", -- 1485 - 0x5cd  :  128 - 0x80
    "00000001", -- 1486 - 0x5ce  :    1 - 0x1
    "00000010", -- 1487 - 0x5cf  :    2 - 0x2
    "11110000", -- 1488 - 0x5d0  :  240 - 0xf0 -- Sprite 0xba
    "00000000", -- 1489 - 0x5d1  :    0 - 0x0
    "00100000", -- 1490 - 0x5d2  :   32 - 0x20
    "00100000", -- 1491 - 0x5d3  :   32 - 0x20
    "00000000", -- 1492 - 0x5d4  :    0 - 0x0
    "11110000", -- 1493 - 0x5d5  :  240 - 0xf0
    "00000000", -- 1494 - 0x5d6  :    0 - 0x0
    "00000000", -- 1495 - 0x5d7  :    0 - 0x0
    "00000000", -- 1496 - 0x5d8  :    0 - 0x0 -- Sprite 0xbb
    "00000000", -- 1497 - 0x5d9  :    0 - 0x0
    "00000000", -- 1498 - 0x5da  :    0 - 0x0
    "00000000", -- 1499 - 0x5db  :    0 - 0x0
    "00000000", -- 1500 - 0x5dc  :    0 - 0x0
    "01100000", -- 1501 - 0x5dd  :   96 - 0x60
    "01100000", -- 1502 - 0x5de  :   96 - 0x60
    "00000000", -- 1503 - 0x5df  :    0 - 0x0
    "00001100", -- 1504 - 0x5e0  :   12 - 0xc -- Sprite 0xbc
    "00000000", -- 1505 - 0x5e1  :    0 - 0x0
    "00000000", -- 1506 - 0x5e2  :    0 - 0x0
    "00000000", -- 1507 - 0x5e3  :    0 - 0x0
    "00000000", -- 1508 - 0x5e4  :    0 - 0x0
    "00000110", -- 1509 - 0x5e5  :    6 - 0x6
    "00000110", -- 1510 - 0x5e6  :    6 - 0x6
    "00000000", -- 1511 - 0x5e7  :    0 - 0x0
    "00000000", -- 1512 - 0x5e8  :    0 - 0x0 -- Sprite 0xbd
    "10000011", -- 1513 - 0x5e9  :  131 - 0x83
    "00000111", -- 1514 - 0x5ea  :    7 - 0x7
    "00000111", -- 1515 - 0x5eb  :    7 - 0x7
    "00000111", -- 1516 - 0x5ec  :    7 - 0x7
    "00000011", -- 1517 - 0x5ed  :    3 - 0x3
    "00000000", -- 1518 - 0x5ee  :    0 - 0x0
    "00000000", -- 1519 - 0x5ef  :    0 - 0x0
    "00000000", -- 1520 - 0x5f0  :    0 - 0x0 -- Sprite 0xbe
    "11000100", -- 1521 - 0x5f1  :  196 - 0xc4
    "11100000", -- 1522 - 0x5f2  :  224 - 0xe0
    "11000000", -- 1523 - 0x5f3  :  192 - 0xc0
    "11000000", -- 1524 - 0x5f4  :  192 - 0xc0
    "10000000", -- 1525 - 0x5f5  :  128 - 0x80
    "00000000", -- 1526 - 0x5f6  :    0 - 0x0
    "00000000", -- 1527 - 0x5f7  :    0 - 0x0
    "00000000", -- 1528 - 0x5f8  :    0 - 0x0 -- Sprite 0xbf
    "00000000", -- 1529 - 0x5f9  :    0 - 0x0
    "00000000", -- 1530 - 0x5fa  :    0 - 0x0
    "00000000", -- 1531 - 0x5fb  :    0 - 0x0
    "00001000", -- 1532 - 0x5fc  :    8 - 0x8
    "10001000", -- 1533 - 0x5fd  :  136 - 0x88
    "00001011", -- 1534 - 0x5fe  :   11 - 0xb
    "00001000", -- 1535 - 0x5ff  :    8 - 0x8
    "00000000", -- 1536 - 0x600  :    0 - 0x0 -- Sprite 0xc0
    "00000000", -- 1537 - 0x601  :    0 - 0x0
    "00000000", -- 1538 - 0x602  :    0 - 0x0
    "00000000", -- 1539 - 0x603  :    0 - 0x0
    "00100000", -- 1540 - 0x604  :   32 - 0x20
    "00100100", -- 1541 - 0x605  :   36 - 0x24
    "10100000", -- 1542 - 0x606  :  160 - 0xa0
    "00100000", -- 1543 - 0x607  :   32 - 0x20
    "00000000", -- 1544 - 0x608  :    0 - 0x0 -- Sprite 0xc1
    "00000000", -- 1545 - 0x609  :    0 - 0x0
    "00000000", -- 1546 - 0x60a  :    0 - 0x0
    "00000000", -- 1547 - 0x60b  :    0 - 0x0
    "00000000", -- 1548 - 0x60c  :    0 - 0x0
    "00000000", -- 1549 - 0x60d  :    0 - 0x0
    "00000000", -- 1550 - 0x60e  :    0 - 0x0
    "00000000", -- 1551 - 0x60f  :    0 - 0x0
    "00000000", -- 1552 - 0x610  :    0 - 0x0 -- Sprite 0xc2
    "00000000", -- 1553 - 0x611  :    0 - 0x0
    "00000000", -- 1554 - 0x612  :    0 - 0x0
    "00000000", -- 1555 - 0x613  :    0 - 0x0
    "00000000", -- 1556 - 0x614  :    0 - 0x0
    "00000000", -- 1557 - 0x615  :    0 - 0x0
    "00000000", -- 1558 - 0x616  :    0 - 0x0
    "00000000", -- 1559 - 0x617  :    0 - 0x0
    "00000000", -- 1560 - 0x618  :    0 - 0x0 -- Sprite 0xc3
    "00000000", -- 1561 - 0x619  :    0 - 0x0
    "00001000", -- 1562 - 0x61a  :    8 - 0x8
    "00001011", -- 1563 - 0x61b  :   11 - 0xb
    "00001000", -- 1564 - 0x61c  :    8 - 0x8
    "00001000", -- 1565 - 0x61d  :    8 - 0x8
    "00001000", -- 1566 - 0x61e  :    8 - 0x8
    "00001000", -- 1567 - 0x61f  :    8 - 0x8
    "00000000", -- 1568 - 0x620  :    0 - 0x0 -- Sprite 0xc4
    "00000000", -- 1569 - 0x621  :    0 - 0x0
    "00100000", -- 1570 - 0x622  :   32 - 0x20
    "10100000", -- 1571 - 0x623  :  160 - 0xa0
    "00100000", -- 1572 - 0x624  :   32 - 0x20
    "00100000", -- 1573 - 0x625  :   32 - 0x20
    "00100000", -- 1574 - 0x626  :   32 - 0x20
    "00100000", -- 1575 - 0x627  :   32 - 0x20
    "00001000", -- 1576 - 0x628  :    8 - 0x8 -- Sprite 0xc5
    "11001000", -- 1577 - 0x629  :  200 - 0xc8
    "00000011", -- 1578 - 0x62a  :    3 - 0x3
    "00000111", -- 1579 - 0x62b  :    7 - 0x7
    "00000111", -- 1580 - 0x62c  :    7 - 0x7
    "00000111", -- 1581 - 0x62d  :    7 - 0x7
    "00000011", -- 1582 - 0x62e  :    3 - 0x3
    "00000000", -- 1583 - 0x62f  :    0 - 0x0
    "00100000", -- 1584 - 0x630  :   32 - 0x20 -- Sprite 0xc6
    "00100110", -- 1585 - 0x631  :   38 - 0x26
    "11000000", -- 1586 - 0x632  :  192 - 0xc0
    "11100000", -- 1587 - 0x633  :  224 - 0xe0
    "11000000", -- 1588 - 0x634  :  192 - 0xc0
    "11000000", -- 1589 - 0x635  :  192 - 0xc0
    "10000000", -- 1590 - 0x636  :  128 - 0x80
    "00000000", -- 1591 - 0x637  :    0 - 0x0
    "00000000", -- 1592 - 0x638  :    0 - 0x0 -- Sprite 0xc7
    "00000000", -- 1593 - 0x639  :    0 - 0x0
    "00000000", -- 1594 - 0x63a  :    0 - 0x0
    "00000000", -- 1595 - 0x63b  :    0 - 0x0
    "00000000", -- 1596 - 0x63c  :    0 - 0x0
    "11000000", -- 1597 - 0x63d  :  192 - 0xc0
    "00000000", -- 1598 - 0x63e  :    0 - 0x0
    "00000000", -- 1599 - 0x63f  :    0 - 0x0
    "00000000", -- 1600 - 0x640  :    0 - 0x0 -- Sprite 0xc8
    "00000000", -- 1601 - 0x641  :    0 - 0x0
    "00000000", -- 1602 - 0x642  :    0 - 0x0
    "00000000", -- 1603 - 0x643  :    0 - 0x0
    "00000000", -- 1604 - 0x644  :    0 - 0x0
    "00000110", -- 1605 - 0x645  :    6 - 0x6
    "00000000", -- 1606 - 0x646  :    0 - 0x0
    "00000000", -- 1607 - 0x647  :    0 - 0x0
    "00001111", -- 1608 - 0x648  :   15 - 0xf -- Sprite 0xc9
    "00000000", -- 1609 - 0x649  :    0 - 0x0
    "00001000", -- 1610 - 0x64a  :    8 - 0x8
    "00001000", -- 1611 - 0x64b  :    8 - 0x8
    "00000000", -- 1612 - 0x64c  :    0 - 0x0
    "00001111", -- 1613 - 0x64d  :   15 - 0xf
    "00000000", -- 1614 - 0x64e  :    0 - 0x0
    "00000000", -- 1615 - 0x64f  :    0 - 0x0
    "00000000", -- 1616 - 0x650  :    0 - 0x0 -- Sprite 0xca
    "10000011", -- 1617 - 0x651  :  131 - 0x83
    "01000111", -- 1618 - 0x652  :   71 - 0x47
    "00110111", -- 1619 - 0x653  :   55 - 0x37
    "00000111", -- 1620 - 0x654  :    7 - 0x7
    "00000011", -- 1621 - 0x655  :    3 - 0x3
    "10000000", -- 1622 - 0x656  :  128 - 0x80
    "01000000", -- 1623 - 0x657  :   64 - 0x40
    "00000000", -- 1624 - 0x658  :    0 - 0x0 -- Sprite 0xcb
    "11000000", -- 1625 - 0x659  :  192 - 0xc0
    "11100000", -- 1626 - 0x65a  :  224 - 0xe0
    "11000000", -- 1627 - 0x65b  :  192 - 0xc0
    "11000000", -- 1628 - 0x65c  :  192 - 0xc0
    "10000000", -- 1629 - 0x65d  :  128 - 0x80
    "00000000", -- 1630 - 0x65e  :    0 - 0x0
    "00000000", -- 1631 - 0x65f  :    0 - 0x0
    "00110000", -- 1632 - 0x660  :   48 - 0x30 -- Sprite 0xcc
    "00000000", -- 1633 - 0x661  :    0 - 0x0
    "00000000", -- 1634 - 0x662  :    0 - 0x0
    "00000000", -- 1635 - 0x663  :    0 - 0x0
    "00000000", -- 1636 - 0x664  :    0 - 0x0
    "01100000", -- 1637 - 0x665  :   96 - 0x60
    "01100000", -- 1638 - 0x666  :   96 - 0x60
    "00000000", -- 1639 - 0x667  :    0 - 0x0
    "00000000", -- 1640 - 0x668  :    0 - 0x0 -- Sprite 0xcd
    "00000000", -- 1641 - 0x669  :    0 - 0x0
    "00000000", -- 1642 - 0x66a  :    0 - 0x0
    "00000000", -- 1643 - 0x66b  :    0 - 0x0
    "00000000", -- 1644 - 0x66c  :    0 - 0x0
    "00000110", -- 1645 - 0x66d  :    6 - 0x6
    "00000110", -- 1646 - 0x66e  :    6 - 0x6
    "00000000", -- 1647 - 0x66f  :    0 - 0x0
    "00000000", -- 1648 - 0x670  :    0 - 0x0 -- Sprite 0xce
    "00000001", -- 1649 - 0x671  :    1 - 0x1
    "00011011", -- 1650 - 0x672  :   27 - 0x1b
    "00010011", -- 1651 - 0x673  :   19 - 0x13
    "00011111", -- 1652 - 0x674  :   31 - 0x1f
    "00111111", -- 1653 - 0x675  :   63 - 0x3f
    "00111111", -- 1654 - 0x676  :   63 - 0x3f
    "00111111", -- 1655 - 0x677  :   63 - 0x3f
    "00000000", -- 1656 - 0x678  :    0 - 0x0 -- Sprite 0xcf
    "11111000", -- 1657 - 0x679  :  248 - 0xf8
    "00001000", -- 1658 - 0x67a  :    8 - 0x8
    "00001000", -- 1659 - 0x67b  :    8 - 0x8
    "00001000", -- 1660 - 0x67c  :    8 - 0x8
    "11111000", -- 1661 - 0x67d  :  248 - 0xf8
    "11110000", -- 1662 - 0x67e  :  240 - 0xf0
    "11010000", -- 1663 - 0x67f  :  208 - 0xd0
    "00000000", -- 1664 - 0x680  :    0 - 0x0 -- Sprite 0xd0
    "00000000", -- 1665 - 0x681  :    0 - 0x0
    "01111100", -- 1666 - 0x682  :  124 - 0x7c
    "11111110", -- 1667 - 0x683  :  254 - 0xfe
    "11101110", -- 1668 - 0x684  :  238 - 0xee
    "11101110", -- 1669 - 0x685  :  238 - 0xee
    "11101110", -- 1670 - 0x686  :  238 - 0xee
    "11101110", -- 1671 - 0x687  :  238 - 0xee
    "00000000", -- 1672 - 0x688  :    0 - 0x0 -- Sprite 0xd1
    "00000000", -- 1673 - 0x689  :    0 - 0x0
    "00111000", -- 1674 - 0x68a  :   56 - 0x38
    "01111000", -- 1675 - 0x68b  :  120 - 0x78
    "01111000", -- 1676 - 0x68c  :  120 - 0x78
    "00111000", -- 1677 - 0x68d  :   56 - 0x38
    "00111000", -- 1678 - 0x68e  :   56 - 0x38
    "00111000", -- 1679 - 0x68f  :   56 - 0x38
    "00000000", -- 1680 - 0x690  :    0 - 0x0 -- Sprite 0xd2
    "00000000", -- 1681 - 0x691  :    0 - 0x0
    "01111100", -- 1682 - 0x692  :  124 - 0x7c
    "11111110", -- 1683 - 0x693  :  254 - 0xfe
    "11101110", -- 1684 - 0x694  :  238 - 0xee
    "00001110", -- 1685 - 0x695  :   14 - 0xe
    "00001110", -- 1686 - 0x696  :   14 - 0xe
    "01111110", -- 1687 - 0x697  :  126 - 0x7e
    "00000000", -- 1688 - 0x698  :    0 - 0x0 -- Sprite 0xd3
    "00000000", -- 1689 - 0x699  :    0 - 0x0
    "01111100", -- 1690 - 0x69a  :  124 - 0x7c
    "11111110", -- 1691 - 0x69b  :  254 - 0xfe
    "11101110", -- 1692 - 0x69c  :  238 - 0xee
    "00001110", -- 1693 - 0x69d  :   14 - 0xe
    "00111100", -- 1694 - 0x69e  :   60 - 0x3c
    "00111100", -- 1695 - 0x69f  :   60 - 0x3c
    "00000000", -- 1696 - 0x6a0  :    0 - 0x0 -- Sprite 0xd4
    "00000000", -- 1697 - 0x6a1  :    0 - 0x0
    "00111110", -- 1698 - 0x6a2  :   62 - 0x3e
    "01111110", -- 1699 - 0x6a3  :  126 - 0x7e
    "11101110", -- 1700 - 0x6a4  :  238 - 0xee
    "11101110", -- 1701 - 0x6a5  :  238 - 0xee
    "11101110", -- 1702 - 0x6a6  :  238 - 0xee
    "11101110", -- 1703 - 0x6a7  :  238 - 0xee
    "00000000", -- 1704 - 0x6a8  :    0 - 0x0 -- Sprite 0xd5
    "00000000", -- 1705 - 0x6a9  :    0 - 0x0
    "11111100", -- 1706 - 0x6aa  :  252 - 0xfc
    "11111100", -- 1707 - 0x6ab  :  252 - 0xfc
    "11100000", -- 1708 - 0x6ac  :  224 - 0xe0
    "11100000", -- 1709 - 0x6ad  :  224 - 0xe0
    "11111100", -- 1710 - 0x6ae  :  252 - 0xfc
    "11111110", -- 1711 - 0x6af  :  254 - 0xfe
    "00000000", -- 1712 - 0x6b0  :    0 - 0x0 -- Sprite 0xd6
    "00000000", -- 1713 - 0x6b1  :    0 - 0x0
    "01111100", -- 1714 - 0x6b2  :  124 - 0x7c
    "11111100", -- 1715 - 0x6b3  :  252 - 0xfc
    "11100000", -- 1716 - 0x6b4  :  224 - 0xe0
    "11100000", -- 1717 - 0x6b5  :  224 - 0xe0
    "11111100", -- 1718 - 0x6b6  :  252 - 0xfc
    "11111110", -- 1719 - 0x6b7  :  254 - 0xfe
    "00000000", -- 1720 - 0x6b8  :    0 - 0x0 -- Sprite 0xd7
    "00000000", -- 1721 - 0x6b9  :    0 - 0x0
    "11111110", -- 1722 - 0x6ba  :  254 - 0xfe
    "11111110", -- 1723 - 0x6bb  :  254 - 0xfe
    "11101110", -- 1724 - 0x6bc  :  238 - 0xee
    "00001110", -- 1725 - 0x6bd  :   14 - 0xe
    "00001110", -- 1726 - 0x6be  :   14 - 0xe
    "00011100", -- 1727 - 0x6bf  :   28 - 0x1c
    "00000000", -- 1728 - 0x6c0  :    0 - 0x0 -- Sprite 0xd8
    "00000000", -- 1729 - 0x6c1  :    0 - 0x0
    "01111100", -- 1730 - 0x6c2  :  124 - 0x7c
    "11111110", -- 1731 - 0x6c3  :  254 - 0xfe
    "11101110", -- 1732 - 0x6c4  :  238 - 0xee
    "11101110", -- 1733 - 0x6c5  :  238 - 0xee
    "01111100", -- 1734 - 0x6c6  :  124 - 0x7c
    "11111110", -- 1735 - 0x6c7  :  254 - 0xfe
    "00000000", -- 1736 - 0x6c8  :    0 - 0x0 -- Sprite 0xd9
    "00000000", -- 1737 - 0x6c9  :    0 - 0x0
    "01111100", -- 1738 - 0x6ca  :  124 - 0x7c
    "11111110", -- 1739 - 0x6cb  :  254 - 0xfe
    "11101110", -- 1740 - 0x6cc  :  238 - 0xee
    "11101110", -- 1741 - 0x6cd  :  238 - 0xee
    "11101110", -- 1742 - 0x6ce  :  238 - 0xee
    "11101110", -- 1743 - 0x6cf  :  238 - 0xee
    "00000000", -- 1744 - 0x6d0  :    0 - 0x0 -- Sprite 0xda
    "00100000", -- 1745 - 0x6d1  :   32 - 0x20
    "00000000", -- 1746 - 0x6d2  :    0 - 0x0
    "00000010", -- 1747 - 0x6d3  :    2 - 0x2
    "00000000", -- 1748 - 0x6d4  :    0 - 0x0
    "00100000", -- 1749 - 0x6d5  :   32 - 0x20
    "00000000", -- 1750 - 0x6d6  :    0 - 0x0
    "00000000", -- 1751 - 0x6d7  :    0 - 0x0
    "00100000", -- 1752 - 0x6d8  :   32 - 0x20 -- Sprite 0xdb
    "00000000", -- 1753 - 0x6d9  :    0 - 0x0
    "00000000", -- 1754 - 0x6da  :    0 - 0x0
    "00000000", -- 1755 - 0x6db  :    0 - 0x0
    "10000000", -- 1756 - 0x6dc  :  128 - 0x80
    "00000000", -- 1757 - 0x6dd  :    0 - 0x0
    "00000100", -- 1758 - 0x6de  :    4 - 0x4
    "00000000", -- 1759 - 0x6df  :    0 - 0x0
    "00000000", -- 1760 - 0x6e0  :    0 - 0x0 -- Sprite 0xdc
    "00001000", -- 1761 - 0x6e1  :    8 - 0x8
    "00000000", -- 1762 - 0x6e2  :    0 - 0x0
    "00000000", -- 1763 - 0x6e3  :    0 - 0x0
    "00000010", -- 1764 - 0x6e4  :    2 - 0x2
    "00000000", -- 1765 - 0x6e5  :    0 - 0x0
    "01000000", -- 1766 - 0x6e6  :   64 - 0x40
    "00000000", -- 1767 - 0x6e7  :    0 - 0x0
    "00000000", -- 1768 - 0x6e8  :    0 - 0x0 -- Sprite 0xdd
    "01000000", -- 1769 - 0x6e9  :   64 - 0x40
    "00000000", -- 1770 - 0x6ea  :    0 - 0x0
    "00000000", -- 1771 - 0x6eb  :    0 - 0x0
    "00000000", -- 1772 - 0x6ec  :    0 - 0x0
    "00000000", -- 1773 - 0x6ed  :    0 - 0x0
    "00000010", -- 1774 - 0x6ee  :    2 - 0x2
    "00100000", -- 1775 - 0x6ef  :   32 - 0x20
    "00111110", -- 1776 - 0x6f0  :   62 - 0x3e -- Sprite 0xde
    "00111111", -- 1777 - 0x6f1  :   63 - 0x3f
    "00111110", -- 1778 - 0x6f2  :   62 - 0x3e
    "00111100", -- 1779 - 0x6f3  :   60 - 0x3c
    "00111111", -- 1780 - 0x6f4  :   63 - 0x3f
    "00110000", -- 1781 - 0x6f5  :   48 - 0x30
    "00000000", -- 1782 - 0x6f6  :    0 - 0x0
    "00000000", -- 1783 - 0x6f7  :    0 - 0x0
    "00010000", -- 1784 - 0x6f8  :   16 - 0x10 -- Sprite 0xdf
    "10110000", -- 1785 - 0x6f9  :  176 - 0xb0
    "00110000", -- 1786 - 0x6fa  :   48 - 0x30
    "11110000", -- 1787 - 0x6fb  :  240 - 0xf0
    "11110000", -- 1788 - 0x6fc  :  240 - 0xf0
    "00000000", -- 1789 - 0x6fd  :    0 - 0x0
    "00000000", -- 1790 - 0x6fe  :    0 - 0x0
    "00000000", -- 1791 - 0x6ff  :    0 - 0x0
    "11101110", -- 1792 - 0x700  :  238 - 0xee -- Sprite 0xe0
    "11101110", -- 1793 - 0x701  :  238 - 0xee
    "11101110", -- 1794 - 0x702  :  238 - 0xee
    "11101110", -- 1795 - 0x703  :  238 - 0xee
    "11111110", -- 1796 - 0x704  :  254 - 0xfe
    "01111100", -- 1797 - 0x705  :  124 - 0x7c
    "00000000", -- 1798 - 0x706  :    0 - 0x0
    "00000000", -- 1799 - 0x707  :    0 - 0x0
    "00111000", -- 1800 - 0x708  :   56 - 0x38 -- Sprite 0xe1
    "00111000", -- 1801 - 0x709  :   56 - 0x38
    "00111000", -- 1802 - 0x70a  :   56 - 0x38
    "00111000", -- 1803 - 0x70b  :   56 - 0x38
    "01111100", -- 1804 - 0x70c  :  124 - 0x7c
    "01111100", -- 1805 - 0x70d  :  124 - 0x7c
    "00000000", -- 1806 - 0x70e  :    0 - 0x0
    "00000000", -- 1807 - 0x70f  :    0 - 0x0
    "11111100", -- 1808 - 0x710  :  252 - 0xfc -- Sprite 0xe2
    "11100000", -- 1809 - 0x711  :  224 - 0xe0
    "11100000", -- 1810 - 0x712  :  224 - 0xe0
    "11100000", -- 1811 - 0x713  :  224 - 0xe0
    "11111110", -- 1812 - 0x714  :  254 - 0xfe
    "11111110", -- 1813 - 0x715  :  254 - 0xfe
    "00000000", -- 1814 - 0x716  :    0 - 0x0
    "00000000", -- 1815 - 0x717  :    0 - 0x0
    "00001110", -- 1816 - 0x718  :   14 - 0xe -- Sprite 0xe3
    "00001110", -- 1817 - 0x719  :   14 - 0xe
    "00001110", -- 1818 - 0x71a  :   14 - 0xe
    "11101110", -- 1819 - 0x71b  :  238 - 0xee
    "11111110", -- 1820 - 0x71c  :  254 - 0xfe
    "01111100", -- 1821 - 0x71d  :  124 - 0x7c
    "00000000", -- 1822 - 0x71e  :    0 - 0x0
    "00000000", -- 1823 - 0x71f  :    0 - 0x0
    "11101110", -- 1824 - 0x720  :  238 - 0xee -- Sprite 0xe4
    "11101110", -- 1825 - 0x721  :  238 - 0xee
    "11111110", -- 1826 - 0x722  :  254 - 0xfe
    "11111110", -- 1827 - 0x723  :  254 - 0xfe
    "00001110", -- 1828 - 0x724  :   14 - 0xe
    "00001110", -- 1829 - 0x725  :   14 - 0xe
    "00000000", -- 1830 - 0x726  :    0 - 0x0
    "00000000", -- 1831 - 0x727  :    0 - 0x0
    "00001110", -- 1832 - 0x728  :   14 - 0xe -- Sprite 0xe5
    "00001110", -- 1833 - 0x729  :   14 - 0xe
    "00001110", -- 1834 - 0x72a  :   14 - 0xe
    "11101110", -- 1835 - 0x72b  :  238 - 0xee
    "11111110", -- 1836 - 0x72c  :  254 - 0xfe
    "01111100", -- 1837 - 0x72d  :  124 - 0x7c
    "00000000", -- 1838 - 0x72e  :    0 - 0x0
    "00000000", -- 1839 - 0x72f  :    0 - 0x0
    "11101110", -- 1840 - 0x730  :  238 - 0xee -- Sprite 0xe6
    "11101110", -- 1841 - 0x731  :  238 - 0xee
    "11101110", -- 1842 - 0x732  :  238 - 0xee
    "11101110", -- 1843 - 0x733  :  238 - 0xee
    "11111110", -- 1844 - 0x734  :  254 - 0xfe
    "01111100", -- 1845 - 0x735  :  124 - 0x7c
    "00000000", -- 1846 - 0x736  :    0 - 0x0
    "00000000", -- 1847 - 0x737  :    0 - 0x0
    "00011100", -- 1848 - 0x738  :   28 - 0x1c -- Sprite 0xe7
    "00011100", -- 1849 - 0x739  :   28 - 0x1c
    "00111000", -- 1850 - 0x73a  :   56 - 0x38
    "00111000", -- 1851 - 0x73b  :   56 - 0x38
    "00111000", -- 1852 - 0x73c  :   56 - 0x38
    "00111000", -- 1853 - 0x73d  :   56 - 0x38
    "00000000", -- 1854 - 0x73e  :    0 - 0x0
    "00000000", -- 1855 - 0x73f  :    0 - 0x0
    "11101110", -- 1856 - 0x740  :  238 - 0xee -- Sprite 0xe8
    "11101110", -- 1857 - 0x741  :  238 - 0xee
    "11101110", -- 1858 - 0x742  :  238 - 0xee
    "11101110", -- 1859 - 0x743  :  238 - 0xee
    "11111110", -- 1860 - 0x744  :  254 - 0xfe
    "01111100", -- 1861 - 0x745  :  124 - 0x7c
    "00000000", -- 1862 - 0x746  :    0 - 0x0
    "00000000", -- 1863 - 0x747  :    0 - 0x0
    "11111110", -- 1864 - 0x748  :  254 - 0xfe -- Sprite 0xe9
    "01111110", -- 1865 - 0x749  :  126 - 0x7e
    "00001110", -- 1866 - 0x74a  :   14 - 0xe
    "00001110", -- 1867 - 0x74b  :   14 - 0xe
    "01111110", -- 1868 - 0x74c  :  126 - 0x7e
    "01111100", -- 1869 - 0x74d  :  124 - 0x7c
    "00000000", -- 1870 - 0x74e  :    0 - 0x0
    "00000000", -- 1871 - 0x74f  :    0 - 0x0
    "00000000", -- 1872 - 0x750  :    0 - 0x0 -- Sprite 0xea
    "01110000", -- 1873 - 0x751  :  112 - 0x70
    "00111000", -- 1874 - 0x752  :   56 - 0x38
    "00000000", -- 1875 - 0x753  :    0 - 0x0
    "00000010", -- 1876 - 0x754  :    2 - 0x2
    "00000111", -- 1877 - 0x755  :    7 - 0x7
    "00000011", -- 1878 - 0x756  :    3 - 0x3
    "00000000", -- 1879 - 0x757  :    0 - 0x0
    "00000000", -- 1880 - 0x758  :    0 - 0x0 -- Sprite 0xeb
    "00001100", -- 1881 - 0x759  :   12 - 0xc
    "00000110", -- 1882 - 0x75a  :    6 - 0x6
    "00000110", -- 1883 - 0x75b  :    6 - 0x6
    "01100000", -- 1884 - 0x75c  :   96 - 0x60
    "01110000", -- 1885 - 0x75d  :  112 - 0x70
    "00110000", -- 1886 - 0x75e  :   48 - 0x30
    "00000000", -- 1887 - 0x75f  :    0 - 0x0
    "00000000", -- 1888 - 0x760  :    0 - 0x0 -- Sprite 0xec
    "11000000", -- 1889 - 0x761  :  192 - 0xc0
    "11100000", -- 1890 - 0x762  :  224 - 0xe0
    "01100000", -- 1891 - 0x763  :   96 - 0x60
    "00000000", -- 1892 - 0x764  :    0 - 0x0
    "00001100", -- 1893 - 0x765  :   12 - 0xc
    "00001110", -- 1894 - 0x766  :   14 - 0xe
    "00000110", -- 1895 - 0x767  :    6 - 0x6
    "01100000", -- 1896 - 0x768  :   96 - 0x60 -- Sprite 0xed
    "01110000", -- 1897 - 0x769  :  112 - 0x70
    "00110000", -- 1898 - 0x76a  :   48 - 0x30
    "00000000", -- 1899 - 0x76b  :    0 - 0x0
    "00000000", -- 1900 - 0x76c  :    0 - 0x0
    "00001100", -- 1901 - 0x76d  :   12 - 0xc
    "00001110", -- 1902 - 0x76e  :   14 - 0xe
    "00000110", -- 1903 - 0x76f  :    6 - 0x6
    "00000000", -- 1904 - 0x770  :    0 - 0x0 -- Sprite 0xee
    "00000000", -- 1905 - 0x771  :    0 - 0x0
    "01000010", -- 1906 - 0x772  :   66 - 0x42
    "00000000", -- 1907 - 0x773  :    0 - 0x0
    "00000000", -- 1908 - 0x774  :    0 - 0x0
    "00000100", -- 1909 - 0x775  :    4 - 0x4
    "00000000", -- 1910 - 0x776  :    0 - 0x0
    "00000000", -- 1911 - 0x777  :    0 - 0x0
    "00000000", -- 1912 - 0x778  :    0 - 0x0 -- Sprite 0xef
    "00000000", -- 1913 - 0x779  :    0 - 0x0
    "00000100", -- 1914 - 0x77a  :    4 - 0x4
    "00000000", -- 1915 - 0x77b  :    0 - 0x0
    "00100000", -- 1916 - 0x77c  :   32 - 0x20
    "00000000", -- 1917 - 0x77d  :    0 - 0x0
    "00000000", -- 1918 - 0x77e  :    0 - 0x0
    "00000000", -- 1919 - 0x77f  :    0 - 0x0
    "00000000", -- 1920 - 0x780  :    0 - 0x0 -- Sprite 0xf0
    "00000000", -- 1921 - 0x781  :    0 - 0x0
    "00000000", -- 1922 - 0x782  :    0 - 0x0
    "00000000", -- 1923 - 0x783  :    0 - 0x0
    "00000000", -- 1924 - 0x784  :    0 - 0x0
    "00000000", -- 1925 - 0x785  :    0 - 0x0
    "00000000", -- 1926 - 0x786  :    0 - 0x0
    "00000000", -- 1927 - 0x787  :    0 - 0x0
    "10000000", -- 1928 - 0x788  :  128 - 0x80 -- Sprite 0xf1
    "10000000", -- 1929 - 0x789  :  128 - 0x80
    "10000000", -- 1930 - 0x78a  :  128 - 0x80
    "10000000", -- 1931 - 0x78b  :  128 - 0x80
    "00000000", -- 1932 - 0x78c  :    0 - 0x0
    "00000000", -- 1933 - 0x78d  :    0 - 0x0
    "00000000", -- 1934 - 0x78e  :    0 - 0x0
    "00000000", -- 1935 - 0x78f  :    0 - 0x0
    "11000000", -- 1936 - 0x790  :  192 - 0xc0 -- Sprite 0xf2
    "11000000", -- 1937 - 0x791  :  192 - 0xc0
    "11000000", -- 1938 - 0x792  :  192 - 0xc0
    "11000000", -- 1939 - 0x793  :  192 - 0xc0
    "00000000", -- 1940 - 0x794  :    0 - 0x0
    "00000000", -- 1941 - 0x795  :    0 - 0x0
    "00000000", -- 1942 - 0x796  :    0 - 0x0
    "00000000", -- 1943 - 0x797  :    0 - 0x0
    "11100000", -- 1944 - 0x798  :  224 - 0xe0 -- Sprite 0xf3
    "11100000", -- 1945 - 0x799  :  224 - 0xe0
    "11100000", -- 1946 - 0x79a  :  224 - 0xe0
    "11100000", -- 1947 - 0x79b  :  224 - 0xe0
    "00000000", -- 1948 - 0x79c  :    0 - 0x0
    "00000000", -- 1949 - 0x79d  :    0 - 0x0
    "00000000", -- 1950 - 0x79e  :    0 - 0x0
    "00000000", -- 1951 - 0x79f  :    0 - 0x0
    "11110000", -- 1952 - 0x7a0  :  240 - 0xf0 -- Sprite 0xf4
    "11110000", -- 1953 - 0x7a1  :  240 - 0xf0
    "11110000", -- 1954 - 0x7a2  :  240 - 0xf0
    "11110000", -- 1955 - 0x7a3  :  240 - 0xf0
    "00000000", -- 1956 - 0x7a4  :    0 - 0x0
    "00000000", -- 1957 - 0x7a5  :    0 - 0x0
    "00000000", -- 1958 - 0x7a6  :    0 - 0x0
    "00000000", -- 1959 - 0x7a7  :    0 - 0x0
    "11111000", -- 1960 - 0x7a8  :  248 - 0xf8 -- Sprite 0xf5
    "11111000", -- 1961 - 0x7a9  :  248 - 0xf8
    "11111000", -- 1962 - 0x7aa  :  248 - 0xf8
    "11111000", -- 1963 - 0x7ab  :  248 - 0xf8
    "00000000", -- 1964 - 0x7ac  :    0 - 0x0
    "00000000", -- 1965 - 0x7ad  :    0 - 0x0
    "00000000", -- 1966 - 0x7ae  :    0 - 0x0
    "00000000", -- 1967 - 0x7af  :    0 - 0x0
    "11111100", -- 1968 - 0x7b0  :  252 - 0xfc -- Sprite 0xf6
    "11111100", -- 1969 - 0x7b1  :  252 - 0xfc
    "11111100", -- 1970 - 0x7b2  :  252 - 0xfc
    "11111100", -- 1971 - 0x7b3  :  252 - 0xfc
    "00000000", -- 1972 - 0x7b4  :    0 - 0x0
    "00000000", -- 1973 - 0x7b5  :    0 - 0x0
    "00000000", -- 1974 - 0x7b6  :    0 - 0x0
    "00000000", -- 1975 - 0x7b7  :    0 - 0x0
    "11111110", -- 1976 - 0x7b8  :  254 - 0xfe -- Sprite 0xf7
    "11111110", -- 1977 - 0x7b9  :  254 - 0xfe
    "11111110", -- 1978 - 0x7ba  :  254 - 0xfe
    "11111110", -- 1979 - 0x7bb  :  254 - 0xfe
    "00000000", -- 1980 - 0x7bc  :    0 - 0x0
    "00000000", -- 1981 - 0x7bd  :    0 - 0x0
    "00000000", -- 1982 - 0x7be  :    0 - 0x0
    "00000000", -- 1983 - 0x7bf  :    0 - 0x0
    "11111111", -- 1984 - 0x7c0  :  255 - 0xff -- Sprite 0xf8
    "11111111", -- 1985 - 0x7c1  :  255 - 0xff
    "11111111", -- 1986 - 0x7c2  :  255 - 0xff
    "11111111", -- 1987 - 0x7c3  :  255 - 0xff
    "00000000", -- 1988 - 0x7c4  :    0 - 0x0
    "00000000", -- 1989 - 0x7c5  :    0 - 0x0
    "00000000", -- 1990 - 0x7c6  :    0 - 0x0
    "00000000", -- 1991 - 0x7c7  :    0 - 0x0
    "00000000", -- 1992 - 0x7c8  :    0 - 0x0 -- Sprite 0xf9
    "00000000", -- 1993 - 0x7c9  :    0 - 0x0
    "00000000", -- 1994 - 0x7ca  :    0 - 0x0
    "00000000", -- 1995 - 0x7cb  :    0 - 0x0
    "01111111", -- 1996 - 0x7cc  :  127 - 0x7f
    "01000000", -- 1997 - 0x7cd  :   64 - 0x40
    "01000000", -- 1998 - 0x7ce  :   64 - 0x40
    "01000000", -- 1999 - 0x7cf  :   64 - 0x40
    "00000000", -- 2000 - 0x7d0  :    0 - 0x0 -- Sprite 0xfa
    "00000000", -- 2001 - 0x7d1  :    0 - 0x0
    "00000000", -- 2002 - 0x7d2  :    0 - 0x0
    "00000000", -- 2003 - 0x7d3  :    0 - 0x0
    "11111111", -- 2004 - 0x7d4  :  255 - 0xff
    "00000000", -- 2005 - 0x7d5  :    0 - 0x0
    "00000000", -- 2006 - 0x7d6  :    0 - 0x0
    "00000000", -- 2007 - 0x7d7  :    0 - 0x0
    "00000000", -- 2008 - 0x7d8  :    0 - 0x0 -- Sprite 0xfb
    "00000000", -- 2009 - 0x7d9  :    0 - 0x0
    "00000000", -- 2010 - 0x7da  :    0 - 0x0
    "00000000", -- 2011 - 0x7db  :    0 - 0x0
    "11111110", -- 2012 - 0x7dc  :  254 - 0xfe
    "00000010", -- 2013 - 0x7dd  :    2 - 0x2
    "00000010", -- 2014 - 0x7de  :    2 - 0x2
    "00000010", -- 2015 - 0x7df  :    2 - 0x2
    "01000000", -- 2016 - 0x7e0  :   64 - 0x40 -- Sprite 0xfc
    "01000000", -- 2017 - 0x7e1  :   64 - 0x40
    "01000000", -- 2018 - 0x7e2  :   64 - 0x40
    "01111111", -- 2019 - 0x7e3  :  127 - 0x7f
    "00000000", -- 2020 - 0x7e4  :    0 - 0x0
    "00000000", -- 2021 - 0x7e5  :    0 - 0x0
    "00000000", -- 2022 - 0x7e6  :    0 - 0x0
    "00000000", -- 2023 - 0x7e7  :    0 - 0x0
    "00000000", -- 2024 - 0x7e8  :    0 - 0x0 -- Sprite 0xfd
    "00000000", -- 2025 - 0x7e9  :    0 - 0x0
    "00000000", -- 2026 - 0x7ea  :    0 - 0x0
    "11111111", -- 2027 - 0x7eb  :  255 - 0xff
    "00000000", -- 2028 - 0x7ec  :    0 - 0x0
    "00000000", -- 2029 - 0x7ed  :    0 - 0x0
    "00000000", -- 2030 - 0x7ee  :    0 - 0x0
    "00000000", -- 2031 - 0x7ef  :    0 - 0x0
    "00000010", -- 2032 - 0x7f0  :    2 - 0x2 -- Sprite 0xfe
    "00000010", -- 2033 - 0x7f1  :    2 - 0x2
    "00000010", -- 2034 - 0x7f2  :    2 - 0x2
    "11111110", -- 2035 - 0x7f3  :  254 - 0xfe
    "00000000", -- 2036 - 0x7f4  :    0 - 0x0
    "00000000", -- 2037 - 0x7f5  :    0 - 0x0
    "00000000", -- 2038 - 0x7f6  :    0 - 0x0
    "00000000", -- 2039 - 0x7f7  :    0 - 0x0
    "00000000", -- 2040 - 0x7f8  :    0 - 0x0 -- Sprite 0xff
    "00000000", -- 2041 - 0x7f9  :    0 - 0x0
    "00000000", -- 2042 - 0x7fa  :    0 - 0x0
    "00000000", -- 2043 - 0x7fb  :    0 - 0x0
    "00000000", -- 2044 - 0x7fc  :    0 - 0x0
    "00000000", -- 2045 - 0x7fd  :    0 - 0x0
    "00000000", -- 2046 - 0x7fe  :    0 - 0x0
    "00000000"  -- 2047 - 0x7ff  :    0 - 0x0
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
