--- Autcmatically generated VHDL ROM from a NES memory file----
---   NAME TABLE
-- https://wiki.nesdev.com/w/index.php/PPU_nametables
--- Only the first Name Table: 1KiB


---  Original memory dump file name: smario_traspas_nt.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_NTABLE_SMARIO_TRASPAS is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(10-1 downto 0);  --1024 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_NTABLE_SMARIO_TRASPAS;

architecture BEHAVIORAL of ROM_NTABLE_SMARIO_TRASPAS is
  signal addr_int  : natural range 0 to 2**10-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
     ------- Name Table 0---------
    "00100100", --    0 -  0x0  :   36 - 0x24 -- line 0x0
    "00100100", --    1 -  0x1  :   36 - 0x24
    "00100100", --    2 -  0x2  :   36 - 0x24
    "00100100", --    3 -  0x3  :   36 - 0x24
    "00100100", --    4 -  0x4  :   36 - 0x24
    "00100100", --    5 -  0x5  :   36 - 0x24
    "00100100", --    6 -  0x6  :   36 - 0x24
    "00100100", --    7 -  0x7  :   36 - 0x24
    "00100100", --    8 -  0x8  :   36 - 0x24
    "00100100", --    9 -  0x9  :   36 - 0x24
    "00100100", --   10 -  0xa  :   36 - 0x24
    "00100100", --   11 -  0xb  :   36 - 0x24
    "00100100", --   12 -  0xc  :   36 - 0x24
    "00100100", --   13 -  0xd  :   36 - 0x24
    "00100100", --   14 -  0xe  :   36 - 0x24
    "00100100", --   15 -  0xf  :   36 - 0x24
    "00100100", --   16 - 0x10  :   36 - 0x24
    "00100100", --   17 - 0x11  :   36 - 0x24
    "00100100", --   18 - 0x12  :   36 - 0x24
    "00100100", --   19 - 0x13  :   36 - 0x24
    "00100100", --   20 - 0x14  :   36 - 0x24
    "00100100", --   21 - 0x15  :   36 - 0x24
    "00100100", --   22 - 0x16  :   36 - 0x24
    "00100100", --   23 - 0x17  :   36 - 0x24
    "00100100", --   24 - 0x18  :   36 - 0x24
    "00100100", --   25 - 0x19  :   36 - 0x24
    "00100100", --   26 - 0x1a  :   36 - 0x24
    "00100100", --   27 - 0x1b  :   36 - 0x24
    "00100100", --   28 - 0x1c  :   36 - 0x24
    "00100100", --   29 - 0x1d  :   36 - 0x24
    "00100100", --   30 - 0x1e  :   36 - 0x24
    "00100100", --   31 - 0x1f  :   36 - 0x24
    "00100100", --   32 - 0x20  :   36 - 0x24 -- line 0x1
    "00100100", --   33 - 0x21  :   36 - 0x24
    "00100100", --   34 - 0x22  :   36 - 0x24
    "00100100", --   35 - 0x23  :   36 - 0x24
    "00100100", --   36 - 0x24  :   36 - 0x24
    "00100100", --   37 - 0x25  :   36 - 0x24
    "00100100", --   38 - 0x26  :   36 - 0x24
    "00100100", --   39 - 0x27  :   36 - 0x24
    "00100100", --   40 - 0x28  :   36 - 0x24
    "00100100", --   41 - 0x29  :   36 - 0x24
    "00100100", --   42 - 0x2a  :   36 - 0x24
    "00100100", --   43 - 0x2b  :   36 - 0x24
    "00100100", --   44 - 0x2c  :   36 - 0x24
    "00100100", --   45 - 0x2d  :   36 - 0x24
    "00100100", --   46 - 0x2e  :   36 - 0x24
    "00100100", --   47 - 0x2f  :   36 - 0x24
    "00100100", --   48 - 0x30  :   36 - 0x24
    "00100100", --   49 - 0x31  :   36 - 0x24
    "00100100", --   50 - 0x32  :   36 - 0x24
    "00100100", --   51 - 0x33  :   36 - 0x24
    "00100100", --   52 - 0x34  :   36 - 0x24
    "00100100", --   53 - 0x35  :   36 - 0x24
    "00100100", --   54 - 0x36  :   36 - 0x24
    "00100100", --   55 - 0x37  :   36 - 0x24
    "00100100", --   56 - 0x38  :   36 - 0x24
    "00100100", --   57 - 0x39  :   36 - 0x24
    "00100100", --   58 - 0x3a  :   36 - 0x24
    "00100100", --   59 - 0x3b  :   36 - 0x24
    "00100100", --   60 - 0x3c  :   36 - 0x24
    "00100100", --   61 - 0x3d  :   36 - 0x24
    "00100100", --   62 - 0x3e  :   36 - 0x24
    "00100100", --   63 - 0x3f  :   36 - 0x24
    "00100100", --   64 - 0x40  :   36 - 0x24 -- line 0x2
    "00100100", --   65 - 0x41  :   36 - 0x24
    "00100100", --   66 - 0x42  :   36 - 0x24
    "00010110", --   67 - 0x43  :   22 - 0x16
    "00001010", --   68 - 0x44  :   10 - 0xa
    "00011011", --   69 - 0x45  :   27 - 0x1b
    "00010010", --   70 - 0x46  :   18 - 0x12
    "00011000", --   71 - 0x47  :   24 - 0x18
    "00100100", --   72 - 0x48  :   36 - 0x24
    "00100100", --   73 - 0x49  :   36 - 0x24
    "00100100", --   74 - 0x4a  :   36 - 0x24
    "00100100", --   75 - 0x4b  :   36 - 0x24
    "00100100", --   76 - 0x4c  :   36 - 0x24
    "00100100", --   77 - 0x4d  :   36 - 0x24
    "00100100", --   78 - 0x4e  :   36 - 0x24
    "00100100", --   79 - 0x4f  :   36 - 0x24
    "00100100", --   80 - 0x50  :   36 - 0x24
    "00100100", --   81 - 0x51  :   36 - 0x24
    "00100000", --   82 - 0x52  :   32 - 0x20
    "00011000", --   83 - 0x53  :   24 - 0x18
    "00011011", --   84 - 0x54  :   27 - 0x1b
    "00010101", --   85 - 0x55  :   21 - 0x15
    "00001101", --   86 - 0x56  :   13 - 0xd
    "00100100", --   87 - 0x57  :   36 - 0x24
    "00100100", --   88 - 0x58  :   36 - 0x24
    "00011101", --   89 - 0x59  :   29 - 0x1d
    "00010010", --   90 - 0x5a  :   18 - 0x12
    "00010110", --   91 - 0x5b  :   22 - 0x16
    "00001110", --   92 - 0x5c  :   14 - 0xe
    "00100100", --   93 - 0x5d  :   36 - 0x24
    "00100100", --   94 - 0x5e  :   36 - 0x24
    "00100100", --   95 - 0x5f  :   36 - 0x24
    "00100100", --   96 - 0x60  :   36 - 0x24 -- line 0x3
    "00100100", --   97 - 0x61  :   36 - 0x24
    "00100100", --   98 - 0x62  :   36 - 0x24
    "00000000", --   99 - 0x63  :    0 - 0x0
    "00000000", --  100 - 0x64  :    0 - 0x0
    "00000001", --  101 - 0x65  :    1 - 0x1
    "00000111", --  102 - 0x66  :    7 - 0x7
    "00000000", --  103 - 0x67  :    0 - 0x0
    "00000000", --  104 - 0x68  :    0 - 0x0
    "00100100", --  105 - 0x69  :   36 - 0x24
    "00100100", --  106 - 0x6a  :   36 - 0x24
    "00101110", --  107 - 0x6b  :   46 - 0x2e
    "00101001", --  108 - 0x6c  :   41 - 0x29
    "00000000", --  109 - 0x6d  :    0 - 0x0
    "00000000", --  110 - 0x6e  :    0 - 0x0
    "00100100", --  111 - 0x6f  :   36 - 0x24
    "00100100", --  112 - 0x70  :   36 - 0x24
    "00100100", --  113 - 0x71  :   36 - 0x24
    "00100100", --  114 - 0x72  :   36 - 0x24
    "00000001", --  115 - 0x73  :    1 - 0x1
    "00101000", --  116 - 0x74  :   40 - 0x28
    "00000001", --  117 - 0x75  :    1 - 0x1
    "00100100", --  118 - 0x76  :   36 - 0x24
    "00100100", --  119 - 0x77  :   36 - 0x24
    "00100100", --  120 - 0x78  :   36 - 0x24
    "00100100", --  121 - 0x79  :   36 - 0x24
    "00000011", --  122 - 0x7a  :    3 - 0x3
    "00000010", --  123 - 0x7b  :    2 - 0x2
    "00000011", --  124 - 0x7c  :    3 - 0x3
    "00100100", --  125 - 0x7d  :   36 - 0x24
    "00100100", --  126 - 0x7e  :   36 - 0x24
    "00100100", --  127 - 0x7f  :   36 - 0x24
    "00100100", --  128 - 0x80  :   36 - 0x24 -- line 0x4
    "00100100", --  129 - 0x81  :   36 - 0x24
    "00100100", --  130 - 0x82  :   36 - 0x24
    "00100100", --  131 - 0x83  :   36 - 0x24
    "00100100", --  132 - 0x84  :   36 - 0x24
    "00100100", --  133 - 0x85  :   36 - 0x24
    "00100100", --  134 - 0x86  :   36 - 0x24
    "00100100", --  135 - 0x87  :   36 - 0x24
    "00100100", --  136 - 0x88  :   36 - 0x24
    "00100100", --  137 - 0x89  :   36 - 0x24
    "00100100", --  138 - 0x8a  :   36 - 0x24
    "00100100", --  139 - 0x8b  :   36 - 0x24
    "00100100", --  140 - 0x8c  :   36 - 0x24
    "00100100", --  141 - 0x8d  :   36 - 0x24
    "00100100", --  142 - 0x8e  :   36 - 0x24
    "00100100", --  143 - 0x8f  :   36 - 0x24
    "00100100", --  144 - 0x90  :   36 - 0x24
    "00100100", --  145 - 0x91  :   36 - 0x24
    "00100100", --  146 - 0x92  :   36 - 0x24
    "00100100", --  147 - 0x93  :   36 - 0x24
    "00100100", --  148 - 0x94  :   36 - 0x24
    "00100100", --  149 - 0x95  :   36 - 0x24
    "00100100", --  150 - 0x96  :   36 - 0x24
    "00100100", --  151 - 0x97  :   36 - 0x24
    "00100100", --  152 - 0x98  :   36 - 0x24
    "00100100", --  153 - 0x99  :   36 - 0x24
    "00100100", --  154 - 0x9a  :   36 - 0x24
    "00100100", --  155 - 0x9b  :   36 - 0x24
    "00100100", --  156 - 0x9c  :   36 - 0x24
    "00100100", --  157 - 0x9d  :   36 - 0x24
    "00100100", --  158 - 0x9e  :   36 - 0x24
    "00100100", --  159 - 0x9f  :   36 - 0x24
    "00100100", --  160 - 0xa0  :   36 - 0x24 -- line 0x5
    "00100100", --  161 - 0xa1  :   36 - 0x24
    "00100100", --  162 - 0xa2  :   36 - 0x24
    "00100100", --  163 - 0xa3  :   36 - 0x24
    "00100100", --  164 - 0xa4  :   36 - 0x24
    "00100100", --  165 - 0xa5  :   36 - 0x24
    "00100100", --  166 - 0xa6  :   36 - 0x24
    "00100100", --  167 - 0xa7  :   36 - 0x24
    "00100100", --  168 - 0xa8  :   36 - 0x24
    "00100100", --  169 - 0xa9  :   36 - 0x24
    "00100100", --  170 - 0xaa  :   36 - 0x24
    "00100100", --  171 - 0xab  :   36 - 0x24
    "00100100", --  172 - 0xac  :   36 - 0x24
    "00100100", --  173 - 0xad  :   36 - 0x24
    "00100100", --  174 - 0xae  :   36 - 0x24
    "00100100", --  175 - 0xaf  :   36 - 0x24
    "00100100", --  176 - 0xb0  :   36 - 0x24
    "00100100", --  177 - 0xb1  :   36 - 0x24
    "00100100", --  178 - 0xb2  :   36 - 0x24
    "00100100", --  179 - 0xb3  :   36 - 0x24
    "00100100", --  180 - 0xb4  :   36 - 0x24
    "00100100", --  181 - 0xb5  :   36 - 0x24
    "00100100", --  182 - 0xb6  :   36 - 0x24
    "00100100", --  183 - 0xb7  :   36 - 0x24
    "00100100", --  184 - 0xb8  :   36 - 0x24
    "00100100", --  185 - 0xb9  :   36 - 0x24
    "00100100", --  186 - 0xba  :   36 - 0x24
    "00100100", --  187 - 0xbb  :   36 - 0x24
    "00100100", --  188 - 0xbc  :   36 - 0x24
    "00100100", --  189 - 0xbd  :   36 - 0x24
    "00100100", --  190 - 0xbe  :   36 - 0x24
    "00100100", --  191 - 0xbf  :   36 - 0x24
    "00100100", --  192 - 0xc0  :   36 - 0x24 -- line 0x6
    "00100100", --  193 - 0xc1  :   36 - 0x24
    "00100100", --  194 - 0xc2  :   36 - 0x24
    "00100100", --  195 - 0xc3  :   36 - 0x24
    "00100100", --  196 - 0xc4  :   36 - 0x24
    "00100100", --  197 - 0xc5  :   36 - 0x24
    "00100100", --  198 - 0xc6  :   36 - 0x24
    "00100100", --  199 - 0xc7  :   36 - 0x24
    "00100100", --  200 - 0xc8  :   36 - 0x24
    "00100100", --  201 - 0xc9  :   36 - 0x24
    "00100100", --  202 - 0xca  :   36 - 0x24
    "00100100", --  203 - 0xcb  :   36 - 0x24
    "00100100", --  204 - 0xcc  :   36 - 0x24
    "00100100", --  205 - 0xcd  :   36 - 0x24
    "00100100", --  206 - 0xce  :   36 - 0x24
    "00100100", --  207 - 0xcf  :   36 - 0x24
    "00100100", --  208 - 0xd0  :   36 - 0x24
    "00100100", --  209 - 0xd1  :   36 - 0x24
    "00110110", --  210 - 0xd2  :   54 - 0x36
    "00110111", --  211 - 0xd3  :   55 - 0x37
    "00100100", --  212 - 0xd4  :   36 - 0x24
    "00100100", --  213 - 0xd5  :   36 - 0x24
    "00100100", --  214 - 0xd6  :   36 - 0x24
    "00100100", --  215 - 0xd7  :   36 - 0x24
    "00100100", --  216 - 0xd8  :   36 - 0x24
    "00100100", --  217 - 0xd9  :   36 - 0x24
    "00100100", --  218 - 0xda  :   36 - 0x24
    "00100100", --  219 - 0xdb  :   36 - 0x24
    "00100100", --  220 - 0xdc  :   36 - 0x24
    "00100100", --  221 - 0xdd  :   36 - 0x24
    "00100100", --  222 - 0xde  :   36 - 0x24
    "00100100", --  223 - 0xdf  :   36 - 0x24
    "00100100", --  224 - 0xe0  :   36 - 0x24 -- line 0x7
    "00100100", --  225 - 0xe1  :   36 - 0x24
    "00100100", --  226 - 0xe2  :   36 - 0x24
    "00100100", --  227 - 0xe3  :   36 - 0x24
    "00100100", --  228 - 0xe4  :   36 - 0x24
    "00100100", --  229 - 0xe5  :   36 - 0x24
    "00100100", --  230 - 0xe6  :   36 - 0x24
    "00100100", --  231 - 0xe7  :   36 - 0x24
    "00100100", --  232 - 0xe8  :   36 - 0x24
    "00100100", --  233 - 0xe9  :   36 - 0x24
    "00100100", --  234 - 0xea  :   36 - 0x24
    "00100100", --  235 - 0xeb  :   36 - 0x24
    "00100100", --  236 - 0xec  :   36 - 0x24
    "00100100", --  237 - 0xed  :   36 - 0x24
    "00100100", --  238 - 0xee  :   36 - 0x24
    "00100100", --  239 - 0xef  :   36 - 0x24
    "00100100", --  240 - 0xf0  :   36 - 0x24
    "00110101", --  241 - 0xf1  :   53 - 0x35
    "00100101", --  242 - 0xf2  :   37 - 0x25
    "00100101", --  243 - 0xf3  :   37 - 0x25
    "00111000", --  244 - 0xf4  :   56 - 0x38
    "00100100", --  245 - 0xf5  :   36 - 0x24
    "00100100", --  246 - 0xf6  :   36 - 0x24
    "00100100", --  247 - 0xf7  :   36 - 0x24
    "00100100", --  248 - 0xf8  :   36 - 0x24
    "00100100", --  249 - 0xf9  :   36 - 0x24
    "00100100", --  250 - 0xfa  :   36 - 0x24
    "00100100", --  251 - 0xfb  :   36 - 0x24
    "00100100", --  252 - 0xfc  :   36 - 0x24
    "00100100", --  253 - 0xfd  :   36 - 0x24
    "00100100", --  254 - 0xfe  :   36 - 0x24
    "00100100", --  255 - 0xff  :   36 - 0x24
    "00100100", --  256 - 0x100  :   36 - 0x24 -- line 0x8
    "00100100", --  257 - 0x101  :   36 - 0x24
    "00100100", --  258 - 0x102  :   36 - 0x24
    "00100100", --  259 - 0x103  :   36 - 0x24
    "00100100", --  260 - 0x104  :   36 - 0x24
    "00100100", --  261 - 0x105  :   36 - 0x24
    "00100100", --  262 - 0x106  :   36 - 0x24
    "00100100", --  263 - 0x107  :   36 - 0x24
    "00100100", --  264 - 0x108  :   36 - 0x24
    "00100100", --  265 - 0x109  :   36 - 0x24
    "00100100", --  266 - 0x10a  :   36 - 0x24
    "00100100", --  267 - 0x10b  :   36 - 0x24
    "00100100", --  268 - 0x10c  :   36 - 0x24
    "00100100", --  269 - 0x10d  :   36 - 0x24
    "00100100", --  270 - 0x10e  :   36 - 0x24
    "00100100", --  271 - 0x10f  :   36 - 0x24
    "00100100", --  272 - 0x110  :   36 - 0x24
    "00111001", --  273 - 0x111  :   57 - 0x39
    "00111010", --  274 - 0x112  :   58 - 0x3a
    "00111011", --  275 - 0x113  :   59 - 0x3b
    "00111100", --  276 - 0x114  :   60 - 0x3c
    "00100100", --  277 - 0x115  :   36 - 0x24
    "00100100", --  278 - 0x116  :   36 - 0x24
    "00100100", --  279 - 0x117  :   36 - 0x24
    "00100100", --  280 - 0x118  :   36 - 0x24
    "00100100", --  281 - 0x119  :   36 - 0x24
    "00100100", --  282 - 0x11a  :   36 - 0x24
    "00100100", --  283 - 0x11b  :   36 - 0x24
    "00100100", --  284 - 0x11c  :   36 - 0x24
    "00100100", --  285 - 0x11d  :   36 - 0x24
    "00100100", --  286 - 0x11e  :   36 - 0x24
    "00100100", --  287 - 0x11f  :   36 - 0x24
    "00100100", --  288 - 0x120  :   36 - 0x24 -- line 0x9
    "00100100", --  289 - 0x121  :   36 - 0x24
    "00100100", --  290 - 0x122  :   36 - 0x24
    "00100100", --  291 - 0x123  :   36 - 0x24
    "00100100", --  292 - 0x124  :   36 - 0x24
    "00100100", --  293 - 0x125  :   36 - 0x24
    "00100100", --  294 - 0x126  :   36 - 0x24
    "00100100", --  295 - 0x127  :   36 - 0x24
    "00100100", --  296 - 0x128  :   36 - 0x24
    "00100100", --  297 - 0x129  :   36 - 0x24
    "00100100", --  298 - 0x12a  :   36 - 0x24
    "00100100", --  299 - 0x12b  :   36 - 0x24
    "00100100", --  300 - 0x12c  :   36 - 0x24
    "00100100", --  301 - 0x12d  :   36 - 0x24
    "00100100", --  302 - 0x12e  :   36 - 0x24
    "00100100", --  303 - 0x12f  :   36 - 0x24
    "00100100", --  304 - 0x130  :   36 - 0x24
    "00100100", --  305 - 0x131  :   36 - 0x24
    "00100100", --  306 - 0x132  :   36 - 0x24
    "00100100", --  307 - 0x133  :   36 - 0x24
    "00100100", --  308 - 0x134  :   36 - 0x24
    "00100100", --  309 - 0x135  :   36 - 0x24
    "00100100", --  310 - 0x136  :   36 - 0x24
    "00100100", --  311 - 0x137  :   36 - 0x24
    "00100100", --  312 - 0x138  :   36 - 0x24
    "00100100", --  313 - 0x139  :   36 - 0x24
    "00100100", --  314 - 0x13a  :   36 - 0x24
    "00100100", --  315 - 0x13b  :   36 - 0x24
    "00100100", --  316 - 0x13c  :   36 - 0x24
    "00100100", --  317 - 0x13d  :   36 - 0x24
    "00100100", --  318 - 0x13e  :   36 - 0x24
    "00100100", --  319 - 0x13f  :   36 - 0x24
    "00100100", --  320 - 0x140  :   36 - 0x24 -- line 0xa
    "00100100", --  321 - 0x141  :   36 - 0x24
    "00100100", --  322 - 0x142  :   36 - 0x24
    "00100100", --  323 - 0x143  :   36 - 0x24
    "00100100", --  324 - 0x144  :   36 - 0x24
    "00100100", --  325 - 0x145  :   36 - 0x24
    "00100100", --  326 - 0x146  :   36 - 0x24
    "00100100", --  327 - 0x147  :   36 - 0x24
    "00100100", --  328 - 0x148  :   36 - 0x24
    "00100100", --  329 - 0x149  :   36 - 0x24
    "00100100", --  330 - 0x14a  :   36 - 0x24
    "00100100", --  331 - 0x14b  :   36 - 0x24
    "00100100", --  332 - 0x14c  :   36 - 0x24
    "00100100", --  333 - 0x14d  :   36 - 0x24
    "00100100", --  334 - 0x14e  :   36 - 0x24
    "00100100", --  335 - 0x14f  :   36 - 0x24
    "00100100", --  336 - 0x150  :   36 - 0x24
    "00100100", --  337 - 0x151  :   36 - 0x24
    "00100100", --  338 - 0x152  :   36 - 0x24
    "00100100", --  339 - 0x153  :   36 - 0x24
    "00100100", --  340 - 0x154  :   36 - 0x24
    "00100100", --  341 - 0x155  :   36 - 0x24
    "00100100", --  342 - 0x156  :   36 - 0x24
    "00100100", --  343 - 0x157  :   36 - 0x24
    "00100100", --  344 - 0x158  :   36 - 0x24
    "00100100", --  345 - 0x159  :   36 - 0x24
    "01010011", --  346 - 0x15a  :   83 - 0x53
    "01010100", --  347 - 0x15b  :   84 - 0x54
    "00100100", --  348 - 0x15c  :   36 - 0x24
    "00100100", --  349 - 0x15d  :   36 - 0x24
    "00100100", --  350 - 0x15e  :   36 - 0x24
    "00100100", --  351 - 0x15f  :   36 - 0x24
    "00100100", --  352 - 0x160  :   36 - 0x24 -- line 0xb
    "00100100", --  353 - 0x161  :   36 - 0x24
    "00100100", --  354 - 0x162  :   36 - 0x24
    "00100100", --  355 - 0x163  :   36 - 0x24
    "00100100", --  356 - 0x164  :   36 - 0x24
    "00100100", --  357 - 0x165  :   36 - 0x24
    "00100100", --  358 - 0x166  :   36 - 0x24
    "00100100", --  359 - 0x167  :   36 - 0x24
    "00100100", --  360 - 0x168  :   36 - 0x24
    "00100100", --  361 - 0x169  :   36 - 0x24
    "00100100", --  362 - 0x16a  :   36 - 0x24
    "00100100", --  363 - 0x16b  :   36 - 0x24
    "00100100", --  364 - 0x16c  :   36 - 0x24
    "00100100", --  365 - 0x16d  :   36 - 0x24
    "00100100", --  366 - 0x16e  :   36 - 0x24
    "00100100", --  367 - 0x16f  :   36 - 0x24
    "00100100", --  368 - 0x170  :   36 - 0x24
    "00100100", --  369 - 0x171  :   36 - 0x24
    "00100100", --  370 - 0x172  :   36 - 0x24
    "00100100", --  371 - 0x173  :   36 - 0x24
    "00100100", --  372 - 0x174  :   36 - 0x24
    "00100100", --  373 - 0x175  :   36 - 0x24
    "00100100", --  374 - 0x176  :   36 - 0x24
    "00100100", --  375 - 0x177  :   36 - 0x24
    "00100100", --  376 - 0x178  :   36 - 0x24
    "00100100", --  377 - 0x179  :   36 - 0x24
    "01010101", --  378 - 0x17a  :   85 - 0x55
    "01010110", --  379 - 0x17b  :   86 - 0x56
    "00100100", --  380 - 0x17c  :   36 - 0x24
    "00100100", --  381 - 0x17d  :   36 - 0x24
    "00100100", --  382 - 0x17e  :   36 - 0x24
    "00100100", --  383 - 0x17f  :   36 - 0x24
    "00100100", --  384 - 0x180  :   36 - 0x24 -- line 0xc
    "00100100", --  385 - 0x181  :   36 - 0x24
    "00100100", --  386 - 0x182  :   36 - 0x24
    "00100100", --  387 - 0x183  :   36 - 0x24
    "00100100", --  388 - 0x184  :   36 - 0x24
    "00100100", --  389 - 0x185  :   36 - 0x24
    "00100100", --  390 - 0x186  :   36 - 0x24
    "00100100", --  391 - 0x187  :   36 - 0x24
    "00100100", --  392 - 0x188  :   36 - 0x24
    "00100100", --  393 - 0x189  :   36 - 0x24
    "00100100", --  394 - 0x18a  :   36 - 0x24
    "00100100", --  395 - 0x18b  :   36 - 0x24
    "00100100", --  396 - 0x18c  :   36 - 0x24
    "00100100", --  397 - 0x18d  :   36 - 0x24
    "00100100", --  398 - 0x18e  :   36 - 0x24
    "00100100", --  399 - 0x18f  :   36 - 0x24
    "00100100", --  400 - 0x190  :   36 - 0x24
    "00100100", --  401 - 0x191  :   36 - 0x24
    "00100100", --  402 - 0x192  :   36 - 0x24
    "00100100", --  403 - 0x193  :   36 - 0x24
    "00100100", --  404 - 0x194  :   36 - 0x24
    "00100100", --  405 - 0x195  :   36 - 0x24
    "00100100", --  406 - 0x196  :   36 - 0x24
    "00100100", --  407 - 0x197  :   36 - 0x24
    "00100100", --  408 - 0x198  :   36 - 0x24
    "00100100", --  409 - 0x199  :   36 - 0x24
    "00100100", --  410 - 0x19a  :   36 - 0x24
    "00100100", --  411 - 0x19b  :   36 - 0x24
    "00100100", --  412 - 0x19c  :   36 - 0x24
    "00100100", --  413 - 0x19d  :   36 - 0x24
    "00100100", --  414 - 0x19e  :   36 - 0x24
    "00100100", --  415 - 0x19f  :   36 - 0x24
    "00100100", --  416 - 0x1a0  :   36 - 0x24 -- line 0xd
    "00100100", --  417 - 0x1a1  :   36 - 0x24
    "00100100", --  418 - 0x1a2  :   36 - 0x24
    "00100100", --  419 - 0x1a3  :   36 - 0x24
    "00100100", --  420 - 0x1a4  :   36 - 0x24
    "00100100", --  421 - 0x1a5  :   36 - 0x24
    "00100100", --  422 - 0x1a6  :   36 - 0x24
    "00100100", --  423 - 0x1a7  :   36 - 0x24
    "00100100", --  424 - 0x1a8  :   36 - 0x24
    "00100100", --  425 - 0x1a9  :   36 - 0x24
    "00100100", --  426 - 0x1aa  :   36 - 0x24
    "00100100", --  427 - 0x1ab  :   36 - 0x24
    "00100100", --  428 - 0x1ac  :   36 - 0x24
    "00100100", --  429 - 0x1ad  :   36 - 0x24
    "00100100", --  430 - 0x1ae  :   36 - 0x24
    "00100100", --  431 - 0x1af  :   36 - 0x24
    "00100100", --  432 - 0x1b0  :   36 - 0x24
    "00100100", --  433 - 0x1b1  :   36 - 0x24
    "00100100", --  434 - 0x1b2  :   36 - 0x24
    "00100100", --  435 - 0x1b3  :   36 - 0x24
    "00100100", --  436 - 0x1b4  :   36 - 0x24
    "00100100", --  437 - 0x1b5  :   36 - 0x24
    "00100100", --  438 - 0x1b6  :   36 - 0x24
    "00100100", --  439 - 0x1b7  :   36 - 0x24
    "00100100", --  440 - 0x1b8  :   36 - 0x24
    "00100100", --  441 - 0x1b9  :   36 - 0x24
    "00100100", --  442 - 0x1ba  :   36 - 0x24
    "00100100", --  443 - 0x1bb  :   36 - 0x24
    "00100100", --  444 - 0x1bc  :   36 - 0x24
    "00100100", --  445 - 0x1bd  :   36 - 0x24
    "00100100", --  446 - 0x1be  :   36 - 0x24
    "00100100", --  447 - 0x1bf  :   36 - 0x24
    "00100100", --  448 - 0x1c0  :   36 - 0x24 -- line 0xe
    "00100100", --  449 - 0x1c1  :   36 - 0x24
    "00100100", --  450 - 0x1c2  :   36 - 0x24
    "00100100", --  451 - 0x1c3  :   36 - 0x24
    "00100100", --  452 - 0x1c4  :   36 - 0x24
    "00100100", --  453 - 0x1c5  :   36 - 0x24
    "00100100", --  454 - 0x1c6  :   36 - 0x24
    "00100100", --  455 - 0x1c7  :   36 - 0x24
    "00100100", --  456 - 0x1c8  :   36 - 0x24
    "00100100", --  457 - 0x1c9  :   36 - 0x24
    "00100100", --  458 - 0x1ca  :   36 - 0x24
    "00100100", --  459 - 0x1cb  :   36 - 0x24
    "00100100", --  460 - 0x1cc  :   36 - 0x24
    "00100100", --  461 - 0x1cd  :   36 - 0x24
    "00100100", --  462 - 0x1ce  :   36 - 0x24
    "00100100", --  463 - 0x1cf  :   36 - 0x24
    "00100100", --  464 - 0x1d0  :   36 - 0x24
    "00100100", --  465 - 0x1d1  :   36 - 0x24
    "00100100", --  466 - 0x1d2  :   36 - 0x24
    "00100100", --  467 - 0x1d3  :   36 - 0x24
    "00100100", --  468 - 0x1d4  :   36 - 0x24
    "00100100", --  469 - 0x1d5  :   36 - 0x24
    "00100100", --  470 - 0x1d6  :   36 - 0x24
    "00100100", --  471 - 0x1d7  :   36 - 0x24
    "00100100", --  472 - 0x1d8  :   36 - 0x24
    "00100100", --  473 - 0x1d9  :   36 - 0x24
    "00100100", --  474 - 0x1da  :   36 - 0x24
    "00100100", --  475 - 0x1db  :   36 - 0x24
    "00100100", --  476 - 0x1dc  :   36 - 0x24
    "00100100", --  477 - 0x1dd  :   36 - 0x24
    "00100100", --  478 - 0x1de  :   36 - 0x24
    "00100100", --  479 - 0x1df  :   36 - 0x24
    "00100100", --  480 - 0x1e0  :   36 - 0x24 -- line 0xf
    "00100100", --  481 - 0x1e1  :   36 - 0x24
    "00100100", --  482 - 0x1e2  :   36 - 0x24
    "00100100", --  483 - 0x1e3  :   36 - 0x24
    "00100100", --  484 - 0x1e4  :   36 - 0x24
    "00100100", --  485 - 0x1e5  :   36 - 0x24
    "00100100", --  486 - 0x1e6  :   36 - 0x24
    "00100100", --  487 - 0x1e7  :   36 - 0x24
    "00100100", --  488 - 0x1e8  :   36 - 0x24
    "00100100", --  489 - 0x1e9  :   36 - 0x24
    "00100100", --  490 - 0x1ea  :   36 - 0x24
    "00100100", --  491 - 0x1eb  :   36 - 0x24
    "00100100", --  492 - 0x1ec  :   36 - 0x24
    "00100100", --  493 - 0x1ed  :   36 - 0x24
    "00100100", --  494 - 0x1ee  :   36 - 0x24
    "00100100", --  495 - 0x1ef  :   36 - 0x24
    "00100100", --  496 - 0x1f0  :   36 - 0x24
    "00100100", --  497 - 0x1f1  :   36 - 0x24
    "00100100", --  498 - 0x1f2  :   36 - 0x24
    "00100100", --  499 - 0x1f3  :   36 - 0x24
    "00100100", --  500 - 0x1f4  :   36 - 0x24
    "00100100", --  501 - 0x1f5  :   36 - 0x24
    "00100100", --  502 - 0x1f6  :   36 - 0x24
    "00100100", --  503 - 0x1f7  :   36 - 0x24
    "00100100", --  504 - 0x1f8  :   36 - 0x24
    "00100100", --  505 - 0x1f9  :   36 - 0x24
    "00100100", --  506 - 0x1fa  :   36 - 0x24
    "00100100", --  507 - 0x1fb  :   36 - 0x24
    "00100100", --  508 - 0x1fc  :   36 - 0x24
    "00100100", --  509 - 0x1fd  :   36 - 0x24
    "00100100", --  510 - 0x1fe  :   36 - 0x24
    "00100100", --  511 - 0x1ff  :   36 - 0x24
    "00100100", --  512 - 0x200  :   36 - 0x24 -- line 0x10
    "00100100", --  513 - 0x201  :   36 - 0x24
    "00100100", --  514 - 0x202  :   36 - 0x24
    "00100100", --  515 - 0x203  :   36 - 0x24
    "00100100", --  516 - 0x204  :   36 - 0x24
    "00100100", --  517 - 0x205  :   36 - 0x24
    "00100100", --  518 - 0x206  :   36 - 0x24
    "00100100", --  519 - 0x207  :   36 - 0x24
    "00100100", --  520 - 0x208  :   36 - 0x24
    "00100100", --  521 - 0x209  :   36 - 0x24
    "00100100", --  522 - 0x20a  :   36 - 0x24
    "00100100", --  523 - 0x20b  :   36 - 0x24
    "00100100", --  524 - 0x20c  :   36 - 0x24
    "00100100", --  525 - 0x20d  :   36 - 0x24
    "00100100", --  526 - 0x20e  :   36 - 0x24
    "00100100", --  527 - 0x20f  :   36 - 0x24
    "00100100", --  528 - 0x210  :   36 - 0x24
    "00100100", --  529 - 0x211  :   36 - 0x24
    "00100100", --  530 - 0x212  :   36 - 0x24
    "00100100", --  531 - 0x213  :   36 - 0x24
    "00100100", --  532 - 0x214  :   36 - 0x24
    "00100100", --  533 - 0x215  :   36 - 0x24
    "00100100", --  534 - 0x216  :   36 - 0x24
    "00100100", --  535 - 0x217  :   36 - 0x24
    "00100100", --  536 - 0x218  :   36 - 0x24
    "00100100", --  537 - 0x219  :   36 - 0x24
    "00100100", --  538 - 0x21a  :   36 - 0x24
    "00100100", --  539 - 0x21b  :   36 - 0x24
    "00100100", --  540 - 0x21c  :   36 - 0x24
    "00100100", --  541 - 0x21d  :   36 - 0x24
    "00100100", --  542 - 0x21e  :   36 - 0x24
    "00100100", --  543 - 0x21f  :   36 - 0x24
    "00100100", --  544 - 0x220  :   36 - 0x24 -- line 0x11
    "00100100", --  545 - 0x221  :   36 - 0x24
    "00100100", --  546 - 0x222  :   36 - 0x24
    "00100100", --  547 - 0x223  :   36 - 0x24
    "00100100", --  548 - 0x224  :   36 - 0x24
    "00100100", --  549 - 0x225  :   36 - 0x24
    "00100100", --  550 - 0x226  :   36 - 0x24
    "00100100", --  551 - 0x227  :   36 - 0x24
    "00100100", --  552 - 0x228  :   36 - 0x24
    "00100100", --  553 - 0x229  :   36 - 0x24
    "00100100", --  554 - 0x22a  :   36 - 0x24
    "00100100", --  555 - 0x22b  :   36 - 0x24
    "00100100", --  556 - 0x22c  :   36 - 0x24
    "00100100", --  557 - 0x22d  :   36 - 0x24
    "00100100", --  558 - 0x22e  :   36 - 0x24
    "00100100", --  559 - 0x22f  :   36 - 0x24
    "00100100", --  560 - 0x230  :   36 - 0x24
    "00100100", --  561 - 0x231  :   36 - 0x24
    "00100100", --  562 - 0x232  :   36 - 0x24
    "00100100", --  563 - 0x233  :   36 - 0x24
    "00100100", --  564 - 0x234  :   36 - 0x24
    "00100100", --  565 - 0x235  :   36 - 0x24
    "00100100", --  566 - 0x236  :   36 - 0x24
    "00100100", --  567 - 0x237  :   36 - 0x24
    "00100100", --  568 - 0x238  :   36 - 0x24
    "00100100", --  569 - 0x239  :   36 - 0x24
    "00100100", --  570 - 0x23a  :   36 - 0x24
    "00100100", --  571 - 0x23b  :   36 - 0x24
    "00100100", --  572 - 0x23c  :   36 - 0x24
    "00100100", --  573 - 0x23d  :   36 - 0x24
    "00100100", --  574 - 0x23e  :   36 - 0x24
    "00100100", --  575 - 0x23f  :   36 - 0x24
    "00100100", --  576 - 0x240  :   36 - 0x24 -- line 0x12
    "00100100", --  577 - 0x241  :   36 - 0x24
    "00100100", --  578 - 0x242  :   36 - 0x24
    "00100100", --  579 - 0x243  :   36 - 0x24
    "00100100", --  580 - 0x244  :   36 - 0x24
    "00100100", --  581 - 0x245  :   36 - 0x24
    "00100100", --  582 - 0x246  :   36 - 0x24
    "00100100", --  583 - 0x247  :   36 - 0x24
    "01000101", --  584 - 0x248  :   69 - 0x45
    "01000101", --  585 - 0x249  :   69 - 0x45
    "01000101", --  586 - 0x24a  :   69 - 0x45
    "01000101", --  587 - 0x24b  :   69 - 0x45
    "00100100", --  588 - 0x24c  :   36 - 0x24
    "00100100", --  589 - 0x24d  :   36 - 0x24
    "00100100", --  590 - 0x24e  :   36 - 0x24
    "00100100", --  591 - 0x24f  :   36 - 0x24
    "00100100", --  592 - 0x250  :   36 - 0x24
    "00100100", --  593 - 0x251  :   36 - 0x24
    "00100100", --  594 - 0x252  :   36 - 0x24
    "00100100", --  595 - 0x253  :   36 - 0x24
    "01010011", --  596 - 0x254  :   83 - 0x53
    "01010100", --  597 - 0x255  :   84 - 0x54
    "00100100", --  598 - 0x256  :   36 - 0x24
    "00100100", --  599 - 0x257  :   36 - 0x24
    "00100100", --  600 - 0x258  :   36 - 0x24
    "00100100", --  601 - 0x259  :   36 - 0x24
    "01010011", --  602 - 0x25a  :   83 - 0x53
    "01010100", --  603 - 0x25b  :   84 - 0x54
    "00100100", --  604 - 0x25c  :   36 - 0x24
    "00100100", --  605 - 0x25d  :   36 - 0x24
    "00100100", --  606 - 0x25e  :   36 - 0x24
    "00100100", --  607 - 0x25f  :   36 - 0x24
    "00100100", --  608 - 0x260  :   36 - 0x24 -- line 0x13
    "00100100", --  609 - 0x261  :   36 - 0x24
    "00100100", --  610 - 0x262  :   36 - 0x24
    "00100100", --  611 - 0x263  :   36 - 0x24
    "00100100", --  612 - 0x264  :   36 - 0x24
    "00100100", --  613 - 0x265  :   36 - 0x24
    "00100100", --  614 - 0x266  :   36 - 0x24
    "00100100", --  615 - 0x267  :   36 - 0x24
    "01000111", --  616 - 0x268  :   71 - 0x47
    "01000111", --  617 - 0x269  :   71 - 0x47
    "01000111", --  618 - 0x26a  :   71 - 0x47
    "01000111", --  619 - 0x26b  :   71 - 0x47
    "00100100", --  620 - 0x26c  :   36 - 0x24
    "00100100", --  621 - 0x26d  :   36 - 0x24
    "00100100", --  622 - 0x26e  :   36 - 0x24
    "00100100", --  623 - 0x26f  :   36 - 0x24
    "00100100", --  624 - 0x270  :   36 - 0x24
    "00100100", --  625 - 0x271  :   36 - 0x24
    "00100100", --  626 - 0x272  :   36 - 0x24
    "00100100", --  627 - 0x273  :   36 - 0x24
    "01010101", --  628 - 0x274  :   85 - 0x55
    "01010110", --  629 - 0x275  :   86 - 0x56
    "00100100", --  630 - 0x276  :   36 - 0x24
    "00100100", --  631 - 0x277  :   36 - 0x24
    "00100100", --  632 - 0x278  :   36 - 0x24
    "00100100", --  633 - 0x279  :   36 - 0x24
    "01010101", --  634 - 0x27a  :   85 - 0x55
    "01010110", --  635 - 0x27b  :   86 - 0x56
    "00100100", --  636 - 0x27c  :   36 - 0x24
    "00100100", --  637 - 0x27d  :   36 - 0x24
    "00100100", --  638 - 0x27e  :   36 - 0x24
    "00100100", --  639 - 0x27f  :   36 - 0x24
    "00100100", --  640 - 0x280  :   36 - 0x24 -- line 0x14
    "00100100", --  641 - 0x281  :   36 - 0x24
    "00100100", --  642 - 0x282  :   36 - 0x24
    "00100100", --  643 - 0x283  :   36 - 0x24
    "00100100", --  644 - 0x284  :   36 - 0x24
    "00100100", --  645 - 0x285  :   36 - 0x24
    "00100100", --  646 - 0x286  :   36 - 0x24
    "00100100", --  647 - 0x287  :   36 - 0x24
    "00100100", --  648 - 0x288  :   36 - 0x24
    "00100100", --  649 - 0x289  :   36 - 0x24
    "00100100", --  650 - 0x28a  :   36 - 0x24
    "00100100", --  651 - 0x28b  :   36 - 0x24
    "00100100", --  652 - 0x28c  :   36 - 0x24
    "00100100", --  653 - 0x28d  :   36 - 0x24
    "00100100", --  654 - 0x28e  :   36 - 0x24
    "00100100", --  655 - 0x28f  :   36 - 0x24
    "00100100", --  656 - 0x290  :   36 - 0x24
    "00100100", --  657 - 0x291  :   36 - 0x24
    "00100100", --  658 - 0x292  :   36 - 0x24
    "00100100", --  659 - 0x293  :   36 - 0x24
    "00100100", --  660 - 0x294  :   36 - 0x24
    "00100100", --  661 - 0x295  :   36 - 0x24
    "00100100", --  662 - 0x296  :   36 - 0x24
    "00100100", --  663 - 0x297  :   36 - 0x24
    "00100100", --  664 - 0x298  :   36 - 0x24
    "00100100", --  665 - 0x299  :   36 - 0x24
    "00100100", --  666 - 0x29a  :   36 - 0x24
    "00100100", --  667 - 0x29b  :   36 - 0x24
    "00100100", --  668 - 0x29c  :   36 - 0x24
    "00100100", --  669 - 0x29d  :   36 - 0x24
    "00100100", --  670 - 0x29e  :   36 - 0x24
    "00100100", --  671 - 0x29f  :   36 - 0x24
    "00100100", --  672 - 0x2a0  :   36 - 0x24 -- line 0x15
    "00100100", --  673 - 0x2a1  :   36 - 0x24
    "00100100", --  674 - 0x2a2  :   36 - 0x24
    "00100100", --  675 - 0x2a3  :   36 - 0x24
    "00110001", --  676 - 0x2a4  :   49 - 0x31
    "00110010", --  677 - 0x2a5  :   50 - 0x32
    "00100100", --  678 - 0x2a6  :   36 - 0x24
    "00100100", --  679 - 0x2a7  :   36 - 0x24
    "00100100", --  680 - 0x2a8  :   36 - 0x24
    "00100100", --  681 - 0x2a9  :   36 - 0x24
    "00100100", --  682 - 0x2aa  :   36 - 0x24
    "00100100", --  683 - 0x2ab  :   36 - 0x24
    "00100100", --  684 - 0x2ac  :   36 - 0x24
    "00100100", --  685 - 0x2ad  :   36 - 0x24
    "00100100", --  686 - 0x2ae  :   36 - 0x24
    "00100100", --  687 - 0x2af  :   36 - 0x24
    "00100100", --  688 - 0x2b0  :   36 - 0x24
    "00100100", --  689 - 0x2b1  :   36 - 0x24
    "00100100", --  690 - 0x2b2  :   36 - 0x24
    "00100100", --  691 - 0x2b3  :   36 - 0x24
    "00100100", --  692 - 0x2b4  :   36 - 0x24
    "00100100", --  693 - 0x2b5  :   36 - 0x24
    "00100100", --  694 - 0x2b6  :   36 - 0x24
    "00100100", --  695 - 0x2b7  :   36 - 0x24
    "00100100", --  696 - 0x2b8  :   36 - 0x24
    "00100100", --  697 - 0x2b9  :   36 - 0x24
    "00100100", --  698 - 0x2ba  :   36 - 0x24
    "00100100", --  699 - 0x2bb  :   36 - 0x24
    "00100100", --  700 - 0x2bc  :   36 - 0x24
    "00100100", --  701 - 0x2bd  :   36 - 0x24
    "00100100", --  702 - 0x2be  :   36 - 0x24
    "00100100", --  703 - 0x2bf  :   36 - 0x24
    "00100100", --  704 - 0x2c0  :   36 - 0x24 -- line 0x16
    "00100100", --  705 - 0x2c1  :   36 - 0x24
    "00100100", --  706 - 0x2c2  :   36 - 0x24
    "00110000", --  707 - 0x2c3  :   48 - 0x30
    "00100110", --  708 - 0x2c4  :   38 - 0x26
    "00110100", --  709 - 0x2c5  :   52 - 0x34
    "00110011", --  710 - 0x2c6  :   51 - 0x33
    "00100100", --  711 - 0x2c7  :   36 - 0x24
    "00100100", --  712 - 0x2c8  :   36 - 0x24
    "00100100", --  713 - 0x2c9  :   36 - 0x24
    "00100100", --  714 - 0x2ca  :   36 - 0x24
    "00100100", --  715 - 0x2cb  :   36 - 0x24
    "00100100", --  716 - 0x2cc  :   36 - 0x24
    "00100100", --  717 - 0x2cd  :   36 - 0x24
    "00100100", --  718 - 0x2ce  :   36 - 0x24
    "00100100", --  719 - 0x2cf  :   36 - 0x24
    "00100100", --  720 - 0x2d0  :   36 - 0x24
    "00100100", --  721 - 0x2d1  :   36 - 0x24
    "00100100", --  722 - 0x2d2  :   36 - 0x24
    "00100100", --  723 - 0x2d3  :   36 - 0x24
    "00100100", --  724 - 0x2d4  :   36 - 0x24
    "00100100", --  725 - 0x2d5  :   36 - 0x24
    "00100100", --  726 - 0x2d6  :   36 - 0x24
    "00100100", --  727 - 0x2d7  :   36 - 0x24
    "00100100", --  728 - 0x2d8  :   36 - 0x24
    "00100100", --  729 - 0x2d9  :   36 - 0x24
    "00100100", --  730 - 0x2da  :   36 - 0x24
    "00100100", --  731 - 0x2db  :   36 - 0x24
    "00100100", --  732 - 0x2dc  :   36 - 0x24
    "00100100", --  733 - 0x2dd  :   36 - 0x24
    "00100100", --  734 - 0x2de  :   36 - 0x24
    "00100100", --  735 - 0x2df  :   36 - 0x24
    "00100100", --  736 - 0x2e0  :   36 - 0x24 -- line 0x17
    "00100100", --  737 - 0x2e1  :   36 - 0x24
    "00110000", --  738 - 0x2e2  :   48 - 0x30
    "00100110", --  739 - 0x2e3  :   38 - 0x26
    "00100110", --  740 - 0x2e4  :   38 - 0x26
    "00100110", --  741 - 0x2e5  :   38 - 0x26
    "00100110", --  742 - 0x2e6  :   38 - 0x26
    "00110011", --  743 - 0x2e7  :   51 - 0x33
    "00100100", --  744 - 0x2e8  :   36 - 0x24
    "00100100", --  745 - 0x2e9  :   36 - 0x24
    "00100100", --  746 - 0x2ea  :   36 - 0x24
    "00100100", --  747 - 0x2eb  :   36 - 0x24
    "00100100", --  748 - 0x2ec  :   36 - 0x24
    "00100100", --  749 - 0x2ed  :   36 - 0x24
    "00100100", --  750 - 0x2ee  :   36 - 0x24
    "00100100", --  751 - 0x2ef  :   36 - 0x24
    "00100100", --  752 - 0x2f0  :   36 - 0x24
    "00100100", --  753 - 0x2f1  :   36 - 0x24
    "00100100", --  754 - 0x2f2  :   36 - 0x24
    "00100100", --  755 - 0x2f3  :   36 - 0x24
    "00100100", --  756 - 0x2f4  :   36 - 0x24
    "00100100", --  757 - 0x2f5  :   36 - 0x24
    "00100100", --  758 - 0x2f6  :   36 - 0x24
    "00100100", --  759 - 0x2f7  :   36 - 0x24
    "00100100", --  760 - 0x2f8  :   36 - 0x24
    "00100100", --  761 - 0x2f9  :   36 - 0x24
    "00100100", --  762 - 0x2fa  :   36 - 0x24
    "00100100", --  763 - 0x2fb  :   36 - 0x24
    "00100100", --  764 - 0x2fc  :   36 - 0x24
    "00100100", --  765 - 0x2fd  :   36 - 0x24
    "00100100", --  766 - 0x2fe  :   36 - 0x24
    "00100100", --  767 - 0x2ff  :   36 - 0x24
    "00100100", --  768 - 0x300  :   36 - 0x24 -- line 0x18
    "00110000", --  769 - 0x301  :   48 - 0x30
    "00100110", --  770 - 0x302  :   38 - 0x26
    "00110100", --  771 - 0x303  :   52 - 0x34
    "00100110", --  772 - 0x304  :   38 - 0x26
    "00100110", --  773 - 0x305  :   38 - 0x26
    "00110100", --  774 - 0x306  :   52 - 0x34
    "00100110", --  775 - 0x307  :   38 - 0x26
    "00110011", --  776 - 0x308  :   51 - 0x33
    "00100100", --  777 - 0x309  :   36 - 0x24
    "00100100", --  778 - 0x30a  :   36 - 0x24
    "00100100", --  779 - 0x30b  :   36 - 0x24
    "00100100", --  780 - 0x30c  :   36 - 0x24
    "00100100", --  781 - 0x30d  :   36 - 0x24
    "00100100", --  782 - 0x30e  :   36 - 0x24
    "00100100", --  783 - 0x30f  :   36 - 0x24
    "00100100", --  784 - 0x310  :   36 - 0x24
    "00100100", --  785 - 0x311  :   36 - 0x24
    "00100100", --  786 - 0x312  :   36 - 0x24
    "00100100", --  787 - 0x313  :   36 - 0x24
    "00100100", --  788 - 0x314  :   36 - 0x24
    "00100100", --  789 - 0x315  :   36 - 0x24
    "00100100", --  790 - 0x316  :   36 - 0x24
    "00100100", --  791 - 0x317  :   36 - 0x24
    "00110110", --  792 - 0x318  :   54 - 0x36
    "00110111", --  793 - 0x319  :   55 - 0x37
    "00110110", --  794 - 0x31a  :   54 - 0x36
    "00110111", --  795 - 0x31b  :   55 - 0x37
    "00110110", --  796 - 0x31c  :   54 - 0x36
    "00110111", --  797 - 0x31d  :   55 - 0x37
    "00100100", --  798 - 0x31e  :   36 - 0x24
    "00100100", --  799 - 0x31f  :   36 - 0x24
    "00110000", --  800 - 0x320  :   48 - 0x30 -- line 0x19
    "00100110", --  801 - 0x321  :   38 - 0x26
    "00100110", --  802 - 0x322  :   38 - 0x26
    "00100110", --  803 - 0x323  :   38 - 0x26
    "00100110", --  804 - 0x324  :   38 - 0x26
    "00100110", --  805 - 0x325  :   38 - 0x26
    "00100110", --  806 - 0x326  :   38 - 0x26
    "00100110", --  807 - 0x327  :   38 - 0x26
    "00100110", --  808 - 0x328  :   38 - 0x26
    "00110011", --  809 - 0x329  :   51 - 0x33
    "00100100", --  810 - 0x32a  :   36 - 0x24
    "00100100", --  811 - 0x32b  :   36 - 0x24
    "00100100", --  812 - 0x32c  :   36 - 0x24
    "00100100", --  813 - 0x32d  :   36 - 0x24
    "00100100", --  814 - 0x32e  :   36 - 0x24
    "00100100", --  815 - 0x32f  :   36 - 0x24
    "00100100", --  816 - 0x330  :   36 - 0x24
    "00100100", --  817 - 0x331  :   36 - 0x24
    "00100100", --  818 - 0x332  :   36 - 0x24
    "00100100", --  819 - 0x333  :   36 - 0x24
    "00100100", --  820 - 0x334  :   36 - 0x24
    "00100100", --  821 - 0x335  :   36 - 0x24
    "00100100", --  822 - 0x336  :   36 - 0x24
    "00110101", --  823 - 0x337  :   53 - 0x35
    "00100101", --  824 - 0x338  :   37 - 0x25
    "00100101", --  825 - 0x339  :   37 - 0x25
    "00100101", --  826 - 0x33a  :   37 - 0x25
    "00100101", --  827 - 0x33b  :   37 - 0x25
    "00100101", --  828 - 0x33c  :   37 - 0x25
    "00100101", --  829 - 0x33d  :   37 - 0x25
    "00111000", --  830 - 0x33e  :   56 - 0x38
    "00100100", --  831 - 0x33f  :   36 - 0x24
    "10110100", --  832 - 0x340  :  180 - 0xb4 -- line 0x1a
    "10110101", --  833 - 0x341  :  181 - 0xb5
    "10110100", --  834 - 0x342  :  180 - 0xb4
    "10110101", --  835 - 0x343  :  181 - 0xb5
    "10110100", --  836 - 0x344  :  180 - 0xb4
    "10110101", --  837 - 0x345  :  181 - 0xb5
    "10110100", --  838 - 0x346  :  180 - 0xb4
    "10110101", --  839 - 0x347  :  181 - 0xb5
    "10110100", --  840 - 0x348  :  180 - 0xb4
    "10110101", --  841 - 0x349  :  181 - 0xb5
    "10110100", --  842 - 0x34a  :  180 - 0xb4
    "10110101", --  843 - 0x34b  :  181 - 0xb5
    "10110100", --  844 - 0x34c  :  180 - 0xb4
    "10110101", --  845 - 0x34d  :  181 - 0xb5
    "10110100", --  846 - 0x34e  :  180 - 0xb4
    "10110101", --  847 - 0x34f  :  181 - 0xb5
    "10110100", --  848 - 0x350  :  180 - 0xb4
    "10110101", --  849 - 0x351  :  181 - 0xb5
    "10110100", --  850 - 0x352  :  180 - 0xb4
    "10110101", --  851 - 0x353  :  181 - 0xb5
    "10110100", --  852 - 0x354  :  180 - 0xb4
    "10110101", --  853 - 0x355  :  181 - 0xb5
    "10110100", --  854 - 0x356  :  180 - 0xb4
    "10110101", --  855 - 0x357  :  181 - 0xb5
    "10110100", --  856 - 0x358  :  180 - 0xb4
    "10110101", --  857 - 0x359  :  181 - 0xb5
    "10110100", --  858 - 0x35a  :  180 - 0xb4
    "10110101", --  859 - 0x35b  :  181 - 0xb5
    "10110100", --  860 - 0x35c  :  180 - 0xb4
    "10110101", --  861 - 0x35d  :  181 - 0xb5
    "10110100", --  862 - 0x35e  :  180 - 0xb4
    "10110101", --  863 - 0x35f  :  181 - 0xb5
    "10110110", --  864 - 0x360  :  182 - 0xb6 -- line 0x1b
    "10110111", --  865 - 0x361  :  183 - 0xb7
    "10110110", --  866 - 0x362  :  182 - 0xb6
    "10110111", --  867 - 0x363  :  183 - 0xb7
    "10110110", --  868 - 0x364  :  182 - 0xb6
    "10110111", --  869 - 0x365  :  183 - 0xb7
    "10110110", --  870 - 0x366  :  182 - 0xb6
    "10110111", --  871 - 0x367  :  183 - 0xb7
    "10110110", --  872 - 0x368  :  182 - 0xb6
    "10110111", --  873 - 0x369  :  183 - 0xb7
    "10110110", --  874 - 0x36a  :  182 - 0xb6
    "10110111", --  875 - 0x36b  :  183 - 0xb7
    "10110110", --  876 - 0x36c  :  182 - 0xb6
    "10110111", --  877 - 0x36d  :  183 - 0xb7
    "10110110", --  878 - 0x36e  :  182 - 0xb6
    "10110111", --  879 - 0x36f  :  183 - 0xb7
    "10110110", --  880 - 0x370  :  182 - 0xb6
    "10110111", --  881 - 0x371  :  183 - 0xb7
    "10110110", --  882 - 0x372  :  182 - 0xb6
    "10110111", --  883 - 0x373  :  183 - 0xb7
    "10110110", --  884 - 0x374  :  182 - 0xb6
    "10110111", --  885 - 0x375  :  183 - 0xb7
    "10110110", --  886 - 0x376  :  182 - 0xb6
    "10110111", --  887 - 0x377  :  183 - 0xb7
    "10110110", --  888 - 0x378  :  182 - 0xb6
    "10110111", --  889 - 0x379  :  183 - 0xb7
    "10110110", --  890 - 0x37a  :  182 - 0xb6
    "10110111", --  891 - 0x37b  :  183 - 0xb7
    "10110110", --  892 - 0x37c  :  182 - 0xb6
    "10110111", --  893 - 0x37d  :  183 - 0xb7
    "10110110", --  894 - 0x37e  :  182 - 0xb6
    "10110111", --  895 - 0x37f  :  183 - 0xb7
    "10110100", --  896 - 0x380  :  180 - 0xb4 -- line 0x1c
    "10110101", --  897 - 0x381  :  181 - 0xb5
    "10110100", --  898 - 0x382  :  180 - 0xb4
    "10110101", --  899 - 0x383  :  181 - 0xb5
    "10110100", --  900 - 0x384  :  180 - 0xb4
    "10110101", --  901 - 0x385  :  181 - 0xb5
    "10110100", --  902 - 0x386  :  180 - 0xb4
    "10110101", --  903 - 0x387  :  181 - 0xb5
    "10110100", --  904 - 0x388  :  180 - 0xb4
    "10110101", --  905 - 0x389  :  181 - 0xb5
    "10110100", --  906 - 0x38a  :  180 - 0xb4
    "10110101", --  907 - 0x38b  :  181 - 0xb5
    "10110100", --  908 - 0x38c  :  180 - 0xb4
    "10110101", --  909 - 0x38d  :  181 - 0xb5
    "10110100", --  910 - 0x38e  :  180 - 0xb4
    "10110101", --  911 - 0x38f  :  181 - 0xb5
    "10110100", --  912 - 0x390  :  180 - 0xb4
    "10110101", --  913 - 0x391  :  181 - 0xb5
    "10110100", --  914 - 0x392  :  180 - 0xb4
    "10110101", --  915 - 0x393  :  181 - 0xb5
    "10110100", --  916 - 0x394  :  180 - 0xb4
    "10110101", --  917 - 0x395  :  181 - 0xb5
    "10110100", --  918 - 0x396  :  180 - 0xb4
    "10110101", --  919 - 0x397  :  181 - 0xb5
    "10110100", --  920 - 0x398  :  180 - 0xb4
    "10110101", --  921 - 0x399  :  181 - 0xb5
    "10110100", --  922 - 0x39a  :  180 - 0xb4
    "10110101", --  923 - 0x39b  :  181 - 0xb5
    "10110100", --  924 - 0x39c  :  180 - 0xb4
    "10110101", --  925 - 0x39d  :  181 - 0xb5
    "10110100", --  926 - 0x39e  :  180 - 0xb4
    "10110101", --  927 - 0x39f  :  181 - 0xb5
    "10110110", --  928 - 0x3a0  :  182 - 0xb6 -- line 0x1d
    "10110111", --  929 - 0x3a1  :  183 - 0xb7
    "10110110", --  930 - 0x3a2  :  182 - 0xb6
    "10110111", --  931 - 0x3a3  :  183 - 0xb7
    "10110110", --  932 - 0x3a4  :  182 - 0xb6
    "10110111", --  933 - 0x3a5  :  183 - 0xb7
    "10110110", --  934 - 0x3a6  :  182 - 0xb6
    "10110111", --  935 - 0x3a7  :  183 - 0xb7
    "10110110", --  936 - 0x3a8  :  182 - 0xb6
    "10110111", --  937 - 0x3a9  :  183 - 0xb7
    "10110110", --  938 - 0x3aa  :  182 - 0xb6
    "10110111", --  939 - 0x3ab  :  183 - 0xb7
    "10110110", --  940 - 0x3ac  :  182 - 0xb6
    "10110111", --  941 - 0x3ad  :  183 - 0xb7
    "10110110", --  942 - 0x3ae  :  182 - 0xb6
    "10110111", --  943 - 0x3af  :  183 - 0xb7
    "10110110", --  944 - 0x3b0  :  182 - 0xb6
    "10110111", --  945 - 0x3b1  :  183 - 0xb7
    "10110110", --  946 - 0x3b2  :  182 - 0xb6
    "10110111", --  947 - 0x3b3  :  183 - 0xb7
    "10110110", --  948 - 0x3b4  :  182 - 0xb6
    "10110111", --  949 - 0x3b5  :  183 - 0xb7
    "10110110", --  950 - 0x3b6  :  182 - 0xb6
    "10110111", --  951 - 0x3b7  :  183 - 0xb7
    "10110110", --  952 - 0x3b8  :  182 - 0xb6
    "10110111", --  953 - 0x3b9  :  183 - 0xb7
    "10110110", --  954 - 0x3ba  :  182 - 0xb6
    "10110111", --  955 - 0x3bb  :  183 - 0xb7
    "10110110", --  956 - 0x3bc  :  182 - 0xb6
    "10110111", --  957 - 0x3bd  :  183 - 0xb7
    "10110110", --  958 - 0x3be  :  182 - 0xb6
    "10110111", --  959 - 0x3bf  :  183 - 0xb7
        ---- Attribute Table 0----
    "10101010", --  960 - 0x3c0  :  170 - 0xaa
    "10101010", --  961 - 0x3c1  :  170 - 0xaa
    "11101010", --  962 - 0x3c2  :  234 - 0xea
    "10101010", --  963 - 0x3c3  :  170 - 0xaa
    "10101010", --  964 - 0x3c4  :  170 - 0xaa
    "10101010", --  965 - 0x3c5  :  170 - 0xaa
    "10101010", --  966 - 0x3c6  :  170 - 0xaa
    "10101010", --  967 - 0x3c7  :  170 - 0xaa
    "00000000", --  968 - 0x3c8  :    0 - 0x0
    "00000000", --  969 - 0x3c9  :    0 - 0x0
    "00000000", --  970 - 0x3ca  :    0 - 0x0
    "00000000", --  971 - 0x3cb  :    0 - 0x0
    "10100000", --  972 - 0x3cc  :  160 - 0xa0
    "00100000", --  973 - 0x3cd  :   32 - 0x20
    "00000000", --  974 - 0x3ce  :    0 - 0x0
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "00000000", --  976 - 0x3d0  :    0 - 0x0
    "00000000", --  977 - 0x3d1  :    0 - 0x0
    "00000000", --  978 - 0x3d2  :    0 - 0x0
    "00000000", --  979 - 0x3d3  :    0 - 0x0
    "00001010", --  980 - 0x3d4  :   10 - 0xa
    "00000010", --  981 - 0x3d5  :    2 - 0x2
    "11000000", --  982 - 0x3d6  :  192 - 0xc0
    "00000000", --  983 - 0x3d7  :    0 - 0x0
    "00000000", --  984 - 0x3d8  :    0 - 0x0
    "00000000", --  985 - 0x3d9  :    0 - 0x0
    "00000000", --  986 - 0x3da  :    0 - 0x0
    "00000000", --  987 - 0x3db  :    0 - 0x0
    "00000000", --  988 - 0x3dc  :    0 - 0x0
    "00000000", --  989 - 0x3dd  :    0 - 0x0
    "00000000", --  990 - 0x3de  :    0 - 0x0
    "00000000", --  991 - 0x3df  :    0 - 0x0
    "00000000", --  992 - 0x3e0  :    0 - 0x0
    "00000000", --  993 - 0x3e1  :    0 - 0x0
    "01010000", --  994 - 0x3e2  :   80 - 0x50
    "00000000", --  995 - 0x3e3  :    0 - 0x0
    "00000000", --  996 - 0x3e4  :    0 - 0x0
    "00110000", --  997 - 0x3e5  :   48 - 0x30
    "11000000", --  998 - 0x3e6  :  192 - 0xc0
    "00000000", --  999 - 0x3e7  :    0 - 0x0
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0
    "00000000", -- 1001 - 0x3e9  :    0 - 0x0
    "00000000", -- 1002 - 0x3ea  :    0 - 0x0
    "00000000", -- 1003 - 0x3eb  :    0 - 0x0
    "00000000", -- 1004 - 0x3ec  :    0 - 0x0
    "00000000", -- 1005 - 0x3ed  :    0 - 0x0
    "00000000", -- 1006 - 0x3ee  :    0 - 0x0
    "00000000", -- 1007 - 0x3ef  :    0 - 0x0
    "01010000", -- 1008 - 0x3f0  :   80 - 0x50
    "01010000", -- 1009 - 0x3f1  :   80 - 0x50
    "01010000", -- 1010 - 0x3f2  :   80 - 0x50
    "01010000", -- 1011 - 0x3f3  :   80 - 0x50
    "01010000", -- 1012 - 0x3f4  :   80 - 0x50
    "01010000", -- 1013 - 0x3f5  :   80 - 0x50
    "01010000", -- 1014 - 0x3f6  :   80 - 0x50
    "01010000", -- 1015 - 0x3f7  :   80 - 0x50
    "00000101", -- 1016 - 0x3f8  :    5 - 0x5
    "00000101", -- 1017 - 0x3f9  :    5 - 0x5
    "00000101", -- 1018 - 0x3fa  :    5 - 0x5
    "00000101", -- 1019 - 0x3fb  :    5 - 0x5
    "00000101", -- 1020 - 0x3fc  :    5 - 0x5
    "00000101", -- 1021 - 0x3fd  :    5 - 0x5
    "00000101", -- 1022 - 0x3fe  :    5 - 0x5
    "00000101"  -- 1023 - 0x3ff  :    5 - 0x5
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
