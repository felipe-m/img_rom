--- Autcmatically generated VHDL ROM from a NES memory file----
---   NAME TABLE
-- https://wiki.nesdev.com/w/index.php/PPU_nametables
--- Only the first Name Table: 1KiB


---  Original memory dump file name: lawnmower_ntable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_NTABLE_LAWN_00 is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(10-1 downto 0);  --1024 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_NTABLE_LAWN_00;

architecture BEHAVIORAL of ROM_NTABLE_LAWN_00 is
  signal addr_int  : natural range 0 to 2**10-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
     ------- Name Table 0---------
    "10101001", --    0 -  0x0  :  169 - 0xa9 -- line 0x0
    "10101001", --    1 -  0x1  :  169 - 0xa9
    "10101001", --    2 -  0x2  :  169 - 0xa9
    "10101001", --    3 -  0x3  :  169 - 0xa9
    "10101001", --    4 -  0x4  :  169 - 0xa9
    "10101001", --    5 -  0x5  :  169 - 0xa9
    "10101001", --    6 -  0x6  :  169 - 0xa9
    "10101001", --    7 -  0x7  :  169 - 0xa9
    "10101001", --    8 -  0x8  :  169 - 0xa9
    "10101001", --    9 -  0x9  :  169 - 0xa9
    "10101001", --   10 -  0xa  :  169 - 0xa9
    "10101001", --   11 -  0xb  :  169 - 0xa9
    "10101001", --   12 -  0xc  :  169 - 0xa9
    "10101001", --   13 -  0xd  :  169 - 0xa9
    "10101001", --   14 -  0xe  :  169 - 0xa9
    "10101001", --   15 -  0xf  :  169 - 0xa9
    "10101001", --   16 - 0x10  :  169 - 0xa9
    "10101001", --   17 - 0x11  :  169 - 0xa9
    "10101001", --   18 - 0x12  :  169 - 0xa9
    "10101001", --   19 - 0x13  :  169 - 0xa9
    "10101001", --   20 - 0x14  :  169 - 0xa9
    "10101001", --   21 - 0x15  :  169 - 0xa9
    "10101001", --   22 - 0x16  :  169 - 0xa9
    "10101001", --   23 - 0x17  :  169 - 0xa9
    "10101001", --   24 - 0x18  :  169 - 0xa9
    "10101001", --   25 - 0x19  :  169 - 0xa9
    "10101001", --   26 - 0x1a  :  169 - 0xa9
    "10101001", --   27 - 0x1b  :  169 - 0xa9
    "10101001", --   28 - 0x1c  :  169 - 0xa9
    "10101001", --   29 - 0x1d  :  169 - 0xa9
    "10101001", --   30 - 0x1e  :  169 - 0xa9
    "10101001", --   31 - 0x1f  :  169 - 0xa9
    "10101001", --   32 - 0x20  :  169 - 0xa9 -- line 0x1
    "10101001", --   33 - 0x21  :  169 - 0xa9
    "10101001", --   34 - 0x22  :  169 - 0xa9
    "10101001", --   35 - 0x23  :  169 - 0xa9
    "10101001", --   36 - 0x24  :  169 - 0xa9
    "10101001", --   37 - 0x25  :  169 - 0xa9
    "10101001", --   38 - 0x26  :  169 - 0xa9
    "10101001", --   39 - 0x27  :  169 - 0xa9
    "10101001", --   40 - 0x28  :  169 - 0xa9
    "10101001", --   41 - 0x29  :  169 - 0xa9
    "10101001", --   42 - 0x2a  :  169 - 0xa9
    "10101001", --   43 - 0x2b  :  169 - 0xa9
    "10101001", --   44 - 0x2c  :  169 - 0xa9
    "10101001", --   45 - 0x2d  :  169 - 0xa9
    "10101001", --   46 - 0x2e  :  169 - 0xa9
    "10101001", --   47 - 0x2f  :  169 - 0xa9
    "10101001", --   48 - 0x30  :  169 - 0xa9
    "10101001", --   49 - 0x31  :  169 - 0xa9
    "10101001", --   50 - 0x32  :  169 - 0xa9
    "10101001", --   51 - 0x33  :  169 - 0xa9
    "10101001", --   52 - 0x34  :  169 - 0xa9
    "10101001", --   53 - 0x35  :  169 - 0xa9
    "10101001", --   54 - 0x36  :  169 - 0xa9
    "10101001", --   55 - 0x37  :  169 - 0xa9
    "10101001", --   56 - 0x38  :  169 - 0xa9
    "10101001", --   57 - 0x39  :  169 - 0xa9
    "10101001", --   58 - 0x3a  :  169 - 0xa9
    "10101001", --   59 - 0x3b  :  169 - 0xa9
    "10101001", --   60 - 0x3c  :  169 - 0xa9
    "10101001", --   61 - 0x3d  :  169 - 0xa9
    "10101001", --   62 - 0x3e  :  169 - 0xa9
    "10101001", --   63 - 0x3f  :  169 - 0xa9
    "10101001", --   64 - 0x40  :  169 - 0xa9 -- line 0x2
    "10101001", --   65 - 0x41  :  169 - 0xa9
    "01010110", --   66 - 0x42  :   86 - 0x56
    "01010101", --   67 - 0x43  :   85 - 0x55
    "01010111", --   68 - 0x44  :   87 - 0x57
    "01011000", --   69 - 0x45  :   88 - 0x58
    "11010000", --   70 - 0x46  :  208 - 0xd0
    "11010001", --   71 - 0x47  :  209 - 0xd1
    "10101001", --   72 - 0x48  :  169 - 0xa9
    "01011101", --   73 - 0x49  :   93 - 0x5d
    "01011110", --   74 - 0x4a  :   94 - 0x5e
    "01011011", --   75 - 0x4b  :   91 - 0x5b
    "01010110", --   76 - 0x4c  :   86 - 0x56
    "11111001", --   77 - 0x4d  :  249 - 0xf9
    "11111010", --   78 - 0x4e  :  250 - 0xfa
    "11111010", --   79 - 0x4f  :  250 - 0xfa
    "11111010", --   80 - 0x50  :  250 - 0xfa
    "11111010", --   81 - 0x51  :  250 - 0xfa
    "11111010", --   82 - 0x52  :  250 - 0xfa
    "11111010", --   83 - 0x53  :  250 - 0xfa
    "11111011", --   84 - 0x54  :  251 - 0xfb
    "10101001", --   85 - 0x55  :  169 - 0xa9
    "01011001", --   86 - 0x56  :   89 - 0x59
    "01011010", --   87 - 0x57  :   90 - 0x5a
    "01011000", --   88 - 0x58  :   88 - 0x58
    "01011011", --   89 - 0x59  :   91 - 0x5b
    "11010000", --   90 - 0x5a  :  208 - 0xd0
    "11010000", --   91 - 0x5b  :  208 - 0xd0
    "11010000", --   92 - 0x5c  :  208 - 0xd0
    "01011100", --   93 - 0x5d  :   92 - 0x5c
    "10101001", --   94 - 0x5e  :  169 - 0xa9
    "10101001", --   95 - 0x5f  :  169 - 0xa9
    "10101001", --   96 - 0x60  :  169 - 0xa9 -- line 0x3
    "10101001", --   97 - 0x61  :  169 - 0xa9
    "01100110", --   98 - 0x62  :  102 - 0x66
    "01100101", --   99 - 0x63  :  101 - 0x65
    "01100111", --  100 - 0x64  :  103 - 0x67
    "01101000", --  101 - 0x65  :  104 - 0x68
    "11100000", --  102 - 0x66  :  224 - 0xe0
    "11100001", --  103 - 0x67  :  225 - 0xe1
    "10101001", --  104 - 0x68  :  169 - 0xa9
    "01101101", --  105 - 0x69  :  109 - 0x6d
    "01101110", --  106 - 0x6a  :  110 - 0x6e
    "01101011", --  107 - 0x6b  :  107 - 0x6b
    "01100110", --  108 - 0x6c  :  102 - 0x66
    "11111100", --  109 - 0x6d  :  252 - 0xfc
    "11111101", --  110 - 0x6e  :  253 - 0xfd
    "11111101", --  111 - 0x6f  :  253 - 0xfd
    "11111101", --  112 - 0x70  :  253 - 0xfd
    "11111101", --  113 - 0x71  :  253 - 0xfd
    "11111101", --  114 - 0x72  :  253 - 0xfd
    "11111101", --  115 - 0x73  :  253 - 0xfd
    "11111110", --  116 - 0x74  :  254 - 0xfe
    "10101001", --  117 - 0x75  :  169 - 0xa9
    "01101001", --  118 - 0x76  :  105 - 0x69
    "01101010", --  119 - 0x77  :  106 - 0x6a
    "01101000", --  120 - 0x78  :  104 - 0x68
    "01101011", --  121 - 0x79  :  107 - 0x6b
    "11100000", --  122 - 0x7a  :  224 - 0xe0
    "11100000", --  123 - 0x7b  :  224 - 0xe0
    "11100000", --  124 - 0x7c  :  224 - 0xe0
    "01101100", --  125 - 0x7d  :  108 - 0x6c
    "10101001", --  126 - 0x7e  :  169 - 0xa9
    "10101001", --  127 - 0x7f  :  169 - 0xa9
    "10101010", --  128 - 0x80  :  170 - 0xaa -- line 0x4
    "10101010", --  129 - 0x81  :  170 - 0xaa
    "10101010", --  130 - 0x82  :  170 - 0xaa
    "10101010", --  131 - 0x83  :  170 - 0xaa
    "10101010", --  132 - 0x84  :  170 - 0xaa
    "10101010", --  133 - 0x85  :  170 - 0xaa
    "10101010", --  134 - 0x86  :  170 - 0xaa
    "10101010", --  135 - 0x87  :  170 - 0xaa
    "10101010", --  136 - 0x88  :  170 - 0xaa
    "10101010", --  137 - 0x89  :  170 - 0xaa
    "10101010", --  138 - 0x8a  :  170 - 0xaa
    "10101010", --  139 - 0x8b  :  170 - 0xaa
    "10101010", --  140 - 0x8c  :  170 - 0xaa
    "10101010", --  141 - 0x8d  :  170 - 0xaa
    "10101010", --  142 - 0x8e  :  170 - 0xaa
    "10101010", --  143 - 0x8f  :  170 - 0xaa
    "10101010", --  144 - 0x90  :  170 - 0xaa
    "10101010", --  145 - 0x91  :  170 - 0xaa
    "10101010", --  146 - 0x92  :  170 - 0xaa
    "10101010", --  147 - 0x93  :  170 - 0xaa
    "10101010", --  148 - 0x94  :  170 - 0xaa
    "10101010", --  149 - 0x95  :  170 - 0xaa
    "10101010", --  150 - 0x96  :  170 - 0xaa
    "10101010", --  151 - 0x97  :  170 - 0xaa
    "10101010", --  152 - 0x98  :  170 - 0xaa
    "10101010", --  153 - 0x99  :  170 - 0xaa
    "10101010", --  154 - 0x9a  :  170 - 0xaa
    "10101010", --  155 - 0x9b  :  170 - 0xaa
    "10101010", --  156 - 0x9c  :  170 - 0xaa
    "10101010", --  157 - 0x9d  :  170 - 0xaa
    "10101010", --  158 - 0x9e  :  170 - 0xaa
    "10101010", --  159 - 0x9f  :  170 - 0xaa
    "10100000", --  160 - 0xa0  :  160 - 0xa0 -- line 0x5
    "10100001", --  161 - 0xa1  :  161 - 0xa1
    "10100010", --  162 - 0xa2  :  162 - 0xa2
    "10100010", --  163 - 0xa3  :  162 - 0xa2
    "10100010", --  164 - 0xa4  :  162 - 0xa2
    "10100010", --  165 - 0xa5  :  162 - 0xa2
    "10100010", --  166 - 0xa6  :  162 - 0xa2
    "10100010", --  167 - 0xa7  :  162 - 0xa2
    "10100010", --  168 - 0xa8  :  162 - 0xa2
    "10100010", --  169 - 0xa9  :  162 - 0xa2
    "10100010", --  170 - 0xaa  :  162 - 0xa2
    "10100010", --  171 - 0xab  :  162 - 0xa2
    "10100010", --  172 - 0xac  :  162 - 0xa2
    "10100010", --  173 - 0xad  :  162 - 0xa2
    "10100010", --  174 - 0xae  :  162 - 0xa2
    "10100010", --  175 - 0xaf  :  162 - 0xa2
    "10100010", --  176 - 0xb0  :  162 - 0xa2
    "10100010", --  177 - 0xb1  :  162 - 0xa2
    "10100010", --  178 - 0xb2  :  162 - 0xa2
    "10100010", --  179 - 0xb3  :  162 - 0xa2
    "10100010", --  180 - 0xb4  :  162 - 0xa2
    "10100010", --  181 - 0xb5  :  162 - 0xa2
    "10100010", --  182 - 0xb6  :  162 - 0xa2
    "10100010", --  183 - 0xb7  :  162 - 0xa2
    "10100010", --  184 - 0xb8  :  162 - 0xa2
    "10100010", --  185 - 0xb9  :  162 - 0xa2
    "10100010", --  186 - 0xba  :  162 - 0xa2
    "10100010", --  187 - 0xbb  :  162 - 0xa2
    "10100010", --  188 - 0xbc  :  162 - 0xa2
    "10100010", --  189 - 0xbd  :  162 - 0xa2
    "10100110", --  190 - 0xbe  :  166 - 0xa6
    "10100000", --  191 - 0xbf  :  160 - 0xa0
    "10100000", --  192 - 0xc0  :  160 - 0xa0 -- line 0x6
    "10100011", --  193 - 0xc1  :  163 - 0xa3
    "10000000", --  194 - 0xc2  :  128 - 0x80
    "10000001", --  195 - 0xc3  :  129 - 0x81
    "10000000", --  196 - 0xc4  :  128 - 0x80
    "10000001", --  197 - 0xc5  :  129 - 0x81
    "10000000", --  198 - 0xc6  :  128 - 0x80
    "10000010", --  199 - 0xc7  :  130 - 0x82
    "10000000", --  200 - 0xc8  :  128 - 0x80
    "10000001", --  201 - 0xc9  :  129 - 0x81
    "10000001", --  202 - 0xca  :  129 - 0x81
    "10000000", --  203 - 0xcb  :  128 - 0x80
    "10000000", --  204 - 0xcc  :  128 - 0x80
    "10000001", --  205 - 0xcd  :  129 - 0x81
    "10000010", --  206 - 0xce  :  130 - 0x82
    "10000011", --  207 - 0xcf  :  131 - 0x83
    "10000010", --  208 - 0xd0  :  130 - 0x82
    "10000011", --  209 - 0xd1  :  131 - 0x83
    "10000000", --  210 - 0xd2  :  128 - 0x80
    "10000010", --  211 - 0xd3  :  130 - 0x82
    "10000000", --  212 - 0xd4  :  128 - 0x80
    "10000010", --  213 - 0xd5  :  130 - 0x82
    "10000010", --  214 - 0xd6  :  130 - 0x82
    "10000011", --  215 - 0xd7  :  131 - 0x83
    "10000010", --  216 - 0xd8  :  130 - 0x82
    "10000011", --  217 - 0xd9  :  131 - 0x83
    "10000001", --  218 - 0xda  :  129 - 0x81
    "10000000", --  219 - 0xdb  :  128 - 0x80
    "10000000", --  220 - 0xdc  :  128 - 0x80
    "10000001", --  221 - 0xdd  :  129 - 0x81
    "10100111", --  222 - 0xde  :  167 - 0xa7
    "10100000", --  223 - 0xdf  :  160 - 0xa0
    "10100000", --  224 - 0xe0  :  160 - 0xa0 -- line 0x7
    "10100011", --  225 - 0xe1  :  163 - 0xa3
    "10010000", --  226 - 0xe2  :  144 - 0x90
    "10010001", --  227 - 0xe3  :  145 - 0x91
    "10010000", --  228 - 0xe4  :  144 - 0x90
    "10010001", --  229 - 0xe5  :  145 - 0x91
    "10010010", --  230 - 0xe6  :  146 - 0x92
    "10010001", --  231 - 0xe7  :  145 - 0x91
    "10010000", --  232 - 0xe8  :  144 - 0x90
    "10010001", --  233 - 0xe9  :  145 - 0x91
    "10010011", --  234 - 0xea  :  147 - 0x93
    "10010010", --  235 - 0xeb  :  146 - 0x92
    "10010000", --  236 - 0xec  :  144 - 0x90
    "10010001", --  237 - 0xed  :  145 - 0x91
    "10010010", --  238 - 0xee  :  146 - 0x92
    "10010011", --  239 - 0xef  :  147 - 0x93
    "10010010", --  240 - 0xf0  :  146 - 0x92
    "10010011", --  241 - 0xf1  :  147 - 0x93
    "10010010", --  242 - 0xf2  :  146 - 0x92
    "10010001", --  243 - 0xf3  :  145 - 0x91
    "10010010", --  244 - 0xf4  :  146 - 0x92
    "10010001", --  245 - 0xf5  :  145 - 0x91
    "10010010", --  246 - 0xf6  :  146 - 0x92
    "10010011", --  247 - 0xf7  :  147 - 0x93
    "10010010", --  248 - 0xf8  :  146 - 0x92
    "10010011", --  249 - 0xf9  :  147 - 0x93
    "10010011", --  250 - 0xfa  :  147 - 0x93
    "10010010", --  251 - 0xfb  :  146 - 0x92
    "10010000", --  252 - 0xfc  :  144 - 0x90
    "10010001", --  253 - 0xfd  :  145 - 0x91
    "10100111", --  254 - 0xfe  :  167 - 0xa7
    "10100000", --  255 - 0xff  :  160 - 0xa0
    "10100000", --  256 - 0x100  :  160 - 0xa0 -- line 0x8
    "10100011", --  257 - 0x101  :  163 - 0xa3
    "10000010", --  258 - 0x102  :  130 - 0x82
    "10000011", --  259 - 0x103  :  131 - 0x83
    "10000101", --  260 - 0x104  :  133 - 0x85
    "10000110", --  261 - 0x105  :  134 - 0x86
    "10000101", --  262 - 0x106  :  133 - 0x85
    "10000110", --  263 - 0x107  :  134 - 0x86
    "10000101", --  264 - 0x108  :  133 - 0x85
    "10000110", --  265 - 0x109  :  134 - 0x86
    "10000101", --  266 - 0x10a  :  133 - 0x85
    "10000110", --  267 - 0x10b  :  134 - 0x86
    "10000100", --  268 - 0x10c  :  132 - 0x84
    "10000111", --  269 - 0x10d  :  135 - 0x87
    "10000110", --  270 - 0x10e  :  134 - 0x86
    "10000111", --  271 - 0x10f  :  135 - 0x87
    "10000100", --  272 - 0x110  :  132 - 0x84
    "10000101", --  273 - 0x111  :  133 - 0x85
    "10000101", --  274 - 0x112  :  133 - 0x85
    "10000110", --  275 - 0x113  :  134 - 0x86
    "10000101", --  276 - 0x114  :  133 - 0x85
    "10000110", --  277 - 0x115  :  134 - 0x86
    "10000110", --  278 - 0x116  :  134 - 0x86
    "10000111", --  279 - 0x117  :  135 - 0x87
    "10000110", --  280 - 0x118  :  134 - 0x86
    "10000111", --  281 - 0x119  :  135 - 0x87
    "10000100", --  282 - 0x11a  :  132 - 0x84
    "10000101", --  283 - 0x11b  :  133 - 0x85
    "10000010", --  284 - 0x11c  :  130 - 0x82
    "10000011", --  285 - 0x11d  :  131 - 0x83
    "10100111", --  286 - 0x11e  :  167 - 0xa7
    "10100000", --  287 - 0x11f  :  160 - 0xa0
    "10100000", --  288 - 0x120  :  160 - 0xa0 -- line 0x9
    "10100011", --  289 - 0x121  :  163 - 0xa3
    "10010010", --  290 - 0x122  :  146 - 0x92
    "10010011", --  291 - 0x123  :  147 - 0x93
    "10010111", --  292 - 0x124  :  151 - 0x97
    "10010100", --  293 - 0x125  :  148 - 0x94
    "10010111", --  294 - 0x126  :  151 - 0x97
    "10010100", --  295 - 0x127  :  148 - 0x94
    "10010111", --  296 - 0x128  :  151 - 0x97
    "10010100", --  297 - 0x129  :  148 - 0x94
    "10010111", --  298 - 0x12a  :  151 - 0x97
    "10010100", --  299 - 0x12b  :  148 - 0x94
    "10010110", --  300 - 0x12c  :  150 - 0x96
    "10010101", --  301 - 0x12d  :  149 - 0x95
    "10010110", --  302 - 0x12e  :  150 - 0x96
    "10010111", --  303 - 0x12f  :  151 - 0x97
    "10010100", --  304 - 0x130  :  148 - 0x94
    "10010101", --  305 - 0x131  :  149 - 0x95
    "10010111", --  306 - 0x132  :  151 - 0x97
    "10010100", --  307 - 0x133  :  148 - 0x94
    "10010111", --  308 - 0x134  :  151 - 0x97
    "10010100", --  309 - 0x135  :  148 - 0x94
    "10010110", --  310 - 0x136  :  150 - 0x96
    "10010111", --  311 - 0x137  :  151 - 0x97
    "10010110", --  312 - 0x138  :  150 - 0x96
    "10010111", --  313 - 0x139  :  151 - 0x97
    "10010100", --  314 - 0x13a  :  148 - 0x94
    "10010101", --  315 - 0x13b  :  149 - 0x95
    "10010010", --  316 - 0x13c  :  146 - 0x92
    "10010011", --  317 - 0x13d  :  147 - 0x93
    "10100111", --  318 - 0x13e  :  167 - 0xa7
    "10100000", --  319 - 0x13f  :  160 - 0xa0
    "10100000", --  320 - 0x140  :  160 - 0xa0 -- line 0xa
    "10100011", --  321 - 0x141  :  163 - 0xa3
    "10000000", --  322 - 0x142  :  128 - 0x80
    "10000010", --  323 - 0x143  :  130 - 0x82
    "10000100", --  324 - 0x144  :  132 - 0x84
    "10000111", --  325 - 0x145  :  135 - 0x87
    "10000101", --  326 - 0x146  :  133 - 0x85
    "10000110", --  327 - 0x147  :  134 - 0x86
    "10000100", --  328 - 0x148  :  132 - 0x84
    "10000111", --  329 - 0x149  :  135 - 0x87
    "10000100", --  330 - 0x14a  :  132 - 0x84
    "10000111", --  331 - 0x14b  :  135 - 0x87
    "10000110", --  332 - 0x14c  :  134 - 0x86
    "10000111", --  333 - 0x14d  :  135 - 0x87
    "10000100", --  334 - 0x14e  :  132 - 0x84
    "10000101", --  335 - 0x14f  :  133 - 0x85
    "10000100", --  336 - 0x150  :  132 - 0x84
    "10000101", --  337 - 0x151  :  133 - 0x85
    "10000110", --  338 - 0x152  :  134 - 0x86
    "10000111", --  339 - 0x153  :  135 - 0x87
    "10000100", --  340 - 0x154  :  132 - 0x84
    "10000101", --  341 - 0x155  :  133 - 0x85
    "10000101", --  342 - 0x156  :  133 - 0x85
    "10000110", --  343 - 0x157  :  134 - 0x86
    "10000100", --  344 - 0x158  :  132 - 0x84
    "10000111", --  345 - 0x159  :  135 - 0x87
    "10000100", --  346 - 0x15a  :  132 - 0x84
    "10000111", --  347 - 0x15b  :  135 - 0x87
    "10000000", --  348 - 0x15c  :  128 - 0x80
    "10000001", --  349 - 0x15d  :  129 - 0x81
    "10100111", --  350 - 0x15e  :  167 - 0xa7
    "10100000", --  351 - 0x15f  :  160 - 0xa0
    "10100000", --  352 - 0x160  :  160 - 0xa0 -- line 0xb
    "10100011", --  353 - 0x161  :  163 - 0xa3
    "10010010", --  354 - 0x162  :  146 - 0x92
    "10010001", --  355 - 0x163  :  145 - 0x91
    "10010110", --  356 - 0x164  :  150 - 0x96
    "10010101", --  357 - 0x165  :  149 - 0x95
    "10010111", --  358 - 0x166  :  151 - 0x97
    "10010100", --  359 - 0x167  :  148 - 0x94
    "10010110", --  360 - 0x168  :  150 - 0x96
    "10010101", --  361 - 0x169  :  149 - 0x95
    "10010110", --  362 - 0x16a  :  150 - 0x96
    "10010101", --  363 - 0x16b  :  149 - 0x95
    "10010110", --  364 - 0x16c  :  150 - 0x96
    "10010111", --  365 - 0x16d  :  151 - 0x97
    "10010100", --  366 - 0x16e  :  148 - 0x94
    "10010101", --  367 - 0x16f  :  149 - 0x95
    "10010100", --  368 - 0x170  :  148 - 0x94
    "10010101", --  369 - 0x171  :  149 - 0x95
    "10010110", --  370 - 0x172  :  150 - 0x96
    "10010111", --  371 - 0x173  :  151 - 0x97
    "10010100", --  372 - 0x174  :  148 - 0x94
    "10010101", --  373 - 0x175  :  149 - 0x95
    "10010111", --  374 - 0x176  :  151 - 0x97
    "10010100", --  375 - 0x177  :  148 - 0x94
    "10010110", --  376 - 0x178  :  150 - 0x96
    "10010101", --  377 - 0x179  :  149 - 0x95
    "10010110", --  378 - 0x17a  :  150 - 0x96
    "10010101", --  379 - 0x17b  :  149 - 0x95
    "10010000", --  380 - 0x17c  :  144 - 0x90
    "10010001", --  381 - 0x17d  :  145 - 0x91
    "10100111", --  382 - 0x17e  :  167 - 0xa7
    "10100000", --  383 - 0x17f  :  160 - 0xa0
    "10100000", --  384 - 0x180  :  160 - 0xa0 -- line 0xc
    "10100011", --  385 - 0x181  :  163 - 0xa3
    "10000010", --  386 - 0x182  :  130 - 0x82
    "10000011", --  387 - 0x183  :  131 - 0x83
    "10000110", --  388 - 0x184  :  134 - 0x86
    "10000111", --  389 - 0x185  :  135 - 0x87
    "10000100", --  390 - 0x186  :  132 - 0x84
    "10000101", --  391 - 0x187  :  133 - 0x85
    "10000100", --  392 - 0x188  :  132 - 0x84
    "10000111", --  393 - 0x189  :  135 - 0x87
    "10000100", --  394 - 0x18a  :  132 - 0x84
    "10000111", --  395 - 0x18b  :  135 - 0x87
    "10000110", --  396 - 0x18c  :  134 - 0x86
    "10000111", --  397 - 0x18d  :  135 - 0x87
    "10000100", --  398 - 0x18e  :  132 - 0x84
    "10000111", --  399 - 0x18f  :  135 - 0x87
    "10000110", --  400 - 0x190  :  134 - 0x86
    "10000111", --  401 - 0x191  :  135 - 0x87
    "10000110", --  402 - 0x192  :  134 - 0x86
    "10000111", --  403 - 0x193  :  135 - 0x87
    "10000110", --  404 - 0x194  :  134 - 0x86
    "10000111", --  405 - 0x195  :  135 - 0x87
    "10000110", --  406 - 0x196  :  134 - 0x86
    "10000111", --  407 - 0x197  :  135 - 0x87
    "10000101", --  408 - 0x198  :  133 - 0x85
    "10000110", --  409 - 0x199  :  134 - 0x86
    "10000100", --  410 - 0x19a  :  132 - 0x84
    "10000111", --  411 - 0x19b  :  135 - 0x87
    "10000000", --  412 - 0x19c  :  128 - 0x80
    "10000010", --  413 - 0x19d  :  130 - 0x82
    "10100111", --  414 - 0x19e  :  167 - 0xa7
    "10100000", --  415 - 0x19f  :  160 - 0xa0
    "10100000", --  416 - 0x1a0  :  160 - 0xa0 -- line 0xd
    "10100011", --  417 - 0x1a1  :  163 - 0xa3
    "10010010", --  418 - 0x1a2  :  146 - 0x92
    "10010011", --  419 - 0x1a3  :  147 - 0x93
    "10010110", --  420 - 0x1a4  :  150 - 0x96
    "10010111", --  421 - 0x1a5  :  151 - 0x97
    "10010100", --  422 - 0x1a6  :  148 - 0x94
    "10010101", --  423 - 0x1a7  :  149 - 0x95
    "10010110", --  424 - 0x1a8  :  150 - 0x96
    "10010101", --  425 - 0x1a9  :  149 - 0x95
    "10010110", --  426 - 0x1aa  :  150 - 0x96
    "10010101", --  427 - 0x1ab  :  149 - 0x95
    "10010110", --  428 - 0x1ac  :  150 - 0x96
    "10010111", --  429 - 0x1ad  :  151 - 0x97
    "10010110", --  430 - 0x1ae  :  150 - 0x96
    "10010101", --  431 - 0x1af  :  149 - 0x95
    "10010110", --  432 - 0x1b0  :  150 - 0x96
    "10010111", --  433 - 0x1b1  :  151 - 0x97
    "10010110", --  434 - 0x1b2  :  150 - 0x96
    "10010111", --  435 - 0x1b3  :  151 - 0x97
    "10010110", --  436 - 0x1b4  :  150 - 0x96
    "10010111", --  437 - 0x1b5  :  151 - 0x97
    "10010110", --  438 - 0x1b6  :  150 - 0x96
    "10010111", --  439 - 0x1b7  :  151 - 0x97
    "10010111", --  440 - 0x1b8  :  151 - 0x97
    "10010100", --  441 - 0x1b9  :  148 - 0x94
    "10010110", --  442 - 0x1ba  :  150 - 0x96
    "10010101", --  443 - 0x1bb  :  149 - 0x95
    "10010010", --  444 - 0x1bc  :  146 - 0x92
    "10010001", --  445 - 0x1bd  :  145 - 0x91
    "10100111", --  446 - 0x1be  :  167 - 0xa7
    "10100000", --  447 - 0x1bf  :  160 - 0xa0
    "10100000", --  448 - 0x1c0  :  160 - 0xa0 -- line 0xe
    "10100011", --  449 - 0x1c1  :  163 - 0xa3
    "10000000", --  450 - 0x1c2  :  128 - 0x80
    "10000001", --  451 - 0x1c3  :  129 - 0x81
    "10000101", --  452 - 0x1c4  :  133 - 0x85
    "10000110", --  453 - 0x1c5  :  134 - 0x86
    "10000100", --  454 - 0x1c6  :  132 - 0x84
    "10000101", --  455 - 0x1c7  :  133 - 0x85
    "10000100", --  456 - 0x1c8  :  132 - 0x84
    "10000101", --  457 - 0x1c9  :  133 - 0x85
    "10000100", --  458 - 0x1ca  :  132 - 0x84
    "10000111", --  459 - 0x1cb  :  135 - 0x87
    "10000001", --  460 - 0x1cc  :  129 - 0x81
    "10000000", --  461 - 0x1cd  :  128 - 0x80
    "10000010", --  462 - 0x1ce  :  130 - 0x82
    "10000011", --  463 - 0x1cf  :  131 - 0x83
    "10000010", --  464 - 0x1d0  :  130 - 0x82
    "10000011", --  465 - 0x1d1  :  131 - 0x83
    "10000001", --  466 - 0x1d2  :  129 - 0x81
    "10000000", --  467 - 0x1d3  :  128 - 0x80
    "10000101", --  468 - 0x1d4  :  133 - 0x85
    "10000110", --  469 - 0x1d5  :  134 - 0x86
    "10000110", --  470 - 0x1d6  :  134 - 0x86
    "10000111", --  471 - 0x1d7  :  135 - 0x87
    "10000100", --  472 - 0x1d8  :  132 - 0x84
    "10000111", --  473 - 0x1d9  :  135 - 0x87
    "10000100", --  474 - 0x1da  :  132 - 0x84
    "10000111", --  475 - 0x1db  :  135 - 0x87
    "10000000", --  476 - 0x1dc  :  128 - 0x80
    "10000001", --  477 - 0x1dd  :  129 - 0x81
    "10100111", --  478 - 0x1de  :  167 - 0xa7
    "10100000", --  479 - 0x1df  :  160 - 0xa0
    "10100000", --  480 - 0x1e0  :  160 - 0xa0 -- line 0xf
    "10100011", --  481 - 0x1e1  :  163 - 0xa3
    "10010000", --  482 - 0x1e2  :  144 - 0x90
    "10010001", --  483 - 0x1e3  :  145 - 0x91
    "10010111", --  484 - 0x1e4  :  151 - 0x97
    "10010100", --  485 - 0x1e5  :  148 - 0x94
    "10010100", --  486 - 0x1e6  :  148 - 0x94
    "10010101", --  487 - 0x1e7  :  149 - 0x95
    "10010100", --  488 - 0x1e8  :  148 - 0x94
    "10010101", --  489 - 0x1e9  :  149 - 0x95
    "10010110", --  490 - 0x1ea  :  150 - 0x96
    "10010101", --  491 - 0x1eb  :  149 - 0x95
    "10010011", --  492 - 0x1ec  :  147 - 0x93
    "10010010", --  493 - 0x1ed  :  146 - 0x92
    "10010010", --  494 - 0x1ee  :  146 - 0x92
    "10010011", --  495 - 0x1ef  :  147 - 0x93
    "10010010", --  496 - 0x1f0  :  146 - 0x92
    "10010011", --  497 - 0x1f1  :  147 - 0x93
    "10010011", --  498 - 0x1f2  :  147 - 0x93
    "10010010", --  499 - 0x1f3  :  146 - 0x92
    "10010111", --  500 - 0x1f4  :  151 - 0x97
    "10010100", --  501 - 0x1f5  :  148 - 0x94
    "10010110", --  502 - 0x1f6  :  150 - 0x96
    "10010111", --  503 - 0x1f7  :  151 - 0x97
    "10010110", --  504 - 0x1f8  :  150 - 0x96
    "10010101", --  505 - 0x1f9  :  149 - 0x95
    "10010110", --  506 - 0x1fa  :  150 - 0x96
    "10010101", --  507 - 0x1fb  :  149 - 0x95
    "10010000", --  508 - 0x1fc  :  144 - 0x90
    "10010001", --  509 - 0x1fd  :  145 - 0x91
    "10100111", --  510 - 0x1fe  :  167 - 0xa7
    "10100000", --  511 - 0x1ff  :  160 - 0xa0
    "10100000", --  512 - 0x200  :  160 - 0xa0 -- line 0x10
    "10100011", --  513 - 0x201  :  163 - 0xa3
    "10000010", --  514 - 0x202  :  130 - 0x82
    "10000011", --  515 - 0x203  :  131 - 0x83
    "10000101", --  516 - 0x204  :  133 - 0x85
    "10000110", --  517 - 0x205  :  134 - 0x86
    "10000101", --  518 - 0x206  :  133 - 0x85
    "10000110", --  519 - 0x207  :  134 - 0x86
    "10000101", --  520 - 0x208  :  133 - 0x85
    "10000110", --  521 - 0x209  :  134 - 0x86
    "10000101", --  522 - 0x20a  :  133 - 0x85
    "10000110", --  523 - 0x20b  :  134 - 0x86
    "10000000", --  524 - 0x20c  :  128 - 0x80
    "10000010", --  525 - 0x20d  :  130 - 0x82
    "10000010", --  526 - 0x20e  :  130 - 0x82
    "10000011", --  527 - 0x20f  :  131 - 0x83
    "10000000", --  528 - 0x210  :  128 - 0x80
    "10000001", --  529 - 0x211  :  129 - 0x81
    "10000001", --  530 - 0x212  :  129 - 0x81
    "10000000", --  531 - 0x213  :  128 - 0x80
    "10000101", --  532 - 0x214  :  133 - 0x85
    "10000110", --  533 - 0x215  :  134 - 0x86
    "10000110", --  534 - 0x216  :  134 - 0x86
    "10000111", --  535 - 0x217  :  135 - 0x87
    "10000110", --  536 - 0x218  :  134 - 0x86
    "10000111", --  537 - 0x219  :  135 - 0x87
    "10000100", --  538 - 0x21a  :  132 - 0x84
    "10000101", --  539 - 0x21b  :  133 - 0x85
    "10000010", --  540 - 0x21c  :  130 - 0x82
    "10000011", --  541 - 0x21d  :  131 - 0x83
    "10100111", --  542 - 0x21e  :  167 - 0xa7
    "10100000", --  543 - 0x21f  :  160 - 0xa0
    "10100000", --  544 - 0x220  :  160 - 0xa0 -- line 0x11
    "10100011", --  545 - 0x221  :  163 - 0xa3
    "10010010", --  546 - 0x222  :  146 - 0x92
    "10010011", --  547 - 0x223  :  147 - 0x93
    "10010111", --  548 - 0x224  :  151 - 0x97
    "10010100", --  549 - 0x225  :  148 - 0x94
    "10010111", --  550 - 0x226  :  151 - 0x97
    "10010100", --  551 - 0x227  :  148 - 0x94
    "10010111", --  552 - 0x228  :  151 - 0x97
    "10010100", --  553 - 0x229  :  148 - 0x94
    "10010111", --  554 - 0x22a  :  151 - 0x97
    "10010100", --  555 - 0x22b  :  148 - 0x94
    "10010010", --  556 - 0x22c  :  146 - 0x92
    "10010001", --  557 - 0x22d  :  145 - 0x91
    "10010010", --  558 - 0x22e  :  146 - 0x92
    "10010011", --  559 - 0x22f  :  147 - 0x93
    "10010000", --  560 - 0x230  :  144 - 0x90
    "10010001", --  561 - 0x231  :  145 - 0x91
    "10010011", --  562 - 0x232  :  147 - 0x93
    "10010010", --  563 - 0x233  :  146 - 0x92
    "10010111", --  564 - 0x234  :  151 - 0x97
    "10010100", --  565 - 0x235  :  148 - 0x94
    "10010110", --  566 - 0x236  :  150 - 0x96
    "10010111", --  567 - 0x237  :  151 - 0x97
    "10010110", --  568 - 0x238  :  150 - 0x96
    "10010111", --  569 - 0x239  :  151 - 0x97
    "10010100", --  570 - 0x23a  :  148 - 0x94
    "10010101", --  571 - 0x23b  :  149 - 0x95
    "10010010", --  572 - 0x23c  :  146 - 0x92
    "10010011", --  573 - 0x23d  :  147 - 0x93
    "10100111", --  574 - 0x23e  :  167 - 0xa7
    "10100000", --  575 - 0x23f  :  160 - 0xa0
    "10100000", --  576 - 0x240  :  160 - 0xa0 -- line 0x12
    "10100011", --  577 - 0x241  :  163 - 0xa3
    "10000000", --  578 - 0x242  :  128 - 0x80
    "10000010", --  579 - 0x243  :  130 - 0x82
    "10000100", --  580 - 0x244  :  132 - 0x84
    "10000111", --  581 - 0x245  :  135 - 0x87
    "10000101", --  582 - 0x246  :  133 - 0x85
    "10000110", --  583 - 0x247  :  134 - 0x86
    "10000100", --  584 - 0x248  :  132 - 0x84
    "10000111", --  585 - 0x249  :  135 - 0x87
    "10000100", --  586 - 0x24a  :  132 - 0x84
    "10000111", --  587 - 0x24b  :  135 - 0x87
    "10000010", --  588 - 0x24c  :  130 - 0x82
    "10000011", --  589 - 0x24d  :  131 - 0x83
    "10000000", --  590 - 0x24e  :  128 - 0x80
    "10000001", --  591 - 0x24f  :  129 - 0x81
    "10000000", --  592 - 0x250  :  128 - 0x80
    "10000001", --  593 - 0x251  :  129 - 0x81
    "10000010", --  594 - 0x252  :  130 - 0x82
    "10000011", --  595 - 0x253  :  131 - 0x83
    "10000100", --  596 - 0x254  :  132 - 0x84
    "10000101", --  597 - 0x255  :  133 - 0x85
    "10000101", --  598 - 0x256  :  133 - 0x85
    "10000110", --  599 - 0x257  :  134 - 0x86
    "10000100", --  600 - 0x258  :  132 - 0x84
    "10000111", --  601 - 0x259  :  135 - 0x87
    "10000100", --  602 - 0x25a  :  132 - 0x84
    "10000111", --  603 - 0x25b  :  135 - 0x87
    "10000000", --  604 - 0x25c  :  128 - 0x80
    "10000001", --  605 - 0x25d  :  129 - 0x81
    "10100111", --  606 - 0x25e  :  167 - 0xa7
    "10100000", --  607 - 0x25f  :  160 - 0xa0
    "10100000", --  608 - 0x260  :  160 - 0xa0 -- line 0x13
    "10100011", --  609 - 0x261  :  163 - 0xa3
    "10010010", --  610 - 0x262  :  146 - 0x92
    "10010001", --  611 - 0x263  :  145 - 0x91
    "10010110", --  612 - 0x264  :  150 - 0x96
    "10010101", --  613 - 0x265  :  149 - 0x95
    "10010111", --  614 - 0x266  :  151 - 0x97
    "10010100", --  615 - 0x267  :  148 - 0x94
    "10010110", --  616 - 0x268  :  150 - 0x96
    "10010101", --  617 - 0x269  :  149 - 0x95
    "10010110", --  618 - 0x26a  :  150 - 0x96
    "10010101", --  619 - 0x26b  :  149 - 0x95
    "10010010", --  620 - 0x26c  :  146 - 0x92
    "10010011", --  621 - 0x26d  :  147 - 0x93
    "10010000", --  622 - 0x26e  :  144 - 0x90
    "10010001", --  623 - 0x26f  :  145 - 0x91
    "10010000", --  624 - 0x270  :  144 - 0x90
    "10010001", --  625 - 0x271  :  145 - 0x91
    "10010010", --  626 - 0x272  :  146 - 0x92
    "10010011", --  627 - 0x273  :  147 - 0x93
    "10010100", --  628 - 0x274  :  148 - 0x94
    "10010101", --  629 - 0x275  :  149 - 0x95
    "10010111", --  630 - 0x276  :  151 - 0x97
    "10010100", --  631 - 0x277  :  148 - 0x94
    "10010110", --  632 - 0x278  :  150 - 0x96
    "10010101", --  633 - 0x279  :  149 - 0x95
    "10010110", --  634 - 0x27a  :  150 - 0x96
    "10010101", --  635 - 0x27b  :  149 - 0x95
    "10010000", --  636 - 0x27c  :  144 - 0x90
    "10010001", --  637 - 0x27d  :  145 - 0x91
    "10100111", --  638 - 0x27e  :  167 - 0xa7
    "10100000", --  639 - 0x27f  :  160 - 0xa0
    "10100000", --  640 - 0x280  :  160 - 0xa0 -- line 0x14
    "10100011", --  641 - 0x281  :  163 - 0xa3
    "10000010", --  642 - 0x282  :  130 - 0x82
    "10000011", --  643 - 0x283  :  131 - 0x83
    "10000110", --  644 - 0x284  :  134 - 0x86
    "10000111", --  645 - 0x285  :  135 - 0x87
    "10000100", --  646 - 0x286  :  132 - 0x84
    "10000101", --  647 - 0x287  :  133 - 0x85
    "10000100", --  648 - 0x288  :  132 - 0x84
    "10000111", --  649 - 0x289  :  135 - 0x87
    "10000100", --  650 - 0x28a  :  132 - 0x84
    "10000111", --  651 - 0x28b  :  135 - 0x87
    "10000110", --  652 - 0x28c  :  134 - 0x86
    "10000111", --  653 - 0x28d  :  135 - 0x87
    "10000100", --  654 - 0x28e  :  132 - 0x84
    "10000111", --  655 - 0x28f  :  135 - 0x87
    "10000110", --  656 - 0x290  :  134 - 0x86
    "10000111", --  657 - 0x291  :  135 - 0x87
    "10000110", --  658 - 0x292  :  134 - 0x86
    "10000111", --  659 - 0x293  :  135 - 0x87
    "10000110", --  660 - 0x294  :  134 - 0x86
    "10000111", --  661 - 0x295  :  135 - 0x87
    "10000110", --  662 - 0x296  :  134 - 0x86
    "10000111", --  663 - 0x297  :  135 - 0x87
    "10000101", --  664 - 0x298  :  133 - 0x85
    "10000110", --  665 - 0x299  :  134 - 0x86
    "10000100", --  666 - 0x29a  :  132 - 0x84
    "10000111", --  667 - 0x29b  :  135 - 0x87
    "10000000", --  668 - 0x29c  :  128 - 0x80
    "10000010", --  669 - 0x29d  :  130 - 0x82
    "10100111", --  670 - 0x29e  :  167 - 0xa7
    "10100000", --  671 - 0x29f  :  160 - 0xa0
    "10100000", --  672 - 0x2a0  :  160 - 0xa0 -- line 0x15
    "10100011", --  673 - 0x2a1  :  163 - 0xa3
    "10010010", --  674 - 0x2a2  :  146 - 0x92
    "10010011", --  675 - 0x2a3  :  147 - 0x93
    "10010110", --  676 - 0x2a4  :  150 - 0x96
    "10010111", --  677 - 0x2a5  :  151 - 0x97
    "10010100", --  678 - 0x2a6  :  148 - 0x94
    "10010101", --  679 - 0x2a7  :  149 - 0x95
    "10010110", --  680 - 0x2a8  :  150 - 0x96
    "10010101", --  681 - 0x2a9  :  149 - 0x95
    "10010110", --  682 - 0x2aa  :  150 - 0x96
    "10010101", --  683 - 0x2ab  :  149 - 0x95
    "10010110", --  684 - 0x2ac  :  150 - 0x96
    "10010111", --  685 - 0x2ad  :  151 - 0x97
    "10010110", --  686 - 0x2ae  :  150 - 0x96
    "10010101", --  687 - 0x2af  :  149 - 0x95
    "10010110", --  688 - 0x2b0  :  150 - 0x96
    "10010111", --  689 - 0x2b1  :  151 - 0x97
    "10010110", --  690 - 0x2b2  :  150 - 0x96
    "10010111", --  691 - 0x2b3  :  151 - 0x97
    "10010110", --  692 - 0x2b4  :  150 - 0x96
    "10010111", --  693 - 0x2b5  :  151 - 0x97
    "10010110", --  694 - 0x2b6  :  150 - 0x96
    "10010111", --  695 - 0x2b7  :  151 - 0x97
    "10010111", --  696 - 0x2b8  :  151 - 0x97
    "10010100", --  697 - 0x2b9  :  148 - 0x94
    "10010110", --  698 - 0x2ba  :  150 - 0x96
    "10010101", --  699 - 0x2bb  :  149 - 0x95
    "10010010", --  700 - 0x2bc  :  146 - 0x92
    "10010001", --  701 - 0x2bd  :  145 - 0x91
    "10100111", --  702 - 0x2be  :  167 - 0xa7
    "10100000", --  703 - 0x2bf  :  160 - 0xa0
    "10100000", --  704 - 0x2c0  :  160 - 0xa0 -- line 0x16
    "10100011", --  705 - 0x2c1  :  163 - 0xa3
    "10000000", --  706 - 0x2c2  :  128 - 0x80
    "10000001", --  707 - 0x2c3  :  129 - 0x81
    "10000101", --  708 - 0x2c4  :  133 - 0x85
    "10000110", --  709 - 0x2c5  :  134 - 0x86
    "10000100", --  710 - 0x2c6  :  132 - 0x84
    "10000101", --  711 - 0x2c7  :  133 - 0x85
    "10000100", --  712 - 0x2c8  :  132 - 0x84
    "10000101", --  713 - 0x2c9  :  133 - 0x85
    "10000100", --  714 - 0x2ca  :  132 - 0x84
    "10000111", --  715 - 0x2cb  :  135 - 0x87
    "10000101", --  716 - 0x2cc  :  133 - 0x85
    "10000110", --  717 - 0x2cd  :  134 - 0x86
    "10000110", --  718 - 0x2ce  :  134 - 0x86
    "10000111", --  719 - 0x2cf  :  135 - 0x87
    "10000110", --  720 - 0x2d0  :  134 - 0x86
    "10000111", --  721 - 0x2d1  :  135 - 0x87
    "10000101", --  722 - 0x2d2  :  133 - 0x85
    "10000110", --  723 - 0x2d3  :  134 - 0x86
    "10000101", --  724 - 0x2d4  :  133 - 0x85
    "10000110", --  725 - 0x2d5  :  134 - 0x86
    "10000110", --  726 - 0x2d6  :  134 - 0x86
    "10000111", --  727 - 0x2d7  :  135 - 0x87
    "10000100", --  728 - 0x2d8  :  132 - 0x84
    "10000111", --  729 - 0x2d9  :  135 - 0x87
    "10000100", --  730 - 0x2da  :  132 - 0x84
    "10000111", --  731 - 0x2db  :  135 - 0x87
    "10000000", --  732 - 0x2dc  :  128 - 0x80
    "10000001", --  733 - 0x2dd  :  129 - 0x81
    "10100111", --  734 - 0x2de  :  167 - 0xa7
    "10100000", --  735 - 0x2df  :  160 - 0xa0
    "10100000", --  736 - 0x2e0  :  160 - 0xa0 -- line 0x17
    "10100011", --  737 - 0x2e1  :  163 - 0xa3
    "10010000", --  738 - 0x2e2  :  144 - 0x90
    "10010001", --  739 - 0x2e3  :  145 - 0x91
    "10010111", --  740 - 0x2e4  :  151 - 0x97
    "10010100", --  741 - 0x2e5  :  148 - 0x94
    "10010100", --  742 - 0x2e6  :  148 - 0x94
    "10010101", --  743 - 0x2e7  :  149 - 0x95
    "10010100", --  744 - 0x2e8  :  148 - 0x94
    "10010101", --  745 - 0x2e9  :  149 - 0x95
    "10010110", --  746 - 0x2ea  :  150 - 0x96
    "10010101", --  747 - 0x2eb  :  149 - 0x95
    "10010111", --  748 - 0x2ec  :  151 - 0x97
    "10010100", --  749 - 0x2ed  :  148 - 0x94
    "10010110", --  750 - 0x2ee  :  150 - 0x96
    "10010111", --  751 - 0x2ef  :  151 - 0x97
    "10010110", --  752 - 0x2f0  :  150 - 0x96
    "10010111", --  753 - 0x2f1  :  151 - 0x97
    "10010111", --  754 - 0x2f2  :  151 - 0x97
    "10010100", --  755 - 0x2f3  :  148 - 0x94
    "10010111", --  756 - 0x2f4  :  151 - 0x97
    "10010100", --  757 - 0x2f5  :  148 - 0x94
    "10010110", --  758 - 0x2f6  :  150 - 0x96
    "10010111", --  759 - 0x2f7  :  151 - 0x97
    "10010110", --  760 - 0x2f8  :  150 - 0x96
    "10010101", --  761 - 0x2f9  :  149 - 0x95
    "10010110", --  762 - 0x2fa  :  150 - 0x96
    "10010101", --  763 - 0x2fb  :  149 - 0x95
    "10010000", --  764 - 0x2fc  :  144 - 0x90
    "10010001", --  765 - 0x2fd  :  145 - 0x91
    "10100111", --  766 - 0x2fe  :  167 - 0xa7
    "10100000", --  767 - 0x2ff  :  160 - 0xa0
    "10100000", --  768 - 0x300  :  160 - 0xa0 -- line 0x18
    "10100011", --  769 - 0x301  :  163 - 0xa3
    "10000000", --  770 - 0x302  :  128 - 0x80
    "10000010", --  771 - 0x303  :  130 - 0x82
    "10000100", --  772 - 0x304  :  132 - 0x84
    "10000111", --  773 - 0x305  :  135 - 0x87
    "10000100", --  774 - 0x306  :  132 - 0x84
    "10000111", --  775 - 0x307  :  135 - 0x87
    "10000100", --  776 - 0x308  :  132 - 0x84
    "10000111", --  777 - 0x309  :  135 - 0x87
    "10000110", --  778 - 0x30a  :  134 - 0x86
    "10000111", --  779 - 0x30b  :  135 - 0x87
    "10000101", --  780 - 0x30c  :  133 - 0x85
    "10000110", --  781 - 0x30d  :  134 - 0x86
    "10000100", --  782 - 0x30e  :  132 - 0x84
    "10000111", --  783 - 0x30f  :  135 - 0x87
    "10000100", --  784 - 0x310  :  132 - 0x84
    "10000101", --  785 - 0x311  :  133 - 0x85
    "10000100", --  786 - 0x312  :  132 - 0x84
    "10000111", --  787 - 0x313  :  135 - 0x87
    "10000110", --  788 - 0x314  :  134 - 0x86
    "10000111", --  789 - 0x315  :  135 - 0x87
    "10000110", --  790 - 0x316  :  134 - 0x86
    "10000111", --  791 - 0x317  :  135 - 0x87
    "10000100", --  792 - 0x318  :  132 - 0x84
    "10000111", --  793 - 0x319  :  135 - 0x87
    "10000101", --  794 - 0x31a  :  133 - 0x85
    "10000110", --  795 - 0x31b  :  134 - 0x86
    "10000000", --  796 - 0x31c  :  128 - 0x80
    "10000010", --  797 - 0x31d  :  130 - 0x82
    "10100111", --  798 - 0x31e  :  167 - 0xa7
    "10100000", --  799 - 0x31f  :  160 - 0xa0
    "10100000", --  800 - 0x320  :  160 - 0xa0 -- line 0x19
    "10100011", --  801 - 0x321  :  163 - 0xa3
    "10010010", --  802 - 0x322  :  146 - 0x92
    "10010001", --  803 - 0x323  :  145 - 0x91
    "10010110", --  804 - 0x324  :  150 - 0x96
    "10010101", --  805 - 0x325  :  149 - 0x95
    "10010110", --  806 - 0x326  :  150 - 0x96
    "10010101", --  807 - 0x327  :  149 - 0x95
    "10010110", --  808 - 0x328  :  150 - 0x96
    "10010101", --  809 - 0x329  :  149 - 0x95
    "10010110", --  810 - 0x32a  :  150 - 0x96
    "10010111", --  811 - 0x32b  :  151 - 0x97
    "10010111", --  812 - 0x32c  :  151 - 0x97
    "10010100", --  813 - 0x32d  :  148 - 0x94
    "10010110", --  814 - 0x32e  :  150 - 0x96
    "10010101", --  815 - 0x32f  :  149 - 0x95
    "10010100", --  816 - 0x330  :  148 - 0x94
    "10010101", --  817 - 0x331  :  149 - 0x95
    "10010110", --  818 - 0x332  :  150 - 0x96
    "10010101", --  819 - 0x333  :  149 - 0x95
    "10010110", --  820 - 0x334  :  150 - 0x96
    "10010111", --  821 - 0x335  :  151 - 0x97
    "10010110", --  822 - 0x336  :  150 - 0x96
    "10010111", --  823 - 0x337  :  151 - 0x97
    "10010110", --  824 - 0x338  :  150 - 0x96
    "10010101", --  825 - 0x339  :  149 - 0x95
    "10010111", --  826 - 0x33a  :  151 - 0x97
    "10010100", --  827 - 0x33b  :  148 - 0x94
    "10010010", --  828 - 0x33c  :  146 - 0x92
    "10010001", --  829 - 0x33d  :  145 - 0x91
    "10100111", --  830 - 0x33e  :  167 - 0xa7
    "10100000", --  831 - 0x33f  :  160 - 0xa0
    "10100000", --  832 - 0x340  :  160 - 0xa0 -- line 0x1a
    "10100011", --  833 - 0x341  :  163 - 0xa3
    "10000001", --  834 - 0x342  :  129 - 0x81
    "10000000", --  835 - 0x343  :  128 - 0x80
    "10000000", --  836 - 0x344  :  128 - 0x80
    "10000001", --  837 - 0x345  :  129 - 0x81
    "10000010", --  838 - 0x346  :  130 - 0x82
    "10000011", --  839 - 0x347  :  131 - 0x83
    "10000001", --  840 - 0x348  :  129 - 0x81
    "10000000", --  841 - 0x349  :  128 - 0x80
    "10000001", --  842 - 0x34a  :  129 - 0x81
    "10000000", --  843 - 0x34b  :  128 - 0x80
    "10000000", --  844 - 0x34c  :  128 - 0x80
    "10000010", --  845 - 0x34d  :  130 - 0x82
    "10000000", --  846 - 0x34e  :  128 - 0x80
    "10000001", --  847 - 0x34f  :  129 - 0x81
    "10000001", --  848 - 0x350  :  129 - 0x81
    "10000000", --  849 - 0x351  :  128 - 0x80
    "10000000", --  850 - 0x352  :  128 - 0x80
    "10000010", --  851 - 0x353  :  130 - 0x82
    "10000000", --  852 - 0x354  :  128 - 0x80
    "10000001", --  853 - 0x355  :  129 - 0x81
    "10000010", --  854 - 0x356  :  130 - 0x82
    "10000011", --  855 - 0x357  :  131 - 0x83
    "10000001", --  856 - 0x358  :  129 - 0x81
    "10000000", --  857 - 0x359  :  128 - 0x80
    "10000000", --  858 - 0x35a  :  128 - 0x80
    "10000001", --  859 - 0x35b  :  129 - 0x81
    "10000000", --  860 - 0x35c  :  128 - 0x80
    "10000001", --  861 - 0x35d  :  129 - 0x81
    "10100111", --  862 - 0x35e  :  167 - 0xa7
    "10100000", --  863 - 0x35f  :  160 - 0xa0
    "10100000", --  864 - 0x360  :  160 - 0xa0 -- line 0x1b
    "10100011", --  865 - 0x361  :  163 - 0xa3
    "10010011", --  866 - 0x362  :  147 - 0x93
    "10010010", --  867 - 0x363  :  146 - 0x92
    "10010000", --  868 - 0x364  :  144 - 0x90
    "10010001", --  869 - 0x365  :  145 - 0x91
    "10010010", --  870 - 0x366  :  146 - 0x92
    "10010011", --  871 - 0x367  :  147 - 0x93
    "10010011", --  872 - 0x368  :  147 - 0x93
    "10010010", --  873 - 0x369  :  146 - 0x92
    "10010011", --  874 - 0x36a  :  147 - 0x93
    "10010010", --  875 - 0x36b  :  146 - 0x92
    "10010010", --  876 - 0x36c  :  146 - 0x92
    "10010001", --  877 - 0x36d  :  145 - 0x91
    "10010000", --  878 - 0x36e  :  144 - 0x90
    "10010001", --  879 - 0x36f  :  145 - 0x91
    "10010011", --  880 - 0x370  :  147 - 0x93
    "10010010", --  881 - 0x371  :  146 - 0x92
    "10010010", --  882 - 0x372  :  146 - 0x92
    "10010001", --  883 - 0x373  :  145 - 0x91
    "10010000", --  884 - 0x374  :  144 - 0x90
    "10010001", --  885 - 0x375  :  145 - 0x91
    "10010010", --  886 - 0x376  :  146 - 0x92
    "10010011", --  887 - 0x377  :  147 - 0x93
    "10010011", --  888 - 0x378  :  147 - 0x93
    "10010010", --  889 - 0x379  :  146 - 0x92
    "10010000", --  890 - 0x37a  :  144 - 0x90
    "10010001", --  891 - 0x37b  :  145 - 0x91
    "10010000", --  892 - 0x37c  :  144 - 0x90
    "10010001", --  893 - 0x37d  :  145 - 0x91
    "10100111", --  894 - 0x37e  :  167 - 0xa7
    "10100000", --  895 - 0x37f  :  160 - 0xa0
    "10100000", --  896 - 0x380  :  160 - 0xa0 -- line 0x1c
    "10100100", --  897 - 0x381  :  164 - 0xa4
    "10100101", --  898 - 0x382  :  165 - 0xa5
    "10100101", --  899 - 0x383  :  165 - 0xa5
    "10100101", --  900 - 0x384  :  165 - 0xa5
    "10100101", --  901 - 0x385  :  165 - 0xa5
    "10100101", --  902 - 0x386  :  165 - 0xa5
    "10100101", --  903 - 0x387  :  165 - 0xa5
    "10100101", --  904 - 0x388  :  165 - 0xa5
    "10100101", --  905 - 0x389  :  165 - 0xa5
    "10100101", --  906 - 0x38a  :  165 - 0xa5
    "10100101", --  907 - 0x38b  :  165 - 0xa5
    "10100101", --  908 - 0x38c  :  165 - 0xa5
    "10100101", --  909 - 0x38d  :  165 - 0xa5
    "10100101", --  910 - 0x38e  :  165 - 0xa5
    "10100101", --  911 - 0x38f  :  165 - 0xa5
    "10100101", --  912 - 0x390  :  165 - 0xa5
    "10100101", --  913 - 0x391  :  165 - 0xa5
    "10100101", --  914 - 0x392  :  165 - 0xa5
    "10100101", --  915 - 0x393  :  165 - 0xa5
    "10100101", --  916 - 0x394  :  165 - 0xa5
    "10100101", --  917 - 0x395  :  165 - 0xa5
    "10100101", --  918 - 0x396  :  165 - 0xa5
    "10100101", --  919 - 0x397  :  165 - 0xa5
    "10100101", --  920 - 0x398  :  165 - 0xa5
    "10100101", --  921 - 0x399  :  165 - 0xa5
    "10100101", --  922 - 0x39a  :  165 - 0xa5
    "10100101", --  923 - 0x39b  :  165 - 0xa5
    "10100101", --  924 - 0x39c  :  165 - 0xa5
    "10100101", --  925 - 0x39d  :  165 - 0xa5
    "10101000", --  926 - 0x39e  :  168 - 0xa8
    "10100000", --  927 - 0x39f  :  160 - 0xa0
    "10100000", --  928 - 0x3a0  :  160 - 0xa0 -- line 0x1d
    "10100000", --  929 - 0x3a1  :  160 - 0xa0
    "10100000", --  930 - 0x3a2  :  160 - 0xa0
    "10100000", --  931 - 0x3a3  :  160 - 0xa0
    "10100000", --  932 - 0x3a4  :  160 - 0xa0
    "10100000", --  933 - 0x3a5  :  160 - 0xa0
    "10100000", --  934 - 0x3a6  :  160 - 0xa0
    "10100000", --  935 - 0x3a7  :  160 - 0xa0
    "10100000", --  936 - 0x3a8  :  160 - 0xa0
    "10100000", --  937 - 0x3a9  :  160 - 0xa0
    "10100000", --  938 - 0x3aa  :  160 - 0xa0
    "10100000", --  939 - 0x3ab  :  160 - 0xa0
    "10100000", --  940 - 0x3ac  :  160 - 0xa0
    "10100000", --  941 - 0x3ad  :  160 - 0xa0
    "10100000", --  942 - 0x3ae  :  160 - 0xa0
    "10100000", --  943 - 0x3af  :  160 - 0xa0
    "10100000", --  944 - 0x3b0  :  160 - 0xa0
    "10100000", --  945 - 0x3b1  :  160 - 0xa0
    "10100000", --  946 - 0x3b2  :  160 - 0xa0
    "10100000", --  947 - 0x3b3  :  160 - 0xa0
    "10100000", --  948 - 0x3b4  :  160 - 0xa0
    "10100000", --  949 - 0x3b5  :  160 - 0xa0
    "10100000", --  950 - 0x3b6  :  160 - 0xa0
    "10100000", --  951 - 0x3b7  :  160 - 0xa0
    "10100000", --  952 - 0x3b8  :  160 - 0xa0
    "10100000", --  953 - 0x3b9  :  160 - 0xa0
    "10100000", --  954 - 0x3ba  :  160 - 0xa0
    "10100000", --  955 - 0x3bb  :  160 - 0xa0
    "10100000", --  956 - 0x3bc  :  160 - 0xa0
    "10100000", --  957 - 0x3bd  :  160 - 0xa0
    "10100000", --  958 - 0x3be  :  160 - 0xa0
    "10100000", --  959 - 0x3bf  :  160 - 0xa0
        ---- Attribute Table 0----
    "00000000", --  960 - 0x3c0  :    0 - 0x0
    "00000000", --  961 - 0x3c1  :    0 - 0x0
    "00000000", --  962 - 0x3c2  :    0 - 0x0
    "00000000", --  963 - 0x3c3  :    0 - 0x0
    "00000000", --  964 - 0x3c4  :    0 - 0x0
    "00000000", --  965 - 0x3c5  :    0 - 0x0
    "00000000", --  966 - 0x3c6  :    0 - 0x0
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "10000000", --  968 - 0x3c8  :  128 - 0x80
    "10100000", --  969 - 0x3c9  :  160 - 0xa0
    "10100000", --  970 - 0x3ca  :  160 - 0xa0
    "10100000", --  971 - 0x3cb  :  160 - 0xa0
    "10100000", --  972 - 0x3cc  :  160 - 0xa0
    "10100000", --  973 - 0x3cd  :  160 - 0xa0
    "10100000", --  974 - 0x3ce  :  160 - 0xa0
    "00100000", --  975 - 0x3cf  :   32 - 0x20
    "10001000", --  976 - 0x3d0  :  136 - 0x88
    "10101010", --  977 - 0x3d1  :  170 - 0xaa
    "10101010", --  978 - 0x3d2  :  170 - 0xaa
    "10101010", --  979 - 0x3d3  :  170 - 0xaa
    "10101010", --  980 - 0x3d4  :  170 - 0xaa
    "10101010", --  981 - 0x3d5  :  170 - 0xaa
    "10101010", --  982 - 0x3d6  :  170 - 0xaa
    "00100010", --  983 - 0x3d7  :   34 - 0x22
    "10001000", --  984 - 0x3d8  :  136 - 0x88
    "10101010", --  985 - 0x3d9  :  170 - 0xaa
    "10101010", --  986 - 0x3da  :  170 - 0xaa
    "10101010", --  987 - 0x3db  :  170 - 0xaa
    "10101010", --  988 - 0x3dc  :  170 - 0xaa
    "10101010", --  989 - 0x3dd  :  170 - 0xaa
    "10101010", --  990 - 0x3de  :  170 - 0xaa
    "00100010", --  991 - 0x3df  :   34 - 0x22
    "10001000", --  992 - 0x3e0  :  136 - 0x88
    "10101010", --  993 - 0x3e1  :  170 - 0xaa
    "10101010", --  994 - 0x3e2  :  170 - 0xaa
    "10101010", --  995 - 0x3e3  :  170 - 0xaa
    "10101010", --  996 - 0x3e4  :  170 - 0xaa
    "10101010", --  997 - 0x3e5  :  170 - 0xaa
    "10101010", --  998 - 0x3e6  :  170 - 0xaa
    "00100010", --  999 - 0x3e7  :   34 - 0x22
    "10001000", -- 1000 - 0x3e8  :  136 - 0x88
    "10101010", -- 1001 - 0x3e9  :  170 - 0xaa
    "10101010", -- 1002 - 0x3ea  :  170 - 0xaa
    "10101010", -- 1003 - 0x3eb  :  170 - 0xaa
    "10101010", -- 1004 - 0x3ec  :  170 - 0xaa
    "10101010", -- 1005 - 0x3ed  :  170 - 0xaa
    "10101010", -- 1006 - 0x3ee  :  170 - 0xaa
    "00100010", -- 1007 - 0x3ef  :   34 - 0x22
    "10001000", -- 1008 - 0x3f0  :  136 - 0x88
    "10101010", -- 1009 - 0x3f1  :  170 - 0xaa
    "10101010", -- 1010 - 0x3f2  :  170 - 0xaa
    "10101010", -- 1011 - 0x3f3  :  170 - 0xaa
    "10101010", -- 1012 - 0x3f4  :  170 - 0xaa
    "10101010", -- 1013 - 0x3f5  :  170 - 0xaa
    "10101010", -- 1014 - 0x3f6  :  170 - 0xaa
    "00100010", -- 1015 - 0x3f7  :   34 - 0x22
    "00000000", -- 1016 - 0x3f8  :    0 - 0x0
    "00000000", -- 1017 - 0x3f9  :    0 - 0x0
    "00000000", -- 1018 - 0x3fa  :    0 - 0x0
    "00000000", -- 1019 - 0x3fb  :    0 - 0x0
    "00000000", -- 1020 - 0x3fc  :    0 - 0x0
    "00000000", -- 1021 - 0x3fd  :    0 - 0x0
    "00000000", -- 1022 - 0x3fe  :    0 - 0x0
    "00000000"  -- 1023 - 0x3ff  :    0 - 0x0
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
