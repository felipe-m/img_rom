//-   Sprites Pattern table BOTH COLOR PLANES
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
//- Autcmatically generated verilog ROM from a NES memory file----


//-  Original memory dump file name: nova_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_PTABLE_NOVA_SPR
  (
     //input     clk,   // clock
     input      [12-1:0] addr,  //4096 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Sprite pattern Table both color planes
      12'h0: dout  = 8'b00000000; //    0 :   0 - 0x0 -- Sprite 0x0
      12'h1: dout  = 8'b00001111; //    1 :  15 - 0xf
      12'h2: dout  = 8'b00000100; //    2 :   4 - 0x4
      12'h3: dout  = 8'b00000011; //    3 :   3 - 0x3
      12'h4: dout  = 8'b00000011; //    4 :   3 - 0x3
      12'h5: dout  = 8'b00000011; //    5 :   3 - 0x3
      12'h6: dout  = 8'b00000100; //    6 :   4 - 0x4
      12'h7: dout  = 8'b00111010; //    7 :  58 - 0x3a
      12'h8: dout  = 8'b00000000; //    8 :   0 - 0x0 -- plane 1
      12'h9: dout  = 8'b00000000; //    9 :   0 - 0x0
      12'hA: dout  = 8'b00000011; //   10 :   3 - 0x3
      12'hB: dout  = 8'b00000001; //   11 :   1 - 0x1
      12'hC: dout  = 8'b00000001; //   12 :   1 - 0x1
      12'hD: dout  = 8'b00000000; //   13 :   0 - 0x0
      12'hE: dout  = 8'b00000011; //   14 :   3 - 0x3
      12'hF: dout  = 8'b00000001; //   15 :   1 - 0x1
      12'h10: dout  = 8'b00000000; //   16 :   0 - 0x0 -- Sprite 0x1
      12'h11: dout  = 8'b00111000; //   17 :  56 - 0x38
      12'h12: dout  = 8'b11000110; //   18 : 198 - 0xc6
      12'h13: dout  = 8'b11001011; //   19 : 203 - 0xcb
      12'h14: dout  = 8'b11011100; //   20 : 220 - 0xdc
      12'h15: dout  = 8'b00111010; //   21 :  58 - 0x3a
      12'h16: dout  = 8'b10011010; //   22 : 154 - 0x9a
      12'h17: dout  = 8'b10000001; //   23 : 129 - 0x81
      12'h18: dout  = 8'b00000000; //   24 :   0 - 0x0 -- plane 1
      12'h19: dout  = 8'b00000000; //   25 :   0 - 0x0
      12'h1A: dout  = 8'b00111000; //   26 :  56 - 0x38
      12'h1B: dout  = 8'b10110100; //   27 : 180 - 0xb4
      12'h1C: dout  = 8'b10101000; //   28 : 168 - 0xa8
      12'h1D: dout  = 8'b11010100; //   29 : 212 - 0xd4
      12'h1E: dout  = 8'b01110100; //   30 : 116 - 0x74
      12'h1F: dout  = 8'b01111110; //   31 : 126 - 0x7e
      12'h20: dout  = 8'b01000101; //   32 :  69 - 0x45 -- Sprite 0x2
      12'h21: dout  = 8'b10000111; //   33 : 135 - 0x87
      12'h22: dout  = 8'b10000011; //   34 : 131 - 0x83
      12'h23: dout  = 8'b10000001; //   35 : 129 - 0x81
      12'h24: dout  = 8'b10000001; //   36 : 129 - 0x81
      12'h25: dout  = 8'b10000001; //   37 : 129 - 0x81
      12'h26: dout  = 8'b01000001; //   38 :  65 - 0x41
      12'h27: dout  = 8'b00100001; //   39 :  33 - 0x21
      12'h28: dout  = 8'b00111000; //   40 :  56 - 0x38 -- plane 1
      12'h29: dout  = 8'b01111000; //   41 : 120 - 0x78
      12'h2A: dout  = 8'b01111100; //   42 : 124 - 0x7c
      12'h2B: dout  = 8'b01111110; //   43 : 126 - 0x7e
      12'h2C: dout  = 8'b01111110; //   44 : 126 - 0x7e
      12'h2D: dout  = 8'b01111110; //   45 : 126 - 0x7e
      12'h2E: dout  = 8'b00111110; //   46 :  62 - 0x3e
      12'h2F: dout  = 8'b00011110; //   47 :  30 - 0x1e
      12'h30: dout  = 8'b01111111; //   48 : 127 - 0x7f -- Sprite 0x3
      12'h31: dout  = 8'b01111110; //   49 : 126 - 0x7e
      12'h32: dout  = 8'b11111100; //   50 : 252 - 0xfc
      12'h33: dout  = 8'b00111000; //   51 :  56 - 0x38
      12'h34: dout  = 8'b00011000; //   52 :  24 - 0x18
      12'h35: dout  = 8'b10001100; //   53 : 140 - 0x8c
      12'h36: dout  = 8'b11000100; //   54 : 196 - 0xc4
      12'h37: dout  = 8'b11111100; //   55 : 252 - 0xfc
      12'h38: dout  = 8'b11110110; //   56 : 246 - 0xf6 -- plane 1
      12'h39: dout  = 8'b11110000; //   57 : 240 - 0xf0
      12'h3A: dout  = 8'b00111000; //   58 :  56 - 0x38
      12'h3B: dout  = 8'b11010000; //   59 : 208 - 0xd0
      12'h3C: dout  = 8'b11100000; //   60 : 224 - 0xe0
      12'h3D: dout  = 8'b01110000; //   61 : 112 - 0x70
      12'h3E: dout  = 8'b10111000; //   62 : 184 - 0xb8
      12'h3F: dout  = 8'b01000000; //   63 :  64 - 0x40
      12'h40: dout  = 8'b00100011; //   64 :  35 - 0x23 -- Sprite 0x4
      12'h41: dout  = 8'b00100011; //   65 :  35 - 0x23
      12'h42: dout  = 8'b00100001; //   66 :  33 - 0x21
      12'h43: dout  = 8'b00100000; //   67 :  32 - 0x20
      12'h44: dout  = 8'b00010011; //   68 :  19 - 0x13
      12'h45: dout  = 8'b00001100; //   69 :  12 - 0xc
      12'h46: dout  = 8'b00000000; //   70 :   0 - 0x0
      12'h47: dout  = 8'b00000000; //   71 :   0 - 0x0
      12'h48: dout  = 8'b00011100; //   72 :  28 - 0x1c -- plane 1
      12'h49: dout  = 8'b00011100; //   73 :  28 - 0x1c
      12'h4A: dout  = 8'b00011110; //   74 :  30 - 0x1e
      12'h4B: dout  = 8'b00011111; //   75 :  31 - 0x1f
      12'h4C: dout  = 8'b00001100; //   76 :  12 - 0xc
      12'h4D: dout  = 8'b00000000; //   77 :   0 - 0x0
      12'h4E: dout  = 8'b00000000; //   78 :   0 - 0x0
      12'h4F: dout  = 8'b00000000; //   79 :   0 - 0x0
      12'h50: dout  = 8'b11111100; //   80 : 252 - 0xfc -- Sprite 0x5
      12'h51: dout  = 8'b11111100; //   81 : 252 - 0xfc
      12'h52: dout  = 8'b11111100; //   82 : 252 - 0xfc
      12'h53: dout  = 8'b11111100; //   83 : 252 - 0xfc
      12'h54: dout  = 8'b10010000; //   84 : 144 - 0x90
      12'h55: dout  = 8'b10010000; //   85 : 144 - 0x90
      12'h56: dout  = 8'b10001000; //   86 : 136 - 0x88
      12'h57: dout  = 8'b11111000; //   87 : 248 - 0xf8
      12'h58: dout  = 8'b10101000; //   88 : 168 - 0xa8 -- plane 1
      12'h59: dout  = 8'b01010000; //   89 :  80 - 0x50
      12'h5A: dout  = 8'b10101000; //   90 : 168 - 0xa8
      12'h5B: dout  = 8'b00000000; //   91 :   0 - 0x0
      12'h5C: dout  = 8'b01100000; //   92 :  96 - 0x60
      12'h5D: dout  = 8'b01100000; //   93 :  96 - 0x60
      12'h5E: dout  = 8'b01110000; //   94 : 112 - 0x70
      12'h5F: dout  = 8'b00000000; //   95 :   0 - 0x0
      12'h60: dout  = 8'b00100011; //   96 :  35 - 0x23 -- Sprite 0x6
      12'h61: dout  = 8'b00100011; //   97 :  35 - 0x23
      12'h62: dout  = 8'b00100001; //   98 :  33 - 0x21
      12'h63: dout  = 8'b00100000; //   99 :  32 - 0x20
      12'h64: dout  = 8'b00010011; //  100 :  19 - 0x13
      12'h65: dout  = 8'b00001101; //  101 :  13 - 0xd
      12'h66: dout  = 8'b00000010; //  102 :   2 - 0x2
      12'h67: dout  = 8'b00000001; //  103 :   1 - 0x1
      12'h68: dout  = 8'b00011100; //  104 :  28 - 0x1c -- plane 1
      12'h69: dout  = 8'b00011100; //  105 :  28 - 0x1c
      12'h6A: dout  = 8'b00011110; //  106 :  30 - 0x1e
      12'h6B: dout  = 8'b00011111; //  107 :  31 - 0x1f
      12'h6C: dout  = 8'b00001100; //  108 :  12 - 0xc
      12'h6D: dout  = 8'b00000000; //  109 :   0 - 0x0
      12'h6E: dout  = 8'b00000001; //  110 :   1 - 0x1
      12'h6F: dout  = 8'b00000000; //  111 :   0 - 0x0
      12'h70: dout  = 8'b11111100; //  112 : 252 - 0xfc -- Sprite 0x7
      12'h71: dout  = 8'b11111100; //  113 : 252 - 0xfc
      12'h72: dout  = 8'b11111100; //  114 : 252 - 0xfc
      12'h73: dout  = 8'b11111100; //  115 : 252 - 0xfc
      12'h74: dout  = 8'b10100100; //  116 : 164 - 0xa4
      12'h75: dout  = 8'b00100100; //  117 :  36 - 0x24
      12'h76: dout  = 8'b01010010; //  118 :  82 - 0x52
      12'h77: dout  = 8'b11101110; //  119 : 238 - 0xee
      12'h78: dout  = 8'b10101000; //  120 : 168 - 0xa8 -- plane 1
      12'h79: dout  = 8'b01010000; //  121 :  80 - 0x50
      12'h7A: dout  = 8'b10101000; //  122 : 168 - 0xa8
      12'h7B: dout  = 8'b00000000; //  123 :   0 - 0x0
      12'h7C: dout  = 8'b01011000; //  124 :  88 - 0x58
      12'h7D: dout  = 8'b11011000; //  125 : 216 - 0xd8
      12'h7E: dout  = 8'b10001100; //  126 : 140 - 0x8c
      12'h7F: dout  = 8'b00000000; //  127 :   0 - 0x0
      12'h80: dout  = 8'b00100011; //  128 :  35 - 0x23 -- Sprite 0x8
      12'h81: dout  = 8'b00100011; //  129 :  35 - 0x23
      12'h82: dout  = 8'b00100001; //  130 :  33 - 0x21
      12'h83: dout  = 8'b00100000; //  131 :  32 - 0x20
      12'h84: dout  = 8'b00010011; //  132 :  19 - 0x13
      12'h85: dout  = 8'b00001101; //  133 :  13 - 0xd
      12'h86: dout  = 8'b00000001; //  134 :   1 - 0x1
      12'h87: dout  = 8'b00000001; //  135 :   1 - 0x1
      12'h88: dout  = 8'b00011100; //  136 :  28 - 0x1c -- plane 1
      12'h89: dout  = 8'b00011100; //  137 :  28 - 0x1c
      12'h8A: dout  = 8'b00011110; //  138 :  30 - 0x1e
      12'h8B: dout  = 8'b00011111; //  139 :  31 - 0x1f
      12'h8C: dout  = 8'b00001100; //  140 :  12 - 0xc
      12'h8D: dout  = 8'b00000000; //  141 :   0 - 0x0
      12'h8E: dout  = 8'b00000000; //  142 :   0 - 0x0
      12'h8F: dout  = 8'b00000000; //  143 :   0 - 0x0
      12'h90: dout  = 8'b11111110; //  144 : 254 - 0xfe -- Sprite 0x9
      12'h91: dout  = 8'b11111110; //  145 : 254 - 0xfe
      12'h92: dout  = 8'b11111110; //  146 : 254 - 0xfe
      12'h93: dout  = 8'b11111111; //  147 : 255 - 0xff
      12'h94: dout  = 8'b10010001; //  148 : 145 - 0x91
      12'h95: dout  = 8'b00101111; //  149 :  47 - 0x2f
      12'h96: dout  = 8'b01000000; //  150 :  64 - 0x40
      12'h97: dout  = 8'b11100000; //  151 : 224 - 0xe0
      12'h98: dout  = 8'b10101000; //  152 : 168 - 0xa8 -- plane 1
      12'h99: dout  = 8'b01010100; //  153 :  84 - 0x54
      12'h9A: dout  = 8'b10101000; //  154 : 168 - 0xa8
      12'h9B: dout  = 8'b00000000; //  155 :   0 - 0x0
      12'h9C: dout  = 8'b01101110; //  156 : 110 - 0x6e
      12'h9D: dout  = 8'b11000000; //  157 : 192 - 0xc0
      12'h9E: dout  = 8'b10000000; //  158 : 128 - 0x80
      12'h9F: dout  = 8'b00000000; //  159 :   0 - 0x0
      12'hA0: dout  = 8'b00100011; //  160 :  35 - 0x23 -- Sprite 0xa
      12'hA1: dout  = 8'b00100011; //  161 :  35 - 0x23
      12'hA2: dout  = 8'b00100001; //  162 :  33 - 0x21
      12'hA3: dout  = 8'b00100000; //  163 :  32 - 0x20
      12'hA4: dout  = 8'b00010011; //  164 :  19 - 0x13
      12'hA5: dout  = 8'b00001110; //  165 :  14 - 0xe
      12'hA6: dout  = 8'b00000001; //  166 :   1 - 0x1
      12'hA7: dout  = 8'b00000000; //  167 :   0 - 0x0
      12'hA8: dout  = 8'b00011100; //  168 :  28 - 0x1c -- plane 1
      12'hA9: dout  = 8'b00011100; //  169 :  28 - 0x1c
      12'hAA: dout  = 8'b00011110; //  170 :  30 - 0x1e
      12'hAB: dout  = 8'b00011111; //  171 :  31 - 0x1f
      12'hAC: dout  = 8'b00001100; //  172 :  12 - 0xc
      12'hAD: dout  = 8'b00000001; //  173 :   1 - 0x1
      12'hAE: dout  = 8'b00000000; //  174 :   0 - 0x0
      12'hAF: dout  = 8'b00000000; //  175 :   0 - 0x0
      12'hB0: dout  = 8'b11111110; //  176 : 254 - 0xfe -- Sprite 0xb
      12'hB1: dout  = 8'b11111110; //  177 : 254 - 0xfe
      12'hB2: dout  = 8'b11111110; //  178 : 254 - 0xfe
      12'hB3: dout  = 8'b11111100; //  179 : 252 - 0xfc
      12'hB4: dout  = 8'b00100100; //  180 :  36 - 0x24
      12'hB5: dout  = 8'b00100010; //  181 :  34 - 0x22
      12'hB6: dout  = 8'b11010010; //  182 : 210 - 0xd2
      12'hB7: dout  = 8'b00001111; //  183 :  15 - 0xf
      12'hB8: dout  = 8'b10101000; //  184 : 168 - 0xa8 -- plane 1
      12'hB9: dout  = 8'b01010100; //  185 :  84 - 0x54
      12'hBA: dout  = 8'b10101000; //  186 : 168 - 0xa8
      12'hBB: dout  = 8'b00000000; //  187 :   0 - 0x0
      12'hBC: dout  = 8'b11011000; //  188 : 216 - 0xd8
      12'hBD: dout  = 8'b11011100; //  189 : 220 - 0xdc
      12'hBE: dout  = 8'b00001100; //  190 :  12 - 0xc
      12'hBF: dout  = 8'b00000000; //  191 :   0 - 0x0
      12'hC0: dout  = 8'b01111111; //  192 : 127 - 0x7f -- Sprite 0xc
      12'hC1: dout  = 8'b01111110; //  193 : 126 - 0x7e
      12'hC2: dout  = 8'b11111100; //  194 : 252 - 0xfc
      12'hC3: dout  = 8'b00000010; //  195 :   2 - 0x2
      12'hC4: dout  = 8'b00000100; //  196 :   4 - 0x4
      12'hC5: dout  = 8'b11111100; //  197 : 252 - 0xfc
      12'hC6: dout  = 8'b11111100; //  198 : 252 - 0xfc
      12'hC7: dout  = 8'b11111110; //  199 : 254 - 0xfe
      12'hC8: dout  = 8'b11110110; //  200 : 246 - 0xf6 -- plane 1
      12'hC9: dout  = 8'b11110000; //  201 : 240 - 0xf0
      12'hCA: dout  = 8'b00000000; //  202 :   0 - 0x0
      12'hCB: dout  = 8'b11111100; //  203 : 252 - 0xfc
      12'hCC: dout  = 8'b11111000; //  204 : 248 - 0xf8
      12'hCD: dout  = 8'b00000000; //  205 :   0 - 0x0
      12'hCE: dout  = 8'b10101000; //  206 : 168 - 0xa8
      12'hCF: dout  = 8'b01010100; //  207 :  84 - 0x54
      12'hD0: dout  = 8'b01000101; //  208 :  69 - 0x45 -- Sprite 0xd
      12'hD1: dout  = 8'b10000111; //  209 : 135 - 0x87
      12'hD2: dout  = 8'b10000011; //  210 : 131 - 0x83
      12'hD3: dout  = 8'b10000010; //  211 : 130 - 0x82
      12'hD4: dout  = 8'b10000010; //  212 : 130 - 0x82
      12'hD5: dout  = 8'b10000100; //  213 : 132 - 0x84
      12'hD6: dout  = 8'b01000100; //  214 :  68 - 0x44
      12'hD7: dout  = 8'b00100100; //  215 :  36 - 0x24
      12'hD8: dout  = 8'b00111000; //  216 :  56 - 0x38 -- plane 1
      12'hD9: dout  = 8'b01111000; //  217 : 120 - 0x78
      12'hDA: dout  = 8'b01111100; //  218 : 124 - 0x7c
      12'hDB: dout  = 8'b01111101; //  219 : 125 - 0x7d
      12'hDC: dout  = 8'b01111101; //  220 : 125 - 0x7d
      12'hDD: dout  = 8'b01111011; //  221 : 123 - 0x7b
      12'hDE: dout  = 8'b00111011; //  222 :  59 - 0x3b
      12'hDF: dout  = 8'b00011011; //  223 :  27 - 0x1b
      12'hE0: dout  = 8'b01111111; //  224 : 127 - 0x7f -- Sprite 0xe
      12'hE1: dout  = 8'b01111110; //  225 : 126 - 0x7e
      12'hE2: dout  = 8'b11111100; //  226 : 252 - 0xfc
      12'hE3: dout  = 8'b11111000; //  227 : 248 - 0xf8
      12'hE4: dout  = 8'b01111000; //  228 : 120 - 0x78
      12'hE5: dout  = 8'b01111100; //  229 : 124 - 0x7c
      12'hE6: dout  = 8'b11111100; //  230 : 252 - 0xfc
      12'hE7: dout  = 8'b11111110; //  231 : 254 - 0xfe
      12'hE8: dout  = 8'b11110110; //  232 : 246 - 0xf6 -- plane 1
      12'hE9: dout  = 8'b11110000; //  233 : 240 - 0xf0
      12'hEA: dout  = 8'b01111000; //  234 : 120 - 0x78
      12'hEB: dout  = 8'b01110000; //  235 : 112 - 0x70
      12'hEC: dout  = 8'b10100000; //  236 : 160 - 0xa0
      12'hED: dout  = 8'b10010000; //  237 : 144 - 0x90
      12'hEE: dout  = 8'b00101000; //  238 :  40 - 0x28
      12'hEF: dout  = 8'b01010100; //  239 :  84 - 0x54
      12'hF0: dout  = 8'b00000000; //  240 :   0 - 0x0 -- Sprite 0xf
      12'hF1: dout  = 8'b00001111; //  241 :  15 - 0xf
      12'hF2: dout  = 8'b00000100; //  242 :   4 - 0x4
      12'hF3: dout  = 8'b00000011; //  243 :   3 - 0x3
      12'hF4: dout  = 8'b00000011; //  244 :   3 - 0x3
      12'hF5: dout  = 8'b00000011; //  245 :   3 - 0x3
      12'hF6: dout  = 8'b00000100; //  246 :   4 - 0x4
      12'hF7: dout  = 8'b00000010; //  247 :   2 - 0x2
      12'hF8: dout  = 8'b00000000; //  248 :   0 - 0x0 -- plane 1
      12'hF9: dout  = 8'b00000000; //  249 :   0 - 0x0
      12'hFA: dout  = 8'b00000011; //  250 :   3 - 0x3
      12'hFB: dout  = 8'b00000001; //  251 :   1 - 0x1
      12'hFC: dout  = 8'b00000001; //  252 :   1 - 0x1
      12'hFD: dout  = 8'b00000000; //  253 :   0 - 0x0
      12'hFE: dout  = 8'b00000011; //  254 :   3 - 0x3
      12'hFF: dout  = 8'b00000001; //  255 :   1 - 0x1
      12'h100: dout  = 8'b00000111; //  256 :   7 - 0x7 -- Sprite 0x10
      12'h101: dout  = 8'b00001100; //  257 :  12 - 0xc
      12'h102: dout  = 8'b00010000; //  258 :  16 - 0x10
      12'h103: dout  = 8'b00010000; //  259 :  16 - 0x10
      12'h104: dout  = 8'b00010000; //  260 :  16 - 0x10
      12'h105: dout  = 8'b00100000; //  261 :  32 - 0x20
      12'h106: dout  = 8'b00100000; //  262 :  32 - 0x20
      12'h107: dout  = 8'b00100001; //  263 :  33 - 0x21
      12'h108: dout  = 8'b00000000; //  264 :   0 - 0x0 -- plane 1
      12'h109: dout  = 8'b00000011; //  265 :   3 - 0x3
      12'h10A: dout  = 8'b00001111; //  266 :  15 - 0xf
      12'h10B: dout  = 8'b00001111; //  267 :  15 - 0xf
      12'h10C: dout  = 8'b00001111; //  268 :  15 - 0xf
      12'h10D: dout  = 8'b00011111; //  269 :  31 - 0x1f
      12'h10E: dout  = 8'b00011111; //  270 :  31 - 0x1f
      12'h10F: dout  = 8'b00011110; //  271 :  30 - 0x1e
      12'h110: dout  = 8'b11111111; //  272 : 255 - 0xff -- Sprite 0x11
      12'h111: dout  = 8'b01111110; //  273 : 126 - 0x7e
      12'h112: dout  = 8'b01111100; //  274 : 124 - 0x7c
      12'h113: dout  = 8'b01111000; //  275 : 120 - 0x78
      12'h114: dout  = 8'b01011000; //  276 :  88 - 0x58
      12'h115: dout  = 8'b10001100; //  277 : 140 - 0x8c
      12'h116: dout  = 8'b11000100; //  278 : 196 - 0xc4
      12'h117: dout  = 8'b11111100; //  279 : 252 - 0xfc
      12'h118: dout  = 8'b00110110; //  280 :  54 - 0x36 -- plane 1
      12'h119: dout  = 8'b10110000; //  281 : 176 - 0xb0
      12'h11A: dout  = 8'b10111000; //  282 : 184 - 0xb8
      12'h11B: dout  = 8'b10010000; //  283 : 144 - 0x90
      12'h11C: dout  = 8'b10100000; //  284 : 160 - 0xa0
      12'h11D: dout  = 8'b01110000; //  285 : 112 - 0x70
      12'h11E: dout  = 8'b00111000; //  286 :  56 - 0x38
      12'h11F: dout  = 8'b01000000; //  287 :  64 - 0x40
      12'h120: dout  = 8'b00100011; //  288 :  35 - 0x23 -- Sprite 0x12
      12'h121: dout  = 8'b00100011; //  289 :  35 - 0x23
      12'h122: dout  = 8'b00100001; //  290 :  33 - 0x21
      12'h123: dout  = 8'b00100000; //  291 :  32 - 0x20
      12'h124: dout  = 8'b00010011; //  292 :  19 - 0x13
      12'h125: dout  = 8'b00001100; //  293 :  12 - 0xc
      12'h126: dout  = 8'b00000000; //  294 :   0 - 0x0
      12'h127: dout  = 8'b00000000; //  295 :   0 - 0x0
      12'h128: dout  = 8'b00011100; //  296 :  28 - 0x1c -- plane 1
      12'h129: dout  = 8'b00011100; //  297 :  28 - 0x1c
      12'h12A: dout  = 8'b00011110; //  298 :  30 - 0x1e
      12'h12B: dout  = 8'b00011111; //  299 :  31 - 0x1f
      12'h12C: dout  = 8'b00001100; //  300 :  12 - 0xc
      12'h12D: dout  = 8'b00000000; //  301 :   0 - 0x0
      12'h12E: dout  = 8'b00000000; //  302 :   0 - 0x0
      12'h12F: dout  = 8'b00000000; //  303 :   0 - 0x0
      12'h130: dout  = 8'b00000001; //  304 :   1 - 0x1 -- Sprite 0x13
      12'h131: dout  = 8'b00000001; //  305 :   1 - 0x1
      12'h132: dout  = 8'b00000011; //  306 :   3 - 0x3
      12'h133: dout  = 8'b00000100; //  307 :   4 - 0x4
      12'h134: dout  = 8'b00001000; //  308 :   8 - 0x8
      12'h135: dout  = 8'b00010000; //  309 :  16 - 0x10
      12'h136: dout  = 8'b00010000; //  310 :  16 - 0x10
      12'h137: dout  = 8'b00100000; //  311 :  32 - 0x20
      12'h138: dout  = 8'b00000000; //  312 :   0 - 0x0 -- plane 1
      12'h139: dout  = 8'b00000000; //  313 :   0 - 0x0
      12'h13A: dout  = 8'b00000000; //  314 :   0 - 0x0
      12'h13B: dout  = 8'b00000011; //  315 :   3 - 0x3
      12'h13C: dout  = 8'b00000111; //  316 :   7 - 0x7
      12'h13D: dout  = 8'b00001111; //  317 :  15 - 0xf
      12'h13E: dout  = 8'b00001111; //  318 :  15 - 0xf
      12'h13F: dout  = 8'b00011111; //  319 :  31 - 0x1f
      12'h140: dout  = 8'b01111111; //  320 : 127 - 0x7f -- Sprite 0x14
      12'h141: dout  = 8'b11111110; //  321 : 254 - 0xfe
      12'h142: dout  = 8'b00000110; //  322 :   6 - 0x6
      12'h143: dout  = 8'b00000001; //  323 :   1 - 0x1
      12'h144: dout  = 8'b00000001; //  324 :   1 - 0x1
      12'h145: dout  = 8'b00000001; //  325 :   1 - 0x1
      12'h146: dout  = 8'b00000111; //  326 :   7 - 0x7
      12'h147: dout  = 8'b11111110; //  327 : 254 - 0xfe
      12'h148: dout  = 8'b11110110; //  328 : 246 - 0xf6 -- plane 1
      12'h149: dout  = 8'b00000000; //  329 :   0 - 0x0
      12'h14A: dout  = 8'b11111000; //  330 : 248 - 0xf8
      12'h14B: dout  = 8'b11111110; //  331 : 254 - 0xfe
      12'h14C: dout  = 8'b11111110; //  332 : 254 - 0xfe
      12'h14D: dout  = 8'b11111110; //  333 : 254 - 0xfe
      12'h14E: dout  = 8'b11111000; //  334 : 248 - 0xf8
      12'h14F: dout  = 8'b00000000; //  335 :   0 - 0x0
      12'h150: dout  = 8'b00000101; //  336 :   5 - 0x5 -- Sprite 0x15
      12'h151: dout  = 8'b00000101; //  337 :   5 - 0x5
      12'h152: dout  = 8'b00000111; //  338 :   7 - 0x7
      12'h153: dout  = 8'b00000100; //  339 :   4 - 0x4
      12'h154: dout  = 8'b00000100; //  340 :   4 - 0x4
      12'h155: dout  = 8'b00001111; //  341 :  15 - 0xf
      12'h156: dout  = 8'b00110000; //  342 :  48 - 0x30
      12'h157: dout  = 8'b01000000; //  343 :  64 - 0x40
      12'h158: dout  = 8'b00000011; //  344 :   3 - 0x3 -- plane 1
      12'h159: dout  = 8'b00000011; //  345 :   3 - 0x3
      12'h15A: dout  = 8'b00000000; //  346 :   0 - 0x0
      12'h15B: dout  = 8'b00000011; //  347 :   3 - 0x3
      12'h15C: dout  = 8'b00000011; //  348 :   3 - 0x3
      12'h15D: dout  = 8'b00000000; //  349 :   0 - 0x0
      12'h15E: dout  = 8'b00001111; //  350 :  15 - 0xf
      12'h15F: dout  = 8'b00111111; //  351 :  63 - 0x3f
      12'h160: dout  = 8'b11111100; //  352 : 252 - 0xfc -- Sprite 0x16
      12'h161: dout  = 8'b11111000; //  353 : 248 - 0xf8
      12'h162: dout  = 8'b11110000; //  354 : 240 - 0xf0
      12'h163: dout  = 8'b11100000; //  355 : 224 - 0xe0
      12'h164: dout  = 8'b01100000; //  356 :  96 - 0x60
      12'h165: dout  = 8'b11110000; //  357 : 240 - 0xf0
      12'h166: dout  = 8'b00011100; //  358 :  28 - 0x1c
      12'h167: dout  = 8'b00000010; //  359 :   2 - 0x2
      12'h168: dout  = 8'b11011000; //  360 : 216 - 0xd8 -- plane 1
      12'h169: dout  = 8'b11000000; //  361 : 192 - 0xc0
      12'h16A: dout  = 8'b11100000; //  362 : 224 - 0xe0
      12'h16B: dout  = 8'b01000000; //  363 :  64 - 0x40
      12'h16C: dout  = 8'b10000000; //  364 : 128 - 0x80
      12'h16D: dout  = 8'b00000000; //  365 :   0 - 0x0
      12'h16E: dout  = 8'b11100000; //  366 : 224 - 0xe0
      12'h16F: dout  = 8'b11111100; //  367 : 252 - 0xfc
      12'h170: dout  = 8'b10000000; //  368 : 128 - 0x80 -- Sprite 0x17
      12'h171: dout  = 8'b10000000; //  369 : 128 - 0x80
      12'h172: dout  = 8'b10000000; //  370 : 128 - 0x80
      12'h173: dout  = 8'b10000011; //  371 : 131 - 0x83
      12'h174: dout  = 8'b01001111; //  372 :  79 - 0x4f
      12'h175: dout  = 8'b00110010; //  373 :  50 - 0x32
      12'h176: dout  = 8'b00000010; //  374 :   2 - 0x2
      12'h177: dout  = 8'b00000011; //  375 :   3 - 0x3
      12'h178: dout  = 8'b01111111; //  376 : 127 - 0x7f -- plane 1
      12'h179: dout  = 8'b01111111; //  377 : 127 - 0x7f
      12'h17A: dout  = 8'b01111111; //  378 : 127 - 0x7f
      12'h17B: dout  = 8'b01111100; //  379 : 124 - 0x7c
      12'h17C: dout  = 8'b00110000; //  380 :  48 - 0x30
      12'h17D: dout  = 8'b00000001; //  381 :   1 - 0x1
      12'h17E: dout  = 8'b00000001; //  382 :   1 - 0x1
      12'h17F: dout  = 8'b00000000; //  383 :   0 - 0x0
      12'h180: dout  = 8'b00000010; //  384 :   2 - 0x2 -- Sprite 0x18
      12'h181: dout  = 8'b00000001; //  385 :   1 - 0x1
      12'h182: dout  = 8'b00000010; //  386 :   2 - 0x2
      12'h183: dout  = 8'b11111100; //  387 : 252 - 0xfc
      12'h184: dout  = 8'b11000000; //  388 : 192 - 0xc0
      12'h185: dout  = 8'b01000000; //  389 :  64 - 0x40
      12'h186: dout  = 8'b00100000; //  390 :  32 - 0x20
      12'h187: dout  = 8'b11100000; //  391 : 224 - 0xe0
      12'h188: dout  = 8'b11111100; //  392 : 252 - 0xfc -- plane 1
      12'h189: dout  = 8'b11111110; //  393 : 254 - 0xfe
      12'h18A: dout  = 8'b11111100; //  394 : 252 - 0xfc
      12'h18B: dout  = 8'b00000000; //  395 :   0 - 0x0
      12'h18C: dout  = 8'b00000000; //  396 :   0 - 0x0
      12'h18D: dout  = 8'b10000000; //  397 : 128 - 0x80
      12'h18E: dout  = 8'b11000000; //  398 : 192 - 0xc0
      12'h18F: dout  = 8'b00000000; //  399 :   0 - 0x0
      12'h190: dout  = 8'b00001011; //  400 :  11 - 0xb -- Sprite 0x19
      12'h191: dout  = 8'b00001011; //  401 :  11 - 0xb
      12'h192: dout  = 8'b00001111; //  402 :  15 - 0xf
      12'h193: dout  = 8'b00001001; //  403 :   9 - 0x9
      12'h194: dout  = 8'b00001000; //  404 :   8 - 0x8
      12'h195: dout  = 8'b00001001; //  405 :   9 - 0x9
      12'h196: dout  = 8'b00001111; //  406 :  15 - 0xf
      12'h197: dout  = 8'b00110000; //  407 :  48 - 0x30
      12'h198: dout  = 8'b00000111; //  408 :   7 - 0x7 -- plane 1
      12'h199: dout  = 8'b00000111; //  409 :   7 - 0x7
      12'h19A: dout  = 8'b00000001; //  410 :   1 - 0x1
      12'h19B: dout  = 8'b00000110; //  411 :   6 - 0x6
      12'h19C: dout  = 8'b00000111; //  412 :   7 - 0x7
      12'h19D: dout  = 8'b00000110; //  413 :   6 - 0x6
      12'h19E: dout  = 8'b00000000; //  414 :   0 - 0x0
      12'h19F: dout  = 8'b00001111; //  415 :  15 - 0xf
      12'h1A0: dout  = 8'b11111000; //  416 : 248 - 0xf8 -- Sprite 0x1a
      12'h1A1: dout  = 8'b11110000; //  417 : 240 - 0xf0
      12'h1A2: dout  = 8'b11100000; //  418 : 224 - 0xe0
      12'h1A3: dout  = 8'b11000000; //  419 : 192 - 0xc0
      12'h1A4: dout  = 8'b11000000; //  420 : 192 - 0xc0
      12'h1A5: dout  = 8'b11000000; //  421 : 192 - 0xc0
      12'h1A6: dout  = 8'b11111000; //  422 : 248 - 0xf8
      12'h1A7: dout  = 8'b00011111; //  423 :  31 - 0x1f
      12'h1A8: dout  = 8'b10110000; //  424 : 176 - 0xb0 -- plane 1
      12'h1A9: dout  = 8'b10000000; //  425 : 128 - 0x80
      12'h1AA: dout  = 8'b11000000; //  426 : 192 - 0xc0
      12'h1AB: dout  = 8'b10000000; //  427 : 128 - 0x80
      12'h1AC: dout  = 8'b00000000; //  428 :   0 - 0x0
      12'h1AD: dout  = 8'b00000000; //  429 :   0 - 0x0
      12'h1AE: dout  = 8'b00000000; //  430 :   0 - 0x0
      12'h1AF: dout  = 8'b11100000; //  431 : 224 - 0xe0
      12'h1B0: dout  = 8'b01000000; //  432 :  64 - 0x40 -- Sprite 0x1b
      12'h1B1: dout  = 8'b01000000; //  433 :  64 - 0x40
      12'h1B2: dout  = 8'b10000000; //  434 : 128 - 0x80
      12'h1B3: dout  = 8'b10000000; //  435 : 128 - 0x80
      12'h1B4: dout  = 8'b01000000; //  436 :  64 - 0x40
      12'h1B5: dout  = 8'b00111111; //  437 :  63 - 0x3f
      12'h1B6: dout  = 8'b00000100; //  438 :   4 - 0x4
      12'h1B7: dout  = 8'b00000111; //  439 :   7 - 0x7
      12'h1B8: dout  = 8'b00111111; //  440 :  63 - 0x3f -- plane 1
      12'h1B9: dout  = 8'b00111111; //  441 :  63 - 0x3f
      12'h1BA: dout  = 8'b01111111; //  442 : 127 - 0x7f
      12'h1BB: dout  = 8'b01111111; //  443 : 127 - 0x7f
      12'h1BC: dout  = 8'b00111111; //  444 :  63 - 0x3f
      12'h1BD: dout  = 8'b00000000; //  445 :   0 - 0x0
      12'h1BE: dout  = 8'b00000011; //  446 :   3 - 0x3
      12'h1BF: dout  = 8'b00000000; //  447 :   0 - 0x0
      12'h1C0: dout  = 8'b00000000; //  448 :   0 - 0x0 -- Sprite 0x1c
      12'h1C1: dout  = 8'b00000000; //  449 :   0 - 0x0
      12'h1C2: dout  = 8'b00000000; //  450 :   0 - 0x0
      12'h1C3: dout  = 8'b00000000; //  451 :   0 - 0x0
      12'h1C4: dout  = 8'b00000000; //  452 :   0 - 0x0
      12'h1C5: dout  = 8'b11111111; //  453 : 255 - 0xff
      12'h1C6: dout  = 8'b01000000; //  454 :  64 - 0x40
      12'h1C7: dout  = 8'b11000000; //  455 : 192 - 0xc0
      12'h1C8: dout  = 8'b11111111; //  456 : 255 - 0xff -- plane 1
      12'h1C9: dout  = 8'b11111111; //  457 : 255 - 0xff
      12'h1CA: dout  = 8'b11111111; //  458 : 255 - 0xff
      12'h1CB: dout  = 8'b11111111; //  459 : 255 - 0xff
      12'h1CC: dout  = 8'b11111111; //  460 : 255 - 0xff
      12'h1CD: dout  = 8'b00000000; //  461 :   0 - 0x0
      12'h1CE: dout  = 8'b10000000; //  462 : 128 - 0x80
      12'h1CF: dout  = 8'b00000000; //  463 :   0 - 0x0
      12'h1D0: dout  = 8'b11000000; //  464 : 192 - 0xc0 -- Sprite 0x1d
      12'h1D1: dout  = 8'b00100000; //  465 :  32 - 0x20
      12'h1D2: dout  = 8'b00100000; //  466 :  32 - 0x20
      12'h1D3: dout  = 8'b00100000; //  467 :  32 - 0x20
      12'h1D4: dout  = 8'b01000000; //  468 :  64 - 0x40
      12'h1D5: dout  = 8'b10000000; //  469 : 128 - 0x80
      12'h1D6: dout  = 8'b00000000; //  470 :   0 - 0x0
      12'h1D7: dout  = 8'b00000000; //  471 :   0 - 0x0
      12'h1D8: dout  = 8'b00000000; //  472 :   0 - 0x0 -- plane 1
      12'h1D9: dout  = 8'b11000000; //  473 : 192 - 0xc0
      12'h1DA: dout  = 8'b11000000; //  474 : 192 - 0xc0
      12'h1DB: dout  = 8'b11000000; //  475 : 192 - 0xc0
      12'h1DC: dout  = 8'b10000000; //  476 : 128 - 0x80
      12'h1DD: dout  = 8'b00000000; //  477 :   0 - 0x0
      12'h1DE: dout  = 8'b00000000; //  478 :   0 - 0x0
      12'h1DF: dout  = 8'b00000000; //  479 :   0 - 0x0
      12'h1E0: dout  = 8'b01111111; //  480 : 127 - 0x7f -- Sprite 0x1e
      12'h1E1: dout  = 8'b01100010; //  481 :  98 - 0x62
      12'h1E2: dout  = 8'b11000100; //  482 : 196 - 0xc4
      12'h1E3: dout  = 8'b00011000; //  483 :  24 - 0x18
      12'h1E4: dout  = 8'b00111100; //  484 :  60 - 0x3c
      12'h1E5: dout  = 8'b11111110; //  485 : 254 - 0xfe
      12'h1E6: dout  = 8'b11111110; //  486 : 254 - 0xfe
      12'h1E7: dout  = 8'b11111110; //  487 : 254 - 0xfe
      12'h1E8: dout  = 8'b11100000; //  488 : 224 - 0xe0 -- plane 1
      12'h1E9: dout  = 8'b10011100; //  489 : 156 - 0x9c
      12'h1EA: dout  = 8'b00111000; //  490 :  56 - 0x38
      12'h1EB: dout  = 8'b11100000; //  491 : 224 - 0xe0
      12'h1EC: dout  = 8'b11001000; //  492 : 200 - 0xc8
      12'h1ED: dout  = 8'b00010100; //  493 :  20 - 0x14
      12'h1EE: dout  = 8'b10101000; //  494 : 168 - 0xa8
      12'h1EF: dout  = 8'b01010100; //  495 :  84 - 0x54
      12'h1F0: dout  = 8'b00000000; //  496 :   0 - 0x0 -- Sprite 0x1f
      12'h1F1: dout  = 8'b00111000; //  497 :  56 - 0x38
      12'h1F2: dout  = 8'b11000110; //  498 : 198 - 0xc6
      12'h1F3: dout  = 8'b11001011; //  499 : 203 - 0xcb
      12'h1F4: dout  = 8'b11011100; //  500 : 220 - 0xdc
      12'h1F5: dout  = 8'b00111010; //  501 :  58 - 0x3a
      12'h1F6: dout  = 8'b10011010; //  502 : 154 - 0x9a
      12'h1F7: dout  = 8'b11100001; //  503 : 225 - 0xe1
      12'h1F8: dout  = 8'b00000000; //  504 :   0 - 0x0 -- plane 1
      12'h1F9: dout  = 8'b00000000; //  505 :   0 - 0x0
      12'h1FA: dout  = 8'b00111000; //  506 :  56 - 0x38
      12'h1FB: dout  = 8'b10110100; //  507 : 180 - 0xb4
      12'h1FC: dout  = 8'b10101000; //  508 : 168 - 0xa8
      12'h1FD: dout  = 8'b11010100; //  509 : 212 - 0xd4
      12'h1FE: dout  = 8'b01110100; //  510 : 116 - 0x74
      12'h1FF: dout  = 8'b00011110; //  511 :  30 - 0x1e
      12'h200: dout  = 8'b00000000; //  512 :   0 - 0x0 -- Sprite 0x20
      12'h201: dout  = 8'b00011100; //  513 :  28 - 0x1c
      12'h202: dout  = 8'b00010011; //  514 :  19 - 0x13
      12'h203: dout  = 8'b00001000; //  515 :   8 - 0x8
      12'h204: dout  = 8'b00010000; //  516 :  16 - 0x10
      12'h205: dout  = 8'b00001000; //  517 :   8 - 0x8
      12'h206: dout  = 8'b00010000; //  518 :  16 - 0x10
      12'h207: dout  = 8'b00010000; //  519 :  16 - 0x10
      12'h208: dout  = 8'b00000000; //  520 :   0 - 0x0 -- plane 1
      12'h209: dout  = 8'b00000000; //  521 :   0 - 0x0
      12'h20A: dout  = 8'b00001100; //  522 :  12 - 0xc
      12'h20B: dout  = 8'b00000111; //  523 :   7 - 0x7
      12'h20C: dout  = 8'b00001111; //  524 :  15 - 0xf
      12'h20D: dout  = 8'b00000111; //  525 :   7 - 0x7
      12'h20E: dout  = 8'b00001111; //  526 :  15 - 0xf
      12'h20F: dout  = 8'b00001111; //  527 :  15 - 0xf
      12'h210: dout  = 8'b00000000; //  528 :   0 - 0x0 -- Sprite 0x21
      12'h211: dout  = 8'b00111000; //  529 :  56 - 0x38
      12'h212: dout  = 8'b11001000; //  530 : 200 - 0xc8
      12'h213: dout  = 8'b00010000; //  531 :  16 - 0x10
      12'h214: dout  = 8'b00001000; //  532 :   8 - 0x8
      12'h215: dout  = 8'b00010000; //  533 :  16 - 0x10
      12'h216: dout  = 8'b00001000; //  534 :   8 - 0x8
      12'h217: dout  = 8'b00001000; //  535 :   8 - 0x8
      12'h218: dout  = 8'b00000000; //  536 :   0 - 0x0 -- plane 1
      12'h219: dout  = 8'b00000000; //  537 :   0 - 0x0
      12'h21A: dout  = 8'b00110000; //  538 :  48 - 0x30
      12'h21B: dout  = 8'b11100000; //  539 : 224 - 0xe0
      12'h21C: dout  = 8'b11110000; //  540 : 240 - 0xf0
      12'h21D: dout  = 8'b11100000; //  541 : 224 - 0xe0
      12'h21E: dout  = 8'b11110000; //  542 : 240 - 0xf0
      12'h21F: dout  = 8'b11110000; //  543 : 240 - 0xf0
      12'h220: dout  = 8'b00001000; //  544 :   8 - 0x8 -- Sprite 0x22
      12'h221: dout  = 8'b00011100; //  545 :  28 - 0x1c
      12'h222: dout  = 8'b00100111; //  546 :  39 - 0x27
      12'h223: dout  = 8'b00101111; //  547 :  47 - 0x2f
      12'h224: dout  = 8'b00011111; //  548 :  31 - 0x1f
      12'h225: dout  = 8'b00001111; //  549 :  15 - 0xf
      12'h226: dout  = 8'b00001111; //  550 :  15 - 0xf
      12'h227: dout  = 8'b00001111; //  551 :  15 - 0xf
      12'h228: dout  = 8'b00000111; //  552 :   7 - 0x7 -- plane 1
      12'h229: dout  = 8'b00000011; //  553 :   3 - 0x3
      12'h22A: dout  = 8'b00011000; //  554 :  24 - 0x18
      12'h22B: dout  = 8'b00010101; //  555 :  21 - 0x15
      12'h22C: dout  = 8'b00000010; //  556 :   2 - 0x2
      12'h22D: dout  = 8'b00000101; //  557 :   5 - 0x5
      12'h22E: dout  = 8'b00000010; //  558 :   2 - 0x2
      12'h22F: dout  = 8'b00000100; //  559 :   4 - 0x4
      12'h230: dout  = 8'b00010000; //  560 :  16 - 0x10 -- Sprite 0x23
      12'h231: dout  = 8'b00111100; //  561 :  60 - 0x3c
      12'h232: dout  = 8'b11000010; //  562 : 194 - 0xc2
      12'h233: dout  = 8'b10000010; //  563 : 130 - 0x82
      12'h234: dout  = 8'b10000010; //  564 : 130 - 0x82
      12'h235: dout  = 8'b10000010; //  565 : 130 - 0x82
      12'h236: dout  = 8'b00010010; //  566 :  18 - 0x12
      12'h237: dout  = 8'b00011100; //  567 :  28 - 0x1c
      12'h238: dout  = 8'b11100000; //  568 : 224 - 0xe0 -- plane 1
      12'h239: dout  = 8'b11000000; //  569 : 192 - 0xc0
      12'h23A: dout  = 8'b00111100; //  570 :  60 - 0x3c
      12'h23B: dout  = 8'b01111100; //  571 : 124 - 0x7c
      12'h23C: dout  = 8'b01111100; //  572 : 124 - 0x7c
      12'h23D: dout  = 8'b01111100; //  573 : 124 - 0x7c
      12'h23E: dout  = 8'b11101100; //  574 : 236 - 0xec
      12'h23F: dout  = 8'b11100000; //  575 : 224 - 0xe0
      12'h240: dout  = 8'b00001111; //  576 :  15 - 0xf -- Sprite 0x24
      12'h241: dout  = 8'b00001110; //  577 :  14 - 0xe
      12'h242: dout  = 8'b00010100; //  578 :  20 - 0x14
      12'h243: dout  = 8'b00010100; //  579 :  20 - 0x14
      12'h244: dout  = 8'b00010010; //  580 :  18 - 0x12
      12'h245: dout  = 8'b00100101; //  581 :  37 - 0x25
      12'h246: dout  = 8'b01000100; //  582 :  68 - 0x44
      12'h247: dout  = 8'b00111000; //  583 :  56 - 0x38
      12'h248: dout  = 8'b00000010; //  584 :   2 - 0x2 -- plane 1
      12'h249: dout  = 8'b00000101; //  585 :   5 - 0x5
      12'h24A: dout  = 8'b00001011; //  586 :  11 - 0xb
      12'h24B: dout  = 8'b00001011; //  587 :  11 - 0xb
      12'h24C: dout  = 8'b00001101; //  588 :  13 - 0xd
      12'h24D: dout  = 8'b00011000; //  589 :  24 - 0x18
      12'h24E: dout  = 8'b00111000; //  590 :  56 - 0x38
      12'h24F: dout  = 8'b00000000; //  591 :   0 - 0x0
      12'h250: dout  = 8'b00010000; //  592 :  16 - 0x10 -- Sprite 0x25
      12'h251: dout  = 8'b00010000; //  593 :  16 - 0x10
      12'h252: dout  = 8'b00010000; //  594 :  16 - 0x10
      12'h253: dout  = 8'b00101100; //  595 :  44 - 0x2c
      12'h254: dout  = 8'b01000100; //  596 :  68 - 0x44
      12'h255: dout  = 8'b11000100; //  597 : 196 - 0xc4
      12'h256: dout  = 8'b00111000; //  598 :  56 - 0x38
      12'h257: dout  = 8'b00000000; //  599 :   0 - 0x0
      12'h258: dout  = 8'b11100000; //  600 : 224 - 0xe0 -- plane 1
      12'h259: dout  = 8'b11100000; //  601 : 224 - 0xe0
      12'h25A: dout  = 8'b11100000; //  602 : 224 - 0xe0
      12'h25B: dout  = 8'b11010000; //  603 : 208 - 0xd0
      12'h25C: dout  = 8'b10111000; //  604 : 184 - 0xb8
      12'h25D: dout  = 8'b00111000; //  605 :  56 - 0x38
      12'h25E: dout  = 8'b00000000; //  606 :   0 - 0x0
      12'h25F: dout  = 8'b00000000; //  607 :   0 - 0x0
      12'h260: dout  = 8'b00000000; //  608 :   0 - 0x0 -- Sprite 0x26
      12'h261: dout  = 8'b00000000; //  609 :   0 - 0x0
      12'h262: dout  = 8'b00000000; //  610 :   0 - 0x0
      12'h263: dout  = 8'b00000000; //  611 :   0 - 0x0
      12'h264: dout  = 8'b00000000; //  612 :   0 - 0x0
      12'h265: dout  = 8'b00000000; //  613 :   0 - 0x0
      12'h266: dout  = 8'b00000000; //  614 :   0 - 0x0
      12'h267: dout  = 8'b00000000; //  615 :   0 - 0x0
      12'h268: dout  = 8'b00000000; //  616 :   0 - 0x0 -- plane 1
      12'h269: dout  = 8'b00000000; //  617 :   0 - 0x0
      12'h26A: dout  = 8'b00000000; //  618 :   0 - 0x0
      12'h26B: dout  = 8'b00000000; //  619 :   0 - 0x0
      12'h26C: dout  = 8'b00000000; //  620 :   0 - 0x0
      12'h26D: dout  = 8'b00000000; //  621 :   0 - 0x0
      12'h26E: dout  = 8'b00000000; //  622 :   0 - 0x0
      12'h26F: dout  = 8'b00000000; //  623 :   0 - 0x0
      12'h270: dout  = 8'b00000000; //  624 :   0 - 0x0 -- Sprite 0x27
      12'h271: dout  = 8'b00000000; //  625 :   0 - 0x0
      12'h272: dout  = 8'b00000000; //  626 :   0 - 0x0
      12'h273: dout  = 8'b00000000; //  627 :   0 - 0x0
      12'h274: dout  = 8'b00000000; //  628 :   0 - 0x0
      12'h275: dout  = 8'b00000000; //  629 :   0 - 0x0
      12'h276: dout  = 8'b00000000; //  630 :   0 - 0x0
      12'h277: dout  = 8'b00000000; //  631 :   0 - 0x0
      12'h278: dout  = 8'b00000000; //  632 :   0 - 0x0 -- plane 1
      12'h279: dout  = 8'b00000000; //  633 :   0 - 0x0
      12'h27A: dout  = 8'b00000000; //  634 :   0 - 0x0
      12'h27B: dout  = 8'b00000000; //  635 :   0 - 0x0
      12'h27C: dout  = 8'b00000000; //  636 :   0 - 0x0
      12'h27D: dout  = 8'b00000000; //  637 :   0 - 0x0
      12'h27E: dout  = 8'b00000000; //  638 :   0 - 0x0
      12'h27F: dout  = 8'b00000000; //  639 :   0 - 0x0
      12'h280: dout  = 8'b00000000; //  640 :   0 - 0x0 -- Sprite 0x28
      12'h281: dout  = 8'b00000000; //  641 :   0 - 0x0
      12'h282: dout  = 8'b00000000; //  642 :   0 - 0x0
      12'h283: dout  = 8'b00000000; //  643 :   0 - 0x0
      12'h284: dout  = 8'b00000000; //  644 :   0 - 0x0
      12'h285: dout  = 8'b00000000; //  645 :   0 - 0x0
      12'h286: dout  = 8'b00000000; //  646 :   0 - 0x0
      12'h287: dout  = 8'b00000000; //  647 :   0 - 0x0
      12'h288: dout  = 8'b00000000; //  648 :   0 - 0x0 -- plane 1
      12'h289: dout  = 8'b00000000; //  649 :   0 - 0x0
      12'h28A: dout  = 8'b00000000; //  650 :   0 - 0x0
      12'h28B: dout  = 8'b00000000; //  651 :   0 - 0x0
      12'h28C: dout  = 8'b00000000; //  652 :   0 - 0x0
      12'h28D: dout  = 8'b00000000; //  653 :   0 - 0x0
      12'h28E: dout  = 8'b00000000; //  654 :   0 - 0x0
      12'h28F: dout  = 8'b00000000; //  655 :   0 - 0x0
      12'h290: dout  = 8'b00100000; //  656 :  32 - 0x20 -- Sprite 0x29
      12'h291: dout  = 8'b00100000; //  657 :  32 - 0x20
      12'h292: dout  = 8'b00100000; //  658 :  32 - 0x20
      12'h293: dout  = 8'b00100000; //  659 :  32 - 0x20
      12'h294: dout  = 8'b00010011; //  660 :  19 - 0x13
      12'h295: dout  = 8'b00001101; //  661 :  13 - 0xd
      12'h296: dout  = 8'b00000010; //  662 :   2 - 0x2
      12'h297: dout  = 8'b00000001; //  663 :   1 - 0x1
      12'h298: dout  = 8'b00011111; //  664 :  31 - 0x1f -- plane 1
      12'h299: dout  = 8'b00011111; //  665 :  31 - 0x1f
      12'h29A: dout  = 8'b00011111; //  666 :  31 - 0x1f
      12'h29B: dout  = 8'b00011111; //  667 :  31 - 0x1f
      12'h29C: dout  = 8'b00001100; //  668 :  12 - 0xc
      12'h29D: dout  = 8'b00000000; //  669 :   0 - 0x0
      12'h29E: dout  = 8'b00000001; //  670 :   1 - 0x1
      12'h29F: dout  = 8'b00000000; //  671 :   0 - 0x0
      12'h2A0: dout  = 8'b00100000; //  672 :  32 - 0x20 -- Sprite 0x2a
      12'h2A1: dout  = 8'b00100000; //  673 :  32 - 0x20
      12'h2A2: dout  = 8'b00100000; //  674 :  32 - 0x20
      12'h2A3: dout  = 8'b00100000; //  675 :  32 - 0x20
      12'h2A4: dout  = 8'b00010011; //  676 :  19 - 0x13
      12'h2A5: dout  = 8'b00001101; //  677 :  13 - 0xd
      12'h2A6: dout  = 8'b00000001; //  678 :   1 - 0x1
      12'h2A7: dout  = 8'b00000001; //  679 :   1 - 0x1
      12'h2A8: dout  = 8'b00011111; //  680 :  31 - 0x1f -- plane 1
      12'h2A9: dout  = 8'b00011111; //  681 :  31 - 0x1f
      12'h2AA: dout  = 8'b00011111; //  682 :  31 - 0x1f
      12'h2AB: dout  = 8'b00011111; //  683 :  31 - 0x1f
      12'h2AC: dout  = 8'b00001100; //  684 :  12 - 0xc
      12'h2AD: dout  = 8'b00000000; //  685 :   0 - 0x0
      12'h2AE: dout  = 8'b00000000; //  686 :   0 - 0x0
      12'h2AF: dout  = 8'b00000000; //  687 :   0 - 0x0
      12'h2B0: dout  = 8'b00000000; //  688 :   0 - 0x0 -- Sprite 0x2b
      12'h2B1: dout  = 8'b00000000; //  689 :   0 - 0x0
      12'h2B2: dout  = 8'b00000000; //  690 :   0 - 0x0
      12'h2B3: dout  = 8'b00000000; //  691 :   0 - 0x0
      12'h2B4: dout  = 8'b00000000; //  692 :   0 - 0x0
      12'h2B5: dout  = 8'b00000000; //  693 :   0 - 0x0
      12'h2B6: dout  = 8'b00000000; //  694 :   0 - 0x0
      12'h2B7: dout  = 8'b00000000; //  695 :   0 - 0x0
      12'h2B8: dout  = 8'b00000000; //  696 :   0 - 0x0 -- plane 1
      12'h2B9: dout  = 8'b00000000; //  697 :   0 - 0x0
      12'h2BA: dout  = 8'b00000000; //  698 :   0 - 0x0
      12'h2BB: dout  = 8'b00000000; //  699 :   0 - 0x0
      12'h2BC: dout  = 8'b00000000; //  700 :   0 - 0x0
      12'h2BD: dout  = 8'b00000000; //  701 :   0 - 0x0
      12'h2BE: dout  = 8'b00000000; //  702 :   0 - 0x0
      12'h2BF: dout  = 8'b00000000; //  703 :   0 - 0x0
      12'h2C0: dout  = 8'b00000000; //  704 :   0 - 0x0 -- Sprite 0x2c
      12'h2C1: dout  = 8'b00000000; //  705 :   0 - 0x0
      12'h2C2: dout  = 8'b00000000; //  706 :   0 - 0x0
      12'h2C3: dout  = 8'b00000000; //  707 :   0 - 0x0
      12'h2C4: dout  = 8'b00000000; //  708 :   0 - 0x0
      12'h2C5: dout  = 8'b00000000; //  709 :   0 - 0x0
      12'h2C6: dout  = 8'b00000000; //  710 :   0 - 0x0
      12'h2C7: dout  = 8'b00000000; //  711 :   0 - 0x0
      12'h2C8: dout  = 8'b00000000; //  712 :   0 - 0x0 -- plane 1
      12'h2C9: dout  = 8'b00000000; //  713 :   0 - 0x0
      12'h2CA: dout  = 8'b00000000; //  714 :   0 - 0x0
      12'h2CB: dout  = 8'b00000000; //  715 :   0 - 0x0
      12'h2CC: dout  = 8'b00000000; //  716 :   0 - 0x0
      12'h2CD: dout  = 8'b00000000; //  717 :   0 - 0x0
      12'h2CE: dout  = 8'b00000000; //  718 :   0 - 0x0
      12'h2CF: dout  = 8'b00000000; //  719 :   0 - 0x0
      12'h2D0: dout  = 8'b00111100; //  720 :  60 - 0x3c -- Sprite 0x2d
      12'h2D1: dout  = 8'b00000000; //  721 :   0 - 0x0
      12'h2D2: dout  = 8'b10000001; //  722 : 129 - 0x81
      12'h2D3: dout  = 8'b10011001; //  723 : 153 - 0x99
      12'h2D4: dout  = 8'b10011001; //  724 : 153 - 0x99
      12'h2D5: dout  = 8'b10000001; //  725 : 129 - 0x81
      12'h2D6: dout  = 8'b00000000; //  726 :   0 - 0x0
      12'h2D7: dout  = 8'b00111100; //  727 :  60 - 0x3c
      12'h2D8: dout  = 8'b00000000; //  728 :   0 - 0x0 -- plane 1
      12'h2D9: dout  = 8'b01111110; //  729 : 126 - 0x7e
      12'h2DA: dout  = 8'b01000010; //  730 :  66 - 0x42
      12'h2DB: dout  = 8'b01000010; //  731 :  66 - 0x42
      12'h2DC: dout  = 8'b01000010; //  732 :  66 - 0x42
      12'h2DD: dout  = 8'b01000010; //  733 :  66 - 0x42
      12'h2DE: dout  = 8'b01111110; //  734 : 126 - 0x7e
      12'h2DF: dout  = 8'b00000000; //  735 :   0 - 0x0
      12'h2E0: dout  = 8'b00000000; //  736 :   0 - 0x0 -- Sprite 0x2e
      12'h2E1: dout  = 8'b00000000; //  737 :   0 - 0x0
      12'h2E2: dout  = 8'b00000000; //  738 :   0 - 0x0
      12'h2E3: dout  = 8'b00000000; //  739 :   0 - 0x0
      12'h2E4: dout  = 8'b00000000; //  740 :   0 - 0x0
      12'h2E5: dout  = 8'b00000000; //  741 :   0 - 0x0
      12'h2E6: dout  = 8'b00000000; //  742 :   0 - 0x0
      12'h2E7: dout  = 8'b00000000; //  743 :   0 - 0x0
      12'h2E8: dout  = 8'b00000000; //  744 :   0 - 0x0 -- plane 1
      12'h2E9: dout  = 8'b00000000; //  745 :   0 - 0x0
      12'h2EA: dout  = 8'b00000000; //  746 :   0 - 0x0
      12'h2EB: dout  = 8'b00000000; //  747 :   0 - 0x0
      12'h2EC: dout  = 8'b00000000; //  748 :   0 - 0x0
      12'h2ED: dout  = 8'b00000000; //  749 :   0 - 0x0
      12'h2EE: dout  = 8'b00000000; //  750 :   0 - 0x0
      12'h2EF: dout  = 8'b00000000; //  751 :   0 - 0x0
      12'h2F0: dout  = 8'b10011111; //  752 : 159 - 0x9f -- Sprite 0x2f
      12'h2F1: dout  = 8'b10011110; //  753 : 158 - 0x9e
      12'h2F2: dout  = 8'b10011100; //  754 : 156 - 0x9c
      12'h2F3: dout  = 8'b00011000; //  755 :  24 - 0x18
      12'h2F4: dout  = 8'b00111000; //  756 :  56 - 0x38
      12'h2F5: dout  = 8'b11111100; //  757 : 252 - 0xfc
      12'h2F6: dout  = 8'b11111100; //  758 : 252 - 0xfc
      12'h2F7: dout  = 8'b11111100; //  759 : 252 - 0xfc
      12'h2F8: dout  = 8'b01100110; //  760 : 102 - 0x66 -- plane 1
      12'h2F9: dout  = 8'b01100000; //  761 :  96 - 0x60
      12'h2FA: dout  = 8'b01101000; //  762 : 104 - 0x68
      12'h2FB: dout  = 8'b11100000; //  763 : 224 - 0xe0
      12'h2FC: dout  = 8'b11000000; //  764 : 192 - 0xc0
      12'h2FD: dout  = 8'b00010000; //  765 :  16 - 0x10
      12'h2FE: dout  = 8'b00101000; //  766 :  40 - 0x28
      12'h2FF: dout  = 8'b01010000; //  767 :  80 - 0x50
      12'h300: dout  = 8'b01111111; //  768 : 127 - 0x7f -- Sprite 0x30
      12'h301: dout  = 8'b01111110; //  769 : 126 - 0x7e
      12'h302: dout  = 8'b11111100; //  770 : 252 - 0xfc
      12'h303: dout  = 8'b00111000; //  771 :  56 - 0x38
      12'h304: dout  = 8'b00111000; //  772 :  56 - 0x38
      12'h305: dout  = 8'b00000100; //  773 :   4 - 0x4
      12'h306: dout  = 8'b10000100; //  774 : 132 - 0x84
      12'h307: dout  = 8'b11111100; //  775 : 252 - 0xfc
      12'h308: dout  = 8'b11110110; //  776 : 246 - 0xf6 -- plane 1
      12'h309: dout  = 8'b11110000; //  777 : 240 - 0xf0
      12'h30A: dout  = 8'b00111000; //  778 :  56 - 0x38
      12'h30B: dout  = 8'b11010000; //  779 : 208 - 0xd0
      12'h30C: dout  = 8'b11000000; //  780 : 192 - 0xc0
      12'h30D: dout  = 8'b11111000; //  781 : 248 - 0xf8
      12'h30E: dout  = 8'b01111000; //  782 : 120 - 0x78
      12'h30F: dout  = 8'b00000000; //  783 :   0 - 0x0
      12'h310: dout  = 8'b01111111; //  784 : 127 - 0x7f -- Sprite 0x31
      12'h311: dout  = 8'b01111110; //  785 : 126 - 0x7e
      12'h312: dout  = 8'b11111100; //  786 : 252 - 0xfc
      12'h313: dout  = 8'b00111000; //  787 :  56 - 0x38
      12'h314: dout  = 8'b00111000; //  788 :  56 - 0x38
      12'h315: dout  = 8'b00011100; //  789 :  28 - 0x1c
      12'h316: dout  = 8'b10000100; //  790 : 132 - 0x84
      12'h317: dout  = 8'b11000100; //  791 : 196 - 0xc4
      12'h318: dout  = 8'b11110110; //  792 : 246 - 0xf6 -- plane 1
      12'h319: dout  = 8'b11110000; //  793 : 240 - 0xf0
      12'h31A: dout  = 8'b00111000; //  794 :  56 - 0x38
      12'h31B: dout  = 8'b11010000; //  795 : 208 - 0xd0
      12'h31C: dout  = 8'b11000000; //  796 : 192 - 0xc0
      12'h31D: dout  = 8'b11100000; //  797 : 224 - 0xe0
      12'h31E: dout  = 8'b01111000; //  798 : 120 - 0x78
      12'h31F: dout  = 8'b00111000; //  799 :  56 - 0x38
      12'h320: dout  = 8'b01111111; //  800 : 127 - 0x7f -- Sprite 0x32
      12'h321: dout  = 8'b01111110; //  801 : 126 - 0x7e
      12'h322: dout  = 8'b11111100; //  802 : 252 - 0xfc
      12'h323: dout  = 8'b00111000; //  803 :  56 - 0x38
      12'h324: dout  = 8'b00100100; //  804 :  36 - 0x24
      12'h325: dout  = 8'b00000100; //  805 :   4 - 0x4
      12'h326: dout  = 8'b10011100; //  806 : 156 - 0x9c
      12'h327: dout  = 8'b11111100; //  807 : 252 - 0xfc
      12'h328: dout  = 8'b11110110; //  808 : 246 - 0xf6 -- plane 1
      12'h329: dout  = 8'b11110000; //  809 : 240 - 0xf0
      12'h32A: dout  = 8'b00111000; //  810 :  56 - 0x38
      12'h32B: dout  = 8'b11000000; //  811 : 192 - 0xc0
      12'h32C: dout  = 8'b11011000; //  812 : 216 - 0xd8
      12'h32D: dout  = 8'b11111000; //  813 : 248 - 0xf8
      12'h32E: dout  = 8'b01100000; //  814 :  96 - 0x60
      12'h32F: dout  = 8'b00010000; //  815 :  16 - 0x10
      12'h330: dout  = 8'b00100011; //  816 :  35 - 0x23 -- Sprite 0x33
      12'h331: dout  = 8'b00100011; //  817 :  35 - 0x23
      12'h332: dout  = 8'b00100001; //  818 :  33 - 0x21
      12'h333: dout  = 8'b00100000; //  819 :  32 - 0x20
      12'h334: dout  = 8'b00010011; //  820 :  19 - 0x13
      12'h335: dout  = 8'b00001101; //  821 :  13 - 0xd
      12'h336: dout  = 8'b00000001; //  822 :   1 - 0x1
      12'h337: dout  = 8'b00000001; //  823 :   1 - 0x1
      12'h338: dout  = 8'b00011100; //  824 :  28 - 0x1c -- plane 1
      12'h339: dout  = 8'b00011100; //  825 :  28 - 0x1c
      12'h33A: dout  = 8'b00011110; //  826 :  30 - 0x1e
      12'h33B: dout  = 8'b00011111; //  827 :  31 - 0x1f
      12'h33C: dout  = 8'b00001100; //  828 :  12 - 0xc
      12'h33D: dout  = 8'b00000000; //  829 :   0 - 0x0
      12'h33E: dout  = 8'b00000000; //  830 :   0 - 0x0
      12'h33F: dout  = 8'b00000000; //  831 :   0 - 0x0
      12'h340: dout  = 8'b11111100; //  832 : 252 - 0xfc -- Sprite 0x34
      12'h341: dout  = 8'b11111100; //  833 : 252 - 0xfc
      12'h342: dout  = 8'b11111100; //  834 : 252 - 0xfc
      12'h343: dout  = 8'b11111100; //  835 : 252 - 0xfc
      12'h344: dout  = 8'b10100100; //  836 : 164 - 0xa4
      12'h345: dout  = 8'b00100100; //  837 :  36 - 0x24
      12'h346: dout  = 8'b00010010; //  838 :  18 - 0x12
      12'h347: dout  = 8'b11101110; //  839 : 238 - 0xee
      12'h348: dout  = 8'b10000000; //  840 : 128 - 0x80 -- plane 1
      12'h349: dout  = 8'b01010000; //  841 :  80 - 0x50
      12'h34A: dout  = 8'b10101000; //  842 : 168 - 0xa8
      12'h34B: dout  = 8'b00000000; //  843 :   0 - 0x0
      12'h34C: dout  = 8'b01011000; //  844 :  88 - 0x58
      12'h34D: dout  = 8'b11011000; //  845 : 216 - 0xd8
      12'h34E: dout  = 8'b11101100; //  846 : 236 - 0xec
      12'h34F: dout  = 8'b00000000; //  847 :   0 - 0x0
      12'h350: dout  = 8'b00100011; //  848 :  35 - 0x23 -- Sprite 0x35
      12'h351: dout  = 8'b00100011; //  849 :  35 - 0x23
      12'h352: dout  = 8'b00100001; //  850 :  33 - 0x21
      12'h353: dout  = 8'b00100000; //  851 :  32 - 0x20
      12'h354: dout  = 8'b00010011; //  852 :  19 - 0x13
      12'h355: dout  = 8'b00001110; //  853 :  14 - 0xe
      12'h356: dout  = 8'b00000010; //  854 :   2 - 0x2
      12'h357: dout  = 8'b00000001; //  855 :   1 - 0x1
      12'h358: dout  = 8'b00011100; //  856 :  28 - 0x1c -- plane 1
      12'h359: dout  = 8'b00011100; //  857 :  28 - 0x1c
      12'h35A: dout  = 8'b00011110; //  858 :  30 - 0x1e
      12'h35B: dout  = 8'b00011111; //  859 :  31 - 0x1f
      12'h35C: dout  = 8'b00001100; //  860 :  12 - 0xc
      12'h35D: dout  = 8'b00000001; //  861 :   1 - 0x1
      12'h35E: dout  = 8'b00000001; //  862 :   1 - 0x1
      12'h35F: dout  = 8'b00000000; //  863 :   0 - 0x0
      12'h360: dout  = 8'b11111100; //  864 : 252 - 0xfc -- Sprite 0x36
      12'h361: dout  = 8'b11111100; //  865 : 252 - 0xfc
      12'h362: dout  = 8'b11111100; //  866 : 252 - 0xfc
      12'h363: dout  = 8'b11111100; //  867 : 252 - 0xfc
      12'h364: dout  = 8'b10100110; //  868 : 166 - 0xa6
      12'h365: dout  = 8'b00110001; //  869 :  49 - 0x31
      12'h366: dout  = 8'b01001001; //  870 :  73 - 0x49
      12'h367: dout  = 8'b11000110; //  871 : 198 - 0xc6
      12'h368: dout  = 8'b10101000; //  872 : 168 - 0xa8 -- plane 1
      12'h369: dout  = 8'b01010000; //  873 :  80 - 0x50
      12'h36A: dout  = 8'b10101000; //  874 : 168 - 0xa8
      12'h36B: dout  = 8'b00000000; //  875 :   0 - 0x0
      12'h36C: dout  = 8'b01011000; //  876 :  88 - 0x58
      12'h36D: dout  = 8'b11001110; //  877 : 206 - 0xce
      12'h36E: dout  = 8'b10000110; //  878 : 134 - 0x86
      12'h36F: dout  = 8'b00000000; //  879 :   0 - 0x0
      12'h370: dout  = 8'b11111100; //  880 : 252 - 0xfc -- Sprite 0x37
      12'h371: dout  = 8'b11111100; //  881 : 252 - 0xfc
      12'h372: dout  = 8'b11111100; //  882 : 252 - 0xfc
      12'h373: dout  = 8'b11111100; //  883 : 252 - 0xfc
      12'h374: dout  = 8'b10100100; //  884 : 164 - 0xa4
      12'h375: dout  = 8'b00100100; //  885 :  36 - 0x24
      12'h376: dout  = 8'b00010010; //  886 :  18 - 0x12
      12'h377: dout  = 8'b11101110; //  887 : 238 - 0xee
      12'h378: dout  = 8'b10101000; //  888 : 168 - 0xa8 -- plane 1
      12'h379: dout  = 8'b01010000; //  889 :  80 - 0x50
      12'h37A: dout  = 8'b10101000; //  890 : 168 - 0xa8
      12'h37B: dout  = 8'b00000000; //  891 :   0 - 0x0
      12'h37C: dout  = 8'b01011000; //  892 :  88 - 0x58
      12'h37D: dout  = 8'b11011000; //  893 : 216 - 0xd8
      12'h37E: dout  = 8'b11101100; //  894 : 236 - 0xec
      12'h37F: dout  = 8'b00000000; //  895 :   0 - 0x0
      12'h380: dout  = 8'b00000000; //  896 :   0 - 0x0 -- Sprite 0x38
      12'h381: dout  = 8'b00000000; //  897 :   0 - 0x0
      12'h382: dout  = 8'b00000000; //  898 :   0 - 0x0
      12'h383: dout  = 8'b00000000; //  899 :   0 - 0x0
      12'h384: dout  = 8'b00000000; //  900 :   0 - 0x0
      12'h385: dout  = 8'b00000000; //  901 :   0 - 0x0
      12'h386: dout  = 8'b00000000; //  902 :   0 - 0x0
      12'h387: dout  = 8'b00000000; //  903 :   0 - 0x0
      12'h388: dout  = 8'b00000000; //  904 :   0 - 0x0 -- plane 1
      12'h389: dout  = 8'b00000000; //  905 :   0 - 0x0
      12'h38A: dout  = 8'b00000000; //  906 :   0 - 0x0
      12'h38B: dout  = 8'b00000000; //  907 :   0 - 0x0
      12'h38C: dout  = 8'b00000000; //  908 :   0 - 0x0
      12'h38D: dout  = 8'b00000000; //  909 :   0 - 0x0
      12'h38E: dout  = 8'b00000000; //  910 :   0 - 0x0
      12'h38F: dout  = 8'b00000000; //  911 :   0 - 0x0
      12'h390: dout  = 8'b00000000; //  912 :   0 - 0x0 -- Sprite 0x39
      12'h391: dout  = 8'b00000000; //  913 :   0 - 0x0
      12'h392: dout  = 8'b00000000; //  914 :   0 - 0x0
      12'h393: dout  = 8'b00000000; //  915 :   0 - 0x0
      12'h394: dout  = 8'b00000000; //  916 :   0 - 0x0
      12'h395: dout  = 8'b00000000; //  917 :   0 - 0x0
      12'h396: dout  = 8'b00000000; //  918 :   0 - 0x0
      12'h397: dout  = 8'b00000000; //  919 :   0 - 0x0
      12'h398: dout  = 8'b00000000; //  920 :   0 - 0x0 -- plane 1
      12'h399: dout  = 8'b00000000; //  921 :   0 - 0x0
      12'h39A: dout  = 8'b00000000; //  922 :   0 - 0x0
      12'h39B: dout  = 8'b00000000; //  923 :   0 - 0x0
      12'h39C: dout  = 8'b00000000; //  924 :   0 - 0x0
      12'h39D: dout  = 8'b00000000; //  925 :   0 - 0x0
      12'h39E: dout  = 8'b00000000; //  926 :   0 - 0x0
      12'h39F: dout  = 8'b00000000; //  927 :   0 - 0x0
      12'h3A0: dout  = 8'b00000000; //  928 :   0 - 0x0 -- Sprite 0x3a
      12'h3A1: dout  = 8'b00000000; //  929 :   0 - 0x0
      12'h3A2: dout  = 8'b00000000; //  930 :   0 - 0x0
      12'h3A3: dout  = 8'b00000000; //  931 :   0 - 0x0
      12'h3A4: dout  = 8'b00000000; //  932 :   0 - 0x0
      12'h3A5: dout  = 8'b00000000; //  933 :   0 - 0x0
      12'h3A6: dout  = 8'b00000000; //  934 :   0 - 0x0
      12'h3A7: dout  = 8'b00000000; //  935 :   0 - 0x0
      12'h3A8: dout  = 8'b00000000; //  936 :   0 - 0x0 -- plane 1
      12'h3A9: dout  = 8'b00000000; //  937 :   0 - 0x0
      12'h3AA: dout  = 8'b00000000; //  938 :   0 - 0x0
      12'h3AB: dout  = 8'b00000000; //  939 :   0 - 0x0
      12'h3AC: dout  = 8'b00000000; //  940 :   0 - 0x0
      12'h3AD: dout  = 8'b00000000; //  941 :   0 - 0x0
      12'h3AE: dout  = 8'b00000000; //  942 :   0 - 0x0
      12'h3AF: dout  = 8'b00000000; //  943 :   0 - 0x0
      12'h3B0: dout  = 8'b00000000; //  944 :   0 - 0x0 -- Sprite 0x3b
      12'h3B1: dout  = 8'b00000000; //  945 :   0 - 0x0
      12'h3B2: dout  = 8'b00000000; //  946 :   0 - 0x0
      12'h3B3: dout  = 8'b00000000; //  947 :   0 - 0x0
      12'h3B4: dout  = 8'b00000000; //  948 :   0 - 0x0
      12'h3B5: dout  = 8'b00000000; //  949 :   0 - 0x0
      12'h3B6: dout  = 8'b00000000; //  950 :   0 - 0x0
      12'h3B7: dout  = 8'b00000000; //  951 :   0 - 0x0
      12'h3B8: dout  = 8'b00000000; //  952 :   0 - 0x0 -- plane 1
      12'h3B9: dout  = 8'b00000000; //  953 :   0 - 0x0
      12'h3BA: dout  = 8'b00000000; //  954 :   0 - 0x0
      12'h3BB: dout  = 8'b00000000; //  955 :   0 - 0x0
      12'h3BC: dout  = 8'b00000000; //  956 :   0 - 0x0
      12'h3BD: dout  = 8'b00000000; //  957 :   0 - 0x0
      12'h3BE: dout  = 8'b00000000; //  958 :   0 - 0x0
      12'h3BF: dout  = 8'b00000000; //  959 :   0 - 0x0
      12'h3C0: dout  = 8'b00000000; //  960 :   0 - 0x0 -- Sprite 0x3c
      12'h3C1: dout  = 8'b00000000; //  961 :   0 - 0x0
      12'h3C2: dout  = 8'b00000000; //  962 :   0 - 0x0
      12'h3C3: dout  = 8'b00000000; //  963 :   0 - 0x0
      12'h3C4: dout  = 8'b00000000; //  964 :   0 - 0x0
      12'h3C5: dout  = 8'b00000000; //  965 :   0 - 0x0
      12'h3C6: dout  = 8'b00000000; //  966 :   0 - 0x0
      12'h3C7: dout  = 8'b00000000; //  967 :   0 - 0x0
      12'h3C8: dout  = 8'b00000000; //  968 :   0 - 0x0 -- plane 1
      12'h3C9: dout  = 8'b00000000; //  969 :   0 - 0x0
      12'h3CA: dout  = 8'b00000000; //  970 :   0 - 0x0
      12'h3CB: dout  = 8'b00000000; //  971 :   0 - 0x0
      12'h3CC: dout  = 8'b00000000; //  972 :   0 - 0x0
      12'h3CD: dout  = 8'b00000000; //  973 :   0 - 0x0
      12'h3CE: dout  = 8'b00000000; //  974 :   0 - 0x0
      12'h3CF: dout  = 8'b00000000; //  975 :   0 - 0x0
      12'h3D0: dout  = 8'b00000000; //  976 :   0 - 0x0 -- Sprite 0x3d
      12'h3D1: dout  = 8'b00000000; //  977 :   0 - 0x0
      12'h3D2: dout  = 8'b00000000; //  978 :   0 - 0x0
      12'h3D3: dout  = 8'b00000000; //  979 :   0 - 0x0
      12'h3D4: dout  = 8'b00000000; //  980 :   0 - 0x0
      12'h3D5: dout  = 8'b00000000; //  981 :   0 - 0x0
      12'h3D6: dout  = 8'b00000000; //  982 :   0 - 0x0
      12'h3D7: dout  = 8'b00000000; //  983 :   0 - 0x0
      12'h3D8: dout  = 8'b00000000; //  984 :   0 - 0x0 -- plane 1
      12'h3D9: dout  = 8'b00000000; //  985 :   0 - 0x0
      12'h3DA: dout  = 8'b00000000; //  986 :   0 - 0x0
      12'h3DB: dout  = 8'b00000000; //  987 :   0 - 0x0
      12'h3DC: dout  = 8'b00000000; //  988 :   0 - 0x0
      12'h3DD: dout  = 8'b00000000; //  989 :   0 - 0x0
      12'h3DE: dout  = 8'b00000000; //  990 :   0 - 0x0
      12'h3DF: dout  = 8'b00000000; //  991 :   0 - 0x0
      12'h3E0: dout  = 8'b00000000; //  992 :   0 - 0x0 -- Sprite 0x3e
      12'h3E1: dout  = 8'b00000000; //  993 :   0 - 0x0
      12'h3E2: dout  = 8'b00000000; //  994 :   0 - 0x0
      12'h3E3: dout  = 8'b00000000; //  995 :   0 - 0x0
      12'h3E4: dout  = 8'b00000000; //  996 :   0 - 0x0
      12'h3E5: dout  = 8'b00000000; //  997 :   0 - 0x0
      12'h3E6: dout  = 8'b00000000; //  998 :   0 - 0x0
      12'h3E7: dout  = 8'b00000000; //  999 :   0 - 0x0
      12'h3E8: dout  = 8'b00000000; // 1000 :   0 - 0x0 -- plane 1
      12'h3E9: dout  = 8'b00000000; // 1001 :   0 - 0x0
      12'h3EA: dout  = 8'b00000000; // 1002 :   0 - 0x0
      12'h3EB: dout  = 8'b00000000; // 1003 :   0 - 0x0
      12'h3EC: dout  = 8'b00000000; // 1004 :   0 - 0x0
      12'h3ED: dout  = 8'b00000000; // 1005 :   0 - 0x0
      12'h3EE: dout  = 8'b00000000; // 1006 :   0 - 0x0
      12'h3EF: dout  = 8'b00000000; // 1007 :   0 - 0x0
      12'h3F0: dout  = 8'b00000000; // 1008 :   0 - 0x0 -- Sprite 0x3f
      12'h3F1: dout  = 8'b00000000; // 1009 :   0 - 0x0
      12'h3F2: dout  = 8'b00000000; // 1010 :   0 - 0x0
      12'h3F3: dout  = 8'b00000000; // 1011 :   0 - 0x0
      12'h3F4: dout  = 8'b00000000; // 1012 :   0 - 0x0
      12'h3F5: dout  = 8'b00000000; // 1013 :   0 - 0x0
      12'h3F6: dout  = 8'b00000000; // 1014 :   0 - 0x0
      12'h3F7: dout  = 8'b00000000; // 1015 :   0 - 0x0
      12'h3F8: dout  = 8'b00000000; // 1016 :   0 - 0x0 -- plane 1
      12'h3F9: dout  = 8'b00000000; // 1017 :   0 - 0x0
      12'h3FA: dout  = 8'b00000000; // 1018 :   0 - 0x0
      12'h3FB: dout  = 8'b00000000; // 1019 :   0 - 0x0
      12'h3FC: dout  = 8'b00000000; // 1020 :   0 - 0x0
      12'h3FD: dout  = 8'b00000000; // 1021 :   0 - 0x0
      12'h3FE: dout  = 8'b00000000; // 1022 :   0 - 0x0
      12'h3FF: dout  = 8'b00000000; // 1023 :   0 - 0x0
      12'h400: dout  = 8'b00000000; // 1024 :   0 - 0x0 -- Sprite 0x40
      12'h401: dout  = 8'b00111110; // 1025 :  62 - 0x3e
      12'h402: dout  = 8'b01111111; // 1026 : 127 - 0x7f
      12'h403: dout  = 8'b01111111; // 1027 : 127 - 0x7f
      12'h404: dout  = 8'b01111111; // 1028 : 127 - 0x7f
      12'h405: dout  = 8'b01111111; // 1029 : 127 - 0x7f
      12'h406: dout  = 8'b01111111; // 1030 : 127 - 0x7f
      12'h407: dout  = 8'b00111110; // 1031 :  62 - 0x3e
      12'h408: dout  = 8'b00111100; // 1032 :  60 - 0x3c -- plane 1
      12'h409: dout  = 8'b01111100; // 1033 : 124 - 0x7c
      12'h40A: dout  = 8'b11100110; // 1034 : 230 - 0xe6
      12'h40B: dout  = 8'b11101110; // 1035 : 238 - 0xee
      12'h40C: dout  = 8'b11110110; // 1036 : 246 - 0xf6
      12'h40D: dout  = 8'b11100110; // 1037 : 230 - 0xe6
      12'h40E: dout  = 8'b00111100; // 1038 :  60 - 0x3c
      12'h40F: dout  = 8'b00000000; // 1039 :   0 - 0x0
      12'h410: dout  = 8'b00000000; // 1040 :   0 - 0x0 -- Sprite 0x41
      12'h411: dout  = 8'b00111100; // 1041 :  60 - 0x3c
      12'h412: dout  = 8'b00011100; // 1042 :  28 - 0x1c
      12'h413: dout  = 8'b00011100; // 1043 :  28 - 0x1c
      12'h414: dout  = 8'b00011100; // 1044 :  28 - 0x1c
      12'h415: dout  = 8'b00011100; // 1045 :  28 - 0x1c
      12'h416: dout  = 8'b00011100; // 1046 :  28 - 0x1c
      12'h417: dout  = 8'b00011100; // 1047 :  28 - 0x1c
      12'h418: dout  = 8'b00111000; // 1048 :  56 - 0x38 -- plane 1
      12'h419: dout  = 8'b01111000; // 1049 : 120 - 0x78
      12'h41A: dout  = 8'b00111000; // 1050 :  56 - 0x38
      12'h41B: dout  = 8'b00111000; // 1051 :  56 - 0x38
      12'h41C: dout  = 8'b00111000; // 1052 :  56 - 0x38
      12'h41D: dout  = 8'b00111000; // 1053 :  56 - 0x38
      12'h41E: dout  = 8'b00111000; // 1054 :  56 - 0x38
      12'h41F: dout  = 8'b00000000; // 1055 :   0 - 0x0
      12'h420: dout  = 8'b00000000; // 1056 :   0 - 0x0 -- Sprite 0x42
      12'h421: dout  = 8'b01111100; // 1057 : 124 - 0x7c
      12'h422: dout  = 8'b01111111; // 1058 : 127 - 0x7f
      12'h423: dout  = 8'b01100111; // 1059 : 103 - 0x67
      12'h424: dout  = 8'b00111111; // 1060 :  63 - 0x3f
      12'h425: dout  = 8'b01111110; // 1061 : 126 - 0x7e
      12'h426: dout  = 8'b01111111; // 1062 : 127 - 0x7f
      12'h427: dout  = 8'b01111111; // 1063 : 127 - 0x7f
      12'h428: dout  = 8'b01111100; // 1064 : 124 - 0x7c -- plane 1
      12'h429: dout  = 8'b11111110; // 1065 : 254 - 0xfe
      12'h42A: dout  = 8'b11100110; // 1066 : 230 - 0xe6
      12'h42B: dout  = 8'b00011110; // 1067 :  30 - 0x1e
      12'h42C: dout  = 8'b01111100; // 1068 : 124 - 0x7c
      12'h42D: dout  = 8'b11100000; // 1069 : 224 - 0xe0
      12'h42E: dout  = 8'b11111110; // 1070 : 254 - 0xfe
      12'h42F: dout  = 8'b00000000; // 1071 :   0 - 0x0
      12'h430: dout  = 8'b00000000; // 1072 :   0 - 0x0 -- Sprite 0x43
      12'h431: dout  = 8'b01111110; // 1073 : 126 - 0x7e
      12'h432: dout  = 8'b01111111; // 1074 : 127 - 0x7f
      12'h433: dout  = 8'b01111111; // 1075 : 127 - 0x7f
      12'h434: dout  = 8'b00011111; // 1076 :  31 - 0x1f
      12'h435: dout  = 8'b01110111; // 1077 : 119 - 0x77
      12'h436: dout  = 8'b01111111; // 1078 : 127 - 0x7f
      12'h437: dout  = 8'b01111110; // 1079 : 126 - 0x7e
      12'h438: dout  = 8'b01111100; // 1080 : 124 - 0x7c -- plane 1
      12'h439: dout  = 8'b11111100; // 1081 : 252 - 0xfc
      12'h43A: dout  = 8'b11100110; // 1082 : 230 - 0xe6
      12'h43B: dout  = 8'b00011100; // 1083 :  28 - 0x1c
      12'h43C: dout  = 8'b01100110; // 1084 : 102 - 0x66
      12'h43D: dout  = 8'b11101110; // 1085 : 238 - 0xee
      12'h43E: dout  = 8'b11111100; // 1086 : 252 - 0xfc
      12'h43F: dout  = 8'b00000000; // 1087 :   0 - 0x0
      12'h440: dout  = 8'b00000000; // 1088 :   0 - 0x0 -- Sprite 0x44
      12'h441: dout  = 8'b00001110; // 1089 :  14 - 0xe
      12'h442: dout  = 8'b00011110; // 1090 :  30 - 0x1e
      12'h443: dout  = 8'b00111110; // 1091 :  62 - 0x3e
      12'h444: dout  = 8'b01111110; // 1092 : 126 - 0x7e
      12'h445: dout  = 8'b01111111; // 1093 : 127 - 0x7f
      12'h446: dout  = 8'b01111110; // 1094 : 126 - 0x7e
      12'h447: dout  = 8'b00001100; // 1095 :  12 - 0xc
      12'h448: dout  = 8'b00001100; // 1096 :  12 - 0xc -- plane 1
      12'h449: dout  = 8'b00011100; // 1097 :  28 - 0x1c
      12'h44A: dout  = 8'b00111100; // 1098 :  60 - 0x3c
      12'h44B: dout  = 8'b01111100; // 1099 : 124 - 0x7c
      12'h44C: dout  = 8'b11101100; // 1100 : 236 - 0xec
      12'h44D: dout  = 8'b11111110; // 1101 : 254 - 0xfe
      12'h44E: dout  = 8'b00001100; // 1102 :  12 - 0xc
      12'h44F: dout  = 8'b00000000; // 1103 :   0 - 0x0
      12'h450: dout  = 8'b00000000; // 1104 :   0 - 0x0 -- Sprite 0x45
      12'h451: dout  = 8'b01111111; // 1105 : 127 - 0x7f
      12'h452: dout  = 8'b01111111; // 1106 : 127 - 0x7f
      12'h453: dout  = 8'b01111111; // 1107 : 127 - 0x7f
      12'h454: dout  = 8'b01111111; // 1108 : 127 - 0x7f
      12'h455: dout  = 8'b01110111; // 1109 : 119 - 0x77
      12'h456: dout  = 8'b01111111; // 1110 : 127 - 0x7f
      12'h457: dout  = 8'b01111110; // 1111 : 126 - 0x7e
      12'h458: dout  = 8'b11111110; // 1112 : 254 - 0xfe -- plane 1
      12'h459: dout  = 8'b11111110; // 1113 : 254 - 0xfe
      12'h45A: dout  = 8'b11100000; // 1114 : 224 - 0xe0
      12'h45B: dout  = 8'b11111110; // 1115 : 254 - 0xfe
      12'h45C: dout  = 8'b00000110; // 1116 :   6 - 0x6
      12'h45D: dout  = 8'b11101110; // 1117 : 238 - 0xee
      12'h45E: dout  = 8'b11111100; // 1118 : 252 - 0xfc
      12'h45F: dout  = 8'b00000000; // 1119 :   0 - 0x0
      12'h460: dout  = 8'b00000000; // 1120 :   0 - 0x0 -- Sprite 0x46
      12'h461: dout  = 8'b00111110; // 1121 :  62 - 0x3e
      12'h462: dout  = 8'b01111110; // 1122 : 126 - 0x7e
      12'h463: dout  = 8'b01111111; // 1123 : 127 - 0x7f
      12'h464: dout  = 8'b01111111; // 1124 : 127 - 0x7f
      12'h465: dout  = 8'b01110111; // 1125 : 119 - 0x77
      12'h466: dout  = 8'b01111111; // 1126 : 127 - 0x7f
      12'h467: dout  = 8'b00111110; // 1127 :  62 - 0x3e
      12'h468: dout  = 8'b00111100; // 1128 :  60 - 0x3c -- plane 1
      12'h469: dout  = 8'b01111100; // 1129 : 124 - 0x7c
      12'h46A: dout  = 8'b11100000; // 1130 : 224 - 0xe0
      12'h46B: dout  = 8'b11111110; // 1131 : 254 - 0xfe
      12'h46C: dout  = 8'b11100110; // 1132 : 230 - 0xe6
      12'h46D: dout  = 8'b11101110; // 1133 : 238 - 0xee
      12'h46E: dout  = 8'b00111100; // 1134 :  60 - 0x3c
      12'h46F: dout  = 8'b00000000; // 1135 :   0 - 0x0
      12'h470: dout  = 8'b00000000; // 1136 :   0 - 0x0 -- Sprite 0x47
      12'h471: dout  = 8'b01111110; // 1137 : 126 - 0x7e
      12'h472: dout  = 8'b01111110; // 1138 : 126 - 0x7e
      12'h473: dout  = 8'b00011110; // 1139 :  30 - 0x1e
      12'h474: dout  = 8'b00011100; // 1140 :  28 - 0x1c
      12'h475: dout  = 8'b00111100; // 1141 :  60 - 0x3c
      12'h476: dout  = 8'b00111000; // 1142 :  56 - 0x38
      12'h477: dout  = 8'b00111000; // 1143 :  56 - 0x38
      12'h478: dout  = 8'b11111110; // 1144 : 254 - 0xfe -- plane 1
      12'h479: dout  = 8'b11111100; // 1145 : 252 - 0xfc
      12'h47A: dout  = 8'b00001100; // 1146 :  12 - 0xc
      12'h47B: dout  = 8'b00111000; // 1147 :  56 - 0x38
      12'h47C: dout  = 8'b00111000; // 1148 :  56 - 0x38
      12'h47D: dout  = 8'b01110000; // 1149 : 112 - 0x70
      12'h47E: dout  = 8'b01110000; // 1150 : 112 - 0x70
      12'h47F: dout  = 8'b00000000; // 1151 :   0 - 0x0
      12'h480: dout  = 8'b00000000; // 1152 :   0 - 0x0 -- Sprite 0x48
      12'h481: dout  = 8'b00111110; // 1153 :  62 - 0x3e
      12'h482: dout  = 8'b01111111; // 1154 : 127 - 0x7f
      12'h483: dout  = 8'b01111111; // 1155 : 127 - 0x7f
      12'h484: dout  = 8'b01111111; // 1156 : 127 - 0x7f
      12'h485: dout  = 8'b01111111; // 1157 : 127 - 0x7f
      12'h486: dout  = 8'b01111111; // 1158 : 127 - 0x7f
      12'h487: dout  = 8'b00111110; // 1159 :  62 - 0x3e
      12'h488: dout  = 8'b00111110; // 1160 :  62 - 0x3e -- plane 1
      12'h489: dout  = 8'b01111100; // 1161 : 124 - 0x7c
      12'h48A: dout  = 8'b11100110; // 1162 : 230 - 0xe6
      12'h48B: dout  = 8'b10111100; // 1163 : 188 - 0xbc
      12'h48C: dout  = 8'b11100110; // 1164 : 230 - 0xe6
      12'h48D: dout  = 8'b11101110; // 1165 : 238 - 0xee
      12'h48E: dout  = 8'b00111100; // 1166 :  60 - 0x3c
      12'h48F: dout  = 8'b00000000; // 1167 :   0 - 0x0
      12'h490: dout  = 8'b00000000; // 1168 :   0 - 0x0 -- Sprite 0x49
      12'h491: dout  = 8'b00111110; // 1169 :  62 - 0x3e
      12'h492: dout  = 8'b01111111; // 1170 : 127 - 0x7f
      12'h493: dout  = 8'b01110111; // 1171 : 119 - 0x77
      12'h494: dout  = 8'b01111111; // 1172 : 127 - 0x7f
      12'h495: dout  = 8'b01111111; // 1173 : 127 - 0x7f
      12'h496: dout  = 8'b00111111; // 1174 :  63 - 0x3f
      12'h497: dout  = 8'b00111110; // 1175 :  62 - 0x3e
      12'h498: dout  = 8'b00111100; // 1176 :  60 - 0x3c -- plane 1
      12'h499: dout  = 8'b01111100; // 1177 : 124 - 0x7c
      12'h49A: dout  = 8'b11100110; // 1178 : 230 - 0xe6
      12'h49B: dout  = 8'b11101110; // 1179 : 238 - 0xee
      12'h49C: dout  = 8'b11111110; // 1180 : 254 - 0xfe
      12'h49D: dout  = 8'b10000110; // 1181 : 134 - 0x86
      12'h49E: dout  = 8'b01111100; // 1182 : 124 - 0x7c
      12'h49F: dout  = 8'b01000000; // 1183 :  64 - 0x40
      12'h4A0: dout  = 8'b11111111; // 1184 : 255 - 0xff -- Sprite 0x4a
      12'h4A1: dout  = 8'b10011001; // 1185 : 153 - 0x99
      12'h4A2: dout  = 8'b10011001; // 1186 : 153 - 0x99
      12'h4A3: dout  = 8'b10011001; // 1187 : 153 - 0x99
      12'h4A4: dout  = 8'b10011001; // 1188 : 153 - 0x99
      12'h4A5: dout  = 8'b10011001; // 1189 : 153 - 0x99
      12'h4A6: dout  = 8'b10011001; // 1190 : 153 - 0x99
      12'h4A7: dout  = 8'b11111111; // 1191 : 255 - 0xff
      12'h4A8: dout  = 8'b11101110; // 1192 : 238 - 0xee -- plane 1
      12'h4A9: dout  = 8'b11101110; // 1193 : 238 - 0xee
      12'h4AA: dout  = 8'b11101110; // 1194 : 238 - 0xee
      12'h4AB: dout  = 8'b11101110; // 1195 : 238 - 0xee
      12'h4AC: dout  = 8'b11101110; // 1196 : 238 - 0xee
      12'h4AD: dout  = 8'b11101110; // 1197 : 238 - 0xee
      12'h4AE: dout  = 8'b11101110; // 1198 : 238 - 0xee
      12'h4AF: dout  = 8'b10001000; // 1199 : 136 - 0x88
      12'h4B0: dout  = 8'b11110000; // 1200 : 240 - 0xf0 -- Sprite 0x4b
      12'h4B1: dout  = 8'b10010000; // 1201 : 144 - 0x90
      12'h4B2: dout  = 8'b10010000; // 1202 : 144 - 0x90
      12'h4B3: dout  = 8'b10010000; // 1203 : 144 - 0x90
      12'h4B4: dout  = 8'b10010000; // 1204 : 144 - 0x90
      12'h4B5: dout  = 8'b10010000; // 1205 : 144 - 0x90
      12'h4B6: dout  = 8'b10010000; // 1206 : 144 - 0x90
      12'h4B7: dout  = 8'b11110000; // 1207 : 240 - 0xf0
      12'h4B8: dout  = 8'b11100000; // 1208 : 224 - 0xe0 -- plane 1
      12'h4B9: dout  = 8'b11100000; // 1209 : 224 - 0xe0
      12'h4BA: dout  = 8'b11100000; // 1210 : 224 - 0xe0
      12'h4BB: dout  = 8'b11100000; // 1211 : 224 - 0xe0
      12'h4BC: dout  = 8'b11100000; // 1212 : 224 - 0xe0
      12'h4BD: dout  = 8'b11100000; // 1213 : 224 - 0xe0
      12'h4BE: dout  = 8'b11100000; // 1214 : 224 - 0xe0
      12'h4BF: dout  = 8'b10000000; // 1215 : 128 - 0x80
      12'h4C0: dout  = 8'b11111111; // 1216 : 255 - 0xff -- Sprite 0x4c
      12'h4C1: dout  = 8'b11111111; // 1217 : 255 - 0xff
      12'h4C2: dout  = 8'b11111111; // 1218 : 255 - 0xff
      12'h4C3: dout  = 8'b11111111; // 1219 : 255 - 0xff
      12'h4C4: dout  = 8'b11111111; // 1220 : 255 - 0xff
      12'h4C5: dout  = 8'b11111111; // 1221 : 255 - 0xff
      12'h4C6: dout  = 8'b11111111; // 1222 : 255 - 0xff
      12'h4C7: dout  = 8'b11111111; // 1223 : 255 - 0xff
      12'h4C8: dout  = 8'b00000000; // 1224 :   0 - 0x0 -- plane 1
      12'h4C9: dout  = 8'b01111111; // 1225 : 127 - 0x7f
      12'h4CA: dout  = 8'b01111111; // 1226 : 127 - 0x7f
      12'h4CB: dout  = 8'b01111111; // 1227 : 127 - 0x7f
      12'h4CC: dout  = 8'b01111111; // 1228 : 127 - 0x7f
      12'h4CD: dout  = 8'b01111111; // 1229 : 127 - 0x7f
      12'h4CE: dout  = 8'b01111111; // 1230 : 127 - 0x7f
      12'h4CF: dout  = 8'b01111111; // 1231 : 127 - 0x7f
      12'h4D0: dout  = 8'b11111111; // 1232 : 255 - 0xff -- Sprite 0x4d
      12'h4D1: dout  = 8'b11111111; // 1233 : 255 - 0xff
      12'h4D2: dout  = 8'b11111111; // 1234 : 255 - 0xff
      12'h4D3: dout  = 8'b11111111; // 1235 : 255 - 0xff
      12'h4D4: dout  = 8'b11111111; // 1236 : 255 - 0xff
      12'h4D5: dout  = 8'b11111111; // 1237 : 255 - 0xff
      12'h4D6: dout  = 8'b11111111; // 1238 : 255 - 0xff
      12'h4D7: dout  = 8'b11111111; // 1239 : 255 - 0xff
      12'h4D8: dout  = 8'b01111111; // 1240 : 127 - 0x7f -- plane 1
      12'h4D9: dout  = 8'b01111111; // 1241 : 127 - 0x7f
      12'h4DA: dout  = 8'b01111111; // 1242 : 127 - 0x7f
      12'h4DB: dout  = 8'b01111111; // 1243 : 127 - 0x7f
      12'h4DC: dout  = 8'b01111111; // 1244 : 127 - 0x7f
      12'h4DD: dout  = 8'b01111111; // 1245 : 127 - 0x7f
      12'h4DE: dout  = 8'b01111111; // 1246 : 127 - 0x7f
      12'h4DF: dout  = 8'b00000000; // 1247 :   0 - 0x0
      12'h4E0: dout  = 8'b11111111; // 1248 : 255 - 0xff -- Sprite 0x4e
      12'h4E1: dout  = 8'b11111111; // 1249 : 255 - 0xff
      12'h4E2: dout  = 8'b11111111; // 1250 : 255 - 0xff
      12'h4E3: dout  = 8'b11111111; // 1251 : 255 - 0xff
      12'h4E4: dout  = 8'b11111111; // 1252 : 255 - 0xff
      12'h4E5: dout  = 8'b11111111; // 1253 : 255 - 0xff
      12'h4E6: dout  = 8'b11111111; // 1254 : 255 - 0xff
      12'h4E7: dout  = 8'b11111111; // 1255 : 255 - 0xff
      12'h4E8: dout  = 8'b00000000; // 1256 :   0 - 0x0 -- plane 1
      12'h4E9: dout  = 8'b11111110; // 1257 : 254 - 0xfe
      12'h4EA: dout  = 8'b11111110; // 1258 : 254 - 0xfe
      12'h4EB: dout  = 8'b11111110; // 1259 : 254 - 0xfe
      12'h4EC: dout  = 8'b11111110; // 1260 : 254 - 0xfe
      12'h4ED: dout  = 8'b11111110; // 1261 : 254 - 0xfe
      12'h4EE: dout  = 8'b11111110; // 1262 : 254 - 0xfe
      12'h4EF: dout  = 8'b11111110; // 1263 : 254 - 0xfe
      12'h4F0: dout  = 8'b11111111; // 1264 : 255 - 0xff -- Sprite 0x4f
      12'h4F1: dout  = 8'b11111111; // 1265 : 255 - 0xff
      12'h4F2: dout  = 8'b11111111; // 1266 : 255 - 0xff
      12'h4F3: dout  = 8'b11111111; // 1267 : 255 - 0xff
      12'h4F4: dout  = 8'b11111111; // 1268 : 255 - 0xff
      12'h4F5: dout  = 8'b11111111; // 1269 : 255 - 0xff
      12'h4F6: dout  = 8'b11111111; // 1270 : 255 - 0xff
      12'h4F7: dout  = 8'b11111111; // 1271 : 255 - 0xff
      12'h4F8: dout  = 8'b11111110; // 1272 : 254 - 0xfe -- plane 1
      12'h4F9: dout  = 8'b11111110; // 1273 : 254 - 0xfe
      12'h4FA: dout  = 8'b11111110; // 1274 : 254 - 0xfe
      12'h4FB: dout  = 8'b11111110; // 1275 : 254 - 0xfe
      12'h4FC: dout  = 8'b11111110; // 1276 : 254 - 0xfe
      12'h4FD: dout  = 8'b11111110; // 1277 : 254 - 0xfe
      12'h4FE: dout  = 8'b11111110; // 1278 : 254 - 0xfe
      12'h4FF: dout  = 8'b00000000; // 1279 :   0 - 0x0
      12'h500: dout  = 8'b00010000; // 1280 :  16 - 0x10 -- Sprite 0x50
      12'h501: dout  = 8'b00101000; // 1281 :  40 - 0x28
      12'h502: dout  = 8'b11101110; // 1282 : 238 - 0xee
      12'h503: dout  = 8'b10000010; // 1283 : 130 - 0x82
      12'h504: dout  = 8'b01000100; // 1284 :  68 - 0x44
      12'h505: dout  = 8'b01000100; // 1285 :  68 - 0x44
      12'h506: dout  = 8'b10010010; // 1286 : 146 - 0x92
      12'h507: dout  = 8'b11101110; // 1287 : 238 - 0xee
      12'h508: dout  = 8'b00000000; // 1288 :   0 - 0x0 -- plane 1
      12'h509: dout  = 8'b00000000; // 1289 :   0 - 0x0
      12'h50A: dout  = 8'b00000000; // 1290 :   0 - 0x0
      12'h50B: dout  = 8'b00000000; // 1291 :   0 - 0x0
      12'h50C: dout  = 8'b00000000; // 1292 :   0 - 0x0
      12'h50D: dout  = 8'b00000000; // 1293 :   0 - 0x0
      12'h50E: dout  = 8'b00000000; // 1294 :   0 - 0x0
      12'h50F: dout  = 8'b00000000; // 1295 :   0 - 0x0
      12'h510: dout  = 8'b00010000; // 1296 :  16 - 0x10 -- Sprite 0x51
      12'h511: dout  = 8'b00101000; // 1297 :  40 - 0x28
      12'h512: dout  = 8'b11101110; // 1298 : 238 - 0xee
      12'h513: dout  = 8'b10000010; // 1299 : 130 - 0x82
      12'h514: dout  = 8'b01000100; // 1300 :  68 - 0x44
      12'h515: dout  = 8'b01000100; // 1301 :  68 - 0x44
      12'h516: dout  = 8'b10010010; // 1302 : 146 - 0x92
      12'h517: dout  = 8'b11101110; // 1303 : 238 - 0xee
      12'h518: dout  = 8'b00000000; // 1304 :   0 - 0x0 -- plane 1
      12'h519: dout  = 8'b00010000; // 1305 :  16 - 0x10
      12'h51A: dout  = 8'b00010000; // 1306 :  16 - 0x10
      12'h51B: dout  = 8'b01111100; // 1307 : 124 - 0x7c
      12'h51C: dout  = 8'b00111000; // 1308 :  56 - 0x38
      12'h51D: dout  = 8'b00111000; // 1309 :  56 - 0x38
      12'h51E: dout  = 8'b01101100; // 1310 : 108 - 0x6c
      12'h51F: dout  = 8'b00000000; // 1311 :   0 - 0x0
      12'h520: dout  = 8'b00010000; // 1312 :  16 - 0x10 -- Sprite 0x52
      12'h521: dout  = 8'b00111000; // 1313 :  56 - 0x38
      12'h522: dout  = 8'b11111110; // 1314 : 254 - 0xfe
      12'h523: dout  = 8'b11111110; // 1315 : 254 - 0xfe
      12'h524: dout  = 8'b01111100; // 1316 : 124 - 0x7c
      12'h525: dout  = 8'b01111100; // 1317 : 124 - 0x7c
      12'h526: dout  = 8'b11111110; // 1318 : 254 - 0xfe
      12'h527: dout  = 8'b11101110; // 1319 : 238 - 0xee
      12'h528: dout  = 8'b00000000; // 1320 :   0 - 0x0 -- plane 1
      12'h529: dout  = 8'b00010000; // 1321 :  16 - 0x10
      12'h52A: dout  = 8'b00010000; // 1322 :  16 - 0x10
      12'h52B: dout  = 8'b01111100; // 1323 : 124 - 0x7c
      12'h52C: dout  = 8'b00111000; // 1324 :  56 - 0x38
      12'h52D: dout  = 8'b00111000; // 1325 :  56 - 0x38
      12'h52E: dout  = 8'b01101100; // 1326 : 108 - 0x6c
      12'h52F: dout  = 8'b00000000; // 1327 :   0 - 0x0
      12'h530: dout  = 8'b11111111; // 1328 : 255 - 0xff -- Sprite 0x53
      12'h531: dout  = 8'b11111111; // 1329 : 255 - 0xff
      12'h532: dout  = 8'b11111111; // 1330 : 255 - 0xff
      12'h533: dout  = 8'b11111111; // 1331 : 255 - 0xff
      12'h534: dout  = 8'b11111111; // 1332 : 255 - 0xff
      12'h535: dout  = 8'b11111111; // 1333 : 255 - 0xff
      12'h536: dout  = 8'b11111111; // 1334 : 255 - 0xff
      12'h537: dout  = 8'b11111111; // 1335 : 255 - 0xff
      12'h538: dout  = 8'b00000000; // 1336 :   0 - 0x0 -- plane 1
      12'h539: dout  = 8'b00000000; // 1337 :   0 - 0x0
      12'h53A: dout  = 8'b00000000; // 1338 :   0 - 0x0
      12'h53B: dout  = 8'b00000000; // 1339 :   0 - 0x0
      12'h53C: dout  = 8'b00000000; // 1340 :   0 - 0x0
      12'h53D: dout  = 8'b00000000; // 1341 :   0 - 0x0
      12'h53E: dout  = 8'b00000000; // 1342 :   0 - 0x0
      12'h53F: dout  = 8'b00000000; // 1343 :   0 - 0x0
      12'h540: dout  = 8'b00000000; // 1344 :   0 - 0x0 -- Sprite 0x54
      12'h541: dout  = 8'b00000000; // 1345 :   0 - 0x0
      12'h542: dout  = 8'b00000000; // 1346 :   0 - 0x0
      12'h543: dout  = 8'b00000000; // 1347 :   0 - 0x0
      12'h544: dout  = 8'b00000000; // 1348 :   0 - 0x0
      12'h545: dout  = 8'b00000000; // 1349 :   0 - 0x0
      12'h546: dout  = 8'b00000000; // 1350 :   0 - 0x0
      12'h547: dout  = 8'b00000000; // 1351 :   0 - 0x0
      12'h548: dout  = 8'b11111111; // 1352 : 255 - 0xff -- plane 1
      12'h549: dout  = 8'b11111111; // 1353 : 255 - 0xff
      12'h54A: dout  = 8'b11111111; // 1354 : 255 - 0xff
      12'h54B: dout  = 8'b11111111; // 1355 : 255 - 0xff
      12'h54C: dout  = 8'b11111111; // 1356 : 255 - 0xff
      12'h54D: dout  = 8'b11111111; // 1357 : 255 - 0xff
      12'h54E: dout  = 8'b11111111; // 1358 : 255 - 0xff
      12'h54F: dout  = 8'b11111111; // 1359 : 255 - 0xff
      12'h550: dout  = 8'b11111111; // 1360 : 255 - 0xff -- Sprite 0x55
      12'h551: dout  = 8'b11111111; // 1361 : 255 - 0xff
      12'h552: dout  = 8'b11111111; // 1362 : 255 - 0xff
      12'h553: dout  = 8'b11111111; // 1363 : 255 - 0xff
      12'h554: dout  = 8'b11111111; // 1364 : 255 - 0xff
      12'h555: dout  = 8'b11111111; // 1365 : 255 - 0xff
      12'h556: dout  = 8'b11111111; // 1366 : 255 - 0xff
      12'h557: dout  = 8'b11111111; // 1367 : 255 - 0xff
      12'h558: dout  = 8'b11111111; // 1368 : 255 - 0xff -- plane 1
      12'h559: dout  = 8'b11111111; // 1369 : 255 - 0xff
      12'h55A: dout  = 8'b11111111; // 1370 : 255 - 0xff
      12'h55B: dout  = 8'b11111111; // 1371 : 255 - 0xff
      12'h55C: dout  = 8'b11111111; // 1372 : 255 - 0xff
      12'h55D: dout  = 8'b11111111; // 1373 : 255 - 0xff
      12'h55E: dout  = 8'b11111111; // 1374 : 255 - 0xff
      12'h55F: dout  = 8'b11111111; // 1375 : 255 - 0xff
      12'h560: dout  = 8'b00101010; // 1376 :  42 - 0x2a -- Sprite 0x56
      12'h561: dout  = 8'b01000101; // 1377 :  69 - 0x45
      12'h562: dout  = 8'b00001000; // 1378 :   8 - 0x8
      12'h563: dout  = 8'b00010101; // 1379 :  21 - 0x15
      12'h564: dout  = 8'b00100000; // 1380 :  32 - 0x20
      12'h565: dout  = 8'b01000101; // 1381 :  69 - 0x45
      12'h566: dout  = 8'b10101000; // 1382 : 168 - 0xa8
      12'h567: dout  = 8'b00000000; // 1383 :   0 - 0x0
      12'h568: dout  = 8'b00000010; // 1384 :   2 - 0x2 -- plane 1
      12'h569: dout  = 8'b00000101; // 1385 :   5 - 0x5
      12'h56A: dout  = 8'b10101010; // 1386 : 170 - 0xaa
      12'h56B: dout  = 8'b01010001; // 1387 :  81 - 0x51
      12'h56C: dout  = 8'b10101010; // 1388 : 170 - 0xaa
      12'h56D: dout  = 8'b01010001; // 1389 :  81 - 0x51
      12'h56E: dout  = 8'b10100010; // 1390 : 162 - 0xa2
      12'h56F: dout  = 8'b00000100; // 1391 :   4 - 0x4
      12'h570: dout  = 8'b00001000; // 1392 :   8 - 0x8 -- Sprite 0x57
      12'h571: dout  = 8'b01010101; // 1393 :  85 - 0x55
      12'h572: dout  = 8'b10100000; // 1394 : 160 - 0xa0
      12'h573: dout  = 8'b00010000; // 1395 :  16 - 0x10
      12'h574: dout  = 8'b10000000; // 1396 : 128 - 0x80
      12'h575: dout  = 8'b00010100; // 1397 :  20 - 0x14
      12'h576: dout  = 8'b00100010; // 1398 :  34 - 0x22
      12'h577: dout  = 8'b00000000; // 1399 :   0 - 0x0
      12'h578: dout  = 8'b00001000; // 1400 :   8 - 0x8 -- plane 1
      12'h579: dout  = 8'b01010101; // 1401 :  85 - 0x55
      12'h57A: dout  = 8'b00101010; // 1402 :  42 - 0x2a
      12'h57B: dout  = 8'b01010101; // 1403 :  85 - 0x55
      12'h57C: dout  = 8'b00101010; // 1404 :  42 - 0x2a
      12'h57D: dout  = 8'b01000101; // 1405 :  69 - 0x45
      12'h57E: dout  = 8'b00001010; // 1406 :  10 - 0xa
      12'h57F: dout  = 8'b00010000; // 1407 :  16 - 0x10
      12'h580: dout  = 8'b11111111; // 1408 : 255 - 0xff -- Sprite 0x58
      12'h581: dout  = 8'b11010101; // 1409 : 213 - 0xd5
      12'h582: dout  = 8'b10100000; // 1410 : 160 - 0xa0
      12'h583: dout  = 8'b11010000; // 1411 : 208 - 0xd0
      12'h584: dout  = 8'b10001111; // 1412 : 143 - 0x8f
      12'h585: dout  = 8'b11001000; // 1413 : 200 - 0xc8
      12'h586: dout  = 8'b10001000; // 1414 : 136 - 0x88
      12'h587: dout  = 8'b11001000; // 1415 : 200 - 0xc8
      12'h588: dout  = 8'b00000000; // 1416 :   0 - 0x0 -- plane 1
      12'h589: dout  = 8'b00111111; // 1417 :  63 - 0x3f
      12'h58A: dout  = 8'b01011111; // 1418 :  95 - 0x5f
      12'h58B: dout  = 8'b01101111; // 1419 : 111 - 0x6f
      12'h58C: dout  = 8'b01110000; // 1420 : 112 - 0x70
      12'h58D: dout  = 8'b01110111; // 1421 : 119 - 0x77
      12'h58E: dout  = 8'b01110111; // 1422 : 119 - 0x77
      12'h58F: dout  = 8'b01110111; // 1423 : 119 - 0x77
      12'h590: dout  = 8'b10001000; // 1424 : 136 - 0x88 -- Sprite 0x59
      12'h591: dout  = 8'b11001000; // 1425 : 200 - 0xc8
      12'h592: dout  = 8'b10001000; // 1426 : 136 - 0x88
      12'h593: dout  = 8'b11001111; // 1427 : 207 - 0xcf
      12'h594: dout  = 8'b10010000; // 1428 : 144 - 0x90
      12'h595: dout  = 8'b11100000; // 1429 : 224 - 0xe0
      12'h596: dout  = 8'b11101010; // 1430 : 234 - 0xea
      12'h597: dout  = 8'b11111111; // 1431 : 255 - 0xff
      12'h598: dout  = 8'b01110111; // 1432 : 119 - 0x77 -- plane 1
      12'h599: dout  = 8'b01110111; // 1433 : 119 - 0x77
      12'h59A: dout  = 8'b01110111; // 1434 : 119 - 0x77
      12'h59B: dout  = 8'b01110000; // 1435 : 112 - 0x70
      12'h59C: dout  = 8'b01101111; // 1436 : 111 - 0x6f
      12'h59D: dout  = 8'b01011111; // 1437 :  95 - 0x5f
      12'h59E: dout  = 8'b00010101; // 1438 :  21 - 0x15
      12'h59F: dout  = 8'b00000000; // 1439 :   0 - 0x0
      12'h5A0: dout  = 8'b11111111; // 1440 : 255 - 0xff -- Sprite 0x5a
      12'h5A1: dout  = 8'b01011011; // 1441 :  91 - 0x5b
      12'h5A2: dout  = 8'b00000111; // 1442 :   7 - 0x7
      12'h5A3: dout  = 8'b00001001; // 1443 :   9 - 0x9
      12'h5A4: dout  = 8'b11110011; // 1444 : 243 - 0xf3
      12'h5A5: dout  = 8'b00010001; // 1445 :  17 - 0x11
      12'h5A6: dout  = 8'b00010011; // 1446 :  19 - 0x13
      12'h5A7: dout  = 8'b00010001; // 1447 :  17 - 0x11
      12'h5A8: dout  = 8'b00000000; // 1448 :   0 - 0x0 -- plane 1
      12'h5A9: dout  = 8'b11111100; // 1449 : 252 - 0xfc
      12'h5AA: dout  = 8'b11111000; // 1450 : 248 - 0xf8
      12'h5AB: dout  = 8'b11110110; // 1451 : 246 - 0xf6
      12'h5AC: dout  = 8'b00001100; // 1452 :  12 - 0xc
      12'h5AD: dout  = 8'b11101110; // 1453 : 238 - 0xee
      12'h5AE: dout  = 8'b11101100; // 1454 : 236 - 0xec
      12'h5AF: dout  = 8'b11101110; // 1455 : 238 - 0xee
      12'h5B0: dout  = 8'b00010011; // 1456 :  19 - 0x13 -- Sprite 0x5b
      12'h5B1: dout  = 8'b00010001; // 1457 :  17 - 0x11
      12'h5B2: dout  = 8'b00010011; // 1458 :  19 - 0x13
      12'h5B3: dout  = 8'b11110001; // 1459 : 241 - 0xf1
      12'h5B4: dout  = 8'b00001011; // 1460 :  11 - 0xb
      12'h5B5: dout  = 8'b00000101; // 1461 :   5 - 0x5
      12'h5B6: dout  = 8'b10101011; // 1462 : 171 - 0xab
      12'h5B7: dout  = 8'b11111111; // 1463 : 255 - 0xff
      12'h5B8: dout  = 8'b11101100; // 1464 : 236 - 0xec -- plane 1
      12'h5B9: dout  = 8'b11101110; // 1465 : 238 - 0xee
      12'h5BA: dout  = 8'b11101100; // 1466 : 236 - 0xec
      12'h5BB: dout  = 8'b00001110; // 1467 :  14 - 0xe
      12'h5BC: dout  = 8'b11110100; // 1468 : 244 - 0xf4
      12'h5BD: dout  = 8'b11111010; // 1469 : 250 - 0xfa
      12'h5BE: dout  = 8'b01010100; // 1470 :  84 - 0x54
      12'h5BF: dout  = 8'b00000000; // 1471 :   0 - 0x0
      12'h5C0: dout  = 8'b00011100; // 1472 :  28 - 0x1c -- Sprite 0x5c
      12'h5C1: dout  = 8'b00100010; // 1473 :  34 - 0x22
      12'h5C2: dout  = 8'b01000001; // 1474 :  65 - 0x41
      12'h5C3: dout  = 8'b01000001; // 1475 :  65 - 0x41
      12'h5C4: dout  = 8'b01000001; // 1476 :  65 - 0x41
      12'h5C5: dout  = 8'b00100010; // 1477 :  34 - 0x22
      12'h5C6: dout  = 8'b00100010; // 1478 :  34 - 0x22
      12'h5C7: dout  = 8'b00011100; // 1479 :  28 - 0x1c
      12'h5C8: dout  = 8'b00000000; // 1480 :   0 - 0x0 -- plane 1
      12'h5C9: dout  = 8'b00011100; // 1481 :  28 - 0x1c
      12'h5CA: dout  = 8'b00111110; // 1482 :  62 - 0x3e
      12'h5CB: dout  = 8'b00111110; // 1483 :  62 - 0x3e
      12'h5CC: dout  = 8'b00111110; // 1484 :  62 - 0x3e
      12'h5CD: dout  = 8'b00011100; // 1485 :  28 - 0x1c
      12'h5CE: dout  = 8'b00011100; // 1486 :  28 - 0x1c
      12'h5CF: dout  = 8'b00000000; // 1487 :   0 - 0x0
      12'h5D0: dout  = 8'b00001000; // 1488 :   8 - 0x8 -- Sprite 0x5d
      12'h5D1: dout  = 8'b00010000; // 1489 :  16 - 0x10
      12'h5D2: dout  = 8'b00010000; // 1490 :  16 - 0x10
      12'h5D3: dout  = 8'b00001000; // 1491 :   8 - 0x8
      12'h5D4: dout  = 8'b00000100; // 1492 :   4 - 0x4
      12'h5D5: dout  = 8'b00000100; // 1493 :   4 - 0x4
      12'h5D6: dout  = 8'b00001000; // 1494 :   8 - 0x8
      12'h5D7: dout  = 8'b00010000; // 1495 :  16 - 0x10
      12'h5D8: dout  = 8'b00000000; // 1496 :   0 - 0x0 -- plane 1
      12'h5D9: dout  = 8'b00000000; // 1497 :   0 - 0x0
      12'h5DA: dout  = 8'b00000000; // 1498 :   0 - 0x0
      12'h5DB: dout  = 8'b00000000; // 1499 :   0 - 0x0
      12'h5DC: dout  = 8'b00000000; // 1500 :   0 - 0x0
      12'h5DD: dout  = 8'b00000000; // 1501 :   0 - 0x0
      12'h5DE: dout  = 8'b00000000; // 1502 :   0 - 0x0
      12'h5DF: dout  = 8'b00000000; // 1503 :   0 - 0x0
      12'h5E0: dout  = 8'b00110110; // 1504 :  54 - 0x36 -- Sprite 0x5e
      12'h5E1: dout  = 8'b01101011; // 1505 : 107 - 0x6b
      12'h5E2: dout  = 8'b01001001; // 1506 :  73 - 0x49
      12'h5E3: dout  = 8'b01000001; // 1507 :  65 - 0x41
      12'h5E4: dout  = 8'b01000001; // 1508 :  65 - 0x41
      12'h5E5: dout  = 8'b00100010; // 1509 :  34 - 0x22
      12'h5E6: dout  = 8'b00010100; // 1510 :  20 - 0x14
      12'h5E7: dout  = 8'b00001000; // 1511 :   8 - 0x8
      12'h5E8: dout  = 8'b00000000; // 1512 :   0 - 0x0 -- plane 1
      12'h5E9: dout  = 8'b00010100; // 1513 :  20 - 0x14
      12'h5EA: dout  = 8'b00110110; // 1514 :  54 - 0x36
      12'h5EB: dout  = 8'b00111110; // 1515 :  62 - 0x3e
      12'h5EC: dout  = 8'b00111110; // 1516 :  62 - 0x3e
      12'h5ED: dout  = 8'b00011100; // 1517 :  28 - 0x1c
      12'h5EE: dout  = 8'b00001000; // 1518 :   8 - 0x8
      12'h5EF: dout  = 8'b00000000; // 1519 :   0 - 0x0
      12'h5F0: dout  = 8'b00111110; // 1520 :  62 - 0x3e -- Sprite 0x5f
      12'h5F1: dout  = 8'b01101011; // 1521 : 107 - 0x6b
      12'h5F2: dout  = 8'b00100010; // 1522 :  34 - 0x22
      12'h5F3: dout  = 8'b01100011; // 1523 :  99 - 0x63
      12'h5F4: dout  = 8'b00100010; // 1524 :  34 - 0x22
      12'h5F5: dout  = 8'b01100011; // 1525 :  99 - 0x63
      12'h5F6: dout  = 8'b00100010; // 1526 :  34 - 0x22
      12'h5F7: dout  = 8'b01111111; // 1527 : 127 - 0x7f
      12'h5F8: dout  = 8'b00000000; // 1528 :   0 - 0x0 -- plane 1
      12'h5F9: dout  = 8'b00010100; // 1529 :  20 - 0x14
      12'h5FA: dout  = 8'b00011100; // 1530 :  28 - 0x1c
      12'h5FB: dout  = 8'b00011100; // 1531 :  28 - 0x1c
      12'h5FC: dout  = 8'b00011100; // 1532 :  28 - 0x1c
      12'h5FD: dout  = 8'b00011100; // 1533 :  28 - 0x1c
      12'h5FE: dout  = 8'b00011100; // 1534 :  28 - 0x1c
      12'h5FF: dout  = 8'b00000000; // 1535 :   0 - 0x0
      12'h600: dout  = 8'b11111111; // 1536 : 255 - 0xff -- Sprite 0x60
      12'h601: dout  = 8'b11111111; // 1537 : 255 - 0xff
      12'h602: dout  = 8'b11111111; // 1538 : 255 - 0xff
      12'h603: dout  = 8'b11111111; // 1539 : 255 - 0xff
      12'h604: dout  = 8'b11010101; // 1540 : 213 - 0xd5
      12'h605: dout  = 8'b10101010; // 1541 : 170 - 0xaa
      12'h606: dout  = 8'b11010101; // 1542 : 213 - 0xd5
      12'h607: dout  = 8'b11111111; // 1543 : 255 - 0xff
      12'h608: dout  = 8'b00000000; // 1544 :   0 - 0x0 -- plane 1
      12'h609: dout  = 8'b01111111; // 1545 : 127 - 0x7f
      12'h60A: dout  = 8'b01111111; // 1546 : 127 - 0x7f
      12'h60B: dout  = 8'b01111111; // 1547 : 127 - 0x7f
      12'h60C: dout  = 8'b01111111; // 1548 : 127 - 0x7f
      12'h60D: dout  = 8'b01111111; // 1549 : 127 - 0x7f
      12'h60E: dout  = 8'b00101010; // 1550 :  42 - 0x2a
      12'h60F: dout  = 8'b00000000; // 1551 :   0 - 0x0
      12'h610: dout  = 8'b11111111; // 1552 : 255 - 0xff -- Sprite 0x61
      12'h611: dout  = 8'b11111111; // 1553 : 255 - 0xff
      12'h612: dout  = 8'b11111111; // 1554 : 255 - 0xff
      12'h613: dout  = 8'b11111111; // 1555 : 255 - 0xff
      12'h614: dout  = 8'b01010101; // 1556 :  85 - 0x55
      12'h615: dout  = 8'b10101010; // 1557 : 170 - 0xaa
      12'h616: dout  = 8'b01010101; // 1558 :  85 - 0x55
      12'h617: dout  = 8'b11111111; // 1559 : 255 - 0xff
      12'h618: dout  = 8'b00000000; // 1560 :   0 - 0x0 -- plane 1
      12'h619: dout  = 8'b11111111; // 1561 : 255 - 0xff
      12'h61A: dout  = 8'b11111111; // 1562 : 255 - 0xff
      12'h61B: dout  = 8'b11111111; // 1563 : 255 - 0xff
      12'h61C: dout  = 8'b11111111; // 1564 : 255 - 0xff
      12'h61D: dout  = 8'b11111111; // 1565 : 255 - 0xff
      12'h61E: dout  = 8'b10101010; // 1566 : 170 - 0xaa
      12'h61F: dout  = 8'b00000000; // 1567 :   0 - 0x0
      12'h620: dout  = 8'b11111111; // 1568 : 255 - 0xff -- Sprite 0x62
      12'h621: dout  = 8'b11111111; // 1569 : 255 - 0xff
      12'h622: dout  = 8'b11111111; // 1570 : 255 - 0xff
      12'h623: dout  = 8'b11111111; // 1571 : 255 - 0xff
      12'h624: dout  = 8'b01010101; // 1572 :  85 - 0x55
      12'h625: dout  = 8'b10101011; // 1573 : 171 - 0xab
      12'h626: dout  = 8'b01010101; // 1574 :  85 - 0x55
      12'h627: dout  = 8'b11111111; // 1575 : 255 - 0xff
      12'h628: dout  = 8'b00000000; // 1576 :   0 - 0x0 -- plane 1
      12'h629: dout  = 8'b11111110; // 1577 : 254 - 0xfe
      12'h62A: dout  = 8'b11111110; // 1578 : 254 - 0xfe
      12'h62B: dout  = 8'b11111110; // 1579 : 254 - 0xfe
      12'h62C: dout  = 8'b11111110; // 1580 : 254 - 0xfe
      12'h62D: dout  = 8'b11111110; // 1581 : 254 - 0xfe
      12'h62E: dout  = 8'b10101010; // 1582 : 170 - 0xaa
      12'h62F: dout  = 8'b00000000; // 1583 :   0 - 0x0
      12'h630: dout  = 8'b00000000; // 1584 :   0 - 0x0 -- Sprite 0x63
      12'h631: dout  = 8'b00000000; // 1585 :   0 - 0x0
      12'h632: dout  = 8'b00000000; // 1586 :   0 - 0x0
      12'h633: dout  = 8'b00000000; // 1587 :   0 - 0x0
      12'h634: dout  = 8'b00000000; // 1588 :   0 - 0x0
      12'h635: dout  = 8'b00000000; // 1589 :   0 - 0x0
      12'h636: dout  = 8'b00000000; // 1590 :   0 - 0x0
      12'h637: dout  = 8'b00000000; // 1591 :   0 - 0x0
      12'h638: dout  = 8'b00000000; // 1592 :   0 - 0x0 -- plane 1
      12'h639: dout  = 8'b00000000; // 1593 :   0 - 0x0
      12'h63A: dout  = 8'b00000000; // 1594 :   0 - 0x0
      12'h63B: dout  = 8'b00000000; // 1595 :   0 - 0x0
      12'h63C: dout  = 8'b00000000; // 1596 :   0 - 0x0
      12'h63D: dout  = 8'b00000000; // 1597 :   0 - 0x0
      12'h63E: dout  = 8'b00000000; // 1598 :   0 - 0x0
      12'h63F: dout  = 8'b00000000; // 1599 :   0 - 0x0
      12'h640: dout  = 8'b00000001; // 1600 :   1 - 0x1 -- Sprite 0x64
      12'h641: dout  = 8'b00000001; // 1601 :   1 - 0x1
      12'h642: dout  = 8'b00000011; // 1602 :   3 - 0x3
      12'h643: dout  = 8'b00000011; // 1603 :   3 - 0x3
      12'h644: dout  = 8'b00000110; // 1604 :   6 - 0x6
      12'h645: dout  = 8'b00000110; // 1605 :   6 - 0x6
      12'h646: dout  = 8'b00001100; // 1606 :  12 - 0xc
      12'h647: dout  = 8'b00001100; // 1607 :  12 - 0xc
      12'h648: dout  = 8'b00000000; // 1608 :   0 - 0x0 -- plane 1
      12'h649: dout  = 8'b00000000; // 1609 :   0 - 0x0
      12'h64A: dout  = 8'b00000001; // 1610 :   1 - 0x1
      12'h64B: dout  = 8'b00000001; // 1611 :   1 - 0x1
      12'h64C: dout  = 8'b00000011; // 1612 :   3 - 0x3
      12'h64D: dout  = 8'b00000011; // 1613 :   3 - 0x3
      12'h64E: dout  = 8'b00000111; // 1614 :   7 - 0x7
      12'h64F: dout  = 8'b00000111; // 1615 :   7 - 0x7
      12'h650: dout  = 8'b00011000; // 1616 :  24 - 0x18 -- Sprite 0x65
      12'h651: dout  = 8'b00011000; // 1617 :  24 - 0x18
      12'h652: dout  = 8'b00110000; // 1618 :  48 - 0x30
      12'h653: dout  = 8'b00110000; // 1619 :  48 - 0x30
      12'h654: dout  = 8'b01100000; // 1620 :  96 - 0x60
      12'h655: dout  = 8'b01100000; // 1621 :  96 - 0x60
      12'h656: dout  = 8'b11101010; // 1622 : 234 - 0xea
      12'h657: dout  = 8'b11111111; // 1623 : 255 - 0xff
      12'h658: dout  = 8'b00001111; // 1624 :  15 - 0xf -- plane 1
      12'h659: dout  = 8'b00001111; // 1625 :  15 - 0xf
      12'h65A: dout  = 8'b00011111; // 1626 :  31 - 0x1f
      12'h65B: dout  = 8'b00011111; // 1627 :  31 - 0x1f
      12'h65C: dout  = 8'b00111111; // 1628 :  63 - 0x3f
      12'h65D: dout  = 8'b00111111; // 1629 :  63 - 0x3f
      12'h65E: dout  = 8'b01010101; // 1630 :  85 - 0x55
      12'h65F: dout  = 8'b00000000; // 1631 :   0 - 0x0
      12'h660: dout  = 8'b10000000; // 1632 : 128 - 0x80 -- Sprite 0x66
      12'h661: dout  = 8'b10000000; // 1633 : 128 - 0x80
      12'h662: dout  = 8'b11000000; // 1634 : 192 - 0xc0
      12'h663: dout  = 8'b01000000; // 1635 :  64 - 0x40
      12'h664: dout  = 8'b10100000; // 1636 : 160 - 0xa0
      12'h665: dout  = 8'b01100000; // 1637 :  96 - 0x60
      12'h666: dout  = 8'b00110000; // 1638 :  48 - 0x30
      12'h667: dout  = 8'b00010000; // 1639 :  16 - 0x10
      12'h668: dout  = 8'b00000000; // 1640 :   0 - 0x0 -- plane 1
      12'h669: dout  = 8'b00000000; // 1641 :   0 - 0x0
      12'h66A: dout  = 8'b00000000; // 1642 :   0 - 0x0
      12'h66B: dout  = 8'b10000000; // 1643 : 128 - 0x80
      12'h66C: dout  = 8'b01000000; // 1644 :  64 - 0x40
      12'h66D: dout  = 8'b10000000; // 1645 : 128 - 0x80
      12'h66E: dout  = 8'b11000000; // 1646 : 192 - 0xc0
      12'h66F: dout  = 8'b11100000; // 1647 : 224 - 0xe0
      12'h670: dout  = 8'b00101000; // 1648 :  40 - 0x28 -- Sprite 0x67
      12'h671: dout  = 8'b00011000; // 1649 :  24 - 0x18
      12'h672: dout  = 8'b00001100; // 1650 :  12 - 0xc
      12'h673: dout  = 8'b00010100; // 1651 :  20 - 0x14
      12'h674: dout  = 8'b00001010; // 1652 :  10 - 0xa
      12'h675: dout  = 8'b00000110; // 1653 :   6 - 0x6
      12'h676: dout  = 8'b10101011; // 1654 : 171 - 0xab
      12'h677: dout  = 8'b11111111; // 1655 : 255 - 0xff
      12'h678: dout  = 8'b11010000; // 1656 : 208 - 0xd0 -- plane 1
      12'h679: dout  = 8'b11100000; // 1657 : 224 - 0xe0
      12'h67A: dout  = 8'b11110000; // 1658 : 240 - 0xf0
      12'h67B: dout  = 8'b11101000; // 1659 : 232 - 0xe8
      12'h67C: dout  = 8'b11110100; // 1660 : 244 - 0xf4
      12'h67D: dout  = 8'b11111000; // 1661 : 248 - 0xf8
      12'h67E: dout  = 8'b01010100; // 1662 :  84 - 0x54
      12'h67F: dout  = 8'b00000000; // 1663 :   0 - 0x0
      12'h680: dout  = 8'b00000000; // 1664 :   0 - 0x0 -- Sprite 0x68
      12'h681: dout  = 8'b00000000; // 1665 :   0 - 0x0
      12'h682: dout  = 8'b00000000; // 1666 :   0 - 0x0
      12'h683: dout  = 8'b00000000; // 1667 :   0 - 0x0
      12'h684: dout  = 8'b00000000; // 1668 :   0 - 0x0
      12'h685: dout  = 8'b00000000; // 1669 :   0 - 0x0
      12'h686: dout  = 8'b00000000; // 1670 :   0 - 0x0
      12'h687: dout  = 8'b00000000; // 1671 :   0 - 0x0
      12'h688: dout  = 8'b00000000; // 1672 :   0 - 0x0 -- plane 1
      12'h689: dout  = 8'b00000000; // 1673 :   0 - 0x0
      12'h68A: dout  = 8'b00000000; // 1674 :   0 - 0x0
      12'h68B: dout  = 8'b00000000; // 1675 :   0 - 0x0
      12'h68C: dout  = 8'b00000000; // 1676 :   0 - 0x0
      12'h68D: dout  = 8'b00000000; // 1677 :   0 - 0x0
      12'h68E: dout  = 8'b00000000; // 1678 :   0 - 0x0
      12'h68F: dout  = 8'b00000000; // 1679 :   0 - 0x0
      12'h690: dout  = 8'b00000000; // 1680 :   0 - 0x0 -- Sprite 0x69
      12'h691: dout  = 8'b00000000; // 1681 :   0 - 0x0
      12'h692: dout  = 8'b00000000; // 1682 :   0 - 0x0
      12'h693: dout  = 8'b00000000; // 1683 :   0 - 0x0
      12'h694: dout  = 8'b00000000; // 1684 :   0 - 0x0
      12'h695: dout  = 8'b00000000; // 1685 :   0 - 0x0
      12'h696: dout  = 8'b00000000; // 1686 :   0 - 0x0
      12'h697: dout  = 8'b00000000; // 1687 :   0 - 0x0
      12'h698: dout  = 8'b00000000; // 1688 :   0 - 0x0 -- plane 1
      12'h699: dout  = 8'b00000000; // 1689 :   0 - 0x0
      12'h69A: dout  = 8'b00000000; // 1690 :   0 - 0x0
      12'h69B: dout  = 8'b00000000; // 1691 :   0 - 0x0
      12'h69C: dout  = 8'b00000000; // 1692 :   0 - 0x0
      12'h69D: dout  = 8'b00000000; // 1693 :   0 - 0x0
      12'h69E: dout  = 8'b00000000; // 1694 :   0 - 0x0
      12'h69F: dout  = 8'b00000000; // 1695 :   0 - 0x0
      12'h6A0: dout  = 8'b00000000; // 1696 :   0 - 0x0 -- Sprite 0x6a
      12'h6A1: dout  = 8'b00000000; // 1697 :   0 - 0x0
      12'h6A2: dout  = 8'b00000000; // 1698 :   0 - 0x0
      12'h6A3: dout  = 8'b00000000; // 1699 :   0 - 0x0
      12'h6A4: dout  = 8'b00000000; // 1700 :   0 - 0x0
      12'h6A5: dout  = 8'b00000000; // 1701 :   0 - 0x0
      12'h6A6: dout  = 8'b00000000; // 1702 :   0 - 0x0
      12'h6A7: dout  = 8'b00000000; // 1703 :   0 - 0x0
      12'h6A8: dout  = 8'b00000000; // 1704 :   0 - 0x0 -- plane 1
      12'h6A9: dout  = 8'b00000000; // 1705 :   0 - 0x0
      12'h6AA: dout  = 8'b00000000; // 1706 :   0 - 0x0
      12'h6AB: dout  = 8'b00000000; // 1707 :   0 - 0x0
      12'h6AC: dout  = 8'b00000000; // 1708 :   0 - 0x0
      12'h6AD: dout  = 8'b00000000; // 1709 :   0 - 0x0
      12'h6AE: dout  = 8'b00000000; // 1710 :   0 - 0x0
      12'h6AF: dout  = 8'b00000000; // 1711 :   0 - 0x0
      12'h6B0: dout  = 8'b00000000; // 1712 :   0 - 0x0 -- Sprite 0x6b
      12'h6B1: dout  = 8'b00000000; // 1713 :   0 - 0x0
      12'h6B2: dout  = 8'b00000000; // 1714 :   0 - 0x0
      12'h6B3: dout  = 8'b00000000; // 1715 :   0 - 0x0
      12'h6B4: dout  = 8'b00000000; // 1716 :   0 - 0x0
      12'h6B5: dout  = 8'b00000000; // 1717 :   0 - 0x0
      12'h6B6: dout  = 8'b00000000; // 1718 :   0 - 0x0
      12'h6B7: dout  = 8'b00000000; // 1719 :   0 - 0x0
      12'h6B8: dout  = 8'b00000000; // 1720 :   0 - 0x0 -- plane 1
      12'h6B9: dout  = 8'b00000000; // 1721 :   0 - 0x0
      12'h6BA: dout  = 8'b00000000; // 1722 :   0 - 0x0
      12'h6BB: dout  = 8'b00000000; // 1723 :   0 - 0x0
      12'h6BC: dout  = 8'b00000000; // 1724 :   0 - 0x0
      12'h6BD: dout  = 8'b00000000; // 1725 :   0 - 0x0
      12'h6BE: dout  = 8'b00000000; // 1726 :   0 - 0x0
      12'h6BF: dout  = 8'b00000000; // 1727 :   0 - 0x0
      12'h6C0: dout  = 8'b00000000; // 1728 :   0 - 0x0 -- Sprite 0x6c
      12'h6C1: dout  = 8'b00000000; // 1729 :   0 - 0x0
      12'h6C2: dout  = 8'b00000000; // 1730 :   0 - 0x0
      12'h6C3: dout  = 8'b00000000; // 1731 :   0 - 0x0
      12'h6C4: dout  = 8'b00000000; // 1732 :   0 - 0x0
      12'h6C5: dout  = 8'b00000000; // 1733 :   0 - 0x0
      12'h6C6: dout  = 8'b00000000; // 1734 :   0 - 0x0
      12'h6C7: dout  = 8'b00000000; // 1735 :   0 - 0x0
      12'h6C8: dout  = 8'b00000000; // 1736 :   0 - 0x0 -- plane 1
      12'h6C9: dout  = 8'b00000000; // 1737 :   0 - 0x0
      12'h6CA: dout  = 8'b00000000; // 1738 :   0 - 0x0
      12'h6CB: dout  = 8'b00000000; // 1739 :   0 - 0x0
      12'h6CC: dout  = 8'b00000000; // 1740 :   0 - 0x0
      12'h6CD: dout  = 8'b00000000; // 1741 :   0 - 0x0
      12'h6CE: dout  = 8'b00000000; // 1742 :   0 - 0x0
      12'h6CF: dout  = 8'b00000000; // 1743 :   0 - 0x0
      12'h6D0: dout  = 8'b00000000; // 1744 :   0 - 0x0 -- Sprite 0x6d
      12'h6D1: dout  = 8'b00000000; // 1745 :   0 - 0x0
      12'h6D2: dout  = 8'b00000000; // 1746 :   0 - 0x0
      12'h6D3: dout  = 8'b00000000; // 1747 :   0 - 0x0
      12'h6D4: dout  = 8'b00000000; // 1748 :   0 - 0x0
      12'h6D5: dout  = 8'b00000000; // 1749 :   0 - 0x0
      12'h6D6: dout  = 8'b00000000; // 1750 :   0 - 0x0
      12'h6D7: dout  = 8'b00000000; // 1751 :   0 - 0x0
      12'h6D8: dout  = 8'b00000000; // 1752 :   0 - 0x0 -- plane 1
      12'h6D9: dout  = 8'b00000000; // 1753 :   0 - 0x0
      12'h6DA: dout  = 8'b00000000; // 1754 :   0 - 0x0
      12'h6DB: dout  = 8'b00000000; // 1755 :   0 - 0x0
      12'h6DC: dout  = 8'b00000000; // 1756 :   0 - 0x0
      12'h6DD: dout  = 8'b00000000; // 1757 :   0 - 0x0
      12'h6DE: dout  = 8'b00000000; // 1758 :   0 - 0x0
      12'h6DF: dout  = 8'b00000000; // 1759 :   0 - 0x0
      12'h6E0: dout  = 8'b00000000; // 1760 :   0 - 0x0 -- Sprite 0x6e
      12'h6E1: dout  = 8'b00000000; // 1761 :   0 - 0x0
      12'h6E2: dout  = 8'b00000000; // 1762 :   0 - 0x0
      12'h6E3: dout  = 8'b00000000; // 1763 :   0 - 0x0
      12'h6E4: dout  = 8'b00000000; // 1764 :   0 - 0x0
      12'h6E5: dout  = 8'b00000000; // 1765 :   0 - 0x0
      12'h6E6: dout  = 8'b00000000; // 1766 :   0 - 0x0
      12'h6E7: dout  = 8'b00000000; // 1767 :   0 - 0x0
      12'h6E8: dout  = 8'b00000000; // 1768 :   0 - 0x0 -- plane 1
      12'h6E9: dout  = 8'b00000000; // 1769 :   0 - 0x0
      12'h6EA: dout  = 8'b00000000; // 1770 :   0 - 0x0
      12'h6EB: dout  = 8'b00000000; // 1771 :   0 - 0x0
      12'h6EC: dout  = 8'b00000000; // 1772 :   0 - 0x0
      12'h6ED: dout  = 8'b00000000; // 1773 :   0 - 0x0
      12'h6EE: dout  = 8'b00000000; // 1774 :   0 - 0x0
      12'h6EF: dout  = 8'b00000000; // 1775 :   0 - 0x0
      12'h6F0: dout  = 8'b00000000; // 1776 :   0 - 0x0 -- Sprite 0x6f
      12'h6F1: dout  = 8'b00000000; // 1777 :   0 - 0x0
      12'h6F2: dout  = 8'b00000000; // 1778 :   0 - 0x0
      12'h6F3: dout  = 8'b00000000; // 1779 :   0 - 0x0
      12'h6F4: dout  = 8'b00000000; // 1780 :   0 - 0x0
      12'h6F5: dout  = 8'b00000000; // 1781 :   0 - 0x0
      12'h6F6: dout  = 8'b00000000; // 1782 :   0 - 0x0
      12'h6F7: dout  = 8'b00000000; // 1783 :   0 - 0x0
      12'h6F8: dout  = 8'b00000000; // 1784 :   0 - 0x0 -- plane 1
      12'h6F9: dout  = 8'b00000000; // 1785 :   0 - 0x0
      12'h6FA: dout  = 8'b00000000; // 1786 :   0 - 0x0
      12'h6FB: dout  = 8'b00000000; // 1787 :   0 - 0x0
      12'h6FC: dout  = 8'b00000000; // 1788 :   0 - 0x0
      12'h6FD: dout  = 8'b00000000; // 1789 :   0 - 0x0
      12'h6FE: dout  = 8'b00000000; // 1790 :   0 - 0x0
      12'h6FF: dout  = 8'b00000000; // 1791 :   0 - 0x0
      12'h700: dout  = 8'b00000000; // 1792 :   0 - 0x0 -- Sprite 0x70
      12'h701: dout  = 8'b00000000; // 1793 :   0 - 0x0
      12'h702: dout  = 8'b00000000; // 1794 :   0 - 0x0
      12'h703: dout  = 8'b00000000; // 1795 :   0 - 0x0
      12'h704: dout  = 8'b00000000; // 1796 :   0 - 0x0
      12'h705: dout  = 8'b00000000; // 1797 :   0 - 0x0
      12'h706: dout  = 8'b00000000; // 1798 :   0 - 0x0
      12'h707: dout  = 8'b00000000; // 1799 :   0 - 0x0
      12'h708: dout  = 8'b00000000; // 1800 :   0 - 0x0 -- plane 1
      12'h709: dout  = 8'b00000000; // 1801 :   0 - 0x0
      12'h70A: dout  = 8'b00000000; // 1802 :   0 - 0x0
      12'h70B: dout  = 8'b00000000; // 1803 :   0 - 0x0
      12'h70C: dout  = 8'b00000000; // 1804 :   0 - 0x0
      12'h70D: dout  = 8'b00000000; // 1805 :   0 - 0x0
      12'h70E: dout  = 8'b00000000; // 1806 :   0 - 0x0
      12'h70F: dout  = 8'b00000000; // 1807 :   0 - 0x0
      12'h710: dout  = 8'b00000000; // 1808 :   0 - 0x0 -- Sprite 0x71
      12'h711: dout  = 8'b00000000; // 1809 :   0 - 0x0
      12'h712: dout  = 8'b00000000; // 1810 :   0 - 0x0
      12'h713: dout  = 8'b00000000; // 1811 :   0 - 0x0
      12'h714: dout  = 8'b00000000; // 1812 :   0 - 0x0
      12'h715: dout  = 8'b00000000; // 1813 :   0 - 0x0
      12'h716: dout  = 8'b00000000; // 1814 :   0 - 0x0
      12'h717: dout  = 8'b00000000; // 1815 :   0 - 0x0
      12'h718: dout  = 8'b00000000; // 1816 :   0 - 0x0 -- plane 1
      12'h719: dout  = 8'b00000000; // 1817 :   0 - 0x0
      12'h71A: dout  = 8'b00000000; // 1818 :   0 - 0x0
      12'h71B: dout  = 8'b00000000; // 1819 :   0 - 0x0
      12'h71C: dout  = 8'b00000000; // 1820 :   0 - 0x0
      12'h71D: dout  = 8'b00000000; // 1821 :   0 - 0x0
      12'h71E: dout  = 8'b00000000; // 1822 :   0 - 0x0
      12'h71F: dout  = 8'b00000000; // 1823 :   0 - 0x0
      12'h720: dout  = 8'b00000000; // 1824 :   0 - 0x0 -- Sprite 0x72
      12'h721: dout  = 8'b00000000; // 1825 :   0 - 0x0
      12'h722: dout  = 8'b00000000; // 1826 :   0 - 0x0
      12'h723: dout  = 8'b00000000; // 1827 :   0 - 0x0
      12'h724: dout  = 8'b00000000; // 1828 :   0 - 0x0
      12'h725: dout  = 8'b00000000; // 1829 :   0 - 0x0
      12'h726: dout  = 8'b00000000; // 1830 :   0 - 0x0
      12'h727: dout  = 8'b00000000; // 1831 :   0 - 0x0
      12'h728: dout  = 8'b00000000; // 1832 :   0 - 0x0 -- plane 1
      12'h729: dout  = 8'b00000000; // 1833 :   0 - 0x0
      12'h72A: dout  = 8'b00000000; // 1834 :   0 - 0x0
      12'h72B: dout  = 8'b00000000; // 1835 :   0 - 0x0
      12'h72C: dout  = 8'b00000000; // 1836 :   0 - 0x0
      12'h72D: dout  = 8'b00000000; // 1837 :   0 - 0x0
      12'h72E: dout  = 8'b00000000; // 1838 :   0 - 0x0
      12'h72F: dout  = 8'b00000000; // 1839 :   0 - 0x0
      12'h730: dout  = 8'b00000000; // 1840 :   0 - 0x0 -- Sprite 0x73
      12'h731: dout  = 8'b00000000; // 1841 :   0 - 0x0
      12'h732: dout  = 8'b00000000; // 1842 :   0 - 0x0
      12'h733: dout  = 8'b00000000; // 1843 :   0 - 0x0
      12'h734: dout  = 8'b00000000; // 1844 :   0 - 0x0
      12'h735: dout  = 8'b00000000; // 1845 :   0 - 0x0
      12'h736: dout  = 8'b00000000; // 1846 :   0 - 0x0
      12'h737: dout  = 8'b00000000; // 1847 :   0 - 0x0
      12'h738: dout  = 8'b00000000; // 1848 :   0 - 0x0 -- plane 1
      12'h739: dout  = 8'b00000000; // 1849 :   0 - 0x0
      12'h73A: dout  = 8'b00000000; // 1850 :   0 - 0x0
      12'h73B: dout  = 8'b00000000; // 1851 :   0 - 0x0
      12'h73C: dout  = 8'b00000000; // 1852 :   0 - 0x0
      12'h73D: dout  = 8'b00000000; // 1853 :   0 - 0x0
      12'h73E: dout  = 8'b00000000; // 1854 :   0 - 0x0
      12'h73F: dout  = 8'b00000000; // 1855 :   0 - 0x0
      12'h740: dout  = 8'b00000000; // 1856 :   0 - 0x0 -- Sprite 0x74
      12'h741: dout  = 8'b00000000; // 1857 :   0 - 0x0
      12'h742: dout  = 8'b00000000; // 1858 :   0 - 0x0
      12'h743: dout  = 8'b00000000; // 1859 :   0 - 0x0
      12'h744: dout  = 8'b00000000; // 1860 :   0 - 0x0
      12'h745: dout  = 8'b00000000; // 1861 :   0 - 0x0
      12'h746: dout  = 8'b00000000; // 1862 :   0 - 0x0
      12'h747: dout  = 8'b00000000; // 1863 :   0 - 0x0
      12'h748: dout  = 8'b00000000; // 1864 :   0 - 0x0 -- plane 1
      12'h749: dout  = 8'b00000000; // 1865 :   0 - 0x0
      12'h74A: dout  = 8'b00000000; // 1866 :   0 - 0x0
      12'h74B: dout  = 8'b00000000; // 1867 :   0 - 0x0
      12'h74C: dout  = 8'b00000000; // 1868 :   0 - 0x0
      12'h74D: dout  = 8'b00000000; // 1869 :   0 - 0x0
      12'h74E: dout  = 8'b00000000; // 1870 :   0 - 0x0
      12'h74F: dout  = 8'b00000000; // 1871 :   0 - 0x0
      12'h750: dout  = 8'b00000000; // 1872 :   0 - 0x0 -- Sprite 0x75
      12'h751: dout  = 8'b00000000; // 1873 :   0 - 0x0
      12'h752: dout  = 8'b00000000; // 1874 :   0 - 0x0
      12'h753: dout  = 8'b00000000; // 1875 :   0 - 0x0
      12'h754: dout  = 8'b00000000; // 1876 :   0 - 0x0
      12'h755: dout  = 8'b00000000; // 1877 :   0 - 0x0
      12'h756: dout  = 8'b00000000; // 1878 :   0 - 0x0
      12'h757: dout  = 8'b00000000; // 1879 :   0 - 0x0
      12'h758: dout  = 8'b00000000; // 1880 :   0 - 0x0 -- plane 1
      12'h759: dout  = 8'b00000000; // 1881 :   0 - 0x0
      12'h75A: dout  = 8'b00000000; // 1882 :   0 - 0x0
      12'h75B: dout  = 8'b00000000; // 1883 :   0 - 0x0
      12'h75C: dout  = 8'b00000000; // 1884 :   0 - 0x0
      12'h75D: dout  = 8'b00000000; // 1885 :   0 - 0x0
      12'h75E: dout  = 8'b00000000; // 1886 :   0 - 0x0
      12'h75F: dout  = 8'b00000000; // 1887 :   0 - 0x0
      12'h760: dout  = 8'b00000000; // 1888 :   0 - 0x0 -- Sprite 0x76
      12'h761: dout  = 8'b00000000; // 1889 :   0 - 0x0
      12'h762: dout  = 8'b00000000; // 1890 :   0 - 0x0
      12'h763: dout  = 8'b00000000; // 1891 :   0 - 0x0
      12'h764: dout  = 8'b00000000; // 1892 :   0 - 0x0
      12'h765: dout  = 8'b00000000; // 1893 :   0 - 0x0
      12'h766: dout  = 8'b00000000; // 1894 :   0 - 0x0
      12'h767: dout  = 8'b00000000; // 1895 :   0 - 0x0
      12'h768: dout  = 8'b00000000; // 1896 :   0 - 0x0 -- plane 1
      12'h769: dout  = 8'b00000000; // 1897 :   0 - 0x0
      12'h76A: dout  = 8'b00000000; // 1898 :   0 - 0x0
      12'h76B: dout  = 8'b00000000; // 1899 :   0 - 0x0
      12'h76C: dout  = 8'b00000000; // 1900 :   0 - 0x0
      12'h76D: dout  = 8'b00000000; // 1901 :   0 - 0x0
      12'h76E: dout  = 8'b00000000; // 1902 :   0 - 0x0
      12'h76F: dout  = 8'b00000000; // 1903 :   0 - 0x0
      12'h770: dout  = 8'b00000000; // 1904 :   0 - 0x0 -- Sprite 0x77
      12'h771: dout  = 8'b00000000; // 1905 :   0 - 0x0
      12'h772: dout  = 8'b00000000; // 1906 :   0 - 0x0
      12'h773: dout  = 8'b00000000; // 1907 :   0 - 0x0
      12'h774: dout  = 8'b00000000; // 1908 :   0 - 0x0
      12'h775: dout  = 8'b00000000; // 1909 :   0 - 0x0
      12'h776: dout  = 8'b00000000; // 1910 :   0 - 0x0
      12'h777: dout  = 8'b00000000; // 1911 :   0 - 0x0
      12'h778: dout  = 8'b00000000; // 1912 :   0 - 0x0 -- plane 1
      12'h779: dout  = 8'b00000000; // 1913 :   0 - 0x0
      12'h77A: dout  = 8'b00000000; // 1914 :   0 - 0x0
      12'h77B: dout  = 8'b00000000; // 1915 :   0 - 0x0
      12'h77C: dout  = 8'b00000000; // 1916 :   0 - 0x0
      12'h77D: dout  = 8'b00000000; // 1917 :   0 - 0x0
      12'h77E: dout  = 8'b00000000; // 1918 :   0 - 0x0
      12'h77F: dout  = 8'b00000000; // 1919 :   0 - 0x0
      12'h780: dout  = 8'b00000000; // 1920 :   0 - 0x0 -- Sprite 0x78
      12'h781: dout  = 8'b00000000; // 1921 :   0 - 0x0
      12'h782: dout  = 8'b00000000; // 1922 :   0 - 0x0
      12'h783: dout  = 8'b00000000; // 1923 :   0 - 0x0
      12'h784: dout  = 8'b00000000; // 1924 :   0 - 0x0
      12'h785: dout  = 8'b00000000; // 1925 :   0 - 0x0
      12'h786: dout  = 8'b00000000; // 1926 :   0 - 0x0
      12'h787: dout  = 8'b00000000; // 1927 :   0 - 0x0
      12'h788: dout  = 8'b00000000; // 1928 :   0 - 0x0 -- plane 1
      12'h789: dout  = 8'b00000000; // 1929 :   0 - 0x0
      12'h78A: dout  = 8'b00000000; // 1930 :   0 - 0x0
      12'h78B: dout  = 8'b00000000; // 1931 :   0 - 0x0
      12'h78C: dout  = 8'b00000000; // 1932 :   0 - 0x0
      12'h78D: dout  = 8'b00000000; // 1933 :   0 - 0x0
      12'h78E: dout  = 8'b00000000; // 1934 :   0 - 0x0
      12'h78F: dout  = 8'b00000000; // 1935 :   0 - 0x0
      12'h790: dout  = 8'b00000000; // 1936 :   0 - 0x0 -- Sprite 0x79
      12'h791: dout  = 8'b00000000; // 1937 :   0 - 0x0
      12'h792: dout  = 8'b00000000; // 1938 :   0 - 0x0
      12'h793: dout  = 8'b00000000; // 1939 :   0 - 0x0
      12'h794: dout  = 8'b00000000; // 1940 :   0 - 0x0
      12'h795: dout  = 8'b00000000; // 1941 :   0 - 0x0
      12'h796: dout  = 8'b00000000; // 1942 :   0 - 0x0
      12'h797: dout  = 8'b00000000; // 1943 :   0 - 0x0
      12'h798: dout  = 8'b00000000; // 1944 :   0 - 0x0 -- plane 1
      12'h799: dout  = 8'b00000000; // 1945 :   0 - 0x0
      12'h79A: dout  = 8'b00000000; // 1946 :   0 - 0x0
      12'h79B: dout  = 8'b00000000; // 1947 :   0 - 0x0
      12'h79C: dout  = 8'b00000000; // 1948 :   0 - 0x0
      12'h79D: dout  = 8'b00000000; // 1949 :   0 - 0x0
      12'h79E: dout  = 8'b00000000; // 1950 :   0 - 0x0
      12'h79F: dout  = 8'b00000000; // 1951 :   0 - 0x0
      12'h7A0: dout  = 8'b00000000; // 1952 :   0 - 0x0 -- Sprite 0x7a
      12'h7A1: dout  = 8'b00000000; // 1953 :   0 - 0x0
      12'h7A2: dout  = 8'b00000000; // 1954 :   0 - 0x0
      12'h7A3: dout  = 8'b00000000; // 1955 :   0 - 0x0
      12'h7A4: dout  = 8'b00000000; // 1956 :   0 - 0x0
      12'h7A5: dout  = 8'b00000000; // 1957 :   0 - 0x0
      12'h7A6: dout  = 8'b00000000; // 1958 :   0 - 0x0
      12'h7A7: dout  = 8'b00000000; // 1959 :   0 - 0x0
      12'h7A8: dout  = 8'b00000000; // 1960 :   0 - 0x0 -- plane 1
      12'h7A9: dout  = 8'b00000000; // 1961 :   0 - 0x0
      12'h7AA: dout  = 8'b00000000; // 1962 :   0 - 0x0
      12'h7AB: dout  = 8'b00000000; // 1963 :   0 - 0x0
      12'h7AC: dout  = 8'b00000000; // 1964 :   0 - 0x0
      12'h7AD: dout  = 8'b00000000; // 1965 :   0 - 0x0
      12'h7AE: dout  = 8'b00000000; // 1966 :   0 - 0x0
      12'h7AF: dout  = 8'b00000000; // 1967 :   0 - 0x0
      12'h7B0: dout  = 8'b00000000; // 1968 :   0 - 0x0 -- Sprite 0x7b
      12'h7B1: dout  = 8'b00000000; // 1969 :   0 - 0x0
      12'h7B2: dout  = 8'b00000000; // 1970 :   0 - 0x0
      12'h7B3: dout  = 8'b00000000; // 1971 :   0 - 0x0
      12'h7B4: dout  = 8'b00000000; // 1972 :   0 - 0x0
      12'h7B5: dout  = 8'b00000000; // 1973 :   0 - 0x0
      12'h7B6: dout  = 8'b00000000; // 1974 :   0 - 0x0
      12'h7B7: dout  = 8'b00000000; // 1975 :   0 - 0x0
      12'h7B8: dout  = 8'b00000000; // 1976 :   0 - 0x0 -- plane 1
      12'h7B9: dout  = 8'b00000000; // 1977 :   0 - 0x0
      12'h7BA: dout  = 8'b00000000; // 1978 :   0 - 0x0
      12'h7BB: dout  = 8'b00000000; // 1979 :   0 - 0x0
      12'h7BC: dout  = 8'b00000000; // 1980 :   0 - 0x0
      12'h7BD: dout  = 8'b00000000; // 1981 :   0 - 0x0
      12'h7BE: dout  = 8'b00000000; // 1982 :   0 - 0x0
      12'h7BF: dout  = 8'b00000000; // 1983 :   0 - 0x0
      12'h7C0: dout  = 8'b00000000; // 1984 :   0 - 0x0 -- Sprite 0x7c
      12'h7C1: dout  = 8'b00000000; // 1985 :   0 - 0x0
      12'h7C2: dout  = 8'b00000000; // 1986 :   0 - 0x0
      12'h7C3: dout  = 8'b00000000; // 1987 :   0 - 0x0
      12'h7C4: dout  = 8'b00000000; // 1988 :   0 - 0x0
      12'h7C5: dout  = 8'b00000000; // 1989 :   0 - 0x0
      12'h7C6: dout  = 8'b00000000; // 1990 :   0 - 0x0
      12'h7C7: dout  = 8'b00000000; // 1991 :   0 - 0x0
      12'h7C8: dout  = 8'b00000000; // 1992 :   0 - 0x0 -- plane 1
      12'h7C9: dout  = 8'b00000000; // 1993 :   0 - 0x0
      12'h7CA: dout  = 8'b00000000; // 1994 :   0 - 0x0
      12'h7CB: dout  = 8'b00000000; // 1995 :   0 - 0x0
      12'h7CC: dout  = 8'b00000000; // 1996 :   0 - 0x0
      12'h7CD: dout  = 8'b00000000; // 1997 :   0 - 0x0
      12'h7CE: dout  = 8'b00000000; // 1998 :   0 - 0x0
      12'h7CF: dout  = 8'b00000000; // 1999 :   0 - 0x0
      12'h7D0: dout  = 8'b00000000; // 2000 :   0 - 0x0 -- Sprite 0x7d
      12'h7D1: dout  = 8'b00000000; // 2001 :   0 - 0x0
      12'h7D2: dout  = 8'b00000000; // 2002 :   0 - 0x0
      12'h7D3: dout  = 8'b00000000; // 2003 :   0 - 0x0
      12'h7D4: dout  = 8'b00000000; // 2004 :   0 - 0x0
      12'h7D5: dout  = 8'b00000000; // 2005 :   0 - 0x0
      12'h7D6: dout  = 8'b00000000; // 2006 :   0 - 0x0
      12'h7D7: dout  = 8'b00000000; // 2007 :   0 - 0x0
      12'h7D8: dout  = 8'b00000000; // 2008 :   0 - 0x0 -- plane 1
      12'h7D9: dout  = 8'b00000000; // 2009 :   0 - 0x0
      12'h7DA: dout  = 8'b00000000; // 2010 :   0 - 0x0
      12'h7DB: dout  = 8'b00000000; // 2011 :   0 - 0x0
      12'h7DC: dout  = 8'b00000000; // 2012 :   0 - 0x0
      12'h7DD: dout  = 8'b00000000; // 2013 :   0 - 0x0
      12'h7DE: dout  = 8'b00000000; // 2014 :   0 - 0x0
      12'h7DF: dout  = 8'b00000000; // 2015 :   0 - 0x0
      12'h7E0: dout  = 8'b00000000; // 2016 :   0 - 0x0 -- Sprite 0x7e
      12'h7E1: dout  = 8'b00000000; // 2017 :   0 - 0x0
      12'h7E2: dout  = 8'b00000000; // 2018 :   0 - 0x0
      12'h7E3: dout  = 8'b00000000; // 2019 :   0 - 0x0
      12'h7E4: dout  = 8'b00000000; // 2020 :   0 - 0x0
      12'h7E5: dout  = 8'b00000000; // 2021 :   0 - 0x0
      12'h7E6: dout  = 8'b00000000; // 2022 :   0 - 0x0
      12'h7E7: dout  = 8'b00000000; // 2023 :   0 - 0x0
      12'h7E8: dout  = 8'b00000000; // 2024 :   0 - 0x0 -- plane 1
      12'h7E9: dout  = 8'b00000000; // 2025 :   0 - 0x0
      12'h7EA: dout  = 8'b00000000; // 2026 :   0 - 0x0
      12'h7EB: dout  = 8'b00000000; // 2027 :   0 - 0x0
      12'h7EC: dout  = 8'b00000000; // 2028 :   0 - 0x0
      12'h7ED: dout  = 8'b00000000; // 2029 :   0 - 0x0
      12'h7EE: dout  = 8'b00000000; // 2030 :   0 - 0x0
      12'h7EF: dout  = 8'b00000000; // 2031 :   0 - 0x0
      12'h7F0: dout  = 8'b00000000; // 2032 :   0 - 0x0 -- Sprite 0x7f
      12'h7F1: dout  = 8'b00000000; // 2033 :   0 - 0x0
      12'h7F2: dout  = 8'b00000000; // 2034 :   0 - 0x0
      12'h7F3: dout  = 8'b00000000; // 2035 :   0 - 0x0
      12'h7F4: dout  = 8'b00000000; // 2036 :   0 - 0x0
      12'h7F5: dout  = 8'b00000000; // 2037 :   0 - 0x0
      12'h7F6: dout  = 8'b00000000; // 2038 :   0 - 0x0
      12'h7F7: dout  = 8'b00000000; // 2039 :   0 - 0x0
      12'h7F8: dout  = 8'b00000000; // 2040 :   0 - 0x0 -- plane 1
      12'h7F9: dout  = 8'b00000000; // 2041 :   0 - 0x0
      12'h7FA: dout  = 8'b00000000; // 2042 :   0 - 0x0
      12'h7FB: dout  = 8'b00000000; // 2043 :   0 - 0x0
      12'h7FC: dout  = 8'b00000000; // 2044 :   0 - 0x0
      12'h7FD: dout  = 8'b00000000; // 2045 :   0 - 0x0
      12'h7FE: dout  = 8'b00000000; // 2046 :   0 - 0x0
      12'h7FF: dout  = 8'b00000000; // 2047 :   0 - 0x0
      12'h800: dout  = 8'b00000011; // 2048 :   3 - 0x3 -- Sprite 0x80
      12'h801: dout  = 8'b00001111; // 2049 :  15 - 0xf
      12'h802: dout  = 8'b00011100; // 2050 :  28 - 0x1c
      12'h803: dout  = 8'b00110000; // 2051 :  48 - 0x30
      12'h804: dout  = 8'b00100000; // 2052 :  32 - 0x20
      12'h805: dout  = 8'b01000000; // 2053 :  64 - 0x40
      12'h806: dout  = 8'b01000000; // 2054 :  64 - 0x40
      12'h807: dout  = 8'b01111111; // 2055 : 127 - 0x7f
      12'h808: dout  = 8'b00000000; // 2056 :   0 - 0x0 -- plane 1
      12'h809: dout  = 8'b00000011; // 2057 :   3 - 0x3
      12'h80A: dout  = 8'b00001111; // 2058 :  15 - 0xf
      12'h80B: dout  = 8'b00011111; // 2059 :  31 - 0x1f
      12'h80C: dout  = 8'b00011111; // 2060 :  31 - 0x1f
      12'h80D: dout  = 8'b00111111; // 2061 :  63 - 0x3f
      12'h80E: dout  = 8'b00111111; // 2062 :  63 - 0x3f
      12'h80F: dout  = 8'b00000000; // 2063 :   0 - 0x0
      12'h810: dout  = 8'b00000001; // 2064 :   1 - 0x1 -- Sprite 0x81
      12'h811: dout  = 8'b00000001; // 2065 :   1 - 0x1
      12'h812: dout  = 8'b00000001; // 2066 :   1 - 0x1
      12'h813: dout  = 8'b00000001; // 2067 :   1 - 0x1
      12'h814: dout  = 8'b00000001; // 2068 :   1 - 0x1
      12'h815: dout  = 8'b00000001; // 2069 :   1 - 0x1
      12'h816: dout  = 8'b00000011; // 2070 :   3 - 0x3
      12'h817: dout  = 8'b00000011; // 2071 :   3 - 0x3
      12'h818: dout  = 8'b00000000; // 2072 :   0 - 0x0 -- plane 1
      12'h819: dout  = 8'b00000000; // 2073 :   0 - 0x0
      12'h81A: dout  = 8'b00000000; // 2074 :   0 - 0x0
      12'h81B: dout  = 8'b00000000; // 2075 :   0 - 0x0
      12'h81C: dout  = 8'b00000000; // 2076 :   0 - 0x0
      12'h81D: dout  = 8'b00000000; // 2077 :   0 - 0x0
      12'h81E: dout  = 8'b00000000; // 2078 :   0 - 0x0
      12'h81F: dout  = 8'b00000000; // 2079 :   0 - 0x0
      12'h820: dout  = 8'b11000000; // 2080 : 192 - 0xc0 -- Sprite 0x82
      12'h821: dout  = 8'b11110000; // 2081 : 240 - 0xf0
      12'h822: dout  = 8'b00111000; // 2082 :  56 - 0x38
      12'h823: dout  = 8'b00001110; // 2083 :  14 - 0xe
      12'h824: dout  = 8'b00011110; // 2084 :  30 - 0x1e
      12'h825: dout  = 8'b00011110; // 2085 :  30 - 0x1e
      12'h826: dout  = 8'b00000010; // 2086 :   2 - 0x2
      12'h827: dout  = 8'b11111110; // 2087 : 254 - 0xfe
      12'h828: dout  = 8'b00000000; // 2088 :   0 - 0x0 -- plane 1
      12'h829: dout  = 8'b11000000; // 2089 : 192 - 0xc0
      12'h82A: dout  = 8'b11110000; // 2090 : 240 - 0xf0
      12'h82B: dout  = 8'b11110000; // 2091 : 240 - 0xf0
      12'h82C: dout  = 8'b11101100; // 2092 : 236 - 0xec
      12'h82D: dout  = 8'b11100000; // 2093 : 224 - 0xe0
      12'h82E: dout  = 8'b11111100; // 2094 : 252 - 0xfc
      12'h82F: dout  = 8'b00000000; // 2095 :   0 - 0x0
      12'h830: dout  = 8'b10000000; // 2096 : 128 - 0x80 -- Sprite 0x83
      12'h831: dout  = 8'b10000000; // 2097 : 128 - 0x80
      12'h832: dout  = 8'b10000000; // 2098 : 128 - 0x80
      12'h833: dout  = 8'b10000000; // 2099 : 128 - 0x80
      12'h834: dout  = 8'b10000000; // 2100 : 128 - 0x80
      12'h835: dout  = 8'b11100000; // 2101 : 224 - 0xe0
      12'h836: dout  = 8'b00010000; // 2102 :  16 - 0x10
      12'h837: dout  = 8'b11110000; // 2103 : 240 - 0xf0
      12'h838: dout  = 8'b00000000; // 2104 :   0 - 0x0 -- plane 1
      12'h839: dout  = 8'b00000000; // 2105 :   0 - 0x0
      12'h83A: dout  = 8'b00000000; // 2106 :   0 - 0x0
      12'h83B: dout  = 8'b00000000; // 2107 :   0 - 0x0
      12'h83C: dout  = 8'b00000000; // 2108 :   0 - 0x0
      12'h83D: dout  = 8'b00000000; // 2109 :   0 - 0x0
      12'h83E: dout  = 8'b11100000; // 2110 : 224 - 0xe0
      12'h83F: dout  = 8'b00000000; // 2111 :   0 - 0x0
      12'h840: dout  = 8'b00000011; // 2112 :   3 - 0x3 -- Sprite 0x84
      12'h841: dout  = 8'b00001111; // 2113 :  15 - 0xf
      12'h842: dout  = 8'b00011100; // 2114 :  28 - 0x1c
      12'h843: dout  = 8'b00110000; // 2115 :  48 - 0x30
      12'h844: dout  = 8'b00100000; // 2116 :  32 - 0x20
      12'h845: dout  = 8'b01000000; // 2117 :  64 - 0x40
      12'h846: dout  = 8'b01000000; // 2118 :  64 - 0x40
      12'h847: dout  = 8'b01111111; // 2119 : 127 - 0x7f
      12'h848: dout  = 8'b00000000; // 2120 :   0 - 0x0 -- plane 1
      12'h849: dout  = 8'b00000011; // 2121 :   3 - 0x3
      12'h84A: dout  = 8'b00001111; // 2122 :  15 - 0xf
      12'h84B: dout  = 8'b00011111; // 2123 :  31 - 0x1f
      12'h84C: dout  = 8'b00011111; // 2124 :  31 - 0x1f
      12'h84D: dout  = 8'b00111111; // 2125 :  63 - 0x3f
      12'h84E: dout  = 8'b00111111; // 2126 :  63 - 0x3f
      12'h84F: dout  = 8'b00000000; // 2127 :   0 - 0x0
      12'h850: dout  = 8'b00000011; // 2128 :   3 - 0x3 -- Sprite 0x85
      12'h851: dout  = 8'b00000110; // 2129 :   6 - 0x6
      12'h852: dout  = 8'b00000110; // 2130 :   6 - 0x6
      12'h853: dout  = 8'b00011100; // 2131 :  28 - 0x1c
      12'h854: dout  = 8'b00011000; // 2132 :  24 - 0x18
      12'h855: dout  = 8'b00110110; // 2133 :  54 - 0x36
      12'h856: dout  = 8'b00110001; // 2134 :  49 - 0x31
      12'h857: dout  = 8'b00001111; // 2135 :  15 - 0xf
      12'h858: dout  = 8'b00000000; // 2136 :   0 - 0x0 -- plane 1
      12'h859: dout  = 8'b00000000; // 2137 :   0 - 0x0
      12'h85A: dout  = 8'b00000000; // 2138 :   0 - 0x0
      12'h85B: dout  = 8'b00000000; // 2139 :   0 - 0x0
      12'h85C: dout  = 8'b00000000; // 2140 :   0 - 0x0
      12'h85D: dout  = 8'b00001000; // 2141 :   8 - 0x8
      12'h85E: dout  = 8'b00001110; // 2142 :  14 - 0xe
      12'h85F: dout  = 8'b00000000; // 2143 :   0 - 0x0
      12'h860: dout  = 8'b11000000; // 2144 : 192 - 0xc0 -- Sprite 0x86
      12'h861: dout  = 8'b11110000; // 2145 : 240 - 0xf0
      12'h862: dout  = 8'b00111000; // 2146 :  56 - 0x38
      12'h863: dout  = 8'b00001110; // 2147 :  14 - 0xe
      12'h864: dout  = 8'b00011110; // 2148 :  30 - 0x1e
      12'h865: dout  = 8'b00011110; // 2149 :  30 - 0x1e
      12'h866: dout  = 8'b00000010; // 2150 :   2 - 0x2
      12'h867: dout  = 8'b11111110; // 2151 : 254 - 0xfe
      12'h868: dout  = 8'b00000000; // 2152 :   0 - 0x0 -- plane 1
      12'h869: dout  = 8'b11000000; // 2153 : 192 - 0xc0
      12'h86A: dout  = 8'b11110000; // 2154 : 240 - 0xf0
      12'h86B: dout  = 8'b11110000; // 2155 : 240 - 0xf0
      12'h86C: dout  = 8'b11101100; // 2156 : 236 - 0xec
      12'h86D: dout  = 8'b11100000; // 2157 : 224 - 0xe0
      12'h86E: dout  = 8'b11111100; // 2158 : 252 - 0xfc
      12'h86F: dout  = 8'b00000000; // 2159 :   0 - 0x0
      12'h870: dout  = 8'b11000000; // 2160 : 192 - 0xc0 -- Sprite 0x87
      12'h871: dout  = 8'b01100000; // 2161 :  96 - 0x60
      12'h872: dout  = 8'b01100000; // 2162 :  96 - 0x60
      12'h873: dout  = 8'b00110000; // 2163 :  48 - 0x30
      12'h874: dout  = 8'b00111110; // 2164 :  62 - 0x3e
      12'h875: dout  = 8'b00011001; // 2165 :  25 - 0x19
      12'h876: dout  = 8'b00110011; // 2166 :  51 - 0x33
      12'h877: dout  = 8'b00111100; // 2167 :  60 - 0x3c
      12'h878: dout  = 8'b00000000; // 2168 :   0 - 0x0 -- plane 1
      12'h879: dout  = 8'b00000000; // 2169 :   0 - 0x0
      12'h87A: dout  = 8'b00000000; // 2170 :   0 - 0x0
      12'h87B: dout  = 8'b00000000; // 2171 :   0 - 0x0
      12'h87C: dout  = 8'b00000000; // 2172 :   0 - 0x0
      12'h87D: dout  = 8'b00000110; // 2173 :   6 - 0x6
      12'h87E: dout  = 8'b00001100; // 2174 :  12 - 0xc
      12'h87F: dout  = 8'b00000000; // 2175 :   0 - 0x0
      12'h880: dout  = 8'b00000011; // 2176 :   3 - 0x3 -- Sprite 0x88
      12'h881: dout  = 8'b00000111; // 2177 :   7 - 0x7
      12'h882: dout  = 8'b00000111; // 2178 :   7 - 0x7
      12'h883: dout  = 8'b00001011; // 2179 :  11 - 0xb
      12'h884: dout  = 8'b00010000; // 2180 :  16 - 0x10
      12'h885: dout  = 8'b01100000; // 2181 :  96 - 0x60
      12'h886: dout  = 8'b11110000; // 2182 : 240 - 0xf0
      12'h887: dout  = 8'b11110000; // 2183 : 240 - 0xf0
      12'h888: dout  = 8'b00000000; // 2184 :   0 - 0x0 -- plane 1
      12'h889: dout  = 8'b00000011; // 2185 :   3 - 0x3
      12'h88A: dout  = 8'b00000011; // 2186 :   3 - 0x3
      12'h88B: dout  = 8'b00000100; // 2187 :   4 - 0x4
      12'h88C: dout  = 8'b00001111; // 2188 :  15 - 0xf
      12'h88D: dout  = 8'b00011111; // 2189 :  31 - 0x1f
      12'h88E: dout  = 8'b01101111; // 2190 : 111 - 0x6f
      12'h88F: dout  = 8'b01101111; // 2191 : 111 - 0x6f
      12'h890: dout  = 8'b11110000; // 2192 : 240 - 0xf0 -- Sprite 0x89
      12'h891: dout  = 8'b11110000; // 2193 : 240 - 0xf0
      12'h892: dout  = 8'b01100000; // 2194 :  96 - 0x60
      12'h893: dout  = 8'b00010000; // 2195 :  16 - 0x10
      12'h894: dout  = 8'b00001011; // 2196 :  11 - 0xb
      12'h895: dout  = 8'b00000111; // 2197 :   7 - 0x7
      12'h896: dout  = 8'b00000111; // 2198 :   7 - 0x7
      12'h897: dout  = 8'b00000011; // 2199 :   3 - 0x3
      12'h898: dout  = 8'b01101111; // 2200 : 111 - 0x6f -- plane 1
      12'h899: dout  = 8'b01101111; // 2201 : 111 - 0x6f
      12'h89A: dout  = 8'b00011111; // 2202 :  31 - 0x1f
      12'h89B: dout  = 8'b00001111; // 2203 :  15 - 0xf
      12'h89C: dout  = 8'b00000100; // 2204 :   4 - 0x4
      12'h89D: dout  = 8'b00000011; // 2205 :   3 - 0x3
      12'h89E: dout  = 8'b00000011; // 2206 :   3 - 0x3
      12'h89F: dout  = 8'b00000000; // 2207 :   0 - 0x0
      12'h8A0: dout  = 8'b00000000; // 2208 :   0 - 0x0 -- Sprite 0x8a
      12'h8A1: dout  = 8'b00011100; // 2209 :  28 - 0x1c
      12'h8A2: dout  = 8'b00111111; // 2210 :  63 - 0x3f
      12'h8A3: dout  = 8'b01111000; // 2211 : 120 - 0x78
      12'h8A4: dout  = 8'b01110000; // 2212 : 112 - 0x70
      12'h8A5: dout  = 8'b01100000; // 2213 :  96 - 0x60
      12'h8A6: dout  = 8'b00100000; // 2214 :  32 - 0x20
      12'h8A7: dout  = 8'b00100000; // 2215 :  32 - 0x20
      12'h8A8: dout  = 8'b00000000; // 2216 :   0 - 0x0 -- plane 1
      12'h8A9: dout  = 8'b00000000; // 2217 :   0 - 0x0
      12'h8AA: dout  = 8'b00011000; // 2218 :  24 - 0x18
      12'h8AB: dout  = 8'b00110111; // 2219 :  55 - 0x37
      12'h8AC: dout  = 8'b00101111; // 2220 :  47 - 0x2f
      12'h8AD: dout  = 8'b00011111; // 2221 :  31 - 0x1f
      12'h8AE: dout  = 8'b00011111; // 2222 :  31 - 0x1f
      12'h8AF: dout  = 8'b00011111; // 2223 :  31 - 0x1f
      12'h8B0: dout  = 8'b00100000; // 2224 :  32 - 0x20 -- Sprite 0x8b
      12'h8B1: dout  = 8'b00100000; // 2225 :  32 - 0x20
      12'h8B2: dout  = 8'b01100000; // 2226 :  96 - 0x60
      12'h8B3: dout  = 8'b01110000; // 2227 : 112 - 0x70
      12'h8B4: dout  = 8'b01111000; // 2228 : 120 - 0x78
      12'h8B5: dout  = 8'b00111111; // 2229 :  63 - 0x3f
      12'h8B6: dout  = 8'b00011100; // 2230 :  28 - 0x1c
      12'h8B7: dout  = 8'b00000000; // 2231 :   0 - 0x0
      12'h8B8: dout  = 8'b00011111; // 2232 :  31 - 0x1f -- plane 1
      12'h8B9: dout  = 8'b00011111; // 2233 :  31 - 0x1f
      12'h8BA: dout  = 8'b00011111; // 2234 :  31 - 0x1f
      12'h8BB: dout  = 8'b00101111; // 2235 :  47 - 0x2f
      12'h8BC: dout  = 8'b00110111; // 2236 :  55 - 0x37
      12'h8BD: dout  = 8'b00011000; // 2237 :  24 - 0x18
      12'h8BE: dout  = 8'b00000000; // 2238 :   0 - 0x0
      12'h8BF: dout  = 8'b00000000; // 2239 :   0 - 0x0
      12'h8C0: dout  = 8'b00000011; // 2240 :   3 - 0x3 -- Sprite 0x8c
      12'h8C1: dout  = 8'b00001100; // 2241 :  12 - 0xc
      12'h8C2: dout  = 8'b00011110; // 2242 :  30 - 0x1e
      12'h8C3: dout  = 8'b00100110; // 2243 :  38 - 0x26
      12'h8C4: dout  = 8'b01000110; // 2244 :  70 - 0x46
      12'h8C5: dout  = 8'b01100100; // 2245 : 100 - 0x64
      12'h8C6: dout  = 8'b01110000; // 2246 : 112 - 0x70
      12'h8C7: dout  = 8'b11110000; // 2247 : 240 - 0xf0
      12'h8C8: dout  = 8'b00000000; // 2248 :   0 - 0x0 -- plane 1
      12'h8C9: dout  = 8'b00000011; // 2249 :   3 - 0x3
      12'h8CA: dout  = 8'b00000001; // 2250 :   1 - 0x1
      12'h8CB: dout  = 8'b00011001; // 2251 :  25 - 0x19
      12'h8CC: dout  = 8'b00111001; // 2252 :  57 - 0x39
      12'h8CD: dout  = 8'b00011011; // 2253 :  27 - 0x1b
      12'h8CE: dout  = 8'b00001111; // 2254 :  15 - 0xf
      12'h8CF: dout  = 8'b00001111; // 2255 :  15 - 0xf
      12'h8D0: dout  = 8'b10101010; // 2256 : 170 - 0xaa -- Sprite 0x8d
      12'h8D1: dout  = 8'b11111111; // 2257 : 255 - 0xff
      12'h8D2: dout  = 8'b01111111; // 2258 : 127 - 0x7f
      12'h8D3: dout  = 8'b00111001; // 2259 :  57 - 0x39
      12'h8D4: dout  = 8'b00011001; // 2260 :  25 - 0x19
      12'h8D5: dout  = 8'b00001011; // 2261 :  11 - 0xb
      12'h8D6: dout  = 8'b00001000; // 2262 :   8 - 0x8
      12'h8D7: dout  = 8'b00000111; // 2263 :   7 - 0x7
      12'h8D8: dout  = 8'b01111111; // 2264 : 127 - 0x7f -- plane 1
      12'h8D9: dout  = 8'b01111111; // 2265 : 127 - 0x7f
      12'h8DA: dout  = 8'b00111111; // 2266 :  63 - 0x3f
      12'h8DB: dout  = 8'b00010111; // 2267 :  23 - 0x17
      12'h8DC: dout  = 8'b00000110; // 2268 :   6 - 0x6
      12'h8DD: dout  = 8'b00000100; // 2269 :   4 - 0x4
      12'h8DE: dout  = 8'b00000111; // 2270 :   7 - 0x7
      12'h8DF: dout  = 8'b00000000; // 2271 :   0 - 0x0
      12'h8E0: dout  = 8'b11000000; // 2272 : 192 - 0xc0 -- Sprite 0x8e
      12'h8E1: dout  = 8'b00110000; // 2273 :  48 - 0x30
      12'h8E2: dout  = 8'b00001000; // 2274 :   8 - 0x8
      12'h8E3: dout  = 8'b01000100; // 2275 :  68 - 0x44
      12'h8E4: dout  = 8'b01100010; // 2276 :  98 - 0x62
      12'h8E5: dout  = 8'b01100010; // 2277 :  98 - 0x62
      12'h8E6: dout  = 8'b00000001; // 2278 :   1 - 0x1
      12'h8E7: dout  = 8'b00111111; // 2279 :  63 - 0x3f
      12'h8E8: dout  = 8'b00000000; // 2280 :   0 - 0x0 -- plane 1
      12'h8E9: dout  = 8'b11000000; // 2281 : 192 - 0xc0
      12'h8EA: dout  = 8'b11110000; // 2282 : 240 - 0xf0
      12'h8EB: dout  = 8'b10111000; // 2283 : 184 - 0xb8
      12'h8EC: dout  = 8'b10011100; // 2284 : 156 - 0x9c
      12'h8ED: dout  = 8'b11111100; // 2285 : 252 - 0xfc
      12'h8EE: dout  = 8'b11111110; // 2286 : 254 - 0xfe
      12'h8EF: dout  = 8'b11000000; // 2287 : 192 - 0xc0
      12'h8F0: dout  = 8'b10001011; // 2288 : 139 - 0x8b -- Sprite 0x8f
      12'h8F1: dout  = 8'b11000001; // 2289 : 193 - 0xc1
      12'h8F2: dout  = 8'b11111110; // 2290 : 254 - 0xfe
      12'h8F3: dout  = 8'b11111100; // 2291 : 252 - 0xfc
      12'h8F4: dout  = 8'b11110000; // 2292 : 240 - 0xf0
      12'h8F5: dout  = 8'b11110000; // 2293 : 240 - 0xf0
      12'h8F6: dout  = 8'b11111000; // 2294 : 248 - 0xf8
      12'h8F7: dout  = 8'b11110000; // 2295 : 240 - 0xf0
      12'h8F8: dout  = 8'b11111110; // 2296 : 254 - 0xfe -- plane 1
      12'h8F9: dout  = 8'b11111110; // 2297 : 254 - 0xfe
      12'h8FA: dout  = 8'b11111000; // 2298 : 248 - 0xf8
      12'h8FB: dout  = 8'b11110000; // 2299 : 240 - 0xf0
      12'h8FC: dout  = 8'b11000000; // 2300 : 192 - 0xc0
      12'h8FD: dout  = 8'b00000000; // 2301 :   0 - 0x0
      12'h8FE: dout  = 8'b00000000; // 2302 :   0 - 0x0
      12'h8FF: dout  = 8'b10000000; // 2303 : 128 - 0x80
      12'h900: dout  = 8'b00000011; // 2304 :   3 - 0x3 -- Sprite 0x90
      12'h901: dout  = 8'b00001110; // 2305 :  14 - 0xe
      12'h902: dout  = 8'b00010110; // 2306 :  22 - 0x16
      12'h903: dout  = 8'b00100110; // 2307 :  38 - 0x26
      12'h904: dout  = 8'b01100011; // 2308 :  99 - 0x63
      12'h905: dout  = 8'b01110010; // 2309 : 114 - 0x72
      12'h906: dout  = 8'b01110000; // 2310 : 112 - 0x70
      12'h907: dout  = 8'b11010000; // 2311 : 208 - 0xd0
      12'h908: dout  = 8'b00000000; // 2312 :   0 - 0x0 -- plane 1
      12'h909: dout  = 8'b00000001; // 2313 :   1 - 0x1
      12'h90A: dout  = 8'b00001001; // 2314 :   9 - 0x9
      12'h90B: dout  = 8'b00011001; // 2315 :  25 - 0x19
      12'h90C: dout  = 8'b00011100; // 2316 :  28 - 0x1c
      12'h90D: dout  = 8'b00001101; // 2317 :  13 - 0xd
      12'h90E: dout  = 8'b00001111; // 2318 :  15 - 0xf
      12'h90F: dout  = 8'b00101111; // 2319 :  47 - 0x2f
      12'h910: dout  = 8'b10101010; // 2320 : 170 - 0xaa -- Sprite 0x91
      12'h911: dout  = 8'b11111111; // 2321 : 255 - 0xff
      12'h912: dout  = 8'b01111111; // 2322 : 127 - 0x7f
      12'h913: dout  = 8'b00111100; // 2323 :  60 - 0x3c
      12'h914: dout  = 8'b00011100; // 2324 :  28 - 0x1c
      12'h915: dout  = 8'b00000100; // 2325 :   4 - 0x4
      12'h916: dout  = 8'b00000010; // 2326 :   2 - 0x2
      12'h917: dout  = 8'b00000001; // 2327 :   1 - 0x1
      12'h918: dout  = 8'b01111111; // 2328 : 127 - 0x7f -- plane 1
      12'h919: dout  = 8'b01111111; // 2329 : 127 - 0x7f
      12'h91A: dout  = 8'b00111111; // 2330 :  63 - 0x3f
      12'h91B: dout  = 8'b00011011; // 2331 :  27 - 0x1b
      12'h91C: dout  = 8'b00000011; // 2332 :   3 - 0x3
      12'h91D: dout  = 8'b00000011; // 2333 :   3 - 0x3
      12'h91E: dout  = 8'b00000001; // 2334 :   1 - 0x1
      12'h91F: dout  = 8'b00000000; // 2335 :   0 - 0x0
      12'h920: dout  = 8'b11000000; // 2336 : 192 - 0xc0 -- Sprite 0x92
      12'h921: dout  = 8'b00110000; // 2337 :  48 - 0x30
      12'h922: dout  = 8'b00001000; // 2338 :   8 - 0x8
      12'h923: dout  = 8'b00100100; // 2339 :  36 - 0x24
      12'h924: dout  = 8'b00110010; // 2340 :  50 - 0x32
      12'h925: dout  = 8'b00110010; // 2341 :  50 - 0x32
      12'h926: dout  = 8'b00000001; // 2342 :   1 - 0x1
      12'h927: dout  = 8'b00011111; // 2343 :  31 - 0x1f
      12'h928: dout  = 8'b00000000; // 2344 :   0 - 0x0 -- plane 1
      12'h929: dout  = 8'b11000000; // 2345 : 192 - 0xc0
      12'h92A: dout  = 8'b11110000; // 2346 : 240 - 0xf0
      12'h92B: dout  = 8'b11011000; // 2347 : 216 - 0xd8
      12'h92C: dout  = 8'b11001100; // 2348 : 204 - 0xcc
      12'h92D: dout  = 8'b11111100; // 2349 : 252 - 0xfc
      12'h92E: dout  = 8'b11111110; // 2350 : 254 - 0xfe
      12'h92F: dout  = 8'b11100000; // 2351 : 224 - 0xe0
      12'h930: dout  = 8'b10001011; // 2352 : 139 - 0x8b -- Sprite 0x93
      12'h931: dout  = 8'b11000001; // 2353 : 193 - 0xc1
      12'h932: dout  = 8'b11111110; // 2354 : 254 - 0xfe
      12'h933: dout  = 8'b11111100; // 2355 : 252 - 0xfc
      12'h934: dout  = 8'b11110000; // 2356 : 240 - 0xf0
      12'h935: dout  = 8'b11000000; // 2357 : 192 - 0xc0
      12'h936: dout  = 8'b00100000; // 2358 :  32 - 0x20
      12'h937: dout  = 8'b11100000; // 2359 : 224 - 0xe0
      12'h938: dout  = 8'b11111110; // 2360 : 254 - 0xfe -- plane 1
      12'h939: dout  = 8'b11111110; // 2361 : 254 - 0xfe
      12'h93A: dout  = 8'b11111000; // 2362 : 248 - 0xf8
      12'h93B: dout  = 8'b01110000; // 2363 : 112 - 0x70
      12'h93C: dout  = 8'b01000000; // 2364 :  64 - 0x40
      12'h93D: dout  = 8'b00000000; // 2365 :   0 - 0x0
      12'h93E: dout  = 8'b11000000; // 2366 : 192 - 0xc0
      12'h93F: dout  = 8'b00100000; // 2367 :  32 - 0x20
      12'h940: dout  = 8'b00000011; // 2368 :   3 - 0x3 -- Sprite 0x94
      12'h941: dout  = 8'b00001111; // 2369 :  15 - 0xf
      12'h942: dout  = 8'b00010011; // 2370 :  19 - 0x13
      12'h943: dout  = 8'b00110001; // 2371 :  49 - 0x31
      12'h944: dout  = 8'b01111001; // 2372 : 121 - 0x79
      12'h945: dout  = 8'b01011001; // 2373 :  89 - 0x59
      12'h946: dout  = 8'b01001000; // 2374 :  72 - 0x48
      12'h947: dout  = 8'b11001100; // 2375 : 204 - 0xcc
      12'h948: dout  = 8'b00000000; // 2376 :   0 - 0x0 -- plane 1
      12'h949: dout  = 8'b00000000; // 2377 :   0 - 0x0
      12'h94A: dout  = 8'b00001100; // 2378 :  12 - 0xc
      12'h94B: dout  = 8'b00001110; // 2379 :  14 - 0xe
      12'h94C: dout  = 8'b00000110; // 2380 :   6 - 0x6
      12'h94D: dout  = 8'b00100110; // 2381 :  38 - 0x26
      12'h94E: dout  = 8'b00110111; // 2382 :  55 - 0x37
      12'h94F: dout  = 8'b00110011; // 2383 :  51 - 0x33
      12'h950: dout  = 8'b10010101; // 2384 : 149 - 0x95 -- Sprite 0x95
      12'h951: dout  = 8'b11111111; // 2385 : 255 - 0xff
      12'h952: dout  = 8'b01111111; // 2386 : 127 - 0x7f
      12'h953: dout  = 8'b00111110; // 2387 :  62 - 0x3e
      12'h954: dout  = 8'b00011111; // 2388 :  31 - 0x1f
      12'h955: dout  = 8'b00001111; // 2389 :  15 - 0xf
      12'h956: dout  = 8'b00001111; // 2390 :  15 - 0xf
      12'h957: dout  = 8'b00000111; // 2391 :   7 - 0x7
      12'h958: dout  = 8'b01111111; // 2392 : 127 - 0x7f -- plane 1
      12'h959: dout  = 8'b01111111; // 2393 : 127 - 0x7f
      12'h95A: dout  = 8'b00111111; // 2394 :  63 - 0x3f
      12'h95B: dout  = 8'b00011111; // 2395 :  31 - 0x1f
      12'h95C: dout  = 8'b00001110; // 2396 :  14 - 0xe
      12'h95D: dout  = 8'b00000000; // 2397 :   0 - 0x0
      12'h95E: dout  = 8'b00000000; // 2398 :   0 - 0x0
      12'h95F: dout  = 8'b00000000; // 2399 :   0 - 0x0
      12'h960: dout  = 8'b11000000; // 2400 : 192 - 0xc0 -- Sprite 0x96
      12'h961: dout  = 8'b00110000; // 2401 :  48 - 0x30
      12'h962: dout  = 8'b00001000; // 2402 :   8 - 0x8
      12'h963: dout  = 8'b10010100; // 2403 : 148 - 0x94
      12'h964: dout  = 8'b10011010; // 2404 : 154 - 0x9a
      12'h965: dout  = 8'b00011010; // 2405 :  26 - 0x1a
      12'h966: dout  = 8'b00000001; // 2406 :   1 - 0x1
      12'h967: dout  = 8'b00001111; // 2407 :  15 - 0xf
      12'h968: dout  = 8'b00000000; // 2408 :   0 - 0x0 -- plane 1
      12'h969: dout  = 8'b11000000; // 2409 : 192 - 0xc0
      12'h96A: dout  = 8'b11110000; // 2410 : 240 - 0xf0
      12'h96B: dout  = 8'b01101000; // 2411 : 104 - 0x68
      12'h96C: dout  = 8'b01100100; // 2412 : 100 - 0x64
      12'h96D: dout  = 8'b11111100; // 2413 : 252 - 0xfc
      12'h96E: dout  = 8'b11111110; // 2414 : 254 - 0xfe
      12'h96F: dout  = 8'b11110000; // 2415 : 240 - 0xf0
      12'h970: dout  = 8'b01000101; // 2416 :  69 - 0x45 -- Sprite 0x97
      12'h971: dout  = 8'b11100001; // 2417 : 225 - 0xe1
      12'h972: dout  = 8'b11111110; // 2418 : 254 - 0xfe
      12'h973: dout  = 8'b01111100; // 2419 : 124 - 0x7c
      12'h974: dout  = 8'b00110000; // 2420 :  48 - 0x30
      12'h975: dout  = 8'b00110000; // 2421 :  48 - 0x30
      12'h976: dout  = 8'b10001000; // 2422 : 136 - 0x88
      12'h977: dout  = 8'b01111000; // 2423 : 120 - 0x78
      12'h978: dout  = 8'b11111111; // 2424 : 255 - 0xff -- plane 1
      12'h979: dout  = 8'b11111110; // 2425 : 254 - 0xfe
      12'h97A: dout  = 8'b11111100; // 2426 : 252 - 0xfc
      12'h97B: dout  = 8'b10110000; // 2427 : 176 - 0xb0
      12'h97C: dout  = 8'b11000000; // 2428 : 192 - 0xc0
      12'h97D: dout  = 8'b11000000; // 2429 : 192 - 0xc0
      12'h97E: dout  = 8'b01110000; // 2430 : 112 - 0x70
      12'h97F: dout  = 8'b00001000; // 2431 :   8 - 0x8
      12'h980: dout  = 8'b00000001; // 2432 :   1 - 0x1 -- Sprite 0x98
      12'h981: dout  = 8'b00000000; // 2433 :   0 - 0x0
      12'h982: dout  = 8'b00000000; // 2434 :   0 - 0x0
      12'h983: dout  = 8'b00000000; // 2435 :   0 - 0x0
      12'h984: dout  = 8'b00000001; // 2436 :   1 - 0x1
      12'h985: dout  = 8'b00000001; // 2437 :   1 - 0x1
      12'h986: dout  = 8'b00000010; // 2438 :   2 - 0x2
      12'h987: dout  = 8'b00000110; // 2439 :   6 - 0x6
      12'h988: dout  = 8'b00000000; // 2440 :   0 - 0x0 -- plane 1
      12'h989: dout  = 8'b00000001; // 2441 :   1 - 0x1
      12'h98A: dout  = 8'b00000000; // 2442 :   0 - 0x0
      12'h98B: dout  = 8'b00000000; // 2443 :   0 - 0x0
      12'h98C: dout  = 8'b00000000; // 2444 :   0 - 0x0
      12'h98D: dout  = 8'b00000000; // 2445 :   0 - 0x0
      12'h98E: dout  = 8'b00000001; // 2446 :   1 - 0x1
      12'h98F: dout  = 8'b00000011; // 2447 :   3 - 0x3
      12'h990: dout  = 8'b01111000; // 2448 : 120 - 0x78 -- Sprite 0x99
      12'h991: dout  = 8'b00101010; // 2449 :  42 - 0x2a
      12'h992: dout  = 8'b01010100; // 2450 :  84 - 0x54
      12'h993: dout  = 8'b00101001; // 2451 :  41 - 0x29
      12'h994: dout  = 8'b00101111; // 2452 :  47 - 0x2f
      12'h995: dout  = 8'b00110111; // 2453 :  55 - 0x37
      12'h996: dout  = 8'b00000011; // 2454 :   3 - 0x3
      12'h997: dout  = 8'b00000111; // 2455 :   7 - 0x7
      12'h998: dout  = 8'b00000111; // 2456 :   7 - 0x7 -- plane 1
      12'h999: dout  = 8'b00010111; // 2457 :  23 - 0x17
      12'h99A: dout  = 8'b00101111; // 2458 :  47 - 0x2f
      12'h99B: dout  = 8'b00011110; // 2459 :  30 - 0x1e
      12'h99C: dout  = 8'b00010001; // 2460 :  17 - 0x11
      12'h99D: dout  = 8'b00000000; // 2461 :   0 - 0x0
      12'h99E: dout  = 8'b00000001; // 2462 :   1 - 0x1
      12'h99F: dout  = 8'b00000000; // 2463 :   0 - 0x0
      12'h9A0: dout  = 8'b10110000; // 2464 : 176 - 0xb0 -- Sprite 0x9a
      12'h9A1: dout  = 8'b11101000; // 2465 : 232 - 0xe8
      12'h9A2: dout  = 8'b10001100; // 2466 : 140 - 0x8c
      12'h9A3: dout  = 8'b10011110; // 2467 : 158 - 0x9e
      12'h9A4: dout  = 8'b00011111; // 2468 :  31 - 0x1f
      12'h9A5: dout  = 8'b00001111; // 2469 :  15 - 0xf
      12'h9A6: dout  = 8'b10010110; // 2470 : 150 - 0x96
      12'h9A7: dout  = 8'b00011100; // 2471 :  28 - 0x1c
      12'h9A8: dout  = 8'b00000000; // 2472 :   0 - 0x0 -- plane 1
      12'h9A9: dout  = 8'b00010000; // 2473 :  16 - 0x10
      12'h9AA: dout  = 8'b01111000; // 2474 : 120 - 0x78
      12'h9AB: dout  = 8'b01110100; // 2475 : 116 - 0x74
      12'h9AC: dout  = 8'b11111110; // 2476 : 254 - 0xfe
      12'h9AD: dout  = 8'b11111000; // 2477 : 248 - 0xf8
      12'h9AE: dout  = 8'b11111100; // 2478 : 252 - 0xfc
      12'h9AF: dout  = 8'b11111000; // 2479 : 248 - 0xf8
      12'h9B0: dout  = 8'b00001100; // 2480 :  12 - 0xc -- Sprite 0x9b
      12'h9B1: dout  = 8'b00111000; // 2481 :  56 - 0x38
      12'h9B2: dout  = 8'b11101000; // 2482 : 232 - 0xe8
      12'h9B3: dout  = 8'b11010000; // 2483 : 208 - 0xd0
      12'h9B4: dout  = 8'b11100000; // 2484 : 224 - 0xe0
      12'h9B5: dout  = 8'b10000000; // 2485 : 128 - 0x80
      12'h9B6: dout  = 8'b00000000; // 2486 :   0 - 0x0
      12'h9B7: dout  = 8'b10000000; // 2487 : 128 - 0x80
      12'h9B8: dout  = 8'b11111000; // 2488 : 248 - 0xf8 -- plane 1
      12'h9B9: dout  = 8'b11010000; // 2489 : 208 - 0xd0
      12'h9BA: dout  = 8'b00110000; // 2490 :  48 - 0x30
      12'h9BB: dout  = 8'b01100000; // 2491 :  96 - 0x60
      12'h9BC: dout  = 8'b10000000; // 2492 : 128 - 0x80
      12'h9BD: dout  = 8'b00000000; // 2493 :   0 - 0x0
      12'h9BE: dout  = 8'b00000000; // 2494 :   0 - 0x0
      12'h9BF: dout  = 8'b00000000; // 2495 :   0 - 0x0
      12'h9C0: dout  = 8'b00000001; // 2496 :   1 - 0x1 -- Sprite 0x9c
      12'h9C1: dout  = 8'b00000000; // 2497 :   0 - 0x0
      12'h9C2: dout  = 8'b00000000; // 2498 :   0 - 0x0
      12'h9C3: dout  = 8'b00000000; // 2499 :   0 - 0x0
      12'h9C4: dout  = 8'b00000001; // 2500 :   1 - 0x1
      12'h9C5: dout  = 8'b00000001; // 2501 :   1 - 0x1
      12'h9C6: dout  = 8'b00000010; // 2502 :   2 - 0x2
      12'h9C7: dout  = 8'b00000110; // 2503 :   6 - 0x6
      12'h9C8: dout  = 8'b00000000; // 2504 :   0 - 0x0 -- plane 1
      12'h9C9: dout  = 8'b00000001; // 2505 :   1 - 0x1
      12'h9CA: dout  = 8'b00000000; // 2506 :   0 - 0x0
      12'h9CB: dout  = 8'b00000000; // 2507 :   0 - 0x0
      12'h9CC: dout  = 8'b00000000; // 2508 :   0 - 0x0
      12'h9CD: dout  = 8'b00000000; // 2509 :   0 - 0x0
      12'h9CE: dout  = 8'b00000001; // 2510 :   1 - 0x1
      12'h9CF: dout  = 8'b00000011; // 2511 :   3 - 0x3
      12'h9D0: dout  = 8'b01111000; // 2512 : 120 - 0x78 -- Sprite 0x9d
      12'h9D1: dout  = 8'b00101010; // 2513 :  42 - 0x2a
      12'h9D2: dout  = 8'b01010100; // 2514 :  84 - 0x54
      12'h9D3: dout  = 8'b00101001; // 2515 :  41 - 0x29
      12'h9D4: dout  = 8'b00101111; // 2516 :  47 - 0x2f
      12'h9D5: dout  = 8'b00111100; // 2517 :  60 - 0x3c
      12'h9D6: dout  = 8'b00011110; // 2518 :  30 - 0x1e
      12'h9D7: dout  = 8'b00000000; // 2519 :   0 - 0x0
      12'h9D8: dout  = 8'b00000111; // 2520 :   7 - 0x7 -- plane 1
      12'h9D9: dout  = 8'b00010111; // 2521 :  23 - 0x17
      12'h9DA: dout  = 8'b00101111; // 2522 :  47 - 0x2f
      12'h9DB: dout  = 8'b00011110; // 2523 :  30 - 0x1e
      12'h9DC: dout  = 8'b00010000; // 2524 :  16 - 0x10
      12'h9DD: dout  = 8'b00000100; // 2525 :   4 - 0x4
      12'h9DE: dout  = 8'b00000000; // 2526 :   0 - 0x0
      12'h9DF: dout  = 8'b00000000; // 2527 :   0 - 0x0
      12'h9E0: dout  = 8'b10110000; // 2528 : 176 - 0xb0 -- Sprite 0x9e
      12'h9E1: dout  = 8'b11101000; // 2529 : 232 - 0xe8
      12'h9E2: dout  = 8'b10001100; // 2530 : 140 - 0x8c
      12'h9E3: dout  = 8'b10011110; // 2531 : 158 - 0x9e
      12'h9E4: dout  = 8'b00011111; // 2532 :  31 - 0x1f
      12'h9E5: dout  = 8'b00001111; // 2533 :  15 - 0xf
      12'h9E6: dout  = 8'b10010110; // 2534 : 150 - 0x96
      12'h9E7: dout  = 8'b00011100; // 2535 :  28 - 0x1c
      12'h9E8: dout  = 8'b00000000; // 2536 :   0 - 0x0 -- plane 1
      12'h9E9: dout  = 8'b00010000; // 2537 :  16 - 0x10
      12'h9EA: dout  = 8'b01111000; // 2538 : 120 - 0x78
      12'h9EB: dout  = 8'b01110100; // 2539 : 116 - 0x74
      12'h9EC: dout  = 8'b11111110; // 2540 : 254 - 0xfe
      12'h9ED: dout  = 8'b11111000; // 2541 : 248 - 0xf8
      12'h9EE: dout  = 8'b11111100; // 2542 : 252 - 0xfc
      12'h9EF: dout  = 8'b11111000; // 2543 : 248 - 0xf8
      12'h9F0: dout  = 8'b00001100; // 2544 :  12 - 0xc -- Sprite 0x9f
      12'h9F1: dout  = 8'b00111000; // 2545 :  56 - 0x38
      12'h9F2: dout  = 8'b11101000; // 2546 : 232 - 0xe8
      12'h9F3: dout  = 8'b11110000; // 2547 : 240 - 0xf0
      12'h9F4: dout  = 8'b11000000; // 2548 : 192 - 0xc0
      12'h9F5: dout  = 8'b01110000; // 2549 : 112 - 0x70
      12'h9F6: dout  = 8'b11000000; // 2550 : 192 - 0xc0
      12'h9F7: dout  = 8'b00000000; // 2551 :   0 - 0x0
      12'h9F8: dout  = 8'b11111000; // 2552 : 248 - 0xf8 -- plane 1
      12'h9F9: dout  = 8'b11010000; // 2553 : 208 - 0xd0
      12'h9FA: dout  = 8'b00110000; // 2554 :  48 - 0x30
      12'h9FB: dout  = 8'b11000000; // 2555 : 192 - 0xc0
      12'h9FC: dout  = 8'b00000000; // 2556 :   0 - 0x0
      12'h9FD: dout  = 8'b00000000; // 2557 :   0 - 0x0
      12'h9FE: dout  = 8'b00000000; // 2558 :   0 - 0x0
      12'h9FF: dout  = 8'b00000000; // 2559 :   0 - 0x0
      12'hA00: dout  = 8'b00000011; // 2560 :   3 - 0x3 -- Sprite 0xa0
      12'hA01: dout  = 8'b00001111; // 2561 :  15 - 0xf
      12'hA02: dout  = 8'b00011100; // 2562 :  28 - 0x1c
      12'hA03: dout  = 8'b00110000; // 2563 :  48 - 0x30
      12'hA04: dout  = 8'b01100000; // 2564 :  96 - 0x60
      12'hA05: dout  = 8'b01100000; // 2565 :  96 - 0x60
      12'hA06: dout  = 8'b11000000; // 2566 : 192 - 0xc0
      12'hA07: dout  = 8'b11000000; // 2567 : 192 - 0xc0
      12'hA08: dout  = 8'b00000000; // 2568 :   0 - 0x0 -- plane 1
      12'hA09: dout  = 8'b00000011; // 2569 :   3 - 0x3
      12'hA0A: dout  = 8'b00001111; // 2570 :  15 - 0xf
      12'hA0B: dout  = 8'b00011111; // 2571 :  31 - 0x1f
      12'hA0C: dout  = 8'b00111111; // 2572 :  63 - 0x3f
      12'hA0D: dout  = 8'b00111111; // 2573 :  63 - 0x3f
      12'hA0E: dout  = 8'b01111111; // 2574 : 127 - 0x7f
      12'hA0F: dout  = 8'b01111111; // 2575 : 127 - 0x7f
      12'hA10: dout  = 8'b11000000; // 2576 : 192 - 0xc0 -- Sprite 0xa1
      12'hA11: dout  = 8'b11000000; // 2577 : 192 - 0xc0
      12'hA12: dout  = 8'b01100000; // 2578 :  96 - 0x60
      12'hA13: dout  = 8'b01100000; // 2579 :  96 - 0x60
      12'hA14: dout  = 8'b00110000; // 2580 :  48 - 0x30
      12'hA15: dout  = 8'b00011010; // 2581 :  26 - 0x1a
      12'hA16: dout  = 8'b00001101; // 2582 :  13 - 0xd
      12'hA17: dout  = 8'b00000011; // 2583 :   3 - 0x3
      12'hA18: dout  = 8'b01111111; // 2584 : 127 - 0x7f -- plane 1
      12'hA19: dout  = 8'b01111111; // 2585 : 127 - 0x7f
      12'hA1A: dout  = 8'b00111111; // 2586 :  63 - 0x3f
      12'hA1B: dout  = 8'b00111111; // 2587 :  63 - 0x3f
      12'hA1C: dout  = 8'b00011111; // 2588 :  31 - 0x1f
      12'hA1D: dout  = 8'b00000101; // 2589 :   5 - 0x5
      12'hA1E: dout  = 8'b00000010; // 2590 :   2 - 0x2
      12'hA1F: dout  = 8'b00000000; // 2591 :   0 - 0x0
      12'hA20: dout  = 8'b11000000; // 2592 : 192 - 0xc0 -- Sprite 0xa2
      12'hA21: dout  = 8'b11110000; // 2593 : 240 - 0xf0
      12'hA22: dout  = 8'b00111000; // 2594 :  56 - 0x38
      12'hA23: dout  = 8'b00001100; // 2595 :  12 - 0xc
      12'hA24: dout  = 8'b00000110; // 2596 :   6 - 0x6
      12'hA25: dout  = 8'b00000010; // 2597 :   2 - 0x2
      12'hA26: dout  = 8'b00000101; // 2598 :   5 - 0x5
      12'hA27: dout  = 8'b00000011; // 2599 :   3 - 0x3
      12'hA28: dout  = 8'b00000000; // 2600 :   0 - 0x0 -- plane 1
      12'hA29: dout  = 8'b11000000; // 2601 : 192 - 0xc0
      12'hA2A: dout  = 8'b11110000; // 2602 : 240 - 0xf0
      12'hA2B: dout  = 8'b11111000; // 2603 : 248 - 0xf8
      12'hA2C: dout  = 8'b11111000; // 2604 : 248 - 0xf8
      12'hA2D: dout  = 8'b11111100; // 2605 : 252 - 0xfc
      12'hA2E: dout  = 8'b11111010; // 2606 : 250 - 0xfa
      12'hA2F: dout  = 8'b11111100; // 2607 : 252 - 0xfc
      12'hA30: dout  = 8'b00000101; // 2608 :   5 - 0x5 -- Sprite 0xa3
      12'hA31: dout  = 8'b00001011; // 2609 :  11 - 0xb
      12'hA32: dout  = 8'b00010110; // 2610 :  22 - 0x16
      12'hA33: dout  = 8'b00101010; // 2611 :  42 - 0x2a
      12'hA34: dout  = 8'b01010100; // 2612 :  84 - 0x54
      12'hA35: dout  = 8'b10101000; // 2613 : 168 - 0xa8
      12'hA36: dout  = 8'b01110000; // 2614 : 112 - 0x70
      12'hA37: dout  = 8'b11000000; // 2615 : 192 - 0xc0
      12'hA38: dout  = 8'b11111010; // 2616 : 250 - 0xfa -- plane 1
      12'hA39: dout  = 8'b11110100; // 2617 : 244 - 0xf4
      12'hA3A: dout  = 8'b11101000; // 2618 : 232 - 0xe8
      12'hA3B: dout  = 8'b11010100; // 2619 : 212 - 0xd4
      12'hA3C: dout  = 8'b10101000; // 2620 : 168 - 0xa8
      12'hA3D: dout  = 8'b01010000; // 2621 :  80 - 0x50
      12'hA3E: dout  = 8'b10000000; // 2622 : 128 - 0x80
      12'hA3F: dout  = 8'b00000000; // 2623 :   0 - 0x0
      12'hA40: dout  = 8'b00000000; // 2624 :   0 - 0x0 -- Sprite 0xa4
      12'hA41: dout  = 8'b00001111; // 2625 :  15 - 0xf
      12'hA42: dout  = 8'b00011111; // 2626 :  31 - 0x1f
      12'hA43: dout  = 8'b00110001; // 2627 :  49 - 0x31
      12'hA44: dout  = 8'b00111111; // 2628 :  63 - 0x3f
      12'hA45: dout  = 8'b01111111; // 2629 : 127 - 0x7f
      12'hA46: dout  = 8'b11111111; // 2630 : 255 - 0xff
      12'hA47: dout  = 8'b11011111; // 2631 : 223 - 0xdf
      12'hA48: dout  = 8'b00000000; // 2632 :   0 - 0x0 -- plane 1
      12'hA49: dout  = 8'b00000000; // 2633 :   0 - 0x0
      12'hA4A: dout  = 8'b00000000; // 2634 :   0 - 0x0
      12'hA4B: dout  = 8'b00001110; // 2635 :  14 - 0xe
      12'hA4C: dout  = 8'b00000000; // 2636 :   0 - 0x0
      12'hA4D: dout  = 8'b00001010; // 2637 :  10 - 0xa
      12'hA4E: dout  = 8'b01001010; // 2638 :  74 - 0x4a
      12'hA4F: dout  = 8'b01100000; // 2639 :  96 - 0x60
      12'hA50: dout  = 8'b11000000; // 2640 : 192 - 0xc0 -- Sprite 0xa5
      12'hA51: dout  = 8'b11000111; // 2641 : 199 - 0xc7
      12'hA52: dout  = 8'b01101111; // 2642 : 111 - 0x6f
      12'hA53: dout  = 8'b01100111; // 2643 : 103 - 0x67
      12'hA54: dout  = 8'b01100011; // 2644 :  99 - 0x63
      12'hA55: dout  = 8'b00110000; // 2645 :  48 - 0x30
      12'hA56: dout  = 8'b00011000; // 2646 :  24 - 0x18
      12'hA57: dout  = 8'b00000111; // 2647 :   7 - 0x7
      12'hA58: dout  = 8'b01111111; // 2648 : 127 - 0x7f -- plane 1
      12'hA59: dout  = 8'b01111000; // 2649 : 120 - 0x78
      12'hA5A: dout  = 8'b00110111; // 2650 :  55 - 0x37
      12'hA5B: dout  = 8'b00111011; // 2651 :  59 - 0x3b
      12'hA5C: dout  = 8'b00111100; // 2652 :  60 - 0x3c
      12'hA5D: dout  = 8'b00011111; // 2653 :  31 - 0x1f
      12'hA5E: dout  = 8'b00000111; // 2654 :   7 - 0x7
      12'hA5F: dout  = 8'b00000000; // 2655 :   0 - 0x0
      12'hA60: dout  = 8'b00000000; // 2656 :   0 - 0x0 -- Sprite 0xa6
      12'hA61: dout  = 8'b11110000; // 2657 : 240 - 0xf0
      12'hA62: dout  = 8'b11111000; // 2658 : 248 - 0xf8
      12'hA63: dout  = 8'b10001100; // 2659 : 140 - 0x8c
      12'hA64: dout  = 8'b11111100; // 2660 : 252 - 0xfc
      12'hA65: dout  = 8'b11111110; // 2661 : 254 - 0xfe
      12'hA66: dout  = 8'b11111101; // 2662 : 253 - 0xfd
      12'hA67: dout  = 8'b11111001; // 2663 : 249 - 0xf9
      12'hA68: dout  = 8'b00000000; // 2664 :   0 - 0x0 -- plane 1
      12'hA69: dout  = 8'b00000000; // 2665 :   0 - 0x0
      12'hA6A: dout  = 8'b00000000; // 2666 :   0 - 0x0
      12'hA6B: dout  = 8'b01110000; // 2667 : 112 - 0x70
      12'hA6C: dout  = 8'b00000000; // 2668 :   0 - 0x0
      12'hA6D: dout  = 8'b01010000; // 2669 :  80 - 0x50
      12'hA6E: dout  = 8'b01010010; // 2670 :  82 - 0x52
      12'hA6F: dout  = 8'b00000110; // 2671 :   6 - 0x6
      12'hA70: dout  = 8'b00000011; // 2672 :   3 - 0x3 -- Sprite 0xa7
      12'hA71: dout  = 8'b11100101; // 2673 : 229 - 0xe5
      12'hA72: dout  = 8'b11110010; // 2674 : 242 - 0xf2
      12'hA73: dout  = 8'b11100110; // 2675 : 230 - 0xe6
      12'hA74: dout  = 8'b11001010; // 2676 : 202 - 0xca
      12'hA75: dout  = 8'b00010100; // 2677 :  20 - 0x14
      12'hA76: dout  = 8'b00111000; // 2678 :  56 - 0x38
      12'hA77: dout  = 8'b11100000; // 2679 : 224 - 0xe0
      12'hA78: dout  = 8'b11111100; // 2680 : 252 - 0xfc -- plane 1
      12'hA79: dout  = 8'b00011010; // 2681 :  26 - 0x1a
      12'hA7A: dout  = 8'b11101100; // 2682 : 236 - 0xec
      12'hA7B: dout  = 8'b11011000; // 2683 : 216 - 0xd8
      12'hA7C: dout  = 8'b00110100; // 2684 :  52 - 0x34
      12'hA7D: dout  = 8'b11101000; // 2685 : 232 - 0xe8
      12'hA7E: dout  = 8'b11000000; // 2686 : 192 - 0xc0
      12'hA7F: dout  = 8'b00000000; // 2687 :   0 - 0x0
      12'hA80: dout  = 8'b00000000; // 2688 :   0 - 0x0 -- Sprite 0xa8
      12'hA81: dout  = 8'b00001111; // 2689 :  15 - 0xf
      12'hA82: dout  = 8'b00011111; // 2690 :  31 - 0x1f
      12'hA83: dout  = 8'b00110001; // 2691 :  49 - 0x31
      12'hA84: dout  = 8'b00111111; // 2692 :  63 - 0x3f
      12'hA85: dout  = 8'b01111111; // 2693 : 127 - 0x7f
      12'hA86: dout  = 8'b11111111; // 2694 : 255 - 0xff
      12'hA87: dout  = 8'b11011111; // 2695 : 223 - 0xdf
      12'hA88: dout  = 8'b00000000; // 2696 :   0 - 0x0 -- plane 1
      12'hA89: dout  = 8'b00000000; // 2697 :   0 - 0x0
      12'hA8A: dout  = 8'b00000000; // 2698 :   0 - 0x0
      12'hA8B: dout  = 8'b00001110; // 2699 :  14 - 0xe
      12'hA8C: dout  = 8'b00000000; // 2700 :   0 - 0x0
      12'hA8D: dout  = 8'b00001110; // 2701 :  14 - 0xe
      12'hA8E: dout  = 8'b01001010; // 2702 :  74 - 0x4a
      12'hA8F: dout  = 8'b01100000; // 2703 :  96 - 0x60
      12'hA90: dout  = 8'b11000000; // 2704 : 192 - 0xc0 -- Sprite 0xa9
      12'hA91: dout  = 8'b11000011; // 2705 : 195 - 0xc3
      12'hA92: dout  = 8'b11000111; // 2706 : 199 - 0xc7
      12'hA93: dout  = 8'b11001111; // 2707 : 207 - 0xcf
      12'hA94: dout  = 8'b11000111; // 2708 : 199 - 0xc7
      12'hA95: dout  = 8'b11000000; // 2709 : 192 - 0xc0
      12'hA96: dout  = 8'b11100000; // 2710 : 224 - 0xe0
      12'hA97: dout  = 8'b11111111; // 2711 : 255 - 0xff
      12'hA98: dout  = 8'b01111111; // 2712 : 127 - 0x7f -- plane 1
      12'hA99: dout  = 8'b01111100; // 2713 : 124 - 0x7c
      12'hA9A: dout  = 8'b01111011; // 2714 : 123 - 0x7b
      12'hA9B: dout  = 8'b01110111; // 2715 : 119 - 0x77
      12'hA9C: dout  = 8'b01111000; // 2716 : 120 - 0x78
      12'hA9D: dout  = 8'b01111111; // 2717 : 127 - 0x7f
      12'hA9E: dout  = 8'b01111111; // 2718 : 127 - 0x7f
      12'hA9F: dout  = 8'b00000000; // 2719 :   0 - 0x0
      12'hAA0: dout  = 8'b00000000; // 2720 :   0 - 0x0 -- Sprite 0xaa
      12'hAA1: dout  = 8'b11110000; // 2721 : 240 - 0xf0
      12'hAA2: dout  = 8'b11111000; // 2722 : 248 - 0xf8
      12'hAA3: dout  = 8'b10001100; // 2723 : 140 - 0x8c
      12'hAA4: dout  = 8'b11111100; // 2724 : 252 - 0xfc
      12'hAA5: dout  = 8'b11111110; // 2725 : 254 - 0xfe
      12'hAA6: dout  = 8'b11111101; // 2726 : 253 - 0xfd
      12'hAA7: dout  = 8'b11111001; // 2727 : 249 - 0xf9
      12'hAA8: dout  = 8'b00000000; // 2728 :   0 - 0x0 -- plane 1
      12'hAA9: dout  = 8'b00000000; // 2729 :   0 - 0x0
      12'hAAA: dout  = 8'b00000000; // 2730 :   0 - 0x0
      12'hAAB: dout  = 8'b01110000; // 2731 : 112 - 0x70
      12'hAAC: dout  = 8'b00000000; // 2732 :   0 - 0x0
      12'hAAD: dout  = 8'b01110000; // 2733 : 112 - 0x70
      12'hAAE: dout  = 8'b01010010; // 2734 :  82 - 0x52
      12'hAAF: dout  = 8'b00000110; // 2735 :   6 - 0x6
      12'hAB0: dout  = 8'b00000011; // 2736 :   3 - 0x3 -- Sprite 0xab
      12'hAB1: dout  = 8'b11000101; // 2737 : 197 - 0xc5
      12'hAB2: dout  = 8'b11100011; // 2738 : 227 - 0xe3
      12'hAB3: dout  = 8'b11110101; // 2739 : 245 - 0xf5
      12'hAB4: dout  = 8'b11100011; // 2740 : 227 - 0xe3
      12'hAB5: dout  = 8'b00000101; // 2741 :   5 - 0x5
      12'hAB6: dout  = 8'b00001011; // 2742 :  11 - 0xb
      12'hAB7: dout  = 8'b11111111; // 2743 : 255 - 0xff
      12'hAB8: dout  = 8'b11111100; // 2744 : 252 - 0xfc -- plane 1
      12'hAB9: dout  = 8'b00111010; // 2745 :  58 - 0x3a
      12'hABA: dout  = 8'b11011100; // 2746 : 220 - 0xdc
      12'hABB: dout  = 8'b11101010; // 2747 : 234 - 0xea
      12'hABC: dout  = 8'b00011100; // 2748 :  28 - 0x1c
      12'hABD: dout  = 8'b11111010; // 2749 : 250 - 0xfa
      12'hABE: dout  = 8'b11110100; // 2750 : 244 - 0xf4
      12'hABF: dout  = 8'b00000000; // 2751 :   0 - 0x0
      12'hAC0: dout  = 8'b10000011; // 2752 : 131 - 0x83 -- Sprite 0xac
      12'hAC1: dout  = 8'b10001100; // 2753 : 140 - 0x8c
      12'hAC2: dout  = 8'b10010000; // 2754 : 144 - 0x90
      12'hAC3: dout  = 8'b10010000; // 2755 : 144 - 0x90
      12'hAC4: dout  = 8'b11100000; // 2756 : 224 - 0xe0
      12'hAC5: dout  = 8'b10100000; // 2757 : 160 - 0xa0
      12'hAC6: dout  = 8'b10101111; // 2758 : 175 - 0xaf
      12'hAC7: dout  = 8'b01101111; // 2759 : 111 - 0x6f
      12'hAC8: dout  = 8'b00000000; // 2760 :   0 - 0x0 -- plane 1
      12'hAC9: dout  = 8'b00000011; // 2761 :   3 - 0x3
      12'hACA: dout  = 8'b00001111; // 2762 :  15 - 0xf
      12'hACB: dout  = 8'b00001111; // 2763 :  15 - 0xf
      12'hACC: dout  = 8'b00011111; // 2764 :  31 - 0x1f
      12'hACD: dout  = 8'b01011111; // 2765 :  95 - 0x5f
      12'hACE: dout  = 8'b01010000; // 2766 :  80 - 0x50
      12'hACF: dout  = 8'b00010000; // 2767 :  16 - 0x10
      12'hAD0: dout  = 8'b11111011; // 2768 : 251 - 0xfb -- Sprite 0xad
      12'hAD1: dout  = 8'b00000101; // 2769 :   5 - 0x5
      12'hAD2: dout  = 8'b00000101; // 2770 :   5 - 0x5
      12'hAD3: dout  = 8'b00000101; // 2771 :   5 - 0x5
      12'hAD4: dout  = 8'b01000101; // 2772 :  69 - 0x45
      12'hAD5: dout  = 8'b01100101; // 2773 : 101 - 0x65
      12'hAD6: dout  = 8'b11110101; // 2774 : 245 - 0xf5
      12'hAD7: dout  = 8'b11111101; // 2775 : 253 - 0xfd
      12'hAD8: dout  = 8'b00000000; // 2776 :   0 - 0x0 -- plane 1
      12'hAD9: dout  = 8'b11111010; // 2777 : 250 - 0xfa
      12'hADA: dout  = 8'b11111010; // 2778 : 250 - 0xfa
      12'hADB: dout  = 8'b11111010; // 2779 : 250 - 0xfa
      12'hADC: dout  = 8'b10111010; // 2780 : 186 - 0xba
      12'hADD: dout  = 8'b10011010; // 2781 : 154 - 0x9a
      12'hADE: dout  = 8'b00001010; // 2782 :  10 - 0xa
      12'hADF: dout  = 8'b00000010; // 2783 :   2 - 0x2
      12'hAE0: dout  = 8'b10000011; // 2784 : 131 - 0x83 -- Sprite 0xae
      12'hAE1: dout  = 8'b10001100; // 2785 : 140 - 0x8c
      12'hAE2: dout  = 8'b10010000; // 2786 : 144 - 0x90
      12'hAE3: dout  = 8'b10010000; // 2787 : 144 - 0x90
      12'hAE4: dout  = 8'b11100000; // 2788 : 224 - 0xe0
      12'hAE5: dout  = 8'b10100000; // 2789 : 160 - 0xa0
      12'hAE6: dout  = 8'b10101111; // 2790 : 175 - 0xaf
      12'hAE7: dout  = 8'b01101111; // 2791 : 111 - 0x6f
      12'hAE8: dout  = 8'b00000000; // 2792 :   0 - 0x0 -- plane 1
      12'hAE9: dout  = 8'b00000011; // 2793 :   3 - 0x3
      12'hAEA: dout  = 8'b00001111; // 2794 :  15 - 0xf
      12'hAEB: dout  = 8'b00001111; // 2795 :  15 - 0xf
      12'hAEC: dout  = 8'b00011111; // 2796 :  31 - 0x1f
      12'hAED: dout  = 8'b01011111; // 2797 :  95 - 0x5f
      12'hAEE: dout  = 8'b01010000; // 2798 :  80 - 0x50
      12'hAEF: dout  = 8'b00010111; // 2799 :  23 - 0x17
      12'hAF0: dout  = 8'b11111011; // 2800 : 251 - 0xfb -- Sprite 0xaf
      12'hAF1: dout  = 8'b00000101; // 2801 :   5 - 0x5
      12'hAF2: dout  = 8'b00000101; // 2802 :   5 - 0x5
      12'hAF3: dout  = 8'b00000101; // 2803 :   5 - 0x5
      12'hAF4: dout  = 8'b11000101; // 2804 : 197 - 0xc5
      12'hAF5: dout  = 8'b11100101; // 2805 : 229 - 0xe5
      12'hAF6: dout  = 8'b11110101; // 2806 : 245 - 0xf5
      12'hAF7: dout  = 8'b11111101; // 2807 : 253 - 0xfd
      12'hAF8: dout  = 8'b00000000; // 2808 :   0 - 0x0 -- plane 1
      12'hAF9: dout  = 8'b11111010; // 2809 : 250 - 0xfa
      12'hAFA: dout  = 8'b11111010; // 2810 : 250 - 0xfa
      12'hAFB: dout  = 8'b11111010; // 2811 : 250 - 0xfa
      12'hAFC: dout  = 8'b00111010; // 2812 :  58 - 0x3a
      12'hAFD: dout  = 8'b01011010; // 2813 :  90 - 0x5a
      12'hAFE: dout  = 8'b01101010; // 2814 : 106 - 0x6a
      12'hAFF: dout  = 8'b11110010; // 2815 : 242 - 0xf2
      12'hB00: dout  = 8'b00000000; // 2816 :   0 - 0x0 -- Sprite 0xb0
      12'hB01: dout  = 8'b00000011; // 2817 :   3 - 0x3
      12'hB02: dout  = 8'b00001111; // 2818 :  15 - 0xf
      12'hB03: dout  = 8'b00111111; // 2819 :  63 - 0x3f
      12'hB04: dout  = 8'b01111111; // 2820 : 127 - 0x7f
      12'hB05: dout  = 8'b01111111; // 2821 : 127 - 0x7f
      12'hB06: dout  = 8'b11111111; // 2822 : 255 - 0xff
      12'hB07: dout  = 8'b11111111; // 2823 : 255 - 0xff
      12'hB08: dout  = 8'b00000000; // 2824 :   0 - 0x0 -- plane 1
      12'hB09: dout  = 8'b00000000; // 2825 :   0 - 0x0
      12'hB0A: dout  = 8'b00000011; // 2826 :   3 - 0x3
      12'hB0B: dout  = 8'b00001111; // 2827 :  15 - 0xf
      12'hB0C: dout  = 8'b00111011; // 2828 :  59 - 0x3b
      12'hB0D: dout  = 8'b00111111; // 2829 :  63 - 0x3f
      12'hB0E: dout  = 8'b01101111; // 2830 : 111 - 0x6f
      12'hB0F: dout  = 8'b01111101; // 2831 : 125 - 0x7d
      12'hB10: dout  = 8'b11111111; // 2832 : 255 - 0xff -- Sprite 0xb1
      12'hB11: dout  = 8'b10001111; // 2833 : 143 - 0x8f
      12'hB12: dout  = 8'b10000000; // 2834 : 128 - 0x80
      12'hB13: dout  = 8'b11110000; // 2835 : 240 - 0xf0
      12'hB14: dout  = 8'b11111111; // 2836 : 255 - 0xff
      12'hB15: dout  = 8'b11111111; // 2837 : 255 - 0xff
      12'hB16: dout  = 8'b01111111; // 2838 : 127 - 0x7f
      12'hB17: dout  = 8'b00001111; // 2839 :  15 - 0xf
      12'hB18: dout  = 8'b00001111; // 2840 :  15 - 0xf -- plane 1
      12'hB19: dout  = 8'b01110000; // 2841 : 112 - 0x70
      12'hB1A: dout  = 8'b01111111; // 2842 : 127 - 0x7f
      12'hB1B: dout  = 8'b00001111; // 2843 :  15 - 0xf
      12'hB1C: dout  = 8'b01110000; // 2844 : 112 - 0x70
      12'hB1D: dout  = 8'b01111111; // 2845 : 127 - 0x7f
      12'hB1E: dout  = 8'b00001111; // 2846 :  15 - 0xf
      12'hB1F: dout  = 8'b00000000; // 2847 :   0 - 0x0
      12'hB20: dout  = 8'b00000000; // 2848 :   0 - 0x0 -- Sprite 0xb2
      12'hB21: dout  = 8'b11000000; // 2849 : 192 - 0xc0
      12'hB22: dout  = 8'b11110000; // 2850 : 240 - 0xf0
      12'hB23: dout  = 8'b11111100; // 2851 : 252 - 0xfc
      12'hB24: dout  = 8'b11111110; // 2852 : 254 - 0xfe
      12'hB25: dout  = 8'b11111110; // 2853 : 254 - 0xfe
      12'hB26: dout  = 8'b11111111; // 2854 : 255 - 0xff
      12'hB27: dout  = 8'b11111111; // 2855 : 255 - 0xff
      12'hB28: dout  = 8'b00000000; // 2856 :   0 - 0x0 -- plane 1
      12'hB29: dout  = 8'b00000000; // 2857 :   0 - 0x0
      12'hB2A: dout  = 8'b11000000; // 2858 : 192 - 0xc0
      12'hB2B: dout  = 8'b11110000; // 2859 : 240 - 0xf0
      12'hB2C: dout  = 8'b10111100; // 2860 : 188 - 0xbc
      12'hB2D: dout  = 8'b11110100; // 2861 : 244 - 0xf4
      12'hB2E: dout  = 8'b11111110; // 2862 : 254 - 0xfe
      12'hB2F: dout  = 8'b11011110; // 2863 : 222 - 0xde
      12'hB30: dout  = 8'b11111111; // 2864 : 255 - 0xff -- Sprite 0xb3
      12'hB31: dout  = 8'b11110001; // 2865 : 241 - 0xf1
      12'hB32: dout  = 8'b00000001; // 2866 :   1 - 0x1
      12'hB33: dout  = 8'b00001111; // 2867 :  15 - 0xf
      12'hB34: dout  = 8'b11111111; // 2868 : 255 - 0xff
      12'hB35: dout  = 8'b11111111; // 2869 : 255 - 0xff
      12'hB36: dout  = 8'b11111110; // 2870 : 254 - 0xfe
      12'hB37: dout  = 8'b11110000; // 2871 : 240 - 0xf0
      12'hB38: dout  = 8'b11110000; // 2872 : 240 - 0xf0 -- plane 1
      12'hB39: dout  = 8'b00001110; // 2873 :  14 - 0xe
      12'hB3A: dout  = 8'b11111110; // 2874 : 254 - 0xfe
      12'hB3B: dout  = 8'b11110000; // 2875 : 240 - 0xf0
      12'hB3C: dout  = 8'b00001110; // 2876 :  14 - 0xe
      12'hB3D: dout  = 8'b11111110; // 2877 : 254 - 0xfe
      12'hB3E: dout  = 8'b11110000; // 2878 : 240 - 0xf0
      12'hB3F: dout  = 8'b00000000; // 2879 :   0 - 0x0
      12'hB40: dout  = 8'b00000000; // 2880 :   0 - 0x0 -- Sprite 0xb4
      12'hB41: dout  = 8'b00000011; // 2881 :   3 - 0x3
      12'hB42: dout  = 8'b00001110; // 2882 :  14 - 0xe
      12'hB43: dout  = 8'b00110101; // 2883 :  53 - 0x35
      12'hB44: dout  = 8'b01101110; // 2884 : 110 - 0x6e
      12'hB45: dout  = 8'b01010101; // 2885 :  85 - 0x55
      12'hB46: dout  = 8'b10111010; // 2886 : 186 - 0xba
      12'hB47: dout  = 8'b11010111; // 2887 : 215 - 0xd7
      12'hB48: dout  = 8'b00000000; // 2888 :   0 - 0x0 -- plane 1
      12'hB49: dout  = 8'b00000000; // 2889 :   0 - 0x0
      12'hB4A: dout  = 8'b00000011; // 2890 :   3 - 0x3
      12'hB4B: dout  = 8'b00001111; // 2891 :  15 - 0xf
      12'hB4C: dout  = 8'b00111011; // 2892 :  59 - 0x3b
      12'hB4D: dout  = 8'b00111111; // 2893 :  63 - 0x3f
      12'hB4E: dout  = 8'b01101111; // 2894 : 111 - 0x6f
      12'hB4F: dout  = 8'b01111101; // 2895 : 125 - 0x7d
      12'hB50: dout  = 8'b11111010; // 2896 : 250 - 0xfa -- Sprite 0xb5
      12'hB51: dout  = 8'b10001111; // 2897 : 143 - 0x8f
      12'hB52: dout  = 8'b10000000; // 2898 : 128 - 0x80
      12'hB53: dout  = 8'b11110000; // 2899 : 240 - 0xf0
      12'hB54: dout  = 8'b10101111; // 2900 : 175 - 0xaf
      12'hB55: dout  = 8'b11010101; // 2901 : 213 - 0xd5
      12'hB56: dout  = 8'b01111010; // 2902 : 122 - 0x7a
      12'hB57: dout  = 8'b00001111; // 2903 :  15 - 0xf
      12'hB58: dout  = 8'b00001111; // 2904 :  15 - 0xf -- plane 1
      12'hB59: dout  = 8'b01110000; // 2905 : 112 - 0x70
      12'hB5A: dout  = 8'b01111111; // 2906 : 127 - 0x7f
      12'hB5B: dout  = 8'b00001111; // 2907 :  15 - 0xf
      12'hB5C: dout  = 8'b01110000; // 2908 : 112 - 0x70
      12'hB5D: dout  = 8'b01111111; // 2909 : 127 - 0x7f
      12'hB5E: dout  = 8'b00001111; // 2910 :  15 - 0xf
      12'hB5F: dout  = 8'b00000000; // 2911 :   0 - 0x0
      12'hB60: dout  = 8'b00000000; // 2912 :   0 - 0x0 -- Sprite 0xb6
      12'hB61: dout  = 8'b11000000; // 2913 : 192 - 0xc0
      12'hB62: dout  = 8'b10110000; // 2914 : 176 - 0xb0
      12'hB63: dout  = 8'b01011100; // 2915 :  92 - 0x5c
      12'hB64: dout  = 8'b11101010; // 2916 : 234 - 0xea
      12'hB65: dout  = 8'b01011110; // 2917 :  94 - 0x5e
      12'hB66: dout  = 8'b10101011; // 2918 : 171 - 0xab
      12'hB67: dout  = 8'b01110101; // 2919 : 117 - 0x75
      12'hB68: dout  = 8'b00000000; // 2920 :   0 - 0x0 -- plane 1
      12'hB69: dout  = 8'b00000000; // 2921 :   0 - 0x0
      12'hB6A: dout  = 8'b11000000; // 2922 : 192 - 0xc0
      12'hB6B: dout  = 8'b11110000; // 2923 : 240 - 0xf0
      12'hB6C: dout  = 8'b10111100; // 2924 : 188 - 0xbc
      12'hB6D: dout  = 8'b11110100; // 2925 : 244 - 0xf4
      12'hB6E: dout  = 8'b11111110; // 2926 : 254 - 0xfe
      12'hB6F: dout  = 8'b11011110; // 2927 : 222 - 0xde
      12'hB70: dout  = 8'b10101111; // 2928 : 175 - 0xaf -- Sprite 0xb7
      12'hB71: dout  = 8'b11110001; // 2929 : 241 - 0xf1
      12'hB72: dout  = 8'b00000001; // 2930 :   1 - 0x1
      12'hB73: dout  = 8'b00001111; // 2931 :  15 - 0xf
      12'hB74: dout  = 8'b11111011; // 2932 : 251 - 0xfb
      12'hB75: dout  = 8'b01010101; // 2933 :  85 - 0x55
      12'hB76: dout  = 8'b10101110; // 2934 : 174 - 0xae
      12'hB77: dout  = 8'b11110000; // 2935 : 240 - 0xf0
      12'hB78: dout  = 8'b11110000; // 2936 : 240 - 0xf0 -- plane 1
      12'hB79: dout  = 8'b00001110; // 2937 :  14 - 0xe
      12'hB7A: dout  = 8'b11111110; // 2938 : 254 - 0xfe
      12'hB7B: dout  = 8'b11110000; // 2939 : 240 - 0xf0
      12'hB7C: dout  = 8'b00001110; // 2940 :  14 - 0xe
      12'hB7D: dout  = 8'b11111110; // 2941 : 254 - 0xfe
      12'hB7E: dout  = 8'b11110000; // 2942 : 240 - 0xf0
      12'hB7F: dout  = 8'b00000000; // 2943 :   0 - 0x0
      12'hB80: dout  = 8'b00000000; // 2944 :   0 - 0x0 -- Sprite 0xb8
      12'hB81: dout  = 8'b00000011; // 2945 :   3 - 0x3
      12'hB82: dout  = 8'b00001100; // 2946 :  12 - 0xc
      12'hB83: dout  = 8'b00110000; // 2947 :  48 - 0x30
      12'hB84: dout  = 8'b01000100; // 2948 :  68 - 0x44
      12'hB85: dout  = 8'b01000000; // 2949 :  64 - 0x40
      12'hB86: dout  = 8'b10010000; // 2950 : 144 - 0x90
      12'hB87: dout  = 8'b10000010; // 2951 : 130 - 0x82
      12'hB88: dout  = 8'b00000000; // 2952 :   0 - 0x0 -- plane 1
      12'hB89: dout  = 8'b00000000; // 2953 :   0 - 0x0
      12'hB8A: dout  = 8'b00000011; // 2954 :   3 - 0x3
      12'hB8B: dout  = 8'b00001111; // 2955 :  15 - 0xf
      12'hB8C: dout  = 8'b00111011; // 2956 :  59 - 0x3b
      12'hB8D: dout  = 8'b00111111; // 2957 :  63 - 0x3f
      12'hB8E: dout  = 8'b01101111; // 2958 : 111 - 0x6f
      12'hB8F: dout  = 8'b01111101; // 2959 : 125 - 0x7d
      12'hB90: dout  = 8'b11110000; // 2960 : 240 - 0xf0 -- Sprite 0xb9
      12'hB91: dout  = 8'b11111111; // 2961 : 255 - 0xff
      12'hB92: dout  = 8'b11111111; // 2962 : 255 - 0xff
      12'hB93: dout  = 8'b11111111; // 2963 : 255 - 0xff
      12'hB94: dout  = 8'b10001111; // 2964 : 143 - 0x8f
      12'hB95: dout  = 8'b10000000; // 2965 : 128 - 0x80
      12'hB96: dout  = 8'b01110000; // 2966 : 112 - 0x70
      12'hB97: dout  = 8'b00001111; // 2967 :  15 - 0xf
      12'hB98: dout  = 8'b00001111; // 2968 :  15 - 0xf -- plane 1
      12'hB99: dout  = 8'b00100000; // 2969 :  32 - 0x20
      12'hB9A: dout  = 8'b01010101; // 2970 :  85 - 0x55
      12'hB9B: dout  = 8'b00001010; // 2971 :  10 - 0xa
      12'hB9C: dout  = 8'b01110000; // 2972 : 112 - 0x70
      12'hB9D: dout  = 8'b01111111; // 2973 : 127 - 0x7f
      12'hB9E: dout  = 8'b00001111; // 2974 :  15 - 0xf
      12'hB9F: dout  = 8'b00000000; // 2975 :   0 - 0x0
      12'hBA0: dout  = 8'b00000000; // 2976 :   0 - 0x0 -- Sprite 0xba
      12'hBA1: dout  = 8'b11000000; // 2977 : 192 - 0xc0
      12'hBA2: dout  = 8'b00110000; // 2978 :  48 - 0x30
      12'hBA3: dout  = 8'b00001100; // 2979 :  12 - 0xc
      12'hBA4: dout  = 8'b01000010; // 2980 :  66 - 0x42
      12'hBA5: dout  = 8'b00001010; // 2981 :  10 - 0xa
      12'hBA6: dout  = 8'b00000001; // 2982 :   1 - 0x1
      12'hBA7: dout  = 8'b00100001; // 2983 :  33 - 0x21
      12'hBA8: dout  = 8'b00000000; // 2984 :   0 - 0x0 -- plane 1
      12'hBA9: dout  = 8'b00000000; // 2985 :   0 - 0x0
      12'hBAA: dout  = 8'b11000000; // 2986 : 192 - 0xc0
      12'hBAB: dout  = 8'b11110000; // 2987 : 240 - 0xf0
      12'hBAC: dout  = 8'b10111100; // 2988 : 188 - 0xbc
      12'hBAD: dout  = 8'b11110100; // 2989 : 244 - 0xf4
      12'hBAE: dout  = 8'b11111110; // 2990 : 254 - 0xfe
      12'hBAF: dout  = 8'b11011110; // 2991 : 222 - 0xde
      12'hBB0: dout  = 8'b00001111; // 2992 :  15 - 0xf -- Sprite 0xbb
      12'hBB1: dout  = 8'b11111111; // 2993 : 255 - 0xff
      12'hBB2: dout  = 8'b11111111; // 2994 : 255 - 0xff
      12'hBB3: dout  = 8'b11111111; // 2995 : 255 - 0xff
      12'hBB4: dout  = 8'b11110001; // 2996 : 241 - 0xf1
      12'hBB5: dout  = 8'b00000001; // 2997 :   1 - 0x1
      12'hBB6: dout  = 8'b00001110; // 2998 :  14 - 0xe
      12'hBB7: dout  = 8'b11110000; // 2999 : 240 - 0xf0
      12'hBB8: dout  = 8'b11110000; // 3000 : 240 - 0xf0 -- plane 1
      12'hBB9: dout  = 8'b00001010; // 3001 :  10 - 0xa
      12'hBBA: dout  = 8'b01010100; // 3002 :  84 - 0x54
      12'hBBB: dout  = 8'b10100000; // 3003 : 160 - 0xa0
      12'hBBC: dout  = 8'b00001110; // 3004 :  14 - 0xe
      12'hBBD: dout  = 8'b11111110; // 3005 : 254 - 0xfe
      12'hBBE: dout  = 8'b11110000; // 3006 : 240 - 0xf0
      12'hBBF: dout  = 8'b00000000; // 3007 :   0 - 0x0
      12'hBC0: dout  = 8'b11110011; // 3008 : 243 - 0xf3 -- Sprite 0xbc
      12'hBC1: dout  = 8'b11111111; // 3009 : 255 - 0xff
      12'hBC2: dout  = 8'b11000100; // 3010 : 196 - 0xc4
      12'hBC3: dout  = 8'b11000000; // 3011 : 192 - 0xc0
      12'hBC4: dout  = 8'b01000000; // 3012 :  64 - 0x40
      12'hBC5: dout  = 8'b01100011; // 3013 :  99 - 0x63
      12'hBC6: dout  = 8'b11000111; // 3014 : 199 - 0xc7
      12'hBC7: dout  = 8'b11000110; // 3015 : 198 - 0xc6
      12'hBC8: dout  = 8'b00000000; // 3016 :   0 - 0x0 -- plane 1
      12'hBC9: dout  = 8'b01110011; // 3017 : 115 - 0x73
      12'hBCA: dout  = 8'b01111011; // 3018 : 123 - 0x7b
      12'hBCB: dout  = 8'b01111111; // 3019 : 127 - 0x7f
      12'hBCC: dout  = 8'b00111111; // 3020 :  63 - 0x3f
      12'hBCD: dout  = 8'b00011100; // 3021 :  28 - 0x1c
      12'hBCE: dout  = 8'b01111011; // 3022 : 123 - 0x7b
      12'hBCF: dout  = 8'b01111011; // 3023 : 123 - 0x7b
      12'hBD0: dout  = 8'b11000110; // 3024 : 198 - 0xc6 -- Sprite 0xbd
      12'hBD1: dout  = 8'b11000110; // 3025 : 198 - 0xc6
      12'hBD2: dout  = 8'b01100011; // 3026 :  99 - 0x63
      12'hBD3: dout  = 8'b01000000; // 3027 :  64 - 0x40
      12'hBD4: dout  = 8'b11000000; // 3028 : 192 - 0xc0
      12'hBD5: dout  = 8'b11000100; // 3029 : 196 - 0xc4
      12'hBD6: dout  = 8'b11001100; // 3030 : 204 - 0xcc
      12'hBD7: dout  = 8'b11110011; // 3031 : 243 - 0xf3
      12'hBD8: dout  = 8'b01111011; // 3032 : 123 - 0x7b -- plane 1
      12'hBD9: dout  = 8'b01111011; // 3033 : 123 - 0x7b
      12'hBDA: dout  = 8'b00011100; // 3034 :  28 - 0x1c
      12'hBDB: dout  = 8'b00111111; // 3035 :  63 - 0x3f
      12'hBDC: dout  = 8'b01111111; // 3036 : 127 - 0x7f
      12'hBDD: dout  = 8'b01111011; // 3037 : 123 - 0x7b
      12'hBDE: dout  = 8'b01110011; // 3038 : 115 - 0x73
      12'hBDF: dout  = 8'b00000000; // 3039 :   0 - 0x0
      12'hBE0: dout  = 8'b11001111; // 3040 : 207 - 0xcf -- Sprite 0xbe
      12'hBE1: dout  = 8'b11111111; // 3041 : 255 - 0xff
      12'hBE2: dout  = 8'b00100001; // 3042 :  33 - 0x21
      12'hBE3: dout  = 8'b00000001; // 3043 :   1 - 0x1
      12'hBE4: dout  = 8'b00000010; // 3044 :   2 - 0x2
      12'hBE5: dout  = 8'b11000110; // 3045 : 198 - 0xc6
      12'hBE6: dout  = 8'b11100001; // 3046 : 225 - 0xe1
      12'hBE7: dout  = 8'b00100001; // 3047 :  33 - 0x21
      12'hBE8: dout  = 8'b00000000; // 3048 :   0 - 0x0 -- plane 1
      12'hBE9: dout  = 8'b11001110; // 3049 : 206 - 0xce
      12'hBEA: dout  = 8'b11011110; // 3050 : 222 - 0xde
      12'hBEB: dout  = 8'b11111110; // 3051 : 254 - 0xfe
      12'hBEC: dout  = 8'b11111100; // 3052 : 252 - 0xfc
      12'hBED: dout  = 8'b00111000; // 3053 :  56 - 0x38
      12'hBEE: dout  = 8'b11011110; // 3054 : 222 - 0xde
      12'hBEF: dout  = 8'b11011110; // 3055 : 222 - 0xde
      12'hBF0: dout  = 8'b00100001; // 3056 :  33 - 0x21 -- Sprite 0xbf
      12'hBF1: dout  = 8'b00100001; // 3057 :  33 - 0x21
      12'hBF2: dout  = 8'b11000110; // 3058 : 198 - 0xc6
      12'hBF3: dout  = 8'b00000010; // 3059 :   2 - 0x2
      12'hBF4: dout  = 8'b00000001; // 3060 :   1 - 0x1
      12'hBF5: dout  = 8'b00100001; // 3061 :  33 - 0x21
      12'hBF6: dout  = 8'b00110001; // 3062 :  49 - 0x31
      12'hBF7: dout  = 8'b11001111; // 3063 : 207 - 0xcf
      12'hBF8: dout  = 8'b11011110; // 3064 : 222 - 0xde -- plane 1
      12'hBF9: dout  = 8'b11011110; // 3065 : 222 - 0xde
      12'hBFA: dout  = 8'b00111000; // 3066 :  56 - 0x38
      12'hBFB: dout  = 8'b11111100; // 3067 : 252 - 0xfc
      12'hBFC: dout  = 8'b11111110; // 3068 : 254 - 0xfe
      12'hBFD: dout  = 8'b11011110; // 3069 : 222 - 0xde
      12'hBFE: dout  = 8'b11001110; // 3070 : 206 - 0xce
      12'hBFF: dout  = 8'b00000000; // 3071 :   0 - 0x0
      12'hC00: dout  = 8'b00000000; // 3072 :   0 - 0x0 -- Sprite 0xc0
      12'hC01: dout  = 8'b01010000; // 3073 :  80 - 0x50
      12'hC02: dout  = 8'b10110011; // 3074 : 179 - 0xb3
      12'hC03: dout  = 8'b10010111; // 3075 : 151 - 0x97
      12'hC04: dout  = 8'b10011111; // 3076 : 159 - 0x9f
      12'hC05: dout  = 8'b01101111; // 3077 : 111 - 0x6f
      12'hC06: dout  = 8'b00011111; // 3078 :  31 - 0x1f
      12'hC07: dout  = 8'b00011111; // 3079 :  31 - 0x1f
      12'hC08: dout  = 8'b00000000; // 3080 :   0 - 0x0 -- plane 1
      12'hC09: dout  = 8'b00000000; // 3081 :   0 - 0x0
      12'hC0A: dout  = 8'b01000000; // 3082 :  64 - 0x40
      12'hC0B: dout  = 8'b01100000; // 3083 :  96 - 0x60
      12'hC0C: dout  = 8'b01100001; // 3084 :  97 - 0x61
      12'hC0D: dout  = 8'b00000010; // 3085 :   2 - 0x2
      12'hC0E: dout  = 8'b00000010; // 3086 :   2 - 0x2
      12'hC0F: dout  = 8'b00000111; // 3087 :   7 - 0x7
      12'hC10: dout  = 8'b00011111; // 3088 :  31 - 0x1f -- Sprite 0xc1
      12'hC11: dout  = 8'b00011111; // 3089 :  31 - 0x1f
      12'hC12: dout  = 8'b00001111; // 3090 :  15 - 0xf
      12'hC13: dout  = 8'b00000111; // 3091 :   7 - 0x7
      12'hC14: dout  = 8'b00011101; // 3092 :  29 - 0x1d
      12'hC15: dout  = 8'b00101100; // 3093 :  44 - 0x2c
      12'hC16: dout  = 8'b01010100; // 3094 :  84 - 0x54
      12'hC17: dout  = 8'b01111100; // 3095 : 124 - 0x7c
      12'hC18: dout  = 8'b00000111; // 3096 :   7 - 0x7 -- plane 1
      12'hC19: dout  = 8'b00000100; // 3097 :   4 - 0x4
      12'hC1A: dout  = 8'b00000111; // 3098 :   7 - 0x7
      12'hC1B: dout  = 8'b00000001; // 3099 :   1 - 0x1
      12'hC1C: dout  = 8'b00000000; // 3100 :   0 - 0x0
      12'hC1D: dout  = 8'b00010000; // 3101 :  16 - 0x10
      12'hC1E: dout  = 8'b00101000; // 3102 :  40 - 0x28
      12'hC1F: dout  = 8'b00000000; // 3103 :   0 - 0x0
      12'hC20: dout  = 8'b00000000; // 3104 :   0 - 0x0 -- Sprite 0xc2
      12'hC21: dout  = 8'b00001010; // 3105 :  10 - 0xa
      12'hC22: dout  = 8'b11001101; // 3106 : 205 - 0xcd
      12'hC23: dout  = 8'b11101001; // 3107 : 233 - 0xe9
      12'hC24: dout  = 8'b11111001; // 3108 : 249 - 0xf9
      12'hC25: dout  = 8'b11110110; // 3109 : 246 - 0xf6
      12'hC26: dout  = 8'b11110000; // 3110 : 240 - 0xf0
      12'hC27: dout  = 8'b11111000; // 3111 : 248 - 0xf8
      12'hC28: dout  = 8'b00000000; // 3112 :   0 - 0x0 -- plane 1
      12'hC29: dout  = 8'b00000000; // 3113 :   0 - 0x0
      12'hC2A: dout  = 8'b00000010; // 3114 :   2 - 0x2
      12'hC2B: dout  = 8'b00000110; // 3115 :   6 - 0x6
      12'hC2C: dout  = 8'b11100110; // 3116 : 230 - 0xe6
      12'hC2D: dout  = 8'b10100000; // 3117 : 160 - 0xa0
      12'hC2E: dout  = 8'b10100000; // 3118 : 160 - 0xa0
      12'hC2F: dout  = 8'b11110000; // 3119 : 240 - 0xf0
      12'hC30: dout  = 8'b11111000; // 3120 : 248 - 0xf8 -- Sprite 0xc3
      12'hC31: dout  = 8'b11111000; // 3121 : 248 - 0xf8
      12'hC32: dout  = 8'b11110000; // 3122 : 240 - 0xf0
      12'hC33: dout  = 8'b11000000; // 3123 : 192 - 0xc0
      12'hC34: dout  = 8'b10111000; // 3124 : 184 - 0xb8
      12'hC35: dout  = 8'b00110100; // 3125 :  52 - 0x34
      12'hC36: dout  = 8'b00101010; // 3126 :  42 - 0x2a
      12'hC37: dout  = 8'b00111110; // 3127 :  62 - 0x3e
      12'hC38: dout  = 8'b11110000; // 3128 : 240 - 0xf0 -- plane 1
      12'hC39: dout  = 8'b00110000; // 3129 :  48 - 0x30
      12'hC3A: dout  = 8'b11000000; // 3130 : 192 - 0xc0
      12'hC3B: dout  = 8'b10000000; // 3131 : 128 - 0x80
      12'hC3C: dout  = 8'b00000000; // 3132 :   0 - 0x0
      12'hC3D: dout  = 8'b00001000; // 3133 :   8 - 0x8
      12'hC3E: dout  = 8'b00010100; // 3134 :  20 - 0x14
      12'hC3F: dout  = 8'b00000000; // 3135 :   0 - 0x0
      12'hC40: dout  = 8'b00000101; // 3136 :   5 - 0x5 -- Sprite 0xc4
      12'hC41: dout  = 8'b00001010; // 3137 :  10 - 0xa
      12'hC42: dout  = 8'b00001000; // 3138 :   8 - 0x8
      12'hC43: dout  = 8'b00001111; // 3139 :  15 - 0xf
      12'hC44: dout  = 8'b00000001; // 3140 :   1 - 0x1
      12'hC45: dout  = 8'b00000011; // 3141 :   3 - 0x3
      12'hC46: dout  = 8'b00000111; // 3142 :   7 - 0x7
      12'hC47: dout  = 8'b00001111; // 3143 :  15 - 0xf
      12'hC48: dout  = 8'b00000000; // 3144 :   0 - 0x0 -- plane 1
      12'hC49: dout  = 8'b00000101; // 3145 :   5 - 0x5
      12'hC4A: dout  = 8'b00000111; // 3146 :   7 - 0x7
      12'hC4B: dout  = 8'b00000000; // 3147 :   0 - 0x0
      12'hC4C: dout  = 8'b00000000; // 3148 :   0 - 0x0
      12'hC4D: dout  = 8'b00000000; // 3149 :   0 - 0x0
      12'hC4E: dout  = 8'b00000000; // 3150 :   0 - 0x0
      12'hC4F: dout  = 8'b00000001; // 3151 :   1 - 0x1
      12'hC50: dout  = 8'b00001111; // 3152 :  15 - 0xf -- Sprite 0xc5
      12'hC51: dout  = 8'b11101111; // 3153 : 239 - 0xef
      12'hC52: dout  = 8'b11011111; // 3154 : 223 - 0xdf
      12'hC53: dout  = 8'b10101111; // 3155 : 175 - 0xaf
      12'hC54: dout  = 8'b01100111; // 3156 : 103 - 0x67
      12'hC55: dout  = 8'b00001101; // 3157 :  13 - 0xd
      12'hC56: dout  = 8'b00001010; // 3158 :  10 - 0xa
      12'hC57: dout  = 8'b00000111; // 3159 :   7 - 0x7
      12'hC58: dout  = 8'b00000010; // 3160 :   2 - 0x2 -- plane 1
      12'hC59: dout  = 8'b00000111; // 3161 :   7 - 0x7
      12'hC5A: dout  = 8'b00100111; // 3162 :  39 - 0x27
      12'hC5B: dout  = 8'b01010011; // 3163 :  83 - 0x53
      12'hC5C: dout  = 8'b00000000; // 3164 :   0 - 0x0
      12'hC5D: dout  = 8'b00000010; // 3165 :   2 - 0x2
      12'hC5E: dout  = 8'b00000101; // 3166 :   5 - 0x5
      12'hC5F: dout  = 8'b00000000; // 3167 :   0 - 0x0
      12'hC60: dout  = 8'b00000000; // 3168 :   0 - 0x0 -- Sprite 0xc6
      12'hC61: dout  = 8'b10000000; // 3169 : 128 - 0x80
      12'hC62: dout  = 8'b10000000; // 3170 : 128 - 0x80
      12'hC63: dout  = 8'b11110000; // 3171 : 240 - 0xf0
      12'hC64: dout  = 8'b11111000; // 3172 : 248 - 0xf8
      12'hC65: dout  = 8'b11111100; // 3173 : 252 - 0xfc
      12'hC66: dout  = 8'b11111100; // 3174 : 252 - 0xfc
      12'hC67: dout  = 8'b11111100; // 3175 : 252 - 0xfc
      12'hC68: dout  = 8'b00000000; // 3176 :   0 - 0x0 -- plane 1
      12'hC69: dout  = 8'b00000000; // 3177 :   0 - 0x0
      12'hC6A: dout  = 8'b00000000; // 3178 :   0 - 0x0
      12'hC6B: dout  = 8'b00000000; // 3179 :   0 - 0x0
      12'hC6C: dout  = 8'b00000000; // 3180 :   0 - 0x0
      12'hC6D: dout  = 8'b01100000; // 3181 :  96 - 0x60
      12'hC6E: dout  = 8'b11011000; // 3182 : 216 - 0xd8
      12'hC6F: dout  = 8'b10110000; // 3183 : 176 - 0xb0
      12'hC70: dout  = 8'b11111100; // 3184 : 252 - 0xfc -- Sprite 0xc7
      12'hC71: dout  = 8'b11111110; // 3185 : 254 - 0xfe
      12'hC72: dout  = 8'b11111001; // 3186 : 249 - 0xf9
      12'hC73: dout  = 8'b11111010; // 3187 : 250 - 0xfa
      12'hC74: dout  = 8'b11101001; // 3188 : 233 - 0xe9
      12'hC75: dout  = 8'b00001110; // 3189 :  14 - 0xe
      12'hC76: dout  = 8'b10000000; // 3190 : 128 - 0x80
      12'hC77: dout  = 8'b00000000; // 3191 :   0 - 0x0
      12'hC78: dout  = 8'b11101000; // 3192 : 232 - 0xe8 -- plane 1
      12'hC79: dout  = 8'b01111000; // 3193 : 120 - 0x78
      12'hC7A: dout  = 8'b10110110; // 3194 : 182 - 0xb6
      12'hC7B: dout  = 8'b11100100; // 3195 : 228 - 0xe4
      12'hC7C: dout  = 8'b00000110; // 3196 :   6 - 0x6
      12'hC7D: dout  = 8'b00000000; // 3197 :   0 - 0x0
      12'hC7E: dout  = 8'b00000000; // 3198 :   0 - 0x0
      12'hC7F: dout  = 8'b00000000; // 3199 :   0 - 0x0
      12'hC80: dout  = 8'b00000000; // 3200 :   0 - 0x0 -- Sprite 0xc8
      12'hC81: dout  = 8'b11000000; // 3201 : 192 - 0xc0
      12'hC82: dout  = 8'b10100000; // 3202 : 160 - 0xa0
      12'hC83: dout  = 8'b11010011; // 3203 : 211 - 0xd3
      12'hC84: dout  = 8'b10110111; // 3204 : 183 - 0xb7
      12'hC85: dout  = 8'b11111111; // 3205 : 255 - 0xff
      12'hC86: dout  = 8'b00001111; // 3206 :  15 - 0xf
      12'hC87: dout  = 8'b00011111; // 3207 :  31 - 0x1f
      12'hC88: dout  = 8'b00000000; // 3208 :   0 - 0x0 -- plane 1
      12'hC89: dout  = 8'b00000000; // 3209 :   0 - 0x0
      12'hC8A: dout  = 8'b01000000; // 3210 :  64 - 0x40
      12'hC8B: dout  = 8'b00100000; // 3211 :  32 - 0x20
      12'hC8C: dout  = 8'b01000000; // 3212 :  64 - 0x40
      12'hC8D: dout  = 8'b00000111; // 3213 :   7 - 0x7
      12'hC8E: dout  = 8'b00000101; // 3214 :   5 - 0x5
      12'hC8F: dout  = 8'b00001101; // 3215 :  13 - 0xd
      12'hC90: dout  = 8'b00011111; // 3216 :  31 - 0x1f -- Sprite 0xc9
      12'hC91: dout  = 8'b00001111; // 3217 :  15 - 0xf
      12'hC92: dout  = 8'b11110111; // 3218 : 247 - 0xf7
      12'hC93: dout  = 8'b10110111; // 3219 : 183 - 0xb7
      12'hC94: dout  = 8'b11010011; // 3220 : 211 - 0xd3
      12'hC95: dout  = 8'b10100000; // 3221 : 160 - 0xa0
      12'hC96: dout  = 8'b11000000; // 3222 : 192 - 0xc0
      12'hC97: dout  = 8'b00000000; // 3223 :   0 - 0x0
      12'hC98: dout  = 8'b00001101; // 3224 :  13 - 0xd -- plane 1
      12'hC99: dout  = 8'b00000101; // 3225 :   5 - 0x5
      12'hC9A: dout  = 8'b00000011; // 3226 :   3 - 0x3
      12'hC9B: dout  = 8'b01000011; // 3227 :  67 - 0x43
      12'hC9C: dout  = 8'b00100000; // 3228 :  32 - 0x20
      12'hC9D: dout  = 8'b01000000; // 3229 :  64 - 0x40
      12'hC9E: dout  = 8'b00000000; // 3230 :   0 - 0x0
      12'hC9F: dout  = 8'b00000000; // 3231 :   0 - 0x0
      12'hCA0: dout  = 8'b00011100; // 3232 :  28 - 0x1c -- Sprite 0xca
      12'hCA1: dout  = 8'b00100010; // 3233 :  34 - 0x22
      12'hCA2: dout  = 8'b00100100; // 3234 :  36 - 0x24
      12'hCA3: dout  = 8'b11011110; // 3235 : 222 - 0xde
      12'hCA4: dout  = 8'b11110000; // 3236 : 240 - 0xf0
      12'hCA5: dout  = 8'b11111000; // 3237 : 248 - 0xf8
      12'hCA6: dout  = 8'b11111100; // 3238 : 252 - 0xfc
      12'hCA7: dout  = 8'b11111100; // 3239 : 252 - 0xfc
      12'hCA8: dout  = 8'b00000000; // 3240 :   0 - 0x0 -- plane 1
      12'hCA9: dout  = 8'b00011100; // 3241 :  28 - 0x1c
      12'hCAA: dout  = 8'b00011000; // 3242 :  24 - 0x18
      12'hCAB: dout  = 8'b00000000; // 3243 :   0 - 0x0
      12'hCAC: dout  = 8'b00000000; // 3244 :   0 - 0x0
      12'hCAD: dout  = 8'b10000000; // 3245 : 128 - 0x80
      12'hCAE: dout  = 8'b11100000; // 3246 : 224 - 0xe0
      12'hCAF: dout  = 8'b10010000; // 3247 : 144 - 0x90
      12'hCB0: dout  = 8'b11111100; // 3248 : 252 - 0xfc -- Sprite 0xcb
      12'hCB1: dout  = 8'b11111100; // 3249 : 252 - 0xfc
      12'hCB2: dout  = 8'b11111000; // 3250 : 248 - 0xf8
      12'hCB3: dout  = 8'b11110000; // 3251 : 240 - 0xf0
      12'hCB4: dout  = 8'b10011110; // 3252 : 158 - 0x9e
      12'hCB5: dout  = 8'b00100100; // 3253 :  36 - 0x24
      12'hCB6: dout  = 8'b00100010; // 3254 :  34 - 0x22
      12'hCB7: dout  = 8'b00011100; // 3255 :  28 - 0x1c
      12'hCB8: dout  = 8'b11110000; // 3256 : 240 - 0xf0 -- plane 1
      12'hCB9: dout  = 8'b10010000; // 3257 : 144 - 0x90
      12'hCBA: dout  = 8'b11110000; // 3258 : 240 - 0xf0
      12'hCBB: dout  = 8'b10000000; // 3259 : 128 - 0x80
      12'hCBC: dout  = 8'b00000000; // 3260 :   0 - 0x0
      12'hCBD: dout  = 8'b00011000; // 3261 :  24 - 0x18
      12'hCBE: dout  = 8'b00011100; // 3262 :  28 - 0x1c
      12'hCBF: dout  = 8'b00000000; // 3263 :   0 - 0x0
      12'hCC0: dout  = 8'b00001110; // 3264 :  14 - 0xe -- Sprite 0xcc
      12'hCC1: dout  = 8'b00010110; // 3265 :  22 - 0x16
      12'hCC2: dout  = 8'b00011010; // 3266 :  26 - 0x1a
      12'hCC3: dout  = 8'b00000100; // 3267 :   4 - 0x4
      12'hCC4: dout  = 8'b01101111; // 3268 : 111 - 0x6f
      12'hCC5: dout  = 8'b10111111; // 3269 : 191 - 0xbf
      12'hCC6: dout  = 8'b11011111; // 3270 : 223 - 0xdf
      12'hCC7: dout  = 8'b10111111; // 3271 : 191 - 0xbf
      12'hCC8: dout  = 8'b00000000; // 3272 :   0 - 0x0 -- plane 1
      12'hCC9: dout  = 8'b00001000; // 3273 :   8 - 0x8
      12'hCCA: dout  = 8'b00000100; // 3274 :   4 - 0x4
      12'hCCB: dout  = 8'b00001000; // 3275 :   8 - 0x8
      12'hCCC: dout  = 8'b00000000; // 3276 :   0 - 0x0
      12'hCCD: dout  = 8'b01000110; // 3277 :  70 - 0x46
      12'hCCE: dout  = 8'b00101111; // 3278 :  47 - 0x2f
      12'hCCF: dout  = 8'b01001110; // 3279 :  78 - 0x4e
      12'hCD0: dout  = 8'b01011111; // 3280 :  95 - 0x5f -- Sprite 0xcd
      12'hCD1: dout  = 8'b00011111; // 3281 :  31 - 0x1f
      12'hCD2: dout  = 8'b00011111; // 3282 :  31 - 0x1f
      12'hCD3: dout  = 8'b00001111; // 3283 :  15 - 0xf
      12'hCD4: dout  = 8'b00111111; // 3284 :  63 - 0x3f
      12'hCD5: dout  = 8'b00100011; // 3285 :  35 - 0x23
      12'hCD6: dout  = 8'b00101010; // 3286 :  42 - 0x2a
      12'hCD7: dout  = 8'b00010100; // 3287 :  20 - 0x14
      12'hCD8: dout  = 8'b00001101; // 3288 :  13 - 0xd -- plane 1
      12'hCD9: dout  = 8'b00001011; // 3289 :  11 - 0xb
      12'hCDA: dout  = 8'b00001111; // 3290 :  15 - 0xf
      12'hCDB: dout  = 8'b00000110; // 3291 :   6 - 0x6
      12'hCDC: dout  = 8'b00000011; // 3292 :   3 - 0x3
      12'hCDD: dout  = 8'b00011100; // 3293 :  28 - 0x1c
      12'hCDE: dout  = 8'b00010100; // 3294 :  20 - 0x14
      12'hCDF: dout  = 8'b00000000; // 3295 :   0 - 0x0
      12'hCE0: dout  = 8'b00000000; // 3296 :   0 - 0x0 -- Sprite 0xce
      12'hCE1: dout  = 8'b00000000; // 3297 :   0 - 0x0
      12'hCE2: dout  = 8'b00000000; // 3298 :   0 - 0x0
      12'hCE3: dout  = 8'b00000000; // 3299 :   0 - 0x0
      12'hCE4: dout  = 8'b10001110; // 3300 : 142 - 0x8e
      12'hCE5: dout  = 8'b11001001; // 3301 : 201 - 0xc9
      12'hCE6: dout  = 8'b11101010; // 3302 : 234 - 0xea
      12'hCE7: dout  = 8'b11111001; // 3303 : 249 - 0xf9
      12'hCE8: dout  = 8'b00000000; // 3304 :   0 - 0x0 -- plane 1
      12'hCE9: dout  = 8'b00000000; // 3305 :   0 - 0x0
      12'hCEA: dout  = 8'b00000000; // 3306 :   0 - 0x0
      12'hCEB: dout  = 8'b00000000; // 3307 :   0 - 0x0
      12'hCEC: dout  = 8'b00000000; // 3308 :   0 - 0x0
      12'hCED: dout  = 8'b00000110; // 3309 :   6 - 0x6
      12'hCEE: dout  = 8'b00000100; // 3310 :   4 - 0x4
      12'hCEF: dout  = 8'b10000110; // 3311 : 134 - 0x86
      12'hCF0: dout  = 8'b11111110; // 3312 : 254 - 0xfe -- Sprite 0xcf
      12'hCF1: dout  = 8'b11111000; // 3313 : 248 - 0xf8
      12'hCF2: dout  = 8'b11111000; // 3314 : 248 - 0xf8
      12'hCF3: dout  = 8'b11111000; // 3315 : 248 - 0xf8
      12'hCF4: dout  = 8'b11110000; // 3316 : 240 - 0xf0
      12'hCF5: dout  = 8'b11100000; // 3317 : 224 - 0xe0
      12'hCF6: dout  = 8'b00000000; // 3318 :   0 - 0x0
      12'hCF7: dout  = 8'b00000000; // 3319 :   0 - 0x0
      12'hCF8: dout  = 8'b11000000; // 3320 : 192 - 0xc0 -- plane 1
      12'hCF9: dout  = 8'b01100000; // 3321 :  96 - 0x60
      12'hCFA: dout  = 8'b10100000; // 3322 : 160 - 0xa0
      12'hCFB: dout  = 8'b11000000; // 3323 : 192 - 0xc0
      12'hCFC: dout  = 8'b01000000; // 3324 :  64 - 0x40
      12'hCFD: dout  = 8'b00000000; // 3325 :   0 - 0x0
      12'hCFE: dout  = 8'b00000000; // 3326 :   0 - 0x0
      12'hCFF: dout  = 8'b00000000; // 3327 :   0 - 0x0
      12'hD00: dout  = 8'b00000000; // 3328 :   0 - 0x0 -- Sprite 0xd0
      12'hD01: dout  = 8'b00000000; // 3329 :   0 - 0x0
      12'hD02: dout  = 8'b00000100; // 3330 :   4 - 0x4
      12'hD03: dout  = 8'b00100110; // 3331 :  38 - 0x26
      12'hD04: dout  = 8'b00101011; // 3332 :  43 - 0x2b
      12'hD05: dout  = 8'b01110001; // 3333 : 113 - 0x71
      12'hD06: dout  = 8'b01000000; // 3334 :  64 - 0x40
      12'hD07: dout  = 8'b01000111; // 3335 :  71 - 0x47
      12'hD08: dout  = 8'b00000000; // 3336 :   0 - 0x0 -- plane 1
      12'hD09: dout  = 8'b00000000; // 3337 :   0 - 0x0
      12'hD0A: dout  = 8'b00000000; // 3338 :   0 - 0x0
      12'hD0B: dout  = 8'b00000000; // 3339 :   0 - 0x0
      12'hD0C: dout  = 8'b00000100; // 3340 :   4 - 0x4
      12'hD0D: dout  = 8'b00001110; // 3341 :  14 - 0xe
      12'hD0E: dout  = 8'b00111111; // 3342 :  63 - 0x3f
      12'hD0F: dout  = 8'b00111001; // 3343 :  57 - 0x39
      12'hD10: dout  = 8'b10001111; // 3344 : 143 - 0x8f -- Sprite 0xd1
      12'hD11: dout  = 8'b10001111; // 3345 : 143 - 0x8f
      12'hD12: dout  = 8'b01001111; // 3346 :  79 - 0x4f
      12'hD13: dout  = 8'b01001111; // 3347 :  79 - 0x4f
      12'hD14: dout  = 8'b00111111; // 3348 :  63 - 0x3f
      12'hD15: dout  = 8'b00010011; // 3349 :  19 - 0x13
      12'hD16: dout  = 8'b00010001; // 3350 :  17 - 0x11
      12'hD17: dout  = 8'b00011111; // 3351 :  31 - 0x1f
      12'hD18: dout  = 8'b01110000; // 3352 : 112 - 0x70 -- plane 1
      12'hD19: dout  = 8'b01111000; // 3353 : 120 - 0x78
      12'hD1A: dout  = 8'b00111111; // 3354 :  63 - 0x3f
      12'hD1B: dout  = 8'b00111111; // 3355 :  63 - 0x3f
      12'hD1C: dout  = 8'b00000011; // 3356 :   3 - 0x3
      12'hD1D: dout  = 8'b00001100; // 3357 :  12 - 0xc
      12'hD1E: dout  = 8'b00001110; // 3358 :  14 - 0xe
      12'hD1F: dout  = 8'b00000000; // 3359 :   0 - 0x0
      12'hD20: dout  = 8'b00000000; // 3360 :   0 - 0x0 -- Sprite 0xd2
      12'hD21: dout  = 8'b10000000; // 3361 : 128 - 0x80
      12'hD22: dout  = 8'b11001000; // 3362 : 200 - 0xc8
      12'hD23: dout  = 8'b11010100; // 3363 : 212 - 0xd4
      12'hD24: dout  = 8'b00100100; // 3364 :  36 - 0x24
      12'hD25: dout  = 8'b00000010; // 3365 :   2 - 0x2
      12'hD26: dout  = 8'b00000010; // 3366 :   2 - 0x2
      12'hD27: dout  = 8'b11110010; // 3367 : 242 - 0xf2
      12'hD28: dout  = 8'b00000000; // 3368 :   0 - 0x0 -- plane 1
      12'hD29: dout  = 8'b00000000; // 3369 :   0 - 0x0
      12'hD2A: dout  = 8'b00000000; // 3370 :   0 - 0x0
      12'hD2B: dout  = 8'b00001000; // 3371 :   8 - 0x8
      12'hD2C: dout  = 8'b11011000; // 3372 : 216 - 0xd8
      12'hD2D: dout  = 8'b11111100; // 3373 : 252 - 0xfc
      12'hD2E: dout  = 8'b11111100; // 3374 : 252 - 0xfc
      12'hD2F: dout  = 8'b10011100; // 3375 : 156 - 0x9c
      12'hD30: dout  = 8'b11110010; // 3376 : 242 - 0xf2 -- Sprite 0xd3
      12'hD31: dout  = 8'b11110010; // 3377 : 242 - 0xf2
      12'hD32: dout  = 8'b11110100; // 3378 : 244 - 0xf4
      12'hD33: dout  = 8'b11110100; // 3379 : 244 - 0xf4
      12'hD34: dout  = 8'b11110100; // 3380 : 244 - 0xf4
      12'hD35: dout  = 8'b11001000; // 3381 : 200 - 0xc8
      12'hD36: dout  = 8'b01000100; // 3382 :  68 - 0x44
      12'hD37: dout  = 8'b01111100; // 3383 : 124 - 0x7c
      12'hD38: dout  = 8'b00001100; // 3384 :  12 - 0xc -- plane 1
      12'hD39: dout  = 8'b10011100; // 3385 : 156 - 0x9c
      12'hD3A: dout  = 8'b11111000; // 3386 : 248 - 0xf8
      12'hD3B: dout  = 8'b01111000; // 3387 : 120 - 0x78
      12'hD3C: dout  = 8'b10001000; // 3388 : 136 - 0x88
      12'hD3D: dout  = 8'b00110000; // 3389 :  48 - 0x30
      12'hD3E: dout  = 8'b00111000; // 3390 :  56 - 0x38
      12'hD3F: dout  = 8'b00000000; // 3391 :   0 - 0x0
      12'hD40: dout  = 8'b00000000; // 3392 :   0 - 0x0 -- Sprite 0xd4
      12'hD41: dout  = 8'b00000000; // 3393 :   0 - 0x0
      12'hD42: dout  = 8'b00000000; // 3394 :   0 - 0x0
      12'hD43: dout  = 8'b00001001; // 3395 :   9 - 0x9
      12'hD44: dout  = 8'b00011010; // 3396 :  26 - 0x1a
      12'hD45: dout  = 8'b00010100; // 3397 :  20 - 0x14
      12'hD46: dout  = 8'b00100000; // 3398 :  32 - 0x20
      12'hD47: dout  = 8'b01000111; // 3399 :  71 - 0x47
      12'hD48: dout  = 8'b00000000; // 3400 :   0 - 0x0 -- plane 1
      12'hD49: dout  = 8'b00000000; // 3401 :   0 - 0x0
      12'hD4A: dout  = 8'b00000000; // 3402 :   0 - 0x0
      12'hD4B: dout  = 8'b00000000; // 3403 :   0 - 0x0
      12'hD4C: dout  = 8'b00000001; // 3404 :   1 - 0x1
      12'hD4D: dout  = 8'b00001011; // 3405 :  11 - 0xb
      12'hD4E: dout  = 8'b00011111; // 3406 :  31 - 0x1f
      12'hD4F: dout  = 8'b00111001; // 3407 :  57 - 0x39
      12'hD50: dout  = 8'b10001111; // 3408 : 143 - 0x8f -- Sprite 0xd5
      12'hD51: dout  = 8'b10001111; // 3409 : 143 - 0x8f
      12'hD52: dout  = 8'b01001111; // 3410 :  79 - 0x4f
      12'hD53: dout  = 8'b01001111; // 3411 :  79 - 0x4f
      12'hD54: dout  = 8'b00111111; // 3412 :  63 - 0x3f
      12'hD55: dout  = 8'b01000111; // 3413 :  71 - 0x47
      12'hD56: dout  = 8'b00100010; // 3414 :  34 - 0x22
      12'hD57: dout  = 8'b00011100; // 3415 :  28 - 0x1c
      12'hD58: dout  = 8'b01110000; // 3416 : 112 - 0x70 -- plane 1
      12'hD59: dout  = 8'b01111000; // 3417 : 120 - 0x78
      12'hD5A: dout  = 8'b00111111; // 3418 :  63 - 0x3f
      12'hD5B: dout  = 8'b00111111; // 3419 :  63 - 0x3f
      12'hD5C: dout  = 8'b00000011; // 3420 :   3 - 0x3
      12'hD5D: dout  = 8'b00111000; // 3421 :  56 - 0x38
      12'hD5E: dout  = 8'b00011100; // 3422 :  28 - 0x1c
      12'hD5F: dout  = 8'b00000000; // 3423 :   0 - 0x0
      12'hD60: dout  = 8'b00000000; // 3424 :   0 - 0x0 -- Sprite 0xd6
      12'hD61: dout  = 8'b01000000; // 3425 :  64 - 0x40
      12'hD62: dout  = 8'b11000000; // 3426 : 192 - 0xc0
      12'hD63: dout  = 8'b00101100; // 3427 :  44 - 0x2c
      12'hD64: dout  = 8'b00110100; // 3428 :  52 - 0x34
      12'hD65: dout  = 8'b00000100; // 3429 :   4 - 0x4
      12'hD66: dout  = 8'b00000010; // 3430 :   2 - 0x2
      12'hD67: dout  = 8'b11110010; // 3431 : 242 - 0xf2
      12'hD68: dout  = 8'b00000000; // 3432 :   0 - 0x0 -- plane 1
      12'hD69: dout  = 8'b00000000; // 3433 :   0 - 0x0
      12'hD6A: dout  = 8'b00000000; // 3434 :   0 - 0x0
      12'hD6B: dout  = 8'b11000000; // 3435 : 192 - 0xc0
      12'hD6C: dout  = 8'b11001000; // 3436 : 200 - 0xc8
      12'hD6D: dout  = 8'b11111000; // 3437 : 248 - 0xf8
      12'hD6E: dout  = 8'b11111100; // 3438 : 252 - 0xfc
      12'hD6F: dout  = 8'b10011100; // 3439 : 156 - 0x9c
      12'hD70: dout  = 8'b11110010; // 3440 : 242 - 0xf2 -- Sprite 0xd7
      12'hD71: dout  = 8'b11110010; // 3441 : 242 - 0xf2
      12'hD72: dout  = 8'b11110100; // 3442 : 244 - 0xf4
      12'hD73: dout  = 8'b11110111; // 3443 : 247 - 0xf7
      12'hD74: dout  = 8'b11111101; // 3444 : 253 - 0xfd
      12'hD75: dout  = 8'b11100001; // 3445 : 225 - 0xe1
      12'hD76: dout  = 8'b00010010; // 3446 :  18 - 0x12
      12'hD77: dout  = 8'b00001100; // 3447 :  12 - 0xc
      12'hD78: dout  = 8'b00001100; // 3448 :  12 - 0xc -- plane 1
      12'hD79: dout  = 8'b10011100; // 3449 : 156 - 0x9c
      12'hD7A: dout  = 8'b11111000; // 3450 : 248 - 0xf8
      12'hD7B: dout  = 8'b01111000; // 3451 : 120 - 0x78
      12'hD7C: dout  = 8'b11100010; // 3452 : 226 - 0xe2
      12'hD7D: dout  = 8'b00011110; // 3453 :  30 - 0x1e
      12'hD7E: dout  = 8'b00001100; // 3454 :  12 - 0xc
      12'hD7F: dout  = 8'b00000000; // 3455 :   0 - 0x0
      12'hD80: dout  = 8'b01111000; // 3456 : 120 - 0x78 -- Sprite 0xd8
      12'hD81: dout  = 8'b01001110; // 3457 :  78 - 0x4e
      12'hD82: dout  = 8'b11000010; // 3458 : 194 - 0xc2
      12'hD83: dout  = 8'b10011010; // 3459 : 154 - 0x9a
      12'hD84: dout  = 8'b10011011; // 3460 : 155 - 0x9b
      12'hD85: dout  = 8'b11011001; // 3461 : 217 - 0xd9
      12'hD86: dout  = 8'b01100011; // 3462 :  99 - 0x63
      12'hD87: dout  = 8'b00111110; // 3463 :  62 - 0x3e
      12'hD88: dout  = 8'b00000000; // 3464 :   0 - 0x0 -- plane 1
      12'hD89: dout  = 8'b00110000; // 3465 :  48 - 0x30
      12'hD8A: dout  = 8'b00111100; // 3466 :  60 - 0x3c
      12'hD8B: dout  = 8'b01111100; // 3467 : 124 - 0x7c
      12'hD8C: dout  = 8'b01111100; // 3468 : 124 - 0x7c
      12'hD8D: dout  = 8'b00111110; // 3469 :  62 - 0x3e
      12'hD8E: dout  = 8'b00011100; // 3470 :  28 - 0x1c
      12'hD8F: dout  = 8'b00000000; // 3471 :   0 - 0x0
      12'hD90: dout  = 8'b00011110; // 3472 :  30 - 0x1e -- Sprite 0xd9
      12'hD91: dout  = 8'b01110001; // 3473 : 113 - 0x71
      12'hD92: dout  = 8'b01001001; // 3474 :  73 - 0x49
      12'hD93: dout  = 8'b10111001; // 3475 : 185 - 0xb9
      12'hD94: dout  = 8'b10011101; // 3476 : 157 - 0x9d
      12'hD95: dout  = 8'b01010010; // 3477 :  82 - 0x52
      12'hD96: dout  = 8'b01110010; // 3478 : 114 - 0x72
      12'hD97: dout  = 8'b00011110; // 3479 :  30 - 0x1e
      12'hD98: dout  = 8'b00000000; // 3480 :   0 - 0x0 -- plane 1
      12'hD99: dout  = 8'b00001110; // 3481 :  14 - 0xe
      12'hD9A: dout  = 8'b00111110; // 3482 :  62 - 0x3e
      12'hD9B: dout  = 8'b01111110; // 3483 : 126 - 0x7e
      12'hD9C: dout  = 8'b01111110; // 3484 : 126 - 0x7e
      12'hD9D: dout  = 8'b00111100; // 3485 :  60 - 0x3c
      12'hD9E: dout  = 8'b00001100; // 3486 :  12 - 0xc
      12'hD9F: dout  = 8'b00000000; // 3487 :   0 - 0x0
      12'hDA0: dout  = 8'b01100000; // 3488 :  96 - 0x60 -- Sprite 0xda
      12'hDA1: dout  = 8'b01011110; // 3489 :  94 - 0x5e
      12'hDA2: dout  = 8'b10001001; // 3490 : 137 - 0x89
      12'hDA3: dout  = 8'b10111101; // 3491 : 189 - 0xbd
      12'hDA4: dout  = 8'b10011101; // 3492 : 157 - 0x9d
      12'hDA5: dout  = 8'b11010011; // 3493 : 211 - 0xd3
      12'hDA6: dout  = 8'b01000110; // 3494 :  70 - 0x46
      12'hDA7: dout  = 8'b01111100; // 3495 : 124 - 0x7c
      12'hDA8: dout  = 8'b00000000; // 3496 :   0 - 0x0 -- plane 1
      12'hDA9: dout  = 8'b00100000; // 3497 :  32 - 0x20
      12'hDAA: dout  = 8'b01111110; // 3498 : 126 - 0x7e
      12'hDAB: dout  = 8'b01111110; // 3499 : 126 - 0x7e
      12'hDAC: dout  = 8'b01111110; // 3500 : 126 - 0x7e
      12'hDAD: dout  = 8'b00111100; // 3501 :  60 - 0x3c
      12'hDAE: dout  = 8'b00111000; // 3502 :  56 - 0x38
      12'hDAF: dout  = 8'b00000000; // 3503 :   0 - 0x0
      12'hDB0: dout  = 8'b00011110; // 3504 :  30 - 0x1e -- Sprite 0xdb
      12'hDB1: dout  = 8'b00100011; // 3505 :  35 - 0x23
      12'hDB2: dout  = 8'b01001001; // 3506 :  73 - 0x49
      12'hDB3: dout  = 8'b10111101; // 3507 : 189 - 0xbd
      12'hDB4: dout  = 8'b10011001; // 3508 : 153 - 0x99
      12'hDB5: dout  = 8'b01000011; // 3509 :  67 - 0x43
      12'hDB6: dout  = 8'b01101110; // 3510 : 110 - 0x6e
      12'hDB7: dout  = 8'b00011000; // 3511 :  24 - 0x18
      12'hDB8: dout  = 8'b00000000; // 3512 :   0 - 0x0 -- plane 1
      12'hDB9: dout  = 8'b00011100; // 3513 :  28 - 0x1c
      12'hDBA: dout  = 8'b00111110; // 3514 :  62 - 0x3e
      12'hDBB: dout  = 8'b01111110; // 3515 : 126 - 0x7e
      12'hDBC: dout  = 8'b01111110; // 3516 : 126 - 0x7e
      12'hDBD: dout  = 8'b00111100; // 3517 :  60 - 0x3c
      12'hDBE: dout  = 8'b00010000; // 3518 :  16 - 0x10
      12'hDBF: dout  = 8'b00000000; // 3519 :   0 - 0x0
      12'hDC0: dout  = 8'b00000000; // 3520 :   0 - 0x0 -- Sprite 0xdc
      12'hDC1: dout  = 8'b00000000; // 3521 :   0 - 0x0
      12'hDC2: dout  = 8'b00000001; // 3522 :   1 - 0x1
      12'hDC3: dout  = 8'b00000010; // 3523 :   2 - 0x2
      12'hDC4: dout  = 8'b00000100; // 3524 :   4 - 0x4
      12'hDC5: dout  = 8'b00000010; // 3525 :   2 - 0x2
      12'hDC6: dout  = 8'b00011110; // 3526 :  30 - 0x1e
      12'hDC7: dout  = 8'b00010000; // 3527 :  16 - 0x10
      12'hDC8: dout  = 8'b00000000; // 3528 :   0 - 0x0 -- plane 1
      12'hDC9: dout  = 8'b00000000; // 3529 :   0 - 0x0
      12'hDCA: dout  = 8'b00000000; // 3530 :   0 - 0x0
      12'hDCB: dout  = 8'b00000001; // 3531 :   1 - 0x1
      12'hDCC: dout  = 8'b00000011; // 3532 :   3 - 0x3
      12'hDCD: dout  = 8'b00000001; // 3533 :   1 - 0x1
      12'hDCE: dout  = 8'b00000001; // 3534 :   1 - 0x1
      12'hDCF: dout  = 8'b00001111; // 3535 :  15 - 0xf
      12'hDD0: dout  = 8'b00001000; // 3536 :   8 - 0x8 -- Sprite 0xdd
      12'hDD1: dout  = 8'b00001101; // 3537 :  13 - 0xd
      12'hDD2: dout  = 8'b00111010; // 3538 :  58 - 0x3a
      12'hDD3: dout  = 8'b00100101; // 3539 :  37 - 0x25
      12'hDD4: dout  = 8'b00011011; // 3540 :  27 - 0x1b
      12'hDD5: dout  = 8'b00001111; // 3541 :  15 - 0xf
      12'hDD6: dout  = 8'b00000111; // 3542 :   7 - 0x7
      12'hDD7: dout  = 8'b00000011; // 3543 :   3 - 0x3
      12'hDD8: dout  = 8'b00000111; // 3544 :   7 - 0x7 -- plane 1
      12'hDD9: dout  = 8'b00000111; // 3545 :   7 - 0x7
      12'hDDA: dout  = 8'b00000111; // 3546 :   7 - 0x7
      12'hDDB: dout  = 8'b00011111; // 3547 :  31 - 0x1f
      12'hDDC: dout  = 8'b00001111; // 3548 :  15 - 0xf
      12'hDDD: dout  = 8'b00000111; // 3549 :   7 - 0x7
      12'hDDE: dout  = 8'b00000011; // 3550 :   3 - 0x3
      12'hDDF: dout  = 8'b00000000; // 3551 :   0 - 0x0
      12'hDE0: dout  = 8'b00000000; // 3552 :   0 - 0x0 -- Sprite 0xde
      12'hDE1: dout  = 8'b00000000; // 3553 :   0 - 0x0
      12'hDE2: dout  = 8'b00000000; // 3554 :   0 - 0x0
      12'hDE3: dout  = 8'b11000000; // 3555 : 192 - 0xc0
      12'hDE4: dout  = 8'b01000000; // 3556 :  64 - 0x40
      12'hDE5: dout  = 8'b01011000; // 3557 :  88 - 0x58
      12'hDE6: dout  = 8'b01101000; // 3558 : 104 - 0x68
      12'hDE7: dout  = 8'b00001000; // 3559 :   8 - 0x8
      12'hDE8: dout  = 8'b00000000; // 3560 :   0 - 0x0 -- plane 1
      12'hDE9: dout  = 8'b00000000; // 3561 :   0 - 0x0
      12'hDEA: dout  = 8'b00000000; // 3562 :   0 - 0x0
      12'hDEB: dout  = 8'b00000000; // 3563 :   0 - 0x0
      12'hDEC: dout  = 8'b10000000; // 3564 : 128 - 0x80
      12'hDED: dout  = 8'b10000000; // 3565 : 128 - 0x80
      12'hDEE: dout  = 8'b10010000; // 3566 : 144 - 0x90
      12'hDEF: dout  = 8'b11110000; // 3567 : 240 - 0xf0
      12'hDF0: dout  = 8'b00010000; // 3568 :  16 - 0x10 -- Sprite 0xdf
      12'hDF1: dout  = 8'b01011100; // 3569 :  92 - 0x5c
      12'hDF2: dout  = 8'b10101000; // 3570 : 168 - 0xa8
      12'hDF3: dout  = 8'b11011000; // 3571 : 216 - 0xd8
      12'hDF4: dout  = 8'b10111000; // 3572 : 184 - 0xb8
      12'hDF5: dout  = 8'b11110000; // 3573 : 240 - 0xf0
      12'hDF6: dout  = 8'b11100000; // 3574 : 224 - 0xe0
      12'hDF7: dout  = 8'b11000000; // 3575 : 192 - 0xc0
      12'hDF8: dout  = 8'b11100000; // 3576 : 224 - 0xe0 -- plane 1
      12'hDF9: dout  = 8'b11100000; // 3577 : 224 - 0xe0
      12'hDFA: dout  = 8'b11110000; // 3578 : 240 - 0xf0
      12'hDFB: dout  = 8'b11110000; // 3579 : 240 - 0xf0
      12'hDFC: dout  = 8'b11100000; // 3580 : 224 - 0xe0
      12'hDFD: dout  = 8'b11000000; // 3581 : 192 - 0xc0
      12'hDFE: dout  = 8'b11000000; // 3582 : 192 - 0xc0
      12'hDFF: dout  = 8'b00000000; // 3583 :   0 - 0x0
      12'hE00: dout  = 8'b00000000; // 3584 :   0 - 0x0 -- Sprite 0xe0
      12'hE01: dout  = 8'b00000000; // 3585 :   0 - 0x0
      12'hE02: dout  = 8'b00000000; // 3586 :   0 - 0x0
      12'hE03: dout  = 8'b00010011; // 3587 :  19 - 0x13
      12'hE04: dout  = 8'b00010011; // 3588 :  19 - 0x13
      12'hE05: dout  = 8'b00110111; // 3589 :  55 - 0x37
      12'hE06: dout  = 8'b00110111; // 3590 :  55 - 0x37
      12'hE07: dout  = 8'b00000111; // 3591 :   7 - 0x7
      12'hE08: dout  = 8'b00001111; // 3592 :  15 - 0xf -- plane 1
      12'hE09: dout  = 8'b00011111; // 3593 :  31 - 0x1f
      12'hE0A: dout  = 8'b00011111; // 3594 :  31 - 0x1f
      12'hE0B: dout  = 8'b00111111; // 3595 :  63 - 0x3f
      12'hE0C: dout  = 8'b01111111; // 3596 : 127 - 0x7f
      12'hE0D: dout  = 8'b11111111; // 3597 : 255 - 0xff
      12'hE0E: dout  = 8'b11111111; // 3598 : 255 - 0xff
      12'hE0F: dout  = 8'b11111111; // 3599 : 255 - 0xff
      12'hE10: dout  = 8'b00000111; // 3600 :   7 - 0x7 -- Sprite 0xe1
      12'hE11: dout  = 8'b00000100; // 3601 :   4 - 0x4
      12'hE12: dout  = 8'b00000000; // 3602 :   0 - 0x0
      12'hE13: dout  = 8'b00000000; // 3603 :   0 - 0x0
      12'hE14: dout  = 8'b00000000; // 3604 :   0 - 0x0
      12'hE15: dout  = 8'b00100000; // 3605 :  32 - 0x20
      12'hE16: dout  = 8'b01110000; // 3606 : 112 - 0x70
      12'hE17: dout  = 8'b11111000; // 3607 : 248 - 0xf8
      12'hE18: dout  = 8'b11111111; // 3608 : 255 - 0xff -- plane 1
      12'hE19: dout  = 8'b11111111; // 3609 : 255 - 0xff
      12'hE1A: dout  = 8'b01111111; // 3610 : 127 - 0x7f
      12'hE1B: dout  = 8'b00111111; // 3611 :  63 - 0x3f
      12'hE1C: dout  = 8'b00111111; // 3612 :  63 - 0x3f
      12'hE1D: dout  = 8'b00011111; // 3613 :  31 - 0x1f
      12'hE1E: dout  = 8'b00001111; // 3614 :  15 - 0xf
      12'hE1F: dout  = 8'b00000111; // 3615 :   7 - 0x7
      12'hE20: dout  = 8'b00000000; // 3616 :   0 - 0x0 -- Sprite 0xe2
      12'hE21: dout  = 8'b00000000; // 3617 :   0 - 0x0
      12'hE22: dout  = 8'b00000000; // 3618 :   0 - 0x0
      12'hE23: dout  = 8'b11111000; // 3619 : 248 - 0xf8
      12'hE24: dout  = 8'b11111100; // 3620 : 252 - 0xfc
      12'hE25: dout  = 8'b11111100; // 3621 : 252 - 0xfc
      12'hE26: dout  = 8'b11111100; // 3622 : 252 - 0xfc
      12'hE27: dout  = 8'b11111101; // 3623 : 253 - 0xfd
      12'hE28: dout  = 8'b11111110; // 3624 : 254 - 0xfe -- plane 1
      12'hE29: dout  = 8'b11111111; // 3625 : 255 - 0xff
      12'hE2A: dout  = 8'b11111111; // 3626 : 255 - 0xff
      12'hE2B: dout  = 8'b00001111; // 3627 :  15 - 0xf
      12'hE2C: dout  = 8'b10111111; // 3628 : 191 - 0xbf
      12'hE2D: dout  = 8'b10100011; // 3629 : 163 - 0xa3
      12'hE2E: dout  = 8'b11110111; // 3630 : 247 - 0xf7
      12'hE2F: dout  = 8'b11110111; // 3631 : 247 - 0xf7
      12'hE30: dout  = 8'b11111100; // 3632 : 252 - 0xfc -- Sprite 0xe3
      12'hE31: dout  = 8'b00011100; // 3633 :  28 - 0x1c
      12'hE32: dout  = 8'b11000000; // 3634 : 192 - 0xc0
      12'hE33: dout  = 8'b11100000; // 3635 : 224 - 0xe0
      12'hE34: dout  = 8'b00000000; // 3636 :   0 - 0x0
      12'hE35: dout  = 8'b00000000; // 3637 :   0 - 0x0
      12'hE36: dout  = 8'b00000110; // 3638 :   6 - 0x6
      12'hE37: dout  = 8'b00001111; // 3639 :  15 - 0xf
      12'hE38: dout  = 8'b11111111; // 3640 : 255 - 0xff -- plane 1
      12'hE39: dout  = 8'b11111111; // 3641 : 255 - 0xff
      12'hE3A: dout  = 8'b00111111; // 3642 :  63 - 0x3f
      12'hE3B: dout  = 8'b00011111; // 3643 :  31 - 0x1f
      12'hE3C: dout  = 8'b11111110; // 3644 : 254 - 0xfe
      12'hE3D: dout  = 8'b11111100; // 3645 : 252 - 0xfc
      12'hE3E: dout  = 8'b11111000; // 3646 : 248 - 0xf8
      12'hE3F: dout  = 8'b11110000; // 3647 : 240 - 0xf0
      12'hE40: dout  = 8'b00000000; // 3648 :   0 - 0x0 -- Sprite 0xe4
      12'hE41: dout  = 8'b00000000; // 3649 :   0 - 0x0
      12'hE42: dout  = 8'b00000000; // 3650 :   0 - 0x0
      12'hE43: dout  = 8'b00010011; // 3651 :  19 - 0x13
      12'hE44: dout  = 8'b00010011; // 3652 :  19 - 0x13
      12'hE45: dout  = 8'b00110111; // 3653 :  55 - 0x37
      12'hE46: dout  = 8'b00110111; // 3654 :  55 - 0x37
      12'hE47: dout  = 8'b00000111; // 3655 :   7 - 0x7
      12'hE48: dout  = 8'b00001111; // 3656 :  15 - 0xf -- plane 1
      12'hE49: dout  = 8'b00011111; // 3657 :  31 - 0x1f
      12'hE4A: dout  = 8'b00011111; // 3658 :  31 - 0x1f
      12'hE4B: dout  = 8'b00111111; // 3659 :  63 - 0x3f
      12'hE4C: dout  = 8'b01111111; // 3660 : 127 - 0x7f
      12'hE4D: dout  = 8'b11111111; // 3661 : 255 - 0xff
      12'hE4E: dout  = 8'b11111111; // 3662 : 255 - 0xff
      12'hE4F: dout  = 8'b11111111; // 3663 : 255 - 0xff
      12'hE50: dout  = 8'b00000111; // 3664 :   7 - 0x7 -- Sprite 0xe5
      12'hE51: dout  = 8'b00000100; // 3665 :   4 - 0x4
      12'hE52: dout  = 8'b00000001; // 3666 :   1 - 0x1
      12'hE53: dout  = 8'b00000000; // 3667 :   0 - 0x0
      12'hE54: dout  = 8'b00000000; // 3668 :   0 - 0x0
      12'hE55: dout  = 8'b00100000; // 3669 :  32 - 0x20
      12'hE56: dout  = 8'b01110000; // 3670 : 112 - 0x70
      12'hE57: dout  = 8'b11111000; // 3671 : 248 - 0xf8
      12'hE58: dout  = 8'b11111111; // 3672 : 255 - 0xff -- plane 1
      12'hE59: dout  = 8'b11111111; // 3673 : 255 - 0xff
      12'hE5A: dout  = 8'b01111110; // 3674 : 126 - 0x7e
      12'hE5B: dout  = 8'b00111111; // 3675 :  63 - 0x3f
      12'hE5C: dout  = 8'b00111111; // 3676 :  63 - 0x3f
      12'hE5D: dout  = 8'b00011111; // 3677 :  31 - 0x1f
      12'hE5E: dout  = 8'b00001111; // 3678 :  15 - 0xf
      12'hE5F: dout  = 8'b00000111; // 3679 :   7 - 0x7
      12'hE60: dout  = 8'b00000000; // 3680 :   0 - 0x0 -- Sprite 0xe6
      12'hE61: dout  = 8'b00000000; // 3681 :   0 - 0x0
      12'hE62: dout  = 8'b00000000; // 3682 :   0 - 0x0
      12'hE63: dout  = 8'b11111100; // 3683 : 252 - 0xfc
      12'hE64: dout  = 8'b11111100; // 3684 : 252 - 0xfc
      12'hE65: dout  = 8'b11111100; // 3685 : 252 - 0xfc
      12'hE66: dout  = 8'b11111100; // 3686 : 252 - 0xfc
      12'hE67: dout  = 8'b11111101; // 3687 : 253 - 0xfd
      12'hE68: dout  = 8'b11111110; // 3688 : 254 - 0xfe -- plane 1
      12'hE69: dout  = 8'b11111111; // 3689 : 255 - 0xff
      12'hE6A: dout  = 8'b11111111; // 3690 : 255 - 0xff
      12'hE6B: dout  = 8'b11100011; // 3691 : 227 - 0xe3
      12'hE6C: dout  = 8'b00010111; // 3692 :  23 - 0x17
      12'hE6D: dout  = 8'b10110111; // 3693 : 183 - 0xb7
      12'hE6E: dout  = 8'b10111111; // 3694 : 191 - 0xbf
      12'hE6F: dout  = 8'b11111111; // 3695 : 255 - 0xff
      12'hE70: dout  = 8'b11111100; // 3696 : 252 - 0xfc -- Sprite 0xe7
      12'hE71: dout  = 8'b00001100; // 3697 :  12 - 0xc
      12'hE72: dout  = 8'b11000000; // 3698 : 192 - 0xc0
      12'hE73: dout  = 8'b11110000; // 3699 : 240 - 0xf0
      12'hE74: dout  = 8'b11110000; // 3700 : 240 - 0xf0
      12'hE75: dout  = 8'b00000000; // 3701 :   0 - 0x0
      12'hE76: dout  = 8'b00000110; // 3702 :   6 - 0x6
      12'hE77: dout  = 8'b00001111; // 3703 :  15 - 0xf
      12'hE78: dout  = 8'b11111111; // 3704 : 255 - 0xff -- plane 1
      12'hE79: dout  = 8'b11111111; // 3705 : 255 - 0xff
      12'hE7A: dout  = 8'b00111111; // 3706 :  63 - 0x3f
      12'hE7B: dout  = 8'b00001111; // 3707 :  15 - 0xf
      12'hE7C: dout  = 8'b00001110; // 3708 :  14 - 0xe
      12'hE7D: dout  = 8'b11111100; // 3709 : 252 - 0xfc
      12'hE7E: dout  = 8'b11111000; // 3710 : 248 - 0xf8
      12'hE7F: dout  = 8'b11110000; // 3711 : 240 - 0xf0
      12'hE80: dout  = 8'b11111111; // 3712 : 255 - 0xff -- Sprite 0xe8
      12'hE81: dout  = 8'b11111111; // 3713 : 255 - 0xff
      12'hE82: dout  = 8'b01111111; // 3714 : 127 - 0x7f
      12'hE83: dout  = 8'b01111111; // 3715 : 127 - 0x7f
      12'hE84: dout  = 8'b01111111; // 3716 : 127 - 0x7f
      12'hE85: dout  = 8'b00111111; // 3717 :  63 - 0x3f
      12'hE86: dout  = 8'b00111111; // 3718 :  63 - 0x3f
      12'hE87: dout  = 8'b00111111; // 3719 :  63 - 0x3f
      12'hE88: dout  = 8'b00000000; // 3720 :   0 - 0x0 -- plane 1
      12'hE89: dout  = 8'b00000101; // 3721 :   5 - 0x5
      12'hE8A: dout  = 8'b00000111; // 3722 :   7 - 0x7
      12'hE8B: dout  = 8'b00000011; // 3723 :   3 - 0x3
      12'hE8C: dout  = 8'b00000000; // 3724 :   0 - 0x0
      12'hE8D: dout  = 8'b00000000; // 3725 :   0 - 0x0
      12'hE8E: dout  = 8'b00000000; // 3726 :   0 - 0x0
      12'hE8F: dout  = 8'b00000000; // 3727 :   0 - 0x0
      12'hE90: dout  = 8'b00111100; // 3728 :  60 - 0x3c -- Sprite 0xe9
      12'hE91: dout  = 8'b00111110; // 3729 :  62 - 0x3e
      12'hE92: dout  = 8'b00011111; // 3730 :  31 - 0x1f
      12'hE93: dout  = 8'b00001111; // 3731 :  15 - 0xf
      12'hE94: dout  = 8'b00000111; // 3732 :   7 - 0x7
      12'hE95: dout  = 8'b00000000; // 3733 :   0 - 0x0
      12'hE96: dout  = 8'b00000000; // 3734 :   0 - 0x0
      12'hE97: dout  = 8'b00000000; // 3735 :   0 - 0x0
      12'hE98: dout  = 8'b00000000; // 3736 :   0 - 0x0 -- plane 1
      12'hE99: dout  = 8'b00000000; // 3737 :   0 - 0x0
      12'hE9A: dout  = 8'b00000000; // 3738 :   0 - 0x0
      12'hE9B: dout  = 8'b00000000; // 3739 :   0 - 0x0
      12'hE9C: dout  = 8'b00000000; // 3740 :   0 - 0x0
      12'hE9D: dout  = 8'b00000000; // 3741 :   0 - 0x0
      12'hE9E: dout  = 8'b00000000; // 3742 :   0 - 0x0
      12'hE9F: dout  = 8'b00000000; // 3743 :   0 - 0x0
      12'hEA0: dout  = 8'b11111111; // 3744 : 255 - 0xff -- Sprite 0xea
      12'hEA1: dout  = 8'b11111110; // 3745 : 254 - 0xfe
      12'hEA2: dout  = 8'b11111110; // 3746 : 254 - 0xfe
      12'hEA3: dout  = 8'b11111100; // 3747 : 252 - 0xfc
      12'hEA4: dout  = 8'b11111000; // 3748 : 248 - 0xf8
      12'hEA5: dout  = 8'b11110000; // 3749 : 240 - 0xf0
      12'hEA6: dout  = 8'b10110000; // 3750 : 176 - 0xb0
      12'hEA7: dout  = 8'b00111001; // 3751 :  57 - 0x39
      12'hEA8: dout  = 8'b00000011; // 3752 :   3 - 0x3 -- plane 1
      12'hEA9: dout  = 8'b10011110; // 3753 : 158 - 0x9e
      12'hEAA: dout  = 8'b00001110; // 3754 :  14 - 0xe
      12'hEAB: dout  = 8'b00000000; // 3755 :   0 - 0x0
      12'hEAC: dout  = 8'b00000000; // 3756 :   0 - 0x0
      12'hEAD: dout  = 8'b00000000; // 3757 :   0 - 0x0
      12'hEAE: dout  = 8'b00000000; // 3758 :   0 - 0x0
      12'hEAF: dout  = 8'b00000000; // 3759 :   0 - 0x0
      12'hEB0: dout  = 8'b00011111; // 3760 :  31 - 0x1f -- Sprite 0xeb
      12'hEB1: dout  = 8'b11001111; // 3761 : 207 - 0xcf
      12'hEB2: dout  = 8'b11000110; // 3762 : 198 - 0xc6
      12'hEB3: dout  = 8'b10000000; // 3763 : 128 - 0x80
      12'hEB4: dout  = 8'b00000000; // 3764 :   0 - 0x0
      12'hEB5: dout  = 8'b00000000; // 3765 :   0 - 0x0
      12'hEB6: dout  = 8'b00000000; // 3766 :   0 - 0x0
      12'hEB7: dout  = 8'b00000000; // 3767 :   0 - 0x0
      12'hEB8: dout  = 8'b00000000; // 3768 :   0 - 0x0 -- plane 1
      12'hEB9: dout  = 8'b00000000; // 3769 :   0 - 0x0
      12'hEBA: dout  = 8'b00000000; // 3770 :   0 - 0x0
      12'hEBB: dout  = 8'b00000000; // 3771 :   0 - 0x0
      12'hEBC: dout  = 8'b00000000; // 3772 :   0 - 0x0
      12'hEBD: dout  = 8'b00000000; // 3773 :   0 - 0x0
      12'hEBE: dout  = 8'b00000000; // 3774 :   0 - 0x0
      12'hEBF: dout  = 8'b00000000; // 3775 :   0 - 0x0
      12'hEC0: dout  = 8'b00000000; // 3776 :   0 - 0x0 -- Sprite 0xec
      12'hEC1: dout  = 8'b00000000; // 3777 :   0 - 0x0
      12'hEC2: dout  = 8'b00000000; // 3778 :   0 - 0x0
      12'hEC3: dout  = 8'b00000000; // 3779 :   0 - 0x0
      12'hEC4: dout  = 8'b00000000; // 3780 :   0 - 0x0
      12'hEC5: dout  = 8'b00000000; // 3781 :   0 - 0x0
      12'hEC6: dout  = 8'b00001100; // 3782 :  12 - 0xc
      12'hEC7: dout  = 8'b00001100; // 3783 :  12 - 0xc
      12'hEC8: dout  = 8'b00000000; // 3784 :   0 - 0x0 -- plane 1
      12'hEC9: dout  = 8'b00000000; // 3785 :   0 - 0x0
      12'hECA: dout  = 8'b00000000; // 3786 :   0 - 0x0
      12'hECB: dout  = 8'b00000000; // 3787 :   0 - 0x0
      12'hECC: dout  = 8'b00000100; // 3788 :   4 - 0x4
      12'hECD: dout  = 8'b00001110; // 3789 :  14 - 0xe
      12'hECE: dout  = 8'b00001111; // 3790 :  15 - 0xf
      12'hECF: dout  = 8'b00001011; // 3791 :  11 - 0xb
      12'hED0: dout  = 8'b00110000; // 3792 :  48 - 0x30 -- Sprite 0xed
      12'hED1: dout  = 8'b01000011; // 3793 :  67 - 0x43
      12'hED2: dout  = 8'b01000000; // 3794 :  64 - 0x40
      12'hED3: dout  = 8'b01100000; // 3795 :  96 - 0x60
      12'hED4: dout  = 8'b00000011; // 3796 :   3 - 0x3
      12'hED5: dout  = 8'b00000000; // 3797 :   0 - 0x0
      12'hED6: dout  = 8'b01111111; // 3798 : 127 - 0x7f
      12'hED7: dout  = 8'b00000000; // 3799 :   0 - 0x0
      12'hED8: dout  = 8'b00001111; // 3800 :  15 - 0xf -- plane 1
      12'hED9: dout  = 8'b00001100; // 3801 :  12 - 0xc
      12'hEDA: dout  = 8'b00001111; // 3802 :  15 - 0xf
      12'hEDB: dout  = 8'b00001111; // 3803 :  15 - 0xf
      12'hEDC: dout  = 8'b00000000; // 3804 :   0 - 0x0
      12'hEDD: dout  = 8'b01111111; // 3805 : 127 - 0x7f
      12'hEDE: dout  = 8'b11010101; // 3806 : 213 - 0xd5
      12'hEDF: dout  = 8'b01111111; // 3807 : 127 - 0x7f
      12'hEE0: dout  = 8'b00000000; // 3808 :   0 - 0x0 -- Sprite 0xee
      12'hEE1: dout  = 8'b00000000; // 3809 :   0 - 0x0
      12'hEE2: dout  = 8'b00000000; // 3810 :   0 - 0x0
      12'hEE3: dout  = 8'b00000000; // 3811 :   0 - 0x0
      12'hEE4: dout  = 8'b00000000; // 3812 :   0 - 0x0
      12'hEE5: dout  = 8'b00000000; // 3813 :   0 - 0x0
      12'hEE6: dout  = 8'b00110000; // 3814 :  48 - 0x30
      12'hEE7: dout  = 8'b00110000; // 3815 :  48 - 0x30
      12'hEE8: dout  = 8'b00000000; // 3816 :   0 - 0x0 -- plane 1
      12'hEE9: dout  = 8'b00000000; // 3817 :   0 - 0x0
      12'hEEA: dout  = 8'b00000000; // 3818 :   0 - 0x0
      12'hEEB: dout  = 8'b00000000; // 3819 :   0 - 0x0
      12'hEEC: dout  = 8'b00100000; // 3820 :  32 - 0x20
      12'hEED: dout  = 8'b01110000; // 3821 : 112 - 0x70
      12'hEEE: dout  = 8'b11110000; // 3822 : 240 - 0xf0
      12'hEEF: dout  = 8'b11100000; // 3823 : 224 - 0xe0
      12'hEF0: dout  = 8'b00001110; // 3824 :  14 - 0xe -- Sprite 0xef
      12'hEF1: dout  = 8'b11001011; // 3825 : 203 - 0xcb
      12'hEF2: dout  = 8'b00000000; // 3826 :   0 - 0x0
      12'hEF3: dout  = 8'b00000000; // 3827 :   0 - 0x0
      12'hEF4: dout  = 8'b11000000; // 3828 : 192 - 0xc0
      12'hEF5: dout  = 8'b00000000; // 3829 :   0 - 0x0
      12'hEF6: dout  = 8'b11111110; // 3830 : 254 - 0xfe
      12'hEF7: dout  = 8'b00000000; // 3831 :   0 - 0x0
      12'hEF8: dout  = 8'b11110000; // 3832 : 240 - 0xf0 -- plane 1
      12'hEF9: dout  = 8'b00110000; // 3833 :  48 - 0x30
      12'hEFA: dout  = 8'b11110000; // 3834 : 240 - 0xf0
      12'hEFB: dout  = 8'b11110000; // 3835 : 240 - 0xf0
      12'hEFC: dout  = 8'b00000000; // 3836 :   0 - 0x0
      12'hEFD: dout  = 8'b11111110; // 3837 : 254 - 0xfe
      12'hEFE: dout  = 8'b01010101; // 3838 :  85 - 0x55
      12'hEFF: dout  = 8'b11111110; // 3839 : 254 - 0xfe
      12'hF00: dout  = 8'b00000000; // 3840 :   0 - 0x0 -- Sprite 0xf0
      12'hF01: dout  = 8'b00000000; // 3841 :   0 - 0x0
      12'hF02: dout  = 8'b00000000; // 3842 :   0 - 0x0
      12'hF03: dout  = 8'b00000000; // 3843 :   0 - 0x0
      12'hF04: dout  = 8'b00000000; // 3844 :   0 - 0x0
      12'hF05: dout  = 8'b00000000; // 3845 :   0 - 0x0
      12'hF06: dout  = 8'b00001100; // 3846 :  12 - 0xc
      12'hF07: dout  = 8'b00001100; // 3847 :  12 - 0xc
      12'hF08: dout  = 8'b00000000; // 3848 :   0 - 0x0 -- plane 1
      12'hF09: dout  = 8'b00000000; // 3849 :   0 - 0x0
      12'hF0A: dout  = 8'b00000000; // 3850 :   0 - 0x0
      12'hF0B: dout  = 8'b00000000; // 3851 :   0 - 0x0
      12'hF0C: dout  = 8'b00000100; // 3852 :   4 - 0x4
      12'hF0D: dout  = 8'b00001110; // 3853 :  14 - 0xe
      12'hF0E: dout  = 8'b00001111; // 3854 :  15 - 0xf
      12'hF0F: dout  = 8'b00001011; // 3855 :  11 - 0xb
      12'hF10: dout  = 8'b00110000; // 3856 :  48 - 0x30 -- Sprite 0xf1
      12'hF11: dout  = 8'b00100011; // 3857 :  35 - 0x23
      12'hF12: dout  = 8'b00100000; // 3858 :  32 - 0x20
      12'hF13: dout  = 8'b01100000; // 3859 :  96 - 0x60
      12'hF14: dout  = 8'b00000011; // 3860 :   3 - 0x3
      12'hF15: dout  = 8'b00000000; // 3861 :   0 - 0x0
      12'hF16: dout  = 8'b01111111; // 3862 : 127 - 0x7f
      12'hF17: dout  = 8'b00000000; // 3863 :   0 - 0x0
      12'hF18: dout  = 8'b00001111; // 3864 :  15 - 0xf -- plane 1
      12'hF19: dout  = 8'b00001100; // 3865 :  12 - 0xc
      12'hF1A: dout  = 8'b00001111; // 3866 :  15 - 0xf
      12'hF1B: dout  = 8'b00001111; // 3867 :  15 - 0xf
      12'hF1C: dout  = 8'b00000000; // 3868 :   0 - 0x0
      12'hF1D: dout  = 8'b01111111; // 3869 : 127 - 0x7f
      12'hF1E: dout  = 8'b10101010; // 3870 : 170 - 0xaa
      12'hF1F: dout  = 8'b01111111; // 3871 : 127 - 0x7f
      12'hF20: dout  = 8'b00000000; // 3872 :   0 - 0x0 -- Sprite 0xf2
      12'hF21: dout  = 8'b00000000; // 3873 :   0 - 0x0
      12'hF22: dout  = 8'b00000000; // 3874 :   0 - 0x0
      12'hF23: dout  = 8'b00000000; // 3875 :   0 - 0x0
      12'hF24: dout  = 8'b00000000; // 3876 :   0 - 0x0
      12'hF25: dout  = 8'b00000000; // 3877 :   0 - 0x0
      12'hF26: dout  = 8'b00110000; // 3878 :  48 - 0x30
      12'hF27: dout  = 8'b00110000; // 3879 :  48 - 0x30
      12'hF28: dout  = 8'b00000000; // 3880 :   0 - 0x0 -- plane 1
      12'hF29: dout  = 8'b00000000; // 3881 :   0 - 0x0
      12'hF2A: dout  = 8'b00000000; // 3882 :   0 - 0x0
      12'hF2B: dout  = 8'b00000000; // 3883 :   0 - 0x0
      12'hF2C: dout  = 8'b00100000; // 3884 :  32 - 0x20
      12'hF2D: dout  = 8'b01110000; // 3885 : 112 - 0x70
      12'hF2E: dout  = 8'b11110000; // 3886 : 240 - 0xf0
      12'hF2F: dout  = 8'b11100000; // 3887 : 224 - 0xe0
      12'hF30: dout  = 8'b00001001; // 3888 :   9 - 0x9 -- Sprite 0xf3
      12'hF31: dout  = 8'b11001111; // 3889 : 207 - 0xcf
      12'hF32: dout  = 8'b00000000; // 3890 :   0 - 0x0
      12'hF33: dout  = 8'b00000000; // 3891 :   0 - 0x0
      12'hF34: dout  = 8'b11000000; // 3892 : 192 - 0xc0
      12'hF35: dout  = 8'b00000000; // 3893 :   0 - 0x0
      12'hF36: dout  = 8'b11111110; // 3894 : 254 - 0xfe
      12'hF37: dout  = 8'b00000000; // 3895 :   0 - 0x0
      12'hF38: dout  = 8'b11110000; // 3896 : 240 - 0xf0 -- plane 1
      12'hF39: dout  = 8'b00110000; // 3897 :  48 - 0x30
      12'hF3A: dout  = 8'b11110000; // 3898 : 240 - 0xf0
      12'hF3B: dout  = 8'b11110000; // 3899 : 240 - 0xf0
      12'hF3C: dout  = 8'b00000000; // 3900 :   0 - 0x0
      12'hF3D: dout  = 8'b11111110; // 3901 : 254 - 0xfe
      12'hF3E: dout  = 8'b10101011; // 3902 : 171 - 0xab
      12'hF3F: dout  = 8'b11111110; // 3903 : 254 - 0xfe
      12'hF40: dout  = 8'b00111111; // 3904 :  63 - 0x3f -- Sprite 0xf4
      12'hF41: dout  = 8'b00110101; // 3905 :  53 - 0x35
      12'hF42: dout  = 8'b00011010; // 3906 :  26 - 0x1a
      12'hF43: dout  = 8'b00001101; // 3907 :  13 - 0xd
      12'hF44: dout  = 8'b00001010; // 3908 :  10 - 0xa
      12'hF45: dout  = 8'b00001101; // 3909 :  13 - 0xd
      12'hF46: dout  = 8'b00001000; // 3910 :   8 - 0x8
      12'hF47: dout  = 8'b00111000; // 3911 :  56 - 0x38
      12'hF48: dout  = 8'b00000000; // 3912 :   0 - 0x0 -- plane 1
      12'hF49: dout  = 8'b00010101; // 3913 :  21 - 0x15
      12'hF4A: dout  = 8'b00001010; // 3914 :  10 - 0xa
      12'hF4B: dout  = 8'b00000101; // 3915 :   5 - 0x5
      12'hF4C: dout  = 8'b00000010; // 3916 :   2 - 0x2
      12'hF4D: dout  = 8'b00000101; // 3917 :   5 - 0x5
      12'hF4E: dout  = 8'b00000111; // 3918 :   7 - 0x7
      12'hF4F: dout  = 8'b00000111; // 3919 :   7 - 0x7
      12'hF50: dout  = 8'b01110011; // 3920 : 115 - 0x73 -- Sprite 0xf5
      12'hF51: dout  = 8'b11000100; // 3921 : 196 - 0xc4
      12'hF52: dout  = 8'b11000100; // 3922 : 196 - 0xc4
      12'hF53: dout  = 8'b11000000; // 3923 : 192 - 0xc0
      12'hF54: dout  = 8'b11000001; // 3924 : 193 - 0xc1
      12'hF55: dout  = 8'b11000000; // 3925 : 192 - 0xc0
      12'hF56: dout  = 8'b01100001; // 3926 :  97 - 0x61
      12'hF57: dout  = 8'b00111111; // 3927 :  63 - 0x3f
      12'hF58: dout  = 8'b00111100; // 3928 :  60 - 0x3c -- plane 1
      12'hF59: dout  = 8'b01111011; // 3929 : 123 - 0x7b
      12'hF5A: dout  = 8'b01111011; // 3930 : 123 - 0x7b
      12'hF5B: dout  = 8'b01111111; // 3931 : 127 - 0x7f
      12'hF5C: dout  = 8'b01111110; // 3932 : 126 - 0x7e
      12'hF5D: dout  = 8'b01111111; // 3933 : 127 - 0x7f
      12'hF5E: dout  = 8'b00111110; // 3934 :  62 - 0x3e
      12'hF5F: dout  = 8'b00000000; // 3935 :   0 - 0x0
      12'hF60: dout  = 8'b11111100; // 3936 : 252 - 0xfc -- Sprite 0xf6
      12'hF61: dout  = 8'b01010100; // 3937 :  84 - 0x54
      12'hF62: dout  = 8'b10101000; // 3938 : 168 - 0xa8
      12'hF63: dout  = 8'b01010000; // 3939 :  80 - 0x50
      12'hF64: dout  = 8'b10110000; // 3940 : 176 - 0xb0
      12'hF65: dout  = 8'b01010000; // 3941 :  80 - 0x50
      12'hF66: dout  = 8'b10010000; // 3942 : 144 - 0x90
      12'hF67: dout  = 8'b00011100; // 3943 :  28 - 0x1c
      12'hF68: dout  = 8'b00000000; // 3944 :   0 - 0x0 -- plane 1
      12'hF69: dout  = 8'b01010000; // 3945 :  80 - 0x50
      12'hF6A: dout  = 8'b10100000; // 3946 : 160 - 0xa0
      12'hF6B: dout  = 8'b01000000; // 3947 :  64 - 0x40
      12'hF6C: dout  = 8'b10100000; // 3948 : 160 - 0xa0
      12'hF6D: dout  = 8'b01000000; // 3949 :  64 - 0x40
      12'hF6E: dout  = 8'b11100000; // 3950 : 224 - 0xe0
      12'hF6F: dout  = 8'b11100000; // 3951 : 224 - 0xe0
      12'hF70: dout  = 8'b10000110; // 3952 : 134 - 0x86 -- Sprite 0xf7
      12'hF71: dout  = 8'b01000010; // 3953 :  66 - 0x42
      12'hF72: dout  = 8'b01000111; // 3954 :  71 - 0x47
      12'hF73: dout  = 8'b01000001; // 3955 :  65 - 0x41
      12'hF74: dout  = 8'b10000011; // 3956 : 131 - 0x83
      12'hF75: dout  = 8'b00000001; // 3957 :   1 - 0x1
      12'hF76: dout  = 8'b10000110; // 3958 : 134 - 0x86
      12'hF77: dout  = 8'b11111100; // 3959 : 252 - 0xfc
      12'hF78: dout  = 8'b01111000; // 3960 : 120 - 0x78 -- plane 1
      12'hF79: dout  = 8'b10111100; // 3961 : 188 - 0xbc
      12'hF7A: dout  = 8'b10111000; // 3962 : 184 - 0xb8
      12'hF7B: dout  = 8'b10111110; // 3963 : 190 - 0xbe
      12'hF7C: dout  = 8'b01111100; // 3964 : 124 - 0x7c
      12'hF7D: dout  = 8'b11111110; // 3965 : 254 - 0xfe
      12'hF7E: dout  = 8'b01111000; // 3966 : 120 - 0x78
      12'hF7F: dout  = 8'b00000000; // 3967 :   0 - 0x0
      12'hF80: dout  = 8'b11100100; // 3968 : 228 - 0xe4 -- Sprite 0xf8
      12'hF81: dout  = 8'b11100100; // 3969 : 228 - 0xe4
      12'hF82: dout  = 8'b11101111; // 3970 : 239 - 0xef
      12'hF83: dout  = 8'b11101111; // 3971 : 239 - 0xef
      12'hF84: dout  = 8'b11111111; // 3972 : 255 - 0xff
      12'hF85: dout  = 8'b11111111; // 3973 : 255 - 0xff
      12'hF86: dout  = 8'b01111111; // 3974 : 127 - 0x7f
      12'hF87: dout  = 8'b01111111; // 3975 : 127 - 0x7f
      12'hF88: dout  = 8'b00000011; // 3976 :   3 - 0x3 -- plane 1
      12'hF89: dout  = 8'b00000011; // 3977 :   3 - 0x3
      12'hF8A: dout  = 8'b00000000; // 3978 :   0 - 0x0
      12'hF8B: dout  = 8'b00000011; // 3979 :   3 - 0x3
      12'hF8C: dout  = 8'b00000111; // 3980 :   7 - 0x7
      12'hF8D: dout  = 8'b00000110; // 3981 :   6 - 0x6
      12'hF8E: dout  = 8'b00000111; // 3982 :   7 - 0x7
      12'hF8F: dout  = 8'b00000000; // 3983 :   0 - 0x0
      12'hF90: dout  = 8'b00111111; // 3984 :  63 - 0x3f -- Sprite 0xf9
      12'hF91: dout  = 8'b01111111; // 3985 : 127 - 0x7f
      12'hF92: dout  = 8'b01111111; // 3986 : 127 - 0x7f
      12'hF93: dout  = 8'b11111111; // 3987 : 255 - 0xff
      12'hF94: dout  = 8'b11111111; // 3988 : 255 - 0xff
      12'hF95: dout  = 8'b11111111; // 3989 : 255 - 0xff
      12'hF96: dout  = 8'b11111111; // 3990 : 255 - 0xff
      12'hF97: dout  = 8'b11111111; // 3991 : 255 - 0xff
      12'hF98: dout  = 8'b00000000; // 3992 :   0 - 0x0 -- plane 1
      12'hF99: dout  = 8'b00011111; // 3993 :  31 - 0x1f
      12'hF9A: dout  = 8'b00011111; // 3994 :  31 - 0x1f
      12'hF9B: dout  = 8'b00001111; // 3995 :  15 - 0xf
      12'hF9C: dout  = 8'b00000011; // 3996 :   3 - 0x3
      12'hF9D: dout  = 8'b00000000; // 3997 :   0 - 0x0
      12'hF9E: dout  = 8'b00000000; // 3998 :   0 - 0x0
      12'hF9F: dout  = 8'b00000000; // 3999 :   0 - 0x0
      12'hFA0: dout  = 8'b00010011; // 4000 :  19 - 0x13 -- Sprite 0xfa
      12'hFA1: dout  = 8'b00010011; // 4001 :  19 - 0x13
      12'hFA2: dout  = 8'b11111011; // 4002 : 251 - 0xfb
      12'hFA3: dout  = 8'b11111011; // 4003 : 251 - 0xfb
      12'hFA4: dout  = 8'b11111111; // 4004 : 255 - 0xff
      12'hFA5: dout  = 8'b11111111; // 4005 : 255 - 0xff
      12'hFA6: dout  = 8'b11111110; // 4006 : 254 - 0xfe
      12'hFA7: dout  = 8'b11111110; // 4007 : 254 - 0xfe
      12'hFA8: dout  = 8'b11100000; // 4008 : 224 - 0xe0 -- plane 1
      12'hFA9: dout  = 8'b11100000; // 4009 : 224 - 0xe0
      12'hFAA: dout  = 8'b00000000; // 4010 :   0 - 0x0
      12'hFAB: dout  = 8'b00110000; // 4011 :  48 - 0x30
      12'hFAC: dout  = 8'b01110000; // 4012 : 112 - 0x70
      12'hFAD: dout  = 8'b01100000; // 4013 :  96 - 0x60
      12'hFAE: dout  = 8'b01110000; // 4014 : 112 - 0x70
      12'hFAF: dout  = 8'b00000000; // 4015 :   0 - 0x0
      12'hFB0: dout  = 8'b11111110; // 4016 : 254 - 0xfe -- Sprite 0xfb
      12'hFB1: dout  = 8'b11111111; // 4017 : 255 - 0xff
      12'hFB2: dout  = 8'b11111111; // 4018 : 255 - 0xff
      12'hFB3: dout  = 8'b11111111; // 4019 : 255 - 0xff
      12'hFB4: dout  = 8'b11111111; // 4020 : 255 - 0xff
      12'hFB5: dout  = 8'b11111111; // 4021 : 255 - 0xff
      12'hFB6: dout  = 8'b11111111; // 4022 : 255 - 0xff
      12'hFB7: dout  = 8'b11111111; // 4023 : 255 - 0xff
      12'hFB8: dout  = 8'b00000000; // 4024 :   0 - 0x0 -- plane 1
      12'hFB9: dout  = 8'b11111000; // 4025 : 248 - 0xf8
      12'hFBA: dout  = 8'b11111000; // 4026 : 248 - 0xf8
      12'hFBB: dout  = 8'b11110000; // 4027 : 240 - 0xf0
      12'hFBC: dout  = 8'b11000000; // 4028 : 192 - 0xc0
      12'hFBD: dout  = 8'b00000000; // 4029 :   0 - 0x0
      12'hFBE: dout  = 8'b00000000; // 4030 :   0 - 0x0
      12'hFBF: dout  = 8'b00000000; // 4031 :   0 - 0x0
      12'hFC0: dout  = 8'b00000000; // 4032 :   0 - 0x0 -- Sprite 0xfc
      12'hFC1: dout  = 8'b00000000; // 4033 :   0 - 0x0
      12'hFC2: dout  = 8'b01111100; // 4034 : 124 - 0x7c
      12'hFC3: dout  = 8'b11111110; // 4035 : 254 - 0xfe
      12'hFC4: dout  = 8'b11111110; // 4036 : 254 - 0xfe
      12'hFC5: dout  = 8'b01111100; // 4037 : 124 - 0x7c
      12'hFC6: dout  = 8'b01000100; // 4038 :  68 - 0x44
      12'hFC7: dout  = 8'b10000010; // 4039 : 130 - 0x82
      12'hFC8: dout  = 8'b00111000; // 4040 :  56 - 0x38 -- plane 1
      12'hFC9: dout  = 8'b00111000; // 4041 :  56 - 0x38
      12'hFCA: dout  = 8'b00000000; // 4042 :   0 - 0x0
      12'hFCB: dout  = 8'b01111100; // 4043 : 124 - 0x7c
      12'hFCC: dout  = 8'b00000000; // 4044 :   0 - 0x0
      12'hFCD: dout  = 8'b00111000; // 4045 :  56 - 0x38
      12'hFCE: dout  = 8'b00111000; // 4046 :  56 - 0x38
      12'hFCF: dout  = 8'b01111100; // 4047 : 124 - 0x7c
      12'hFD0: dout  = 8'b10000010; // 4048 : 130 - 0x82 -- Sprite 0xfd
      12'hFD1: dout  = 8'b10000010; // 4049 : 130 - 0x82
      12'hFD2: dout  = 8'b10000010; // 4050 : 130 - 0x82
      12'hFD3: dout  = 8'b11000110; // 4051 : 198 - 0xc6
      12'hFD4: dout  = 8'b11111110; // 4052 : 254 - 0xfe
      12'hFD5: dout  = 8'b11111110; // 4053 : 254 - 0xfe
      12'hFD6: dout  = 8'b10111010; // 4054 : 186 - 0xba
      12'hFD7: dout  = 8'b01111100; // 4055 : 124 - 0x7c
      12'hFD8: dout  = 8'b01111100; // 4056 : 124 - 0x7c -- plane 1
      12'hFD9: dout  = 8'b01111100; // 4057 : 124 - 0x7c
      12'hFDA: dout  = 8'b01111100; // 4058 : 124 - 0x7c
      12'hFDB: dout  = 8'b00111000; // 4059 :  56 - 0x38
      12'hFDC: dout  = 8'b00000000; // 4060 :   0 - 0x0
      12'hFDD: dout  = 8'b01111100; // 4061 : 124 - 0x7c
      12'hFDE: dout  = 8'b01111100; // 4062 : 124 - 0x7c
      12'hFDF: dout  = 8'b00000000; // 4063 :   0 - 0x0
      12'hFE0: dout  = 8'b00000000; // 4064 :   0 - 0x0 -- Sprite 0xfe
      12'hFE1: dout  = 8'b00011001; // 4065 :  25 - 0x19
      12'hFE2: dout  = 8'b00111110; // 4066 :  62 - 0x3e
      12'hFE3: dout  = 8'b00111100; // 4067 :  60 - 0x3c
      12'hFE4: dout  = 8'b00111100; // 4068 :  60 - 0x3c
      12'hFE5: dout  = 8'b00111100; // 4069 :  60 - 0x3c
      12'hFE6: dout  = 8'b00111110; // 4070 :  62 - 0x3e
      12'hFE7: dout  = 8'b00011001; // 4071 :  25 - 0x19
      12'hFE8: dout  = 8'b00000000; // 4072 :   0 - 0x0 -- plane 1
      12'hFE9: dout  = 8'b00000000; // 4073 :   0 - 0x0
      12'hFEA: dout  = 8'b00010001; // 4074 :  17 - 0x11
      12'hFEB: dout  = 8'b11010111; // 4075 : 215 - 0xd7
      12'hFEC: dout  = 8'b11010111; // 4076 : 215 - 0xd7
      12'hFED: dout  = 8'b11010111; // 4077 : 215 - 0xd7
      12'hFEE: dout  = 8'b00010001; // 4078 :  17 - 0x11
      12'hFEF: dout  = 8'b00000000; // 4079 :   0 - 0x0
      12'hFF0: dout  = 8'b00000000; // 4080 :   0 - 0x0 -- Sprite 0xff
      12'hFF1: dout  = 8'b11111110; // 4081 : 254 - 0xfe
      12'hFF2: dout  = 8'b00011101; // 4082 :  29 - 0x1d
      12'hFF3: dout  = 8'b00001111; // 4083 :  15 - 0xf
      12'hFF4: dout  = 8'b00001111; // 4084 :  15 - 0xf
      12'hFF5: dout  = 8'b00001111; // 4085 :  15 - 0xf
      12'hFF6: dout  = 8'b00011101; // 4086 :  29 - 0x1d
      12'hFF7: dout  = 8'b11111110; // 4087 : 254 - 0xfe
      12'hFF8: dout  = 8'b00000000; // 4088 :   0 - 0x0 -- plane 1
      12'hFF9: dout  = 8'b00000000; // 4089 :   0 - 0x0
      12'hFFA: dout  = 8'b11100110; // 4090 : 230 - 0xe6
      12'hFFB: dout  = 8'b11110110; // 4091 : 246 - 0xf6
      12'hFFC: dout  = 8'b11110110; // 4092 : 246 - 0xf6
      12'hFFD: dout  = 8'b11110110; // 4093 : 246 - 0xf6
      12'hFFE: dout  = 8'b11100110; // 4094 : 230 - 0xe6
      12'hFFF: dout  = 8'b00000000; // 4095 :   0 - 0x0
    endcase
  end

endmodule
