//- Autcmatically generated verilog ROM from a NES memory file----
//-   NAME TABLE
// https://wiki.nesdev.com/w/index.php/PPU_nametables
//- Only the first Name Table: 1KiB


//-  Original memory dump file name: smario_ntable_01.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_NTABLE_SMARIO_01
  (
     //input     clk,   // clock
     input      [10-1:0] addr,  //1024 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
     //----- Name Table 0---------
      10'h0: dout  = 8'b00100100; //    0 :  36 - 0x24 -- line 0x0
      10'h1: dout  = 8'b00100100; //    1 :  36 - 0x24
      10'h2: dout  = 8'b00100100; //    2 :  36 - 0x24
      10'h3: dout  = 8'b00100100; //    3 :  36 - 0x24
      10'h4: dout  = 8'b00100100; //    4 :  36 - 0x24
      10'h5: dout  = 8'b00100100; //    5 :  36 - 0x24
      10'h6: dout  = 8'b00100100; //    6 :  36 - 0x24
      10'h7: dout  = 8'b00100100; //    7 :  36 - 0x24
      10'h8: dout  = 8'b00100100; //    8 :  36 - 0x24
      10'h9: dout  = 8'b00100100; //    9 :  36 - 0x24
      10'hA: dout  = 8'b00100100; //   10 :  36 - 0x24
      10'hB: dout  = 8'b00100100; //   11 :  36 - 0x24
      10'hC: dout  = 8'b00100100; //   12 :  36 - 0x24
      10'hD: dout  = 8'b00100100; //   13 :  36 - 0x24
      10'hE: dout  = 8'b00100100; //   14 :  36 - 0x24
      10'hF: dout  = 8'b00100100; //   15 :  36 - 0x24
      10'h10: dout  = 8'b00100100; //   16 :  36 - 0x24
      10'h11: dout  = 8'b00100100; //   17 :  36 - 0x24
      10'h12: dout  = 8'b00100100; //   18 :  36 - 0x24
      10'h13: dout  = 8'b00100100; //   19 :  36 - 0x24
      10'h14: dout  = 8'b00100100; //   20 :  36 - 0x24
      10'h15: dout  = 8'b00100100; //   21 :  36 - 0x24
      10'h16: dout  = 8'b00100100; //   22 :  36 - 0x24
      10'h17: dout  = 8'b00100100; //   23 :  36 - 0x24
      10'h18: dout  = 8'b00100100; //   24 :  36 - 0x24
      10'h19: dout  = 8'b00100100; //   25 :  36 - 0x24
      10'h1A: dout  = 8'b00100100; //   26 :  36 - 0x24
      10'h1B: dout  = 8'b00100100; //   27 :  36 - 0x24
      10'h1C: dout  = 8'b00100100; //   28 :  36 - 0x24
      10'h1D: dout  = 8'b00100100; //   29 :  36 - 0x24
      10'h1E: dout  = 8'b00100100; //   30 :  36 - 0x24
      10'h1F: dout  = 8'b00100100; //   31 :  36 - 0x24
      10'h20: dout  = 8'b00100100; //   32 :  36 - 0x24 -- line 0x1
      10'h21: dout  = 8'b00100100; //   33 :  36 - 0x24
      10'h22: dout  = 8'b00100100; //   34 :  36 - 0x24
      10'h23: dout  = 8'b00100100; //   35 :  36 - 0x24
      10'h24: dout  = 8'b00100100; //   36 :  36 - 0x24
      10'h25: dout  = 8'b00100100; //   37 :  36 - 0x24
      10'h26: dout  = 8'b00100100; //   38 :  36 - 0x24
      10'h27: dout  = 8'b00100100; //   39 :  36 - 0x24
      10'h28: dout  = 8'b00100100; //   40 :  36 - 0x24
      10'h29: dout  = 8'b00100100; //   41 :  36 - 0x24
      10'h2A: dout  = 8'b00100100; //   42 :  36 - 0x24
      10'h2B: dout  = 8'b00100100; //   43 :  36 - 0x24
      10'h2C: dout  = 8'b00100100; //   44 :  36 - 0x24
      10'h2D: dout  = 8'b00100100; //   45 :  36 - 0x24
      10'h2E: dout  = 8'b00100100; //   46 :  36 - 0x24
      10'h2F: dout  = 8'b00100100; //   47 :  36 - 0x24
      10'h30: dout  = 8'b00100100; //   48 :  36 - 0x24
      10'h31: dout  = 8'b00100100; //   49 :  36 - 0x24
      10'h32: dout  = 8'b00100100; //   50 :  36 - 0x24
      10'h33: dout  = 8'b00100100; //   51 :  36 - 0x24
      10'h34: dout  = 8'b00100100; //   52 :  36 - 0x24
      10'h35: dout  = 8'b00100100; //   53 :  36 - 0x24
      10'h36: dout  = 8'b00100100; //   54 :  36 - 0x24
      10'h37: dout  = 8'b00100100; //   55 :  36 - 0x24
      10'h38: dout  = 8'b00100100; //   56 :  36 - 0x24
      10'h39: dout  = 8'b00100100; //   57 :  36 - 0x24
      10'h3A: dout  = 8'b00100100; //   58 :  36 - 0x24
      10'h3B: dout  = 8'b00100100; //   59 :  36 - 0x24
      10'h3C: dout  = 8'b00100100; //   60 :  36 - 0x24
      10'h3D: dout  = 8'b00100100; //   61 :  36 - 0x24
      10'h3E: dout  = 8'b00100100; //   62 :  36 - 0x24
      10'h3F: dout  = 8'b00100100; //   63 :  36 - 0x24
      10'h40: dout  = 8'b00100100; //   64 :  36 - 0x24 -- line 0x2
      10'h41: dout  = 8'b00100100; //   65 :  36 - 0x24
      10'h42: dout  = 8'b00100100; //   66 :  36 - 0x24
      10'h43: dout  = 8'b00010110; //   67 :  22 - 0x16
      10'h44: dout  = 8'b00001010; //   68 :  10 - 0xa
      10'h45: dout  = 8'b00011011; //   69 :  27 - 0x1b
      10'h46: dout  = 8'b00010010; //   70 :  18 - 0x12
      10'h47: dout  = 8'b00011000; //   71 :  24 - 0x18
      10'h48: dout  = 8'b00100100; //   72 :  36 - 0x24
      10'h49: dout  = 8'b00100100; //   73 :  36 - 0x24
      10'h4A: dout  = 8'b00100100; //   74 :  36 - 0x24
      10'h4B: dout  = 8'b00100100; //   75 :  36 - 0x24
      10'h4C: dout  = 8'b00100100; //   76 :  36 - 0x24
      10'h4D: dout  = 8'b00100100; //   77 :  36 - 0x24
      10'h4E: dout  = 8'b00100100; //   78 :  36 - 0x24
      10'h4F: dout  = 8'b00100100; //   79 :  36 - 0x24
      10'h50: dout  = 8'b00100100; //   80 :  36 - 0x24
      10'h51: dout  = 8'b00100100; //   81 :  36 - 0x24
      10'h52: dout  = 8'b00100000; //   82 :  32 - 0x20
      10'h53: dout  = 8'b00011000; //   83 :  24 - 0x18
      10'h54: dout  = 8'b00011011; //   84 :  27 - 0x1b
      10'h55: dout  = 8'b00010101; //   85 :  21 - 0x15
      10'h56: dout  = 8'b00001101; //   86 :  13 - 0xd
      10'h57: dout  = 8'b00100100; //   87 :  36 - 0x24
      10'h58: dout  = 8'b00100100; //   88 :  36 - 0x24
      10'h59: dout  = 8'b00011101; //   89 :  29 - 0x1d
      10'h5A: dout  = 8'b00010010; //   90 :  18 - 0x12
      10'h5B: dout  = 8'b00010110; //   91 :  22 - 0x16
      10'h5C: dout  = 8'b00001110; //   92 :  14 - 0xe
      10'h5D: dout  = 8'b00100100; //   93 :  36 - 0x24
      10'h5E: dout  = 8'b00100100; //   94 :  36 - 0x24
      10'h5F: dout  = 8'b00100100; //   95 :  36 - 0x24
      10'h60: dout  = 8'b00100100; //   96 :  36 - 0x24 -- line 0x3
      10'h61: dout  = 8'b00100100; //   97 :  36 - 0x24
      10'h62: dout  = 8'b00100100; //   98 :  36 - 0x24
      10'h63: dout  = 8'b00000000; //   99 :   0 - 0x0
      10'h64: dout  = 8'b00000000; //  100 :   0 - 0x0
      10'h65: dout  = 8'b00000000; //  101 :   0 - 0x0
      10'h66: dout  = 8'b00000000; //  102 :   0 - 0x0
      10'h67: dout  = 8'b00000000; //  103 :   0 - 0x0
      10'h68: dout  = 8'b00000000; //  104 :   0 - 0x0
      10'h69: dout  = 8'b00100100; //  105 :  36 - 0x24
      10'h6A: dout  = 8'b00100100; //  106 :  36 - 0x24
      10'h6B: dout  = 8'b00101110; //  107 :  46 - 0x2e
      10'h6C: dout  = 8'b00101001; //  108 :  41 - 0x29
      10'h6D: dout  = 8'b00000000; //  109 :   0 - 0x0
      10'h6E: dout  = 8'b00000000; //  110 :   0 - 0x0
      10'h6F: dout  = 8'b00100100; //  111 :  36 - 0x24
      10'h70: dout  = 8'b00100100; //  112 :  36 - 0x24
      10'h71: dout  = 8'b00100100; //  113 :  36 - 0x24
      10'h72: dout  = 8'b00100100; //  114 :  36 - 0x24
      10'h73: dout  = 8'b00000001; //  115 :   1 - 0x1
      10'h74: dout  = 8'b00101000; //  116 :  40 - 0x28
      10'h75: dout  = 8'b00000001; //  117 :   1 - 0x1
      10'h76: dout  = 8'b00100100; //  118 :  36 - 0x24
      10'h77: dout  = 8'b00100100; //  119 :  36 - 0x24
      10'h78: dout  = 8'b00100100; //  120 :  36 - 0x24
      10'h79: dout  = 8'b00100100; //  121 :  36 - 0x24
      10'h7A: dout  = 8'b00100100; //  122 :  36 - 0x24
      10'h7B: dout  = 8'b00100100; //  123 :  36 - 0x24
      10'h7C: dout  = 8'b00100100; //  124 :  36 - 0x24
      10'h7D: dout  = 8'b00100100; //  125 :  36 - 0x24
      10'h7E: dout  = 8'b00100100; //  126 :  36 - 0x24
      10'h7F: dout  = 8'b00100100; //  127 :  36 - 0x24
      10'h80: dout  = 8'b00100100; //  128 :  36 - 0x24 -- line 0x4
      10'h81: dout  = 8'b00100100; //  129 :  36 - 0x24
      10'h82: dout  = 8'b00100100; //  130 :  36 - 0x24
      10'h83: dout  = 8'b00100100; //  131 :  36 - 0x24
      10'h84: dout  = 8'b00100100; //  132 :  36 - 0x24
      10'h85: dout  = 8'b01000100; //  133 :  68 - 0x44
      10'h86: dout  = 8'b01001000; //  134 :  72 - 0x48
      10'h87: dout  = 8'b01001000; //  135 :  72 - 0x48
      10'h88: dout  = 8'b01001000; //  136 :  72 - 0x48
      10'h89: dout  = 8'b01001000; //  137 :  72 - 0x48
      10'h8A: dout  = 8'b01001000; //  138 :  72 - 0x48
      10'h8B: dout  = 8'b01001000; //  139 :  72 - 0x48
      10'h8C: dout  = 8'b01001000; //  140 :  72 - 0x48
      10'h8D: dout  = 8'b01001000; //  141 :  72 - 0x48
      10'h8E: dout  = 8'b01001000; //  142 :  72 - 0x48
      10'h8F: dout  = 8'b01001000; //  143 :  72 - 0x48
      10'h90: dout  = 8'b01001000; //  144 :  72 - 0x48
      10'h91: dout  = 8'b01001000; //  145 :  72 - 0x48
      10'h92: dout  = 8'b01001000; //  146 :  72 - 0x48
      10'h93: dout  = 8'b01001000; //  147 :  72 - 0x48
      10'h94: dout  = 8'b01001000; //  148 :  72 - 0x48
      10'h95: dout  = 8'b01001000; //  149 :  72 - 0x48
      10'h96: dout  = 8'b01001000; //  150 :  72 - 0x48
      10'h97: dout  = 8'b01001000; //  151 :  72 - 0x48
      10'h98: dout  = 8'b01001000; //  152 :  72 - 0x48
      10'h99: dout  = 8'b01001000; //  153 :  72 - 0x48
      10'h9A: dout  = 8'b01001001; //  154 :  73 - 0x49
      10'h9B: dout  = 8'b00100100; //  155 :  36 - 0x24
      10'h9C: dout  = 8'b00100100; //  156 :  36 - 0x24
      10'h9D: dout  = 8'b00100100; //  157 :  36 - 0x24
      10'h9E: dout  = 8'b00100100; //  158 :  36 - 0x24
      10'h9F: dout  = 8'b00100100; //  159 :  36 - 0x24
      10'hA0: dout  = 8'b00100100; //  160 :  36 - 0x24 -- line 0x5
      10'hA1: dout  = 8'b00100100; //  161 :  36 - 0x24
      10'hA2: dout  = 8'b00100100; //  162 :  36 - 0x24
      10'hA3: dout  = 8'b00100100; //  163 :  36 - 0x24
      10'hA4: dout  = 8'b00100100; //  164 :  36 - 0x24
      10'hA5: dout  = 8'b01000110; //  165 :  70 - 0x46
      10'hA6: dout  = 8'b11010000; //  166 : 208 - 0xd0
      10'hA7: dout  = 8'b11010001; //  167 : 209 - 0xd1
      10'hA8: dout  = 8'b11011000; //  168 : 216 - 0xd8
      10'hA9: dout  = 8'b11011000; //  169 : 216 - 0xd8
      10'hAA: dout  = 8'b11011110; //  170 : 222 - 0xde
      10'hAB: dout  = 8'b11010001; //  171 : 209 - 0xd1
      10'hAC: dout  = 8'b11010000; //  172 : 208 - 0xd0
      10'hAD: dout  = 8'b11011010; //  173 : 218 - 0xda
      10'hAE: dout  = 8'b11011110; //  174 : 222 - 0xde
      10'hAF: dout  = 8'b11010001; //  175 : 209 - 0xd1
      10'hB0: dout  = 8'b00100110; //  176 :  38 - 0x26
      10'hB1: dout  = 8'b00100110; //  177 :  38 - 0x26
      10'hB2: dout  = 8'b00100110; //  178 :  38 - 0x26
      10'hB3: dout  = 8'b00100110; //  179 :  38 - 0x26
      10'hB4: dout  = 8'b00100110; //  180 :  38 - 0x26
      10'hB5: dout  = 8'b00100110; //  181 :  38 - 0x26
      10'hB6: dout  = 8'b00100110; //  182 :  38 - 0x26
      10'hB7: dout  = 8'b00100110; //  183 :  38 - 0x26
      10'hB8: dout  = 8'b00100110; //  184 :  38 - 0x26
      10'hB9: dout  = 8'b00100110; //  185 :  38 - 0x26
      10'hBA: dout  = 8'b01001010; //  186 :  74 - 0x4a
      10'hBB: dout  = 8'b00100100; //  187 :  36 - 0x24
      10'hBC: dout  = 8'b00100100; //  188 :  36 - 0x24
      10'hBD: dout  = 8'b00100100; //  189 :  36 - 0x24
      10'hBE: dout  = 8'b00100100; //  190 :  36 - 0x24
      10'hBF: dout  = 8'b00100100; //  191 :  36 - 0x24
      10'hC0: dout  = 8'b00100100; //  192 :  36 - 0x24 -- line 0x6
      10'hC1: dout  = 8'b00100100; //  193 :  36 - 0x24
      10'hC2: dout  = 8'b00100100; //  194 :  36 - 0x24
      10'hC3: dout  = 8'b00100100; //  195 :  36 - 0x24
      10'hC4: dout  = 8'b00100100; //  196 :  36 - 0x24
      10'hC5: dout  = 8'b01000110; //  197 :  70 - 0x46
      10'hC6: dout  = 8'b11010010; //  198 : 210 - 0xd2
      10'hC7: dout  = 8'b11010011; //  199 : 211 - 0xd3
      10'hC8: dout  = 8'b11011011; //  200 : 219 - 0xdb
      10'hC9: dout  = 8'b11011011; //  201 : 219 - 0xdb
      10'hCA: dout  = 8'b11011011; //  202 : 219 - 0xdb
      10'hCB: dout  = 8'b11011001; //  203 : 217 - 0xd9
      10'hCC: dout  = 8'b11011011; //  204 : 219 - 0xdb
      10'hCD: dout  = 8'b11011100; //  205 : 220 - 0xdc
      10'hCE: dout  = 8'b11011011; //  206 : 219 - 0xdb
      10'hCF: dout  = 8'b11011111; //  207 : 223 - 0xdf
      10'hD0: dout  = 8'b00100110; //  208 :  38 - 0x26
      10'hD1: dout  = 8'b00100110; //  209 :  38 - 0x26
      10'hD2: dout  = 8'b00100110; //  210 :  38 - 0x26
      10'hD3: dout  = 8'b00100110; //  211 :  38 - 0x26
      10'hD4: dout  = 8'b00100110; //  212 :  38 - 0x26
      10'hD5: dout  = 8'b00100110; //  213 :  38 - 0x26
      10'hD6: dout  = 8'b00100110; //  214 :  38 - 0x26
      10'hD7: dout  = 8'b00100110; //  215 :  38 - 0x26
      10'hD8: dout  = 8'b00100110; //  216 :  38 - 0x26
      10'hD9: dout  = 8'b00100110; //  217 :  38 - 0x26
      10'hDA: dout  = 8'b01001010; //  218 :  74 - 0x4a
      10'hDB: dout  = 8'b00100100; //  219 :  36 - 0x24
      10'hDC: dout  = 8'b00100100; //  220 :  36 - 0x24
      10'hDD: dout  = 8'b00100100; //  221 :  36 - 0x24
      10'hDE: dout  = 8'b00100100; //  222 :  36 - 0x24
      10'hDF: dout  = 8'b00100100; //  223 :  36 - 0x24
      10'hE0: dout  = 8'b00100100; //  224 :  36 - 0x24 -- line 0x7
      10'hE1: dout  = 8'b00100100; //  225 :  36 - 0x24
      10'hE2: dout  = 8'b00100100; //  226 :  36 - 0x24
      10'hE3: dout  = 8'b00100100; //  227 :  36 - 0x24
      10'hE4: dout  = 8'b00100100; //  228 :  36 - 0x24
      10'hE5: dout  = 8'b01000110; //  229 :  70 - 0x46
      10'hE6: dout  = 8'b11010100; //  230 : 212 - 0xd4
      10'hE7: dout  = 8'b11010101; //  231 : 213 - 0xd5
      10'hE8: dout  = 8'b11010100; //  232 : 212 - 0xd4
      10'hE9: dout  = 8'b11011001; //  233 : 217 - 0xd9
      10'hEA: dout  = 8'b11011011; //  234 : 219 - 0xdb
      10'hEB: dout  = 8'b11100010; //  235 : 226 - 0xe2
      10'hEC: dout  = 8'b11010100; //  236 : 212 - 0xd4
      10'hED: dout  = 8'b11011010; //  237 : 218 - 0xda
      10'hEE: dout  = 8'b11011011; //  238 : 219 - 0xdb
      10'hEF: dout  = 8'b11100000; //  239 : 224 - 0xe0
      10'hF0: dout  = 8'b00100110; //  240 :  38 - 0x26
      10'hF1: dout  = 8'b00100110; //  241 :  38 - 0x26
      10'hF2: dout  = 8'b00100110; //  242 :  38 - 0x26
      10'hF3: dout  = 8'b00100110; //  243 :  38 - 0x26
      10'hF4: dout  = 8'b00100110; //  244 :  38 - 0x26
      10'hF5: dout  = 8'b00100110; //  245 :  38 - 0x26
      10'hF6: dout  = 8'b00100110; //  246 :  38 - 0x26
      10'hF7: dout  = 8'b00100110; //  247 :  38 - 0x26
      10'hF8: dout  = 8'b00100110; //  248 :  38 - 0x26
      10'hF9: dout  = 8'b00100110; //  249 :  38 - 0x26
      10'hFA: dout  = 8'b01001010; //  250 :  74 - 0x4a
      10'hFB: dout  = 8'b00100100; //  251 :  36 - 0x24
      10'hFC: dout  = 8'b00100100; //  252 :  36 - 0x24
      10'hFD: dout  = 8'b00100100; //  253 :  36 - 0x24
      10'hFE: dout  = 8'b00100100; //  254 :  36 - 0x24
      10'hFF: dout  = 8'b00100100; //  255 :  36 - 0x24
      10'h100: dout  = 8'b00100100; //  256 :  36 - 0x24 -- line 0x8
      10'h101: dout  = 8'b00100100; //  257 :  36 - 0x24
      10'h102: dout  = 8'b00100100; //  258 :  36 - 0x24
      10'h103: dout  = 8'b00100100; //  259 :  36 - 0x24
      10'h104: dout  = 8'b00100100; //  260 :  36 - 0x24
      10'h105: dout  = 8'b01000110; //  261 :  70 - 0x46
      10'h106: dout  = 8'b11010110; //  262 : 214 - 0xd6
      10'h107: dout  = 8'b11010111; //  263 : 215 - 0xd7
      10'h108: dout  = 8'b11010110; //  264 : 214 - 0xd6
      10'h109: dout  = 8'b11010111; //  265 : 215 - 0xd7
      10'h10A: dout  = 8'b11100001; //  266 : 225 - 0xe1
      10'h10B: dout  = 8'b00100110; //  267 :  38 - 0x26
      10'h10C: dout  = 8'b11010110; //  268 : 214 - 0xd6
      10'h10D: dout  = 8'b11011101; //  269 : 221 - 0xdd
      10'h10E: dout  = 8'b11100001; //  270 : 225 - 0xe1
      10'h10F: dout  = 8'b11100001; //  271 : 225 - 0xe1
      10'h110: dout  = 8'b00100110; //  272 :  38 - 0x26
      10'h111: dout  = 8'b00100110; //  273 :  38 - 0x26
      10'h112: dout  = 8'b00100110; //  274 :  38 - 0x26
      10'h113: dout  = 8'b00100110; //  275 :  38 - 0x26
      10'h114: dout  = 8'b00100110; //  276 :  38 - 0x26
      10'h115: dout  = 8'b00100110; //  277 :  38 - 0x26
      10'h116: dout  = 8'b00100110; //  278 :  38 - 0x26
      10'h117: dout  = 8'b00100110; //  279 :  38 - 0x26
      10'h118: dout  = 8'b00100110; //  280 :  38 - 0x26
      10'h119: dout  = 8'b00100110; //  281 :  38 - 0x26
      10'h11A: dout  = 8'b01001010; //  282 :  74 - 0x4a
      10'h11B: dout  = 8'b00100100; //  283 :  36 - 0x24
      10'h11C: dout  = 8'b00100100; //  284 :  36 - 0x24
      10'h11D: dout  = 8'b00100100; //  285 :  36 - 0x24
      10'h11E: dout  = 8'b00100100; //  286 :  36 - 0x24
      10'h11F: dout  = 8'b00100100; //  287 :  36 - 0x24
      10'h120: dout  = 8'b00100100; //  288 :  36 - 0x24 -- line 0x9
      10'h121: dout  = 8'b00100100; //  289 :  36 - 0x24
      10'h122: dout  = 8'b00100100; //  290 :  36 - 0x24
      10'h123: dout  = 8'b00100100; //  291 :  36 - 0x24
      10'h124: dout  = 8'b00100100; //  292 :  36 - 0x24
      10'h125: dout  = 8'b01000110; //  293 :  70 - 0x46
      10'h126: dout  = 8'b11010000; //  294 : 208 - 0xd0
      10'h127: dout  = 8'b11101000; //  295 : 232 - 0xe8
      10'h128: dout  = 8'b11010001; //  296 : 209 - 0xd1
      10'h129: dout  = 8'b11010000; //  297 : 208 - 0xd0
      10'h12A: dout  = 8'b11010001; //  298 : 209 - 0xd1
      10'h12B: dout  = 8'b11011110; //  299 : 222 - 0xde
      10'h12C: dout  = 8'b11010001; //  300 : 209 - 0xd1
      10'h12D: dout  = 8'b11011000; //  301 : 216 - 0xd8
      10'h12E: dout  = 8'b11010000; //  302 : 208 - 0xd0
      10'h12F: dout  = 8'b11010001; //  303 : 209 - 0xd1
      10'h130: dout  = 8'b00100110; //  304 :  38 - 0x26
      10'h131: dout  = 8'b11011110; //  305 : 222 - 0xde
      10'h132: dout  = 8'b11010001; //  306 : 209 - 0xd1
      10'h133: dout  = 8'b11011110; //  307 : 222 - 0xde
      10'h134: dout  = 8'b11010001; //  308 : 209 - 0xd1
      10'h135: dout  = 8'b11010000; //  309 : 208 - 0xd0
      10'h136: dout  = 8'b11010001; //  310 : 209 - 0xd1
      10'h137: dout  = 8'b11010000; //  311 : 208 - 0xd0
      10'h138: dout  = 8'b11010001; //  312 : 209 - 0xd1
      10'h139: dout  = 8'b00100110; //  313 :  38 - 0x26
      10'h13A: dout  = 8'b01001010; //  314 :  74 - 0x4a
      10'h13B: dout  = 8'b00100100; //  315 :  36 - 0x24
      10'h13C: dout  = 8'b00100100; //  316 :  36 - 0x24
      10'h13D: dout  = 8'b00100100; //  317 :  36 - 0x24
      10'h13E: dout  = 8'b00100100; //  318 :  36 - 0x24
      10'h13F: dout  = 8'b00100100; //  319 :  36 - 0x24
      10'h140: dout  = 8'b00100100; //  320 :  36 - 0x24 -- line 0xa
      10'h141: dout  = 8'b00100100; //  321 :  36 - 0x24
      10'h142: dout  = 8'b00100100; //  322 :  36 - 0x24
      10'h143: dout  = 8'b00100100; //  323 :  36 - 0x24
      10'h144: dout  = 8'b00100100; //  324 :  36 - 0x24
      10'h145: dout  = 8'b01000110; //  325 :  70 - 0x46
      10'h146: dout  = 8'b11011011; //  326 : 219 - 0xdb
      10'h147: dout  = 8'b01000010; //  327 :  66 - 0x42
      10'h148: dout  = 8'b01000010; //  328 :  66 - 0x42
      10'h149: dout  = 8'b11011011; //  329 : 219 - 0xdb
      10'h14A: dout  = 8'b01000010; //  330 :  66 - 0x42
      10'h14B: dout  = 8'b11011011; //  331 : 219 - 0xdb
      10'h14C: dout  = 8'b01000010; //  332 :  66 - 0x42
      10'h14D: dout  = 8'b11011011; //  333 : 219 - 0xdb
      10'h14E: dout  = 8'b11011011; //  334 : 219 - 0xdb
      10'h14F: dout  = 8'b01000010; //  335 :  66 - 0x42
      10'h150: dout  = 8'b00100110; //  336 :  38 - 0x26
      10'h151: dout  = 8'b11011011; //  337 : 219 - 0xdb
      10'h152: dout  = 8'b01000010; //  338 :  66 - 0x42
      10'h153: dout  = 8'b11011011; //  339 : 219 - 0xdb
      10'h154: dout  = 8'b01000010; //  340 :  66 - 0x42
      10'h155: dout  = 8'b11011011; //  341 : 219 - 0xdb
      10'h156: dout  = 8'b01000010; //  342 :  66 - 0x42
      10'h157: dout  = 8'b11011011; //  343 : 219 - 0xdb
      10'h158: dout  = 8'b01000010; //  344 :  66 - 0x42
      10'h159: dout  = 8'b00100110; //  345 :  38 - 0x26
      10'h15A: dout  = 8'b01001010; //  346 :  74 - 0x4a
      10'h15B: dout  = 8'b00100100; //  347 :  36 - 0x24
      10'h15C: dout  = 8'b00100100; //  348 :  36 - 0x24
      10'h15D: dout  = 8'b00100100; //  349 :  36 - 0x24
      10'h15E: dout  = 8'b00100100; //  350 :  36 - 0x24
      10'h15F: dout  = 8'b00100100; //  351 :  36 - 0x24
      10'h160: dout  = 8'b00100100; //  352 :  36 - 0x24 -- line 0xb
      10'h161: dout  = 8'b00100100; //  353 :  36 - 0x24
      10'h162: dout  = 8'b00100100; //  354 :  36 - 0x24
      10'h163: dout  = 8'b00100100; //  355 :  36 - 0x24
      10'h164: dout  = 8'b00100100; //  356 :  36 - 0x24
      10'h165: dout  = 8'b01000110; //  357 :  70 - 0x46
      10'h166: dout  = 8'b11011011; //  358 : 219 - 0xdb
      10'h167: dout  = 8'b11011011; //  359 : 219 - 0xdb
      10'h168: dout  = 8'b11011011; //  360 : 219 - 0xdb
      10'h169: dout  = 8'b11011011; //  361 : 219 - 0xdb
      10'h16A: dout  = 8'b11011011; //  362 : 219 - 0xdb
      10'h16B: dout  = 8'b11011011; //  363 : 219 - 0xdb
      10'h16C: dout  = 8'b11011111; //  364 : 223 - 0xdf
      10'h16D: dout  = 8'b11011011; //  365 : 219 - 0xdb
      10'h16E: dout  = 8'b11011011; //  366 : 219 - 0xdb
      10'h16F: dout  = 8'b11011011; //  367 : 219 - 0xdb
      10'h170: dout  = 8'b00100110; //  368 :  38 - 0x26
      10'h171: dout  = 8'b11011011; //  369 : 219 - 0xdb
      10'h172: dout  = 8'b11011111; //  370 : 223 - 0xdf
      10'h173: dout  = 8'b11011011; //  371 : 219 - 0xdb
      10'h174: dout  = 8'b11011111; //  372 : 223 - 0xdf
      10'h175: dout  = 8'b11011011; //  373 : 219 - 0xdb
      10'h176: dout  = 8'b11011011; //  374 : 219 - 0xdb
      10'h177: dout  = 8'b11100100; //  375 : 228 - 0xe4
      10'h178: dout  = 8'b11100101; //  376 : 229 - 0xe5
      10'h179: dout  = 8'b00100110; //  377 :  38 - 0x26
      10'h17A: dout  = 8'b01001010; //  378 :  74 - 0x4a
      10'h17B: dout  = 8'b00100100; //  379 :  36 - 0x24
      10'h17C: dout  = 8'b00100100; //  380 :  36 - 0x24
      10'h17D: dout  = 8'b00100100; //  381 :  36 - 0x24
      10'h17E: dout  = 8'b00100100; //  382 :  36 - 0x24
      10'h17F: dout  = 8'b00100100; //  383 :  36 - 0x24
      10'h180: dout  = 8'b00100100; //  384 :  36 - 0x24 -- line 0xc
      10'h181: dout  = 8'b00100100; //  385 :  36 - 0x24
      10'h182: dout  = 8'b00100100; //  386 :  36 - 0x24
      10'h183: dout  = 8'b00100100; //  387 :  36 - 0x24
      10'h184: dout  = 8'b00100100; //  388 :  36 - 0x24
      10'h185: dout  = 8'b01000110; //  389 :  70 - 0x46
      10'h186: dout  = 8'b11011011; //  390 : 219 - 0xdb
      10'h187: dout  = 8'b11011011; //  391 : 219 - 0xdb
      10'h188: dout  = 8'b11011011; //  392 : 219 - 0xdb
      10'h189: dout  = 8'b11011110; //  393 : 222 - 0xde
      10'h18A: dout  = 8'b01000011; //  394 :  67 - 0x43
      10'h18B: dout  = 8'b11011011; //  395 : 219 - 0xdb
      10'h18C: dout  = 8'b11100000; //  396 : 224 - 0xe0
      10'h18D: dout  = 8'b11011011; //  397 : 219 - 0xdb
      10'h18E: dout  = 8'b11011011; //  398 : 219 - 0xdb
      10'h18F: dout  = 8'b11011011; //  399 : 219 - 0xdb
      10'h190: dout  = 8'b00100110; //  400 :  38 - 0x26
      10'h191: dout  = 8'b11011011; //  401 : 219 - 0xdb
      10'h192: dout  = 8'b11100011; //  402 : 227 - 0xe3
      10'h193: dout  = 8'b11011011; //  403 : 219 - 0xdb
      10'h194: dout  = 8'b11100000; //  404 : 224 - 0xe0
      10'h195: dout  = 8'b11011011; //  405 : 219 - 0xdb
      10'h196: dout  = 8'b11011011; //  406 : 219 - 0xdb
      10'h197: dout  = 8'b11100110; //  407 : 230 - 0xe6
      10'h198: dout  = 8'b11100011; //  408 : 227 - 0xe3
      10'h199: dout  = 8'b00100110; //  409 :  38 - 0x26
      10'h19A: dout  = 8'b01001010; //  410 :  74 - 0x4a
      10'h19B: dout  = 8'b00100100; //  411 :  36 - 0x24
      10'h19C: dout  = 8'b00100100; //  412 :  36 - 0x24
      10'h19D: dout  = 8'b00100100; //  413 :  36 - 0x24
      10'h19E: dout  = 8'b00100100; //  414 :  36 - 0x24
      10'h19F: dout  = 8'b00100100; //  415 :  36 - 0x24
      10'h1A0: dout  = 8'b00100100; //  416 :  36 - 0x24 -- line 0xd
      10'h1A1: dout  = 8'b00100100; //  417 :  36 - 0x24
      10'h1A2: dout  = 8'b00100100; //  418 :  36 - 0x24
      10'h1A3: dout  = 8'b00100100; //  419 :  36 - 0x24
      10'h1A4: dout  = 8'b00100100; //  420 :  36 - 0x24
      10'h1A5: dout  = 8'b01000110; //  421 :  70 - 0x46
      10'h1A6: dout  = 8'b11011011; //  422 : 219 - 0xdb
      10'h1A7: dout  = 8'b11011011; //  423 : 219 - 0xdb
      10'h1A8: dout  = 8'b11011011; //  424 : 219 - 0xdb
      10'h1A9: dout  = 8'b11011011; //  425 : 219 - 0xdb
      10'h1AA: dout  = 8'b01000010; //  426 :  66 - 0x42
      10'h1AB: dout  = 8'b11011011; //  427 : 219 - 0xdb
      10'h1AC: dout  = 8'b11011011; //  428 : 219 - 0xdb
      10'h1AD: dout  = 8'b11011011; //  429 : 219 - 0xdb
      10'h1AE: dout  = 8'b11010100; //  430 : 212 - 0xd4
      10'h1AF: dout  = 8'b11011001; //  431 : 217 - 0xd9
      10'h1B0: dout  = 8'b00100110; //  432 :  38 - 0x26
      10'h1B1: dout  = 8'b11011011; //  433 : 219 - 0xdb
      10'h1B2: dout  = 8'b11011001; //  434 : 217 - 0xd9
      10'h1B3: dout  = 8'b11011011; //  435 : 219 - 0xdb
      10'h1B4: dout  = 8'b11011011; //  436 : 219 - 0xdb
      10'h1B5: dout  = 8'b11010100; //  437 : 212 - 0xd4
      10'h1B6: dout  = 8'b11011001; //  438 : 217 - 0xd9
      10'h1B7: dout  = 8'b11010100; //  439 : 212 - 0xd4
      10'h1B8: dout  = 8'b11011001; //  440 : 217 - 0xd9
      10'h1B9: dout  = 8'b11100111; //  441 : 231 - 0xe7
      10'h1BA: dout  = 8'b01001010; //  442 :  74 - 0x4a
      10'h1BB: dout  = 8'b00100100; //  443 :  36 - 0x24
      10'h1BC: dout  = 8'b00100100; //  444 :  36 - 0x24
      10'h1BD: dout  = 8'b00100100; //  445 :  36 - 0x24
      10'h1BE: dout  = 8'b00100100; //  446 :  36 - 0x24
      10'h1BF: dout  = 8'b00100100; //  447 :  36 - 0x24
      10'h1C0: dout  = 8'b00100100; //  448 :  36 - 0x24 -- line 0xe
      10'h1C1: dout  = 8'b00100100; //  449 :  36 - 0x24
      10'h1C2: dout  = 8'b00100100; //  450 :  36 - 0x24
      10'h1C3: dout  = 8'b00100100; //  451 :  36 - 0x24
      10'h1C4: dout  = 8'b00100100; //  452 :  36 - 0x24
      10'h1C5: dout  = 8'b01011111; //  453 :  95 - 0x5f
      10'h1C6: dout  = 8'b10010101; //  454 : 149 - 0x95
      10'h1C7: dout  = 8'b10010101; //  455 : 149 - 0x95
      10'h1C8: dout  = 8'b10010101; //  456 : 149 - 0x95
      10'h1C9: dout  = 8'b10010101; //  457 : 149 - 0x95
      10'h1CA: dout  = 8'b10010101; //  458 : 149 - 0x95
      10'h1CB: dout  = 8'b10010101; //  459 : 149 - 0x95
      10'h1CC: dout  = 8'b10010101; //  460 : 149 - 0x95
      10'h1CD: dout  = 8'b10010101; //  461 : 149 - 0x95
      10'h1CE: dout  = 8'b10010111; //  462 : 151 - 0x97
      10'h1CF: dout  = 8'b10011000; //  463 : 152 - 0x98
      10'h1D0: dout  = 8'b01111000; //  464 : 120 - 0x78
      10'h1D1: dout  = 8'b10010101; //  465 : 149 - 0x95
      10'h1D2: dout  = 8'b10010110; //  466 : 150 - 0x96
      10'h1D3: dout  = 8'b10010101; //  467 : 149 - 0x95
      10'h1D4: dout  = 8'b10010101; //  468 : 149 - 0x95
      10'h1D5: dout  = 8'b10010111; //  469 : 151 - 0x97
      10'h1D6: dout  = 8'b10011000; //  470 : 152 - 0x98
      10'h1D7: dout  = 8'b10010111; //  471 : 151 - 0x97
      10'h1D8: dout  = 8'b10011000; //  472 : 152 - 0x98
      10'h1D9: dout  = 8'b10010101; //  473 : 149 - 0x95
      10'h1DA: dout  = 8'b01111010; //  474 : 122 - 0x7a
      10'h1DB: dout  = 8'b00100100; //  475 :  36 - 0x24
      10'h1DC: dout  = 8'b00100100; //  476 :  36 - 0x24
      10'h1DD: dout  = 8'b00100100; //  477 :  36 - 0x24
      10'h1DE: dout  = 8'b00100100; //  478 :  36 - 0x24
      10'h1DF: dout  = 8'b00100100; //  479 :  36 - 0x24
      10'h1E0: dout  = 8'b00100100; //  480 :  36 - 0x24 -- line 0xf
      10'h1E1: dout  = 8'b00100100; //  481 :  36 - 0x24
      10'h1E2: dout  = 8'b00100100; //  482 :  36 - 0x24
      10'h1E3: dout  = 8'b00100100; //  483 :  36 - 0x24
      10'h1E4: dout  = 8'b00100100; //  484 :  36 - 0x24
      10'h1E5: dout  = 8'b00100100; //  485 :  36 - 0x24
      10'h1E6: dout  = 8'b00100100; //  486 :  36 - 0x24
      10'h1E7: dout  = 8'b00100100; //  487 :  36 - 0x24
      10'h1E8: dout  = 8'b00100100; //  488 :  36 - 0x24
      10'h1E9: dout  = 8'b00100100; //  489 :  36 - 0x24
      10'h1EA: dout  = 8'b00100100; //  490 :  36 - 0x24
      10'h1EB: dout  = 8'b00100100; //  491 :  36 - 0x24
      10'h1EC: dout  = 8'b00100100; //  492 :  36 - 0x24
      10'h1ED: dout  = 8'b11001111; //  493 : 207 - 0xcf
      10'h1EE: dout  = 8'b00000001; //  494 :   1 - 0x1
      10'h1EF: dout  = 8'b00001001; //  495 :   9 - 0x9
      10'h1F0: dout  = 8'b00001000; //  496 :   8 - 0x8
      10'h1F1: dout  = 8'b00000101; //  497 :   5 - 0x5
      10'h1F2: dout  = 8'b00100100; //  498 :  36 - 0x24
      10'h1F3: dout  = 8'b00010111; //  499 :  23 - 0x17
      10'h1F4: dout  = 8'b00010010; //  500 :  18 - 0x12
      10'h1F5: dout  = 8'b00010111; //  501 :  23 - 0x17
      10'h1F6: dout  = 8'b00011101; //  502 :  29 - 0x1d
      10'h1F7: dout  = 8'b00001110; //  503 :  14 - 0xe
      10'h1F8: dout  = 8'b00010111; //  504 :  23 - 0x17
      10'h1F9: dout  = 8'b00001101; //  505 :  13 - 0xd
      10'h1FA: dout  = 8'b00011000; //  506 :  24 - 0x18
      10'h1FB: dout  = 8'b00100100; //  507 :  36 - 0x24
      10'h1FC: dout  = 8'b00100100; //  508 :  36 - 0x24
      10'h1FD: dout  = 8'b00100100; //  509 :  36 - 0x24
      10'h1FE: dout  = 8'b00100100; //  510 :  36 - 0x24
      10'h1FF: dout  = 8'b00100100; //  511 :  36 - 0x24
      10'h200: dout  = 8'b00100100; //  512 :  36 - 0x24 -- line 0x10
      10'h201: dout  = 8'b00100100; //  513 :  36 - 0x24
      10'h202: dout  = 8'b00100100; //  514 :  36 - 0x24
      10'h203: dout  = 8'b00100100; //  515 :  36 - 0x24
      10'h204: dout  = 8'b00100100; //  516 :  36 - 0x24
      10'h205: dout  = 8'b00100100; //  517 :  36 - 0x24
      10'h206: dout  = 8'b00100100; //  518 :  36 - 0x24
      10'h207: dout  = 8'b00100100; //  519 :  36 - 0x24
      10'h208: dout  = 8'b00100100; //  520 :  36 - 0x24
      10'h209: dout  = 8'b00100100; //  521 :  36 - 0x24
      10'h20A: dout  = 8'b00100100; //  522 :  36 - 0x24
      10'h20B: dout  = 8'b00100100; //  523 :  36 - 0x24
      10'h20C: dout  = 8'b00100100; //  524 :  36 - 0x24
      10'h20D: dout  = 8'b00100100; //  525 :  36 - 0x24
      10'h20E: dout  = 8'b00100100; //  526 :  36 - 0x24
      10'h20F: dout  = 8'b00100100; //  527 :  36 - 0x24
      10'h210: dout  = 8'b00100100; //  528 :  36 - 0x24
      10'h211: dout  = 8'b00100100; //  529 :  36 - 0x24
      10'h212: dout  = 8'b00100100; //  530 :  36 - 0x24
      10'h213: dout  = 8'b00100100; //  531 :  36 - 0x24
      10'h214: dout  = 8'b00100100; //  532 :  36 - 0x24
      10'h215: dout  = 8'b00100100; //  533 :  36 - 0x24
      10'h216: dout  = 8'b00100100; //  534 :  36 - 0x24
      10'h217: dout  = 8'b00100100; //  535 :  36 - 0x24
      10'h218: dout  = 8'b00100100; //  536 :  36 - 0x24
      10'h219: dout  = 8'b00100100; //  537 :  36 - 0x24
      10'h21A: dout  = 8'b00100100; //  538 :  36 - 0x24
      10'h21B: dout  = 8'b00100100; //  539 :  36 - 0x24
      10'h21C: dout  = 8'b00100100; //  540 :  36 - 0x24
      10'h21D: dout  = 8'b00100100; //  541 :  36 - 0x24
      10'h21E: dout  = 8'b00100100; //  542 :  36 - 0x24
      10'h21F: dout  = 8'b00100100; //  543 :  36 - 0x24
      10'h220: dout  = 8'b00100100; //  544 :  36 - 0x24 -- line 0x11
      10'h221: dout  = 8'b00100100; //  545 :  36 - 0x24
      10'h222: dout  = 8'b00100100; //  546 :  36 - 0x24
      10'h223: dout  = 8'b00100100; //  547 :  36 - 0x24
      10'h224: dout  = 8'b00100100; //  548 :  36 - 0x24
      10'h225: dout  = 8'b00100100; //  549 :  36 - 0x24
      10'h226: dout  = 8'b00100100; //  550 :  36 - 0x24
      10'h227: dout  = 8'b00100100; //  551 :  36 - 0x24
      10'h228: dout  = 8'b00100100; //  552 :  36 - 0x24
      10'h229: dout  = 8'b00100100; //  553 :  36 - 0x24
      10'h22A: dout  = 8'b00100100; //  554 :  36 - 0x24
      10'h22B: dout  = 8'b00100100; //  555 :  36 - 0x24
      10'h22C: dout  = 8'b00100100; //  556 :  36 - 0x24
      10'h22D: dout  = 8'b00100100; //  557 :  36 - 0x24
      10'h22E: dout  = 8'b00100100; //  558 :  36 - 0x24
      10'h22F: dout  = 8'b00100100; //  559 :  36 - 0x24
      10'h230: dout  = 8'b00100100; //  560 :  36 - 0x24
      10'h231: dout  = 8'b00100100; //  561 :  36 - 0x24
      10'h232: dout  = 8'b00100100; //  562 :  36 - 0x24
      10'h233: dout  = 8'b00100100; //  563 :  36 - 0x24
      10'h234: dout  = 8'b00100100; //  564 :  36 - 0x24
      10'h235: dout  = 8'b00100100; //  565 :  36 - 0x24
      10'h236: dout  = 8'b00100100; //  566 :  36 - 0x24
      10'h237: dout  = 8'b00100100; //  567 :  36 - 0x24
      10'h238: dout  = 8'b00100100; //  568 :  36 - 0x24
      10'h239: dout  = 8'b00100100; //  569 :  36 - 0x24
      10'h23A: dout  = 8'b00100100; //  570 :  36 - 0x24
      10'h23B: dout  = 8'b00100100; //  571 :  36 - 0x24
      10'h23C: dout  = 8'b00100100; //  572 :  36 - 0x24
      10'h23D: dout  = 8'b00100100; //  573 :  36 - 0x24
      10'h23E: dout  = 8'b00100100; //  574 :  36 - 0x24
      10'h23F: dout  = 8'b00100100; //  575 :  36 - 0x24
      10'h240: dout  = 8'b00100100; //  576 :  36 - 0x24 -- line 0x12
      10'h241: dout  = 8'b00100100; //  577 :  36 - 0x24
      10'h242: dout  = 8'b00100100; //  578 :  36 - 0x24
      10'h243: dout  = 8'b00100100; //  579 :  36 - 0x24
      10'h244: dout  = 8'b00100100; //  580 :  36 - 0x24
      10'h245: dout  = 8'b00100100; //  581 :  36 - 0x24
      10'h246: dout  = 8'b00100100; //  582 :  36 - 0x24
      10'h247: dout  = 8'b00100100; //  583 :  36 - 0x24
      10'h248: dout  = 8'b00100100; //  584 :  36 - 0x24
      10'h249: dout  = 8'b11001110; //  585 : 206 - 0xce
      10'h24A: dout  = 8'b00100100; //  586 :  36 - 0x24
      10'h24B: dout  = 8'b00000001; //  587 :   1 - 0x1
      10'h24C: dout  = 8'b00100100; //  588 :  36 - 0x24
      10'h24D: dout  = 8'b00011001; //  589 :  25 - 0x19
      10'h24E: dout  = 8'b00010101; //  590 :  21 - 0x15
      10'h24F: dout  = 8'b00001010; //  591 :  10 - 0xa
      10'h250: dout  = 8'b00100010; //  592 :  34 - 0x22
      10'h251: dout  = 8'b00001110; //  593 :  14 - 0xe
      10'h252: dout  = 8'b00011011; //  594 :  27 - 0x1b
      10'h253: dout  = 8'b00100100; //  595 :  36 - 0x24
      10'h254: dout  = 8'b00010000; //  596 :  16 - 0x10
      10'h255: dout  = 8'b00001010; //  597 :  10 - 0xa
      10'h256: dout  = 8'b00010110; //  598 :  22 - 0x16
      10'h257: dout  = 8'b00001110; //  599 :  14 - 0xe
      10'h258: dout  = 8'b00100100; //  600 :  36 - 0x24
      10'h259: dout  = 8'b00100100; //  601 :  36 - 0x24
      10'h25A: dout  = 8'b00100100; //  602 :  36 - 0x24
      10'h25B: dout  = 8'b00100100; //  603 :  36 - 0x24
      10'h25C: dout  = 8'b00100100; //  604 :  36 - 0x24
      10'h25D: dout  = 8'b00100100; //  605 :  36 - 0x24
      10'h25E: dout  = 8'b00100100; //  606 :  36 - 0x24
      10'h25F: dout  = 8'b00100100; //  607 :  36 - 0x24
      10'h260: dout  = 8'b00100100; //  608 :  36 - 0x24 -- line 0x13
      10'h261: dout  = 8'b00100100; //  609 :  36 - 0x24
      10'h262: dout  = 8'b00100100; //  610 :  36 - 0x24
      10'h263: dout  = 8'b00100100; //  611 :  36 - 0x24
      10'h264: dout  = 8'b00100100; //  612 :  36 - 0x24
      10'h265: dout  = 8'b00100100; //  613 :  36 - 0x24
      10'h266: dout  = 8'b00100100; //  614 :  36 - 0x24
      10'h267: dout  = 8'b00100100; //  615 :  36 - 0x24
      10'h268: dout  = 8'b00100100; //  616 :  36 - 0x24
      10'h269: dout  = 8'b00100100; //  617 :  36 - 0x24
      10'h26A: dout  = 8'b00100100; //  618 :  36 - 0x24
      10'h26B: dout  = 8'b00100100; //  619 :  36 - 0x24
      10'h26C: dout  = 8'b00100100; //  620 :  36 - 0x24
      10'h26D: dout  = 8'b00100100; //  621 :  36 - 0x24
      10'h26E: dout  = 8'b00100100; //  622 :  36 - 0x24
      10'h26F: dout  = 8'b00100100; //  623 :  36 - 0x24
      10'h270: dout  = 8'b00100100; //  624 :  36 - 0x24
      10'h271: dout  = 8'b00100100; //  625 :  36 - 0x24
      10'h272: dout  = 8'b00100100; //  626 :  36 - 0x24
      10'h273: dout  = 8'b00100100; //  627 :  36 - 0x24
      10'h274: dout  = 8'b00100100; //  628 :  36 - 0x24
      10'h275: dout  = 8'b00100100; //  629 :  36 - 0x24
      10'h276: dout  = 8'b00100100; //  630 :  36 - 0x24
      10'h277: dout  = 8'b00100100; //  631 :  36 - 0x24
      10'h278: dout  = 8'b00100100; //  632 :  36 - 0x24
      10'h279: dout  = 8'b00100100; //  633 :  36 - 0x24
      10'h27A: dout  = 8'b00100100; //  634 :  36 - 0x24
      10'h27B: dout  = 8'b00100100; //  635 :  36 - 0x24
      10'h27C: dout  = 8'b00100100; //  636 :  36 - 0x24
      10'h27D: dout  = 8'b00100100; //  637 :  36 - 0x24
      10'h27E: dout  = 8'b00100100; //  638 :  36 - 0x24
      10'h27F: dout  = 8'b00100100; //  639 :  36 - 0x24
      10'h280: dout  = 8'b00100100; //  640 :  36 - 0x24 -- line 0x14
      10'h281: dout  = 8'b00100100; //  641 :  36 - 0x24
      10'h282: dout  = 8'b00100100; //  642 :  36 - 0x24
      10'h283: dout  = 8'b00100100; //  643 :  36 - 0x24
      10'h284: dout  = 8'b00100100; //  644 :  36 - 0x24
      10'h285: dout  = 8'b00100100; //  645 :  36 - 0x24
      10'h286: dout  = 8'b00100100; //  646 :  36 - 0x24
      10'h287: dout  = 8'b00100100; //  647 :  36 - 0x24
      10'h288: dout  = 8'b00100100; //  648 :  36 - 0x24
      10'h289: dout  = 8'b00100100; //  649 :  36 - 0x24
      10'h28A: dout  = 8'b00100100; //  650 :  36 - 0x24
      10'h28B: dout  = 8'b00000010; //  651 :   2 - 0x2
      10'h28C: dout  = 8'b00100100; //  652 :  36 - 0x24
      10'h28D: dout  = 8'b00011001; //  653 :  25 - 0x19
      10'h28E: dout  = 8'b00010101; //  654 :  21 - 0x15
      10'h28F: dout  = 8'b00001010; //  655 :  10 - 0xa
      10'h290: dout  = 8'b00100010; //  656 :  34 - 0x22
      10'h291: dout  = 8'b00001110; //  657 :  14 - 0xe
      10'h292: dout  = 8'b00011011; //  658 :  27 - 0x1b
      10'h293: dout  = 8'b00100100; //  659 :  36 - 0x24
      10'h294: dout  = 8'b00010000; //  660 :  16 - 0x10
      10'h295: dout  = 8'b00001010; //  661 :  10 - 0xa
      10'h296: dout  = 8'b00010110; //  662 :  22 - 0x16
      10'h297: dout  = 8'b00001110; //  663 :  14 - 0xe
      10'h298: dout  = 8'b00100100; //  664 :  36 - 0x24
      10'h299: dout  = 8'b00100100; //  665 :  36 - 0x24
      10'h29A: dout  = 8'b00100100; //  666 :  36 - 0x24
      10'h29B: dout  = 8'b00100100; //  667 :  36 - 0x24
      10'h29C: dout  = 8'b00100100; //  668 :  36 - 0x24
      10'h29D: dout  = 8'b00100100; //  669 :  36 - 0x24
      10'h29E: dout  = 8'b00100100; //  670 :  36 - 0x24
      10'h29F: dout  = 8'b00100100; //  671 :  36 - 0x24
      10'h2A0: dout  = 8'b00100100; //  672 :  36 - 0x24 -- line 0x15
      10'h2A1: dout  = 8'b00100100; //  673 :  36 - 0x24
      10'h2A2: dout  = 8'b00100100; //  674 :  36 - 0x24
      10'h2A3: dout  = 8'b00100100; //  675 :  36 - 0x24
      10'h2A4: dout  = 8'b00110001; //  676 :  49 - 0x31
      10'h2A5: dout  = 8'b00110010; //  677 :  50 - 0x32
      10'h2A6: dout  = 8'b00100100; //  678 :  36 - 0x24
      10'h2A7: dout  = 8'b00100100; //  679 :  36 - 0x24
      10'h2A8: dout  = 8'b00100100; //  680 :  36 - 0x24
      10'h2A9: dout  = 8'b00100100; //  681 :  36 - 0x24
      10'h2AA: dout  = 8'b00100100; //  682 :  36 - 0x24
      10'h2AB: dout  = 8'b00100100; //  683 :  36 - 0x24
      10'h2AC: dout  = 8'b00100100; //  684 :  36 - 0x24
      10'h2AD: dout  = 8'b00100100; //  685 :  36 - 0x24
      10'h2AE: dout  = 8'b00100100; //  686 :  36 - 0x24
      10'h2AF: dout  = 8'b00100100; //  687 :  36 - 0x24
      10'h2B0: dout  = 8'b00100100; //  688 :  36 - 0x24
      10'h2B1: dout  = 8'b00100100; //  689 :  36 - 0x24
      10'h2B2: dout  = 8'b00100100; //  690 :  36 - 0x24
      10'h2B3: dout  = 8'b00100100; //  691 :  36 - 0x24
      10'h2B4: dout  = 8'b00100100; //  692 :  36 - 0x24
      10'h2B5: dout  = 8'b00100100; //  693 :  36 - 0x24
      10'h2B6: dout  = 8'b00100100; //  694 :  36 - 0x24
      10'h2B7: dout  = 8'b00100100; //  695 :  36 - 0x24
      10'h2B8: dout  = 8'b00100100; //  696 :  36 - 0x24
      10'h2B9: dout  = 8'b00100100; //  697 :  36 - 0x24
      10'h2BA: dout  = 8'b00100100; //  698 :  36 - 0x24
      10'h2BB: dout  = 8'b00100100; //  699 :  36 - 0x24
      10'h2BC: dout  = 8'b00100100; //  700 :  36 - 0x24
      10'h2BD: dout  = 8'b00100100; //  701 :  36 - 0x24
      10'h2BE: dout  = 8'b00100100; //  702 :  36 - 0x24
      10'h2BF: dout  = 8'b00100100; //  703 :  36 - 0x24
      10'h2C0: dout  = 8'b00100100; //  704 :  36 - 0x24 -- line 0x16
      10'h2C1: dout  = 8'b00100100; //  705 :  36 - 0x24
      10'h2C2: dout  = 8'b00100100; //  706 :  36 - 0x24
      10'h2C3: dout  = 8'b00110000; //  707 :  48 - 0x30
      10'h2C4: dout  = 8'b00100110; //  708 :  38 - 0x26
      10'h2C5: dout  = 8'b00110100; //  709 :  52 - 0x34
      10'h2C6: dout  = 8'b00110011; //  710 :  51 - 0x33
      10'h2C7: dout  = 8'b00100100; //  711 :  36 - 0x24
      10'h2C8: dout  = 8'b00100100; //  712 :  36 - 0x24
      10'h2C9: dout  = 8'b00100100; //  713 :  36 - 0x24
      10'h2CA: dout  = 8'b00100100; //  714 :  36 - 0x24
      10'h2CB: dout  = 8'b00100100; //  715 :  36 - 0x24
      10'h2CC: dout  = 8'b00100100; //  716 :  36 - 0x24
      10'h2CD: dout  = 8'b00100100; //  717 :  36 - 0x24
      10'h2CE: dout  = 8'b00100100; //  718 :  36 - 0x24
      10'h2CF: dout  = 8'b00100100; //  719 :  36 - 0x24
      10'h2D0: dout  = 8'b00100100; //  720 :  36 - 0x24
      10'h2D1: dout  = 8'b00100100; //  721 :  36 - 0x24
      10'h2D2: dout  = 8'b00100100; //  722 :  36 - 0x24
      10'h2D3: dout  = 8'b00100100; //  723 :  36 - 0x24
      10'h2D4: dout  = 8'b00100100; //  724 :  36 - 0x24
      10'h2D5: dout  = 8'b00100100; //  725 :  36 - 0x24
      10'h2D6: dout  = 8'b00100100; //  726 :  36 - 0x24
      10'h2D7: dout  = 8'b00100100; //  727 :  36 - 0x24
      10'h2D8: dout  = 8'b00100100; //  728 :  36 - 0x24
      10'h2D9: dout  = 8'b00100100; //  729 :  36 - 0x24
      10'h2DA: dout  = 8'b00100100; //  730 :  36 - 0x24
      10'h2DB: dout  = 8'b00100100; //  731 :  36 - 0x24
      10'h2DC: dout  = 8'b00100100; //  732 :  36 - 0x24
      10'h2DD: dout  = 8'b00100100; //  733 :  36 - 0x24
      10'h2DE: dout  = 8'b00100100; //  734 :  36 - 0x24
      10'h2DF: dout  = 8'b00100100; //  735 :  36 - 0x24
      10'h2E0: dout  = 8'b00100100; //  736 :  36 - 0x24 -- line 0x17
      10'h2E1: dout  = 8'b00100100; //  737 :  36 - 0x24
      10'h2E2: dout  = 8'b00110000; //  738 :  48 - 0x30
      10'h2E3: dout  = 8'b00100110; //  739 :  38 - 0x26
      10'h2E4: dout  = 8'b00100110; //  740 :  38 - 0x26
      10'h2E5: dout  = 8'b00100110; //  741 :  38 - 0x26
      10'h2E6: dout  = 8'b00100110; //  742 :  38 - 0x26
      10'h2E7: dout  = 8'b00110011; //  743 :  51 - 0x33
      10'h2E8: dout  = 8'b00100100; //  744 :  36 - 0x24
      10'h2E9: dout  = 8'b00100100; //  745 :  36 - 0x24
      10'h2EA: dout  = 8'b00100100; //  746 :  36 - 0x24
      10'h2EB: dout  = 8'b00100100; //  747 :  36 - 0x24
      10'h2EC: dout  = 8'b00011101; //  748 :  29 - 0x1d
      10'h2ED: dout  = 8'b00011000; //  749 :  24 - 0x18
      10'h2EE: dout  = 8'b00011001; //  750 :  25 - 0x19
      10'h2EF: dout  = 8'b00101000; //  751 :  40 - 0x28
      10'h2F0: dout  = 8'b00100100; //  752 :  36 - 0x24
      10'h2F1: dout  = 8'b00000000; //  753 :   0 - 0x0
      10'h2F2: dout  = 8'b00000000; //  754 :   0 - 0x0
      10'h2F3: dout  = 8'b00000000; //  755 :   0 - 0x0
      10'h2F4: dout  = 8'b00000000; //  756 :   0 - 0x0
      10'h2F5: dout  = 8'b00000000; //  757 :   0 - 0x0
      10'h2F6: dout  = 8'b00000000; //  758 :   0 - 0x0
      10'h2F7: dout  = 8'b00100100; //  759 :  36 - 0x24
      10'h2F8: dout  = 8'b00100100; //  760 :  36 - 0x24
      10'h2F9: dout  = 8'b00100100; //  761 :  36 - 0x24
      10'h2FA: dout  = 8'b00100100; //  762 :  36 - 0x24
      10'h2FB: dout  = 8'b00100100; //  763 :  36 - 0x24
      10'h2FC: dout  = 8'b00100100; //  764 :  36 - 0x24
      10'h2FD: dout  = 8'b00100100; //  765 :  36 - 0x24
      10'h2FE: dout  = 8'b00100100; //  766 :  36 - 0x24
      10'h2FF: dout  = 8'b00100100; //  767 :  36 - 0x24
      10'h300: dout  = 8'b00100100; //  768 :  36 - 0x24 -- line 0x18
      10'h301: dout  = 8'b00110000; //  769 :  48 - 0x30
      10'h302: dout  = 8'b00100110; //  770 :  38 - 0x26
      10'h303: dout  = 8'b00110100; //  771 :  52 - 0x34
      10'h304: dout  = 8'b00100110; //  772 :  38 - 0x26
      10'h305: dout  = 8'b00100110; //  773 :  38 - 0x26
      10'h306: dout  = 8'b00110100; //  774 :  52 - 0x34
      10'h307: dout  = 8'b00100110; //  775 :  38 - 0x26
      10'h308: dout  = 8'b00110011; //  776 :  51 - 0x33
      10'h309: dout  = 8'b00100100; //  777 :  36 - 0x24
      10'h30A: dout  = 8'b00100100; //  778 :  36 - 0x24
      10'h30B: dout  = 8'b00100100; //  779 :  36 - 0x24
      10'h30C: dout  = 8'b00100100; //  780 :  36 - 0x24
      10'h30D: dout  = 8'b00100100; //  781 :  36 - 0x24
      10'h30E: dout  = 8'b00100100; //  782 :  36 - 0x24
      10'h30F: dout  = 8'b00100100; //  783 :  36 - 0x24
      10'h310: dout  = 8'b00100100; //  784 :  36 - 0x24
      10'h311: dout  = 8'b00100100; //  785 :  36 - 0x24
      10'h312: dout  = 8'b00100100; //  786 :  36 - 0x24
      10'h313: dout  = 8'b00100100; //  787 :  36 - 0x24
      10'h314: dout  = 8'b00100100; //  788 :  36 - 0x24
      10'h315: dout  = 8'b00100100; //  789 :  36 - 0x24
      10'h316: dout  = 8'b00100100; //  790 :  36 - 0x24
      10'h317: dout  = 8'b00100100; //  791 :  36 - 0x24
      10'h318: dout  = 8'b00110110; //  792 :  54 - 0x36
      10'h319: dout  = 8'b00110111; //  793 :  55 - 0x37
      10'h31A: dout  = 8'b00110110; //  794 :  54 - 0x36
      10'h31B: dout  = 8'b00110111; //  795 :  55 - 0x37
      10'h31C: dout  = 8'b00110110; //  796 :  54 - 0x36
      10'h31D: dout  = 8'b00110111; //  797 :  55 - 0x37
      10'h31E: dout  = 8'b00100100; //  798 :  36 - 0x24
      10'h31F: dout  = 8'b00100100; //  799 :  36 - 0x24
      10'h320: dout  = 8'b00110000; //  800 :  48 - 0x30 -- line 0x19
      10'h321: dout  = 8'b00100110; //  801 :  38 - 0x26
      10'h322: dout  = 8'b00100110; //  802 :  38 - 0x26
      10'h323: dout  = 8'b00100110; //  803 :  38 - 0x26
      10'h324: dout  = 8'b00100110; //  804 :  38 - 0x26
      10'h325: dout  = 8'b00100110; //  805 :  38 - 0x26
      10'h326: dout  = 8'b00100110; //  806 :  38 - 0x26
      10'h327: dout  = 8'b00100110; //  807 :  38 - 0x26
      10'h328: dout  = 8'b00100110; //  808 :  38 - 0x26
      10'h329: dout  = 8'b00110011; //  809 :  51 - 0x33
      10'h32A: dout  = 8'b00100100; //  810 :  36 - 0x24
      10'h32B: dout  = 8'b00100100; //  811 :  36 - 0x24
      10'h32C: dout  = 8'b00100100; //  812 :  36 - 0x24
      10'h32D: dout  = 8'b00100100; //  813 :  36 - 0x24
      10'h32E: dout  = 8'b00100100; //  814 :  36 - 0x24
      10'h32F: dout  = 8'b00100100; //  815 :  36 - 0x24
      10'h330: dout  = 8'b00100100; //  816 :  36 - 0x24
      10'h331: dout  = 8'b00100100; //  817 :  36 - 0x24
      10'h332: dout  = 8'b00100100; //  818 :  36 - 0x24
      10'h333: dout  = 8'b00100100; //  819 :  36 - 0x24
      10'h334: dout  = 8'b00100100; //  820 :  36 - 0x24
      10'h335: dout  = 8'b00100100; //  821 :  36 - 0x24
      10'h336: dout  = 8'b00100100; //  822 :  36 - 0x24
      10'h337: dout  = 8'b00110101; //  823 :  53 - 0x35
      10'h338: dout  = 8'b00100101; //  824 :  37 - 0x25
      10'h339: dout  = 8'b00100101; //  825 :  37 - 0x25
      10'h33A: dout  = 8'b00100101; //  826 :  37 - 0x25
      10'h33B: dout  = 8'b00100101; //  827 :  37 - 0x25
      10'h33C: dout  = 8'b00100101; //  828 :  37 - 0x25
      10'h33D: dout  = 8'b00100101; //  829 :  37 - 0x25
      10'h33E: dout  = 8'b00111000; //  830 :  56 - 0x38
      10'h33F: dout  = 8'b00100100; //  831 :  36 - 0x24
      10'h340: dout  = 8'b10110100; //  832 : 180 - 0xb4 -- line 0x1a
      10'h341: dout  = 8'b10110101; //  833 : 181 - 0xb5
      10'h342: dout  = 8'b10110100; //  834 : 180 - 0xb4
      10'h343: dout  = 8'b10110101; //  835 : 181 - 0xb5
      10'h344: dout  = 8'b10110100; //  836 : 180 - 0xb4
      10'h345: dout  = 8'b10110101; //  837 : 181 - 0xb5
      10'h346: dout  = 8'b10110100; //  838 : 180 - 0xb4
      10'h347: dout  = 8'b10110101; //  839 : 181 - 0xb5
      10'h348: dout  = 8'b10110100; //  840 : 180 - 0xb4
      10'h349: dout  = 8'b10110101; //  841 : 181 - 0xb5
      10'h34A: dout  = 8'b10110100; //  842 : 180 - 0xb4
      10'h34B: dout  = 8'b10110101; //  843 : 181 - 0xb5
      10'h34C: dout  = 8'b10110100; //  844 : 180 - 0xb4
      10'h34D: dout  = 8'b10110101; //  845 : 181 - 0xb5
      10'h34E: dout  = 8'b10110100; //  846 : 180 - 0xb4
      10'h34F: dout  = 8'b10110101; //  847 : 181 - 0xb5
      10'h350: dout  = 8'b10110100; //  848 : 180 - 0xb4
      10'h351: dout  = 8'b10110101; //  849 : 181 - 0xb5
      10'h352: dout  = 8'b10110100; //  850 : 180 - 0xb4
      10'h353: dout  = 8'b10110101; //  851 : 181 - 0xb5
      10'h354: dout  = 8'b10110100; //  852 : 180 - 0xb4
      10'h355: dout  = 8'b10110101; //  853 : 181 - 0xb5
      10'h356: dout  = 8'b10110100; //  854 : 180 - 0xb4
      10'h357: dout  = 8'b10110101; //  855 : 181 - 0xb5
      10'h358: dout  = 8'b10110100; //  856 : 180 - 0xb4
      10'h359: dout  = 8'b10110101; //  857 : 181 - 0xb5
      10'h35A: dout  = 8'b10110100; //  858 : 180 - 0xb4
      10'h35B: dout  = 8'b10110101; //  859 : 181 - 0xb5
      10'h35C: dout  = 8'b10110100; //  860 : 180 - 0xb4
      10'h35D: dout  = 8'b10110101; //  861 : 181 - 0xb5
      10'h35E: dout  = 8'b10110100; //  862 : 180 - 0xb4
      10'h35F: dout  = 8'b10110101; //  863 : 181 - 0xb5
      10'h360: dout  = 8'b10110110; //  864 : 182 - 0xb6 -- line 0x1b
      10'h361: dout  = 8'b10110111; //  865 : 183 - 0xb7
      10'h362: dout  = 8'b10110110; //  866 : 182 - 0xb6
      10'h363: dout  = 8'b10110111; //  867 : 183 - 0xb7
      10'h364: dout  = 8'b10110110; //  868 : 182 - 0xb6
      10'h365: dout  = 8'b10110111; //  869 : 183 - 0xb7
      10'h366: dout  = 8'b10110110; //  870 : 182 - 0xb6
      10'h367: dout  = 8'b10110111; //  871 : 183 - 0xb7
      10'h368: dout  = 8'b10110110; //  872 : 182 - 0xb6
      10'h369: dout  = 8'b10110111; //  873 : 183 - 0xb7
      10'h36A: dout  = 8'b10110110; //  874 : 182 - 0xb6
      10'h36B: dout  = 8'b10110111; //  875 : 183 - 0xb7
      10'h36C: dout  = 8'b10110110; //  876 : 182 - 0xb6
      10'h36D: dout  = 8'b10110111; //  877 : 183 - 0xb7
      10'h36E: dout  = 8'b10110110; //  878 : 182 - 0xb6
      10'h36F: dout  = 8'b10110111; //  879 : 183 - 0xb7
      10'h370: dout  = 8'b10110110; //  880 : 182 - 0xb6
      10'h371: dout  = 8'b10110111; //  881 : 183 - 0xb7
      10'h372: dout  = 8'b10110110; //  882 : 182 - 0xb6
      10'h373: dout  = 8'b10110111; //  883 : 183 - 0xb7
      10'h374: dout  = 8'b10110110; //  884 : 182 - 0xb6
      10'h375: dout  = 8'b10110111; //  885 : 183 - 0xb7
      10'h376: dout  = 8'b10110110; //  886 : 182 - 0xb6
      10'h377: dout  = 8'b10110111; //  887 : 183 - 0xb7
      10'h378: dout  = 8'b10110110; //  888 : 182 - 0xb6
      10'h379: dout  = 8'b10110111; //  889 : 183 - 0xb7
      10'h37A: dout  = 8'b10110110; //  890 : 182 - 0xb6
      10'h37B: dout  = 8'b10110111; //  891 : 183 - 0xb7
      10'h37C: dout  = 8'b10110110; //  892 : 182 - 0xb6
      10'h37D: dout  = 8'b10110111; //  893 : 183 - 0xb7
      10'h37E: dout  = 8'b10110110; //  894 : 182 - 0xb6
      10'h37F: dout  = 8'b10110111; //  895 : 183 - 0xb7
      10'h380: dout  = 8'b10110100; //  896 : 180 - 0xb4 -- line 0x1c
      10'h381: dout  = 8'b10110101; //  897 : 181 - 0xb5
      10'h382: dout  = 8'b10110100; //  898 : 180 - 0xb4
      10'h383: dout  = 8'b10110101; //  899 : 181 - 0xb5
      10'h384: dout  = 8'b10110100; //  900 : 180 - 0xb4
      10'h385: dout  = 8'b10110101; //  901 : 181 - 0xb5
      10'h386: dout  = 8'b10110100; //  902 : 180 - 0xb4
      10'h387: dout  = 8'b10110101; //  903 : 181 - 0xb5
      10'h388: dout  = 8'b10110100; //  904 : 180 - 0xb4
      10'h389: dout  = 8'b10110101; //  905 : 181 - 0xb5
      10'h38A: dout  = 8'b10110100; //  906 : 180 - 0xb4
      10'h38B: dout  = 8'b10110101; //  907 : 181 - 0xb5
      10'h38C: dout  = 8'b10110100; //  908 : 180 - 0xb4
      10'h38D: dout  = 8'b10110101; //  909 : 181 - 0xb5
      10'h38E: dout  = 8'b10110100; //  910 : 180 - 0xb4
      10'h38F: dout  = 8'b10110101; //  911 : 181 - 0xb5
      10'h390: dout  = 8'b10110100; //  912 : 180 - 0xb4
      10'h391: dout  = 8'b10110101; //  913 : 181 - 0xb5
      10'h392: dout  = 8'b10110100; //  914 : 180 - 0xb4
      10'h393: dout  = 8'b10110101; //  915 : 181 - 0xb5
      10'h394: dout  = 8'b10110100; //  916 : 180 - 0xb4
      10'h395: dout  = 8'b10110101; //  917 : 181 - 0xb5
      10'h396: dout  = 8'b10110100; //  918 : 180 - 0xb4
      10'h397: dout  = 8'b10110101; //  919 : 181 - 0xb5
      10'h398: dout  = 8'b10110100; //  920 : 180 - 0xb4
      10'h399: dout  = 8'b10110101; //  921 : 181 - 0xb5
      10'h39A: dout  = 8'b10110100; //  922 : 180 - 0xb4
      10'h39B: dout  = 8'b10110101; //  923 : 181 - 0xb5
      10'h39C: dout  = 8'b10110100; //  924 : 180 - 0xb4
      10'h39D: dout  = 8'b10110101; //  925 : 181 - 0xb5
      10'h39E: dout  = 8'b10110100; //  926 : 180 - 0xb4
      10'h39F: dout  = 8'b10110101; //  927 : 181 - 0xb5
      10'h3A0: dout  = 8'b10110110; //  928 : 182 - 0xb6 -- line 0x1d
      10'h3A1: dout  = 8'b10110111; //  929 : 183 - 0xb7
      10'h3A2: dout  = 8'b10110110; //  930 : 182 - 0xb6
      10'h3A3: dout  = 8'b10110111; //  931 : 183 - 0xb7
      10'h3A4: dout  = 8'b10110110; //  932 : 182 - 0xb6
      10'h3A5: dout  = 8'b10110111; //  933 : 183 - 0xb7
      10'h3A6: dout  = 8'b10110110; //  934 : 182 - 0xb6
      10'h3A7: dout  = 8'b10110111; //  935 : 183 - 0xb7
      10'h3A8: dout  = 8'b10110110; //  936 : 182 - 0xb6
      10'h3A9: dout  = 8'b10110111; //  937 : 183 - 0xb7
      10'h3AA: dout  = 8'b10110110; //  938 : 182 - 0xb6
      10'h3AB: dout  = 8'b10110111; //  939 : 183 - 0xb7
      10'h3AC: dout  = 8'b10110110; //  940 : 182 - 0xb6
      10'h3AD: dout  = 8'b10110111; //  941 : 183 - 0xb7
      10'h3AE: dout  = 8'b10110110; //  942 : 182 - 0xb6
      10'h3AF: dout  = 8'b10110111; //  943 : 183 - 0xb7
      10'h3B0: dout  = 8'b10110110; //  944 : 182 - 0xb6
      10'h3B1: dout  = 8'b10110111; //  945 : 183 - 0xb7
      10'h3B2: dout  = 8'b10110110; //  946 : 182 - 0xb6
      10'h3B3: dout  = 8'b10110111; //  947 : 183 - 0xb7
      10'h3B4: dout  = 8'b10110110; //  948 : 182 - 0xb6
      10'h3B5: dout  = 8'b10110111; //  949 : 183 - 0xb7
      10'h3B6: dout  = 8'b10110110; //  950 : 182 - 0xb6
      10'h3B7: dout  = 8'b10110111; //  951 : 183 - 0xb7
      10'h3B8: dout  = 8'b10110110; //  952 : 182 - 0xb6
      10'h3B9: dout  = 8'b10110111; //  953 : 183 - 0xb7
      10'h3BA: dout  = 8'b10110110; //  954 : 182 - 0xb6
      10'h3BB: dout  = 8'b10110111; //  955 : 183 - 0xb7
      10'h3BC: dout  = 8'b10110110; //  956 : 182 - 0xb6
      10'h3BD: dout  = 8'b10110111; //  957 : 183 - 0xb7
      10'h3BE: dout  = 8'b10110110; //  958 : 182 - 0xb6
      10'h3BF: dout  = 8'b10110111; //  959 : 183 - 0xb7
        //-- Attribute Table 0----
      10'h3C0: dout  = 8'b10101010; //  960 : 170 - 0xaa
      10'h3C1: dout  = 8'b10101010; //  961 : 170 - 0xaa
      10'h3C2: dout  = 8'b11101010; //  962 : 234 - 0xea
      10'h3C3: dout  = 8'b10101010; //  963 : 170 - 0xaa
      10'h3C4: dout  = 8'b10101010; //  964 : 170 - 0xaa
      10'h3C5: dout  = 8'b10101010; //  965 : 170 - 0xaa
      10'h3C6: dout  = 8'b10101010; //  966 : 170 - 0xaa
      10'h3C7: dout  = 8'b10101010; //  967 : 170 - 0xaa
      10'h3C8: dout  = 8'b00000000; //  968 :   0 - 0x0
      10'h3C9: dout  = 8'b01010101; //  969 :  85 - 0x55
      10'h3CA: dout  = 8'b01010101; //  970 :  85 - 0x55
      10'h3CB: dout  = 8'b01010101; //  971 :  85 - 0x55
      10'h3CC: dout  = 8'b01010101; //  972 :  85 - 0x55
      10'h3CD: dout  = 8'b01010101; //  973 :  85 - 0x55
      10'h3CE: dout  = 8'b01010101; //  974 :  85 - 0x55
      10'h3CF: dout  = 8'b01010101; //  975 :  85 - 0x55
      10'h3D0: dout  = 8'b01010101; //  976 :  85 - 0x55
      10'h3D1: dout  = 8'b01010101; //  977 :  85 - 0x55
      10'h3D2: dout  = 8'b01010101; //  978 :  85 - 0x55
      10'h3D3: dout  = 8'b01010101; //  979 :  85 - 0x55
      10'h3D4: dout  = 8'b01010101; //  980 :  85 - 0x55
      10'h3D5: dout  = 8'b01010101; //  981 :  85 - 0x55
      10'h3D6: dout  = 8'b01010101; //  982 :  85 - 0x55
      10'h3D7: dout  = 8'b01010101; //  983 :  85 - 0x55
      10'h3D8: dout  = 8'b01010101; //  984 :  85 - 0x55
      10'h3D9: dout  = 8'b01010101; //  985 :  85 - 0x55
      10'h3DA: dout  = 8'b01010101; //  986 :  85 - 0x55
      10'h3DB: dout  = 8'b01010101; //  987 :  85 - 0x55
      10'h3DC: dout  = 8'b01010101; //  988 :  85 - 0x55
      10'h3DD: dout  = 8'b01010101; //  989 :  85 - 0x55
      10'h3DE: dout  = 8'b01010101; //  990 :  85 - 0x55
      10'h3DF: dout  = 8'b00000000; //  991 :   0 - 0x0
      10'h3E0: dout  = 8'b00000000; //  992 :   0 - 0x0
      10'h3E1: dout  = 8'b00000000; //  993 :   0 - 0x0
      10'h3E2: dout  = 8'b10011001; //  994 : 153 - 0x99
      10'h3E3: dout  = 8'b10101010; //  995 : 170 - 0xaa
      10'h3E4: dout  = 8'b10101010; //  996 : 170 - 0xaa
      10'h3E5: dout  = 8'b10101010; //  997 : 170 - 0xaa
      10'h3E6: dout  = 8'b00000000; //  998 :   0 - 0x0
      10'h3E7: dout  = 8'b00000000; //  999 :   0 - 0x0
      10'h3E8: dout  = 8'b00000000; // 1000 :   0 - 0x0
      10'h3E9: dout  = 8'b00000000; // 1001 :   0 - 0x0
      10'h3EA: dout  = 8'b10011001; // 1002 : 153 - 0x99
      10'h3EB: dout  = 8'b10101010; // 1003 : 170 - 0xaa
      10'h3EC: dout  = 8'b10101010; // 1004 : 170 - 0xaa
      10'h3ED: dout  = 8'b10101010; // 1005 : 170 - 0xaa
      10'h3EE: dout  = 8'b00000000; // 1006 :   0 - 0x0
      10'h3EF: dout  = 8'b00000000; // 1007 :   0 - 0x0
      10'h3F0: dout  = 8'b01010000; // 1008 :  80 - 0x50
      10'h3F1: dout  = 8'b01010000; // 1009 :  80 - 0x50
      10'h3F2: dout  = 8'b01010000; // 1010 :  80 - 0x50
      10'h3F3: dout  = 8'b01010000; // 1011 :  80 - 0x50
      10'h3F4: dout  = 8'b01010000; // 1012 :  80 - 0x50
      10'h3F5: dout  = 8'b01010000; // 1013 :  80 - 0x50
      10'h3F6: dout  = 8'b01010000; // 1014 :  80 - 0x50
      10'h3F7: dout  = 8'b01010000; // 1015 :  80 - 0x50
      10'h3F8: dout  = 8'b00000101; // 1016 :   5 - 0x5
      10'h3F9: dout  = 8'b00000101; // 1017 :   5 - 0x5
      10'h3FA: dout  = 8'b00000101; // 1018 :   5 - 0x5
      10'h3FB: dout  = 8'b00000101; // 1019 :   5 - 0x5
      10'h3FC: dout  = 8'b00000101; // 1020 :   5 - 0x5
      10'h3FD: dout  = 8'b00000101; // 1021 :   5 - 0x5
      10'h3FE: dout  = 8'b00000101; // 1022 :   5 - 0x5
      10'h3FF: dout  = 8'b00000101; // 1023 :   5 - 0x5
    endcase
  end

endmodule
