--- Autcmatically generated VHDL ROM from a NES memory file----
---   SPRITEs MEMORY (OAM)
-- https://wiki.nesdev.com/w/index.php/PPU_OAM


---  Original memory dump file name: pacman_oam_00.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_OAM_PACMAN_00 is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(8-1 downto 0);  --256 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_OAM_PACMAN_00;

architecture BEHAVIORAL of ROM_OAM_PACMAN_00 is
  signal addr_int  : natural range 0 to 2**8-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
    "10101011", --    0 -  0x0  :  171 - 0xab -- Sprite 0x0
    "00000010", --    1 -  0x1  :    2 - 0x2
    "00000000", --    2 -  0x2  :    0 - 0x0
    "01001111", --    3 -  0x3  :   79 - 0x4f
    "10101011", --    4 -  0x4  :  171 - 0xab -- Sprite 0x1
    "00000001", --    5 -  0x5  :    1 - 0x1
    "00000000", --    6 -  0x6  :    0 - 0x0
    "01010111", --    7 -  0x7  :   87 - 0x57
    "10110011", --    8 -  0x8  :  179 - 0xb3 -- Sprite 0x2
    "00000010", --    9 -  0x9  :    2 - 0x2
    "10000000", --   10 -  0xa  :  128 - 0x80
    "01001111", --   11 -  0xb  :   79 - 0x4f
    "10110011", --   12 -  0xc  :  179 - 0xb3 -- Sprite 0x3
    "00000001", --   13 -  0xd  :    1 - 0x1
    "10000000", --   14 -  0xe  :  128 - 0x80
    "01010111", --   15 -  0xf  :   87 - 0x57
    "01011011", --   16 - 0x10  :   91 - 0x5b -- Sprite 0x4
    "00011011", --   17 - 0x11  :   27 - 0x1b
    "00000000", --   18 - 0x12  :    0 - 0x0
    "01010000", --   19 - 0x13  :   80 - 0x50
    "01011011", --   20 - 0x14  :   91 - 0x5b -- Sprite 0x5
    "00011100", --   21 - 0x15  :   28 - 0x1c
    "00000000", --   22 - 0x16  :    0 - 0x0
    "01011000", --   23 - 0x17  :   88 - 0x58
    "01100011", --   24 - 0x18  :   99 - 0x63 -- Sprite 0x6
    "00011101", --   25 - 0x19  :   29 - 0x1d
    "00000000", --   26 - 0x1a  :    0 - 0x0
    "01010000", --   27 - 0x1b  :   80 - 0x50
    "01100011", --   28 - 0x1c  :   99 - 0x63 -- Sprite 0x7
    "00011111", --   29 - 0x1d  :   31 - 0x1f
    "00000000", --   30 - 0x1e  :    0 - 0x0
    "01011000", --   31 - 0x1f  :   88 - 0x58
    "01101111", --   32 - 0x20  :  111 - 0x6f -- Sprite 0x8
    "00011000", --   33 - 0x21  :   24 - 0x18
    "00000001", --   34 - 0x22  :    1 - 0x1
    "01010100", --   35 - 0x23  :   84 - 0x54
    "01101111", --   36 - 0x24  :  111 - 0x6f -- Sprite 0x9
    "00011000", --   37 - 0x25  :   24 - 0x18
    "01000001", --   38 - 0x26  :   65 - 0x41
    "01011100", --   39 - 0x27  :   92 - 0x5c
    "01110111", --   40 - 0x28  :  119 - 0x77 -- Sprite 0xa
    "00011001", --   41 - 0x29  :   25 - 0x19
    "00000001", --   42 - 0x2a  :    1 - 0x1
    "01010100", --   43 - 0x2b  :   84 - 0x54
    "01110111", --   44 - 0x2c  :  119 - 0x77 -- Sprite 0xb
    "00011001", --   45 - 0x2d  :   25 - 0x19
    "01000001", --   46 - 0x2e  :   65 - 0x41
    "01011100", --   47 - 0x2f  :   92 - 0x5c
    "01101111", --   48 - 0x30  :  111 - 0x6f -- Sprite 0xc
    "00011000", --   49 - 0x31  :   24 - 0x18
    "00000010", --   50 - 0x32  :    2 - 0x2
    "01001100", --   51 - 0x33  :   76 - 0x4c
    "01101111", --   52 - 0x34  :  111 - 0x6f -- Sprite 0xd
    "00011000", --   53 - 0x35  :   24 - 0x18
    "01000010", --   54 - 0x36  :   66 - 0x42
    "01010100", --   55 - 0x37  :   84 - 0x54
    "01110111", --   56 - 0x38  :  119 - 0x77 -- Sprite 0xe
    "00011001", --   57 - 0x39  :   25 - 0x19
    "00000010", --   58 - 0x3a  :    2 - 0x2
    "01001100", --   59 - 0x3b  :   76 - 0x4c
    "01110111", --   60 - 0x3c  :  119 - 0x77 -- Sprite 0xf
    "00011001", --   61 - 0x3d  :   25 - 0x19
    "01000010", --   62 - 0x3e  :   66 - 0x42
    "01010100", --   63 - 0x3f  :   84 - 0x54
    "01101111", --   64 - 0x40  :  111 - 0x6f -- Sprite 0x10
    "00011000", --   65 - 0x41  :   24 - 0x18
    "00000011", --   66 - 0x42  :    3 - 0x3
    "01011100", --   67 - 0x43  :   92 - 0x5c
    "01101111", --   68 - 0x44  :  111 - 0x6f -- Sprite 0x11
    "00011000", --   69 - 0x45  :   24 - 0x18
    "01000011", --   70 - 0x46  :   67 - 0x43
    "01100100", --   71 - 0x47  :  100 - 0x64
    "01110111", --   72 - 0x48  :  119 - 0x77 -- Sprite 0x12
    "00011001", --   73 - 0x49  :   25 - 0x19
    "00000011", --   74 - 0x4a  :    3 - 0x3
    "01011100", --   75 - 0x4b  :   92 - 0x5c
    "01110111", --   76 - 0x4c  :  119 - 0x77 -- Sprite 0x13
    "00011001", --   77 - 0x4d  :   25 - 0x19
    "01000011", --   78 - 0x4e  :   67 - 0x43
    "01100100", --   79 - 0x4f  :  100 - 0x64
    "11111111", --   80 - 0x50  :  255 - 0xff -- Sprite 0x14
    "01001100", --   81 - 0x51  :   76 - 0x4c
    "00000000", --   82 - 0x52  :    0 - 0x0
    "11111111", --   83 - 0x53  :  255 - 0xff
    "11111111", --   84 - 0x54  :  255 - 0xff -- Sprite 0x15
    "01001100", --   85 - 0x55  :   76 - 0x4c
    "00000000", --   86 - 0x56  :    0 - 0x0
    "11111111", --   87 - 0x57  :  255 - 0xff
    "11111111", --   88 - 0x58  :  255 - 0xff -- Sprite 0x16
    "01001100", --   89 - 0x59  :   76 - 0x4c
    "00000000", --   90 - 0x5a  :    0 - 0x0
    "11111111", --   91 - 0x5b  :  255 - 0xff
    "11111111", --   92 - 0x5c  :  255 - 0xff -- Sprite 0x17
    "01001100", --   93 - 0x5d  :   76 - 0x4c
    "00000000", --   94 - 0x5e  :    0 - 0x0
    "11111111", --   95 - 0x5f  :  255 - 0xff
    "00000000", --   96 - 0x60  :    0 - 0x0 -- Sprite 0x18
    "00000000", --   97 - 0x61  :    0 - 0x0
    "00000000", --   98 - 0x62  :    0 - 0x0
    "00000000", --   99 - 0x63  :    0 - 0x0
    "00000000", --  100 - 0x64  :    0 - 0x0 -- Sprite 0x19
    "00000000", --  101 - 0x65  :    0 - 0x0
    "00000000", --  102 - 0x66  :    0 - 0x0
    "00000000", --  103 - 0x67  :    0 - 0x0
    "00000000", --  104 - 0x68  :    0 - 0x0 -- Sprite 0x1a
    "00000000", --  105 - 0x69  :    0 - 0x0
    "00000000", --  106 - 0x6a  :    0 - 0x0
    "00000000", --  107 - 0x6b  :    0 - 0x0
    "00000000", --  108 - 0x6c  :    0 - 0x0 -- Sprite 0x1b
    "00000000", --  109 - 0x6d  :    0 - 0x0
    "00000000", --  110 - 0x6e  :    0 - 0x0
    "00000000", --  111 - 0x6f  :    0 - 0x0
    "00000000", --  112 - 0x70  :    0 - 0x0 -- Sprite 0x1c
    "00000000", --  113 - 0x71  :    0 - 0x0
    "00000000", --  114 - 0x72  :    0 - 0x0
    "00000000", --  115 - 0x73  :    0 - 0x0
    "00000000", --  116 - 0x74  :    0 - 0x0 -- Sprite 0x1d
    "00000000", --  117 - 0x75  :    0 - 0x0
    "00000000", --  118 - 0x76  :    0 - 0x0
    "00000000", --  119 - 0x77  :    0 - 0x0
    "00000000", --  120 - 0x78  :    0 - 0x0 -- Sprite 0x1e
    "00000000", --  121 - 0x79  :    0 - 0x0
    "00000000", --  122 - 0x7a  :    0 - 0x0
    "00000000", --  123 - 0x7b  :    0 - 0x0
    "00000000", --  124 - 0x7c  :    0 - 0x0 -- Sprite 0x1f
    "00000000", --  125 - 0x7d  :    0 - 0x0
    "00000000", --  126 - 0x7e  :    0 - 0x0
    "00000000", --  127 - 0x7f  :    0 - 0x0
    "00000000", --  128 - 0x80  :    0 - 0x0 -- Sprite 0x20
    "00000000", --  129 - 0x81  :    0 - 0x0
    "00000000", --  130 - 0x82  :    0 - 0x0
    "00000000", --  131 - 0x83  :    0 - 0x0
    "00000000", --  132 - 0x84  :    0 - 0x0 -- Sprite 0x21
    "00000000", --  133 - 0x85  :    0 - 0x0
    "00000000", --  134 - 0x86  :    0 - 0x0
    "00000000", --  135 - 0x87  :    0 - 0x0
    "00000000", --  136 - 0x88  :    0 - 0x0 -- Sprite 0x22
    "00000000", --  137 - 0x89  :    0 - 0x0
    "00000000", --  138 - 0x8a  :    0 - 0x0
    "00000000", --  139 - 0x8b  :    0 - 0x0
    "00000000", --  140 - 0x8c  :    0 - 0x0 -- Sprite 0x23
    "00000000", --  141 - 0x8d  :    0 - 0x0
    "00000000", --  142 - 0x8e  :    0 - 0x0
    "00000000", --  143 - 0x8f  :    0 - 0x0
    "00000000", --  144 - 0x90  :    0 - 0x0 -- Sprite 0x24
    "00000000", --  145 - 0x91  :    0 - 0x0
    "00000000", --  146 - 0x92  :    0 - 0x0
    "00000000", --  147 - 0x93  :    0 - 0x0
    "00000000", --  148 - 0x94  :    0 - 0x0 -- Sprite 0x25
    "00000000", --  149 - 0x95  :    0 - 0x0
    "00000000", --  150 - 0x96  :    0 - 0x0
    "00000000", --  151 - 0x97  :    0 - 0x0
    "00000000", --  152 - 0x98  :    0 - 0x0 -- Sprite 0x26
    "00000000", --  153 - 0x99  :    0 - 0x0
    "00000000", --  154 - 0x9a  :    0 - 0x0
    "00000000", --  155 - 0x9b  :    0 - 0x0
    "00000000", --  156 - 0x9c  :    0 - 0x0 -- Sprite 0x27
    "00000000", --  157 - 0x9d  :    0 - 0x0
    "00000000", --  158 - 0x9e  :    0 - 0x0
    "00000000", --  159 - 0x9f  :    0 - 0x0
    "00000000", --  160 - 0xa0  :    0 - 0x0 -- Sprite 0x28
    "00000000", --  161 - 0xa1  :    0 - 0x0
    "00000000", --  162 - 0xa2  :    0 - 0x0
    "00000000", --  163 - 0xa3  :    0 - 0x0
    "00000000", --  164 - 0xa4  :    0 - 0x0 -- Sprite 0x29
    "00000000", --  165 - 0xa5  :    0 - 0x0
    "00000000", --  166 - 0xa6  :    0 - 0x0
    "00000000", --  167 - 0xa7  :    0 - 0x0
    "00000000", --  168 - 0xa8  :    0 - 0x0 -- Sprite 0x2a
    "00000000", --  169 - 0xa9  :    0 - 0x0
    "00000000", --  170 - 0xaa  :    0 - 0x0
    "00000000", --  171 - 0xab  :    0 - 0x0
    "00000000", --  172 - 0xac  :    0 - 0x0 -- Sprite 0x2b
    "00000000", --  173 - 0xad  :    0 - 0x0
    "00000000", --  174 - 0xae  :    0 - 0x0
    "00000000", --  175 - 0xaf  :    0 - 0x0
    "00000000", --  176 - 0xb0  :    0 - 0x0 -- Sprite 0x2c
    "00000000", --  177 - 0xb1  :    0 - 0x0
    "00000000", --  178 - 0xb2  :    0 - 0x0
    "00000000", --  179 - 0xb3  :    0 - 0x0
    "00000000", --  180 - 0xb4  :    0 - 0x0 -- Sprite 0x2d
    "00000000", --  181 - 0xb5  :    0 - 0x0
    "00000000", --  182 - 0xb6  :    0 - 0x0
    "00000000", --  183 - 0xb7  :    0 - 0x0
    "00000000", --  184 - 0xb8  :    0 - 0x0 -- Sprite 0x2e
    "00000000", --  185 - 0xb9  :    0 - 0x0
    "00000000", --  186 - 0xba  :    0 - 0x0
    "00000000", --  187 - 0xbb  :    0 - 0x0
    "00000000", --  188 - 0xbc  :    0 - 0x0 -- Sprite 0x2f
    "00000000", --  189 - 0xbd  :    0 - 0x0
    "00000000", --  190 - 0xbe  :    0 - 0x0
    "00000000", --  191 - 0xbf  :    0 - 0x0
    "00000000", --  192 - 0xc0  :    0 - 0x0 -- Sprite 0x30
    "00000000", --  193 - 0xc1  :    0 - 0x0
    "00000000", --  194 - 0xc2  :    0 - 0x0
    "00000000", --  195 - 0xc3  :    0 - 0x0
    "00000000", --  196 - 0xc4  :    0 - 0x0 -- Sprite 0x31
    "00000000", --  197 - 0xc5  :    0 - 0x0
    "00000000", --  198 - 0xc6  :    0 - 0x0
    "00000000", --  199 - 0xc7  :    0 - 0x0
    "00000000", --  200 - 0xc8  :    0 - 0x0 -- Sprite 0x32
    "00000000", --  201 - 0xc9  :    0 - 0x0
    "00000000", --  202 - 0xca  :    0 - 0x0
    "00000000", --  203 - 0xcb  :    0 - 0x0
    "00000000", --  204 - 0xcc  :    0 - 0x0 -- Sprite 0x33
    "00000000", --  205 - 0xcd  :    0 - 0x0
    "00000000", --  206 - 0xce  :    0 - 0x0
    "00000000", --  207 - 0xcf  :    0 - 0x0
    "00000000", --  208 - 0xd0  :    0 - 0x0 -- Sprite 0x34
    "00000000", --  209 - 0xd1  :    0 - 0x0
    "00000000", --  210 - 0xd2  :    0 - 0x0
    "00000000", --  211 - 0xd3  :    0 - 0x0
    "00000000", --  212 - 0xd4  :    0 - 0x0 -- Sprite 0x35
    "00000000", --  213 - 0xd5  :    0 - 0x0
    "00000000", --  214 - 0xd6  :    0 - 0x0
    "00000000", --  215 - 0xd7  :    0 - 0x0
    "00000000", --  216 - 0xd8  :    0 - 0x0 -- Sprite 0x36
    "00000000", --  217 - 0xd9  :    0 - 0x0
    "00000000", --  218 - 0xda  :    0 - 0x0
    "00000000", --  219 - 0xdb  :    0 - 0x0
    "00000000", --  220 - 0xdc  :    0 - 0x0 -- Sprite 0x37
    "00000000", --  221 - 0xdd  :    0 - 0x0
    "00000000", --  222 - 0xde  :    0 - 0x0
    "00000000", --  223 - 0xdf  :    0 - 0x0
    "00000000", --  224 - 0xe0  :    0 - 0x0 -- Sprite 0x38
    "00000000", --  225 - 0xe1  :    0 - 0x0
    "00000000", --  226 - 0xe2  :    0 - 0x0
    "00000000", --  227 - 0xe3  :    0 - 0x0
    "00000000", --  228 - 0xe4  :    0 - 0x0 -- Sprite 0x39
    "00000000", --  229 - 0xe5  :    0 - 0x0
    "00000000", --  230 - 0xe6  :    0 - 0x0
    "00000000", --  231 - 0xe7  :    0 - 0x0
    "00000000", --  232 - 0xe8  :    0 - 0x0 -- Sprite 0x3a
    "00000000", --  233 - 0xe9  :    0 - 0x0
    "00000000", --  234 - 0xea  :    0 - 0x0
    "00000000", --  235 - 0xeb  :    0 - 0x0
    "00000000", --  236 - 0xec  :    0 - 0x0 -- Sprite 0x3b
    "00000000", --  237 - 0xed  :    0 - 0x0
    "00000000", --  238 - 0xee  :    0 - 0x0
    "00000000", --  239 - 0xef  :    0 - 0x0
    "00000000", --  240 - 0xf0  :    0 - 0x0 -- Sprite 0x3c
    "00000000", --  241 - 0xf1  :    0 - 0x0
    "00000000", --  242 - 0xf2  :    0 - 0x0
    "00000000", --  243 - 0xf3  :    0 - 0x0
    "00000000", --  244 - 0xf4  :    0 - 0x0 -- Sprite 0x3d
    "00000000", --  245 - 0xf5  :    0 - 0x0
    "00000000", --  246 - 0xf6  :    0 - 0x0
    "00000000", --  247 - 0xf7  :    0 - 0x0
    "00000000", --  248 - 0xf8  :    0 - 0x0 -- Sprite 0x3e
    "00000000", --  249 - 0xf9  :    0 - 0x0
    "00000000", --  250 - 0xfa  :    0 - 0x0
    "00000000", --  251 - 0xfb  :    0 - 0x0
    "00000000", --  252 - 0xfc  :    0 - 0x0 -- Sprite 0x3f
    "00000000", --  253 - 0xfd  :    0 - 0x0
    "00000000", --  254 - 0xfe  :    0 - 0x0
    "00000000"  --  255 - 0xff  :    0 - 0x0
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
