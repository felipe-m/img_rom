//- Autcmatically generated verilog ROM from a NES memory file----
//-   NAME TABLE
// https://wiki.nesdev.com/w/index.php/PPU_nametables
//- Only the first Name Table: 1KiB


//-  Original memory dump file name: lawnmower_ntable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_NTABLE_LAWN_00
  (
     input     clk,   // clock
     input      [10-1:0] addr,  //1024 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
     //----- Name Table 0---------
      10'h0: dout <= 8'b10101001; //    0 : 169 - 0xa9 -- line 0x0
      10'h1: dout <= 8'b10101001; //    1 : 169 - 0xa9
      10'h2: dout <= 8'b10101001; //    2 : 169 - 0xa9
      10'h3: dout <= 8'b10101001; //    3 : 169 - 0xa9
      10'h4: dout <= 8'b10101001; //    4 : 169 - 0xa9
      10'h5: dout <= 8'b10101001; //    5 : 169 - 0xa9
      10'h6: dout <= 8'b10101001; //    6 : 169 - 0xa9
      10'h7: dout <= 8'b10101001; //    7 : 169 - 0xa9
      10'h8: dout <= 8'b10101001; //    8 : 169 - 0xa9
      10'h9: dout <= 8'b10101001; //    9 : 169 - 0xa9
      10'hA: dout <= 8'b10101001; //   10 : 169 - 0xa9
      10'hB: dout <= 8'b10101001; //   11 : 169 - 0xa9
      10'hC: dout <= 8'b10101001; //   12 : 169 - 0xa9
      10'hD: dout <= 8'b10101001; //   13 : 169 - 0xa9
      10'hE: dout <= 8'b10101001; //   14 : 169 - 0xa9
      10'hF: dout <= 8'b10101001; //   15 : 169 - 0xa9
      10'h10: dout <= 8'b10101001; //   16 : 169 - 0xa9
      10'h11: dout <= 8'b10101001; //   17 : 169 - 0xa9
      10'h12: dout <= 8'b10101001; //   18 : 169 - 0xa9
      10'h13: dout <= 8'b10101001; //   19 : 169 - 0xa9
      10'h14: dout <= 8'b10101001; //   20 : 169 - 0xa9
      10'h15: dout <= 8'b10101001; //   21 : 169 - 0xa9
      10'h16: dout <= 8'b10101001; //   22 : 169 - 0xa9
      10'h17: dout <= 8'b10101001; //   23 : 169 - 0xa9
      10'h18: dout <= 8'b10101001; //   24 : 169 - 0xa9
      10'h19: dout <= 8'b10101001; //   25 : 169 - 0xa9
      10'h1A: dout <= 8'b10101001; //   26 : 169 - 0xa9
      10'h1B: dout <= 8'b10101001; //   27 : 169 - 0xa9
      10'h1C: dout <= 8'b10101001; //   28 : 169 - 0xa9
      10'h1D: dout <= 8'b10101001; //   29 : 169 - 0xa9
      10'h1E: dout <= 8'b10101001; //   30 : 169 - 0xa9
      10'h1F: dout <= 8'b10101001; //   31 : 169 - 0xa9
      10'h20: dout <= 8'b10101001; //   32 : 169 - 0xa9 -- line 0x1
      10'h21: dout <= 8'b10101001; //   33 : 169 - 0xa9
      10'h22: dout <= 8'b10101001; //   34 : 169 - 0xa9
      10'h23: dout <= 8'b10101001; //   35 : 169 - 0xa9
      10'h24: dout <= 8'b10101001; //   36 : 169 - 0xa9
      10'h25: dout <= 8'b10101001; //   37 : 169 - 0xa9
      10'h26: dout <= 8'b10101001; //   38 : 169 - 0xa9
      10'h27: dout <= 8'b10101001; //   39 : 169 - 0xa9
      10'h28: dout <= 8'b10101001; //   40 : 169 - 0xa9
      10'h29: dout <= 8'b10101001; //   41 : 169 - 0xa9
      10'h2A: dout <= 8'b10101001; //   42 : 169 - 0xa9
      10'h2B: dout <= 8'b10101001; //   43 : 169 - 0xa9
      10'h2C: dout <= 8'b10101001; //   44 : 169 - 0xa9
      10'h2D: dout <= 8'b10101001; //   45 : 169 - 0xa9
      10'h2E: dout <= 8'b10101001; //   46 : 169 - 0xa9
      10'h2F: dout <= 8'b10101001; //   47 : 169 - 0xa9
      10'h30: dout <= 8'b10101001; //   48 : 169 - 0xa9
      10'h31: dout <= 8'b10101001; //   49 : 169 - 0xa9
      10'h32: dout <= 8'b10101001; //   50 : 169 - 0xa9
      10'h33: dout <= 8'b10101001; //   51 : 169 - 0xa9
      10'h34: dout <= 8'b10101001; //   52 : 169 - 0xa9
      10'h35: dout <= 8'b10101001; //   53 : 169 - 0xa9
      10'h36: dout <= 8'b10101001; //   54 : 169 - 0xa9
      10'h37: dout <= 8'b10101001; //   55 : 169 - 0xa9
      10'h38: dout <= 8'b10101001; //   56 : 169 - 0xa9
      10'h39: dout <= 8'b10101001; //   57 : 169 - 0xa9
      10'h3A: dout <= 8'b10101001; //   58 : 169 - 0xa9
      10'h3B: dout <= 8'b10101001; //   59 : 169 - 0xa9
      10'h3C: dout <= 8'b10101001; //   60 : 169 - 0xa9
      10'h3D: dout <= 8'b10101001; //   61 : 169 - 0xa9
      10'h3E: dout <= 8'b10101001; //   62 : 169 - 0xa9
      10'h3F: dout <= 8'b10101001; //   63 : 169 - 0xa9
      10'h40: dout <= 8'b10101001; //   64 : 169 - 0xa9 -- line 0x2
      10'h41: dout <= 8'b10101001; //   65 : 169 - 0xa9
      10'h42: dout <= 8'b01010110; //   66 :  86 - 0x56
      10'h43: dout <= 8'b01010101; //   67 :  85 - 0x55
      10'h44: dout <= 8'b01010111; //   68 :  87 - 0x57
      10'h45: dout <= 8'b01011000; //   69 :  88 - 0x58
      10'h46: dout <= 8'b11010000; //   70 : 208 - 0xd0
      10'h47: dout <= 8'b11010001; //   71 : 209 - 0xd1
      10'h48: dout <= 8'b10101001; //   72 : 169 - 0xa9
      10'h49: dout <= 8'b01011101; //   73 :  93 - 0x5d
      10'h4A: dout <= 8'b01011110; //   74 :  94 - 0x5e
      10'h4B: dout <= 8'b01011011; //   75 :  91 - 0x5b
      10'h4C: dout <= 8'b01010110; //   76 :  86 - 0x56
      10'h4D: dout <= 8'b11111001; //   77 : 249 - 0xf9
      10'h4E: dout <= 8'b11111010; //   78 : 250 - 0xfa
      10'h4F: dout <= 8'b11111010; //   79 : 250 - 0xfa
      10'h50: dout <= 8'b11111010; //   80 : 250 - 0xfa
      10'h51: dout <= 8'b11111010; //   81 : 250 - 0xfa
      10'h52: dout <= 8'b11111010; //   82 : 250 - 0xfa
      10'h53: dout <= 8'b11111010; //   83 : 250 - 0xfa
      10'h54: dout <= 8'b11111011; //   84 : 251 - 0xfb
      10'h55: dout <= 8'b10101001; //   85 : 169 - 0xa9
      10'h56: dout <= 8'b01011001; //   86 :  89 - 0x59
      10'h57: dout <= 8'b01011010; //   87 :  90 - 0x5a
      10'h58: dout <= 8'b01011000; //   88 :  88 - 0x58
      10'h59: dout <= 8'b01011011; //   89 :  91 - 0x5b
      10'h5A: dout <= 8'b11010000; //   90 : 208 - 0xd0
      10'h5B: dout <= 8'b11010000; //   91 : 208 - 0xd0
      10'h5C: dout <= 8'b11010000; //   92 : 208 - 0xd0
      10'h5D: dout <= 8'b01011100; //   93 :  92 - 0x5c
      10'h5E: dout <= 8'b10101001; //   94 : 169 - 0xa9
      10'h5F: dout <= 8'b10101001; //   95 : 169 - 0xa9
      10'h60: dout <= 8'b10101001; //   96 : 169 - 0xa9 -- line 0x3
      10'h61: dout <= 8'b10101001; //   97 : 169 - 0xa9
      10'h62: dout <= 8'b01100110; //   98 : 102 - 0x66
      10'h63: dout <= 8'b01100101; //   99 : 101 - 0x65
      10'h64: dout <= 8'b01100111; //  100 : 103 - 0x67
      10'h65: dout <= 8'b01101000; //  101 : 104 - 0x68
      10'h66: dout <= 8'b11100000; //  102 : 224 - 0xe0
      10'h67: dout <= 8'b11100001; //  103 : 225 - 0xe1
      10'h68: dout <= 8'b10101001; //  104 : 169 - 0xa9
      10'h69: dout <= 8'b01101101; //  105 : 109 - 0x6d
      10'h6A: dout <= 8'b01101110; //  106 : 110 - 0x6e
      10'h6B: dout <= 8'b01101011; //  107 : 107 - 0x6b
      10'h6C: dout <= 8'b01100110; //  108 : 102 - 0x66
      10'h6D: dout <= 8'b11111100; //  109 : 252 - 0xfc
      10'h6E: dout <= 8'b11111101; //  110 : 253 - 0xfd
      10'h6F: dout <= 8'b11111101; //  111 : 253 - 0xfd
      10'h70: dout <= 8'b11111101; //  112 : 253 - 0xfd
      10'h71: dout <= 8'b11111101; //  113 : 253 - 0xfd
      10'h72: dout <= 8'b11111101; //  114 : 253 - 0xfd
      10'h73: dout <= 8'b11111101; //  115 : 253 - 0xfd
      10'h74: dout <= 8'b11111110; //  116 : 254 - 0xfe
      10'h75: dout <= 8'b10101001; //  117 : 169 - 0xa9
      10'h76: dout <= 8'b01101001; //  118 : 105 - 0x69
      10'h77: dout <= 8'b01101010; //  119 : 106 - 0x6a
      10'h78: dout <= 8'b01101000; //  120 : 104 - 0x68
      10'h79: dout <= 8'b01101011; //  121 : 107 - 0x6b
      10'h7A: dout <= 8'b11100000; //  122 : 224 - 0xe0
      10'h7B: dout <= 8'b11100000; //  123 : 224 - 0xe0
      10'h7C: dout <= 8'b11100000; //  124 : 224 - 0xe0
      10'h7D: dout <= 8'b01101100; //  125 : 108 - 0x6c
      10'h7E: dout <= 8'b10101001; //  126 : 169 - 0xa9
      10'h7F: dout <= 8'b10101001; //  127 : 169 - 0xa9
      10'h80: dout <= 8'b10101010; //  128 : 170 - 0xaa -- line 0x4
      10'h81: dout <= 8'b10101010; //  129 : 170 - 0xaa
      10'h82: dout <= 8'b10101010; //  130 : 170 - 0xaa
      10'h83: dout <= 8'b10101010; //  131 : 170 - 0xaa
      10'h84: dout <= 8'b10101010; //  132 : 170 - 0xaa
      10'h85: dout <= 8'b10101010; //  133 : 170 - 0xaa
      10'h86: dout <= 8'b10101010; //  134 : 170 - 0xaa
      10'h87: dout <= 8'b10101010; //  135 : 170 - 0xaa
      10'h88: dout <= 8'b10101010; //  136 : 170 - 0xaa
      10'h89: dout <= 8'b10101010; //  137 : 170 - 0xaa
      10'h8A: dout <= 8'b10101010; //  138 : 170 - 0xaa
      10'h8B: dout <= 8'b10101010; //  139 : 170 - 0xaa
      10'h8C: dout <= 8'b10101010; //  140 : 170 - 0xaa
      10'h8D: dout <= 8'b10101010; //  141 : 170 - 0xaa
      10'h8E: dout <= 8'b10101010; //  142 : 170 - 0xaa
      10'h8F: dout <= 8'b10101010; //  143 : 170 - 0xaa
      10'h90: dout <= 8'b10101010; //  144 : 170 - 0xaa
      10'h91: dout <= 8'b10101010; //  145 : 170 - 0xaa
      10'h92: dout <= 8'b10101010; //  146 : 170 - 0xaa
      10'h93: dout <= 8'b10101010; //  147 : 170 - 0xaa
      10'h94: dout <= 8'b10101010; //  148 : 170 - 0xaa
      10'h95: dout <= 8'b10101010; //  149 : 170 - 0xaa
      10'h96: dout <= 8'b10101010; //  150 : 170 - 0xaa
      10'h97: dout <= 8'b10101010; //  151 : 170 - 0xaa
      10'h98: dout <= 8'b10101010; //  152 : 170 - 0xaa
      10'h99: dout <= 8'b10101010; //  153 : 170 - 0xaa
      10'h9A: dout <= 8'b10101010; //  154 : 170 - 0xaa
      10'h9B: dout <= 8'b10101010; //  155 : 170 - 0xaa
      10'h9C: dout <= 8'b10101010; //  156 : 170 - 0xaa
      10'h9D: dout <= 8'b10101010; //  157 : 170 - 0xaa
      10'h9E: dout <= 8'b10101010; //  158 : 170 - 0xaa
      10'h9F: dout <= 8'b10101010; //  159 : 170 - 0xaa
      10'hA0: dout <= 8'b10100000; //  160 : 160 - 0xa0 -- line 0x5
      10'hA1: dout <= 8'b10100001; //  161 : 161 - 0xa1
      10'hA2: dout <= 8'b10100010; //  162 : 162 - 0xa2
      10'hA3: dout <= 8'b10100010; //  163 : 162 - 0xa2
      10'hA4: dout <= 8'b10100010; //  164 : 162 - 0xa2
      10'hA5: dout <= 8'b10100010; //  165 : 162 - 0xa2
      10'hA6: dout <= 8'b10100010; //  166 : 162 - 0xa2
      10'hA7: dout <= 8'b10100010; //  167 : 162 - 0xa2
      10'hA8: dout <= 8'b10100010; //  168 : 162 - 0xa2
      10'hA9: dout <= 8'b10100010; //  169 : 162 - 0xa2
      10'hAA: dout <= 8'b10100010; //  170 : 162 - 0xa2
      10'hAB: dout <= 8'b10100010; //  171 : 162 - 0xa2
      10'hAC: dout <= 8'b10100010; //  172 : 162 - 0xa2
      10'hAD: dout <= 8'b10100010; //  173 : 162 - 0xa2
      10'hAE: dout <= 8'b10100010; //  174 : 162 - 0xa2
      10'hAF: dout <= 8'b10100010; //  175 : 162 - 0xa2
      10'hB0: dout <= 8'b10100010; //  176 : 162 - 0xa2
      10'hB1: dout <= 8'b10100010; //  177 : 162 - 0xa2
      10'hB2: dout <= 8'b10100010; //  178 : 162 - 0xa2
      10'hB3: dout <= 8'b10100010; //  179 : 162 - 0xa2
      10'hB4: dout <= 8'b10100010; //  180 : 162 - 0xa2
      10'hB5: dout <= 8'b10100010; //  181 : 162 - 0xa2
      10'hB6: dout <= 8'b10100010; //  182 : 162 - 0xa2
      10'hB7: dout <= 8'b10100010; //  183 : 162 - 0xa2
      10'hB8: dout <= 8'b10100010; //  184 : 162 - 0xa2
      10'hB9: dout <= 8'b10100010; //  185 : 162 - 0xa2
      10'hBA: dout <= 8'b10100010; //  186 : 162 - 0xa2
      10'hBB: dout <= 8'b10100010; //  187 : 162 - 0xa2
      10'hBC: dout <= 8'b10100010; //  188 : 162 - 0xa2
      10'hBD: dout <= 8'b10100010; //  189 : 162 - 0xa2
      10'hBE: dout <= 8'b10100110; //  190 : 166 - 0xa6
      10'hBF: dout <= 8'b10100000; //  191 : 160 - 0xa0
      10'hC0: dout <= 8'b10100000; //  192 : 160 - 0xa0 -- line 0x6
      10'hC1: dout <= 8'b10100011; //  193 : 163 - 0xa3
      10'hC2: dout <= 8'b10000000; //  194 : 128 - 0x80
      10'hC3: dout <= 8'b10000001; //  195 : 129 - 0x81
      10'hC4: dout <= 8'b10000000; //  196 : 128 - 0x80
      10'hC5: dout <= 8'b10000001; //  197 : 129 - 0x81
      10'hC6: dout <= 8'b10000000; //  198 : 128 - 0x80
      10'hC7: dout <= 8'b10000010; //  199 : 130 - 0x82
      10'hC8: dout <= 8'b10000000; //  200 : 128 - 0x80
      10'hC9: dout <= 8'b10000001; //  201 : 129 - 0x81
      10'hCA: dout <= 8'b10000001; //  202 : 129 - 0x81
      10'hCB: dout <= 8'b10000000; //  203 : 128 - 0x80
      10'hCC: dout <= 8'b10000000; //  204 : 128 - 0x80
      10'hCD: dout <= 8'b10000001; //  205 : 129 - 0x81
      10'hCE: dout <= 8'b10000010; //  206 : 130 - 0x82
      10'hCF: dout <= 8'b10000011; //  207 : 131 - 0x83
      10'hD0: dout <= 8'b10000010; //  208 : 130 - 0x82
      10'hD1: dout <= 8'b10000011; //  209 : 131 - 0x83
      10'hD2: dout <= 8'b10000000; //  210 : 128 - 0x80
      10'hD3: dout <= 8'b10000010; //  211 : 130 - 0x82
      10'hD4: dout <= 8'b10000000; //  212 : 128 - 0x80
      10'hD5: dout <= 8'b10000010; //  213 : 130 - 0x82
      10'hD6: dout <= 8'b10000010; //  214 : 130 - 0x82
      10'hD7: dout <= 8'b10000011; //  215 : 131 - 0x83
      10'hD8: dout <= 8'b10000010; //  216 : 130 - 0x82
      10'hD9: dout <= 8'b10000011; //  217 : 131 - 0x83
      10'hDA: dout <= 8'b10000001; //  218 : 129 - 0x81
      10'hDB: dout <= 8'b10000000; //  219 : 128 - 0x80
      10'hDC: dout <= 8'b10000000; //  220 : 128 - 0x80
      10'hDD: dout <= 8'b10000001; //  221 : 129 - 0x81
      10'hDE: dout <= 8'b10100111; //  222 : 167 - 0xa7
      10'hDF: dout <= 8'b10100000; //  223 : 160 - 0xa0
      10'hE0: dout <= 8'b10100000; //  224 : 160 - 0xa0 -- line 0x7
      10'hE1: dout <= 8'b10100011; //  225 : 163 - 0xa3
      10'hE2: dout <= 8'b10010000; //  226 : 144 - 0x90
      10'hE3: dout <= 8'b10010001; //  227 : 145 - 0x91
      10'hE4: dout <= 8'b10010000; //  228 : 144 - 0x90
      10'hE5: dout <= 8'b10010001; //  229 : 145 - 0x91
      10'hE6: dout <= 8'b10010010; //  230 : 146 - 0x92
      10'hE7: dout <= 8'b10010001; //  231 : 145 - 0x91
      10'hE8: dout <= 8'b10010000; //  232 : 144 - 0x90
      10'hE9: dout <= 8'b10010001; //  233 : 145 - 0x91
      10'hEA: dout <= 8'b10010011; //  234 : 147 - 0x93
      10'hEB: dout <= 8'b10010010; //  235 : 146 - 0x92
      10'hEC: dout <= 8'b10010000; //  236 : 144 - 0x90
      10'hED: dout <= 8'b10010001; //  237 : 145 - 0x91
      10'hEE: dout <= 8'b10010010; //  238 : 146 - 0x92
      10'hEF: dout <= 8'b10010011; //  239 : 147 - 0x93
      10'hF0: dout <= 8'b10010010; //  240 : 146 - 0x92
      10'hF1: dout <= 8'b10010011; //  241 : 147 - 0x93
      10'hF2: dout <= 8'b10010010; //  242 : 146 - 0x92
      10'hF3: dout <= 8'b10010001; //  243 : 145 - 0x91
      10'hF4: dout <= 8'b10010010; //  244 : 146 - 0x92
      10'hF5: dout <= 8'b10010001; //  245 : 145 - 0x91
      10'hF6: dout <= 8'b10010010; //  246 : 146 - 0x92
      10'hF7: dout <= 8'b10010011; //  247 : 147 - 0x93
      10'hF8: dout <= 8'b10010010; //  248 : 146 - 0x92
      10'hF9: dout <= 8'b10010011; //  249 : 147 - 0x93
      10'hFA: dout <= 8'b10010011; //  250 : 147 - 0x93
      10'hFB: dout <= 8'b10010010; //  251 : 146 - 0x92
      10'hFC: dout <= 8'b10010000; //  252 : 144 - 0x90
      10'hFD: dout <= 8'b10010001; //  253 : 145 - 0x91
      10'hFE: dout <= 8'b10100111; //  254 : 167 - 0xa7
      10'hFF: dout <= 8'b10100000; //  255 : 160 - 0xa0
      10'h100: dout <= 8'b10100000; //  256 : 160 - 0xa0 -- line 0x8
      10'h101: dout <= 8'b10100011; //  257 : 163 - 0xa3
      10'h102: dout <= 8'b10000010; //  258 : 130 - 0x82
      10'h103: dout <= 8'b10000011; //  259 : 131 - 0x83
      10'h104: dout <= 8'b10000101; //  260 : 133 - 0x85
      10'h105: dout <= 8'b10000110; //  261 : 134 - 0x86
      10'h106: dout <= 8'b10000101; //  262 : 133 - 0x85
      10'h107: dout <= 8'b10000110; //  263 : 134 - 0x86
      10'h108: dout <= 8'b10000101; //  264 : 133 - 0x85
      10'h109: dout <= 8'b10000110; //  265 : 134 - 0x86
      10'h10A: dout <= 8'b10000101; //  266 : 133 - 0x85
      10'h10B: dout <= 8'b10000110; //  267 : 134 - 0x86
      10'h10C: dout <= 8'b10000100; //  268 : 132 - 0x84
      10'h10D: dout <= 8'b10000111; //  269 : 135 - 0x87
      10'h10E: dout <= 8'b10000110; //  270 : 134 - 0x86
      10'h10F: dout <= 8'b10000111; //  271 : 135 - 0x87
      10'h110: dout <= 8'b10000100; //  272 : 132 - 0x84
      10'h111: dout <= 8'b10000101; //  273 : 133 - 0x85
      10'h112: dout <= 8'b10000101; //  274 : 133 - 0x85
      10'h113: dout <= 8'b10000110; //  275 : 134 - 0x86
      10'h114: dout <= 8'b10000101; //  276 : 133 - 0x85
      10'h115: dout <= 8'b10000110; //  277 : 134 - 0x86
      10'h116: dout <= 8'b10000110; //  278 : 134 - 0x86
      10'h117: dout <= 8'b10000111; //  279 : 135 - 0x87
      10'h118: dout <= 8'b10000110; //  280 : 134 - 0x86
      10'h119: dout <= 8'b10000111; //  281 : 135 - 0x87
      10'h11A: dout <= 8'b10000100; //  282 : 132 - 0x84
      10'h11B: dout <= 8'b10000101; //  283 : 133 - 0x85
      10'h11C: dout <= 8'b10000010; //  284 : 130 - 0x82
      10'h11D: dout <= 8'b10000011; //  285 : 131 - 0x83
      10'h11E: dout <= 8'b10100111; //  286 : 167 - 0xa7
      10'h11F: dout <= 8'b10100000; //  287 : 160 - 0xa0
      10'h120: dout <= 8'b10100000; //  288 : 160 - 0xa0 -- line 0x9
      10'h121: dout <= 8'b10100011; //  289 : 163 - 0xa3
      10'h122: dout <= 8'b10010010; //  290 : 146 - 0x92
      10'h123: dout <= 8'b10010011; //  291 : 147 - 0x93
      10'h124: dout <= 8'b10010111; //  292 : 151 - 0x97
      10'h125: dout <= 8'b10010100; //  293 : 148 - 0x94
      10'h126: dout <= 8'b10010111; //  294 : 151 - 0x97
      10'h127: dout <= 8'b10010100; //  295 : 148 - 0x94
      10'h128: dout <= 8'b10010111; //  296 : 151 - 0x97
      10'h129: dout <= 8'b10010100; //  297 : 148 - 0x94
      10'h12A: dout <= 8'b10010111; //  298 : 151 - 0x97
      10'h12B: dout <= 8'b10010100; //  299 : 148 - 0x94
      10'h12C: dout <= 8'b10010110; //  300 : 150 - 0x96
      10'h12D: dout <= 8'b10010101; //  301 : 149 - 0x95
      10'h12E: dout <= 8'b10010110; //  302 : 150 - 0x96
      10'h12F: dout <= 8'b10010111; //  303 : 151 - 0x97
      10'h130: dout <= 8'b10010100; //  304 : 148 - 0x94
      10'h131: dout <= 8'b10010101; //  305 : 149 - 0x95
      10'h132: dout <= 8'b10010111; //  306 : 151 - 0x97
      10'h133: dout <= 8'b10010100; //  307 : 148 - 0x94
      10'h134: dout <= 8'b10010111; //  308 : 151 - 0x97
      10'h135: dout <= 8'b10010100; //  309 : 148 - 0x94
      10'h136: dout <= 8'b10010110; //  310 : 150 - 0x96
      10'h137: dout <= 8'b10010111; //  311 : 151 - 0x97
      10'h138: dout <= 8'b10010110; //  312 : 150 - 0x96
      10'h139: dout <= 8'b10010111; //  313 : 151 - 0x97
      10'h13A: dout <= 8'b10010100; //  314 : 148 - 0x94
      10'h13B: dout <= 8'b10010101; //  315 : 149 - 0x95
      10'h13C: dout <= 8'b10010010; //  316 : 146 - 0x92
      10'h13D: dout <= 8'b10010011; //  317 : 147 - 0x93
      10'h13E: dout <= 8'b10100111; //  318 : 167 - 0xa7
      10'h13F: dout <= 8'b10100000; //  319 : 160 - 0xa0
      10'h140: dout <= 8'b10100000; //  320 : 160 - 0xa0 -- line 0xa
      10'h141: dout <= 8'b10100011; //  321 : 163 - 0xa3
      10'h142: dout <= 8'b10000000; //  322 : 128 - 0x80
      10'h143: dout <= 8'b10000010; //  323 : 130 - 0x82
      10'h144: dout <= 8'b10000100; //  324 : 132 - 0x84
      10'h145: dout <= 8'b10000111; //  325 : 135 - 0x87
      10'h146: dout <= 8'b10000101; //  326 : 133 - 0x85
      10'h147: dout <= 8'b10000110; //  327 : 134 - 0x86
      10'h148: dout <= 8'b10000100; //  328 : 132 - 0x84
      10'h149: dout <= 8'b10000111; //  329 : 135 - 0x87
      10'h14A: dout <= 8'b10000100; //  330 : 132 - 0x84
      10'h14B: dout <= 8'b10000111; //  331 : 135 - 0x87
      10'h14C: dout <= 8'b10000110; //  332 : 134 - 0x86
      10'h14D: dout <= 8'b10000111; //  333 : 135 - 0x87
      10'h14E: dout <= 8'b10000100; //  334 : 132 - 0x84
      10'h14F: dout <= 8'b10000101; //  335 : 133 - 0x85
      10'h150: dout <= 8'b10000100; //  336 : 132 - 0x84
      10'h151: dout <= 8'b10000101; //  337 : 133 - 0x85
      10'h152: dout <= 8'b10000110; //  338 : 134 - 0x86
      10'h153: dout <= 8'b10000111; //  339 : 135 - 0x87
      10'h154: dout <= 8'b10000100; //  340 : 132 - 0x84
      10'h155: dout <= 8'b10000101; //  341 : 133 - 0x85
      10'h156: dout <= 8'b10000101; //  342 : 133 - 0x85
      10'h157: dout <= 8'b10000110; //  343 : 134 - 0x86
      10'h158: dout <= 8'b10000100; //  344 : 132 - 0x84
      10'h159: dout <= 8'b10000111; //  345 : 135 - 0x87
      10'h15A: dout <= 8'b10000100; //  346 : 132 - 0x84
      10'h15B: dout <= 8'b10000111; //  347 : 135 - 0x87
      10'h15C: dout <= 8'b10000000; //  348 : 128 - 0x80
      10'h15D: dout <= 8'b10000001; //  349 : 129 - 0x81
      10'h15E: dout <= 8'b10100111; //  350 : 167 - 0xa7
      10'h15F: dout <= 8'b10100000; //  351 : 160 - 0xa0
      10'h160: dout <= 8'b10100000; //  352 : 160 - 0xa0 -- line 0xb
      10'h161: dout <= 8'b10100011; //  353 : 163 - 0xa3
      10'h162: dout <= 8'b10010010; //  354 : 146 - 0x92
      10'h163: dout <= 8'b10010001; //  355 : 145 - 0x91
      10'h164: dout <= 8'b10010110; //  356 : 150 - 0x96
      10'h165: dout <= 8'b10010101; //  357 : 149 - 0x95
      10'h166: dout <= 8'b10010111; //  358 : 151 - 0x97
      10'h167: dout <= 8'b10010100; //  359 : 148 - 0x94
      10'h168: dout <= 8'b10010110; //  360 : 150 - 0x96
      10'h169: dout <= 8'b10010101; //  361 : 149 - 0x95
      10'h16A: dout <= 8'b10010110; //  362 : 150 - 0x96
      10'h16B: dout <= 8'b10010101; //  363 : 149 - 0x95
      10'h16C: dout <= 8'b10010110; //  364 : 150 - 0x96
      10'h16D: dout <= 8'b10010111; //  365 : 151 - 0x97
      10'h16E: dout <= 8'b10010100; //  366 : 148 - 0x94
      10'h16F: dout <= 8'b10010101; //  367 : 149 - 0x95
      10'h170: dout <= 8'b10010100; //  368 : 148 - 0x94
      10'h171: dout <= 8'b10010101; //  369 : 149 - 0x95
      10'h172: dout <= 8'b10010110; //  370 : 150 - 0x96
      10'h173: dout <= 8'b10010111; //  371 : 151 - 0x97
      10'h174: dout <= 8'b10010100; //  372 : 148 - 0x94
      10'h175: dout <= 8'b10010101; //  373 : 149 - 0x95
      10'h176: dout <= 8'b10010111; //  374 : 151 - 0x97
      10'h177: dout <= 8'b10010100; //  375 : 148 - 0x94
      10'h178: dout <= 8'b10010110; //  376 : 150 - 0x96
      10'h179: dout <= 8'b10010101; //  377 : 149 - 0x95
      10'h17A: dout <= 8'b10010110; //  378 : 150 - 0x96
      10'h17B: dout <= 8'b10010101; //  379 : 149 - 0x95
      10'h17C: dout <= 8'b10010000; //  380 : 144 - 0x90
      10'h17D: dout <= 8'b10010001; //  381 : 145 - 0x91
      10'h17E: dout <= 8'b10100111; //  382 : 167 - 0xa7
      10'h17F: dout <= 8'b10100000; //  383 : 160 - 0xa0
      10'h180: dout <= 8'b10100000; //  384 : 160 - 0xa0 -- line 0xc
      10'h181: dout <= 8'b10100011; //  385 : 163 - 0xa3
      10'h182: dout <= 8'b10000010; //  386 : 130 - 0x82
      10'h183: dout <= 8'b10000011; //  387 : 131 - 0x83
      10'h184: dout <= 8'b10000110; //  388 : 134 - 0x86
      10'h185: dout <= 8'b10000111; //  389 : 135 - 0x87
      10'h186: dout <= 8'b10000100; //  390 : 132 - 0x84
      10'h187: dout <= 8'b10000101; //  391 : 133 - 0x85
      10'h188: dout <= 8'b10000100; //  392 : 132 - 0x84
      10'h189: dout <= 8'b10000111; //  393 : 135 - 0x87
      10'h18A: dout <= 8'b10000100; //  394 : 132 - 0x84
      10'h18B: dout <= 8'b10000111; //  395 : 135 - 0x87
      10'h18C: dout <= 8'b10000110; //  396 : 134 - 0x86
      10'h18D: dout <= 8'b10000111; //  397 : 135 - 0x87
      10'h18E: dout <= 8'b10000100; //  398 : 132 - 0x84
      10'h18F: dout <= 8'b10000111; //  399 : 135 - 0x87
      10'h190: dout <= 8'b10000110; //  400 : 134 - 0x86
      10'h191: dout <= 8'b10000111; //  401 : 135 - 0x87
      10'h192: dout <= 8'b10000110; //  402 : 134 - 0x86
      10'h193: dout <= 8'b10000111; //  403 : 135 - 0x87
      10'h194: dout <= 8'b10000110; //  404 : 134 - 0x86
      10'h195: dout <= 8'b10000111; //  405 : 135 - 0x87
      10'h196: dout <= 8'b10000110; //  406 : 134 - 0x86
      10'h197: dout <= 8'b10000111; //  407 : 135 - 0x87
      10'h198: dout <= 8'b10000101; //  408 : 133 - 0x85
      10'h199: dout <= 8'b10000110; //  409 : 134 - 0x86
      10'h19A: dout <= 8'b10000100; //  410 : 132 - 0x84
      10'h19B: dout <= 8'b10000111; //  411 : 135 - 0x87
      10'h19C: dout <= 8'b10000000; //  412 : 128 - 0x80
      10'h19D: dout <= 8'b10000010; //  413 : 130 - 0x82
      10'h19E: dout <= 8'b10100111; //  414 : 167 - 0xa7
      10'h19F: dout <= 8'b10100000; //  415 : 160 - 0xa0
      10'h1A0: dout <= 8'b10100000; //  416 : 160 - 0xa0 -- line 0xd
      10'h1A1: dout <= 8'b10100011; //  417 : 163 - 0xa3
      10'h1A2: dout <= 8'b10010010; //  418 : 146 - 0x92
      10'h1A3: dout <= 8'b10010011; //  419 : 147 - 0x93
      10'h1A4: dout <= 8'b10010110; //  420 : 150 - 0x96
      10'h1A5: dout <= 8'b10010111; //  421 : 151 - 0x97
      10'h1A6: dout <= 8'b10010100; //  422 : 148 - 0x94
      10'h1A7: dout <= 8'b10010101; //  423 : 149 - 0x95
      10'h1A8: dout <= 8'b10010110; //  424 : 150 - 0x96
      10'h1A9: dout <= 8'b10010101; //  425 : 149 - 0x95
      10'h1AA: dout <= 8'b10010110; //  426 : 150 - 0x96
      10'h1AB: dout <= 8'b10010101; //  427 : 149 - 0x95
      10'h1AC: dout <= 8'b10010110; //  428 : 150 - 0x96
      10'h1AD: dout <= 8'b10010111; //  429 : 151 - 0x97
      10'h1AE: dout <= 8'b10010110; //  430 : 150 - 0x96
      10'h1AF: dout <= 8'b10010101; //  431 : 149 - 0x95
      10'h1B0: dout <= 8'b10010110; //  432 : 150 - 0x96
      10'h1B1: dout <= 8'b10010111; //  433 : 151 - 0x97
      10'h1B2: dout <= 8'b10010110; //  434 : 150 - 0x96
      10'h1B3: dout <= 8'b10010111; //  435 : 151 - 0x97
      10'h1B4: dout <= 8'b10010110; //  436 : 150 - 0x96
      10'h1B5: dout <= 8'b10010111; //  437 : 151 - 0x97
      10'h1B6: dout <= 8'b10010110; //  438 : 150 - 0x96
      10'h1B7: dout <= 8'b10010111; //  439 : 151 - 0x97
      10'h1B8: dout <= 8'b10010111; //  440 : 151 - 0x97
      10'h1B9: dout <= 8'b10010100; //  441 : 148 - 0x94
      10'h1BA: dout <= 8'b10010110; //  442 : 150 - 0x96
      10'h1BB: dout <= 8'b10010101; //  443 : 149 - 0x95
      10'h1BC: dout <= 8'b10010010; //  444 : 146 - 0x92
      10'h1BD: dout <= 8'b10010001; //  445 : 145 - 0x91
      10'h1BE: dout <= 8'b10100111; //  446 : 167 - 0xa7
      10'h1BF: dout <= 8'b10100000; //  447 : 160 - 0xa0
      10'h1C0: dout <= 8'b10100000; //  448 : 160 - 0xa0 -- line 0xe
      10'h1C1: dout <= 8'b10100011; //  449 : 163 - 0xa3
      10'h1C2: dout <= 8'b10000000; //  450 : 128 - 0x80
      10'h1C3: dout <= 8'b10000001; //  451 : 129 - 0x81
      10'h1C4: dout <= 8'b10000101; //  452 : 133 - 0x85
      10'h1C5: dout <= 8'b10000110; //  453 : 134 - 0x86
      10'h1C6: dout <= 8'b10000100; //  454 : 132 - 0x84
      10'h1C7: dout <= 8'b10000101; //  455 : 133 - 0x85
      10'h1C8: dout <= 8'b10000100; //  456 : 132 - 0x84
      10'h1C9: dout <= 8'b10000101; //  457 : 133 - 0x85
      10'h1CA: dout <= 8'b10000100; //  458 : 132 - 0x84
      10'h1CB: dout <= 8'b10000111; //  459 : 135 - 0x87
      10'h1CC: dout <= 8'b10000001; //  460 : 129 - 0x81
      10'h1CD: dout <= 8'b10000000; //  461 : 128 - 0x80
      10'h1CE: dout <= 8'b10000010; //  462 : 130 - 0x82
      10'h1CF: dout <= 8'b10000011; //  463 : 131 - 0x83
      10'h1D0: dout <= 8'b10000010; //  464 : 130 - 0x82
      10'h1D1: dout <= 8'b10000011; //  465 : 131 - 0x83
      10'h1D2: dout <= 8'b10000001; //  466 : 129 - 0x81
      10'h1D3: dout <= 8'b10000000; //  467 : 128 - 0x80
      10'h1D4: dout <= 8'b10000101; //  468 : 133 - 0x85
      10'h1D5: dout <= 8'b10000110; //  469 : 134 - 0x86
      10'h1D6: dout <= 8'b10000110; //  470 : 134 - 0x86
      10'h1D7: dout <= 8'b10000111; //  471 : 135 - 0x87
      10'h1D8: dout <= 8'b10000100; //  472 : 132 - 0x84
      10'h1D9: dout <= 8'b10000111; //  473 : 135 - 0x87
      10'h1DA: dout <= 8'b10000100; //  474 : 132 - 0x84
      10'h1DB: dout <= 8'b10000111; //  475 : 135 - 0x87
      10'h1DC: dout <= 8'b10000000; //  476 : 128 - 0x80
      10'h1DD: dout <= 8'b10000001; //  477 : 129 - 0x81
      10'h1DE: dout <= 8'b10100111; //  478 : 167 - 0xa7
      10'h1DF: dout <= 8'b10100000; //  479 : 160 - 0xa0
      10'h1E0: dout <= 8'b10100000; //  480 : 160 - 0xa0 -- line 0xf
      10'h1E1: dout <= 8'b10100011; //  481 : 163 - 0xa3
      10'h1E2: dout <= 8'b10010000; //  482 : 144 - 0x90
      10'h1E3: dout <= 8'b10010001; //  483 : 145 - 0x91
      10'h1E4: dout <= 8'b10010111; //  484 : 151 - 0x97
      10'h1E5: dout <= 8'b10010100; //  485 : 148 - 0x94
      10'h1E6: dout <= 8'b10010100; //  486 : 148 - 0x94
      10'h1E7: dout <= 8'b10010101; //  487 : 149 - 0x95
      10'h1E8: dout <= 8'b10010100; //  488 : 148 - 0x94
      10'h1E9: dout <= 8'b10010101; //  489 : 149 - 0x95
      10'h1EA: dout <= 8'b10010110; //  490 : 150 - 0x96
      10'h1EB: dout <= 8'b10010101; //  491 : 149 - 0x95
      10'h1EC: dout <= 8'b10010011; //  492 : 147 - 0x93
      10'h1ED: dout <= 8'b10010010; //  493 : 146 - 0x92
      10'h1EE: dout <= 8'b10010010; //  494 : 146 - 0x92
      10'h1EF: dout <= 8'b10010011; //  495 : 147 - 0x93
      10'h1F0: dout <= 8'b10010010; //  496 : 146 - 0x92
      10'h1F1: dout <= 8'b10010011; //  497 : 147 - 0x93
      10'h1F2: dout <= 8'b10010011; //  498 : 147 - 0x93
      10'h1F3: dout <= 8'b10010010; //  499 : 146 - 0x92
      10'h1F4: dout <= 8'b10010111; //  500 : 151 - 0x97
      10'h1F5: dout <= 8'b10010100; //  501 : 148 - 0x94
      10'h1F6: dout <= 8'b10010110; //  502 : 150 - 0x96
      10'h1F7: dout <= 8'b10010111; //  503 : 151 - 0x97
      10'h1F8: dout <= 8'b10010110; //  504 : 150 - 0x96
      10'h1F9: dout <= 8'b10010101; //  505 : 149 - 0x95
      10'h1FA: dout <= 8'b10010110; //  506 : 150 - 0x96
      10'h1FB: dout <= 8'b10010101; //  507 : 149 - 0x95
      10'h1FC: dout <= 8'b10010000; //  508 : 144 - 0x90
      10'h1FD: dout <= 8'b10010001; //  509 : 145 - 0x91
      10'h1FE: dout <= 8'b10100111; //  510 : 167 - 0xa7
      10'h1FF: dout <= 8'b10100000; //  511 : 160 - 0xa0
      10'h200: dout <= 8'b10100000; //  512 : 160 - 0xa0 -- line 0x10
      10'h201: dout <= 8'b10100011; //  513 : 163 - 0xa3
      10'h202: dout <= 8'b10000010; //  514 : 130 - 0x82
      10'h203: dout <= 8'b10000011; //  515 : 131 - 0x83
      10'h204: dout <= 8'b10000101; //  516 : 133 - 0x85
      10'h205: dout <= 8'b10000110; //  517 : 134 - 0x86
      10'h206: dout <= 8'b10000101; //  518 : 133 - 0x85
      10'h207: dout <= 8'b10000110; //  519 : 134 - 0x86
      10'h208: dout <= 8'b10000101; //  520 : 133 - 0x85
      10'h209: dout <= 8'b10000110; //  521 : 134 - 0x86
      10'h20A: dout <= 8'b10000101; //  522 : 133 - 0x85
      10'h20B: dout <= 8'b10000110; //  523 : 134 - 0x86
      10'h20C: dout <= 8'b10000000; //  524 : 128 - 0x80
      10'h20D: dout <= 8'b10000010; //  525 : 130 - 0x82
      10'h20E: dout <= 8'b10000010; //  526 : 130 - 0x82
      10'h20F: dout <= 8'b10000011; //  527 : 131 - 0x83
      10'h210: dout <= 8'b10000000; //  528 : 128 - 0x80
      10'h211: dout <= 8'b10000001; //  529 : 129 - 0x81
      10'h212: dout <= 8'b10000001; //  530 : 129 - 0x81
      10'h213: dout <= 8'b10000000; //  531 : 128 - 0x80
      10'h214: dout <= 8'b10000101; //  532 : 133 - 0x85
      10'h215: dout <= 8'b10000110; //  533 : 134 - 0x86
      10'h216: dout <= 8'b10000110; //  534 : 134 - 0x86
      10'h217: dout <= 8'b10000111; //  535 : 135 - 0x87
      10'h218: dout <= 8'b10000110; //  536 : 134 - 0x86
      10'h219: dout <= 8'b10000111; //  537 : 135 - 0x87
      10'h21A: dout <= 8'b10000100; //  538 : 132 - 0x84
      10'h21B: dout <= 8'b10000101; //  539 : 133 - 0x85
      10'h21C: dout <= 8'b10000010; //  540 : 130 - 0x82
      10'h21D: dout <= 8'b10000011; //  541 : 131 - 0x83
      10'h21E: dout <= 8'b10100111; //  542 : 167 - 0xa7
      10'h21F: dout <= 8'b10100000; //  543 : 160 - 0xa0
      10'h220: dout <= 8'b10100000; //  544 : 160 - 0xa0 -- line 0x11
      10'h221: dout <= 8'b10100011; //  545 : 163 - 0xa3
      10'h222: dout <= 8'b10010010; //  546 : 146 - 0x92
      10'h223: dout <= 8'b10010011; //  547 : 147 - 0x93
      10'h224: dout <= 8'b10010111; //  548 : 151 - 0x97
      10'h225: dout <= 8'b10010100; //  549 : 148 - 0x94
      10'h226: dout <= 8'b10010111; //  550 : 151 - 0x97
      10'h227: dout <= 8'b10010100; //  551 : 148 - 0x94
      10'h228: dout <= 8'b10010111; //  552 : 151 - 0x97
      10'h229: dout <= 8'b10010100; //  553 : 148 - 0x94
      10'h22A: dout <= 8'b10010111; //  554 : 151 - 0x97
      10'h22B: dout <= 8'b10010100; //  555 : 148 - 0x94
      10'h22C: dout <= 8'b10010010; //  556 : 146 - 0x92
      10'h22D: dout <= 8'b10010001; //  557 : 145 - 0x91
      10'h22E: dout <= 8'b10010010; //  558 : 146 - 0x92
      10'h22F: dout <= 8'b10010011; //  559 : 147 - 0x93
      10'h230: dout <= 8'b10010000; //  560 : 144 - 0x90
      10'h231: dout <= 8'b10010001; //  561 : 145 - 0x91
      10'h232: dout <= 8'b10010011; //  562 : 147 - 0x93
      10'h233: dout <= 8'b10010010; //  563 : 146 - 0x92
      10'h234: dout <= 8'b10010111; //  564 : 151 - 0x97
      10'h235: dout <= 8'b10010100; //  565 : 148 - 0x94
      10'h236: dout <= 8'b10010110; //  566 : 150 - 0x96
      10'h237: dout <= 8'b10010111; //  567 : 151 - 0x97
      10'h238: dout <= 8'b10010110; //  568 : 150 - 0x96
      10'h239: dout <= 8'b10010111; //  569 : 151 - 0x97
      10'h23A: dout <= 8'b10010100; //  570 : 148 - 0x94
      10'h23B: dout <= 8'b10010101; //  571 : 149 - 0x95
      10'h23C: dout <= 8'b10010010; //  572 : 146 - 0x92
      10'h23D: dout <= 8'b10010011; //  573 : 147 - 0x93
      10'h23E: dout <= 8'b10100111; //  574 : 167 - 0xa7
      10'h23F: dout <= 8'b10100000; //  575 : 160 - 0xa0
      10'h240: dout <= 8'b10100000; //  576 : 160 - 0xa0 -- line 0x12
      10'h241: dout <= 8'b10100011; //  577 : 163 - 0xa3
      10'h242: dout <= 8'b10000000; //  578 : 128 - 0x80
      10'h243: dout <= 8'b10000010; //  579 : 130 - 0x82
      10'h244: dout <= 8'b10000100; //  580 : 132 - 0x84
      10'h245: dout <= 8'b10000111; //  581 : 135 - 0x87
      10'h246: dout <= 8'b10000101; //  582 : 133 - 0x85
      10'h247: dout <= 8'b10000110; //  583 : 134 - 0x86
      10'h248: dout <= 8'b10000100; //  584 : 132 - 0x84
      10'h249: dout <= 8'b10000111; //  585 : 135 - 0x87
      10'h24A: dout <= 8'b10000100; //  586 : 132 - 0x84
      10'h24B: dout <= 8'b10000111; //  587 : 135 - 0x87
      10'h24C: dout <= 8'b10000010; //  588 : 130 - 0x82
      10'h24D: dout <= 8'b10000011; //  589 : 131 - 0x83
      10'h24E: dout <= 8'b10000000; //  590 : 128 - 0x80
      10'h24F: dout <= 8'b10000001; //  591 : 129 - 0x81
      10'h250: dout <= 8'b10000000; //  592 : 128 - 0x80
      10'h251: dout <= 8'b10000001; //  593 : 129 - 0x81
      10'h252: dout <= 8'b10000010; //  594 : 130 - 0x82
      10'h253: dout <= 8'b10000011; //  595 : 131 - 0x83
      10'h254: dout <= 8'b10000100; //  596 : 132 - 0x84
      10'h255: dout <= 8'b10000101; //  597 : 133 - 0x85
      10'h256: dout <= 8'b10000101; //  598 : 133 - 0x85
      10'h257: dout <= 8'b10000110; //  599 : 134 - 0x86
      10'h258: dout <= 8'b10000100; //  600 : 132 - 0x84
      10'h259: dout <= 8'b10000111; //  601 : 135 - 0x87
      10'h25A: dout <= 8'b10000100; //  602 : 132 - 0x84
      10'h25B: dout <= 8'b10000111; //  603 : 135 - 0x87
      10'h25C: dout <= 8'b10000000; //  604 : 128 - 0x80
      10'h25D: dout <= 8'b10000001; //  605 : 129 - 0x81
      10'h25E: dout <= 8'b10100111; //  606 : 167 - 0xa7
      10'h25F: dout <= 8'b10100000; //  607 : 160 - 0xa0
      10'h260: dout <= 8'b10100000; //  608 : 160 - 0xa0 -- line 0x13
      10'h261: dout <= 8'b10100011; //  609 : 163 - 0xa3
      10'h262: dout <= 8'b10010010; //  610 : 146 - 0x92
      10'h263: dout <= 8'b10010001; //  611 : 145 - 0x91
      10'h264: dout <= 8'b10010110; //  612 : 150 - 0x96
      10'h265: dout <= 8'b10010101; //  613 : 149 - 0x95
      10'h266: dout <= 8'b10010111; //  614 : 151 - 0x97
      10'h267: dout <= 8'b10010100; //  615 : 148 - 0x94
      10'h268: dout <= 8'b10010110; //  616 : 150 - 0x96
      10'h269: dout <= 8'b10010101; //  617 : 149 - 0x95
      10'h26A: dout <= 8'b10010110; //  618 : 150 - 0x96
      10'h26B: dout <= 8'b10010101; //  619 : 149 - 0x95
      10'h26C: dout <= 8'b10010010; //  620 : 146 - 0x92
      10'h26D: dout <= 8'b10010011; //  621 : 147 - 0x93
      10'h26E: dout <= 8'b10010000; //  622 : 144 - 0x90
      10'h26F: dout <= 8'b10010001; //  623 : 145 - 0x91
      10'h270: dout <= 8'b10010000; //  624 : 144 - 0x90
      10'h271: dout <= 8'b10010001; //  625 : 145 - 0x91
      10'h272: dout <= 8'b10010010; //  626 : 146 - 0x92
      10'h273: dout <= 8'b10010011; //  627 : 147 - 0x93
      10'h274: dout <= 8'b10010100; //  628 : 148 - 0x94
      10'h275: dout <= 8'b10010101; //  629 : 149 - 0x95
      10'h276: dout <= 8'b10010111; //  630 : 151 - 0x97
      10'h277: dout <= 8'b10010100; //  631 : 148 - 0x94
      10'h278: dout <= 8'b10010110; //  632 : 150 - 0x96
      10'h279: dout <= 8'b10010101; //  633 : 149 - 0x95
      10'h27A: dout <= 8'b10010110; //  634 : 150 - 0x96
      10'h27B: dout <= 8'b10010101; //  635 : 149 - 0x95
      10'h27C: dout <= 8'b10010000; //  636 : 144 - 0x90
      10'h27D: dout <= 8'b10010001; //  637 : 145 - 0x91
      10'h27E: dout <= 8'b10100111; //  638 : 167 - 0xa7
      10'h27F: dout <= 8'b10100000; //  639 : 160 - 0xa0
      10'h280: dout <= 8'b10100000; //  640 : 160 - 0xa0 -- line 0x14
      10'h281: dout <= 8'b10100011; //  641 : 163 - 0xa3
      10'h282: dout <= 8'b10000010; //  642 : 130 - 0x82
      10'h283: dout <= 8'b10000011; //  643 : 131 - 0x83
      10'h284: dout <= 8'b10000110; //  644 : 134 - 0x86
      10'h285: dout <= 8'b10000111; //  645 : 135 - 0x87
      10'h286: dout <= 8'b10000100; //  646 : 132 - 0x84
      10'h287: dout <= 8'b10000101; //  647 : 133 - 0x85
      10'h288: dout <= 8'b10000100; //  648 : 132 - 0x84
      10'h289: dout <= 8'b10000111; //  649 : 135 - 0x87
      10'h28A: dout <= 8'b10000100; //  650 : 132 - 0x84
      10'h28B: dout <= 8'b10000111; //  651 : 135 - 0x87
      10'h28C: dout <= 8'b10000110; //  652 : 134 - 0x86
      10'h28D: dout <= 8'b10000111; //  653 : 135 - 0x87
      10'h28E: dout <= 8'b10000100; //  654 : 132 - 0x84
      10'h28F: dout <= 8'b10000111; //  655 : 135 - 0x87
      10'h290: dout <= 8'b10000110; //  656 : 134 - 0x86
      10'h291: dout <= 8'b10000111; //  657 : 135 - 0x87
      10'h292: dout <= 8'b10000110; //  658 : 134 - 0x86
      10'h293: dout <= 8'b10000111; //  659 : 135 - 0x87
      10'h294: dout <= 8'b10000110; //  660 : 134 - 0x86
      10'h295: dout <= 8'b10000111; //  661 : 135 - 0x87
      10'h296: dout <= 8'b10000110; //  662 : 134 - 0x86
      10'h297: dout <= 8'b10000111; //  663 : 135 - 0x87
      10'h298: dout <= 8'b10000101; //  664 : 133 - 0x85
      10'h299: dout <= 8'b10000110; //  665 : 134 - 0x86
      10'h29A: dout <= 8'b10000100; //  666 : 132 - 0x84
      10'h29B: dout <= 8'b10000111; //  667 : 135 - 0x87
      10'h29C: dout <= 8'b10000000; //  668 : 128 - 0x80
      10'h29D: dout <= 8'b10000010; //  669 : 130 - 0x82
      10'h29E: dout <= 8'b10100111; //  670 : 167 - 0xa7
      10'h29F: dout <= 8'b10100000; //  671 : 160 - 0xa0
      10'h2A0: dout <= 8'b10100000; //  672 : 160 - 0xa0 -- line 0x15
      10'h2A1: dout <= 8'b10100011; //  673 : 163 - 0xa3
      10'h2A2: dout <= 8'b10010010; //  674 : 146 - 0x92
      10'h2A3: dout <= 8'b10010011; //  675 : 147 - 0x93
      10'h2A4: dout <= 8'b10010110; //  676 : 150 - 0x96
      10'h2A5: dout <= 8'b10010111; //  677 : 151 - 0x97
      10'h2A6: dout <= 8'b10010100; //  678 : 148 - 0x94
      10'h2A7: dout <= 8'b10010101; //  679 : 149 - 0x95
      10'h2A8: dout <= 8'b10010110; //  680 : 150 - 0x96
      10'h2A9: dout <= 8'b10010101; //  681 : 149 - 0x95
      10'h2AA: dout <= 8'b10010110; //  682 : 150 - 0x96
      10'h2AB: dout <= 8'b10010101; //  683 : 149 - 0x95
      10'h2AC: dout <= 8'b10010110; //  684 : 150 - 0x96
      10'h2AD: dout <= 8'b10010111; //  685 : 151 - 0x97
      10'h2AE: dout <= 8'b10010110; //  686 : 150 - 0x96
      10'h2AF: dout <= 8'b10010101; //  687 : 149 - 0x95
      10'h2B0: dout <= 8'b10010110; //  688 : 150 - 0x96
      10'h2B1: dout <= 8'b10010111; //  689 : 151 - 0x97
      10'h2B2: dout <= 8'b10010110; //  690 : 150 - 0x96
      10'h2B3: dout <= 8'b10010111; //  691 : 151 - 0x97
      10'h2B4: dout <= 8'b10010110; //  692 : 150 - 0x96
      10'h2B5: dout <= 8'b10010111; //  693 : 151 - 0x97
      10'h2B6: dout <= 8'b10010110; //  694 : 150 - 0x96
      10'h2B7: dout <= 8'b10010111; //  695 : 151 - 0x97
      10'h2B8: dout <= 8'b10010111; //  696 : 151 - 0x97
      10'h2B9: dout <= 8'b10010100; //  697 : 148 - 0x94
      10'h2BA: dout <= 8'b10010110; //  698 : 150 - 0x96
      10'h2BB: dout <= 8'b10010101; //  699 : 149 - 0x95
      10'h2BC: dout <= 8'b10010010; //  700 : 146 - 0x92
      10'h2BD: dout <= 8'b10010001; //  701 : 145 - 0x91
      10'h2BE: dout <= 8'b10100111; //  702 : 167 - 0xa7
      10'h2BF: dout <= 8'b10100000; //  703 : 160 - 0xa0
      10'h2C0: dout <= 8'b10100000; //  704 : 160 - 0xa0 -- line 0x16
      10'h2C1: dout <= 8'b10100011; //  705 : 163 - 0xa3
      10'h2C2: dout <= 8'b10000000; //  706 : 128 - 0x80
      10'h2C3: dout <= 8'b10000001; //  707 : 129 - 0x81
      10'h2C4: dout <= 8'b10000101; //  708 : 133 - 0x85
      10'h2C5: dout <= 8'b10000110; //  709 : 134 - 0x86
      10'h2C6: dout <= 8'b10000100; //  710 : 132 - 0x84
      10'h2C7: dout <= 8'b10000101; //  711 : 133 - 0x85
      10'h2C8: dout <= 8'b10000100; //  712 : 132 - 0x84
      10'h2C9: dout <= 8'b10000101; //  713 : 133 - 0x85
      10'h2CA: dout <= 8'b10000100; //  714 : 132 - 0x84
      10'h2CB: dout <= 8'b10000111; //  715 : 135 - 0x87
      10'h2CC: dout <= 8'b10000101; //  716 : 133 - 0x85
      10'h2CD: dout <= 8'b10000110; //  717 : 134 - 0x86
      10'h2CE: dout <= 8'b10000110; //  718 : 134 - 0x86
      10'h2CF: dout <= 8'b10000111; //  719 : 135 - 0x87
      10'h2D0: dout <= 8'b10000110; //  720 : 134 - 0x86
      10'h2D1: dout <= 8'b10000111; //  721 : 135 - 0x87
      10'h2D2: dout <= 8'b10000101; //  722 : 133 - 0x85
      10'h2D3: dout <= 8'b10000110; //  723 : 134 - 0x86
      10'h2D4: dout <= 8'b10000101; //  724 : 133 - 0x85
      10'h2D5: dout <= 8'b10000110; //  725 : 134 - 0x86
      10'h2D6: dout <= 8'b10000110; //  726 : 134 - 0x86
      10'h2D7: dout <= 8'b10000111; //  727 : 135 - 0x87
      10'h2D8: dout <= 8'b10000100; //  728 : 132 - 0x84
      10'h2D9: dout <= 8'b10000111; //  729 : 135 - 0x87
      10'h2DA: dout <= 8'b10000100; //  730 : 132 - 0x84
      10'h2DB: dout <= 8'b10000111; //  731 : 135 - 0x87
      10'h2DC: dout <= 8'b10000000; //  732 : 128 - 0x80
      10'h2DD: dout <= 8'b10000001; //  733 : 129 - 0x81
      10'h2DE: dout <= 8'b10100111; //  734 : 167 - 0xa7
      10'h2DF: dout <= 8'b10100000; //  735 : 160 - 0xa0
      10'h2E0: dout <= 8'b10100000; //  736 : 160 - 0xa0 -- line 0x17
      10'h2E1: dout <= 8'b10100011; //  737 : 163 - 0xa3
      10'h2E2: dout <= 8'b10010000; //  738 : 144 - 0x90
      10'h2E3: dout <= 8'b10010001; //  739 : 145 - 0x91
      10'h2E4: dout <= 8'b10010111; //  740 : 151 - 0x97
      10'h2E5: dout <= 8'b10010100; //  741 : 148 - 0x94
      10'h2E6: dout <= 8'b10010100; //  742 : 148 - 0x94
      10'h2E7: dout <= 8'b10010101; //  743 : 149 - 0x95
      10'h2E8: dout <= 8'b10010100; //  744 : 148 - 0x94
      10'h2E9: dout <= 8'b10010101; //  745 : 149 - 0x95
      10'h2EA: dout <= 8'b10010110; //  746 : 150 - 0x96
      10'h2EB: dout <= 8'b10010101; //  747 : 149 - 0x95
      10'h2EC: dout <= 8'b10010111; //  748 : 151 - 0x97
      10'h2ED: dout <= 8'b10010100; //  749 : 148 - 0x94
      10'h2EE: dout <= 8'b10010110; //  750 : 150 - 0x96
      10'h2EF: dout <= 8'b10010111; //  751 : 151 - 0x97
      10'h2F0: dout <= 8'b10010110; //  752 : 150 - 0x96
      10'h2F1: dout <= 8'b10010111; //  753 : 151 - 0x97
      10'h2F2: dout <= 8'b10010111; //  754 : 151 - 0x97
      10'h2F3: dout <= 8'b10010100; //  755 : 148 - 0x94
      10'h2F4: dout <= 8'b10010111; //  756 : 151 - 0x97
      10'h2F5: dout <= 8'b10010100; //  757 : 148 - 0x94
      10'h2F6: dout <= 8'b10010110; //  758 : 150 - 0x96
      10'h2F7: dout <= 8'b10010111; //  759 : 151 - 0x97
      10'h2F8: dout <= 8'b10010110; //  760 : 150 - 0x96
      10'h2F9: dout <= 8'b10010101; //  761 : 149 - 0x95
      10'h2FA: dout <= 8'b10010110; //  762 : 150 - 0x96
      10'h2FB: dout <= 8'b10010101; //  763 : 149 - 0x95
      10'h2FC: dout <= 8'b10010000; //  764 : 144 - 0x90
      10'h2FD: dout <= 8'b10010001; //  765 : 145 - 0x91
      10'h2FE: dout <= 8'b10100111; //  766 : 167 - 0xa7
      10'h2FF: dout <= 8'b10100000; //  767 : 160 - 0xa0
      10'h300: dout <= 8'b10100000; //  768 : 160 - 0xa0 -- line 0x18
      10'h301: dout <= 8'b10100011; //  769 : 163 - 0xa3
      10'h302: dout <= 8'b10000000; //  770 : 128 - 0x80
      10'h303: dout <= 8'b10000010; //  771 : 130 - 0x82
      10'h304: dout <= 8'b10000100; //  772 : 132 - 0x84
      10'h305: dout <= 8'b10000111; //  773 : 135 - 0x87
      10'h306: dout <= 8'b10000100; //  774 : 132 - 0x84
      10'h307: dout <= 8'b10000111; //  775 : 135 - 0x87
      10'h308: dout <= 8'b10000100; //  776 : 132 - 0x84
      10'h309: dout <= 8'b10000111; //  777 : 135 - 0x87
      10'h30A: dout <= 8'b10000110; //  778 : 134 - 0x86
      10'h30B: dout <= 8'b10000111; //  779 : 135 - 0x87
      10'h30C: dout <= 8'b10000101; //  780 : 133 - 0x85
      10'h30D: dout <= 8'b10000110; //  781 : 134 - 0x86
      10'h30E: dout <= 8'b10000100; //  782 : 132 - 0x84
      10'h30F: dout <= 8'b10000111; //  783 : 135 - 0x87
      10'h310: dout <= 8'b10000100; //  784 : 132 - 0x84
      10'h311: dout <= 8'b10000101; //  785 : 133 - 0x85
      10'h312: dout <= 8'b10000100; //  786 : 132 - 0x84
      10'h313: dout <= 8'b10000111; //  787 : 135 - 0x87
      10'h314: dout <= 8'b10000110; //  788 : 134 - 0x86
      10'h315: dout <= 8'b10000111; //  789 : 135 - 0x87
      10'h316: dout <= 8'b10000110; //  790 : 134 - 0x86
      10'h317: dout <= 8'b10000111; //  791 : 135 - 0x87
      10'h318: dout <= 8'b10000100; //  792 : 132 - 0x84
      10'h319: dout <= 8'b10000111; //  793 : 135 - 0x87
      10'h31A: dout <= 8'b10000101; //  794 : 133 - 0x85
      10'h31B: dout <= 8'b10000110; //  795 : 134 - 0x86
      10'h31C: dout <= 8'b10000000; //  796 : 128 - 0x80
      10'h31D: dout <= 8'b10000010; //  797 : 130 - 0x82
      10'h31E: dout <= 8'b10100111; //  798 : 167 - 0xa7
      10'h31F: dout <= 8'b10100000; //  799 : 160 - 0xa0
      10'h320: dout <= 8'b10100000; //  800 : 160 - 0xa0 -- line 0x19
      10'h321: dout <= 8'b10100011; //  801 : 163 - 0xa3
      10'h322: dout <= 8'b10010010; //  802 : 146 - 0x92
      10'h323: dout <= 8'b10010001; //  803 : 145 - 0x91
      10'h324: dout <= 8'b10010110; //  804 : 150 - 0x96
      10'h325: dout <= 8'b10010101; //  805 : 149 - 0x95
      10'h326: dout <= 8'b10010110; //  806 : 150 - 0x96
      10'h327: dout <= 8'b10010101; //  807 : 149 - 0x95
      10'h328: dout <= 8'b10010110; //  808 : 150 - 0x96
      10'h329: dout <= 8'b10010101; //  809 : 149 - 0x95
      10'h32A: dout <= 8'b10010110; //  810 : 150 - 0x96
      10'h32B: dout <= 8'b10010111; //  811 : 151 - 0x97
      10'h32C: dout <= 8'b10010111; //  812 : 151 - 0x97
      10'h32D: dout <= 8'b10010100; //  813 : 148 - 0x94
      10'h32E: dout <= 8'b10010110; //  814 : 150 - 0x96
      10'h32F: dout <= 8'b10010101; //  815 : 149 - 0x95
      10'h330: dout <= 8'b10010100; //  816 : 148 - 0x94
      10'h331: dout <= 8'b10010101; //  817 : 149 - 0x95
      10'h332: dout <= 8'b10010110; //  818 : 150 - 0x96
      10'h333: dout <= 8'b10010101; //  819 : 149 - 0x95
      10'h334: dout <= 8'b10010110; //  820 : 150 - 0x96
      10'h335: dout <= 8'b10010111; //  821 : 151 - 0x97
      10'h336: dout <= 8'b10010110; //  822 : 150 - 0x96
      10'h337: dout <= 8'b10010111; //  823 : 151 - 0x97
      10'h338: dout <= 8'b10010110; //  824 : 150 - 0x96
      10'h339: dout <= 8'b10010101; //  825 : 149 - 0x95
      10'h33A: dout <= 8'b10010111; //  826 : 151 - 0x97
      10'h33B: dout <= 8'b10010100; //  827 : 148 - 0x94
      10'h33C: dout <= 8'b10010010; //  828 : 146 - 0x92
      10'h33D: dout <= 8'b10010001; //  829 : 145 - 0x91
      10'h33E: dout <= 8'b10100111; //  830 : 167 - 0xa7
      10'h33F: dout <= 8'b10100000; //  831 : 160 - 0xa0
      10'h340: dout <= 8'b10100000; //  832 : 160 - 0xa0 -- line 0x1a
      10'h341: dout <= 8'b10100011; //  833 : 163 - 0xa3
      10'h342: dout <= 8'b10000001; //  834 : 129 - 0x81
      10'h343: dout <= 8'b10000000; //  835 : 128 - 0x80
      10'h344: dout <= 8'b10000000; //  836 : 128 - 0x80
      10'h345: dout <= 8'b10000001; //  837 : 129 - 0x81
      10'h346: dout <= 8'b10000010; //  838 : 130 - 0x82
      10'h347: dout <= 8'b10000011; //  839 : 131 - 0x83
      10'h348: dout <= 8'b10000001; //  840 : 129 - 0x81
      10'h349: dout <= 8'b10000000; //  841 : 128 - 0x80
      10'h34A: dout <= 8'b10000001; //  842 : 129 - 0x81
      10'h34B: dout <= 8'b10000000; //  843 : 128 - 0x80
      10'h34C: dout <= 8'b10000000; //  844 : 128 - 0x80
      10'h34D: dout <= 8'b10000010; //  845 : 130 - 0x82
      10'h34E: dout <= 8'b10000000; //  846 : 128 - 0x80
      10'h34F: dout <= 8'b10000001; //  847 : 129 - 0x81
      10'h350: dout <= 8'b10000001; //  848 : 129 - 0x81
      10'h351: dout <= 8'b10000000; //  849 : 128 - 0x80
      10'h352: dout <= 8'b10000000; //  850 : 128 - 0x80
      10'h353: dout <= 8'b10000010; //  851 : 130 - 0x82
      10'h354: dout <= 8'b10000000; //  852 : 128 - 0x80
      10'h355: dout <= 8'b10000001; //  853 : 129 - 0x81
      10'h356: dout <= 8'b10000010; //  854 : 130 - 0x82
      10'h357: dout <= 8'b10000011; //  855 : 131 - 0x83
      10'h358: dout <= 8'b10000001; //  856 : 129 - 0x81
      10'h359: dout <= 8'b10000000; //  857 : 128 - 0x80
      10'h35A: dout <= 8'b10000000; //  858 : 128 - 0x80
      10'h35B: dout <= 8'b10000001; //  859 : 129 - 0x81
      10'h35C: dout <= 8'b10000000; //  860 : 128 - 0x80
      10'h35D: dout <= 8'b10000001; //  861 : 129 - 0x81
      10'h35E: dout <= 8'b10100111; //  862 : 167 - 0xa7
      10'h35F: dout <= 8'b10100000; //  863 : 160 - 0xa0
      10'h360: dout <= 8'b10100000; //  864 : 160 - 0xa0 -- line 0x1b
      10'h361: dout <= 8'b10100011; //  865 : 163 - 0xa3
      10'h362: dout <= 8'b10010011; //  866 : 147 - 0x93
      10'h363: dout <= 8'b10010010; //  867 : 146 - 0x92
      10'h364: dout <= 8'b10010000; //  868 : 144 - 0x90
      10'h365: dout <= 8'b10010001; //  869 : 145 - 0x91
      10'h366: dout <= 8'b10010010; //  870 : 146 - 0x92
      10'h367: dout <= 8'b10010011; //  871 : 147 - 0x93
      10'h368: dout <= 8'b10010011; //  872 : 147 - 0x93
      10'h369: dout <= 8'b10010010; //  873 : 146 - 0x92
      10'h36A: dout <= 8'b10010011; //  874 : 147 - 0x93
      10'h36B: dout <= 8'b10010010; //  875 : 146 - 0x92
      10'h36C: dout <= 8'b10010010; //  876 : 146 - 0x92
      10'h36D: dout <= 8'b10010001; //  877 : 145 - 0x91
      10'h36E: dout <= 8'b10010000; //  878 : 144 - 0x90
      10'h36F: dout <= 8'b10010001; //  879 : 145 - 0x91
      10'h370: dout <= 8'b10010011; //  880 : 147 - 0x93
      10'h371: dout <= 8'b10010010; //  881 : 146 - 0x92
      10'h372: dout <= 8'b10010010; //  882 : 146 - 0x92
      10'h373: dout <= 8'b10010001; //  883 : 145 - 0x91
      10'h374: dout <= 8'b10010000; //  884 : 144 - 0x90
      10'h375: dout <= 8'b10010001; //  885 : 145 - 0x91
      10'h376: dout <= 8'b10010010; //  886 : 146 - 0x92
      10'h377: dout <= 8'b10010011; //  887 : 147 - 0x93
      10'h378: dout <= 8'b10010011; //  888 : 147 - 0x93
      10'h379: dout <= 8'b10010010; //  889 : 146 - 0x92
      10'h37A: dout <= 8'b10010000; //  890 : 144 - 0x90
      10'h37B: dout <= 8'b10010001; //  891 : 145 - 0x91
      10'h37C: dout <= 8'b10010000; //  892 : 144 - 0x90
      10'h37D: dout <= 8'b10010001; //  893 : 145 - 0x91
      10'h37E: dout <= 8'b10100111; //  894 : 167 - 0xa7
      10'h37F: dout <= 8'b10100000; //  895 : 160 - 0xa0
      10'h380: dout <= 8'b10100000; //  896 : 160 - 0xa0 -- line 0x1c
      10'h381: dout <= 8'b10100100; //  897 : 164 - 0xa4
      10'h382: dout <= 8'b10100101; //  898 : 165 - 0xa5
      10'h383: dout <= 8'b10100101; //  899 : 165 - 0xa5
      10'h384: dout <= 8'b10100101; //  900 : 165 - 0xa5
      10'h385: dout <= 8'b10100101; //  901 : 165 - 0xa5
      10'h386: dout <= 8'b10100101; //  902 : 165 - 0xa5
      10'h387: dout <= 8'b10100101; //  903 : 165 - 0xa5
      10'h388: dout <= 8'b10100101; //  904 : 165 - 0xa5
      10'h389: dout <= 8'b10100101; //  905 : 165 - 0xa5
      10'h38A: dout <= 8'b10100101; //  906 : 165 - 0xa5
      10'h38B: dout <= 8'b10100101; //  907 : 165 - 0xa5
      10'h38C: dout <= 8'b10100101; //  908 : 165 - 0xa5
      10'h38D: dout <= 8'b10100101; //  909 : 165 - 0xa5
      10'h38E: dout <= 8'b10100101; //  910 : 165 - 0xa5
      10'h38F: dout <= 8'b10100101; //  911 : 165 - 0xa5
      10'h390: dout <= 8'b10100101; //  912 : 165 - 0xa5
      10'h391: dout <= 8'b10100101; //  913 : 165 - 0xa5
      10'h392: dout <= 8'b10100101; //  914 : 165 - 0xa5
      10'h393: dout <= 8'b10100101; //  915 : 165 - 0xa5
      10'h394: dout <= 8'b10100101; //  916 : 165 - 0xa5
      10'h395: dout <= 8'b10100101; //  917 : 165 - 0xa5
      10'h396: dout <= 8'b10100101; //  918 : 165 - 0xa5
      10'h397: dout <= 8'b10100101; //  919 : 165 - 0xa5
      10'h398: dout <= 8'b10100101; //  920 : 165 - 0xa5
      10'h399: dout <= 8'b10100101; //  921 : 165 - 0xa5
      10'h39A: dout <= 8'b10100101; //  922 : 165 - 0xa5
      10'h39B: dout <= 8'b10100101; //  923 : 165 - 0xa5
      10'h39C: dout <= 8'b10100101; //  924 : 165 - 0xa5
      10'h39D: dout <= 8'b10100101; //  925 : 165 - 0xa5
      10'h39E: dout <= 8'b10101000; //  926 : 168 - 0xa8
      10'h39F: dout <= 8'b10100000; //  927 : 160 - 0xa0
      10'h3A0: dout <= 8'b10100000; //  928 : 160 - 0xa0 -- line 0x1d
      10'h3A1: dout <= 8'b10100000; //  929 : 160 - 0xa0
      10'h3A2: dout <= 8'b10100000; //  930 : 160 - 0xa0
      10'h3A3: dout <= 8'b10100000; //  931 : 160 - 0xa0
      10'h3A4: dout <= 8'b10100000; //  932 : 160 - 0xa0
      10'h3A5: dout <= 8'b10100000; //  933 : 160 - 0xa0
      10'h3A6: dout <= 8'b10100000; //  934 : 160 - 0xa0
      10'h3A7: dout <= 8'b10100000; //  935 : 160 - 0xa0
      10'h3A8: dout <= 8'b10100000; //  936 : 160 - 0xa0
      10'h3A9: dout <= 8'b10100000; //  937 : 160 - 0xa0
      10'h3AA: dout <= 8'b10100000; //  938 : 160 - 0xa0
      10'h3AB: dout <= 8'b10100000; //  939 : 160 - 0xa0
      10'h3AC: dout <= 8'b10100000; //  940 : 160 - 0xa0
      10'h3AD: dout <= 8'b10100000; //  941 : 160 - 0xa0
      10'h3AE: dout <= 8'b10100000; //  942 : 160 - 0xa0
      10'h3AF: dout <= 8'b10100000; //  943 : 160 - 0xa0
      10'h3B0: dout <= 8'b10100000; //  944 : 160 - 0xa0
      10'h3B1: dout <= 8'b10100000; //  945 : 160 - 0xa0
      10'h3B2: dout <= 8'b10100000; //  946 : 160 - 0xa0
      10'h3B3: dout <= 8'b10100000; //  947 : 160 - 0xa0
      10'h3B4: dout <= 8'b10100000; //  948 : 160 - 0xa0
      10'h3B5: dout <= 8'b10100000; //  949 : 160 - 0xa0
      10'h3B6: dout <= 8'b10100000; //  950 : 160 - 0xa0
      10'h3B7: dout <= 8'b10100000; //  951 : 160 - 0xa0
      10'h3B8: dout <= 8'b10100000; //  952 : 160 - 0xa0
      10'h3B9: dout <= 8'b10100000; //  953 : 160 - 0xa0
      10'h3BA: dout <= 8'b10100000; //  954 : 160 - 0xa0
      10'h3BB: dout <= 8'b10100000; //  955 : 160 - 0xa0
      10'h3BC: dout <= 8'b10100000; //  956 : 160 - 0xa0
      10'h3BD: dout <= 8'b10100000; //  957 : 160 - 0xa0
      10'h3BE: dout <= 8'b10100000; //  958 : 160 - 0xa0
      10'h3BF: dout <= 8'b10100000; //  959 : 160 - 0xa0
        //-- Attribute Table 0----
      10'h3C0: dout <= 8'b00000000; //  960 :   0 - 0x0
      10'h3C1: dout <= 8'b00000000; //  961 :   0 - 0x0
      10'h3C2: dout <= 8'b00000000; //  962 :   0 - 0x0
      10'h3C3: dout <= 8'b00000000; //  963 :   0 - 0x0
      10'h3C4: dout <= 8'b00000000; //  964 :   0 - 0x0
      10'h3C5: dout <= 8'b00000000; //  965 :   0 - 0x0
      10'h3C6: dout <= 8'b00000000; //  966 :   0 - 0x0
      10'h3C7: dout <= 8'b00000000; //  967 :   0 - 0x0
      10'h3C8: dout <= 8'b10000000; //  968 : 128 - 0x80
      10'h3C9: dout <= 8'b10100000; //  969 : 160 - 0xa0
      10'h3CA: dout <= 8'b10100000; //  970 : 160 - 0xa0
      10'h3CB: dout <= 8'b10100000; //  971 : 160 - 0xa0
      10'h3CC: dout <= 8'b10100000; //  972 : 160 - 0xa0
      10'h3CD: dout <= 8'b10100000; //  973 : 160 - 0xa0
      10'h3CE: dout <= 8'b10100000; //  974 : 160 - 0xa0
      10'h3CF: dout <= 8'b00100000; //  975 :  32 - 0x20
      10'h3D0: dout <= 8'b10001000; //  976 : 136 - 0x88
      10'h3D1: dout <= 8'b10101010; //  977 : 170 - 0xaa
      10'h3D2: dout <= 8'b10101010; //  978 : 170 - 0xaa
      10'h3D3: dout <= 8'b10101010; //  979 : 170 - 0xaa
      10'h3D4: dout <= 8'b10101010; //  980 : 170 - 0xaa
      10'h3D5: dout <= 8'b10101010; //  981 : 170 - 0xaa
      10'h3D6: dout <= 8'b10101010; //  982 : 170 - 0xaa
      10'h3D7: dout <= 8'b00100010; //  983 :  34 - 0x22
      10'h3D8: dout <= 8'b10001000; //  984 : 136 - 0x88
      10'h3D9: dout <= 8'b10101010; //  985 : 170 - 0xaa
      10'h3DA: dout <= 8'b10101010; //  986 : 170 - 0xaa
      10'h3DB: dout <= 8'b10101010; //  987 : 170 - 0xaa
      10'h3DC: dout <= 8'b10101010; //  988 : 170 - 0xaa
      10'h3DD: dout <= 8'b10101010; //  989 : 170 - 0xaa
      10'h3DE: dout <= 8'b10101010; //  990 : 170 - 0xaa
      10'h3DF: dout <= 8'b00100010; //  991 :  34 - 0x22
      10'h3E0: dout <= 8'b10001000; //  992 : 136 - 0x88
      10'h3E1: dout <= 8'b10101010; //  993 : 170 - 0xaa
      10'h3E2: dout <= 8'b10101010; //  994 : 170 - 0xaa
      10'h3E3: dout <= 8'b10101010; //  995 : 170 - 0xaa
      10'h3E4: dout <= 8'b10101010; //  996 : 170 - 0xaa
      10'h3E5: dout <= 8'b10101010; //  997 : 170 - 0xaa
      10'h3E6: dout <= 8'b10101010; //  998 : 170 - 0xaa
      10'h3E7: dout <= 8'b00100010; //  999 :  34 - 0x22
      10'h3E8: dout <= 8'b10001000; // 1000 : 136 - 0x88
      10'h3E9: dout <= 8'b10101010; // 1001 : 170 - 0xaa
      10'h3EA: dout <= 8'b10101010; // 1002 : 170 - 0xaa
      10'h3EB: dout <= 8'b10101010; // 1003 : 170 - 0xaa
      10'h3EC: dout <= 8'b10101010; // 1004 : 170 - 0xaa
      10'h3ED: dout <= 8'b10101010; // 1005 : 170 - 0xaa
      10'h3EE: dout <= 8'b10101010; // 1006 : 170 - 0xaa
      10'h3EF: dout <= 8'b00100010; // 1007 :  34 - 0x22
      10'h3F0: dout <= 8'b10001000; // 1008 : 136 - 0x88
      10'h3F1: dout <= 8'b10101010; // 1009 : 170 - 0xaa
      10'h3F2: dout <= 8'b10101010; // 1010 : 170 - 0xaa
      10'h3F3: dout <= 8'b10101010; // 1011 : 170 - 0xaa
      10'h3F4: dout <= 8'b10101010; // 1012 : 170 - 0xaa
      10'h3F5: dout <= 8'b10101010; // 1013 : 170 - 0xaa
      10'h3F6: dout <= 8'b10101010; // 1014 : 170 - 0xaa
      10'h3F7: dout <= 8'b00100010; // 1015 :  34 - 0x22
      10'h3F8: dout <= 8'b00000000; // 1016 :   0 - 0x0
      10'h3F9: dout <= 8'b00000000; // 1017 :   0 - 0x0
      10'h3FA: dout <= 8'b00000000; // 1018 :   0 - 0x0
      10'h3FB: dout <= 8'b00000000; // 1019 :   0 - 0x0
      10'h3FC: dout <= 8'b00000000; // 1020 :   0 - 0x0
      10'h3FD: dout <= 8'b00000000; // 1021 :   0 - 0x0
      10'h3FE: dout <= 8'b00000000; // 1022 :   0 - 0x0
      10'h3FF: dout <= 8'b00000000; // 1023 :   0 - 0x0
    endcase
  end

endmodule
