--- Autcmatically generated VHDL ROM from a NES memory file----
---   ATTRIBUTE TABLE SEPARATED FROM NAME TABLE
-- https://wiki.nesdev.com/w/index.php/PPU_attribute_tables


---  Original memory dump file name: lawnmower_ntable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory with clock ------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_ATABLE_LAWN_00 is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(7-1 downto 0);  --128 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_ATABLE_LAWN_00;

architecture BEHAVIORAL of ROM_ATABLE_LAWN_00 is
  signal addr_int  : natural range 0 to 2**7-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
    "00000000", --    0 -  0x0  :    0 - 0x0
    "00000000", --    1 -  0x1  :    0 - 0x0
    "00000000", --    2 -  0x2  :    0 - 0x0
    "00000000", --    3 -  0x3  :    0 - 0x0
    "00000000", --    4 -  0x4  :    0 - 0x0
    "00000000", --    5 -  0x5  :    0 - 0x0
    "00000000", --    6 -  0x6  :    0 - 0x0
    "00000000", --    7 -  0x7  :    0 - 0x0
    "10000000", --    8 -  0x8  :  128 - 0x80
    "10100000", --    9 -  0x9  :  160 - 0xa0
    "10100000", --   10 -  0xa  :  160 - 0xa0
    "10100000", --   11 -  0xb  :  160 - 0xa0
    "10100000", --   12 -  0xc  :  160 - 0xa0
    "10100000", --   13 -  0xd  :  160 - 0xa0
    "10100000", --   14 -  0xe  :  160 - 0xa0
    "00100000", --   15 -  0xf  :   32 - 0x20
    "10001000", --   16 - 0x10  :  136 - 0x88
    "10101010", --   17 - 0x11  :  170 - 0xaa
    "10101010", --   18 - 0x12  :  170 - 0xaa
    "10101010", --   19 - 0x13  :  170 - 0xaa
    "10101010", --   20 - 0x14  :  170 - 0xaa
    "10101010", --   21 - 0x15  :  170 - 0xaa
    "10101010", --   22 - 0x16  :  170 - 0xaa
    "00100010", --   23 - 0x17  :   34 - 0x22
    "10001000", --   24 - 0x18  :  136 - 0x88
    "10101010", --   25 - 0x19  :  170 - 0xaa
    "10101010", --   26 - 0x1a  :  170 - 0xaa
    "10101010", --   27 - 0x1b  :  170 - 0xaa
    "10101010", --   28 - 0x1c  :  170 - 0xaa
    "10101010", --   29 - 0x1d  :  170 - 0xaa
    "10101010", --   30 - 0x1e  :  170 - 0xaa
    "00100010", --   31 - 0x1f  :   34 - 0x22
    "10001000", --   32 - 0x20  :  136 - 0x88
    "10101010", --   33 - 0x21  :  170 - 0xaa
    "10101010", --   34 - 0x22  :  170 - 0xaa
    "10101010", --   35 - 0x23  :  170 - 0xaa
    "10101010", --   36 - 0x24  :  170 - 0xaa
    "10101010", --   37 - 0x25  :  170 - 0xaa
    "10101010", --   38 - 0x26  :  170 - 0xaa
    "00100010", --   39 - 0x27  :   34 - 0x22
    "10001000", --   40 - 0x28  :  136 - 0x88
    "10101010", --   41 - 0x29  :  170 - 0xaa
    "10101010", --   42 - 0x2a  :  170 - 0xaa
    "10101010", --   43 - 0x2b  :  170 - 0xaa
    "10101010", --   44 - 0x2c  :  170 - 0xaa
    "10101010", --   45 - 0x2d  :  170 - 0xaa
    "10101010", --   46 - 0x2e  :  170 - 0xaa
    "00100010", --   47 - 0x2f  :   34 - 0x22
    "10001000", --   48 - 0x30  :  136 - 0x88
    "10101010", --   49 - 0x31  :  170 - 0xaa
    "10101010", --   50 - 0x32  :  170 - 0xaa
    "10101010", --   51 - 0x33  :  170 - 0xaa
    "10101010", --   52 - 0x34  :  170 - 0xaa
    "10101010", --   53 - 0x35  :  170 - 0xaa
    "10101010", --   54 - 0x36  :  170 - 0xaa
    "00100010", --   55 - 0x37  :   34 - 0x22
    "00000000", --   56 - 0x38  :    0 - 0x0
    "00000000", --   57 - 0x39  :    0 - 0x0
    "00000000", --   58 - 0x3a  :    0 - 0x0
    "00000000", --   59 - 0x3b  :    0 - 0x0
    "00000000", --   60 - 0x3c  :    0 - 0x0
    "00000000", --   61 - 0x3d  :    0 - 0x0
    "00000000", --   62 - 0x3e  :    0 - 0x0
    "00000000", --   63 - 0x3f  :    0 - 0x0
    "00000000", --   64 - 0x40  :    0 - 0x0
    "00000000", --   65 - 0x41  :    0 - 0x0
    "00000000", --   66 - 0x42  :    0 - 0x0
    "00000000", --   67 - 0x43  :    0 - 0x0
    "00000000", --   68 - 0x44  :    0 - 0x0
    "00000000", --   69 - 0x45  :    0 - 0x0
    "00000000", --   70 - 0x46  :    0 - 0x0
    "00000000", --   71 - 0x47  :    0 - 0x0
    "00000000", --   72 - 0x48  :    0 - 0x0
    "00000000", --   73 - 0x49  :    0 - 0x0
    "00000000", --   74 - 0x4a  :    0 - 0x0
    "00000000", --   75 - 0x4b  :    0 - 0x0
    "00000000", --   76 - 0x4c  :    0 - 0x0
    "00000000", --   77 - 0x4d  :    0 - 0x0
    "00000000", --   78 - 0x4e  :    0 - 0x0
    "00000000", --   79 - 0x4f  :    0 - 0x0
    "00000000", --   80 - 0x50  :    0 - 0x0
    "00000000", --   81 - 0x51  :    0 - 0x0
    "00000000", --   82 - 0x52  :    0 - 0x0
    "00000000", --   83 - 0x53  :    0 - 0x0
    "00000000", --   84 - 0x54  :    0 - 0x0
    "00000000", --   85 - 0x55  :    0 - 0x0
    "00000000", --   86 - 0x56  :    0 - 0x0
    "00000000", --   87 - 0x57  :    0 - 0x0
    "00000000", --   88 - 0x58  :    0 - 0x0
    "00000000", --   89 - 0x59  :    0 - 0x0
    "00000000", --   90 - 0x5a  :    0 - 0x0
    "00000000", --   91 - 0x5b  :    0 - 0x0
    "00000000", --   92 - 0x5c  :    0 - 0x0
    "00000000", --   93 - 0x5d  :    0 - 0x0
    "00000000", --   94 - 0x5e  :    0 - 0x0
    "00000000", --   95 - 0x5f  :    0 - 0x0
    "00000000", --   96 - 0x60  :    0 - 0x0
    "00000000", --   97 - 0x61  :    0 - 0x0
    "00000000", --   98 - 0x62  :    0 - 0x0
    "00000000", --   99 - 0x63  :    0 - 0x0
    "00000000", --  100 - 0x64  :    0 - 0x0
    "00000000", --  101 - 0x65  :    0 - 0x0
    "00000000", --  102 - 0x66  :    0 - 0x0
    "00000000", --  103 - 0x67  :    0 - 0x0
    "00000000", --  104 - 0x68  :    0 - 0x0
    "00000000", --  105 - 0x69  :    0 - 0x0
    "00000000", --  106 - 0x6a  :    0 - 0x0
    "00000000", --  107 - 0x6b  :    0 - 0x0
    "00000000", --  108 - 0x6c  :    0 - 0x0
    "00000000", --  109 - 0x6d  :    0 - 0x0
    "00000000", --  110 - 0x6e  :    0 - 0x0
    "00000000", --  111 - 0x6f  :    0 - 0x0
    "00000000", --  112 - 0x70  :    0 - 0x0
    "00000000", --  113 - 0x71  :    0 - 0x0
    "00000000", --  114 - 0x72  :    0 - 0x0
    "00000000", --  115 - 0x73  :    0 - 0x0
    "00000000", --  116 - 0x74  :    0 - 0x0
    "00000000", --  117 - 0x75  :    0 - 0x0
    "00000000", --  118 - 0x76  :    0 - 0x0
    "00000000", --  119 - 0x77  :    0 - 0x0
    "00000000", --  120 - 0x78  :    0 - 0x0
    "00000000", --  121 - 0x79  :    0 - 0x0
    "00000000", --  122 - 0x7a  :    0 - 0x0
    "00000000", --  123 - 0x7b  :    0 - 0x0
    "00000000", --  124 - 0x7c  :    0 - 0x0
    "00000000", --  125 - 0x7d  :    0 - 0x0
    "00000000", --  126 - 0x7e  :    0 - 0x0
    "00000000"  --  127 - 0x7f  :    0 - 0x0
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
