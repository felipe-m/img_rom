//- Autcmatically generated verilog ROM from a NES memory file----
//-   PATTERN TABLE
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


//-  Original memory dump file name: sprilo_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_PTABLE_SPRILO
  (
     //input     clk,   // clock
     input      [13-1:0] addr,  //8192 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Pattern Table 0---------
      13'h0: dout  = 8'b00000000; //    0 :   0 - 0x0 -- Sprite 0x0
      13'h1: dout  = 8'b00000000; //    1 :   0 - 0x0
      13'h2: dout  = 8'b00000000; //    2 :   0 - 0x0
      13'h3: dout  = 8'b00000000; //    3 :   0 - 0x0
      13'h4: dout  = 8'b00000000; //    4 :   0 - 0x0
      13'h5: dout  = 8'b00000000; //    5 :   0 - 0x0
      13'h6: dout  = 8'b00000000; //    6 :   0 - 0x0
      13'h7: dout  = 8'b00000000; //    7 :   0 - 0x0
      13'h8: dout  = 8'b00000000; //    8 :   0 - 0x0
      13'h9: dout  = 8'b00000000; //    9 :   0 - 0x0
      13'hA: dout  = 8'b00000000; //   10 :   0 - 0x0
      13'hB: dout  = 8'b00000000; //   11 :   0 - 0x0
      13'hC: dout  = 8'b00000000; //   12 :   0 - 0x0
      13'hD: dout  = 8'b00000000; //   13 :   0 - 0x0
      13'hE: dout  = 8'b00000000; //   14 :   0 - 0x0
      13'hF: dout  = 8'b00000000; //   15 :   0 - 0x0
      13'h10: dout  = 8'b00000000; //   16 :   0 - 0x0 -- Sprite 0x1
      13'h11: dout  = 8'b00000000; //   17 :   0 - 0x0
      13'h12: dout  = 8'b00000000; //   18 :   0 - 0x0
      13'h13: dout  = 8'b00000000; //   19 :   0 - 0x0
      13'h14: dout  = 8'b00000000; //   20 :   0 - 0x0
      13'h15: dout  = 8'b00000000; //   21 :   0 - 0x0
      13'h16: dout  = 8'b00000000; //   22 :   0 - 0x0
      13'h17: dout  = 8'b00000000; //   23 :   0 - 0x0
      13'h18: dout  = 8'b00000000; //   24 :   0 - 0x0
      13'h19: dout  = 8'b00000000; //   25 :   0 - 0x0
      13'h1A: dout  = 8'b00000000; //   26 :   0 - 0x0
      13'h1B: dout  = 8'b00000000; //   27 :   0 - 0x0
      13'h1C: dout  = 8'b00000000; //   28 :   0 - 0x0
      13'h1D: dout  = 8'b00000000; //   29 :   0 - 0x0
      13'h1E: dout  = 8'b00000000; //   30 :   0 - 0x0
      13'h1F: dout  = 8'b00000000; //   31 :   0 - 0x0
      13'h20: dout  = 8'b00000000; //   32 :   0 - 0x0 -- Sprite 0x2
      13'h21: dout  = 8'b00000000; //   33 :   0 - 0x0
      13'h22: dout  = 8'b00000000; //   34 :   0 - 0x0
      13'h23: dout  = 8'b00000000; //   35 :   0 - 0x0
      13'h24: dout  = 8'b00000000; //   36 :   0 - 0x0
      13'h25: dout  = 8'b00000000; //   37 :   0 - 0x0
      13'h26: dout  = 8'b00000000; //   38 :   0 - 0x0
      13'h27: dout  = 8'b00000000; //   39 :   0 - 0x0
      13'h28: dout  = 8'b00000000; //   40 :   0 - 0x0
      13'h29: dout  = 8'b00000000; //   41 :   0 - 0x0
      13'h2A: dout  = 8'b00000000; //   42 :   0 - 0x0
      13'h2B: dout  = 8'b00000000; //   43 :   0 - 0x0
      13'h2C: dout  = 8'b00000000; //   44 :   0 - 0x0
      13'h2D: dout  = 8'b00000000; //   45 :   0 - 0x0
      13'h2E: dout  = 8'b00000000; //   46 :   0 - 0x0
      13'h2F: dout  = 8'b00000000; //   47 :   0 - 0x0
      13'h30: dout  = 8'b00000000; //   48 :   0 - 0x0 -- Sprite 0x3
      13'h31: dout  = 8'b00000000; //   49 :   0 - 0x0
      13'h32: dout  = 8'b00000000; //   50 :   0 - 0x0
      13'h33: dout  = 8'b00000000; //   51 :   0 - 0x0
      13'h34: dout  = 8'b00000000; //   52 :   0 - 0x0
      13'h35: dout  = 8'b00000000; //   53 :   0 - 0x0
      13'h36: dout  = 8'b00000000; //   54 :   0 - 0x0
      13'h37: dout  = 8'b00000000; //   55 :   0 - 0x0
      13'h38: dout  = 8'b00000000; //   56 :   0 - 0x0
      13'h39: dout  = 8'b00000000; //   57 :   0 - 0x0
      13'h3A: dout  = 8'b00000000; //   58 :   0 - 0x0
      13'h3B: dout  = 8'b00000000; //   59 :   0 - 0x0
      13'h3C: dout  = 8'b00000000; //   60 :   0 - 0x0
      13'h3D: dout  = 8'b00000000; //   61 :   0 - 0x0
      13'h3E: dout  = 8'b00000000; //   62 :   0 - 0x0
      13'h3F: dout  = 8'b00000000; //   63 :   0 - 0x0
      13'h40: dout  = 8'b00000000; //   64 :   0 - 0x0 -- Sprite 0x4
      13'h41: dout  = 8'b00000000; //   65 :   0 - 0x0
      13'h42: dout  = 8'b00000000; //   66 :   0 - 0x0
      13'h43: dout  = 8'b00000000; //   67 :   0 - 0x0
      13'h44: dout  = 8'b00000000; //   68 :   0 - 0x0
      13'h45: dout  = 8'b00000000; //   69 :   0 - 0x0
      13'h46: dout  = 8'b00000000; //   70 :   0 - 0x0
      13'h47: dout  = 8'b00000000; //   71 :   0 - 0x0
      13'h48: dout  = 8'b00000000; //   72 :   0 - 0x0
      13'h49: dout  = 8'b00000000; //   73 :   0 - 0x0
      13'h4A: dout  = 8'b00000000; //   74 :   0 - 0x0
      13'h4B: dout  = 8'b00000000; //   75 :   0 - 0x0
      13'h4C: dout  = 8'b00000000; //   76 :   0 - 0x0
      13'h4D: dout  = 8'b00000000; //   77 :   0 - 0x0
      13'h4E: dout  = 8'b00000000; //   78 :   0 - 0x0
      13'h4F: dout  = 8'b00000000; //   79 :   0 - 0x0
      13'h50: dout  = 8'b00000000; //   80 :   0 - 0x0 -- Sprite 0x5
      13'h51: dout  = 8'b00000000; //   81 :   0 - 0x0
      13'h52: dout  = 8'b00000000; //   82 :   0 - 0x0
      13'h53: dout  = 8'b00000000; //   83 :   0 - 0x0
      13'h54: dout  = 8'b00000000; //   84 :   0 - 0x0
      13'h55: dout  = 8'b00000000; //   85 :   0 - 0x0
      13'h56: dout  = 8'b00000000; //   86 :   0 - 0x0
      13'h57: dout  = 8'b00000000; //   87 :   0 - 0x0
      13'h58: dout  = 8'b00000000; //   88 :   0 - 0x0
      13'h59: dout  = 8'b00000000; //   89 :   0 - 0x0
      13'h5A: dout  = 8'b00000000; //   90 :   0 - 0x0
      13'h5B: dout  = 8'b00000000; //   91 :   0 - 0x0
      13'h5C: dout  = 8'b00000000; //   92 :   0 - 0x0
      13'h5D: dout  = 8'b00000000; //   93 :   0 - 0x0
      13'h5E: dout  = 8'b00000000; //   94 :   0 - 0x0
      13'h5F: dout  = 8'b00000000; //   95 :   0 - 0x0
      13'h60: dout  = 8'b00000000; //   96 :   0 - 0x0 -- Sprite 0x6
      13'h61: dout  = 8'b00000000; //   97 :   0 - 0x0
      13'h62: dout  = 8'b00000000; //   98 :   0 - 0x0
      13'h63: dout  = 8'b00000000; //   99 :   0 - 0x0
      13'h64: dout  = 8'b00000000; //  100 :   0 - 0x0
      13'h65: dout  = 8'b00000000; //  101 :   0 - 0x0
      13'h66: dout  = 8'b00000000; //  102 :   0 - 0x0
      13'h67: dout  = 8'b00000000; //  103 :   0 - 0x0
      13'h68: dout  = 8'b00000000; //  104 :   0 - 0x0
      13'h69: dout  = 8'b00000000; //  105 :   0 - 0x0
      13'h6A: dout  = 8'b00000000; //  106 :   0 - 0x0
      13'h6B: dout  = 8'b00000000; //  107 :   0 - 0x0
      13'h6C: dout  = 8'b00000000; //  108 :   0 - 0x0
      13'h6D: dout  = 8'b00000000; //  109 :   0 - 0x0
      13'h6E: dout  = 8'b00000000; //  110 :   0 - 0x0
      13'h6F: dout  = 8'b00000000; //  111 :   0 - 0x0
      13'h70: dout  = 8'b00000000; //  112 :   0 - 0x0 -- Sprite 0x7
      13'h71: dout  = 8'b00000000; //  113 :   0 - 0x0
      13'h72: dout  = 8'b00000000; //  114 :   0 - 0x0
      13'h73: dout  = 8'b00000000; //  115 :   0 - 0x0
      13'h74: dout  = 8'b00000000; //  116 :   0 - 0x0
      13'h75: dout  = 8'b00000000; //  117 :   0 - 0x0
      13'h76: dout  = 8'b00000000; //  118 :   0 - 0x0
      13'h77: dout  = 8'b00000000; //  119 :   0 - 0x0
      13'h78: dout  = 8'b00000000; //  120 :   0 - 0x0
      13'h79: dout  = 8'b00000000; //  121 :   0 - 0x0
      13'h7A: dout  = 8'b00000000; //  122 :   0 - 0x0
      13'h7B: dout  = 8'b00000000; //  123 :   0 - 0x0
      13'h7C: dout  = 8'b00000000; //  124 :   0 - 0x0
      13'h7D: dout  = 8'b00000000; //  125 :   0 - 0x0
      13'h7E: dout  = 8'b00000000; //  126 :   0 - 0x0
      13'h7F: dout  = 8'b00000000; //  127 :   0 - 0x0
      13'h80: dout  = 8'b00000000; //  128 :   0 - 0x0 -- Sprite 0x8
      13'h81: dout  = 8'b01111110; //  129 : 126 - 0x7e
      13'h82: dout  = 8'b01111110; //  130 : 126 - 0x7e
      13'h83: dout  = 8'b00111100; //  131 :  60 - 0x3c
      13'h84: dout  = 8'b00111100; //  132 :  60 - 0x3c
      13'h85: dout  = 8'b01111110; //  133 : 126 - 0x7e
      13'h86: dout  = 8'b01011010; //  134 :  90 - 0x5a
      13'h87: dout  = 8'b00000000; //  135 :   0 - 0x0
      13'h88: dout  = 8'b00000000; //  136 :   0 - 0x0
      13'h89: dout  = 8'b01000010; //  137 :  66 - 0x42
      13'h8A: dout  = 8'b01000010; //  138 :  66 - 0x42
      13'h8B: dout  = 8'b00000000; //  139 :   0 - 0x0
      13'h8C: dout  = 8'b00000000; //  140 :   0 - 0x0
      13'h8D: dout  = 8'b01000010; //  141 :  66 - 0x42
      13'h8E: dout  = 8'b01100110; //  142 : 102 - 0x66
      13'h8F: dout  = 8'b00000000; //  143 :   0 - 0x0
      13'h90: dout  = 8'b00000000; //  144 :   0 - 0x0 -- Sprite 0x9
      13'h91: dout  = 8'b01100110; //  145 : 102 - 0x66
      13'h92: dout  = 8'b01111100; //  146 : 124 - 0x7c
      13'h93: dout  = 8'b01111110; //  147 : 126 - 0x7e
      13'h94: dout  = 8'b01111110; //  148 : 126 - 0x7e
      13'h95: dout  = 8'b01111100; //  149 : 124 - 0x7c
      13'h96: dout  = 8'b01100110; //  150 : 102 - 0x66
      13'h97: dout  = 8'b00000000; //  151 :   0 - 0x0
      13'h98: dout  = 8'b00000000; //  152 :   0 - 0x0
      13'h99: dout  = 8'b01100110; //  153 : 102 - 0x66
      13'h9A: dout  = 8'b00000010; //  154 :   2 - 0x2
      13'h9B: dout  = 8'b00000000; //  155 :   0 - 0x0
      13'h9C: dout  = 8'b00000000; //  156 :   0 - 0x0
      13'h9D: dout  = 8'b00000010; //  157 :   2 - 0x2
      13'h9E: dout  = 8'b01100110; //  158 : 102 - 0x66
      13'h9F: dout  = 8'b00000000; //  159 :   0 - 0x0
      13'hA0: dout  = 8'b00010000; //  160 :  16 - 0x10 -- Sprite 0xa
      13'hA1: dout  = 8'b00011000; //  161 :  24 - 0x18
      13'hA2: dout  = 8'b00111000; //  162 :  56 - 0x38
      13'hA3: dout  = 8'b11111110; //  163 : 254 - 0xfe
      13'hA4: dout  = 8'b01111101; //  164 : 125 - 0x7d
      13'hA5: dout  = 8'b00011100; //  165 :  28 - 0x1c
      13'hA6: dout  = 8'b00010000; //  166 :  16 - 0x10
      13'hA7: dout  = 8'b00001000; //  167 :   8 - 0x8
      13'hA8: dout  = 8'b00010000; //  168 :  16 - 0x10
      13'hA9: dout  = 8'b00001000; //  169 :   8 - 0x8
      13'hAA: dout  = 8'b00000000; //  170 :   0 - 0x0
      13'hAB: dout  = 8'b10000010; //  171 : 130 - 0x82
      13'hAC: dout  = 8'b01000011; //  172 :  67 - 0x43
      13'hAD: dout  = 8'b00000000; //  173 :   0 - 0x0
      13'hAE: dout  = 8'b00011000; //  174 :  24 - 0x18
      13'hAF: dout  = 8'b00001000; //  175 :   8 - 0x8
      13'hB0: dout  = 8'b00000000; //  176 :   0 - 0x0 -- Sprite 0xb
      13'hB1: dout  = 8'b00000000; //  177 :   0 - 0x0
      13'hB2: dout  = 8'b00000000; //  178 :   0 - 0x0
      13'hB3: dout  = 8'b00000000; //  179 :   0 - 0x0
      13'hB4: dout  = 8'b00000000; //  180 :   0 - 0x0
      13'hB5: dout  = 8'b00000000; //  181 :   0 - 0x0
      13'hB6: dout  = 8'b00000000; //  182 :   0 - 0x0
      13'hB7: dout  = 8'b00000000; //  183 :   0 - 0x0
      13'hB8: dout  = 8'b00000000; //  184 :   0 - 0x0
      13'hB9: dout  = 8'b00000000; //  185 :   0 - 0x0
      13'hBA: dout  = 8'b00000000; //  186 :   0 - 0x0
      13'hBB: dout  = 8'b00000000; //  187 :   0 - 0x0
      13'hBC: dout  = 8'b00000000; //  188 :   0 - 0x0
      13'hBD: dout  = 8'b00000000; //  189 :   0 - 0x0
      13'hBE: dout  = 8'b00000000; //  190 :   0 - 0x0
      13'hBF: dout  = 8'b00000000; //  191 :   0 - 0x0
      13'hC0: dout  = 8'b00000000; //  192 :   0 - 0x0 -- Sprite 0xc
      13'hC1: dout  = 8'b00000000; //  193 :   0 - 0x0
      13'hC2: dout  = 8'b00000000; //  194 :   0 - 0x0
      13'hC3: dout  = 8'b00000000; //  195 :   0 - 0x0
      13'hC4: dout  = 8'b00000000; //  196 :   0 - 0x0
      13'hC5: dout  = 8'b00000000; //  197 :   0 - 0x0
      13'hC6: dout  = 8'b00000000; //  198 :   0 - 0x0
      13'hC7: dout  = 8'b00000000; //  199 :   0 - 0x0
      13'hC8: dout  = 8'b00000000; //  200 :   0 - 0x0
      13'hC9: dout  = 8'b00000000; //  201 :   0 - 0x0
      13'hCA: dout  = 8'b00000000; //  202 :   0 - 0x0
      13'hCB: dout  = 8'b00000000; //  203 :   0 - 0x0
      13'hCC: dout  = 8'b00000000; //  204 :   0 - 0x0
      13'hCD: dout  = 8'b00000000; //  205 :   0 - 0x0
      13'hCE: dout  = 8'b00000000; //  206 :   0 - 0x0
      13'hCF: dout  = 8'b00000000; //  207 :   0 - 0x0
      13'hD0: dout  = 8'b00000000; //  208 :   0 - 0x0 -- Sprite 0xd
      13'hD1: dout  = 8'b00000000; //  209 :   0 - 0x0
      13'hD2: dout  = 8'b00000000; //  210 :   0 - 0x0
      13'hD3: dout  = 8'b00000000; //  211 :   0 - 0x0
      13'hD4: dout  = 8'b00000000; //  212 :   0 - 0x0
      13'hD5: dout  = 8'b00000000; //  213 :   0 - 0x0
      13'hD6: dout  = 8'b00000000; //  214 :   0 - 0x0
      13'hD7: dout  = 8'b00000000; //  215 :   0 - 0x0
      13'hD8: dout  = 8'b00000000; //  216 :   0 - 0x0
      13'hD9: dout  = 8'b00000000; //  217 :   0 - 0x0
      13'hDA: dout  = 8'b00000000; //  218 :   0 - 0x0
      13'hDB: dout  = 8'b00000000; //  219 :   0 - 0x0
      13'hDC: dout  = 8'b00000000; //  220 :   0 - 0x0
      13'hDD: dout  = 8'b00000000; //  221 :   0 - 0x0
      13'hDE: dout  = 8'b00000000; //  222 :   0 - 0x0
      13'hDF: dout  = 8'b00000000; //  223 :   0 - 0x0
      13'hE0: dout  = 8'b00000000; //  224 :   0 - 0x0 -- Sprite 0xe
      13'hE1: dout  = 8'b00000000; //  225 :   0 - 0x0
      13'hE2: dout  = 8'b00000000; //  226 :   0 - 0x0
      13'hE3: dout  = 8'b00000000; //  227 :   0 - 0x0
      13'hE4: dout  = 8'b00000000; //  228 :   0 - 0x0
      13'hE5: dout  = 8'b00000000; //  229 :   0 - 0x0
      13'hE6: dout  = 8'b00000000; //  230 :   0 - 0x0
      13'hE7: dout  = 8'b00000000; //  231 :   0 - 0x0
      13'hE8: dout  = 8'b00000000; //  232 :   0 - 0x0
      13'hE9: dout  = 8'b00000000; //  233 :   0 - 0x0
      13'hEA: dout  = 8'b00000000; //  234 :   0 - 0x0
      13'hEB: dout  = 8'b00000000; //  235 :   0 - 0x0
      13'hEC: dout  = 8'b00000000; //  236 :   0 - 0x0
      13'hED: dout  = 8'b00000000; //  237 :   0 - 0x0
      13'hEE: dout  = 8'b00000000; //  238 :   0 - 0x0
      13'hEF: dout  = 8'b00000000; //  239 :   0 - 0x0
      13'hF0: dout  = 8'b00000000; //  240 :   0 - 0x0 -- Sprite 0xf
      13'hF1: dout  = 8'b00000000; //  241 :   0 - 0x0
      13'hF2: dout  = 8'b00000000; //  242 :   0 - 0x0
      13'hF3: dout  = 8'b00000000; //  243 :   0 - 0x0
      13'hF4: dout  = 8'b00000000; //  244 :   0 - 0x0
      13'hF5: dout  = 8'b00000000; //  245 :   0 - 0x0
      13'hF6: dout  = 8'b00000000; //  246 :   0 - 0x0
      13'hF7: dout  = 8'b00000000; //  247 :   0 - 0x0
      13'hF8: dout  = 8'b00000000; //  248 :   0 - 0x0
      13'hF9: dout  = 8'b00000000; //  249 :   0 - 0x0
      13'hFA: dout  = 8'b00000000; //  250 :   0 - 0x0
      13'hFB: dout  = 8'b00000000; //  251 :   0 - 0x0
      13'hFC: dout  = 8'b00000000; //  252 :   0 - 0x0
      13'hFD: dout  = 8'b00000000; //  253 :   0 - 0x0
      13'hFE: dout  = 8'b00000000; //  254 :   0 - 0x0
      13'hFF: dout  = 8'b00000000; //  255 :   0 - 0x0
      13'h100: dout  = 8'b00000000; //  256 :   0 - 0x0 -- Sprite 0x10
      13'h101: dout  = 8'b00000000; //  257 :   0 - 0x0
      13'h102: dout  = 8'b00000000; //  258 :   0 - 0x0
      13'h103: dout  = 8'b00000000; //  259 :   0 - 0x0
      13'h104: dout  = 8'b00000000; //  260 :   0 - 0x0
      13'h105: dout  = 8'b00000000; //  261 :   0 - 0x0
      13'h106: dout  = 8'b00000000; //  262 :   0 - 0x0
      13'h107: dout  = 8'b00000000; //  263 :   0 - 0x0
      13'h108: dout  = 8'b00000000; //  264 :   0 - 0x0
      13'h109: dout  = 8'b00000000; //  265 :   0 - 0x0
      13'h10A: dout  = 8'b00000000; //  266 :   0 - 0x0
      13'h10B: dout  = 8'b00000000; //  267 :   0 - 0x0
      13'h10C: dout  = 8'b00000000; //  268 :   0 - 0x0
      13'h10D: dout  = 8'b00000000; //  269 :   0 - 0x0
      13'h10E: dout  = 8'b00000000; //  270 :   0 - 0x0
      13'h10F: dout  = 8'b00000000; //  271 :   0 - 0x0
      13'h110: dout  = 8'b00000000; //  272 :   0 - 0x0 -- Sprite 0x11
      13'h111: dout  = 8'b00000000; //  273 :   0 - 0x0
      13'h112: dout  = 8'b00000000; //  274 :   0 - 0x0
      13'h113: dout  = 8'b00000000; //  275 :   0 - 0x0
      13'h114: dout  = 8'b00000000; //  276 :   0 - 0x0
      13'h115: dout  = 8'b00000000; //  277 :   0 - 0x0
      13'h116: dout  = 8'b00000000; //  278 :   0 - 0x0
      13'h117: dout  = 8'b00000000; //  279 :   0 - 0x0
      13'h118: dout  = 8'b00000000; //  280 :   0 - 0x0
      13'h119: dout  = 8'b00000000; //  281 :   0 - 0x0
      13'h11A: dout  = 8'b00000000; //  282 :   0 - 0x0
      13'h11B: dout  = 8'b00000000; //  283 :   0 - 0x0
      13'h11C: dout  = 8'b00000000; //  284 :   0 - 0x0
      13'h11D: dout  = 8'b00000000; //  285 :   0 - 0x0
      13'h11E: dout  = 8'b00000000; //  286 :   0 - 0x0
      13'h11F: dout  = 8'b00000000; //  287 :   0 - 0x0
      13'h120: dout  = 8'b00000000; //  288 :   0 - 0x0 -- Sprite 0x12
      13'h121: dout  = 8'b00000000; //  289 :   0 - 0x0
      13'h122: dout  = 8'b00000000; //  290 :   0 - 0x0
      13'h123: dout  = 8'b00000000; //  291 :   0 - 0x0
      13'h124: dout  = 8'b00000000; //  292 :   0 - 0x0
      13'h125: dout  = 8'b00000000; //  293 :   0 - 0x0
      13'h126: dout  = 8'b00000000; //  294 :   0 - 0x0
      13'h127: dout  = 8'b00000000; //  295 :   0 - 0x0
      13'h128: dout  = 8'b00000000; //  296 :   0 - 0x0
      13'h129: dout  = 8'b00000000; //  297 :   0 - 0x0
      13'h12A: dout  = 8'b00000000; //  298 :   0 - 0x0
      13'h12B: dout  = 8'b00000000; //  299 :   0 - 0x0
      13'h12C: dout  = 8'b00000000; //  300 :   0 - 0x0
      13'h12D: dout  = 8'b00000000; //  301 :   0 - 0x0
      13'h12E: dout  = 8'b00000000; //  302 :   0 - 0x0
      13'h12F: dout  = 8'b00000000; //  303 :   0 - 0x0
      13'h130: dout  = 8'b00000000; //  304 :   0 - 0x0 -- Sprite 0x13
      13'h131: dout  = 8'b00000000; //  305 :   0 - 0x0
      13'h132: dout  = 8'b00000000; //  306 :   0 - 0x0
      13'h133: dout  = 8'b00000000; //  307 :   0 - 0x0
      13'h134: dout  = 8'b00000000; //  308 :   0 - 0x0
      13'h135: dout  = 8'b00000000; //  309 :   0 - 0x0
      13'h136: dout  = 8'b00000000; //  310 :   0 - 0x0
      13'h137: dout  = 8'b00000000; //  311 :   0 - 0x0
      13'h138: dout  = 8'b00000000; //  312 :   0 - 0x0
      13'h139: dout  = 8'b00000000; //  313 :   0 - 0x0
      13'h13A: dout  = 8'b00000000; //  314 :   0 - 0x0
      13'h13B: dout  = 8'b00000000; //  315 :   0 - 0x0
      13'h13C: dout  = 8'b00000000; //  316 :   0 - 0x0
      13'h13D: dout  = 8'b00000000; //  317 :   0 - 0x0
      13'h13E: dout  = 8'b00000000; //  318 :   0 - 0x0
      13'h13F: dout  = 8'b00000000; //  319 :   0 - 0x0
      13'h140: dout  = 8'b00000000; //  320 :   0 - 0x0 -- Sprite 0x14
      13'h141: dout  = 8'b00000000; //  321 :   0 - 0x0
      13'h142: dout  = 8'b00000000; //  322 :   0 - 0x0
      13'h143: dout  = 8'b00000000; //  323 :   0 - 0x0
      13'h144: dout  = 8'b00000000; //  324 :   0 - 0x0
      13'h145: dout  = 8'b00000000; //  325 :   0 - 0x0
      13'h146: dout  = 8'b00000000; //  326 :   0 - 0x0
      13'h147: dout  = 8'b00000000; //  327 :   0 - 0x0
      13'h148: dout  = 8'b00000000; //  328 :   0 - 0x0
      13'h149: dout  = 8'b00000000; //  329 :   0 - 0x0
      13'h14A: dout  = 8'b00000000; //  330 :   0 - 0x0
      13'h14B: dout  = 8'b00000000; //  331 :   0 - 0x0
      13'h14C: dout  = 8'b00000000; //  332 :   0 - 0x0
      13'h14D: dout  = 8'b00000000; //  333 :   0 - 0x0
      13'h14E: dout  = 8'b00000000; //  334 :   0 - 0x0
      13'h14F: dout  = 8'b00000000; //  335 :   0 - 0x0
      13'h150: dout  = 8'b00000000; //  336 :   0 - 0x0 -- Sprite 0x15
      13'h151: dout  = 8'b00000000; //  337 :   0 - 0x0
      13'h152: dout  = 8'b00000000; //  338 :   0 - 0x0
      13'h153: dout  = 8'b00000000; //  339 :   0 - 0x0
      13'h154: dout  = 8'b00000000; //  340 :   0 - 0x0
      13'h155: dout  = 8'b00000000; //  341 :   0 - 0x0
      13'h156: dout  = 8'b00000000; //  342 :   0 - 0x0
      13'h157: dout  = 8'b00000000; //  343 :   0 - 0x0
      13'h158: dout  = 8'b00000000; //  344 :   0 - 0x0
      13'h159: dout  = 8'b00000000; //  345 :   0 - 0x0
      13'h15A: dout  = 8'b00000000; //  346 :   0 - 0x0
      13'h15B: dout  = 8'b00000000; //  347 :   0 - 0x0
      13'h15C: dout  = 8'b00000000; //  348 :   0 - 0x0
      13'h15D: dout  = 8'b00000000; //  349 :   0 - 0x0
      13'h15E: dout  = 8'b00000000; //  350 :   0 - 0x0
      13'h15F: dout  = 8'b00000000; //  351 :   0 - 0x0
      13'h160: dout  = 8'b00000000; //  352 :   0 - 0x0 -- Sprite 0x16
      13'h161: dout  = 8'b00000000; //  353 :   0 - 0x0
      13'h162: dout  = 8'b00000000; //  354 :   0 - 0x0
      13'h163: dout  = 8'b00000000; //  355 :   0 - 0x0
      13'h164: dout  = 8'b00000000; //  356 :   0 - 0x0
      13'h165: dout  = 8'b00000000; //  357 :   0 - 0x0
      13'h166: dout  = 8'b00000000; //  358 :   0 - 0x0
      13'h167: dout  = 8'b00000000; //  359 :   0 - 0x0
      13'h168: dout  = 8'b00000000; //  360 :   0 - 0x0
      13'h169: dout  = 8'b00000000; //  361 :   0 - 0x0
      13'h16A: dout  = 8'b00000000; //  362 :   0 - 0x0
      13'h16B: dout  = 8'b00000000; //  363 :   0 - 0x0
      13'h16C: dout  = 8'b00000000; //  364 :   0 - 0x0
      13'h16D: dout  = 8'b00000000; //  365 :   0 - 0x0
      13'h16E: dout  = 8'b00000000; //  366 :   0 - 0x0
      13'h16F: dout  = 8'b00000000; //  367 :   0 - 0x0
      13'h170: dout  = 8'b00000000; //  368 :   0 - 0x0 -- Sprite 0x17
      13'h171: dout  = 8'b00000000; //  369 :   0 - 0x0
      13'h172: dout  = 8'b00000000; //  370 :   0 - 0x0
      13'h173: dout  = 8'b00000000; //  371 :   0 - 0x0
      13'h174: dout  = 8'b00000000; //  372 :   0 - 0x0
      13'h175: dout  = 8'b00000000; //  373 :   0 - 0x0
      13'h176: dout  = 8'b00000000; //  374 :   0 - 0x0
      13'h177: dout  = 8'b00000000; //  375 :   0 - 0x0
      13'h178: dout  = 8'b00000000; //  376 :   0 - 0x0
      13'h179: dout  = 8'b00000000; //  377 :   0 - 0x0
      13'h17A: dout  = 8'b00000000; //  378 :   0 - 0x0
      13'h17B: dout  = 8'b00000000; //  379 :   0 - 0x0
      13'h17C: dout  = 8'b00000000; //  380 :   0 - 0x0
      13'h17D: dout  = 8'b00000000; //  381 :   0 - 0x0
      13'h17E: dout  = 8'b00000000; //  382 :   0 - 0x0
      13'h17F: dout  = 8'b00000000; //  383 :   0 - 0x0
      13'h180: dout  = 8'b00000000; //  384 :   0 - 0x0 -- Sprite 0x18
      13'h181: dout  = 8'b00000000; //  385 :   0 - 0x0
      13'h182: dout  = 8'b00000000; //  386 :   0 - 0x0
      13'h183: dout  = 8'b00000000; //  387 :   0 - 0x0
      13'h184: dout  = 8'b00000000; //  388 :   0 - 0x0
      13'h185: dout  = 8'b00000000; //  389 :   0 - 0x0
      13'h186: dout  = 8'b00000000; //  390 :   0 - 0x0
      13'h187: dout  = 8'b00000000; //  391 :   0 - 0x0
      13'h188: dout  = 8'b00000000; //  392 :   0 - 0x0
      13'h189: dout  = 8'b00000000; //  393 :   0 - 0x0
      13'h18A: dout  = 8'b00000000; //  394 :   0 - 0x0
      13'h18B: dout  = 8'b00000000; //  395 :   0 - 0x0
      13'h18C: dout  = 8'b00000000; //  396 :   0 - 0x0
      13'h18D: dout  = 8'b00000000; //  397 :   0 - 0x0
      13'h18E: dout  = 8'b00000000; //  398 :   0 - 0x0
      13'h18F: dout  = 8'b00000000; //  399 :   0 - 0x0
      13'h190: dout  = 8'b00000000; //  400 :   0 - 0x0 -- Sprite 0x19
      13'h191: dout  = 8'b00000000; //  401 :   0 - 0x0
      13'h192: dout  = 8'b00000000; //  402 :   0 - 0x0
      13'h193: dout  = 8'b00000000; //  403 :   0 - 0x0
      13'h194: dout  = 8'b00000000; //  404 :   0 - 0x0
      13'h195: dout  = 8'b00000000; //  405 :   0 - 0x0
      13'h196: dout  = 8'b00000000; //  406 :   0 - 0x0
      13'h197: dout  = 8'b00000000; //  407 :   0 - 0x0
      13'h198: dout  = 8'b00000000; //  408 :   0 - 0x0
      13'h199: dout  = 8'b00000000; //  409 :   0 - 0x0
      13'h19A: dout  = 8'b00000000; //  410 :   0 - 0x0
      13'h19B: dout  = 8'b00000000; //  411 :   0 - 0x0
      13'h19C: dout  = 8'b00000000; //  412 :   0 - 0x0
      13'h19D: dout  = 8'b00000000; //  413 :   0 - 0x0
      13'h19E: dout  = 8'b00000000; //  414 :   0 - 0x0
      13'h19F: dout  = 8'b00000000; //  415 :   0 - 0x0
      13'h1A0: dout  = 8'b00000000; //  416 :   0 - 0x0 -- Sprite 0x1a
      13'h1A1: dout  = 8'b00000000; //  417 :   0 - 0x0
      13'h1A2: dout  = 8'b00000000; //  418 :   0 - 0x0
      13'h1A3: dout  = 8'b00000000; //  419 :   0 - 0x0
      13'h1A4: dout  = 8'b00000000; //  420 :   0 - 0x0
      13'h1A5: dout  = 8'b00000000; //  421 :   0 - 0x0
      13'h1A6: dout  = 8'b00000000; //  422 :   0 - 0x0
      13'h1A7: dout  = 8'b00000000; //  423 :   0 - 0x0
      13'h1A8: dout  = 8'b00000000; //  424 :   0 - 0x0
      13'h1A9: dout  = 8'b00000000; //  425 :   0 - 0x0
      13'h1AA: dout  = 8'b00000000; //  426 :   0 - 0x0
      13'h1AB: dout  = 8'b00000000; //  427 :   0 - 0x0
      13'h1AC: dout  = 8'b00000000; //  428 :   0 - 0x0
      13'h1AD: dout  = 8'b00000000; //  429 :   0 - 0x0
      13'h1AE: dout  = 8'b00000000; //  430 :   0 - 0x0
      13'h1AF: dout  = 8'b00000000; //  431 :   0 - 0x0
      13'h1B0: dout  = 8'b00000000; //  432 :   0 - 0x0 -- Sprite 0x1b
      13'h1B1: dout  = 8'b00000000; //  433 :   0 - 0x0
      13'h1B2: dout  = 8'b00000000; //  434 :   0 - 0x0
      13'h1B3: dout  = 8'b00000000; //  435 :   0 - 0x0
      13'h1B4: dout  = 8'b00000000; //  436 :   0 - 0x0
      13'h1B5: dout  = 8'b00000000; //  437 :   0 - 0x0
      13'h1B6: dout  = 8'b00000000; //  438 :   0 - 0x0
      13'h1B7: dout  = 8'b00000000; //  439 :   0 - 0x0
      13'h1B8: dout  = 8'b00000000; //  440 :   0 - 0x0
      13'h1B9: dout  = 8'b00000000; //  441 :   0 - 0x0
      13'h1BA: dout  = 8'b00000000; //  442 :   0 - 0x0
      13'h1BB: dout  = 8'b00000000; //  443 :   0 - 0x0
      13'h1BC: dout  = 8'b00000000; //  444 :   0 - 0x0
      13'h1BD: dout  = 8'b00000000; //  445 :   0 - 0x0
      13'h1BE: dout  = 8'b00000000; //  446 :   0 - 0x0
      13'h1BF: dout  = 8'b00000000; //  447 :   0 - 0x0
      13'h1C0: dout  = 8'b00000000; //  448 :   0 - 0x0 -- Sprite 0x1c
      13'h1C1: dout  = 8'b00000000; //  449 :   0 - 0x0
      13'h1C2: dout  = 8'b00000000; //  450 :   0 - 0x0
      13'h1C3: dout  = 8'b00000000; //  451 :   0 - 0x0
      13'h1C4: dout  = 8'b00000000; //  452 :   0 - 0x0
      13'h1C5: dout  = 8'b00000000; //  453 :   0 - 0x0
      13'h1C6: dout  = 8'b00000000; //  454 :   0 - 0x0
      13'h1C7: dout  = 8'b00000000; //  455 :   0 - 0x0
      13'h1C8: dout  = 8'b00000000; //  456 :   0 - 0x0
      13'h1C9: dout  = 8'b00000000; //  457 :   0 - 0x0
      13'h1CA: dout  = 8'b00000000; //  458 :   0 - 0x0
      13'h1CB: dout  = 8'b00000000; //  459 :   0 - 0x0
      13'h1CC: dout  = 8'b00000000; //  460 :   0 - 0x0
      13'h1CD: dout  = 8'b00000000; //  461 :   0 - 0x0
      13'h1CE: dout  = 8'b00000000; //  462 :   0 - 0x0
      13'h1CF: dout  = 8'b00000000; //  463 :   0 - 0x0
      13'h1D0: dout  = 8'b00000000; //  464 :   0 - 0x0 -- Sprite 0x1d
      13'h1D1: dout  = 8'b00000000; //  465 :   0 - 0x0
      13'h1D2: dout  = 8'b00000000; //  466 :   0 - 0x0
      13'h1D3: dout  = 8'b00000000; //  467 :   0 - 0x0
      13'h1D4: dout  = 8'b00000000; //  468 :   0 - 0x0
      13'h1D5: dout  = 8'b00000000; //  469 :   0 - 0x0
      13'h1D6: dout  = 8'b00000000; //  470 :   0 - 0x0
      13'h1D7: dout  = 8'b00000000; //  471 :   0 - 0x0
      13'h1D8: dout  = 8'b00000000; //  472 :   0 - 0x0
      13'h1D9: dout  = 8'b00000000; //  473 :   0 - 0x0
      13'h1DA: dout  = 8'b00000000; //  474 :   0 - 0x0
      13'h1DB: dout  = 8'b00000000; //  475 :   0 - 0x0
      13'h1DC: dout  = 8'b00000000; //  476 :   0 - 0x0
      13'h1DD: dout  = 8'b00000000; //  477 :   0 - 0x0
      13'h1DE: dout  = 8'b00000000; //  478 :   0 - 0x0
      13'h1DF: dout  = 8'b00000000; //  479 :   0 - 0x0
      13'h1E0: dout  = 8'b00000000; //  480 :   0 - 0x0 -- Sprite 0x1e
      13'h1E1: dout  = 8'b00000000; //  481 :   0 - 0x0
      13'h1E2: dout  = 8'b00000000; //  482 :   0 - 0x0
      13'h1E3: dout  = 8'b00000000; //  483 :   0 - 0x0
      13'h1E4: dout  = 8'b00000000; //  484 :   0 - 0x0
      13'h1E5: dout  = 8'b00000000; //  485 :   0 - 0x0
      13'h1E6: dout  = 8'b00000000; //  486 :   0 - 0x0
      13'h1E7: dout  = 8'b00000000; //  487 :   0 - 0x0
      13'h1E8: dout  = 8'b00000000; //  488 :   0 - 0x0
      13'h1E9: dout  = 8'b00000000; //  489 :   0 - 0x0
      13'h1EA: dout  = 8'b00000000; //  490 :   0 - 0x0
      13'h1EB: dout  = 8'b00000000; //  491 :   0 - 0x0
      13'h1EC: dout  = 8'b00000000; //  492 :   0 - 0x0
      13'h1ED: dout  = 8'b00000000; //  493 :   0 - 0x0
      13'h1EE: dout  = 8'b00000000; //  494 :   0 - 0x0
      13'h1EF: dout  = 8'b00000000; //  495 :   0 - 0x0
      13'h1F0: dout  = 8'b00000000; //  496 :   0 - 0x0 -- Sprite 0x1f
      13'h1F1: dout  = 8'b00000000; //  497 :   0 - 0x0
      13'h1F2: dout  = 8'b00000000; //  498 :   0 - 0x0
      13'h1F3: dout  = 8'b00000000; //  499 :   0 - 0x0
      13'h1F4: dout  = 8'b00000000; //  500 :   0 - 0x0
      13'h1F5: dout  = 8'b00000000; //  501 :   0 - 0x0
      13'h1F6: dout  = 8'b00000000; //  502 :   0 - 0x0
      13'h1F7: dout  = 8'b00000000; //  503 :   0 - 0x0
      13'h1F8: dout  = 8'b00000000; //  504 :   0 - 0x0
      13'h1F9: dout  = 8'b00000000; //  505 :   0 - 0x0
      13'h1FA: dout  = 8'b00000000; //  506 :   0 - 0x0
      13'h1FB: dout  = 8'b00000000; //  507 :   0 - 0x0
      13'h1FC: dout  = 8'b00000000; //  508 :   0 - 0x0
      13'h1FD: dout  = 8'b00000000; //  509 :   0 - 0x0
      13'h1FE: dout  = 8'b00000000; //  510 :   0 - 0x0
      13'h1FF: dout  = 8'b00000000; //  511 :   0 - 0x0
      13'h200: dout  = 8'b00000000; //  512 :   0 - 0x0 -- Sprite 0x20
      13'h201: dout  = 8'b00000000; //  513 :   0 - 0x0
      13'h202: dout  = 8'b00000000; //  514 :   0 - 0x0
      13'h203: dout  = 8'b00000000; //  515 :   0 - 0x0
      13'h204: dout  = 8'b00000000; //  516 :   0 - 0x0
      13'h205: dout  = 8'b00000000; //  517 :   0 - 0x0
      13'h206: dout  = 8'b00000000; //  518 :   0 - 0x0
      13'h207: dout  = 8'b00000000; //  519 :   0 - 0x0
      13'h208: dout  = 8'b00000000; //  520 :   0 - 0x0
      13'h209: dout  = 8'b00000000; //  521 :   0 - 0x0
      13'h20A: dout  = 8'b00000000; //  522 :   0 - 0x0
      13'h20B: dout  = 8'b00000000; //  523 :   0 - 0x0
      13'h20C: dout  = 8'b00000000; //  524 :   0 - 0x0
      13'h20D: dout  = 8'b00000000; //  525 :   0 - 0x0
      13'h20E: dout  = 8'b00000000; //  526 :   0 - 0x0
      13'h20F: dout  = 8'b00000000; //  527 :   0 - 0x0
      13'h210: dout  = 8'b00000000; //  528 :   0 - 0x0 -- Sprite 0x21
      13'h211: dout  = 8'b00000000; //  529 :   0 - 0x0
      13'h212: dout  = 8'b00000000; //  530 :   0 - 0x0
      13'h213: dout  = 8'b00000000; //  531 :   0 - 0x0
      13'h214: dout  = 8'b00000000; //  532 :   0 - 0x0
      13'h215: dout  = 8'b00000000; //  533 :   0 - 0x0
      13'h216: dout  = 8'b00000000; //  534 :   0 - 0x0
      13'h217: dout  = 8'b00000000; //  535 :   0 - 0x0
      13'h218: dout  = 8'b00000000; //  536 :   0 - 0x0
      13'h219: dout  = 8'b00000000; //  537 :   0 - 0x0
      13'h21A: dout  = 8'b00000000; //  538 :   0 - 0x0
      13'h21B: dout  = 8'b00000000; //  539 :   0 - 0x0
      13'h21C: dout  = 8'b00000000; //  540 :   0 - 0x0
      13'h21D: dout  = 8'b00000000; //  541 :   0 - 0x0
      13'h21E: dout  = 8'b00000000; //  542 :   0 - 0x0
      13'h21F: dout  = 8'b00000000; //  543 :   0 - 0x0
      13'h220: dout  = 8'b00000000; //  544 :   0 - 0x0 -- Sprite 0x22
      13'h221: dout  = 8'b00000000; //  545 :   0 - 0x0
      13'h222: dout  = 8'b00000000; //  546 :   0 - 0x0
      13'h223: dout  = 8'b00000000; //  547 :   0 - 0x0
      13'h224: dout  = 8'b00000000; //  548 :   0 - 0x0
      13'h225: dout  = 8'b00000000; //  549 :   0 - 0x0
      13'h226: dout  = 8'b00000000; //  550 :   0 - 0x0
      13'h227: dout  = 8'b00000000; //  551 :   0 - 0x0
      13'h228: dout  = 8'b00000000; //  552 :   0 - 0x0
      13'h229: dout  = 8'b00000000; //  553 :   0 - 0x0
      13'h22A: dout  = 8'b00000000; //  554 :   0 - 0x0
      13'h22B: dout  = 8'b00000000; //  555 :   0 - 0x0
      13'h22C: dout  = 8'b00000000; //  556 :   0 - 0x0
      13'h22D: dout  = 8'b00000000; //  557 :   0 - 0x0
      13'h22E: dout  = 8'b00000000; //  558 :   0 - 0x0
      13'h22F: dout  = 8'b00000000; //  559 :   0 - 0x0
      13'h230: dout  = 8'b00000000; //  560 :   0 - 0x0 -- Sprite 0x23
      13'h231: dout  = 8'b00000000; //  561 :   0 - 0x0
      13'h232: dout  = 8'b00000000; //  562 :   0 - 0x0
      13'h233: dout  = 8'b00000000; //  563 :   0 - 0x0
      13'h234: dout  = 8'b00000000; //  564 :   0 - 0x0
      13'h235: dout  = 8'b00000000; //  565 :   0 - 0x0
      13'h236: dout  = 8'b00000000; //  566 :   0 - 0x0
      13'h237: dout  = 8'b00000000; //  567 :   0 - 0x0
      13'h238: dout  = 8'b00000000; //  568 :   0 - 0x0
      13'h239: dout  = 8'b00000000; //  569 :   0 - 0x0
      13'h23A: dout  = 8'b00000000; //  570 :   0 - 0x0
      13'h23B: dout  = 8'b00000000; //  571 :   0 - 0x0
      13'h23C: dout  = 8'b00000000; //  572 :   0 - 0x0
      13'h23D: dout  = 8'b00000000; //  573 :   0 - 0x0
      13'h23E: dout  = 8'b00000000; //  574 :   0 - 0x0
      13'h23F: dout  = 8'b00000000; //  575 :   0 - 0x0
      13'h240: dout  = 8'b00000000; //  576 :   0 - 0x0 -- Sprite 0x24
      13'h241: dout  = 8'b00000000; //  577 :   0 - 0x0
      13'h242: dout  = 8'b00000000; //  578 :   0 - 0x0
      13'h243: dout  = 8'b00000000; //  579 :   0 - 0x0
      13'h244: dout  = 8'b00000000; //  580 :   0 - 0x0
      13'h245: dout  = 8'b00000000; //  581 :   0 - 0x0
      13'h246: dout  = 8'b00000000; //  582 :   0 - 0x0
      13'h247: dout  = 8'b00000000; //  583 :   0 - 0x0
      13'h248: dout  = 8'b00000000; //  584 :   0 - 0x0
      13'h249: dout  = 8'b00000000; //  585 :   0 - 0x0
      13'h24A: dout  = 8'b00000000; //  586 :   0 - 0x0
      13'h24B: dout  = 8'b00000000; //  587 :   0 - 0x0
      13'h24C: dout  = 8'b00000000; //  588 :   0 - 0x0
      13'h24D: dout  = 8'b00000000; //  589 :   0 - 0x0
      13'h24E: dout  = 8'b00000000; //  590 :   0 - 0x0
      13'h24F: dout  = 8'b00000000; //  591 :   0 - 0x0
      13'h250: dout  = 8'b00000000; //  592 :   0 - 0x0 -- Sprite 0x25
      13'h251: dout  = 8'b00000000; //  593 :   0 - 0x0
      13'h252: dout  = 8'b00000000; //  594 :   0 - 0x0
      13'h253: dout  = 8'b00000000; //  595 :   0 - 0x0
      13'h254: dout  = 8'b00000000; //  596 :   0 - 0x0
      13'h255: dout  = 8'b00000000; //  597 :   0 - 0x0
      13'h256: dout  = 8'b00000000; //  598 :   0 - 0x0
      13'h257: dout  = 8'b00000000; //  599 :   0 - 0x0
      13'h258: dout  = 8'b00000000; //  600 :   0 - 0x0
      13'h259: dout  = 8'b00000000; //  601 :   0 - 0x0
      13'h25A: dout  = 8'b00000000; //  602 :   0 - 0x0
      13'h25B: dout  = 8'b00000000; //  603 :   0 - 0x0
      13'h25C: dout  = 8'b00000000; //  604 :   0 - 0x0
      13'h25D: dout  = 8'b00000000; //  605 :   0 - 0x0
      13'h25E: dout  = 8'b00000000; //  606 :   0 - 0x0
      13'h25F: dout  = 8'b00000000; //  607 :   0 - 0x0
      13'h260: dout  = 8'b00000000; //  608 :   0 - 0x0 -- Sprite 0x26
      13'h261: dout  = 8'b00000000; //  609 :   0 - 0x0
      13'h262: dout  = 8'b00000000; //  610 :   0 - 0x0
      13'h263: dout  = 8'b00000000; //  611 :   0 - 0x0
      13'h264: dout  = 8'b00000000; //  612 :   0 - 0x0
      13'h265: dout  = 8'b00000000; //  613 :   0 - 0x0
      13'h266: dout  = 8'b00000000; //  614 :   0 - 0x0
      13'h267: dout  = 8'b00000000; //  615 :   0 - 0x0
      13'h268: dout  = 8'b00000000; //  616 :   0 - 0x0
      13'h269: dout  = 8'b00000000; //  617 :   0 - 0x0
      13'h26A: dout  = 8'b00000000; //  618 :   0 - 0x0
      13'h26B: dout  = 8'b00000000; //  619 :   0 - 0x0
      13'h26C: dout  = 8'b00000000; //  620 :   0 - 0x0
      13'h26D: dout  = 8'b00000000; //  621 :   0 - 0x0
      13'h26E: dout  = 8'b00000000; //  622 :   0 - 0x0
      13'h26F: dout  = 8'b00000000; //  623 :   0 - 0x0
      13'h270: dout  = 8'b00000000; //  624 :   0 - 0x0 -- Sprite 0x27
      13'h271: dout  = 8'b00000000; //  625 :   0 - 0x0
      13'h272: dout  = 8'b00000000; //  626 :   0 - 0x0
      13'h273: dout  = 8'b00000000; //  627 :   0 - 0x0
      13'h274: dout  = 8'b00000000; //  628 :   0 - 0x0
      13'h275: dout  = 8'b00000000; //  629 :   0 - 0x0
      13'h276: dout  = 8'b00000000; //  630 :   0 - 0x0
      13'h277: dout  = 8'b00000000; //  631 :   0 - 0x0
      13'h278: dout  = 8'b00000000; //  632 :   0 - 0x0
      13'h279: dout  = 8'b00000000; //  633 :   0 - 0x0
      13'h27A: dout  = 8'b00000000; //  634 :   0 - 0x0
      13'h27B: dout  = 8'b00000000; //  635 :   0 - 0x0
      13'h27C: dout  = 8'b00000000; //  636 :   0 - 0x0
      13'h27D: dout  = 8'b00000000; //  637 :   0 - 0x0
      13'h27E: dout  = 8'b00000000; //  638 :   0 - 0x0
      13'h27F: dout  = 8'b00000000; //  639 :   0 - 0x0
      13'h280: dout  = 8'b00000000; //  640 :   0 - 0x0 -- Sprite 0x28
      13'h281: dout  = 8'b00000000; //  641 :   0 - 0x0
      13'h282: dout  = 8'b00000000; //  642 :   0 - 0x0
      13'h283: dout  = 8'b00000000; //  643 :   0 - 0x0
      13'h284: dout  = 8'b00000000; //  644 :   0 - 0x0
      13'h285: dout  = 8'b00000000; //  645 :   0 - 0x0
      13'h286: dout  = 8'b00000000; //  646 :   0 - 0x0
      13'h287: dout  = 8'b00000000; //  647 :   0 - 0x0
      13'h288: dout  = 8'b00000000; //  648 :   0 - 0x0
      13'h289: dout  = 8'b00000000; //  649 :   0 - 0x0
      13'h28A: dout  = 8'b00000000; //  650 :   0 - 0x0
      13'h28B: dout  = 8'b00000000; //  651 :   0 - 0x0
      13'h28C: dout  = 8'b00000000; //  652 :   0 - 0x0
      13'h28D: dout  = 8'b00000000; //  653 :   0 - 0x0
      13'h28E: dout  = 8'b00000000; //  654 :   0 - 0x0
      13'h28F: dout  = 8'b00000000; //  655 :   0 - 0x0
      13'h290: dout  = 8'b00000000; //  656 :   0 - 0x0 -- Sprite 0x29
      13'h291: dout  = 8'b00000000; //  657 :   0 - 0x0
      13'h292: dout  = 8'b00000000; //  658 :   0 - 0x0
      13'h293: dout  = 8'b00000000; //  659 :   0 - 0x0
      13'h294: dout  = 8'b00000000; //  660 :   0 - 0x0
      13'h295: dout  = 8'b00000000; //  661 :   0 - 0x0
      13'h296: dout  = 8'b00000000; //  662 :   0 - 0x0
      13'h297: dout  = 8'b00000000; //  663 :   0 - 0x0
      13'h298: dout  = 8'b00000000; //  664 :   0 - 0x0
      13'h299: dout  = 8'b00000000; //  665 :   0 - 0x0
      13'h29A: dout  = 8'b00000000; //  666 :   0 - 0x0
      13'h29B: dout  = 8'b00000000; //  667 :   0 - 0x0
      13'h29C: dout  = 8'b00000000; //  668 :   0 - 0x0
      13'h29D: dout  = 8'b00000000; //  669 :   0 - 0x0
      13'h29E: dout  = 8'b00000000; //  670 :   0 - 0x0
      13'h29F: dout  = 8'b00000000; //  671 :   0 - 0x0
      13'h2A0: dout  = 8'b00000000; //  672 :   0 - 0x0 -- Sprite 0x2a
      13'h2A1: dout  = 8'b00000000; //  673 :   0 - 0x0
      13'h2A2: dout  = 8'b00000000; //  674 :   0 - 0x0
      13'h2A3: dout  = 8'b00000000; //  675 :   0 - 0x0
      13'h2A4: dout  = 8'b00000000; //  676 :   0 - 0x0
      13'h2A5: dout  = 8'b00000000; //  677 :   0 - 0x0
      13'h2A6: dout  = 8'b00000000; //  678 :   0 - 0x0
      13'h2A7: dout  = 8'b00000000; //  679 :   0 - 0x0
      13'h2A8: dout  = 8'b00000000; //  680 :   0 - 0x0
      13'h2A9: dout  = 8'b00000000; //  681 :   0 - 0x0
      13'h2AA: dout  = 8'b00000000; //  682 :   0 - 0x0
      13'h2AB: dout  = 8'b00000000; //  683 :   0 - 0x0
      13'h2AC: dout  = 8'b00000000; //  684 :   0 - 0x0
      13'h2AD: dout  = 8'b00000000; //  685 :   0 - 0x0
      13'h2AE: dout  = 8'b00000000; //  686 :   0 - 0x0
      13'h2AF: dout  = 8'b00000000; //  687 :   0 - 0x0
      13'h2B0: dout  = 8'b00000000; //  688 :   0 - 0x0 -- Sprite 0x2b
      13'h2B1: dout  = 8'b00000000; //  689 :   0 - 0x0
      13'h2B2: dout  = 8'b00000000; //  690 :   0 - 0x0
      13'h2B3: dout  = 8'b00000000; //  691 :   0 - 0x0
      13'h2B4: dout  = 8'b00000000; //  692 :   0 - 0x0
      13'h2B5: dout  = 8'b00000000; //  693 :   0 - 0x0
      13'h2B6: dout  = 8'b00000000; //  694 :   0 - 0x0
      13'h2B7: dout  = 8'b00000000; //  695 :   0 - 0x0
      13'h2B8: dout  = 8'b00000000; //  696 :   0 - 0x0
      13'h2B9: dout  = 8'b00000000; //  697 :   0 - 0x0
      13'h2BA: dout  = 8'b00000000; //  698 :   0 - 0x0
      13'h2BB: dout  = 8'b00000000; //  699 :   0 - 0x0
      13'h2BC: dout  = 8'b00000000; //  700 :   0 - 0x0
      13'h2BD: dout  = 8'b00000000; //  701 :   0 - 0x0
      13'h2BE: dout  = 8'b00000000; //  702 :   0 - 0x0
      13'h2BF: dout  = 8'b00000000; //  703 :   0 - 0x0
      13'h2C0: dout  = 8'b00000000; //  704 :   0 - 0x0 -- Sprite 0x2c
      13'h2C1: dout  = 8'b00000000; //  705 :   0 - 0x0
      13'h2C2: dout  = 8'b00000000; //  706 :   0 - 0x0
      13'h2C3: dout  = 8'b00000000; //  707 :   0 - 0x0
      13'h2C4: dout  = 8'b00000000; //  708 :   0 - 0x0
      13'h2C5: dout  = 8'b00000000; //  709 :   0 - 0x0
      13'h2C6: dout  = 8'b00000000; //  710 :   0 - 0x0
      13'h2C7: dout  = 8'b00000000; //  711 :   0 - 0x0
      13'h2C8: dout  = 8'b00000000; //  712 :   0 - 0x0
      13'h2C9: dout  = 8'b00000000; //  713 :   0 - 0x0
      13'h2CA: dout  = 8'b00000000; //  714 :   0 - 0x0
      13'h2CB: dout  = 8'b00000000; //  715 :   0 - 0x0
      13'h2CC: dout  = 8'b00000000; //  716 :   0 - 0x0
      13'h2CD: dout  = 8'b00000000; //  717 :   0 - 0x0
      13'h2CE: dout  = 8'b00000000; //  718 :   0 - 0x0
      13'h2CF: dout  = 8'b00000000; //  719 :   0 - 0x0
      13'h2D0: dout  = 8'b00000000; //  720 :   0 - 0x0 -- Sprite 0x2d
      13'h2D1: dout  = 8'b00000000; //  721 :   0 - 0x0
      13'h2D2: dout  = 8'b00000000; //  722 :   0 - 0x0
      13'h2D3: dout  = 8'b00000000; //  723 :   0 - 0x0
      13'h2D4: dout  = 8'b00000000; //  724 :   0 - 0x0
      13'h2D5: dout  = 8'b00000000; //  725 :   0 - 0x0
      13'h2D6: dout  = 8'b00000000; //  726 :   0 - 0x0
      13'h2D7: dout  = 8'b00000000; //  727 :   0 - 0x0
      13'h2D8: dout  = 8'b00000000; //  728 :   0 - 0x0
      13'h2D9: dout  = 8'b00000000; //  729 :   0 - 0x0
      13'h2DA: dout  = 8'b00000000; //  730 :   0 - 0x0
      13'h2DB: dout  = 8'b00000000; //  731 :   0 - 0x0
      13'h2DC: dout  = 8'b00000000; //  732 :   0 - 0x0
      13'h2DD: dout  = 8'b00000000; //  733 :   0 - 0x0
      13'h2DE: dout  = 8'b00000000; //  734 :   0 - 0x0
      13'h2DF: dout  = 8'b00000000; //  735 :   0 - 0x0
      13'h2E0: dout  = 8'b00000000; //  736 :   0 - 0x0 -- Sprite 0x2e
      13'h2E1: dout  = 8'b00000000; //  737 :   0 - 0x0
      13'h2E2: dout  = 8'b00000000; //  738 :   0 - 0x0
      13'h2E3: dout  = 8'b00000000; //  739 :   0 - 0x0
      13'h2E4: dout  = 8'b00000000; //  740 :   0 - 0x0
      13'h2E5: dout  = 8'b00000000; //  741 :   0 - 0x0
      13'h2E6: dout  = 8'b00000000; //  742 :   0 - 0x0
      13'h2E7: dout  = 8'b00000000; //  743 :   0 - 0x0
      13'h2E8: dout  = 8'b00000000; //  744 :   0 - 0x0
      13'h2E9: dout  = 8'b00000000; //  745 :   0 - 0x0
      13'h2EA: dout  = 8'b00000000; //  746 :   0 - 0x0
      13'h2EB: dout  = 8'b00000000; //  747 :   0 - 0x0
      13'h2EC: dout  = 8'b00000000; //  748 :   0 - 0x0
      13'h2ED: dout  = 8'b00000000; //  749 :   0 - 0x0
      13'h2EE: dout  = 8'b00000000; //  750 :   0 - 0x0
      13'h2EF: dout  = 8'b00000000; //  751 :   0 - 0x0
      13'h2F0: dout  = 8'b00000000; //  752 :   0 - 0x0 -- Sprite 0x2f
      13'h2F1: dout  = 8'b00000000; //  753 :   0 - 0x0
      13'h2F2: dout  = 8'b00000000; //  754 :   0 - 0x0
      13'h2F3: dout  = 8'b00000000; //  755 :   0 - 0x0
      13'h2F4: dout  = 8'b00000000; //  756 :   0 - 0x0
      13'h2F5: dout  = 8'b00000000; //  757 :   0 - 0x0
      13'h2F6: dout  = 8'b00000000; //  758 :   0 - 0x0
      13'h2F7: dout  = 8'b00000000; //  759 :   0 - 0x0
      13'h2F8: dout  = 8'b00000000; //  760 :   0 - 0x0
      13'h2F9: dout  = 8'b00000000; //  761 :   0 - 0x0
      13'h2FA: dout  = 8'b00000000; //  762 :   0 - 0x0
      13'h2FB: dout  = 8'b00000000; //  763 :   0 - 0x0
      13'h2FC: dout  = 8'b00000000; //  764 :   0 - 0x0
      13'h2FD: dout  = 8'b00000000; //  765 :   0 - 0x0
      13'h2FE: dout  = 8'b00000000; //  766 :   0 - 0x0
      13'h2FF: dout  = 8'b00000000; //  767 :   0 - 0x0
      13'h300: dout  = 8'b00000000; //  768 :   0 - 0x0 -- Sprite 0x30
      13'h301: dout  = 8'b00000000; //  769 :   0 - 0x0
      13'h302: dout  = 8'b00000000; //  770 :   0 - 0x0
      13'h303: dout  = 8'b00000000; //  771 :   0 - 0x0
      13'h304: dout  = 8'b00000000; //  772 :   0 - 0x0
      13'h305: dout  = 8'b00000000; //  773 :   0 - 0x0
      13'h306: dout  = 8'b00000000; //  774 :   0 - 0x0
      13'h307: dout  = 8'b00000000; //  775 :   0 - 0x0
      13'h308: dout  = 8'b00000000; //  776 :   0 - 0x0
      13'h309: dout  = 8'b00000000; //  777 :   0 - 0x0
      13'h30A: dout  = 8'b00000000; //  778 :   0 - 0x0
      13'h30B: dout  = 8'b00000000; //  779 :   0 - 0x0
      13'h30C: dout  = 8'b00000000; //  780 :   0 - 0x0
      13'h30D: dout  = 8'b00000000; //  781 :   0 - 0x0
      13'h30E: dout  = 8'b00000000; //  782 :   0 - 0x0
      13'h30F: dout  = 8'b00000000; //  783 :   0 - 0x0
      13'h310: dout  = 8'b00000000; //  784 :   0 - 0x0 -- Sprite 0x31
      13'h311: dout  = 8'b00000000; //  785 :   0 - 0x0
      13'h312: dout  = 8'b00000000; //  786 :   0 - 0x0
      13'h313: dout  = 8'b00000000; //  787 :   0 - 0x0
      13'h314: dout  = 8'b00000000; //  788 :   0 - 0x0
      13'h315: dout  = 8'b00000000; //  789 :   0 - 0x0
      13'h316: dout  = 8'b00000000; //  790 :   0 - 0x0
      13'h317: dout  = 8'b00000000; //  791 :   0 - 0x0
      13'h318: dout  = 8'b00000000; //  792 :   0 - 0x0
      13'h319: dout  = 8'b00000000; //  793 :   0 - 0x0
      13'h31A: dout  = 8'b00000000; //  794 :   0 - 0x0
      13'h31B: dout  = 8'b00000000; //  795 :   0 - 0x0
      13'h31C: dout  = 8'b00000000; //  796 :   0 - 0x0
      13'h31D: dout  = 8'b00000000; //  797 :   0 - 0x0
      13'h31E: dout  = 8'b00000000; //  798 :   0 - 0x0
      13'h31F: dout  = 8'b00000000; //  799 :   0 - 0x0
      13'h320: dout  = 8'b00000000; //  800 :   0 - 0x0 -- Sprite 0x32
      13'h321: dout  = 8'b00000000; //  801 :   0 - 0x0
      13'h322: dout  = 8'b00000000; //  802 :   0 - 0x0
      13'h323: dout  = 8'b00000000; //  803 :   0 - 0x0
      13'h324: dout  = 8'b00000000; //  804 :   0 - 0x0
      13'h325: dout  = 8'b00000000; //  805 :   0 - 0x0
      13'h326: dout  = 8'b00000000; //  806 :   0 - 0x0
      13'h327: dout  = 8'b00000000; //  807 :   0 - 0x0
      13'h328: dout  = 8'b00000000; //  808 :   0 - 0x0
      13'h329: dout  = 8'b00000000; //  809 :   0 - 0x0
      13'h32A: dout  = 8'b00000000; //  810 :   0 - 0x0
      13'h32B: dout  = 8'b00000000; //  811 :   0 - 0x0
      13'h32C: dout  = 8'b00000000; //  812 :   0 - 0x0
      13'h32D: dout  = 8'b00000000; //  813 :   0 - 0x0
      13'h32E: dout  = 8'b00000000; //  814 :   0 - 0x0
      13'h32F: dout  = 8'b00000000; //  815 :   0 - 0x0
      13'h330: dout  = 8'b00000000; //  816 :   0 - 0x0 -- Sprite 0x33
      13'h331: dout  = 8'b00000000; //  817 :   0 - 0x0
      13'h332: dout  = 8'b00000000; //  818 :   0 - 0x0
      13'h333: dout  = 8'b00000000; //  819 :   0 - 0x0
      13'h334: dout  = 8'b00000000; //  820 :   0 - 0x0
      13'h335: dout  = 8'b00000000; //  821 :   0 - 0x0
      13'h336: dout  = 8'b00000000; //  822 :   0 - 0x0
      13'h337: dout  = 8'b00000000; //  823 :   0 - 0x0
      13'h338: dout  = 8'b00000000; //  824 :   0 - 0x0
      13'h339: dout  = 8'b00000000; //  825 :   0 - 0x0
      13'h33A: dout  = 8'b00000000; //  826 :   0 - 0x0
      13'h33B: dout  = 8'b00000000; //  827 :   0 - 0x0
      13'h33C: dout  = 8'b00000000; //  828 :   0 - 0x0
      13'h33D: dout  = 8'b00000000; //  829 :   0 - 0x0
      13'h33E: dout  = 8'b00000000; //  830 :   0 - 0x0
      13'h33F: dout  = 8'b00000000; //  831 :   0 - 0x0
      13'h340: dout  = 8'b00000000; //  832 :   0 - 0x0 -- Sprite 0x34
      13'h341: dout  = 8'b00000000; //  833 :   0 - 0x0
      13'h342: dout  = 8'b00000000; //  834 :   0 - 0x0
      13'h343: dout  = 8'b00000000; //  835 :   0 - 0x0
      13'h344: dout  = 8'b00000000; //  836 :   0 - 0x0
      13'h345: dout  = 8'b00000000; //  837 :   0 - 0x0
      13'h346: dout  = 8'b00000000; //  838 :   0 - 0x0
      13'h347: dout  = 8'b00000000; //  839 :   0 - 0x0
      13'h348: dout  = 8'b00000000; //  840 :   0 - 0x0
      13'h349: dout  = 8'b00000000; //  841 :   0 - 0x0
      13'h34A: dout  = 8'b00000000; //  842 :   0 - 0x0
      13'h34B: dout  = 8'b00000000; //  843 :   0 - 0x0
      13'h34C: dout  = 8'b00000000; //  844 :   0 - 0x0
      13'h34D: dout  = 8'b00000000; //  845 :   0 - 0x0
      13'h34E: dout  = 8'b00000000; //  846 :   0 - 0x0
      13'h34F: dout  = 8'b00000000; //  847 :   0 - 0x0
      13'h350: dout  = 8'b00000000; //  848 :   0 - 0x0 -- Sprite 0x35
      13'h351: dout  = 8'b00000000; //  849 :   0 - 0x0
      13'h352: dout  = 8'b00000000; //  850 :   0 - 0x0
      13'h353: dout  = 8'b00000000; //  851 :   0 - 0x0
      13'h354: dout  = 8'b00000000; //  852 :   0 - 0x0
      13'h355: dout  = 8'b00000000; //  853 :   0 - 0x0
      13'h356: dout  = 8'b00000000; //  854 :   0 - 0x0
      13'h357: dout  = 8'b00000000; //  855 :   0 - 0x0
      13'h358: dout  = 8'b00000000; //  856 :   0 - 0x0
      13'h359: dout  = 8'b00000000; //  857 :   0 - 0x0
      13'h35A: dout  = 8'b00000000; //  858 :   0 - 0x0
      13'h35B: dout  = 8'b00000000; //  859 :   0 - 0x0
      13'h35C: dout  = 8'b00000000; //  860 :   0 - 0x0
      13'h35D: dout  = 8'b00000000; //  861 :   0 - 0x0
      13'h35E: dout  = 8'b00000000; //  862 :   0 - 0x0
      13'h35F: dout  = 8'b00000000; //  863 :   0 - 0x0
      13'h360: dout  = 8'b00000000; //  864 :   0 - 0x0 -- Sprite 0x36
      13'h361: dout  = 8'b00000000; //  865 :   0 - 0x0
      13'h362: dout  = 8'b00000000; //  866 :   0 - 0x0
      13'h363: dout  = 8'b00000000; //  867 :   0 - 0x0
      13'h364: dout  = 8'b00000000; //  868 :   0 - 0x0
      13'h365: dout  = 8'b00000000; //  869 :   0 - 0x0
      13'h366: dout  = 8'b00000000; //  870 :   0 - 0x0
      13'h367: dout  = 8'b00000000; //  871 :   0 - 0x0
      13'h368: dout  = 8'b00000000; //  872 :   0 - 0x0
      13'h369: dout  = 8'b00000000; //  873 :   0 - 0x0
      13'h36A: dout  = 8'b00000000; //  874 :   0 - 0x0
      13'h36B: dout  = 8'b00000000; //  875 :   0 - 0x0
      13'h36C: dout  = 8'b00000000; //  876 :   0 - 0x0
      13'h36D: dout  = 8'b00000000; //  877 :   0 - 0x0
      13'h36E: dout  = 8'b00000000; //  878 :   0 - 0x0
      13'h36F: dout  = 8'b00000000; //  879 :   0 - 0x0
      13'h370: dout  = 8'b00000000; //  880 :   0 - 0x0 -- Sprite 0x37
      13'h371: dout  = 8'b00000000; //  881 :   0 - 0x0
      13'h372: dout  = 8'b00000000; //  882 :   0 - 0x0
      13'h373: dout  = 8'b00000000; //  883 :   0 - 0x0
      13'h374: dout  = 8'b00000000; //  884 :   0 - 0x0
      13'h375: dout  = 8'b00000000; //  885 :   0 - 0x0
      13'h376: dout  = 8'b00000000; //  886 :   0 - 0x0
      13'h377: dout  = 8'b00000000; //  887 :   0 - 0x0
      13'h378: dout  = 8'b00000000; //  888 :   0 - 0x0
      13'h379: dout  = 8'b00000000; //  889 :   0 - 0x0
      13'h37A: dout  = 8'b00000000; //  890 :   0 - 0x0
      13'h37B: dout  = 8'b00000000; //  891 :   0 - 0x0
      13'h37C: dout  = 8'b00000000; //  892 :   0 - 0x0
      13'h37D: dout  = 8'b00000000; //  893 :   0 - 0x0
      13'h37E: dout  = 8'b00000000; //  894 :   0 - 0x0
      13'h37F: dout  = 8'b00000000; //  895 :   0 - 0x0
      13'h380: dout  = 8'b00000000; //  896 :   0 - 0x0 -- Sprite 0x38
      13'h381: dout  = 8'b00000000; //  897 :   0 - 0x0
      13'h382: dout  = 8'b00000000; //  898 :   0 - 0x0
      13'h383: dout  = 8'b00000000; //  899 :   0 - 0x0
      13'h384: dout  = 8'b00000000; //  900 :   0 - 0x0
      13'h385: dout  = 8'b00000000; //  901 :   0 - 0x0
      13'h386: dout  = 8'b00000000; //  902 :   0 - 0x0
      13'h387: dout  = 8'b00000000; //  903 :   0 - 0x0
      13'h388: dout  = 8'b00000000; //  904 :   0 - 0x0
      13'h389: dout  = 8'b00000000; //  905 :   0 - 0x0
      13'h38A: dout  = 8'b00000000; //  906 :   0 - 0x0
      13'h38B: dout  = 8'b00000000; //  907 :   0 - 0x0
      13'h38C: dout  = 8'b00000000; //  908 :   0 - 0x0
      13'h38D: dout  = 8'b00000000; //  909 :   0 - 0x0
      13'h38E: dout  = 8'b00000000; //  910 :   0 - 0x0
      13'h38F: dout  = 8'b00000000; //  911 :   0 - 0x0
      13'h390: dout  = 8'b00000000; //  912 :   0 - 0x0 -- Sprite 0x39
      13'h391: dout  = 8'b00000000; //  913 :   0 - 0x0
      13'h392: dout  = 8'b00000000; //  914 :   0 - 0x0
      13'h393: dout  = 8'b00000000; //  915 :   0 - 0x0
      13'h394: dout  = 8'b00000000; //  916 :   0 - 0x0
      13'h395: dout  = 8'b00000000; //  917 :   0 - 0x0
      13'h396: dout  = 8'b00000000; //  918 :   0 - 0x0
      13'h397: dout  = 8'b00000000; //  919 :   0 - 0x0
      13'h398: dout  = 8'b00000000; //  920 :   0 - 0x0
      13'h399: dout  = 8'b00000000; //  921 :   0 - 0x0
      13'h39A: dout  = 8'b00000000; //  922 :   0 - 0x0
      13'h39B: dout  = 8'b00000000; //  923 :   0 - 0x0
      13'h39C: dout  = 8'b00000000; //  924 :   0 - 0x0
      13'h39D: dout  = 8'b00000000; //  925 :   0 - 0x0
      13'h39E: dout  = 8'b00000000; //  926 :   0 - 0x0
      13'h39F: dout  = 8'b00000000; //  927 :   0 - 0x0
      13'h3A0: dout  = 8'b00000000; //  928 :   0 - 0x0 -- Sprite 0x3a
      13'h3A1: dout  = 8'b00000000; //  929 :   0 - 0x0
      13'h3A2: dout  = 8'b00000000; //  930 :   0 - 0x0
      13'h3A3: dout  = 8'b00000000; //  931 :   0 - 0x0
      13'h3A4: dout  = 8'b00000000; //  932 :   0 - 0x0
      13'h3A5: dout  = 8'b00000000; //  933 :   0 - 0x0
      13'h3A6: dout  = 8'b00000000; //  934 :   0 - 0x0
      13'h3A7: dout  = 8'b00000000; //  935 :   0 - 0x0
      13'h3A8: dout  = 8'b00000000; //  936 :   0 - 0x0
      13'h3A9: dout  = 8'b00000000; //  937 :   0 - 0x0
      13'h3AA: dout  = 8'b00000000; //  938 :   0 - 0x0
      13'h3AB: dout  = 8'b00000000; //  939 :   0 - 0x0
      13'h3AC: dout  = 8'b00000000; //  940 :   0 - 0x0
      13'h3AD: dout  = 8'b00000000; //  941 :   0 - 0x0
      13'h3AE: dout  = 8'b00000000; //  942 :   0 - 0x0
      13'h3AF: dout  = 8'b00000000; //  943 :   0 - 0x0
      13'h3B0: dout  = 8'b00000000; //  944 :   0 - 0x0 -- Sprite 0x3b
      13'h3B1: dout  = 8'b00000000; //  945 :   0 - 0x0
      13'h3B2: dout  = 8'b00000000; //  946 :   0 - 0x0
      13'h3B3: dout  = 8'b00000000; //  947 :   0 - 0x0
      13'h3B4: dout  = 8'b00000000; //  948 :   0 - 0x0
      13'h3B5: dout  = 8'b00000000; //  949 :   0 - 0x0
      13'h3B6: dout  = 8'b00000000; //  950 :   0 - 0x0
      13'h3B7: dout  = 8'b00000000; //  951 :   0 - 0x0
      13'h3B8: dout  = 8'b00000000; //  952 :   0 - 0x0
      13'h3B9: dout  = 8'b00000000; //  953 :   0 - 0x0
      13'h3BA: dout  = 8'b00000000; //  954 :   0 - 0x0
      13'h3BB: dout  = 8'b00000000; //  955 :   0 - 0x0
      13'h3BC: dout  = 8'b00000000; //  956 :   0 - 0x0
      13'h3BD: dout  = 8'b00000000; //  957 :   0 - 0x0
      13'h3BE: dout  = 8'b00000000; //  958 :   0 - 0x0
      13'h3BF: dout  = 8'b00000000; //  959 :   0 - 0x0
      13'h3C0: dout  = 8'b00000000; //  960 :   0 - 0x0 -- Sprite 0x3c
      13'h3C1: dout  = 8'b00000000; //  961 :   0 - 0x0
      13'h3C2: dout  = 8'b00000000; //  962 :   0 - 0x0
      13'h3C3: dout  = 8'b00000000; //  963 :   0 - 0x0
      13'h3C4: dout  = 8'b00000000; //  964 :   0 - 0x0
      13'h3C5: dout  = 8'b00000000; //  965 :   0 - 0x0
      13'h3C6: dout  = 8'b00000000; //  966 :   0 - 0x0
      13'h3C7: dout  = 8'b00000000; //  967 :   0 - 0x0
      13'h3C8: dout  = 8'b00000000; //  968 :   0 - 0x0
      13'h3C9: dout  = 8'b00000000; //  969 :   0 - 0x0
      13'h3CA: dout  = 8'b00000000; //  970 :   0 - 0x0
      13'h3CB: dout  = 8'b00000000; //  971 :   0 - 0x0
      13'h3CC: dout  = 8'b00000000; //  972 :   0 - 0x0
      13'h3CD: dout  = 8'b00000000; //  973 :   0 - 0x0
      13'h3CE: dout  = 8'b00000000; //  974 :   0 - 0x0
      13'h3CF: dout  = 8'b00000000; //  975 :   0 - 0x0
      13'h3D0: dout  = 8'b00000000; //  976 :   0 - 0x0 -- Sprite 0x3d
      13'h3D1: dout  = 8'b00000000; //  977 :   0 - 0x0
      13'h3D2: dout  = 8'b00000000; //  978 :   0 - 0x0
      13'h3D3: dout  = 8'b00000000; //  979 :   0 - 0x0
      13'h3D4: dout  = 8'b00000000; //  980 :   0 - 0x0
      13'h3D5: dout  = 8'b00000000; //  981 :   0 - 0x0
      13'h3D6: dout  = 8'b00000000; //  982 :   0 - 0x0
      13'h3D7: dout  = 8'b00000000; //  983 :   0 - 0x0
      13'h3D8: dout  = 8'b00000000; //  984 :   0 - 0x0
      13'h3D9: dout  = 8'b00000000; //  985 :   0 - 0x0
      13'h3DA: dout  = 8'b00000000; //  986 :   0 - 0x0
      13'h3DB: dout  = 8'b00000000; //  987 :   0 - 0x0
      13'h3DC: dout  = 8'b00000000; //  988 :   0 - 0x0
      13'h3DD: dout  = 8'b00000000; //  989 :   0 - 0x0
      13'h3DE: dout  = 8'b00000000; //  990 :   0 - 0x0
      13'h3DF: dout  = 8'b00000000; //  991 :   0 - 0x0
      13'h3E0: dout  = 8'b00000000; //  992 :   0 - 0x0 -- Sprite 0x3e
      13'h3E1: dout  = 8'b00000000; //  993 :   0 - 0x0
      13'h3E2: dout  = 8'b00000000; //  994 :   0 - 0x0
      13'h3E3: dout  = 8'b00000000; //  995 :   0 - 0x0
      13'h3E4: dout  = 8'b00000000; //  996 :   0 - 0x0
      13'h3E5: dout  = 8'b00000000; //  997 :   0 - 0x0
      13'h3E6: dout  = 8'b00000000; //  998 :   0 - 0x0
      13'h3E7: dout  = 8'b00000000; //  999 :   0 - 0x0
      13'h3E8: dout  = 8'b00000000; // 1000 :   0 - 0x0
      13'h3E9: dout  = 8'b00000000; // 1001 :   0 - 0x0
      13'h3EA: dout  = 8'b00000000; // 1002 :   0 - 0x0
      13'h3EB: dout  = 8'b00000000; // 1003 :   0 - 0x0
      13'h3EC: dout  = 8'b00000000; // 1004 :   0 - 0x0
      13'h3ED: dout  = 8'b00000000; // 1005 :   0 - 0x0
      13'h3EE: dout  = 8'b00000000; // 1006 :   0 - 0x0
      13'h3EF: dout  = 8'b00000000; // 1007 :   0 - 0x0
      13'h3F0: dout  = 8'b00000000; // 1008 :   0 - 0x0 -- Sprite 0x3f
      13'h3F1: dout  = 8'b00000000; // 1009 :   0 - 0x0
      13'h3F2: dout  = 8'b00000000; // 1010 :   0 - 0x0
      13'h3F3: dout  = 8'b00000000; // 1011 :   0 - 0x0
      13'h3F4: dout  = 8'b00000000; // 1012 :   0 - 0x0
      13'h3F5: dout  = 8'b00000000; // 1013 :   0 - 0x0
      13'h3F6: dout  = 8'b00000000; // 1014 :   0 - 0x0
      13'h3F7: dout  = 8'b00000000; // 1015 :   0 - 0x0
      13'h3F8: dout  = 8'b00000000; // 1016 :   0 - 0x0
      13'h3F9: dout  = 8'b00000000; // 1017 :   0 - 0x0
      13'h3FA: dout  = 8'b00000000; // 1018 :   0 - 0x0
      13'h3FB: dout  = 8'b00000000; // 1019 :   0 - 0x0
      13'h3FC: dout  = 8'b00000000; // 1020 :   0 - 0x0
      13'h3FD: dout  = 8'b00000000; // 1021 :   0 - 0x0
      13'h3FE: dout  = 8'b00000000; // 1022 :   0 - 0x0
      13'h3FF: dout  = 8'b00000000; // 1023 :   0 - 0x0
      13'h400: dout  = 8'b00000000; // 1024 :   0 - 0x0 -- Sprite 0x40
      13'h401: dout  = 8'b00000000; // 1025 :   0 - 0x0
      13'h402: dout  = 8'b00000000; // 1026 :   0 - 0x0
      13'h403: dout  = 8'b00000000; // 1027 :   0 - 0x0
      13'h404: dout  = 8'b00000000; // 1028 :   0 - 0x0
      13'h405: dout  = 8'b00000000; // 1029 :   0 - 0x0
      13'h406: dout  = 8'b00000000; // 1030 :   0 - 0x0
      13'h407: dout  = 8'b00000000; // 1031 :   0 - 0x0
      13'h408: dout  = 8'b00000000; // 1032 :   0 - 0x0
      13'h409: dout  = 8'b00000000; // 1033 :   0 - 0x0
      13'h40A: dout  = 8'b00000000; // 1034 :   0 - 0x0
      13'h40B: dout  = 8'b00000000; // 1035 :   0 - 0x0
      13'h40C: dout  = 8'b00000000; // 1036 :   0 - 0x0
      13'h40D: dout  = 8'b00000000; // 1037 :   0 - 0x0
      13'h40E: dout  = 8'b00000000; // 1038 :   0 - 0x0
      13'h40F: dout  = 8'b00000000; // 1039 :   0 - 0x0
      13'h410: dout  = 8'b00000000; // 1040 :   0 - 0x0 -- Sprite 0x41
      13'h411: dout  = 8'b00000000; // 1041 :   0 - 0x0
      13'h412: dout  = 8'b00000000; // 1042 :   0 - 0x0
      13'h413: dout  = 8'b00000000; // 1043 :   0 - 0x0
      13'h414: dout  = 8'b00000000; // 1044 :   0 - 0x0
      13'h415: dout  = 8'b00000000; // 1045 :   0 - 0x0
      13'h416: dout  = 8'b00000000; // 1046 :   0 - 0x0
      13'h417: dout  = 8'b00000000; // 1047 :   0 - 0x0
      13'h418: dout  = 8'b00000000; // 1048 :   0 - 0x0
      13'h419: dout  = 8'b00000000; // 1049 :   0 - 0x0
      13'h41A: dout  = 8'b00000000; // 1050 :   0 - 0x0
      13'h41B: dout  = 8'b00000000; // 1051 :   0 - 0x0
      13'h41C: dout  = 8'b00000000; // 1052 :   0 - 0x0
      13'h41D: dout  = 8'b00000000; // 1053 :   0 - 0x0
      13'h41E: dout  = 8'b00000000; // 1054 :   0 - 0x0
      13'h41F: dout  = 8'b00000000; // 1055 :   0 - 0x0
      13'h420: dout  = 8'b00000000; // 1056 :   0 - 0x0 -- Sprite 0x42
      13'h421: dout  = 8'b00000000; // 1057 :   0 - 0x0
      13'h422: dout  = 8'b00000000; // 1058 :   0 - 0x0
      13'h423: dout  = 8'b00000000; // 1059 :   0 - 0x0
      13'h424: dout  = 8'b00000000; // 1060 :   0 - 0x0
      13'h425: dout  = 8'b00000000; // 1061 :   0 - 0x0
      13'h426: dout  = 8'b00000000; // 1062 :   0 - 0x0
      13'h427: dout  = 8'b00000000; // 1063 :   0 - 0x0
      13'h428: dout  = 8'b00000000; // 1064 :   0 - 0x0
      13'h429: dout  = 8'b00000000; // 1065 :   0 - 0x0
      13'h42A: dout  = 8'b00000000; // 1066 :   0 - 0x0
      13'h42B: dout  = 8'b00000000; // 1067 :   0 - 0x0
      13'h42C: dout  = 8'b00000000; // 1068 :   0 - 0x0
      13'h42D: dout  = 8'b00000000; // 1069 :   0 - 0x0
      13'h42E: dout  = 8'b00000000; // 1070 :   0 - 0x0
      13'h42F: dout  = 8'b00000000; // 1071 :   0 - 0x0
      13'h430: dout  = 8'b00000000; // 1072 :   0 - 0x0 -- Sprite 0x43
      13'h431: dout  = 8'b00000000; // 1073 :   0 - 0x0
      13'h432: dout  = 8'b00000000; // 1074 :   0 - 0x0
      13'h433: dout  = 8'b00000000; // 1075 :   0 - 0x0
      13'h434: dout  = 8'b00000000; // 1076 :   0 - 0x0
      13'h435: dout  = 8'b00000000; // 1077 :   0 - 0x0
      13'h436: dout  = 8'b00000000; // 1078 :   0 - 0x0
      13'h437: dout  = 8'b00000000; // 1079 :   0 - 0x0
      13'h438: dout  = 8'b00000000; // 1080 :   0 - 0x0
      13'h439: dout  = 8'b00000000; // 1081 :   0 - 0x0
      13'h43A: dout  = 8'b00000000; // 1082 :   0 - 0x0
      13'h43B: dout  = 8'b00000000; // 1083 :   0 - 0x0
      13'h43C: dout  = 8'b00000000; // 1084 :   0 - 0x0
      13'h43D: dout  = 8'b00000000; // 1085 :   0 - 0x0
      13'h43E: dout  = 8'b00000000; // 1086 :   0 - 0x0
      13'h43F: dout  = 8'b00000000; // 1087 :   0 - 0x0
      13'h440: dout  = 8'b00000000; // 1088 :   0 - 0x0 -- Sprite 0x44
      13'h441: dout  = 8'b00000000; // 1089 :   0 - 0x0
      13'h442: dout  = 8'b00000000; // 1090 :   0 - 0x0
      13'h443: dout  = 8'b00000000; // 1091 :   0 - 0x0
      13'h444: dout  = 8'b00000000; // 1092 :   0 - 0x0
      13'h445: dout  = 8'b00000000; // 1093 :   0 - 0x0
      13'h446: dout  = 8'b00000000; // 1094 :   0 - 0x0
      13'h447: dout  = 8'b00000000; // 1095 :   0 - 0x0
      13'h448: dout  = 8'b00000000; // 1096 :   0 - 0x0
      13'h449: dout  = 8'b00000000; // 1097 :   0 - 0x0
      13'h44A: dout  = 8'b00000000; // 1098 :   0 - 0x0
      13'h44B: dout  = 8'b00000000; // 1099 :   0 - 0x0
      13'h44C: dout  = 8'b00000000; // 1100 :   0 - 0x0
      13'h44D: dout  = 8'b00000000; // 1101 :   0 - 0x0
      13'h44E: dout  = 8'b00000000; // 1102 :   0 - 0x0
      13'h44F: dout  = 8'b00000000; // 1103 :   0 - 0x0
      13'h450: dout  = 8'b00000000; // 1104 :   0 - 0x0 -- Sprite 0x45
      13'h451: dout  = 8'b00000000; // 1105 :   0 - 0x0
      13'h452: dout  = 8'b00000000; // 1106 :   0 - 0x0
      13'h453: dout  = 8'b00000000; // 1107 :   0 - 0x0
      13'h454: dout  = 8'b00000000; // 1108 :   0 - 0x0
      13'h455: dout  = 8'b00000000; // 1109 :   0 - 0x0
      13'h456: dout  = 8'b00000000; // 1110 :   0 - 0x0
      13'h457: dout  = 8'b00000000; // 1111 :   0 - 0x0
      13'h458: dout  = 8'b00000000; // 1112 :   0 - 0x0
      13'h459: dout  = 8'b00000000; // 1113 :   0 - 0x0
      13'h45A: dout  = 8'b00000000; // 1114 :   0 - 0x0
      13'h45B: dout  = 8'b00000000; // 1115 :   0 - 0x0
      13'h45C: dout  = 8'b00000000; // 1116 :   0 - 0x0
      13'h45D: dout  = 8'b00000000; // 1117 :   0 - 0x0
      13'h45E: dout  = 8'b00000000; // 1118 :   0 - 0x0
      13'h45F: dout  = 8'b00000000; // 1119 :   0 - 0x0
      13'h460: dout  = 8'b00000000; // 1120 :   0 - 0x0 -- Sprite 0x46
      13'h461: dout  = 8'b00000000; // 1121 :   0 - 0x0
      13'h462: dout  = 8'b00000000; // 1122 :   0 - 0x0
      13'h463: dout  = 8'b00000000; // 1123 :   0 - 0x0
      13'h464: dout  = 8'b00000000; // 1124 :   0 - 0x0
      13'h465: dout  = 8'b00000000; // 1125 :   0 - 0x0
      13'h466: dout  = 8'b00000000; // 1126 :   0 - 0x0
      13'h467: dout  = 8'b00000000; // 1127 :   0 - 0x0
      13'h468: dout  = 8'b00000000; // 1128 :   0 - 0x0
      13'h469: dout  = 8'b00000000; // 1129 :   0 - 0x0
      13'h46A: dout  = 8'b00000000; // 1130 :   0 - 0x0
      13'h46B: dout  = 8'b00000000; // 1131 :   0 - 0x0
      13'h46C: dout  = 8'b00000000; // 1132 :   0 - 0x0
      13'h46D: dout  = 8'b00000000; // 1133 :   0 - 0x0
      13'h46E: dout  = 8'b00000000; // 1134 :   0 - 0x0
      13'h46F: dout  = 8'b00000000; // 1135 :   0 - 0x0
      13'h470: dout  = 8'b00000000; // 1136 :   0 - 0x0 -- Sprite 0x47
      13'h471: dout  = 8'b00000000; // 1137 :   0 - 0x0
      13'h472: dout  = 8'b00000000; // 1138 :   0 - 0x0
      13'h473: dout  = 8'b00000000; // 1139 :   0 - 0x0
      13'h474: dout  = 8'b00000000; // 1140 :   0 - 0x0
      13'h475: dout  = 8'b00000000; // 1141 :   0 - 0x0
      13'h476: dout  = 8'b00000000; // 1142 :   0 - 0x0
      13'h477: dout  = 8'b00000000; // 1143 :   0 - 0x0
      13'h478: dout  = 8'b00000000; // 1144 :   0 - 0x0
      13'h479: dout  = 8'b00000000; // 1145 :   0 - 0x0
      13'h47A: dout  = 8'b00000000; // 1146 :   0 - 0x0
      13'h47B: dout  = 8'b00000000; // 1147 :   0 - 0x0
      13'h47C: dout  = 8'b00000000; // 1148 :   0 - 0x0
      13'h47D: dout  = 8'b00000000; // 1149 :   0 - 0x0
      13'h47E: dout  = 8'b00000000; // 1150 :   0 - 0x0
      13'h47F: dout  = 8'b00000000; // 1151 :   0 - 0x0
      13'h480: dout  = 8'b00000000; // 1152 :   0 - 0x0 -- Sprite 0x48
      13'h481: dout  = 8'b00000000; // 1153 :   0 - 0x0
      13'h482: dout  = 8'b00000000; // 1154 :   0 - 0x0
      13'h483: dout  = 8'b00000000; // 1155 :   0 - 0x0
      13'h484: dout  = 8'b00000000; // 1156 :   0 - 0x0
      13'h485: dout  = 8'b00000000; // 1157 :   0 - 0x0
      13'h486: dout  = 8'b00000000; // 1158 :   0 - 0x0
      13'h487: dout  = 8'b00000000; // 1159 :   0 - 0x0
      13'h488: dout  = 8'b00000000; // 1160 :   0 - 0x0
      13'h489: dout  = 8'b00000000; // 1161 :   0 - 0x0
      13'h48A: dout  = 8'b00000000; // 1162 :   0 - 0x0
      13'h48B: dout  = 8'b00000000; // 1163 :   0 - 0x0
      13'h48C: dout  = 8'b00000000; // 1164 :   0 - 0x0
      13'h48D: dout  = 8'b00000000; // 1165 :   0 - 0x0
      13'h48E: dout  = 8'b00000000; // 1166 :   0 - 0x0
      13'h48F: dout  = 8'b00000000; // 1167 :   0 - 0x0
      13'h490: dout  = 8'b00000000; // 1168 :   0 - 0x0 -- Sprite 0x49
      13'h491: dout  = 8'b00000000; // 1169 :   0 - 0x0
      13'h492: dout  = 8'b00000000; // 1170 :   0 - 0x0
      13'h493: dout  = 8'b00000000; // 1171 :   0 - 0x0
      13'h494: dout  = 8'b00000000; // 1172 :   0 - 0x0
      13'h495: dout  = 8'b00000000; // 1173 :   0 - 0x0
      13'h496: dout  = 8'b00000000; // 1174 :   0 - 0x0
      13'h497: dout  = 8'b00000000; // 1175 :   0 - 0x0
      13'h498: dout  = 8'b00000000; // 1176 :   0 - 0x0
      13'h499: dout  = 8'b00000000; // 1177 :   0 - 0x0
      13'h49A: dout  = 8'b00000000; // 1178 :   0 - 0x0
      13'h49B: dout  = 8'b00000000; // 1179 :   0 - 0x0
      13'h49C: dout  = 8'b00000000; // 1180 :   0 - 0x0
      13'h49D: dout  = 8'b00000000; // 1181 :   0 - 0x0
      13'h49E: dout  = 8'b00000000; // 1182 :   0 - 0x0
      13'h49F: dout  = 8'b00000000; // 1183 :   0 - 0x0
      13'h4A0: dout  = 8'b00000000; // 1184 :   0 - 0x0 -- Sprite 0x4a
      13'h4A1: dout  = 8'b00000000; // 1185 :   0 - 0x0
      13'h4A2: dout  = 8'b00000000; // 1186 :   0 - 0x0
      13'h4A3: dout  = 8'b00000000; // 1187 :   0 - 0x0
      13'h4A4: dout  = 8'b00000000; // 1188 :   0 - 0x0
      13'h4A5: dout  = 8'b00000000; // 1189 :   0 - 0x0
      13'h4A6: dout  = 8'b00000000; // 1190 :   0 - 0x0
      13'h4A7: dout  = 8'b00000000; // 1191 :   0 - 0x0
      13'h4A8: dout  = 8'b00000000; // 1192 :   0 - 0x0
      13'h4A9: dout  = 8'b00000000; // 1193 :   0 - 0x0
      13'h4AA: dout  = 8'b00000000; // 1194 :   0 - 0x0
      13'h4AB: dout  = 8'b00000000; // 1195 :   0 - 0x0
      13'h4AC: dout  = 8'b00000000; // 1196 :   0 - 0x0
      13'h4AD: dout  = 8'b00000000; // 1197 :   0 - 0x0
      13'h4AE: dout  = 8'b00000000; // 1198 :   0 - 0x0
      13'h4AF: dout  = 8'b00000000; // 1199 :   0 - 0x0
      13'h4B0: dout  = 8'b00000000; // 1200 :   0 - 0x0 -- Sprite 0x4b
      13'h4B1: dout  = 8'b00000000; // 1201 :   0 - 0x0
      13'h4B2: dout  = 8'b00000000; // 1202 :   0 - 0x0
      13'h4B3: dout  = 8'b00000000; // 1203 :   0 - 0x0
      13'h4B4: dout  = 8'b00000000; // 1204 :   0 - 0x0
      13'h4B5: dout  = 8'b00000000; // 1205 :   0 - 0x0
      13'h4B6: dout  = 8'b00000000; // 1206 :   0 - 0x0
      13'h4B7: dout  = 8'b00000000; // 1207 :   0 - 0x0
      13'h4B8: dout  = 8'b00000000; // 1208 :   0 - 0x0
      13'h4B9: dout  = 8'b00000000; // 1209 :   0 - 0x0
      13'h4BA: dout  = 8'b00000000; // 1210 :   0 - 0x0
      13'h4BB: dout  = 8'b00000000; // 1211 :   0 - 0x0
      13'h4BC: dout  = 8'b00000000; // 1212 :   0 - 0x0
      13'h4BD: dout  = 8'b00000000; // 1213 :   0 - 0x0
      13'h4BE: dout  = 8'b00000000; // 1214 :   0 - 0x0
      13'h4BF: dout  = 8'b00000000; // 1215 :   0 - 0x0
      13'h4C0: dout  = 8'b00000000; // 1216 :   0 - 0x0 -- Sprite 0x4c
      13'h4C1: dout  = 8'b00000000; // 1217 :   0 - 0x0
      13'h4C2: dout  = 8'b00000000; // 1218 :   0 - 0x0
      13'h4C3: dout  = 8'b00000000; // 1219 :   0 - 0x0
      13'h4C4: dout  = 8'b00000000; // 1220 :   0 - 0x0
      13'h4C5: dout  = 8'b00000000; // 1221 :   0 - 0x0
      13'h4C6: dout  = 8'b00000000; // 1222 :   0 - 0x0
      13'h4C7: dout  = 8'b00000000; // 1223 :   0 - 0x0
      13'h4C8: dout  = 8'b00000000; // 1224 :   0 - 0x0
      13'h4C9: dout  = 8'b00000000; // 1225 :   0 - 0x0
      13'h4CA: dout  = 8'b00000000; // 1226 :   0 - 0x0
      13'h4CB: dout  = 8'b00000000; // 1227 :   0 - 0x0
      13'h4CC: dout  = 8'b00000000; // 1228 :   0 - 0x0
      13'h4CD: dout  = 8'b00000000; // 1229 :   0 - 0x0
      13'h4CE: dout  = 8'b00000000; // 1230 :   0 - 0x0
      13'h4CF: dout  = 8'b00000000; // 1231 :   0 - 0x0
      13'h4D0: dout  = 8'b00000000; // 1232 :   0 - 0x0 -- Sprite 0x4d
      13'h4D1: dout  = 8'b00000000; // 1233 :   0 - 0x0
      13'h4D2: dout  = 8'b00000000; // 1234 :   0 - 0x0
      13'h4D3: dout  = 8'b00000000; // 1235 :   0 - 0x0
      13'h4D4: dout  = 8'b00000000; // 1236 :   0 - 0x0
      13'h4D5: dout  = 8'b00000000; // 1237 :   0 - 0x0
      13'h4D6: dout  = 8'b00000000; // 1238 :   0 - 0x0
      13'h4D7: dout  = 8'b00000000; // 1239 :   0 - 0x0
      13'h4D8: dout  = 8'b00000000; // 1240 :   0 - 0x0
      13'h4D9: dout  = 8'b00000000; // 1241 :   0 - 0x0
      13'h4DA: dout  = 8'b00000000; // 1242 :   0 - 0x0
      13'h4DB: dout  = 8'b00000000; // 1243 :   0 - 0x0
      13'h4DC: dout  = 8'b00000000; // 1244 :   0 - 0x0
      13'h4DD: dout  = 8'b00000000; // 1245 :   0 - 0x0
      13'h4DE: dout  = 8'b00000000; // 1246 :   0 - 0x0
      13'h4DF: dout  = 8'b00000000; // 1247 :   0 - 0x0
      13'h4E0: dout  = 8'b00000000; // 1248 :   0 - 0x0 -- Sprite 0x4e
      13'h4E1: dout  = 8'b00000000; // 1249 :   0 - 0x0
      13'h4E2: dout  = 8'b00000000; // 1250 :   0 - 0x0
      13'h4E3: dout  = 8'b00000000; // 1251 :   0 - 0x0
      13'h4E4: dout  = 8'b00000000; // 1252 :   0 - 0x0
      13'h4E5: dout  = 8'b00000000; // 1253 :   0 - 0x0
      13'h4E6: dout  = 8'b00000000; // 1254 :   0 - 0x0
      13'h4E7: dout  = 8'b00000000; // 1255 :   0 - 0x0
      13'h4E8: dout  = 8'b00000000; // 1256 :   0 - 0x0
      13'h4E9: dout  = 8'b00000000; // 1257 :   0 - 0x0
      13'h4EA: dout  = 8'b00000000; // 1258 :   0 - 0x0
      13'h4EB: dout  = 8'b00000000; // 1259 :   0 - 0x0
      13'h4EC: dout  = 8'b00000000; // 1260 :   0 - 0x0
      13'h4ED: dout  = 8'b00000000; // 1261 :   0 - 0x0
      13'h4EE: dout  = 8'b00000000; // 1262 :   0 - 0x0
      13'h4EF: dout  = 8'b00000000; // 1263 :   0 - 0x0
      13'h4F0: dout  = 8'b00000000; // 1264 :   0 - 0x0 -- Sprite 0x4f
      13'h4F1: dout  = 8'b00000000; // 1265 :   0 - 0x0
      13'h4F2: dout  = 8'b00000000; // 1266 :   0 - 0x0
      13'h4F3: dout  = 8'b00000000; // 1267 :   0 - 0x0
      13'h4F4: dout  = 8'b00000000; // 1268 :   0 - 0x0
      13'h4F5: dout  = 8'b00000000; // 1269 :   0 - 0x0
      13'h4F6: dout  = 8'b00000000; // 1270 :   0 - 0x0
      13'h4F7: dout  = 8'b00000000; // 1271 :   0 - 0x0
      13'h4F8: dout  = 8'b00000000; // 1272 :   0 - 0x0
      13'h4F9: dout  = 8'b00000000; // 1273 :   0 - 0x0
      13'h4FA: dout  = 8'b00000000; // 1274 :   0 - 0x0
      13'h4FB: dout  = 8'b00000000; // 1275 :   0 - 0x0
      13'h4FC: dout  = 8'b00000000; // 1276 :   0 - 0x0
      13'h4FD: dout  = 8'b00000000; // 1277 :   0 - 0x0
      13'h4FE: dout  = 8'b00000000; // 1278 :   0 - 0x0
      13'h4FF: dout  = 8'b00000000; // 1279 :   0 - 0x0
      13'h500: dout  = 8'b00000000; // 1280 :   0 - 0x0 -- Sprite 0x50
      13'h501: dout  = 8'b00000000; // 1281 :   0 - 0x0
      13'h502: dout  = 8'b00000000; // 1282 :   0 - 0x0
      13'h503: dout  = 8'b00000000; // 1283 :   0 - 0x0
      13'h504: dout  = 8'b00000000; // 1284 :   0 - 0x0
      13'h505: dout  = 8'b00000000; // 1285 :   0 - 0x0
      13'h506: dout  = 8'b00000000; // 1286 :   0 - 0x0
      13'h507: dout  = 8'b00000000; // 1287 :   0 - 0x0
      13'h508: dout  = 8'b00000000; // 1288 :   0 - 0x0
      13'h509: dout  = 8'b00000000; // 1289 :   0 - 0x0
      13'h50A: dout  = 8'b00000000; // 1290 :   0 - 0x0
      13'h50B: dout  = 8'b00000000; // 1291 :   0 - 0x0
      13'h50C: dout  = 8'b00000000; // 1292 :   0 - 0x0
      13'h50D: dout  = 8'b00000000; // 1293 :   0 - 0x0
      13'h50E: dout  = 8'b00000000; // 1294 :   0 - 0x0
      13'h50F: dout  = 8'b00000000; // 1295 :   0 - 0x0
      13'h510: dout  = 8'b00000000; // 1296 :   0 - 0x0 -- Sprite 0x51
      13'h511: dout  = 8'b00000000; // 1297 :   0 - 0x0
      13'h512: dout  = 8'b00000000; // 1298 :   0 - 0x0
      13'h513: dout  = 8'b00000000; // 1299 :   0 - 0x0
      13'h514: dout  = 8'b00000000; // 1300 :   0 - 0x0
      13'h515: dout  = 8'b00000000; // 1301 :   0 - 0x0
      13'h516: dout  = 8'b00000000; // 1302 :   0 - 0x0
      13'h517: dout  = 8'b00000000; // 1303 :   0 - 0x0
      13'h518: dout  = 8'b00000000; // 1304 :   0 - 0x0
      13'h519: dout  = 8'b00000000; // 1305 :   0 - 0x0
      13'h51A: dout  = 8'b00000000; // 1306 :   0 - 0x0
      13'h51B: dout  = 8'b00000000; // 1307 :   0 - 0x0
      13'h51C: dout  = 8'b00000000; // 1308 :   0 - 0x0
      13'h51D: dout  = 8'b00000000; // 1309 :   0 - 0x0
      13'h51E: dout  = 8'b00000000; // 1310 :   0 - 0x0
      13'h51F: dout  = 8'b00000000; // 1311 :   0 - 0x0
      13'h520: dout  = 8'b00000000; // 1312 :   0 - 0x0 -- Sprite 0x52
      13'h521: dout  = 8'b00000000; // 1313 :   0 - 0x0
      13'h522: dout  = 8'b00000000; // 1314 :   0 - 0x0
      13'h523: dout  = 8'b00000000; // 1315 :   0 - 0x0
      13'h524: dout  = 8'b00000000; // 1316 :   0 - 0x0
      13'h525: dout  = 8'b00000000; // 1317 :   0 - 0x0
      13'h526: dout  = 8'b00000000; // 1318 :   0 - 0x0
      13'h527: dout  = 8'b00000000; // 1319 :   0 - 0x0
      13'h528: dout  = 8'b00000000; // 1320 :   0 - 0x0
      13'h529: dout  = 8'b00000000; // 1321 :   0 - 0x0
      13'h52A: dout  = 8'b00000000; // 1322 :   0 - 0x0
      13'h52B: dout  = 8'b00000000; // 1323 :   0 - 0x0
      13'h52C: dout  = 8'b00000000; // 1324 :   0 - 0x0
      13'h52D: dout  = 8'b00000000; // 1325 :   0 - 0x0
      13'h52E: dout  = 8'b00000000; // 1326 :   0 - 0x0
      13'h52F: dout  = 8'b00000000; // 1327 :   0 - 0x0
      13'h530: dout  = 8'b00000000; // 1328 :   0 - 0x0 -- Sprite 0x53
      13'h531: dout  = 8'b00000000; // 1329 :   0 - 0x0
      13'h532: dout  = 8'b00000000; // 1330 :   0 - 0x0
      13'h533: dout  = 8'b00000000; // 1331 :   0 - 0x0
      13'h534: dout  = 8'b00000000; // 1332 :   0 - 0x0
      13'h535: dout  = 8'b00000000; // 1333 :   0 - 0x0
      13'h536: dout  = 8'b00000000; // 1334 :   0 - 0x0
      13'h537: dout  = 8'b00000000; // 1335 :   0 - 0x0
      13'h538: dout  = 8'b00000000; // 1336 :   0 - 0x0
      13'h539: dout  = 8'b00000000; // 1337 :   0 - 0x0
      13'h53A: dout  = 8'b00000000; // 1338 :   0 - 0x0
      13'h53B: dout  = 8'b00000000; // 1339 :   0 - 0x0
      13'h53C: dout  = 8'b00000000; // 1340 :   0 - 0x0
      13'h53D: dout  = 8'b00000000; // 1341 :   0 - 0x0
      13'h53E: dout  = 8'b00000000; // 1342 :   0 - 0x0
      13'h53F: dout  = 8'b00000000; // 1343 :   0 - 0x0
      13'h540: dout  = 8'b00000000; // 1344 :   0 - 0x0 -- Sprite 0x54
      13'h541: dout  = 8'b00000000; // 1345 :   0 - 0x0
      13'h542: dout  = 8'b00000000; // 1346 :   0 - 0x0
      13'h543: dout  = 8'b00000000; // 1347 :   0 - 0x0
      13'h544: dout  = 8'b00000000; // 1348 :   0 - 0x0
      13'h545: dout  = 8'b00000000; // 1349 :   0 - 0x0
      13'h546: dout  = 8'b00000000; // 1350 :   0 - 0x0
      13'h547: dout  = 8'b00000000; // 1351 :   0 - 0x0
      13'h548: dout  = 8'b00000000; // 1352 :   0 - 0x0
      13'h549: dout  = 8'b00000000; // 1353 :   0 - 0x0
      13'h54A: dout  = 8'b00000000; // 1354 :   0 - 0x0
      13'h54B: dout  = 8'b00000000; // 1355 :   0 - 0x0
      13'h54C: dout  = 8'b00000000; // 1356 :   0 - 0x0
      13'h54D: dout  = 8'b00000000; // 1357 :   0 - 0x0
      13'h54E: dout  = 8'b00000000; // 1358 :   0 - 0x0
      13'h54F: dout  = 8'b00000000; // 1359 :   0 - 0x0
      13'h550: dout  = 8'b00000000; // 1360 :   0 - 0x0 -- Sprite 0x55
      13'h551: dout  = 8'b00000000; // 1361 :   0 - 0x0
      13'h552: dout  = 8'b00000000; // 1362 :   0 - 0x0
      13'h553: dout  = 8'b00000000; // 1363 :   0 - 0x0
      13'h554: dout  = 8'b00000000; // 1364 :   0 - 0x0
      13'h555: dout  = 8'b00000000; // 1365 :   0 - 0x0
      13'h556: dout  = 8'b00000000; // 1366 :   0 - 0x0
      13'h557: dout  = 8'b00000000; // 1367 :   0 - 0x0
      13'h558: dout  = 8'b00000000; // 1368 :   0 - 0x0
      13'h559: dout  = 8'b00000000; // 1369 :   0 - 0x0
      13'h55A: dout  = 8'b00000000; // 1370 :   0 - 0x0
      13'h55B: dout  = 8'b00000000; // 1371 :   0 - 0x0
      13'h55C: dout  = 8'b00000000; // 1372 :   0 - 0x0
      13'h55D: dout  = 8'b00000000; // 1373 :   0 - 0x0
      13'h55E: dout  = 8'b00000000; // 1374 :   0 - 0x0
      13'h55F: dout  = 8'b00000000; // 1375 :   0 - 0x0
      13'h560: dout  = 8'b00000000; // 1376 :   0 - 0x0 -- Sprite 0x56
      13'h561: dout  = 8'b00000000; // 1377 :   0 - 0x0
      13'h562: dout  = 8'b00000000; // 1378 :   0 - 0x0
      13'h563: dout  = 8'b00000000; // 1379 :   0 - 0x0
      13'h564: dout  = 8'b00000000; // 1380 :   0 - 0x0
      13'h565: dout  = 8'b00000000; // 1381 :   0 - 0x0
      13'h566: dout  = 8'b00000000; // 1382 :   0 - 0x0
      13'h567: dout  = 8'b00000000; // 1383 :   0 - 0x0
      13'h568: dout  = 8'b00000000; // 1384 :   0 - 0x0
      13'h569: dout  = 8'b00000000; // 1385 :   0 - 0x0
      13'h56A: dout  = 8'b00000000; // 1386 :   0 - 0x0
      13'h56B: dout  = 8'b00000000; // 1387 :   0 - 0x0
      13'h56C: dout  = 8'b00000000; // 1388 :   0 - 0x0
      13'h56D: dout  = 8'b00000000; // 1389 :   0 - 0x0
      13'h56E: dout  = 8'b00000000; // 1390 :   0 - 0x0
      13'h56F: dout  = 8'b00000000; // 1391 :   0 - 0x0
      13'h570: dout  = 8'b00000000; // 1392 :   0 - 0x0 -- Sprite 0x57
      13'h571: dout  = 8'b00000000; // 1393 :   0 - 0x0
      13'h572: dout  = 8'b00000000; // 1394 :   0 - 0x0
      13'h573: dout  = 8'b00000000; // 1395 :   0 - 0x0
      13'h574: dout  = 8'b00000000; // 1396 :   0 - 0x0
      13'h575: dout  = 8'b00000000; // 1397 :   0 - 0x0
      13'h576: dout  = 8'b00000000; // 1398 :   0 - 0x0
      13'h577: dout  = 8'b00000000; // 1399 :   0 - 0x0
      13'h578: dout  = 8'b00000000; // 1400 :   0 - 0x0
      13'h579: dout  = 8'b00000000; // 1401 :   0 - 0x0
      13'h57A: dout  = 8'b00000000; // 1402 :   0 - 0x0
      13'h57B: dout  = 8'b00000000; // 1403 :   0 - 0x0
      13'h57C: dout  = 8'b00000000; // 1404 :   0 - 0x0
      13'h57D: dout  = 8'b00000000; // 1405 :   0 - 0x0
      13'h57E: dout  = 8'b00000000; // 1406 :   0 - 0x0
      13'h57F: dout  = 8'b00000000; // 1407 :   0 - 0x0
      13'h580: dout  = 8'b00000000; // 1408 :   0 - 0x0 -- Sprite 0x58
      13'h581: dout  = 8'b00000000; // 1409 :   0 - 0x0
      13'h582: dout  = 8'b00000000; // 1410 :   0 - 0x0
      13'h583: dout  = 8'b00000000; // 1411 :   0 - 0x0
      13'h584: dout  = 8'b00000000; // 1412 :   0 - 0x0
      13'h585: dout  = 8'b00000000; // 1413 :   0 - 0x0
      13'h586: dout  = 8'b00000000; // 1414 :   0 - 0x0
      13'h587: dout  = 8'b00000000; // 1415 :   0 - 0x0
      13'h588: dout  = 8'b00000000; // 1416 :   0 - 0x0
      13'h589: dout  = 8'b00000000; // 1417 :   0 - 0x0
      13'h58A: dout  = 8'b00000000; // 1418 :   0 - 0x0
      13'h58B: dout  = 8'b00000000; // 1419 :   0 - 0x0
      13'h58C: dout  = 8'b00000000; // 1420 :   0 - 0x0
      13'h58D: dout  = 8'b00000000; // 1421 :   0 - 0x0
      13'h58E: dout  = 8'b00000000; // 1422 :   0 - 0x0
      13'h58F: dout  = 8'b00000000; // 1423 :   0 - 0x0
      13'h590: dout  = 8'b00000000; // 1424 :   0 - 0x0 -- Sprite 0x59
      13'h591: dout  = 8'b00000000; // 1425 :   0 - 0x0
      13'h592: dout  = 8'b00000000; // 1426 :   0 - 0x0
      13'h593: dout  = 8'b00000000; // 1427 :   0 - 0x0
      13'h594: dout  = 8'b00000000; // 1428 :   0 - 0x0
      13'h595: dout  = 8'b00000000; // 1429 :   0 - 0x0
      13'h596: dout  = 8'b00000000; // 1430 :   0 - 0x0
      13'h597: dout  = 8'b00000000; // 1431 :   0 - 0x0
      13'h598: dout  = 8'b00000000; // 1432 :   0 - 0x0
      13'h599: dout  = 8'b00000000; // 1433 :   0 - 0x0
      13'h59A: dout  = 8'b00000000; // 1434 :   0 - 0x0
      13'h59B: dout  = 8'b00000000; // 1435 :   0 - 0x0
      13'h59C: dout  = 8'b00000000; // 1436 :   0 - 0x0
      13'h59D: dout  = 8'b00000000; // 1437 :   0 - 0x0
      13'h59E: dout  = 8'b00000000; // 1438 :   0 - 0x0
      13'h59F: dout  = 8'b00000000; // 1439 :   0 - 0x0
      13'h5A0: dout  = 8'b00000000; // 1440 :   0 - 0x0 -- Sprite 0x5a
      13'h5A1: dout  = 8'b00000000; // 1441 :   0 - 0x0
      13'h5A2: dout  = 8'b00000000; // 1442 :   0 - 0x0
      13'h5A3: dout  = 8'b00000000; // 1443 :   0 - 0x0
      13'h5A4: dout  = 8'b00000000; // 1444 :   0 - 0x0
      13'h5A5: dout  = 8'b00000000; // 1445 :   0 - 0x0
      13'h5A6: dout  = 8'b00000000; // 1446 :   0 - 0x0
      13'h5A7: dout  = 8'b00000000; // 1447 :   0 - 0x0
      13'h5A8: dout  = 8'b00000000; // 1448 :   0 - 0x0
      13'h5A9: dout  = 8'b00000000; // 1449 :   0 - 0x0
      13'h5AA: dout  = 8'b00000000; // 1450 :   0 - 0x0
      13'h5AB: dout  = 8'b00000000; // 1451 :   0 - 0x0
      13'h5AC: dout  = 8'b00000000; // 1452 :   0 - 0x0
      13'h5AD: dout  = 8'b00000000; // 1453 :   0 - 0x0
      13'h5AE: dout  = 8'b00000000; // 1454 :   0 - 0x0
      13'h5AF: dout  = 8'b00000000; // 1455 :   0 - 0x0
      13'h5B0: dout  = 8'b00000000; // 1456 :   0 - 0x0 -- Sprite 0x5b
      13'h5B1: dout  = 8'b00000000; // 1457 :   0 - 0x0
      13'h5B2: dout  = 8'b00000000; // 1458 :   0 - 0x0
      13'h5B3: dout  = 8'b00000000; // 1459 :   0 - 0x0
      13'h5B4: dout  = 8'b00000000; // 1460 :   0 - 0x0
      13'h5B5: dout  = 8'b00000000; // 1461 :   0 - 0x0
      13'h5B6: dout  = 8'b00000000; // 1462 :   0 - 0x0
      13'h5B7: dout  = 8'b00000000; // 1463 :   0 - 0x0
      13'h5B8: dout  = 8'b00000000; // 1464 :   0 - 0x0
      13'h5B9: dout  = 8'b00000000; // 1465 :   0 - 0x0
      13'h5BA: dout  = 8'b00000000; // 1466 :   0 - 0x0
      13'h5BB: dout  = 8'b00000000; // 1467 :   0 - 0x0
      13'h5BC: dout  = 8'b00000000; // 1468 :   0 - 0x0
      13'h5BD: dout  = 8'b00000000; // 1469 :   0 - 0x0
      13'h5BE: dout  = 8'b00000000; // 1470 :   0 - 0x0
      13'h5BF: dout  = 8'b00000000; // 1471 :   0 - 0x0
      13'h5C0: dout  = 8'b00000000; // 1472 :   0 - 0x0 -- Sprite 0x5c
      13'h5C1: dout  = 8'b00000000; // 1473 :   0 - 0x0
      13'h5C2: dout  = 8'b00000000; // 1474 :   0 - 0x0
      13'h5C3: dout  = 8'b00000000; // 1475 :   0 - 0x0
      13'h5C4: dout  = 8'b00000000; // 1476 :   0 - 0x0
      13'h5C5: dout  = 8'b00000000; // 1477 :   0 - 0x0
      13'h5C6: dout  = 8'b00000000; // 1478 :   0 - 0x0
      13'h5C7: dout  = 8'b00000000; // 1479 :   0 - 0x0
      13'h5C8: dout  = 8'b00000000; // 1480 :   0 - 0x0
      13'h5C9: dout  = 8'b00000000; // 1481 :   0 - 0x0
      13'h5CA: dout  = 8'b00000000; // 1482 :   0 - 0x0
      13'h5CB: dout  = 8'b00000000; // 1483 :   0 - 0x0
      13'h5CC: dout  = 8'b00000000; // 1484 :   0 - 0x0
      13'h5CD: dout  = 8'b00000000; // 1485 :   0 - 0x0
      13'h5CE: dout  = 8'b00000000; // 1486 :   0 - 0x0
      13'h5CF: dout  = 8'b00000000; // 1487 :   0 - 0x0
      13'h5D0: dout  = 8'b00000000; // 1488 :   0 - 0x0 -- Sprite 0x5d
      13'h5D1: dout  = 8'b00000000; // 1489 :   0 - 0x0
      13'h5D2: dout  = 8'b00000000; // 1490 :   0 - 0x0
      13'h5D3: dout  = 8'b00000000; // 1491 :   0 - 0x0
      13'h5D4: dout  = 8'b00000000; // 1492 :   0 - 0x0
      13'h5D5: dout  = 8'b00000000; // 1493 :   0 - 0x0
      13'h5D6: dout  = 8'b00000000; // 1494 :   0 - 0x0
      13'h5D7: dout  = 8'b00000000; // 1495 :   0 - 0x0
      13'h5D8: dout  = 8'b00000000; // 1496 :   0 - 0x0
      13'h5D9: dout  = 8'b00000000; // 1497 :   0 - 0x0
      13'h5DA: dout  = 8'b00000000; // 1498 :   0 - 0x0
      13'h5DB: dout  = 8'b00000000; // 1499 :   0 - 0x0
      13'h5DC: dout  = 8'b00000000; // 1500 :   0 - 0x0
      13'h5DD: dout  = 8'b00000000; // 1501 :   0 - 0x0
      13'h5DE: dout  = 8'b00000000; // 1502 :   0 - 0x0
      13'h5DF: dout  = 8'b00000000; // 1503 :   0 - 0x0
      13'h5E0: dout  = 8'b00000000; // 1504 :   0 - 0x0 -- Sprite 0x5e
      13'h5E1: dout  = 8'b00000000; // 1505 :   0 - 0x0
      13'h5E2: dout  = 8'b00000000; // 1506 :   0 - 0x0
      13'h5E3: dout  = 8'b00000000; // 1507 :   0 - 0x0
      13'h5E4: dout  = 8'b00000000; // 1508 :   0 - 0x0
      13'h5E5: dout  = 8'b00000000; // 1509 :   0 - 0x0
      13'h5E6: dout  = 8'b00000000; // 1510 :   0 - 0x0
      13'h5E7: dout  = 8'b00000000; // 1511 :   0 - 0x0
      13'h5E8: dout  = 8'b00000000; // 1512 :   0 - 0x0
      13'h5E9: dout  = 8'b00000000; // 1513 :   0 - 0x0
      13'h5EA: dout  = 8'b00000000; // 1514 :   0 - 0x0
      13'h5EB: dout  = 8'b00000000; // 1515 :   0 - 0x0
      13'h5EC: dout  = 8'b00000000; // 1516 :   0 - 0x0
      13'h5ED: dout  = 8'b00000000; // 1517 :   0 - 0x0
      13'h5EE: dout  = 8'b00000000; // 1518 :   0 - 0x0
      13'h5EF: dout  = 8'b00000000; // 1519 :   0 - 0x0
      13'h5F0: dout  = 8'b00000000; // 1520 :   0 - 0x0 -- Sprite 0x5f
      13'h5F1: dout  = 8'b00000000; // 1521 :   0 - 0x0
      13'h5F2: dout  = 8'b00000000; // 1522 :   0 - 0x0
      13'h5F3: dout  = 8'b00000000; // 1523 :   0 - 0x0
      13'h5F4: dout  = 8'b00000000; // 1524 :   0 - 0x0
      13'h5F5: dout  = 8'b00000000; // 1525 :   0 - 0x0
      13'h5F6: dout  = 8'b00000000; // 1526 :   0 - 0x0
      13'h5F7: dout  = 8'b00000000; // 1527 :   0 - 0x0
      13'h5F8: dout  = 8'b00000000; // 1528 :   0 - 0x0
      13'h5F9: dout  = 8'b00000000; // 1529 :   0 - 0x0
      13'h5FA: dout  = 8'b00000000; // 1530 :   0 - 0x0
      13'h5FB: dout  = 8'b00000000; // 1531 :   0 - 0x0
      13'h5FC: dout  = 8'b00000000; // 1532 :   0 - 0x0
      13'h5FD: dout  = 8'b00000000; // 1533 :   0 - 0x0
      13'h5FE: dout  = 8'b00000000; // 1534 :   0 - 0x0
      13'h5FF: dout  = 8'b00000000; // 1535 :   0 - 0x0
      13'h600: dout  = 8'b00000000; // 1536 :   0 - 0x0 -- Sprite 0x60
      13'h601: dout  = 8'b00000000; // 1537 :   0 - 0x0
      13'h602: dout  = 8'b00000000; // 1538 :   0 - 0x0
      13'h603: dout  = 8'b00000000; // 1539 :   0 - 0x0
      13'h604: dout  = 8'b00000000; // 1540 :   0 - 0x0
      13'h605: dout  = 8'b00000000; // 1541 :   0 - 0x0
      13'h606: dout  = 8'b00000000; // 1542 :   0 - 0x0
      13'h607: dout  = 8'b00000000; // 1543 :   0 - 0x0
      13'h608: dout  = 8'b00000000; // 1544 :   0 - 0x0
      13'h609: dout  = 8'b00000000; // 1545 :   0 - 0x0
      13'h60A: dout  = 8'b00000000; // 1546 :   0 - 0x0
      13'h60B: dout  = 8'b00000000; // 1547 :   0 - 0x0
      13'h60C: dout  = 8'b00000000; // 1548 :   0 - 0x0
      13'h60D: dout  = 8'b00000000; // 1549 :   0 - 0x0
      13'h60E: dout  = 8'b00000000; // 1550 :   0 - 0x0
      13'h60F: dout  = 8'b00000000; // 1551 :   0 - 0x0
      13'h610: dout  = 8'b00000000; // 1552 :   0 - 0x0 -- Sprite 0x61
      13'h611: dout  = 8'b00000000; // 1553 :   0 - 0x0
      13'h612: dout  = 8'b00000000; // 1554 :   0 - 0x0
      13'h613: dout  = 8'b00000000; // 1555 :   0 - 0x0
      13'h614: dout  = 8'b00000000; // 1556 :   0 - 0x0
      13'h615: dout  = 8'b00000000; // 1557 :   0 - 0x0
      13'h616: dout  = 8'b00000000; // 1558 :   0 - 0x0
      13'h617: dout  = 8'b00000000; // 1559 :   0 - 0x0
      13'h618: dout  = 8'b00000000; // 1560 :   0 - 0x0
      13'h619: dout  = 8'b00000000; // 1561 :   0 - 0x0
      13'h61A: dout  = 8'b00000000; // 1562 :   0 - 0x0
      13'h61B: dout  = 8'b00000000; // 1563 :   0 - 0x0
      13'h61C: dout  = 8'b00000000; // 1564 :   0 - 0x0
      13'h61D: dout  = 8'b00000000; // 1565 :   0 - 0x0
      13'h61E: dout  = 8'b00000000; // 1566 :   0 - 0x0
      13'h61F: dout  = 8'b00000000; // 1567 :   0 - 0x0
      13'h620: dout  = 8'b00000000; // 1568 :   0 - 0x0 -- Sprite 0x62
      13'h621: dout  = 8'b00000000; // 1569 :   0 - 0x0
      13'h622: dout  = 8'b00000000; // 1570 :   0 - 0x0
      13'h623: dout  = 8'b00000000; // 1571 :   0 - 0x0
      13'h624: dout  = 8'b00000000; // 1572 :   0 - 0x0
      13'h625: dout  = 8'b00000000; // 1573 :   0 - 0x0
      13'h626: dout  = 8'b00000000; // 1574 :   0 - 0x0
      13'h627: dout  = 8'b00000000; // 1575 :   0 - 0x0
      13'h628: dout  = 8'b00000000; // 1576 :   0 - 0x0
      13'h629: dout  = 8'b00000000; // 1577 :   0 - 0x0
      13'h62A: dout  = 8'b00000000; // 1578 :   0 - 0x0
      13'h62B: dout  = 8'b00000000; // 1579 :   0 - 0x0
      13'h62C: dout  = 8'b00000000; // 1580 :   0 - 0x0
      13'h62D: dout  = 8'b00000000; // 1581 :   0 - 0x0
      13'h62E: dout  = 8'b00000000; // 1582 :   0 - 0x0
      13'h62F: dout  = 8'b00000000; // 1583 :   0 - 0x0
      13'h630: dout  = 8'b00000000; // 1584 :   0 - 0x0 -- Sprite 0x63
      13'h631: dout  = 8'b00000000; // 1585 :   0 - 0x0
      13'h632: dout  = 8'b00000000; // 1586 :   0 - 0x0
      13'h633: dout  = 8'b00000000; // 1587 :   0 - 0x0
      13'h634: dout  = 8'b00000000; // 1588 :   0 - 0x0
      13'h635: dout  = 8'b00000000; // 1589 :   0 - 0x0
      13'h636: dout  = 8'b00000000; // 1590 :   0 - 0x0
      13'h637: dout  = 8'b00000000; // 1591 :   0 - 0x0
      13'h638: dout  = 8'b00000000; // 1592 :   0 - 0x0
      13'h639: dout  = 8'b00000000; // 1593 :   0 - 0x0
      13'h63A: dout  = 8'b00000000; // 1594 :   0 - 0x0
      13'h63B: dout  = 8'b00000000; // 1595 :   0 - 0x0
      13'h63C: dout  = 8'b00000000; // 1596 :   0 - 0x0
      13'h63D: dout  = 8'b00000000; // 1597 :   0 - 0x0
      13'h63E: dout  = 8'b00000000; // 1598 :   0 - 0x0
      13'h63F: dout  = 8'b00000000; // 1599 :   0 - 0x0
      13'h640: dout  = 8'b00000000; // 1600 :   0 - 0x0 -- Sprite 0x64
      13'h641: dout  = 8'b00000000; // 1601 :   0 - 0x0
      13'h642: dout  = 8'b00000000; // 1602 :   0 - 0x0
      13'h643: dout  = 8'b00000000; // 1603 :   0 - 0x0
      13'h644: dout  = 8'b00000000; // 1604 :   0 - 0x0
      13'h645: dout  = 8'b00000000; // 1605 :   0 - 0x0
      13'h646: dout  = 8'b00000000; // 1606 :   0 - 0x0
      13'h647: dout  = 8'b00000000; // 1607 :   0 - 0x0
      13'h648: dout  = 8'b00000000; // 1608 :   0 - 0x0
      13'h649: dout  = 8'b00000000; // 1609 :   0 - 0x0
      13'h64A: dout  = 8'b00000000; // 1610 :   0 - 0x0
      13'h64B: dout  = 8'b00000000; // 1611 :   0 - 0x0
      13'h64C: dout  = 8'b00000000; // 1612 :   0 - 0x0
      13'h64D: dout  = 8'b00000000; // 1613 :   0 - 0x0
      13'h64E: dout  = 8'b00000000; // 1614 :   0 - 0x0
      13'h64F: dout  = 8'b00000000; // 1615 :   0 - 0x0
      13'h650: dout  = 8'b00000000; // 1616 :   0 - 0x0 -- Sprite 0x65
      13'h651: dout  = 8'b00000000; // 1617 :   0 - 0x0
      13'h652: dout  = 8'b00000000; // 1618 :   0 - 0x0
      13'h653: dout  = 8'b00000000; // 1619 :   0 - 0x0
      13'h654: dout  = 8'b00000000; // 1620 :   0 - 0x0
      13'h655: dout  = 8'b00000000; // 1621 :   0 - 0x0
      13'h656: dout  = 8'b00000000; // 1622 :   0 - 0x0
      13'h657: dout  = 8'b00000000; // 1623 :   0 - 0x0
      13'h658: dout  = 8'b00000000; // 1624 :   0 - 0x0
      13'h659: dout  = 8'b00000000; // 1625 :   0 - 0x0
      13'h65A: dout  = 8'b00000000; // 1626 :   0 - 0x0
      13'h65B: dout  = 8'b00000000; // 1627 :   0 - 0x0
      13'h65C: dout  = 8'b00000000; // 1628 :   0 - 0x0
      13'h65D: dout  = 8'b00000000; // 1629 :   0 - 0x0
      13'h65E: dout  = 8'b00000000; // 1630 :   0 - 0x0
      13'h65F: dout  = 8'b00000000; // 1631 :   0 - 0x0
      13'h660: dout  = 8'b00000000; // 1632 :   0 - 0x0 -- Sprite 0x66
      13'h661: dout  = 8'b00000000; // 1633 :   0 - 0x0
      13'h662: dout  = 8'b00000000; // 1634 :   0 - 0x0
      13'h663: dout  = 8'b00000000; // 1635 :   0 - 0x0
      13'h664: dout  = 8'b00000000; // 1636 :   0 - 0x0
      13'h665: dout  = 8'b00000000; // 1637 :   0 - 0x0
      13'h666: dout  = 8'b00000000; // 1638 :   0 - 0x0
      13'h667: dout  = 8'b00000000; // 1639 :   0 - 0x0
      13'h668: dout  = 8'b00000000; // 1640 :   0 - 0x0
      13'h669: dout  = 8'b00000000; // 1641 :   0 - 0x0
      13'h66A: dout  = 8'b00000000; // 1642 :   0 - 0x0
      13'h66B: dout  = 8'b00000000; // 1643 :   0 - 0x0
      13'h66C: dout  = 8'b00000000; // 1644 :   0 - 0x0
      13'h66D: dout  = 8'b00000000; // 1645 :   0 - 0x0
      13'h66E: dout  = 8'b00000000; // 1646 :   0 - 0x0
      13'h66F: dout  = 8'b00000000; // 1647 :   0 - 0x0
      13'h670: dout  = 8'b00000000; // 1648 :   0 - 0x0 -- Sprite 0x67
      13'h671: dout  = 8'b00000000; // 1649 :   0 - 0x0
      13'h672: dout  = 8'b00000000; // 1650 :   0 - 0x0
      13'h673: dout  = 8'b00000000; // 1651 :   0 - 0x0
      13'h674: dout  = 8'b00000000; // 1652 :   0 - 0x0
      13'h675: dout  = 8'b00000000; // 1653 :   0 - 0x0
      13'h676: dout  = 8'b00000000; // 1654 :   0 - 0x0
      13'h677: dout  = 8'b00000000; // 1655 :   0 - 0x0
      13'h678: dout  = 8'b00000000; // 1656 :   0 - 0x0
      13'h679: dout  = 8'b00000000; // 1657 :   0 - 0x0
      13'h67A: dout  = 8'b00000000; // 1658 :   0 - 0x0
      13'h67B: dout  = 8'b00000000; // 1659 :   0 - 0x0
      13'h67C: dout  = 8'b00000000; // 1660 :   0 - 0x0
      13'h67D: dout  = 8'b00000000; // 1661 :   0 - 0x0
      13'h67E: dout  = 8'b00000000; // 1662 :   0 - 0x0
      13'h67F: dout  = 8'b00000000; // 1663 :   0 - 0x0
      13'h680: dout  = 8'b00000000; // 1664 :   0 - 0x0 -- Sprite 0x68
      13'h681: dout  = 8'b00000000; // 1665 :   0 - 0x0
      13'h682: dout  = 8'b00000000; // 1666 :   0 - 0x0
      13'h683: dout  = 8'b00000000; // 1667 :   0 - 0x0
      13'h684: dout  = 8'b00000000; // 1668 :   0 - 0x0
      13'h685: dout  = 8'b00000000; // 1669 :   0 - 0x0
      13'h686: dout  = 8'b00000000; // 1670 :   0 - 0x0
      13'h687: dout  = 8'b00000000; // 1671 :   0 - 0x0
      13'h688: dout  = 8'b00000000; // 1672 :   0 - 0x0
      13'h689: dout  = 8'b00000000; // 1673 :   0 - 0x0
      13'h68A: dout  = 8'b00000000; // 1674 :   0 - 0x0
      13'h68B: dout  = 8'b00000000; // 1675 :   0 - 0x0
      13'h68C: dout  = 8'b00000000; // 1676 :   0 - 0x0
      13'h68D: dout  = 8'b00000000; // 1677 :   0 - 0x0
      13'h68E: dout  = 8'b00000000; // 1678 :   0 - 0x0
      13'h68F: dout  = 8'b00000000; // 1679 :   0 - 0x0
      13'h690: dout  = 8'b00000000; // 1680 :   0 - 0x0 -- Sprite 0x69
      13'h691: dout  = 8'b00000000; // 1681 :   0 - 0x0
      13'h692: dout  = 8'b00000000; // 1682 :   0 - 0x0
      13'h693: dout  = 8'b00000000; // 1683 :   0 - 0x0
      13'h694: dout  = 8'b00000000; // 1684 :   0 - 0x0
      13'h695: dout  = 8'b00000000; // 1685 :   0 - 0x0
      13'h696: dout  = 8'b00000000; // 1686 :   0 - 0x0
      13'h697: dout  = 8'b00000000; // 1687 :   0 - 0x0
      13'h698: dout  = 8'b00000000; // 1688 :   0 - 0x0
      13'h699: dout  = 8'b00000000; // 1689 :   0 - 0x0
      13'h69A: dout  = 8'b00000000; // 1690 :   0 - 0x0
      13'h69B: dout  = 8'b00000000; // 1691 :   0 - 0x0
      13'h69C: dout  = 8'b00000000; // 1692 :   0 - 0x0
      13'h69D: dout  = 8'b00000000; // 1693 :   0 - 0x0
      13'h69E: dout  = 8'b00000000; // 1694 :   0 - 0x0
      13'h69F: dout  = 8'b00000000; // 1695 :   0 - 0x0
      13'h6A0: dout  = 8'b00000000; // 1696 :   0 - 0x0 -- Sprite 0x6a
      13'h6A1: dout  = 8'b00000000; // 1697 :   0 - 0x0
      13'h6A2: dout  = 8'b00000000; // 1698 :   0 - 0x0
      13'h6A3: dout  = 8'b00000000; // 1699 :   0 - 0x0
      13'h6A4: dout  = 8'b00000000; // 1700 :   0 - 0x0
      13'h6A5: dout  = 8'b00000000; // 1701 :   0 - 0x0
      13'h6A6: dout  = 8'b00000000; // 1702 :   0 - 0x0
      13'h6A7: dout  = 8'b00000000; // 1703 :   0 - 0x0
      13'h6A8: dout  = 8'b00000000; // 1704 :   0 - 0x0
      13'h6A9: dout  = 8'b00000000; // 1705 :   0 - 0x0
      13'h6AA: dout  = 8'b00000000; // 1706 :   0 - 0x0
      13'h6AB: dout  = 8'b00000000; // 1707 :   0 - 0x0
      13'h6AC: dout  = 8'b00000000; // 1708 :   0 - 0x0
      13'h6AD: dout  = 8'b00000000; // 1709 :   0 - 0x0
      13'h6AE: dout  = 8'b00000000; // 1710 :   0 - 0x0
      13'h6AF: dout  = 8'b00000000; // 1711 :   0 - 0x0
      13'h6B0: dout  = 8'b00000000; // 1712 :   0 - 0x0 -- Sprite 0x6b
      13'h6B1: dout  = 8'b00000000; // 1713 :   0 - 0x0
      13'h6B2: dout  = 8'b00000000; // 1714 :   0 - 0x0
      13'h6B3: dout  = 8'b00000000; // 1715 :   0 - 0x0
      13'h6B4: dout  = 8'b00000000; // 1716 :   0 - 0x0
      13'h6B5: dout  = 8'b00000000; // 1717 :   0 - 0x0
      13'h6B6: dout  = 8'b00000000; // 1718 :   0 - 0x0
      13'h6B7: dout  = 8'b00000000; // 1719 :   0 - 0x0
      13'h6B8: dout  = 8'b00000000; // 1720 :   0 - 0x0
      13'h6B9: dout  = 8'b00000000; // 1721 :   0 - 0x0
      13'h6BA: dout  = 8'b00000000; // 1722 :   0 - 0x0
      13'h6BB: dout  = 8'b00000000; // 1723 :   0 - 0x0
      13'h6BC: dout  = 8'b00000000; // 1724 :   0 - 0x0
      13'h6BD: dout  = 8'b00000000; // 1725 :   0 - 0x0
      13'h6BE: dout  = 8'b00000000; // 1726 :   0 - 0x0
      13'h6BF: dout  = 8'b00000000; // 1727 :   0 - 0x0
      13'h6C0: dout  = 8'b00000000; // 1728 :   0 - 0x0 -- Sprite 0x6c
      13'h6C1: dout  = 8'b00000000; // 1729 :   0 - 0x0
      13'h6C2: dout  = 8'b00000000; // 1730 :   0 - 0x0
      13'h6C3: dout  = 8'b00000000; // 1731 :   0 - 0x0
      13'h6C4: dout  = 8'b00000000; // 1732 :   0 - 0x0
      13'h6C5: dout  = 8'b00000000; // 1733 :   0 - 0x0
      13'h6C6: dout  = 8'b00000000; // 1734 :   0 - 0x0
      13'h6C7: dout  = 8'b00000000; // 1735 :   0 - 0x0
      13'h6C8: dout  = 8'b00000000; // 1736 :   0 - 0x0
      13'h6C9: dout  = 8'b00000000; // 1737 :   0 - 0x0
      13'h6CA: dout  = 8'b00000000; // 1738 :   0 - 0x0
      13'h6CB: dout  = 8'b00000000; // 1739 :   0 - 0x0
      13'h6CC: dout  = 8'b00000000; // 1740 :   0 - 0x0
      13'h6CD: dout  = 8'b00000000; // 1741 :   0 - 0x0
      13'h6CE: dout  = 8'b00000000; // 1742 :   0 - 0x0
      13'h6CF: dout  = 8'b00000000; // 1743 :   0 - 0x0
      13'h6D0: dout  = 8'b00000000; // 1744 :   0 - 0x0 -- Sprite 0x6d
      13'h6D1: dout  = 8'b00000000; // 1745 :   0 - 0x0
      13'h6D2: dout  = 8'b00000000; // 1746 :   0 - 0x0
      13'h6D3: dout  = 8'b00000000; // 1747 :   0 - 0x0
      13'h6D4: dout  = 8'b00000000; // 1748 :   0 - 0x0
      13'h6D5: dout  = 8'b00000000; // 1749 :   0 - 0x0
      13'h6D6: dout  = 8'b00000000; // 1750 :   0 - 0x0
      13'h6D7: dout  = 8'b00000000; // 1751 :   0 - 0x0
      13'h6D8: dout  = 8'b00000000; // 1752 :   0 - 0x0
      13'h6D9: dout  = 8'b00000000; // 1753 :   0 - 0x0
      13'h6DA: dout  = 8'b00000000; // 1754 :   0 - 0x0
      13'h6DB: dout  = 8'b00000000; // 1755 :   0 - 0x0
      13'h6DC: dout  = 8'b00000000; // 1756 :   0 - 0x0
      13'h6DD: dout  = 8'b00000000; // 1757 :   0 - 0x0
      13'h6DE: dout  = 8'b00000000; // 1758 :   0 - 0x0
      13'h6DF: dout  = 8'b00000000; // 1759 :   0 - 0x0
      13'h6E0: dout  = 8'b00000000; // 1760 :   0 - 0x0 -- Sprite 0x6e
      13'h6E1: dout  = 8'b00000000; // 1761 :   0 - 0x0
      13'h6E2: dout  = 8'b00000000; // 1762 :   0 - 0x0
      13'h6E3: dout  = 8'b00000000; // 1763 :   0 - 0x0
      13'h6E4: dout  = 8'b00000000; // 1764 :   0 - 0x0
      13'h6E5: dout  = 8'b00000000; // 1765 :   0 - 0x0
      13'h6E6: dout  = 8'b00000000; // 1766 :   0 - 0x0
      13'h6E7: dout  = 8'b00000000; // 1767 :   0 - 0x0
      13'h6E8: dout  = 8'b00000000; // 1768 :   0 - 0x0
      13'h6E9: dout  = 8'b00000000; // 1769 :   0 - 0x0
      13'h6EA: dout  = 8'b00000000; // 1770 :   0 - 0x0
      13'h6EB: dout  = 8'b00000000; // 1771 :   0 - 0x0
      13'h6EC: dout  = 8'b00000000; // 1772 :   0 - 0x0
      13'h6ED: dout  = 8'b00000000; // 1773 :   0 - 0x0
      13'h6EE: dout  = 8'b00000000; // 1774 :   0 - 0x0
      13'h6EF: dout  = 8'b00000000; // 1775 :   0 - 0x0
      13'h6F0: dout  = 8'b00000000; // 1776 :   0 - 0x0 -- Sprite 0x6f
      13'h6F1: dout  = 8'b00000000; // 1777 :   0 - 0x0
      13'h6F2: dout  = 8'b00000000; // 1778 :   0 - 0x0
      13'h6F3: dout  = 8'b00000000; // 1779 :   0 - 0x0
      13'h6F4: dout  = 8'b00000000; // 1780 :   0 - 0x0
      13'h6F5: dout  = 8'b00000000; // 1781 :   0 - 0x0
      13'h6F6: dout  = 8'b00000000; // 1782 :   0 - 0x0
      13'h6F7: dout  = 8'b00000000; // 1783 :   0 - 0x0
      13'h6F8: dout  = 8'b00000000; // 1784 :   0 - 0x0
      13'h6F9: dout  = 8'b00000000; // 1785 :   0 - 0x0
      13'h6FA: dout  = 8'b00000000; // 1786 :   0 - 0x0
      13'h6FB: dout  = 8'b00000000; // 1787 :   0 - 0x0
      13'h6FC: dout  = 8'b00000000; // 1788 :   0 - 0x0
      13'h6FD: dout  = 8'b00000000; // 1789 :   0 - 0x0
      13'h6FE: dout  = 8'b00000000; // 1790 :   0 - 0x0
      13'h6FF: dout  = 8'b00000000; // 1791 :   0 - 0x0
      13'h700: dout  = 8'b00000000; // 1792 :   0 - 0x0 -- Sprite 0x70
      13'h701: dout  = 8'b00000000; // 1793 :   0 - 0x0
      13'h702: dout  = 8'b00000000; // 1794 :   0 - 0x0
      13'h703: dout  = 8'b00000000; // 1795 :   0 - 0x0
      13'h704: dout  = 8'b00000000; // 1796 :   0 - 0x0
      13'h705: dout  = 8'b00000000; // 1797 :   0 - 0x0
      13'h706: dout  = 8'b00000000; // 1798 :   0 - 0x0
      13'h707: dout  = 8'b00000000; // 1799 :   0 - 0x0
      13'h708: dout  = 8'b00000000; // 1800 :   0 - 0x0
      13'h709: dout  = 8'b00000000; // 1801 :   0 - 0x0
      13'h70A: dout  = 8'b00000000; // 1802 :   0 - 0x0
      13'h70B: dout  = 8'b00000000; // 1803 :   0 - 0x0
      13'h70C: dout  = 8'b00000000; // 1804 :   0 - 0x0
      13'h70D: dout  = 8'b00000000; // 1805 :   0 - 0x0
      13'h70E: dout  = 8'b00000000; // 1806 :   0 - 0x0
      13'h70F: dout  = 8'b00000000; // 1807 :   0 - 0x0
      13'h710: dout  = 8'b00000000; // 1808 :   0 - 0x0 -- Sprite 0x71
      13'h711: dout  = 8'b00000000; // 1809 :   0 - 0x0
      13'h712: dout  = 8'b00000000; // 1810 :   0 - 0x0
      13'h713: dout  = 8'b00000000; // 1811 :   0 - 0x0
      13'h714: dout  = 8'b00000000; // 1812 :   0 - 0x0
      13'h715: dout  = 8'b00000000; // 1813 :   0 - 0x0
      13'h716: dout  = 8'b00000000; // 1814 :   0 - 0x0
      13'h717: dout  = 8'b00000000; // 1815 :   0 - 0x0
      13'h718: dout  = 8'b00000000; // 1816 :   0 - 0x0
      13'h719: dout  = 8'b00000000; // 1817 :   0 - 0x0
      13'h71A: dout  = 8'b00000000; // 1818 :   0 - 0x0
      13'h71B: dout  = 8'b00000000; // 1819 :   0 - 0x0
      13'h71C: dout  = 8'b00000000; // 1820 :   0 - 0x0
      13'h71D: dout  = 8'b00000000; // 1821 :   0 - 0x0
      13'h71E: dout  = 8'b00000000; // 1822 :   0 - 0x0
      13'h71F: dout  = 8'b00000000; // 1823 :   0 - 0x0
      13'h720: dout  = 8'b00000000; // 1824 :   0 - 0x0 -- Sprite 0x72
      13'h721: dout  = 8'b00000000; // 1825 :   0 - 0x0
      13'h722: dout  = 8'b00000000; // 1826 :   0 - 0x0
      13'h723: dout  = 8'b00000000; // 1827 :   0 - 0x0
      13'h724: dout  = 8'b00000000; // 1828 :   0 - 0x0
      13'h725: dout  = 8'b00000000; // 1829 :   0 - 0x0
      13'h726: dout  = 8'b00000000; // 1830 :   0 - 0x0
      13'h727: dout  = 8'b00000000; // 1831 :   0 - 0x0
      13'h728: dout  = 8'b00000000; // 1832 :   0 - 0x0
      13'h729: dout  = 8'b00000000; // 1833 :   0 - 0x0
      13'h72A: dout  = 8'b00000000; // 1834 :   0 - 0x0
      13'h72B: dout  = 8'b00000000; // 1835 :   0 - 0x0
      13'h72C: dout  = 8'b00000000; // 1836 :   0 - 0x0
      13'h72D: dout  = 8'b00000000; // 1837 :   0 - 0x0
      13'h72E: dout  = 8'b00000000; // 1838 :   0 - 0x0
      13'h72F: dout  = 8'b00000000; // 1839 :   0 - 0x0
      13'h730: dout  = 8'b00000000; // 1840 :   0 - 0x0 -- Sprite 0x73
      13'h731: dout  = 8'b00000000; // 1841 :   0 - 0x0
      13'h732: dout  = 8'b00000000; // 1842 :   0 - 0x0
      13'h733: dout  = 8'b00000000; // 1843 :   0 - 0x0
      13'h734: dout  = 8'b00000000; // 1844 :   0 - 0x0
      13'h735: dout  = 8'b00000000; // 1845 :   0 - 0x0
      13'h736: dout  = 8'b00000000; // 1846 :   0 - 0x0
      13'h737: dout  = 8'b00000000; // 1847 :   0 - 0x0
      13'h738: dout  = 8'b00000000; // 1848 :   0 - 0x0
      13'h739: dout  = 8'b00000000; // 1849 :   0 - 0x0
      13'h73A: dout  = 8'b00000000; // 1850 :   0 - 0x0
      13'h73B: dout  = 8'b00000000; // 1851 :   0 - 0x0
      13'h73C: dout  = 8'b00000000; // 1852 :   0 - 0x0
      13'h73D: dout  = 8'b00000000; // 1853 :   0 - 0x0
      13'h73E: dout  = 8'b00000000; // 1854 :   0 - 0x0
      13'h73F: dout  = 8'b00000000; // 1855 :   0 - 0x0
      13'h740: dout  = 8'b00000000; // 1856 :   0 - 0x0 -- Sprite 0x74
      13'h741: dout  = 8'b00000000; // 1857 :   0 - 0x0
      13'h742: dout  = 8'b00000000; // 1858 :   0 - 0x0
      13'h743: dout  = 8'b00000000; // 1859 :   0 - 0x0
      13'h744: dout  = 8'b00000000; // 1860 :   0 - 0x0
      13'h745: dout  = 8'b00000000; // 1861 :   0 - 0x0
      13'h746: dout  = 8'b00000000; // 1862 :   0 - 0x0
      13'h747: dout  = 8'b00000000; // 1863 :   0 - 0x0
      13'h748: dout  = 8'b00000000; // 1864 :   0 - 0x0
      13'h749: dout  = 8'b00000000; // 1865 :   0 - 0x0
      13'h74A: dout  = 8'b00000000; // 1866 :   0 - 0x0
      13'h74B: dout  = 8'b00000000; // 1867 :   0 - 0x0
      13'h74C: dout  = 8'b00000000; // 1868 :   0 - 0x0
      13'h74D: dout  = 8'b00000000; // 1869 :   0 - 0x0
      13'h74E: dout  = 8'b00000000; // 1870 :   0 - 0x0
      13'h74F: dout  = 8'b00000000; // 1871 :   0 - 0x0
      13'h750: dout  = 8'b00000000; // 1872 :   0 - 0x0 -- Sprite 0x75
      13'h751: dout  = 8'b00000000; // 1873 :   0 - 0x0
      13'h752: dout  = 8'b00000000; // 1874 :   0 - 0x0
      13'h753: dout  = 8'b00000000; // 1875 :   0 - 0x0
      13'h754: dout  = 8'b00000000; // 1876 :   0 - 0x0
      13'h755: dout  = 8'b00000000; // 1877 :   0 - 0x0
      13'h756: dout  = 8'b00000000; // 1878 :   0 - 0x0
      13'h757: dout  = 8'b00000000; // 1879 :   0 - 0x0
      13'h758: dout  = 8'b00000000; // 1880 :   0 - 0x0
      13'h759: dout  = 8'b00000000; // 1881 :   0 - 0x0
      13'h75A: dout  = 8'b00000000; // 1882 :   0 - 0x0
      13'h75B: dout  = 8'b00000000; // 1883 :   0 - 0x0
      13'h75C: dout  = 8'b00000000; // 1884 :   0 - 0x0
      13'h75D: dout  = 8'b00000000; // 1885 :   0 - 0x0
      13'h75E: dout  = 8'b00000000; // 1886 :   0 - 0x0
      13'h75F: dout  = 8'b00000000; // 1887 :   0 - 0x0
      13'h760: dout  = 8'b00000000; // 1888 :   0 - 0x0 -- Sprite 0x76
      13'h761: dout  = 8'b00000000; // 1889 :   0 - 0x0
      13'h762: dout  = 8'b00000000; // 1890 :   0 - 0x0
      13'h763: dout  = 8'b00000000; // 1891 :   0 - 0x0
      13'h764: dout  = 8'b00000000; // 1892 :   0 - 0x0
      13'h765: dout  = 8'b00000000; // 1893 :   0 - 0x0
      13'h766: dout  = 8'b00000000; // 1894 :   0 - 0x0
      13'h767: dout  = 8'b00000000; // 1895 :   0 - 0x0
      13'h768: dout  = 8'b00000000; // 1896 :   0 - 0x0
      13'h769: dout  = 8'b00000000; // 1897 :   0 - 0x0
      13'h76A: dout  = 8'b00000000; // 1898 :   0 - 0x0
      13'h76B: dout  = 8'b00000000; // 1899 :   0 - 0x0
      13'h76C: dout  = 8'b00000000; // 1900 :   0 - 0x0
      13'h76D: dout  = 8'b00000000; // 1901 :   0 - 0x0
      13'h76E: dout  = 8'b00000000; // 1902 :   0 - 0x0
      13'h76F: dout  = 8'b00000000; // 1903 :   0 - 0x0
      13'h770: dout  = 8'b00000000; // 1904 :   0 - 0x0 -- Sprite 0x77
      13'h771: dout  = 8'b00000000; // 1905 :   0 - 0x0
      13'h772: dout  = 8'b00000000; // 1906 :   0 - 0x0
      13'h773: dout  = 8'b00000000; // 1907 :   0 - 0x0
      13'h774: dout  = 8'b00000000; // 1908 :   0 - 0x0
      13'h775: dout  = 8'b00000000; // 1909 :   0 - 0x0
      13'h776: dout  = 8'b00000000; // 1910 :   0 - 0x0
      13'h777: dout  = 8'b00000000; // 1911 :   0 - 0x0
      13'h778: dout  = 8'b00000000; // 1912 :   0 - 0x0
      13'h779: dout  = 8'b00000000; // 1913 :   0 - 0x0
      13'h77A: dout  = 8'b00000000; // 1914 :   0 - 0x0
      13'h77B: dout  = 8'b00000000; // 1915 :   0 - 0x0
      13'h77C: dout  = 8'b00000000; // 1916 :   0 - 0x0
      13'h77D: dout  = 8'b00000000; // 1917 :   0 - 0x0
      13'h77E: dout  = 8'b00000000; // 1918 :   0 - 0x0
      13'h77F: dout  = 8'b00000000; // 1919 :   0 - 0x0
      13'h780: dout  = 8'b00000000; // 1920 :   0 - 0x0 -- Sprite 0x78
      13'h781: dout  = 8'b00000000; // 1921 :   0 - 0x0
      13'h782: dout  = 8'b00000000; // 1922 :   0 - 0x0
      13'h783: dout  = 8'b00000000; // 1923 :   0 - 0x0
      13'h784: dout  = 8'b00000000; // 1924 :   0 - 0x0
      13'h785: dout  = 8'b00000000; // 1925 :   0 - 0x0
      13'h786: dout  = 8'b00000000; // 1926 :   0 - 0x0
      13'h787: dout  = 8'b00000000; // 1927 :   0 - 0x0
      13'h788: dout  = 8'b00000000; // 1928 :   0 - 0x0
      13'h789: dout  = 8'b00000000; // 1929 :   0 - 0x0
      13'h78A: dout  = 8'b00000000; // 1930 :   0 - 0x0
      13'h78B: dout  = 8'b00000000; // 1931 :   0 - 0x0
      13'h78C: dout  = 8'b00000000; // 1932 :   0 - 0x0
      13'h78D: dout  = 8'b00000000; // 1933 :   0 - 0x0
      13'h78E: dout  = 8'b00000000; // 1934 :   0 - 0x0
      13'h78F: dout  = 8'b00000000; // 1935 :   0 - 0x0
      13'h790: dout  = 8'b00000000; // 1936 :   0 - 0x0 -- Sprite 0x79
      13'h791: dout  = 8'b00000000; // 1937 :   0 - 0x0
      13'h792: dout  = 8'b00000000; // 1938 :   0 - 0x0
      13'h793: dout  = 8'b00000000; // 1939 :   0 - 0x0
      13'h794: dout  = 8'b00000000; // 1940 :   0 - 0x0
      13'h795: dout  = 8'b00000000; // 1941 :   0 - 0x0
      13'h796: dout  = 8'b00000000; // 1942 :   0 - 0x0
      13'h797: dout  = 8'b00000000; // 1943 :   0 - 0x0
      13'h798: dout  = 8'b00000000; // 1944 :   0 - 0x0
      13'h799: dout  = 8'b00000000; // 1945 :   0 - 0x0
      13'h79A: dout  = 8'b00000000; // 1946 :   0 - 0x0
      13'h79B: dout  = 8'b00000000; // 1947 :   0 - 0x0
      13'h79C: dout  = 8'b00000000; // 1948 :   0 - 0x0
      13'h79D: dout  = 8'b00000000; // 1949 :   0 - 0x0
      13'h79E: dout  = 8'b00000000; // 1950 :   0 - 0x0
      13'h79F: dout  = 8'b00000000; // 1951 :   0 - 0x0
      13'h7A0: dout  = 8'b00000000; // 1952 :   0 - 0x0 -- Sprite 0x7a
      13'h7A1: dout  = 8'b00000000; // 1953 :   0 - 0x0
      13'h7A2: dout  = 8'b00000000; // 1954 :   0 - 0x0
      13'h7A3: dout  = 8'b00000000; // 1955 :   0 - 0x0
      13'h7A4: dout  = 8'b00000000; // 1956 :   0 - 0x0
      13'h7A5: dout  = 8'b00000000; // 1957 :   0 - 0x0
      13'h7A6: dout  = 8'b00000000; // 1958 :   0 - 0x0
      13'h7A7: dout  = 8'b00000000; // 1959 :   0 - 0x0
      13'h7A8: dout  = 8'b00000000; // 1960 :   0 - 0x0
      13'h7A9: dout  = 8'b00000000; // 1961 :   0 - 0x0
      13'h7AA: dout  = 8'b00000000; // 1962 :   0 - 0x0
      13'h7AB: dout  = 8'b00000000; // 1963 :   0 - 0x0
      13'h7AC: dout  = 8'b00000000; // 1964 :   0 - 0x0
      13'h7AD: dout  = 8'b00000000; // 1965 :   0 - 0x0
      13'h7AE: dout  = 8'b00000000; // 1966 :   0 - 0x0
      13'h7AF: dout  = 8'b00000000; // 1967 :   0 - 0x0
      13'h7B0: dout  = 8'b00000000; // 1968 :   0 - 0x0 -- Sprite 0x7b
      13'h7B1: dout  = 8'b00000000; // 1969 :   0 - 0x0
      13'h7B2: dout  = 8'b00000000; // 1970 :   0 - 0x0
      13'h7B3: dout  = 8'b00000000; // 1971 :   0 - 0x0
      13'h7B4: dout  = 8'b00000000; // 1972 :   0 - 0x0
      13'h7B5: dout  = 8'b00000000; // 1973 :   0 - 0x0
      13'h7B6: dout  = 8'b00000000; // 1974 :   0 - 0x0
      13'h7B7: dout  = 8'b00000000; // 1975 :   0 - 0x0
      13'h7B8: dout  = 8'b00000000; // 1976 :   0 - 0x0
      13'h7B9: dout  = 8'b00000000; // 1977 :   0 - 0x0
      13'h7BA: dout  = 8'b00000000; // 1978 :   0 - 0x0
      13'h7BB: dout  = 8'b00000000; // 1979 :   0 - 0x0
      13'h7BC: dout  = 8'b00000000; // 1980 :   0 - 0x0
      13'h7BD: dout  = 8'b00000000; // 1981 :   0 - 0x0
      13'h7BE: dout  = 8'b00000000; // 1982 :   0 - 0x0
      13'h7BF: dout  = 8'b00000000; // 1983 :   0 - 0x0
      13'h7C0: dout  = 8'b00000000; // 1984 :   0 - 0x0 -- Sprite 0x7c
      13'h7C1: dout  = 8'b00000000; // 1985 :   0 - 0x0
      13'h7C2: dout  = 8'b00000000; // 1986 :   0 - 0x0
      13'h7C3: dout  = 8'b00000000; // 1987 :   0 - 0x0
      13'h7C4: dout  = 8'b00000000; // 1988 :   0 - 0x0
      13'h7C5: dout  = 8'b00000000; // 1989 :   0 - 0x0
      13'h7C6: dout  = 8'b00000000; // 1990 :   0 - 0x0
      13'h7C7: dout  = 8'b00000000; // 1991 :   0 - 0x0
      13'h7C8: dout  = 8'b00000000; // 1992 :   0 - 0x0
      13'h7C9: dout  = 8'b00000000; // 1993 :   0 - 0x0
      13'h7CA: dout  = 8'b00000000; // 1994 :   0 - 0x0
      13'h7CB: dout  = 8'b00000000; // 1995 :   0 - 0x0
      13'h7CC: dout  = 8'b00000000; // 1996 :   0 - 0x0
      13'h7CD: dout  = 8'b00000000; // 1997 :   0 - 0x0
      13'h7CE: dout  = 8'b00000000; // 1998 :   0 - 0x0
      13'h7CF: dout  = 8'b00000000; // 1999 :   0 - 0x0
      13'h7D0: dout  = 8'b00000000; // 2000 :   0 - 0x0 -- Sprite 0x7d
      13'h7D1: dout  = 8'b00000000; // 2001 :   0 - 0x0
      13'h7D2: dout  = 8'b00000000; // 2002 :   0 - 0x0
      13'h7D3: dout  = 8'b00000000; // 2003 :   0 - 0x0
      13'h7D4: dout  = 8'b00000000; // 2004 :   0 - 0x0
      13'h7D5: dout  = 8'b00000000; // 2005 :   0 - 0x0
      13'h7D6: dout  = 8'b00000000; // 2006 :   0 - 0x0
      13'h7D7: dout  = 8'b00000000; // 2007 :   0 - 0x0
      13'h7D8: dout  = 8'b00000000; // 2008 :   0 - 0x0
      13'h7D9: dout  = 8'b00000000; // 2009 :   0 - 0x0
      13'h7DA: dout  = 8'b00000000; // 2010 :   0 - 0x0
      13'h7DB: dout  = 8'b00000000; // 2011 :   0 - 0x0
      13'h7DC: dout  = 8'b00000000; // 2012 :   0 - 0x0
      13'h7DD: dout  = 8'b00000000; // 2013 :   0 - 0x0
      13'h7DE: dout  = 8'b00000000; // 2014 :   0 - 0x0
      13'h7DF: dout  = 8'b00000000; // 2015 :   0 - 0x0
      13'h7E0: dout  = 8'b00000000; // 2016 :   0 - 0x0 -- Sprite 0x7e
      13'h7E1: dout  = 8'b00000000; // 2017 :   0 - 0x0
      13'h7E2: dout  = 8'b00000000; // 2018 :   0 - 0x0
      13'h7E3: dout  = 8'b00000000; // 2019 :   0 - 0x0
      13'h7E4: dout  = 8'b00000000; // 2020 :   0 - 0x0
      13'h7E5: dout  = 8'b00000000; // 2021 :   0 - 0x0
      13'h7E6: dout  = 8'b00000000; // 2022 :   0 - 0x0
      13'h7E7: dout  = 8'b00000000; // 2023 :   0 - 0x0
      13'h7E8: dout  = 8'b00000000; // 2024 :   0 - 0x0
      13'h7E9: dout  = 8'b00000000; // 2025 :   0 - 0x0
      13'h7EA: dout  = 8'b00000000; // 2026 :   0 - 0x0
      13'h7EB: dout  = 8'b00000000; // 2027 :   0 - 0x0
      13'h7EC: dout  = 8'b00000000; // 2028 :   0 - 0x0
      13'h7ED: dout  = 8'b00000000; // 2029 :   0 - 0x0
      13'h7EE: dout  = 8'b00000000; // 2030 :   0 - 0x0
      13'h7EF: dout  = 8'b00000000; // 2031 :   0 - 0x0
      13'h7F0: dout  = 8'b00000000; // 2032 :   0 - 0x0 -- Sprite 0x7f
      13'h7F1: dout  = 8'b00000000; // 2033 :   0 - 0x0
      13'h7F2: dout  = 8'b00000000; // 2034 :   0 - 0x0
      13'h7F3: dout  = 8'b00000000; // 2035 :   0 - 0x0
      13'h7F4: dout  = 8'b00000000; // 2036 :   0 - 0x0
      13'h7F5: dout  = 8'b00000000; // 2037 :   0 - 0x0
      13'h7F6: dout  = 8'b00000000; // 2038 :   0 - 0x0
      13'h7F7: dout  = 8'b00000000; // 2039 :   0 - 0x0
      13'h7F8: dout  = 8'b00000000; // 2040 :   0 - 0x0
      13'h7F9: dout  = 8'b00000000; // 2041 :   0 - 0x0
      13'h7FA: dout  = 8'b00000000; // 2042 :   0 - 0x0
      13'h7FB: dout  = 8'b00000000; // 2043 :   0 - 0x0
      13'h7FC: dout  = 8'b00000000; // 2044 :   0 - 0x0
      13'h7FD: dout  = 8'b00000000; // 2045 :   0 - 0x0
      13'h7FE: dout  = 8'b00000000; // 2046 :   0 - 0x0
      13'h7FF: dout  = 8'b00000000; // 2047 :   0 - 0x0
      13'h800: dout  = 8'b00000000; // 2048 :   0 - 0x0 -- Sprite 0x80
      13'h801: dout  = 8'b00000000; // 2049 :   0 - 0x0
      13'h802: dout  = 8'b00000000; // 2050 :   0 - 0x0
      13'h803: dout  = 8'b00000000; // 2051 :   0 - 0x0
      13'h804: dout  = 8'b00000000; // 2052 :   0 - 0x0
      13'h805: dout  = 8'b00000000; // 2053 :   0 - 0x0
      13'h806: dout  = 8'b00000000; // 2054 :   0 - 0x0
      13'h807: dout  = 8'b00000000; // 2055 :   0 - 0x0
      13'h808: dout  = 8'b00000000; // 2056 :   0 - 0x0
      13'h809: dout  = 8'b00000000; // 2057 :   0 - 0x0
      13'h80A: dout  = 8'b00000000; // 2058 :   0 - 0x0
      13'h80B: dout  = 8'b00000000; // 2059 :   0 - 0x0
      13'h80C: dout  = 8'b00000000; // 2060 :   0 - 0x0
      13'h80D: dout  = 8'b00000000; // 2061 :   0 - 0x0
      13'h80E: dout  = 8'b00000000; // 2062 :   0 - 0x0
      13'h80F: dout  = 8'b00000000; // 2063 :   0 - 0x0
      13'h810: dout  = 8'b00000000; // 2064 :   0 - 0x0 -- Sprite 0x81
      13'h811: dout  = 8'b00000000; // 2065 :   0 - 0x0
      13'h812: dout  = 8'b00000000; // 2066 :   0 - 0x0
      13'h813: dout  = 8'b00000000; // 2067 :   0 - 0x0
      13'h814: dout  = 8'b00000000; // 2068 :   0 - 0x0
      13'h815: dout  = 8'b00000000; // 2069 :   0 - 0x0
      13'h816: dout  = 8'b00000000; // 2070 :   0 - 0x0
      13'h817: dout  = 8'b00000000; // 2071 :   0 - 0x0
      13'h818: dout  = 8'b00000000; // 2072 :   0 - 0x0
      13'h819: dout  = 8'b00000000; // 2073 :   0 - 0x0
      13'h81A: dout  = 8'b00000000; // 2074 :   0 - 0x0
      13'h81B: dout  = 8'b00000000; // 2075 :   0 - 0x0
      13'h81C: dout  = 8'b00000000; // 2076 :   0 - 0x0
      13'h81D: dout  = 8'b00000000; // 2077 :   0 - 0x0
      13'h81E: dout  = 8'b00000000; // 2078 :   0 - 0x0
      13'h81F: dout  = 8'b00000000; // 2079 :   0 - 0x0
      13'h820: dout  = 8'b00000000; // 2080 :   0 - 0x0 -- Sprite 0x82
      13'h821: dout  = 8'b00000000; // 2081 :   0 - 0x0
      13'h822: dout  = 8'b00000000; // 2082 :   0 - 0x0
      13'h823: dout  = 8'b00000000; // 2083 :   0 - 0x0
      13'h824: dout  = 8'b00000000; // 2084 :   0 - 0x0
      13'h825: dout  = 8'b00000000; // 2085 :   0 - 0x0
      13'h826: dout  = 8'b00000000; // 2086 :   0 - 0x0
      13'h827: dout  = 8'b00000000; // 2087 :   0 - 0x0
      13'h828: dout  = 8'b00000000; // 2088 :   0 - 0x0
      13'h829: dout  = 8'b00000000; // 2089 :   0 - 0x0
      13'h82A: dout  = 8'b00000000; // 2090 :   0 - 0x0
      13'h82B: dout  = 8'b00000000; // 2091 :   0 - 0x0
      13'h82C: dout  = 8'b00000000; // 2092 :   0 - 0x0
      13'h82D: dout  = 8'b00000000; // 2093 :   0 - 0x0
      13'h82E: dout  = 8'b00000000; // 2094 :   0 - 0x0
      13'h82F: dout  = 8'b00000000; // 2095 :   0 - 0x0
      13'h830: dout  = 8'b00000000; // 2096 :   0 - 0x0 -- Sprite 0x83
      13'h831: dout  = 8'b00000000; // 2097 :   0 - 0x0
      13'h832: dout  = 8'b00000000; // 2098 :   0 - 0x0
      13'h833: dout  = 8'b00000000; // 2099 :   0 - 0x0
      13'h834: dout  = 8'b00000000; // 2100 :   0 - 0x0
      13'h835: dout  = 8'b00000000; // 2101 :   0 - 0x0
      13'h836: dout  = 8'b00000000; // 2102 :   0 - 0x0
      13'h837: dout  = 8'b00000000; // 2103 :   0 - 0x0
      13'h838: dout  = 8'b00000000; // 2104 :   0 - 0x0
      13'h839: dout  = 8'b00000000; // 2105 :   0 - 0x0
      13'h83A: dout  = 8'b00000000; // 2106 :   0 - 0x0
      13'h83B: dout  = 8'b00000000; // 2107 :   0 - 0x0
      13'h83C: dout  = 8'b00000000; // 2108 :   0 - 0x0
      13'h83D: dout  = 8'b00000000; // 2109 :   0 - 0x0
      13'h83E: dout  = 8'b00000000; // 2110 :   0 - 0x0
      13'h83F: dout  = 8'b00000000; // 2111 :   0 - 0x0
      13'h840: dout  = 8'b00000000; // 2112 :   0 - 0x0 -- Sprite 0x84
      13'h841: dout  = 8'b00000000; // 2113 :   0 - 0x0
      13'h842: dout  = 8'b00000000; // 2114 :   0 - 0x0
      13'h843: dout  = 8'b00000000; // 2115 :   0 - 0x0
      13'h844: dout  = 8'b00000000; // 2116 :   0 - 0x0
      13'h845: dout  = 8'b00000000; // 2117 :   0 - 0x0
      13'h846: dout  = 8'b00000000; // 2118 :   0 - 0x0
      13'h847: dout  = 8'b00000000; // 2119 :   0 - 0x0
      13'h848: dout  = 8'b00000000; // 2120 :   0 - 0x0
      13'h849: dout  = 8'b00000000; // 2121 :   0 - 0x0
      13'h84A: dout  = 8'b00000000; // 2122 :   0 - 0x0
      13'h84B: dout  = 8'b00000000; // 2123 :   0 - 0x0
      13'h84C: dout  = 8'b00000000; // 2124 :   0 - 0x0
      13'h84D: dout  = 8'b00000000; // 2125 :   0 - 0x0
      13'h84E: dout  = 8'b00000000; // 2126 :   0 - 0x0
      13'h84F: dout  = 8'b00000000; // 2127 :   0 - 0x0
      13'h850: dout  = 8'b00000000; // 2128 :   0 - 0x0 -- Sprite 0x85
      13'h851: dout  = 8'b00000000; // 2129 :   0 - 0x0
      13'h852: dout  = 8'b00000000; // 2130 :   0 - 0x0
      13'h853: dout  = 8'b00000000; // 2131 :   0 - 0x0
      13'h854: dout  = 8'b00000000; // 2132 :   0 - 0x0
      13'h855: dout  = 8'b00000000; // 2133 :   0 - 0x0
      13'h856: dout  = 8'b00000000; // 2134 :   0 - 0x0
      13'h857: dout  = 8'b00000000; // 2135 :   0 - 0x0
      13'h858: dout  = 8'b00000000; // 2136 :   0 - 0x0
      13'h859: dout  = 8'b00000000; // 2137 :   0 - 0x0
      13'h85A: dout  = 8'b00000000; // 2138 :   0 - 0x0
      13'h85B: dout  = 8'b00000000; // 2139 :   0 - 0x0
      13'h85C: dout  = 8'b00000000; // 2140 :   0 - 0x0
      13'h85D: dout  = 8'b00000000; // 2141 :   0 - 0x0
      13'h85E: dout  = 8'b00000000; // 2142 :   0 - 0x0
      13'h85F: dout  = 8'b00000000; // 2143 :   0 - 0x0
      13'h860: dout  = 8'b00000000; // 2144 :   0 - 0x0 -- Sprite 0x86
      13'h861: dout  = 8'b00000000; // 2145 :   0 - 0x0
      13'h862: dout  = 8'b00000000; // 2146 :   0 - 0x0
      13'h863: dout  = 8'b00000000; // 2147 :   0 - 0x0
      13'h864: dout  = 8'b00000000; // 2148 :   0 - 0x0
      13'h865: dout  = 8'b00000000; // 2149 :   0 - 0x0
      13'h866: dout  = 8'b00000000; // 2150 :   0 - 0x0
      13'h867: dout  = 8'b00000000; // 2151 :   0 - 0x0
      13'h868: dout  = 8'b00000000; // 2152 :   0 - 0x0
      13'h869: dout  = 8'b00000000; // 2153 :   0 - 0x0
      13'h86A: dout  = 8'b00000000; // 2154 :   0 - 0x0
      13'h86B: dout  = 8'b00000000; // 2155 :   0 - 0x0
      13'h86C: dout  = 8'b00000000; // 2156 :   0 - 0x0
      13'h86D: dout  = 8'b00000000; // 2157 :   0 - 0x0
      13'h86E: dout  = 8'b00000000; // 2158 :   0 - 0x0
      13'h86F: dout  = 8'b00000000; // 2159 :   0 - 0x0
      13'h870: dout  = 8'b00000000; // 2160 :   0 - 0x0 -- Sprite 0x87
      13'h871: dout  = 8'b00000000; // 2161 :   0 - 0x0
      13'h872: dout  = 8'b00000000; // 2162 :   0 - 0x0
      13'h873: dout  = 8'b00000000; // 2163 :   0 - 0x0
      13'h874: dout  = 8'b00000000; // 2164 :   0 - 0x0
      13'h875: dout  = 8'b00000000; // 2165 :   0 - 0x0
      13'h876: dout  = 8'b00000000; // 2166 :   0 - 0x0
      13'h877: dout  = 8'b00000000; // 2167 :   0 - 0x0
      13'h878: dout  = 8'b00000000; // 2168 :   0 - 0x0
      13'h879: dout  = 8'b00000000; // 2169 :   0 - 0x0
      13'h87A: dout  = 8'b00000000; // 2170 :   0 - 0x0
      13'h87B: dout  = 8'b00000000; // 2171 :   0 - 0x0
      13'h87C: dout  = 8'b00000000; // 2172 :   0 - 0x0
      13'h87D: dout  = 8'b00000000; // 2173 :   0 - 0x0
      13'h87E: dout  = 8'b00000000; // 2174 :   0 - 0x0
      13'h87F: dout  = 8'b00000000; // 2175 :   0 - 0x0
      13'h880: dout  = 8'b00000000; // 2176 :   0 - 0x0 -- Sprite 0x88
      13'h881: dout  = 8'b00000000; // 2177 :   0 - 0x0
      13'h882: dout  = 8'b00000000; // 2178 :   0 - 0x0
      13'h883: dout  = 8'b00000000; // 2179 :   0 - 0x0
      13'h884: dout  = 8'b00000000; // 2180 :   0 - 0x0
      13'h885: dout  = 8'b00000000; // 2181 :   0 - 0x0
      13'h886: dout  = 8'b00000000; // 2182 :   0 - 0x0
      13'h887: dout  = 8'b00000000; // 2183 :   0 - 0x0
      13'h888: dout  = 8'b00000000; // 2184 :   0 - 0x0
      13'h889: dout  = 8'b00000000; // 2185 :   0 - 0x0
      13'h88A: dout  = 8'b00000000; // 2186 :   0 - 0x0
      13'h88B: dout  = 8'b00000000; // 2187 :   0 - 0x0
      13'h88C: dout  = 8'b00000000; // 2188 :   0 - 0x0
      13'h88D: dout  = 8'b00000000; // 2189 :   0 - 0x0
      13'h88E: dout  = 8'b00000000; // 2190 :   0 - 0x0
      13'h88F: dout  = 8'b00000000; // 2191 :   0 - 0x0
      13'h890: dout  = 8'b00000000; // 2192 :   0 - 0x0 -- Sprite 0x89
      13'h891: dout  = 8'b00000000; // 2193 :   0 - 0x0
      13'h892: dout  = 8'b00000000; // 2194 :   0 - 0x0
      13'h893: dout  = 8'b00000000; // 2195 :   0 - 0x0
      13'h894: dout  = 8'b00000000; // 2196 :   0 - 0x0
      13'h895: dout  = 8'b00000000; // 2197 :   0 - 0x0
      13'h896: dout  = 8'b00000000; // 2198 :   0 - 0x0
      13'h897: dout  = 8'b00000000; // 2199 :   0 - 0x0
      13'h898: dout  = 8'b00000000; // 2200 :   0 - 0x0
      13'h899: dout  = 8'b00000000; // 2201 :   0 - 0x0
      13'h89A: dout  = 8'b00000000; // 2202 :   0 - 0x0
      13'h89B: dout  = 8'b00000000; // 2203 :   0 - 0x0
      13'h89C: dout  = 8'b00000000; // 2204 :   0 - 0x0
      13'h89D: dout  = 8'b00000000; // 2205 :   0 - 0x0
      13'h89E: dout  = 8'b00000000; // 2206 :   0 - 0x0
      13'h89F: dout  = 8'b00000000; // 2207 :   0 - 0x0
      13'h8A0: dout  = 8'b00000000; // 2208 :   0 - 0x0 -- Sprite 0x8a
      13'h8A1: dout  = 8'b00000000; // 2209 :   0 - 0x0
      13'h8A2: dout  = 8'b00000000; // 2210 :   0 - 0x0
      13'h8A3: dout  = 8'b00000000; // 2211 :   0 - 0x0
      13'h8A4: dout  = 8'b00000000; // 2212 :   0 - 0x0
      13'h8A5: dout  = 8'b00000000; // 2213 :   0 - 0x0
      13'h8A6: dout  = 8'b00000000; // 2214 :   0 - 0x0
      13'h8A7: dout  = 8'b00000000; // 2215 :   0 - 0x0
      13'h8A8: dout  = 8'b00000000; // 2216 :   0 - 0x0
      13'h8A9: dout  = 8'b00000000; // 2217 :   0 - 0x0
      13'h8AA: dout  = 8'b00000000; // 2218 :   0 - 0x0
      13'h8AB: dout  = 8'b00000000; // 2219 :   0 - 0x0
      13'h8AC: dout  = 8'b00000000; // 2220 :   0 - 0x0
      13'h8AD: dout  = 8'b00000000; // 2221 :   0 - 0x0
      13'h8AE: dout  = 8'b00000000; // 2222 :   0 - 0x0
      13'h8AF: dout  = 8'b00000000; // 2223 :   0 - 0x0
      13'h8B0: dout  = 8'b00000000; // 2224 :   0 - 0x0 -- Sprite 0x8b
      13'h8B1: dout  = 8'b00000000; // 2225 :   0 - 0x0
      13'h8B2: dout  = 8'b00000000; // 2226 :   0 - 0x0
      13'h8B3: dout  = 8'b00000000; // 2227 :   0 - 0x0
      13'h8B4: dout  = 8'b00000000; // 2228 :   0 - 0x0
      13'h8B5: dout  = 8'b00000000; // 2229 :   0 - 0x0
      13'h8B6: dout  = 8'b00000000; // 2230 :   0 - 0x0
      13'h8B7: dout  = 8'b00000000; // 2231 :   0 - 0x0
      13'h8B8: dout  = 8'b00000000; // 2232 :   0 - 0x0
      13'h8B9: dout  = 8'b00000000; // 2233 :   0 - 0x0
      13'h8BA: dout  = 8'b00000000; // 2234 :   0 - 0x0
      13'h8BB: dout  = 8'b00000000; // 2235 :   0 - 0x0
      13'h8BC: dout  = 8'b00000000; // 2236 :   0 - 0x0
      13'h8BD: dout  = 8'b00000000; // 2237 :   0 - 0x0
      13'h8BE: dout  = 8'b00000000; // 2238 :   0 - 0x0
      13'h8BF: dout  = 8'b00000000; // 2239 :   0 - 0x0
      13'h8C0: dout  = 8'b00000000; // 2240 :   0 - 0x0 -- Sprite 0x8c
      13'h8C1: dout  = 8'b00000000; // 2241 :   0 - 0x0
      13'h8C2: dout  = 8'b00000000; // 2242 :   0 - 0x0
      13'h8C3: dout  = 8'b00000000; // 2243 :   0 - 0x0
      13'h8C4: dout  = 8'b00000000; // 2244 :   0 - 0x0
      13'h8C5: dout  = 8'b00000000; // 2245 :   0 - 0x0
      13'h8C6: dout  = 8'b00000000; // 2246 :   0 - 0x0
      13'h8C7: dout  = 8'b00000000; // 2247 :   0 - 0x0
      13'h8C8: dout  = 8'b00000000; // 2248 :   0 - 0x0
      13'h8C9: dout  = 8'b00000000; // 2249 :   0 - 0x0
      13'h8CA: dout  = 8'b00000000; // 2250 :   0 - 0x0
      13'h8CB: dout  = 8'b00000000; // 2251 :   0 - 0x0
      13'h8CC: dout  = 8'b00000000; // 2252 :   0 - 0x0
      13'h8CD: dout  = 8'b00000000; // 2253 :   0 - 0x0
      13'h8CE: dout  = 8'b00000000; // 2254 :   0 - 0x0
      13'h8CF: dout  = 8'b00000000; // 2255 :   0 - 0x0
      13'h8D0: dout  = 8'b00000000; // 2256 :   0 - 0x0 -- Sprite 0x8d
      13'h8D1: dout  = 8'b00000000; // 2257 :   0 - 0x0
      13'h8D2: dout  = 8'b00000000; // 2258 :   0 - 0x0
      13'h8D3: dout  = 8'b00000000; // 2259 :   0 - 0x0
      13'h8D4: dout  = 8'b00000000; // 2260 :   0 - 0x0
      13'h8D5: dout  = 8'b00000000; // 2261 :   0 - 0x0
      13'h8D6: dout  = 8'b00000000; // 2262 :   0 - 0x0
      13'h8D7: dout  = 8'b00000000; // 2263 :   0 - 0x0
      13'h8D8: dout  = 8'b00000000; // 2264 :   0 - 0x0
      13'h8D9: dout  = 8'b00000000; // 2265 :   0 - 0x0
      13'h8DA: dout  = 8'b00000000; // 2266 :   0 - 0x0
      13'h8DB: dout  = 8'b00000000; // 2267 :   0 - 0x0
      13'h8DC: dout  = 8'b00000000; // 2268 :   0 - 0x0
      13'h8DD: dout  = 8'b00000000; // 2269 :   0 - 0x0
      13'h8DE: dout  = 8'b00000000; // 2270 :   0 - 0x0
      13'h8DF: dout  = 8'b00000000; // 2271 :   0 - 0x0
      13'h8E0: dout  = 8'b00000000; // 2272 :   0 - 0x0 -- Sprite 0x8e
      13'h8E1: dout  = 8'b00000000; // 2273 :   0 - 0x0
      13'h8E2: dout  = 8'b00000000; // 2274 :   0 - 0x0
      13'h8E3: dout  = 8'b00000000; // 2275 :   0 - 0x0
      13'h8E4: dout  = 8'b00000000; // 2276 :   0 - 0x0
      13'h8E5: dout  = 8'b00000000; // 2277 :   0 - 0x0
      13'h8E6: dout  = 8'b00000000; // 2278 :   0 - 0x0
      13'h8E7: dout  = 8'b00000000; // 2279 :   0 - 0x0
      13'h8E8: dout  = 8'b00000000; // 2280 :   0 - 0x0
      13'h8E9: dout  = 8'b00000000; // 2281 :   0 - 0x0
      13'h8EA: dout  = 8'b00000000; // 2282 :   0 - 0x0
      13'h8EB: dout  = 8'b00000000; // 2283 :   0 - 0x0
      13'h8EC: dout  = 8'b00000000; // 2284 :   0 - 0x0
      13'h8ED: dout  = 8'b00000000; // 2285 :   0 - 0x0
      13'h8EE: dout  = 8'b00000000; // 2286 :   0 - 0x0
      13'h8EF: dout  = 8'b00000000; // 2287 :   0 - 0x0
      13'h8F0: dout  = 8'b00000000; // 2288 :   0 - 0x0 -- Sprite 0x8f
      13'h8F1: dout  = 8'b00000000; // 2289 :   0 - 0x0
      13'h8F2: dout  = 8'b00000000; // 2290 :   0 - 0x0
      13'h8F3: dout  = 8'b00000000; // 2291 :   0 - 0x0
      13'h8F4: dout  = 8'b00000000; // 2292 :   0 - 0x0
      13'h8F5: dout  = 8'b00000000; // 2293 :   0 - 0x0
      13'h8F6: dout  = 8'b00000000; // 2294 :   0 - 0x0
      13'h8F7: dout  = 8'b00000000; // 2295 :   0 - 0x0
      13'h8F8: dout  = 8'b00000000; // 2296 :   0 - 0x0
      13'h8F9: dout  = 8'b00000000; // 2297 :   0 - 0x0
      13'h8FA: dout  = 8'b00000000; // 2298 :   0 - 0x0
      13'h8FB: dout  = 8'b00000000; // 2299 :   0 - 0x0
      13'h8FC: dout  = 8'b00000000; // 2300 :   0 - 0x0
      13'h8FD: dout  = 8'b00000000; // 2301 :   0 - 0x0
      13'h8FE: dout  = 8'b00000000; // 2302 :   0 - 0x0
      13'h8FF: dout  = 8'b00000000; // 2303 :   0 - 0x0
      13'h900: dout  = 8'b00000000; // 2304 :   0 - 0x0 -- Sprite 0x90
      13'h901: dout  = 8'b00000000; // 2305 :   0 - 0x0
      13'h902: dout  = 8'b00000000; // 2306 :   0 - 0x0
      13'h903: dout  = 8'b00000000; // 2307 :   0 - 0x0
      13'h904: dout  = 8'b00000000; // 2308 :   0 - 0x0
      13'h905: dout  = 8'b00000000; // 2309 :   0 - 0x0
      13'h906: dout  = 8'b00000000; // 2310 :   0 - 0x0
      13'h907: dout  = 8'b00000000; // 2311 :   0 - 0x0
      13'h908: dout  = 8'b00000000; // 2312 :   0 - 0x0
      13'h909: dout  = 8'b00000000; // 2313 :   0 - 0x0
      13'h90A: dout  = 8'b00000000; // 2314 :   0 - 0x0
      13'h90B: dout  = 8'b00000000; // 2315 :   0 - 0x0
      13'h90C: dout  = 8'b00000000; // 2316 :   0 - 0x0
      13'h90D: dout  = 8'b00000000; // 2317 :   0 - 0x0
      13'h90E: dout  = 8'b00000000; // 2318 :   0 - 0x0
      13'h90F: dout  = 8'b00000000; // 2319 :   0 - 0x0
      13'h910: dout  = 8'b00000000; // 2320 :   0 - 0x0 -- Sprite 0x91
      13'h911: dout  = 8'b00000000; // 2321 :   0 - 0x0
      13'h912: dout  = 8'b00000000; // 2322 :   0 - 0x0
      13'h913: dout  = 8'b00000000; // 2323 :   0 - 0x0
      13'h914: dout  = 8'b00000000; // 2324 :   0 - 0x0
      13'h915: dout  = 8'b00000000; // 2325 :   0 - 0x0
      13'h916: dout  = 8'b00000000; // 2326 :   0 - 0x0
      13'h917: dout  = 8'b00000000; // 2327 :   0 - 0x0
      13'h918: dout  = 8'b00000000; // 2328 :   0 - 0x0
      13'h919: dout  = 8'b00000000; // 2329 :   0 - 0x0
      13'h91A: dout  = 8'b00000000; // 2330 :   0 - 0x0
      13'h91B: dout  = 8'b00000000; // 2331 :   0 - 0x0
      13'h91C: dout  = 8'b00000000; // 2332 :   0 - 0x0
      13'h91D: dout  = 8'b00000000; // 2333 :   0 - 0x0
      13'h91E: dout  = 8'b00000000; // 2334 :   0 - 0x0
      13'h91F: dout  = 8'b00000000; // 2335 :   0 - 0x0
      13'h920: dout  = 8'b00000000; // 2336 :   0 - 0x0 -- Sprite 0x92
      13'h921: dout  = 8'b00000000; // 2337 :   0 - 0x0
      13'h922: dout  = 8'b00000000; // 2338 :   0 - 0x0
      13'h923: dout  = 8'b00000000; // 2339 :   0 - 0x0
      13'h924: dout  = 8'b00000000; // 2340 :   0 - 0x0
      13'h925: dout  = 8'b00000000; // 2341 :   0 - 0x0
      13'h926: dout  = 8'b00000000; // 2342 :   0 - 0x0
      13'h927: dout  = 8'b00000000; // 2343 :   0 - 0x0
      13'h928: dout  = 8'b00000000; // 2344 :   0 - 0x0
      13'h929: dout  = 8'b00000000; // 2345 :   0 - 0x0
      13'h92A: dout  = 8'b00000000; // 2346 :   0 - 0x0
      13'h92B: dout  = 8'b00000000; // 2347 :   0 - 0x0
      13'h92C: dout  = 8'b00000000; // 2348 :   0 - 0x0
      13'h92D: dout  = 8'b00000000; // 2349 :   0 - 0x0
      13'h92E: dout  = 8'b00000000; // 2350 :   0 - 0x0
      13'h92F: dout  = 8'b00000000; // 2351 :   0 - 0x0
      13'h930: dout  = 8'b00000000; // 2352 :   0 - 0x0 -- Sprite 0x93
      13'h931: dout  = 8'b00000000; // 2353 :   0 - 0x0
      13'h932: dout  = 8'b00000000; // 2354 :   0 - 0x0
      13'h933: dout  = 8'b00000000; // 2355 :   0 - 0x0
      13'h934: dout  = 8'b00000000; // 2356 :   0 - 0x0
      13'h935: dout  = 8'b00000000; // 2357 :   0 - 0x0
      13'h936: dout  = 8'b00000000; // 2358 :   0 - 0x0
      13'h937: dout  = 8'b00000000; // 2359 :   0 - 0x0
      13'h938: dout  = 8'b00000000; // 2360 :   0 - 0x0
      13'h939: dout  = 8'b00000000; // 2361 :   0 - 0x0
      13'h93A: dout  = 8'b00000000; // 2362 :   0 - 0x0
      13'h93B: dout  = 8'b00000000; // 2363 :   0 - 0x0
      13'h93C: dout  = 8'b00000000; // 2364 :   0 - 0x0
      13'h93D: dout  = 8'b00000000; // 2365 :   0 - 0x0
      13'h93E: dout  = 8'b00000000; // 2366 :   0 - 0x0
      13'h93F: dout  = 8'b00000000; // 2367 :   0 - 0x0
      13'h940: dout  = 8'b00000000; // 2368 :   0 - 0x0 -- Sprite 0x94
      13'h941: dout  = 8'b00000000; // 2369 :   0 - 0x0
      13'h942: dout  = 8'b00000000; // 2370 :   0 - 0x0
      13'h943: dout  = 8'b00000000; // 2371 :   0 - 0x0
      13'h944: dout  = 8'b00000000; // 2372 :   0 - 0x0
      13'h945: dout  = 8'b00000000; // 2373 :   0 - 0x0
      13'h946: dout  = 8'b00000000; // 2374 :   0 - 0x0
      13'h947: dout  = 8'b00000000; // 2375 :   0 - 0x0
      13'h948: dout  = 8'b00000000; // 2376 :   0 - 0x0
      13'h949: dout  = 8'b00000000; // 2377 :   0 - 0x0
      13'h94A: dout  = 8'b00000000; // 2378 :   0 - 0x0
      13'h94B: dout  = 8'b00000000; // 2379 :   0 - 0x0
      13'h94C: dout  = 8'b00000000; // 2380 :   0 - 0x0
      13'h94D: dout  = 8'b00000000; // 2381 :   0 - 0x0
      13'h94E: dout  = 8'b00000000; // 2382 :   0 - 0x0
      13'h94F: dout  = 8'b00000000; // 2383 :   0 - 0x0
      13'h950: dout  = 8'b00000000; // 2384 :   0 - 0x0 -- Sprite 0x95
      13'h951: dout  = 8'b00000000; // 2385 :   0 - 0x0
      13'h952: dout  = 8'b00000000; // 2386 :   0 - 0x0
      13'h953: dout  = 8'b00000000; // 2387 :   0 - 0x0
      13'h954: dout  = 8'b00000000; // 2388 :   0 - 0x0
      13'h955: dout  = 8'b00000000; // 2389 :   0 - 0x0
      13'h956: dout  = 8'b00000000; // 2390 :   0 - 0x0
      13'h957: dout  = 8'b00000000; // 2391 :   0 - 0x0
      13'h958: dout  = 8'b00000000; // 2392 :   0 - 0x0
      13'h959: dout  = 8'b00000000; // 2393 :   0 - 0x0
      13'h95A: dout  = 8'b00000000; // 2394 :   0 - 0x0
      13'h95B: dout  = 8'b00000000; // 2395 :   0 - 0x0
      13'h95C: dout  = 8'b00000000; // 2396 :   0 - 0x0
      13'h95D: dout  = 8'b00000000; // 2397 :   0 - 0x0
      13'h95E: dout  = 8'b00000000; // 2398 :   0 - 0x0
      13'h95F: dout  = 8'b00000000; // 2399 :   0 - 0x0
      13'h960: dout  = 8'b00000000; // 2400 :   0 - 0x0 -- Sprite 0x96
      13'h961: dout  = 8'b00000000; // 2401 :   0 - 0x0
      13'h962: dout  = 8'b00000000; // 2402 :   0 - 0x0
      13'h963: dout  = 8'b00000000; // 2403 :   0 - 0x0
      13'h964: dout  = 8'b00000000; // 2404 :   0 - 0x0
      13'h965: dout  = 8'b00000000; // 2405 :   0 - 0x0
      13'h966: dout  = 8'b00000000; // 2406 :   0 - 0x0
      13'h967: dout  = 8'b00000000; // 2407 :   0 - 0x0
      13'h968: dout  = 8'b00000000; // 2408 :   0 - 0x0
      13'h969: dout  = 8'b00000000; // 2409 :   0 - 0x0
      13'h96A: dout  = 8'b00000000; // 2410 :   0 - 0x0
      13'h96B: dout  = 8'b00000000; // 2411 :   0 - 0x0
      13'h96C: dout  = 8'b00000000; // 2412 :   0 - 0x0
      13'h96D: dout  = 8'b00000000; // 2413 :   0 - 0x0
      13'h96E: dout  = 8'b00000000; // 2414 :   0 - 0x0
      13'h96F: dout  = 8'b00000000; // 2415 :   0 - 0x0
      13'h970: dout  = 8'b00000000; // 2416 :   0 - 0x0 -- Sprite 0x97
      13'h971: dout  = 8'b00000000; // 2417 :   0 - 0x0
      13'h972: dout  = 8'b00000000; // 2418 :   0 - 0x0
      13'h973: dout  = 8'b00000000; // 2419 :   0 - 0x0
      13'h974: dout  = 8'b00000000; // 2420 :   0 - 0x0
      13'h975: dout  = 8'b00000000; // 2421 :   0 - 0x0
      13'h976: dout  = 8'b00000000; // 2422 :   0 - 0x0
      13'h977: dout  = 8'b00000000; // 2423 :   0 - 0x0
      13'h978: dout  = 8'b00000000; // 2424 :   0 - 0x0
      13'h979: dout  = 8'b00000000; // 2425 :   0 - 0x0
      13'h97A: dout  = 8'b00000000; // 2426 :   0 - 0x0
      13'h97B: dout  = 8'b00000000; // 2427 :   0 - 0x0
      13'h97C: dout  = 8'b00000000; // 2428 :   0 - 0x0
      13'h97D: dout  = 8'b00000000; // 2429 :   0 - 0x0
      13'h97E: dout  = 8'b00000000; // 2430 :   0 - 0x0
      13'h97F: dout  = 8'b00000000; // 2431 :   0 - 0x0
      13'h980: dout  = 8'b00000000; // 2432 :   0 - 0x0 -- Sprite 0x98
      13'h981: dout  = 8'b00000000; // 2433 :   0 - 0x0
      13'h982: dout  = 8'b00000000; // 2434 :   0 - 0x0
      13'h983: dout  = 8'b00000000; // 2435 :   0 - 0x0
      13'h984: dout  = 8'b00000000; // 2436 :   0 - 0x0
      13'h985: dout  = 8'b00000000; // 2437 :   0 - 0x0
      13'h986: dout  = 8'b00000000; // 2438 :   0 - 0x0
      13'h987: dout  = 8'b00000000; // 2439 :   0 - 0x0
      13'h988: dout  = 8'b00000000; // 2440 :   0 - 0x0
      13'h989: dout  = 8'b00000000; // 2441 :   0 - 0x0
      13'h98A: dout  = 8'b00000000; // 2442 :   0 - 0x0
      13'h98B: dout  = 8'b00000000; // 2443 :   0 - 0x0
      13'h98C: dout  = 8'b00000000; // 2444 :   0 - 0x0
      13'h98D: dout  = 8'b00000000; // 2445 :   0 - 0x0
      13'h98E: dout  = 8'b00000000; // 2446 :   0 - 0x0
      13'h98F: dout  = 8'b00000000; // 2447 :   0 - 0x0
      13'h990: dout  = 8'b00000000; // 2448 :   0 - 0x0 -- Sprite 0x99
      13'h991: dout  = 8'b00000000; // 2449 :   0 - 0x0
      13'h992: dout  = 8'b00000000; // 2450 :   0 - 0x0
      13'h993: dout  = 8'b00000000; // 2451 :   0 - 0x0
      13'h994: dout  = 8'b00000000; // 2452 :   0 - 0x0
      13'h995: dout  = 8'b00000000; // 2453 :   0 - 0x0
      13'h996: dout  = 8'b00000000; // 2454 :   0 - 0x0
      13'h997: dout  = 8'b00000000; // 2455 :   0 - 0x0
      13'h998: dout  = 8'b00000000; // 2456 :   0 - 0x0
      13'h999: dout  = 8'b00000000; // 2457 :   0 - 0x0
      13'h99A: dout  = 8'b00000000; // 2458 :   0 - 0x0
      13'h99B: dout  = 8'b00000000; // 2459 :   0 - 0x0
      13'h99C: dout  = 8'b00000000; // 2460 :   0 - 0x0
      13'h99D: dout  = 8'b00000000; // 2461 :   0 - 0x0
      13'h99E: dout  = 8'b00000000; // 2462 :   0 - 0x0
      13'h99F: dout  = 8'b00000000; // 2463 :   0 - 0x0
      13'h9A0: dout  = 8'b00000000; // 2464 :   0 - 0x0 -- Sprite 0x9a
      13'h9A1: dout  = 8'b00000000; // 2465 :   0 - 0x0
      13'h9A2: dout  = 8'b00000000; // 2466 :   0 - 0x0
      13'h9A3: dout  = 8'b00000000; // 2467 :   0 - 0x0
      13'h9A4: dout  = 8'b00000000; // 2468 :   0 - 0x0
      13'h9A5: dout  = 8'b00000000; // 2469 :   0 - 0x0
      13'h9A6: dout  = 8'b00000000; // 2470 :   0 - 0x0
      13'h9A7: dout  = 8'b00000000; // 2471 :   0 - 0x0
      13'h9A8: dout  = 8'b00000000; // 2472 :   0 - 0x0
      13'h9A9: dout  = 8'b00000000; // 2473 :   0 - 0x0
      13'h9AA: dout  = 8'b00000000; // 2474 :   0 - 0x0
      13'h9AB: dout  = 8'b00000000; // 2475 :   0 - 0x0
      13'h9AC: dout  = 8'b00000000; // 2476 :   0 - 0x0
      13'h9AD: dout  = 8'b00000000; // 2477 :   0 - 0x0
      13'h9AE: dout  = 8'b00000000; // 2478 :   0 - 0x0
      13'h9AF: dout  = 8'b00000000; // 2479 :   0 - 0x0
      13'h9B0: dout  = 8'b00000000; // 2480 :   0 - 0x0 -- Sprite 0x9b
      13'h9B1: dout  = 8'b00000000; // 2481 :   0 - 0x0
      13'h9B2: dout  = 8'b00000000; // 2482 :   0 - 0x0
      13'h9B3: dout  = 8'b00000000; // 2483 :   0 - 0x0
      13'h9B4: dout  = 8'b00000000; // 2484 :   0 - 0x0
      13'h9B5: dout  = 8'b00000000; // 2485 :   0 - 0x0
      13'h9B6: dout  = 8'b00000000; // 2486 :   0 - 0x0
      13'h9B7: dout  = 8'b00000000; // 2487 :   0 - 0x0
      13'h9B8: dout  = 8'b00000000; // 2488 :   0 - 0x0
      13'h9B9: dout  = 8'b00000000; // 2489 :   0 - 0x0
      13'h9BA: dout  = 8'b00000000; // 2490 :   0 - 0x0
      13'h9BB: dout  = 8'b00000000; // 2491 :   0 - 0x0
      13'h9BC: dout  = 8'b00000000; // 2492 :   0 - 0x0
      13'h9BD: dout  = 8'b00000000; // 2493 :   0 - 0x0
      13'h9BE: dout  = 8'b00000000; // 2494 :   0 - 0x0
      13'h9BF: dout  = 8'b00000000; // 2495 :   0 - 0x0
      13'h9C0: dout  = 8'b00000000; // 2496 :   0 - 0x0 -- Sprite 0x9c
      13'h9C1: dout  = 8'b00000000; // 2497 :   0 - 0x0
      13'h9C2: dout  = 8'b00000000; // 2498 :   0 - 0x0
      13'h9C3: dout  = 8'b00000000; // 2499 :   0 - 0x0
      13'h9C4: dout  = 8'b00000000; // 2500 :   0 - 0x0
      13'h9C5: dout  = 8'b00000000; // 2501 :   0 - 0x0
      13'h9C6: dout  = 8'b00000000; // 2502 :   0 - 0x0
      13'h9C7: dout  = 8'b00000000; // 2503 :   0 - 0x0
      13'h9C8: dout  = 8'b00000000; // 2504 :   0 - 0x0
      13'h9C9: dout  = 8'b00000000; // 2505 :   0 - 0x0
      13'h9CA: dout  = 8'b00000000; // 2506 :   0 - 0x0
      13'h9CB: dout  = 8'b00000000; // 2507 :   0 - 0x0
      13'h9CC: dout  = 8'b00000000; // 2508 :   0 - 0x0
      13'h9CD: dout  = 8'b00000000; // 2509 :   0 - 0x0
      13'h9CE: dout  = 8'b00000000; // 2510 :   0 - 0x0
      13'h9CF: dout  = 8'b00000000; // 2511 :   0 - 0x0
      13'h9D0: dout  = 8'b00000000; // 2512 :   0 - 0x0 -- Sprite 0x9d
      13'h9D1: dout  = 8'b00000000; // 2513 :   0 - 0x0
      13'h9D2: dout  = 8'b00000000; // 2514 :   0 - 0x0
      13'h9D3: dout  = 8'b00000000; // 2515 :   0 - 0x0
      13'h9D4: dout  = 8'b00000000; // 2516 :   0 - 0x0
      13'h9D5: dout  = 8'b00000000; // 2517 :   0 - 0x0
      13'h9D6: dout  = 8'b00000000; // 2518 :   0 - 0x0
      13'h9D7: dout  = 8'b00000000; // 2519 :   0 - 0x0
      13'h9D8: dout  = 8'b00000000; // 2520 :   0 - 0x0
      13'h9D9: dout  = 8'b00000000; // 2521 :   0 - 0x0
      13'h9DA: dout  = 8'b00000000; // 2522 :   0 - 0x0
      13'h9DB: dout  = 8'b00000000; // 2523 :   0 - 0x0
      13'h9DC: dout  = 8'b00000000; // 2524 :   0 - 0x0
      13'h9DD: dout  = 8'b00000000; // 2525 :   0 - 0x0
      13'h9DE: dout  = 8'b00000000; // 2526 :   0 - 0x0
      13'h9DF: dout  = 8'b00000000; // 2527 :   0 - 0x0
      13'h9E0: dout  = 8'b00000000; // 2528 :   0 - 0x0 -- Sprite 0x9e
      13'h9E1: dout  = 8'b00000000; // 2529 :   0 - 0x0
      13'h9E2: dout  = 8'b00000000; // 2530 :   0 - 0x0
      13'h9E3: dout  = 8'b00000000; // 2531 :   0 - 0x0
      13'h9E4: dout  = 8'b00000000; // 2532 :   0 - 0x0
      13'h9E5: dout  = 8'b00000000; // 2533 :   0 - 0x0
      13'h9E6: dout  = 8'b00000000; // 2534 :   0 - 0x0
      13'h9E7: dout  = 8'b00000000; // 2535 :   0 - 0x0
      13'h9E8: dout  = 8'b00000000; // 2536 :   0 - 0x0
      13'h9E9: dout  = 8'b00000000; // 2537 :   0 - 0x0
      13'h9EA: dout  = 8'b00000000; // 2538 :   0 - 0x0
      13'h9EB: dout  = 8'b00000000; // 2539 :   0 - 0x0
      13'h9EC: dout  = 8'b00000000; // 2540 :   0 - 0x0
      13'h9ED: dout  = 8'b00000000; // 2541 :   0 - 0x0
      13'h9EE: dout  = 8'b00000000; // 2542 :   0 - 0x0
      13'h9EF: dout  = 8'b00000000; // 2543 :   0 - 0x0
      13'h9F0: dout  = 8'b00000000; // 2544 :   0 - 0x0 -- Sprite 0x9f
      13'h9F1: dout  = 8'b00000000; // 2545 :   0 - 0x0
      13'h9F2: dout  = 8'b00000000; // 2546 :   0 - 0x0
      13'h9F3: dout  = 8'b00000000; // 2547 :   0 - 0x0
      13'h9F4: dout  = 8'b00000000; // 2548 :   0 - 0x0
      13'h9F5: dout  = 8'b00000000; // 2549 :   0 - 0x0
      13'h9F6: dout  = 8'b00000000; // 2550 :   0 - 0x0
      13'h9F7: dout  = 8'b00000000; // 2551 :   0 - 0x0
      13'h9F8: dout  = 8'b00000000; // 2552 :   0 - 0x0
      13'h9F9: dout  = 8'b00000000; // 2553 :   0 - 0x0
      13'h9FA: dout  = 8'b00000000; // 2554 :   0 - 0x0
      13'h9FB: dout  = 8'b00000000; // 2555 :   0 - 0x0
      13'h9FC: dout  = 8'b00000000; // 2556 :   0 - 0x0
      13'h9FD: dout  = 8'b00000000; // 2557 :   0 - 0x0
      13'h9FE: dout  = 8'b00000000; // 2558 :   0 - 0x0
      13'h9FF: dout  = 8'b00000000; // 2559 :   0 - 0x0
      13'hA00: dout  = 8'b00000000; // 2560 :   0 - 0x0 -- Sprite 0xa0
      13'hA01: dout  = 8'b00000000; // 2561 :   0 - 0x0
      13'hA02: dout  = 8'b00000000; // 2562 :   0 - 0x0
      13'hA03: dout  = 8'b00000000; // 2563 :   0 - 0x0
      13'hA04: dout  = 8'b00000000; // 2564 :   0 - 0x0
      13'hA05: dout  = 8'b00000000; // 2565 :   0 - 0x0
      13'hA06: dout  = 8'b00000000; // 2566 :   0 - 0x0
      13'hA07: dout  = 8'b00000000; // 2567 :   0 - 0x0
      13'hA08: dout  = 8'b00000000; // 2568 :   0 - 0x0
      13'hA09: dout  = 8'b00000000; // 2569 :   0 - 0x0
      13'hA0A: dout  = 8'b00000000; // 2570 :   0 - 0x0
      13'hA0B: dout  = 8'b00000000; // 2571 :   0 - 0x0
      13'hA0C: dout  = 8'b00000000; // 2572 :   0 - 0x0
      13'hA0D: dout  = 8'b00000000; // 2573 :   0 - 0x0
      13'hA0E: dout  = 8'b00000000; // 2574 :   0 - 0x0
      13'hA0F: dout  = 8'b00000000; // 2575 :   0 - 0x0
      13'hA10: dout  = 8'b00000000; // 2576 :   0 - 0x0 -- Sprite 0xa1
      13'hA11: dout  = 8'b00000000; // 2577 :   0 - 0x0
      13'hA12: dout  = 8'b00000000; // 2578 :   0 - 0x0
      13'hA13: dout  = 8'b00000000; // 2579 :   0 - 0x0
      13'hA14: dout  = 8'b00000000; // 2580 :   0 - 0x0
      13'hA15: dout  = 8'b00000000; // 2581 :   0 - 0x0
      13'hA16: dout  = 8'b00000000; // 2582 :   0 - 0x0
      13'hA17: dout  = 8'b00000000; // 2583 :   0 - 0x0
      13'hA18: dout  = 8'b00000000; // 2584 :   0 - 0x0
      13'hA19: dout  = 8'b00000000; // 2585 :   0 - 0x0
      13'hA1A: dout  = 8'b00000000; // 2586 :   0 - 0x0
      13'hA1B: dout  = 8'b00000000; // 2587 :   0 - 0x0
      13'hA1C: dout  = 8'b00000000; // 2588 :   0 - 0x0
      13'hA1D: dout  = 8'b00000000; // 2589 :   0 - 0x0
      13'hA1E: dout  = 8'b00000000; // 2590 :   0 - 0x0
      13'hA1F: dout  = 8'b00000000; // 2591 :   0 - 0x0
      13'hA20: dout  = 8'b00000000; // 2592 :   0 - 0x0 -- Sprite 0xa2
      13'hA21: dout  = 8'b00000000; // 2593 :   0 - 0x0
      13'hA22: dout  = 8'b00000000; // 2594 :   0 - 0x0
      13'hA23: dout  = 8'b00000000; // 2595 :   0 - 0x0
      13'hA24: dout  = 8'b00000000; // 2596 :   0 - 0x0
      13'hA25: dout  = 8'b00000000; // 2597 :   0 - 0x0
      13'hA26: dout  = 8'b00000000; // 2598 :   0 - 0x0
      13'hA27: dout  = 8'b00000000; // 2599 :   0 - 0x0
      13'hA28: dout  = 8'b00000000; // 2600 :   0 - 0x0
      13'hA29: dout  = 8'b00000000; // 2601 :   0 - 0x0
      13'hA2A: dout  = 8'b00000000; // 2602 :   0 - 0x0
      13'hA2B: dout  = 8'b00000000; // 2603 :   0 - 0x0
      13'hA2C: dout  = 8'b00000000; // 2604 :   0 - 0x0
      13'hA2D: dout  = 8'b00000000; // 2605 :   0 - 0x0
      13'hA2E: dout  = 8'b00000000; // 2606 :   0 - 0x0
      13'hA2F: dout  = 8'b00000000; // 2607 :   0 - 0x0
      13'hA30: dout  = 8'b00000000; // 2608 :   0 - 0x0 -- Sprite 0xa3
      13'hA31: dout  = 8'b00000000; // 2609 :   0 - 0x0
      13'hA32: dout  = 8'b00000000; // 2610 :   0 - 0x0
      13'hA33: dout  = 8'b00000000; // 2611 :   0 - 0x0
      13'hA34: dout  = 8'b00000000; // 2612 :   0 - 0x0
      13'hA35: dout  = 8'b00000000; // 2613 :   0 - 0x0
      13'hA36: dout  = 8'b00000000; // 2614 :   0 - 0x0
      13'hA37: dout  = 8'b00000000; // 2615 :   0 - 0x0
      13'hA38: dout  = 8'b00000000; // 2616 :   0 - 0x0
      13'hA39: dout  = 8'b00000000; // 2617 :   0 - 0x0
      13'hA3A: dout  = 8'b00000000; // 2618 :   0 - 0x0
      13'hA3B: dout  = 8'b00000000; // 2619 :   0 - 0x0
      13'hA3C: dout  = 8'b00000000; // 2620 :   0 - 0x0
      13'hA3D: dout  = 8'b00000000; // 2621 :   0 - 0x0
      13'hA3E: dout  = 8'b00000000; // 2622 :   0 - 0x0
      13'hA3F: dout  = 8'b00000000; // 2623 :   0 - 0x0
      13'hA40: dout  = 8'b00000000; // 2624 :   0 - 0x0 -- Sprite 0xa4
      13'hA41: dout  = 8'b00000000; // 2625 :   0 - 0x0
      13'hA42: dout  = 8'b00000000; // 2626 :   0 - 0x0
      13'hA43: dout  = 8'b00000000; // 2627 :   0 - 0x0
      13'hA44: dout  = 8'b00000000; // 2628 :   0 - 0x0
      13'hA45: dout  = 8'b00000000; // 2629 :   0 - 0x0
      13'hA46: dout  = 8'b00000000; // 2630 :   0 - 0x0
      13'hA47: dout  = 8'b00000000; // 2631 :   0 - 0x0
      13'hA48: dout  = 8'b00000000; // 2632 :   0 - 0x0
      13'hA49: dout  = 8'b00000000; // 2633 :   0 - 0x0
      13'hA4A: dout  = 8'b00000000; // 2634 :   0 - 0x0
      13'hA4B: dout  = 8'b00000000; // 2635 :   0 - 0x0
      13'hA4C: dout  = 8'b00000000; // 2636 :   0 - 0x0
      13'hA4D: dout  = 8'b00000000; // 2637 :   0 - 0x0
      13'hA4E: dout  = 8'b00000000; // 2638 :   0 - 0x0
      13'hA4F: dout  = 8'b00000000; // 2639 :   0 - 0x0
      13'hA50: dout  = 8'b00000000; // 2640 :   0 - 0x0 -- Sprite 0xa5
      13'hA51: dout  = 8'b00000000; // 2641 :   0 - 0x0
      13'hA52: dout  = 8'b00000000; // 2642 :   0 - 0x0
      13'hA53: dout  = 8'b00000000; // 2643 :   0 - 0x0
      13'hA54: dout  = 8'b00000000; // 2644 :   0 - 0x0
      13'hA55: dout  = 8'b00000000; // 2645 :   0 - 0x0
      13'hA56: dout  = 8'b00000000; // 2646 :   0 - 0x0
      13'hA57: dout  = 8'b00000000; // 2647 :   0 - 0x0
      13'hA58: dout  = 8'b00000000; // 2648 :   0 - 0x0
      13'hA59: dout  = 8'b00000000; // 2649 :   0 - 0x0
      13'hA5A: dout  = 8'b00000000; // 2650 :   0 - 0x0
      13'hA5B: dout  = 8'b00000000; // 2651 :   0 - 0x0
      13'hA5C: dout  = 8'b00000000; // 2652 :   0 - 0x0
      13'hA5D: dout  = 8'b00000000; // 2653 :   0 - 0x0
      13'hA5E: dout  = 8'b00000000; // 2654 :   0 - 0x0
      13'hA5F: dout  = 8'b00000000; // 2655 :   0 - 0x0
      13'hA60: dout  = 8'b00000000; // 2656 :   0 - 0x0 -- Sprite 0xa6
      13'hA61: dout  = 8'b00000000; // 2657 :   0 - 0x0
      13'hA62: dout  = 8'b00000000; // 2658 :   0 - 0x0
      13'hA63: dout  = 8'b00000000; // 2659 :   0 - 0x0
      13'hA64: dout  = 8'b00000000; // 2660 :   0 - 0x0
      13'hA65: dout  = 8'b00000000; // 2661 :   0 - 0x0
      13'hA66: dout  = 8'b00000000; // 2662 :   0 - 0x0
      13'hA67: dout  = 8'b00000000; // 2663 :   0 - 0x0
      13'hA68: dout  = 8'b00000000; // 2664 :   0 - 0x0
      13'hA69: dout  = 8'b00000000; // 2665 :   0 - 0x0
      13'hA6A: dout  = 8'b00000000; // 2666 :   0 - 0x0
      13'hA6B: dout  = 8'b00000000; // 2667 :   0 - 0x0
      13'hA6C: dout  = 8'b00000000; // 2668 :   0 - 0x0
      13'hA6D: dout  = 8'b00000000; // 2669 :   0 - 0x0
      13'hA6E: dout  = 8'b00000000; // 2670 :   0 - 0x0
      13'hA6F: dout  = 8'b00000000; // 2671 :   0 - 0x0
      13'hA70: dout  = 8'b00000000; // 2672 :   0 - 0x0 -- Sprite 0xa7
      13'hA71: dout  = 8'b00000000; // 2673 :   0 - 0x0
      13'hA72: dout  = 8'b00000000; // 2674 :   0 - 0x0
      13'hA73: dout  = 8'b00000000; // 2675 :   0 - 0x0
      13'hA74: dout  = 8'b00000000; // 2676 :   0 - 0x0
      13'hA75: dout  = 8'b00000000; // 2677 :   0 - 0x0
      13'hA76: dout  = 8'b00000000; // 2678 :   0 - 0x0
      13'hA77: dout  = 8'b00000000; // 2679 :   0 - 0x0
      13'hA78: dout  = 8'b00000000; // 2680 :   0 - 0x0
      13'hA79: dout  = 8'b00000000; // 2681 :   0 - 0x0
      13'hA7A: dout  = 8'b00000000; // 2682 :   0 - 0x0
      13'hA7B: dout  = 8'b00000000; // 2683 :   0 - 0x0
      13'hA7C: dout  = 8'b00000000; // 2684 :   0 - 0x0
      13'hA7D: dout  = 8'b00000000; // 2685 :   0 - 0x0
      13'hA7E: dout  = 8'b00000000; // 2686 :   0 - 0x0
      13'hA7F: dout  = 8'b00000000; // 2687 :   0 - 0x0
      13'hA80: dout  = 8'b00000000; // 2688 :   0 - 0x0 -- Sprite 0xa8
      13'hA81: dout  = 8'b00000000; // 2689 :   0 - 0x0
      13'hA82: dout  = 8'b00000000; // 2690 :   0 - 0x0
      13'hA83: dout  = 8'b00000000; // 2691 :   0 - 0x0
      13'hA84: dout  = 8'b00000000; // 2692 :   0 - 0x0
      13'hA85: dout  = 8'b00000000; // 2693 :   0 - 0x0
      13'hA86: dout  = 8'b00000000; // 2694 :   0 - 0x0
      13'hA87: dout  = 8'b00000000; // 2695 :   0 - 0x0
      13'hA88: dout  = 8'b00000000; // 2696 :   0 - 0x0
      13'hA89: dout  = 8'b00000000; // 2697 :   0 - 0x0
      13'hA8A: dout  = 8'b00000000; // 2698 :   0 - 0x0
      13'hA8B: dout  = 8'b00000000; // 2699 :   0 - 0x0
      13'hA8C: dout  = 8'b00000000; // 2700 :   0 - 0x0
      13'hA8D: dout  = 8'b00000000; // 2701 :   0 - 0x0
      13'hA8E: dout  = 8'b00000000; // 2702 :   0 - 0x0
      13'hA8F: dout  = 8'b00000000; // 2703 :   0 - 0x0
      13'hA90: dout  = 8'b00000000; // 2704 :   0 - 0x0 -- Sprite 0xa9
      13'hA91: dout  = 8'b00000000; // 2705 :   0 - 0x0
      13'hA92: dout  = 8'b00000000; // 2706 :   0 - 0x0
      13'hA93: dout  = 8'b00000000; // 2707 :   0 - 0x0
      13'hA94: dout  = 8'b00000000; // 2708 :   0 - 0x0
      13'hA95: dout  = 8'b00000000; // 2709 :   0 - 0x0
      13'hA96: dout  = 8'b00000000; // 2710 :   0 - 0x0
      13'hA97: dout  = 8'b00000000; // 2711 :   0 - 0x0
      13'hA98: dout  = 8'b00000000; // 2712 :   0 - 0x0
      13'hA99: dout  = 8'b00000000; // 2713 :   0 - 0x0
      13'hA9A: dout  = 8'b00000000; // 2714 :   0 - 0x0
      13'hA9B: dout  = 8'b00000000; // 2715 :   0 - 0x0
      13'hA9C: dout  = 8'b00000000; // 2716 :   0 - 0x0
      13'hA9D: dout  = 8'b00000000; // 2717 :   0 - 0x0
      13'hA9E: dout  = 8'b00000000; // 2718 :   0 - 0x0
      13'hA9F: dout  = 8'b00000000; // 2719 :   0 - 0x0
      13'hAA0: dout  = 8'b00000000; // 2720 :   0 - 0x0 -- Sprite 0xaa
      13'hAA1: dout  = 8'b00000000; // 2721 :   0 - 0x0
      13'hAA2: dout  = 8'b00000000; // 2722 :   0 - 0x0
      13'hAA3: dout  = 8'b00000000; // 2723 :   0 - 0x0
      13'hAA4: dout  = 8'b00000000; // 2724 :   0 - 0x0
      13'hAA5: dout  = 8'b00000000; // 2725 :   0 - 0x0
      13'hAA6: dout  = 8'b00000000; // 2726 :   0 - 0x0
      13'hAA7: dout  = 8'b00000000; // 2727 :   0 - 0x0
      13'hAA8: dout  = 8'b00000000; // 2728 :   0 - 0x0
      13'hAA9: dout  = 8'b00000000; // 2729 :   0 - 0x0
      13'hAAA: dout  = 8'b00000000; // 2730 :   0 - 0x0
      13'hAAB: dout  = 8'b00000000; // 2731 :   0 - 0x0
      13'hAAC: dout  = 8'b00000000; // 2732 :   0 - 0x0
      13'hAAD: dout  = 8'b00000000; // 2733 :   0 - 0x0
      13'hAAE: dout  = 8'b00000000; // 2734 :   0 - 0x0
      13'hAAF: dout  = 8'b00000000; // 2735 :   0 - 0x0
      13'hAB0: dout  = 8'b00000000; // 2736 :   0 - 0x0 -- Sprite 0xab
      13'hAB1: dout  = 8'b00000000; // 2737 :   0 - 0x0
      13'hAB2: dout  = 8'b00000000; // 2738 :   0 - 0x0
      13'hAB3: dout  = 8'b00000000; // 2739 :   0 - 0x0
      13'hAB4: dout  = 8'b00000000; // 2740 :   0 - 0x0
      13'hAB5: dout  = 8'b00000000; // 2741 :   0 - 0x0
      13'hAB6: dout  = 8'b00000000; // 2742 :   0 - 0x0
      13'hAB7: dout  = 8'b00000000; // 2743 :   0 - 0x0
      13'hAB8: dout  = 8'b00000000; // 2744 :   0 - 0x0
      13'hAB9: dout  = 8'b00000000; // 2745 :   0 - 0x0
      13'hABA: dout  = 8'b00000000; // 2746 :   0 - 0x0
      13'hABB: dout  = 8'b00000000; // 2747 :   0 - 0x0
      13'hABC: dout  = 8'b00000000; // 2748 :   0 - 0x0
      13'hABD: dout  = 8'b00000000; // 2749 :   0 - 0x0
      13'hABE: dout  = 8'b00000000; // 2750 :   0 - 0x0
      13'hABF: dout  = 8'b00000000; // 2751 :   0 - 0x0
      13'hAC0: dout  = 8'b00000000; // 2752 :   0 - 0x0 -- Sprite 0xac
      13'hAC1: dout  = 8'b00000000; // 2753 :   0 - 0x0
      13'hAC2: dout  = 8'b00000000; // 2754 :   0 - 0x0
      13'hAC3: dout  = 8'b00000000; // 2755 :   0 - 0x0
      13'hAC4: dout  = 8'b00000000; // 2756 :   0 - 0x0
      13'hAC5: dout  = 8'b00000000; // 2757 :   0 - 0x0
      13'hAC6: dout  = 8'b00000000; // 2758 :   0 - 0x0
      13'hAC7: dout  = 8'b00000000; // 2759 :   0 - 0x0
      13'hAC8: dout  = 8'b00000000; // 2760 :   0 - 0x0
      13'hAC9: dout  = 8'b00000000; // 2761 :   0 - 0x0
      13'hACA: dout  = 8'b00000000; // 2762 :   0 - 0x0
      13'hACB: dout  = 8'b00000000; // 2763 :   0 - 0x0
      13'hACC: dout  = 8'b00000000; // 2764 :   0 - 0x0
      13'hACD: dout  = 8'b00000000; // 2765 :   0 - 0x0
      13'hACE: dout  = 8'b00000000; // 2766 :   0 - 0x0
      13'hACF: dout  = 8'b00000000; // 2767 :   0 - 0x0
      13'hAD0: dout  = 8'b00000000; // 2768 :   0 - 0x0 -- Sprite 0xad
      13'hAD1: dout  = 8'b00000000; // 2769 :   0 - 0x0
      13'hAD2: dout  = 8'b00000000; // 2770 :   0 - 0x0
      13'hAD3: dout  = 8'b00000000; // 2771 :   0 - 0x0
      13'hAD4: dout  = 8'b00000000; // 2772 :   0 - 0x0
      13'hAD5: dout  = 8'b00000000; // 2773 :   0 - 0x0
      13'hAD6: dout  = 8'b00000000; // 2774 :   0 - 0x0
      13'hAD7: dout  = 8'b00000000; // 2775 :   0 - 0x0
      13'hAD8: dout  = 8'b00000000; // 2776 :   0 - 0x0
      13'hAD9: dout  = 8'b00000000; // 2777 :   0 - 0x0
      13'hADA: dout  = 8'b00000000; // 2778 :   0 - 0x0
      13'hADB: dout  = 8'b00000000; // 2779 :   0 - 0x0
      13'hADC: dout  = 8'b00000000; // 2780 :   0 - 0x0
      13'hADD: dout  = 8'b00000000; // 2781 :   0 - 0x0
      13'hADE: dout  = 8'b00000000; // 2782 :   0 - 0x0
      13'hADF: dout  = 8'b00000000; // 2783 :   0 - 0x0
      13'hAE0: dout  = 8'b00000000; // 2784 :   0 - 0x0 -- Sprite 0xae
      13'hAE1: dout  = 8'b00000000; // 2785 :   0 - 0x0
      13'hAE2: dout  = 8'b00000000; // 2786 :   0 - 0x0
      13'hAE3: dout  = 8'b00000000; // 2787 :   0 - 0x0
      13'hAE4: dout  = 8'b00000000; // 2788 :   0 - 0x0
      13'hAE5: dout  = 8'b00000000; // 2789 :   0 - 0x0
      13'hAE6: dout  = 8'b00000000; // 2790 :   0 - 0x0
      13'hAE7: dout  = 8'b00000000; // 2791 :   0 - 0x0
      13'hAE8: dout  = 8'b00000000; // 2792 :   0 - 0x0
      13'hAE9: dout  = 8'b00000000; // 2793 :   0 - 0x0
      13'hAEA: dout  = 8'b00000000; // 2794 :   0 - 0x0
      13'hAEB: dout  = 8'b00000000; // 2795 :   0 - 0x0
      13'hAEC: dout  = 8'b00000000; // 2796 :   0 - 0x0
      13'hAED: dout  = 8'b00000000; // 2797 :   0 - 0x0
      13'hAEE: dout  = 8'b00000000; // 2798 :   0 - 0x0
      13'hAEF: dout  = 8'b00000000; // 2799 :   0 - 0x0
      13'hAF0: dout  = 8'b00000000; // 2800 :   0 - 0x0 -- Sprite 0xaf
      13'hAF1: dout  = 8'b00000000; // 2801 :   0 - 0x0
      13'hAF2: dout  = 8'b00000000; // 2802 :   0 - 0x0
      13'hAF3: dout  = 8'b00000000; // 2803 :   0 - 0x0
      13'hAF4: dout  = 8'b00000000; // 2804 :   0 - 0x0
      13'hAF5: dout  = 8'b00000000; // 2805 :   0 - 0x0
      13'hAF6: dout  = 8'b00000000; // 2806 :   0 - 0x0
      13'hAF7: dout  = 8'b00000000; // 2807 :   0 - 0x0
      13'hAF8: dout  = 8'b00000000; // 2808 :   0 - 0x0
      13'hAF9: dout  = 8'b00000000; // 2809 :   0 - 0x0
      13'hAFA: dout  = 8'b00000000; // 2810 :   0 - 0x0
      13'hAFB: dout  = 8'b00000000; // 2811 :   0 - 0x0
      13'hAFC: dout  = 8'b00000000; // 2812 :   0 - 0x0
      13'hAFD: dout  = 8'b00000000; // 2813 :   0 - 0x0
      13'hAFE: dout  = 8'b00000000; // 2814 :   0 - 0x0
      13'hAFF: dout  = 8'b00000000; // 2815 :   0 - 0x0
      13'hB00: dout  = 8'b00000000; // 2816 :   0 - 0x0 -- Sprite 0xb0
      13'hB01: dout  = 8'b00000000; // 2817 :   0 - 0x0
      13'hB02: dout  = 8'b00000000; // 2818 :   0 - 0x0
      13'hB03: dout  = 8'b00000000; // 2819 :   0 - 0x0
      13'hB04: dout  = 8'b00000000; // 2820 :   0 - 0x0
      13'hB05: dout  = 8'b00000000; // 2821 :   0 - 0x0
      13'hB06: dout  = 8'b00000000; // 2822 :   0 - 0x0
      13'hB07: dout  = 8'b00000000; // 2823 :   0 - 0x0
      13'hB08: dout  = 8'b00000000; // 2824 :   0 - 0x0
      13'hB09: dout  = 8'b00000000; // 2825 :   0 - 0x0
      13'hB0A: dout  = 8'b00000000; // 2826 :   0 - 0x0
      13'hB0B: dout  = 8'b00000000; // 2827 :   0 - 0x0
      13'hB0C: dout  = 8'b00000000; // 2828 :   0 - 0x0
      13'hB0D: dout  = 8'b00000000; // 2829 :   0 - 0x0
      13'hB0E: dout  = 8'b00000000; // 2830 :   0 - 0x0
      13'hB0F: dout  = 8'b00000000; // 2831 :   0 - 0x0
      13'hB10: dout  = 8'b00000000; // 2832 :   0 - 0x0 -- Sprite 0xb1
      13'hB11: dout  = 8'b00000000; // 2833 :   0 - 0x0
      13'hB12: dout  = 8'b00000000; // 2834 :   0 - 0x0
      13'hB13: dout  = 8'b00000000; // 2835 :   0 - 0x0
      13'hB14: dout  = 8'b00000000; // 2836 :   0 - 0x0
      13'hB15: dout  = 8'b00000000; // 2837 :   0 - 0x0
      13'hB16: dout  = 8'b00000000; // 2838 :   0 - 0x0
      13'hB17: dout  = 8'b00000000; // 2839 :   0 - 0x0
      13'hB18: dout  = 8'b00000000; // 2840 :   0 - 0x0
      13'hB19: dout  = 8'b00000000; // 2841 :   0 - 0x0
      13'hB1A: dout  = 8'b00000000; // 2842 :   0 - 0x0
      13'hB1B: dout  = 8'b00000000; // 2843 :   0 - 0x0
      13'hB1C: dout  = 8'b00000000; // 2844 :   0 - 0x0
      13'hB1D: dout  = 8'b00000000; // 2845 :   0 - 0x0
      13'hB1E: dout  = 8'b00000000; // 2846 :   0 - 0x0
      13'hB1F: dout  = 8'b00000000; // 2847 :   0 - 0x0
      13'hB20: dout  = 8'b00000000; // 2848 :   0 - 0x0 -- Sprite 0xb2
      13'hB21: dout  = 8'b00000000; // 2849 :   0 - 0x0
      13'hB22: dout  = 8'b00000000; // 2850 :   0 - 0x0
      13'hB23: dout  = 8'b00000000; // 2851 :   0 - 0x0
      13'hB24: dout  = 8'b00000000; // 2852 :   0 - 0x0
      13'hB25: dout  = 8'b00000000; // 2853 :   0 - 0x0
      13'hB26: dout  = 8'b00000000; // 2854 :   0 - 0x0
      13'hB27: dout  = 8'b00000000; // 2855 :   0 - 0x0
      13'hB28: dout  = 8'b00000000; // 2856 :   0 - 0x0
      13'hB29: dout  = 8'b00000000; // 2857 :   0 - 0x0
      13'hB2A: dout  = 8'b00000000; // 2858 :   0 - 0x0
      13'hB2B: dout  = 8'b00000000; // 2859 :   0 - 0x0
      13'hB2C: dout  = 8'b00000000; // 2860 :   0 - 0x0
      13'hB2D: dout  = 8'b00000000; // 2861 :   0 - 0x0
      13'hB2E: dout  = 8'b00000000; // 2862 :   0 - 0x0
      13'hB2F: dout  = 8'b00000000; // 2863 :   0 - 0x0
      13'hB30: dout  = 8'b00000000; // 2864 :   0 - 0x0 -- Sprite 0xb3
      13'hB31: dout  = 8'b00000000; // 2865 :   0 - 0x0
      13'hB32: dout  = 8'b00000000; // 2866 :   0 - 0x0
      13'hB33: dout  = 8'b00000000; // 2867 :   0 - 0x0
      13'hB34: dout  = 8'b00000000; // 2868 :   0 - 0x0
      13'hB35: dout  = 8'b00000000; // 2869 :   0 - 0x0
      13'hB36: dout  = 8'b00000000; // 2870 :   0 - 0x0
      13'hB37: dout  = 8'b00000000; // 2871 :   0 - 0x0
      13'hB38: dout  = 8'b00000000; // 2872 :   0 - 0x0
      13'hB39: dout  = 8'b00000000; // 2873 :   0 - 0x0
      13'hB3A: dout  = 8'b00000000; // 2874 :   0 - 0x0
      13'hB3B: dout  = 8'b00000000; // 2875 :   0 - 0x0
      13'hB3C: dout  = 8'b00000000; // 2876 :   0 - 0x0
      13'hB3D: dout  = 8'b00000000; // 2877 :   0 - 0x0
      13'hB3E: dout  = 8'b00000000; // 2878 :   0 - 0x0
      13'hB3F: dout  = 8'b00000000; // 2879 :   0 - 0x0
      13'hB40: dout  = 8'b00000000; // 2880 :   0 - 0x0 -- Sprite 0xb4
      13'hB41: dout  = 8'b00000000; // 2881 :   0 - 0x0
      13'hB42: dout  = 8'b00000000; // 2882 :   0 - 0x0
      13'hB43: dout  = 8'b00000000; // 2883 :   0 - 0x0
      13'hB44: dout  = 8'b00000000; // 2884 :   0 - 0x0
      13'hB45: dout  = 8'b00000000; // 2885 :   0 - 0x0
      13'hB46: dout  = 8'b00000000; // 2886 :   0 - 0x0
      13'hB47: dout  = 8'b00000000; // 2887 :   0 - 0x0
      13'hB48: dout  = 8'b00000000; // 2888 :   0 - 0x0
      13'hB49: dout  = 8'b00000000; // 2889 :   0 - 0x0
      13'hB4A: dout  = 8'b00000000; // 2890 :   0 - 0x0
      13'hB4B: dout  = 8'b00000000; // 2891 :   0 - 0x0
      13'hB4C: dout  = 8'b00000000; // 2892 :   0 - 0x0
      13'hB4D: dout  = 8'b00000000; // 2893 :   0 - 0x0
      13'hB4E: dout  = 8'b00000000; // 2894 :   0 - 0x0
      13'hB4F: dout  = 8'b00000000; // 2895 :   0 - 0x0
      13'hB50: dout  = 8'b00000000; // 2896 :   0 - 0x0 -- Sprite 0xb5
      13'hB51: dout  = 8'b00000000; // 2897 :   0 - 0x0
      13'hB52: dout  = 8'b00000000; // 2898 :   0 - 0x0
      13'hB53: dout  = 8'b00000000; // 2899 :   0 - 0x0
      13'hB54: dout  = 8'b00000000; // 2900 :   0 - 0x0
      13'hB55: dout  = 8'b00000000; // 2901 :   0 - 0x0
      13'hB56: dout  = 8'b00000000; // 2902 :   0 - 0x0
      13'hB57: dout  = 8'b00000000; // 2903 :   0 - 0x0
      13'hB58: dout  = 8'b00000000; // 2904 :   0 - 0x0
      13'hB59: dout  = 8'b00000000; // 2905 :   0 - 0x0
      13'hB5A: dout  = 8'b00000000; // 2906 :   0 - 0x0
      13'hB5B: dout  = 8'b00000000; // 2907 :   0 - 0x0
      13'hB5C: dout  = 8'b00000000; // 2908 :   0 - 0x0
      13'hB5D: dout  = 8'b00000000; // 2909 :   0 - 0x0
      13'hB5E: dout  = 8'b00000000; // 2910 :   0 - 0x0
      13'hB5F: dout  = 8'b00000000; // 2911 :   0 - 0x0
      13'hB60: dout  = 8'b00000000; // 2912 :   0 - 0x0 -- Sprite 0xb6
      13'hB61: dout  = 8'b00000000; // 2913 :   0 - 0x0
      13'hB62: dout  = 8'b00000000; // 2914 :   0 - 0x0
      13'hB63: dout  = 8'b00000000; // 2915 :   0 - 0x0
      13'hB64: dout  = 8'b00000000; // 2916 :   0 - 0x0
      13'hB65: dout  = 8'b00000000; // 2917 :   0 - 0x0
      13'hB66: dout  = 8'b00000000; // 2918 :   0 - 0x0
      13'hB67: dout  = 8'b00000000; // 2919 :   0 - 0x0
      13'hB68: dout  = 8'b00000000; // 2920 :   0 - 0x0
      13'hB69: dout  = 8'b00000000; // 2921 :   0 - 0x0
      13'hB6A: dout  = 8'b00000000; // 2922 :   0 - 0x0
      13'hB6B: dout  = 8'b00000000; // 2923 :   0 - 0x0
      13'hB6C: dout  = 8'b00000000; // 2924 :   0 - 0x0
      13'hB6D: dout  = 8'b00000000; // 2925 :   0 - 0x0
      13'hB6E: dout  = 8'b00000000; // 2926 :   0 - 0x0
      13'hB6F: dout  = 8'b00000000; // 2927 :   0 - 0x0
      13'hB70: dout  = 8'b00000000; // 2928 :   0 - 0x0 -- Sprite 0xb7
      13'hB71: dout  = 8'b00000000; // 2929 :   0 - 0x0
      13'hB72: dout  = 8'b00000000; // 2930 :   0 - 0x0
      13'hB73: dout  = 8'b00000000; // 2931 :   0 - 0x0
      13'hB74: dout  = 8'b00000000; // 2932 :   0 - 0x0
      13'hB75: dout  = 8'b00000000; // 2933 :   0 - 0x0
      13'hB76: dout  = 8'b00000000; // 2934 :   0 - 0x0
      13'hB77: dout  = 8'b00000000; // 2935 :   0 - 0x0
      13'hB78: dout  = 8'b00000000; // 2936 :   0 - 0x0
      13'hB79: dout  = 8'b00000000; // 2937 :   0 - 0x0
      13'hB7A: dout  = 8'b00000000; // 2938 :   0 - 0x0
      13'hB7B: dout  = 8'b00000000; // 2939 :   0 - 0x0
      13'hB7C: dout  = 8'b00000000; // 2940 :   0 - 0x0
      13'hB7D: dout  = 8'b00000000; // 2941 :   0 - 0x0
      13'hB7E: dout  = 8'b00000000; // 2942 :   0 - 0x0
      13'hB7F: dout  = 8'b00000000; // 2943 :   0 - 0x0
      13'hB80: dout  = 8'b00000000; // 2944 :   0 - 0x0 -- Sprite 0xb8
      13'hB81: dout  = 8'b00000000; // 2945 :   0 - 0x0
      13'hB82: dout  = 8'b00000000; // 2946 :   0 - 0x0
      13'hB83: dout  = 8'b00000000; // 2947 :   0 - 0x0
      13'hB84: dout  = 8'b00000000; // 2948 :   0 - 0x0
      13'hB85: dout  = 8'b00000000; // 2949 :   0 - 0x0
      13'hB86: dout  = 8'b00000000; // 2950 :   0 - 0x0
      13'hB87: dout  = 8'b00000000; // 2951 :   0 - 0x0
      13'hB88: dout  = 8'b00000000; // 2952 :   0 - 0x0
      13'hB89: dout  = 8'b00000000; // 2953 :   0 - 0x0
      13'hB8A: dout  = 8'b00000000; // 2954 :   0 - 0x0
      13'hB8B: dout  = 8'b00000000; // 2955 :   0 - 0x0
      13'hB8C: dout  = 8'b00000000; // 2956 :   0 - 0x0
      13'hB8D: dout  = 8'b00000000; // 2957 :   0 - 0x0
      13'hB8E: dout  = 8'b00000000; // 2958 :   0 - 0x0
      13'hB8F: dout  = 8'b00000000; // 2959 :   0 - 0x0
      13'hB90: dout  = 8'b00000000; // 2960 :   0 - 0x0 -- Sprite 0xb9
      13'hB91: dout  = 8'b00000000; // 2961 :   0 - 0x0
      13'hB92: dout  = 8'b00000000; // 2962 :   0 - 0x0
      13'hB93: dout  = 8'b00000000; // 2963 :   0 - 0x0
      13'hB94: dout  = 8'b00000000; // 2964 :   0 - 0x0
      13'hB95: dout  = 8'b00000000; // 2965 :   0 - 0x0
      13'hB96: dout  = 8'b00000000; // 2966 :   0 - 0x0
      13'hB97: dout  = 8'b00000000; // 2967 :   0 - 0x0
      13'hB98: dout  = 8'b00000000; // 2968 :   0 - 0x0
      13'hB99: dout  = 8'b00000000; // 2969 :   0 - 0x0
      13'hB9A: dout  = 8'b00000000; // 2970 :   0 - 0x0
      13'hB9B: dout  = 8'b00000000; // 2971 :   0 - 0x0
      13'hB9C: dout  = 8'b00000000; // 2972 :   0 - 0x0
      13'hB9D: dout  = 8'b00000000; // 2973 :   0 - 0x0
      13'hB9E: dout  = 8'b00000000; // 2974 :   0 - 0x0
      13'hB9F: dout  = 8'b00000000; // 2975 :   0 - 0x0
      13'hBA0: dout  = 8'b00000000; // 2976 :   0 - 0x0 -- Sprite 0xba
      13'hBA1: dout  = 8'b00000000; // 2977 :   0 - 0x0
      13'hBA2: dout  = 8'b00000000; // 2978 :   0 - 0x0
      13'hBA3: dout  = 8'b00000000; // 2979 :   0 - 0x0
      13'hBA4: dout  = 8'b00000000; // 2980 :   0 - 0x0
      13'hBA5: dout  = 8'b00000000; // 2981 :   0 - 0x0
      13'hBA6: dout  = 8'b00000000; // 2982 :   0 - 0x0
      13'hBA7: dout  = 8'b00000000; // 2983 :   0 - 0x0
      13'hBA8: dout  = 8'b00000000; // 2984 :   0 - 0x0
      13'hBA9: dout  = 8'b00000000; // 2985 :   0 - 0x0
      13'hBAA: dout  = 8'b00000000; // 2986 :   0 - 0x0
      13'hBAB: dout  = 8'b00000000; // 2987 :   0 - 0x0
      13'hBAC: dout  = 8'b00000000; // 2988 :   0 - 0x0
      13'hBAD: dout  = 8'b00000000; // 2989 :   0 - 0x0
      13'hBAE: dout  = 8'b00000000; // 2990 :   0 - 0x0
      13'hBAF: dout  = 8'b00000000; // 2991 :   0 - 0x0
      13'hBB0: dout  = 8'b00000000; // 2992 :   0 - 0x0 -- Sprite 0xbb
      13'hBB1: dout  = 8'b00000000; // 2993 :   0 - 0x0
      13'hBB2: dout  = 8'b00000000; // 2994 :   0 - 0x0
      13'hBB3: dout  = 8'b00000000; // 2995 :   0 - 0x0
      13'hBB4: dout  = 8'b00000000; // 2996 :   0 - 0x0
      13'hBB5: dout  = 8'b00000000; // 2997 :   0 - 0x0
      13'hBB6: dout  = 8'b00000000; // 2998 :   0 - 0x0
      13'hBB7: dout  = 8'b00000000; // 2999 :   0 - 0x0
      13'hBB8: dout  = 8'b00000000; // 3000 :   0 - 0x0
      13'hBB9: dout  = 8'b00000000; // 3001 :   0 - 0x0
      13'hBBA: dout  = 8'b00000000; // 3002 :   0 - 0x0
      13'hBBB: dout  = 8'b00000000; // 3003 :   0 - 0x0
      13'hBBC: dout  = 8'b00000000; // 3004 :   0 - 0x0
      13'hBBD: dout  = 8'b00000000; // 3005 :   0 - 0x0
      13'hBBE: dout  = 8'b00000000; // 3006 :   0 - 0x0
      13'hBBF: dout  = 8'b00000000; // 3007 :   0 - 0x0
      13'hBC0: dout  = 8'b00000000; // 3008 :   0 - 0x0 -- Sprite 0xbc
      13'hBC1: dout  = 8'b00000000; // 3009 :   0 - 0x0
      13'hBC2: dout  = 8'b00000000; // 3010 :   0 - 0x0
      13'hBC3: dout  = 8'b00000000; // 3011 :   0 - 0x0
      13'hBC4: dout  = 8'b00000000; // 3012 :   0 - 0x0
      13'hBC5: dout  = 8'b00000000; // 3013 :   0 - 0x0
      13'hBC6: dout  = 8'b00000000; // 3014 :   0 - 0x0
      13'hBC7: dout  = 8'b00000000; // 3015 :   0 - 0x0
      13'hBC8: dout  = 8'b00000000; // 3016 :   0 - 0x0
      13'hBC9: dout  = 8'b00000000; // 3017 :   0 - 0x0
      13'hBCA: dout  = 8'b00000000; // 3018 :   0 - 0x0
      13'hBCB: dout  = 8'b00000000; // 3019 :   0 - 0x0
      13'hBCC: dout  = 8'b00000000; // 3020 :   0 - 0x0
      13'hBCD: dout  = 8'b00000000; // 3021 :   0 - 0x0
      13'hBCE: dout  = 8'b00000000; // 3022 :   0 - 0x0
      13'hBCF: dout  = 8'b00000000; // 3023 :   0 - 0x0
      13'hBD0: dout  = 8'b00000000; // 3024 :   0 - 0x0 -- Sprite 0xbd
      13'hBD1: dout  = 8'b00000000; // 3025 :   0 - 0x0
      13'hBD2: dout  = 8'b00000000; // 3026 :   0 - 0x0
      13'hBD3: dout  = 8'b00000000; // 3027 :   0 - 0x0
      13'hBD4: dout  = 8'b00000000; // 3028 :   0 - 0x0
      13'hBD5: dout  = 8'b00000000; // 3029 :   0 - 0x0
      13'hBD6: dout  = 8'b00000000; // 3030 :   0 - 0x0
      13'hBD7: dout  = 8'b00000000; // 3031 :   0 - 0x0
      13'hBD8: dout  = 8'b00000000; // 3032 :   0 - 0x0
      13'hBD9: dout  = 8'b00000000; // 3033 :   0 - 0x0
      13'hBDA: dout  = 8'b00000000; // 3034 :   0 - 0x0
      13'hBDB: dout  = 8'b00000000; // 3035 :   0 - 0x0
      13'hBDC: dout  = 8'b00000000; // 3036 :   0 - 0x0
      13'hBDD: dout  = 8'b00000000; // 3037 :   0 - 0x0
      13'hBDE: dout  = 8'b00000000; // 3038 :   0 - 0x0
      13'hBDF: dout  = 8'b00000000; // 3039 :   0 - 0x0
      13'hBE0: dout  = 8'b00000000; // 3040 :   0 - 0x0 -- Sprite 0xbe
      13'hBE1: dout  = 8'b00000000; // 3041 :   0 - 0x0
      13'hBE2: dout  = 8'b00000000; // 3042 :   0 - 0x0
      13'hBE3: dout  = 8'b00000000; // 3043 :   0 - 0x0
      13'hBE4: dout  = 8'b00000000; // 3044 :   0 - 0x0
      13'hBE5: dout  = 8'b00000000; // 3045 :   0 - 0x0
      13'hBE6: dout  = 8'b00000000; // 3046 :   0 - 0x0
      13'hBE7: dout  = 8'b00000000; // 3047 :   0 - 0x0
      13'hBE8: dout  = 8'b00000000; // 3048 :   0 - 0x0
      13'hBE9: dout  = 8'b00000000; // 3049 :   0 - 0x0
      13'hBEA: dout  = 8'b00000000; // 3050 :   0 - 0x0
      13'hBEB: dout  = 8'b00000000; // 3051 :   0 - 0x0
      13'hBEC: dout  = 8'b00000000; // 3052 :   0 - 0x0
      13'hBED: dout  = 8'b00000000; // 3053 :   0 - 0x0
      13'hBEE: dout  = 8'b00000000; // 3054 :   0 - 0x0
      13'hBEF: dout  = 8'b00000000; // 3055 :   0 - 0x0
      13'hBF0: dout  = 8'b00000000; // 3056 :   0 - 0x0 -- Sprite 0xbf
      13'hBF1: dout  = 8'b00000000; // 3057 :   0 - 0x0
      13'hBF2: dout  = 8'b00000000; // 3058 :   0 - 0x0
      13'hBF3: dout  = 8'b00000000; // 3059 :   0 - 0x0
      13'hBF4: dout  = 8'b00000000; // 3060 :   0 - 0x0
      13'hBF5: dout  = 8'b00000000; // 3061 :   0 - 0x0
      13'hBF6: dout  = 8'b00000000; // 3062 :   0 - 0x0
      13'hBF7: dout  = 8'b00000000; // 3063 :   0 - 0x0
      13'hBF8: dout  = 8'b00000000; // 3064 :   0 - 0x0
      13'hBF9: dout  = 8'b00000000; // 3065 :   0 - 0x0
      13'hBFA: dout  = 8'b00000000; // 3066 :   0 - 0x0
      13'hBFB: dout  = 8'b00000000; // 3067 :   0 - 0x0
      13'hBFC: dout  = 8'b00000000; // 3068 :   0 - 0x0
      13'hBFD: dout  = 8'b00000000; // 3069 :   0 - 0x0
      13'hBFE: dout  = 8'b00000000; // 3070 :   0 - 0x0
      13'hBFF: dout  = 8'b00000000; // 3071 :   0 - 0x0
      13'hC00: dout  = 8'b00000000; // 3072 :   0 - 0x0 -- Sprite 0xc0
      13'hC01: dout  = 8'b00000000; // 3073 :   0 - 0x0
      13'hC02: dout  = 8'b00000000; // 3074 :   0 - 0x0
      13'hC03: dout  = 8'b00000000; // 3075 :   0 - 0x0
      13'hC04: dout  = 8'b00000000; // 3076 :   0 - 0x0
      13'hC05: dout  = 8'b00000000; // 3077 :   0 - 0x0
      13'hC06: dout  = 8'b00000000; // 3078 :   0 - 0x0
      13'hC07: dout  = 8'b00000000; // 3079 :   0 - 0x0
      13'hC08: dout  = 8'b00000000; // 3080 :   0 - 0x0
      13'hC09: dout  = 8'b00000000; // 3081 :   0 - 0x0
      13'hC0A: dout  = 8'b00000000; // 3082 :   0 - 0x0
      13'hC0B: dout  = 8'b00000000; // 3083 :   0 - 0x0
      13'hC0C: dout  = 8'b00000000; // 3084 :   0 - 0x0
      13'hC0D: dout  = 8'b00000000; // 3085 :   0 - 0x0
      13'hC0E: dout  = 8'b00000000; // 3086 :   0 - 0x0
      13'hC0F: dout  = 8'b00000000; // 3087 :   0 - 0x0
      13'hC10: dout  = 8'b00000000; // 3088 :   0 - 0x0 -- Sprite 0xc1
      13'hC11: dout  = 8'b00000000; // 3089 :   0 - 0x0
      13'hC12: dout  = 8'b00000000; // 3090 :   0 - 0x0
      13'hC13: dout  = 8'b00000000; // 3091 :   0 - 0x0
      13'hC14: dout  = 8'b00000000; // 3092 :   0 - 0x0
      13'hC15: dout  = 8'b00000000; // 3093 :   0 - 0x0
      13'hC16: dout  = 8'b00000000; // 3094 :   0 - 0x0
      13'hC17: dout  = 8'b00000000; // 3095 :   0 - 0x0
      13'hC18: dout  = 8'b00000000; // 3096 :   0 - 0x0
      13'hC19: dout  = 8'b00000000; // 3097 :   0 - 0x0
      13'hC1A: dout  = 8'b00000000; // 3098 :   0 - 0x0
      13'hC1B: dout  = 8'b00000000; // 3099 :   0 - 0x0
      13'hC1C: dout  = 8'b00000000; // 3100 :   0 - 0x0
      13'hC1D: dout  = 8'b00000000; // 3101 :   0 - 0x0
      13'hC1E: dout  = 8'b00000000; // 3102 :   0 - 0x0
      13'hC1F: dout  = 8'b00000000; // 3103 :   0 - 0x0
      13'hC20: dout  = 8'b00000000; // 3104 :   0 - 0x0 -- Sprite 0xc2
      13'hC21: dout  = 8'b00000000; // 3105 :   0 - 0x0
      13'hC22: dout  = 8'b00000000; // 3106 :   0 - 0x0
      13'hC23: dout  = 8'b00000000; // 3107 :   0 - 0x0
      13'hC24: dout  = 8'b00000000; // 3108 :   0 - 0x0
      13'hC25: dout  = 8'b00000000; // 3109 :   0 - 0x0
      13'hC26: dout  = 8'b00000000; // 3110 :   0 - 0x0
      13'hC27: dout  = 8'b00000000; // 3111 :   0 - 0x0
      13'hC28: dout  = 8'b00000000; // 3112 :   0 - 0x0
      13'hC29: dout  = 8'b00000000; // 3113 :   0 - 0x0
      13'hC2A: dout  = 8'b00000000; // 3114 :   0 - 0x0
      13'hC2B: dout  = 8'b00000000; // 3115 :   0 - 0x0
      13'hC2C: dout  = 8'b00000000; // 3116 :   0 - 0x0
      13'hC2D: dout  = 8'b00000000; // 3117 :   0 - 0x0
      13'hC2E: dout  = 8'b00000000; // 3118 :   0 - 0x0
      13'hC2F: dout  = 8'b00000000; // 3119 :   0 - 0x0
      13'hC30: dout  = 8'b00000000; // 3120 :   0 - 0x0 -- Sprite 0xc3
      13'hC31: dout  = 8'b00000000; // 3121 :   0 - 0x0
      13'hC32: dout  = 8'b00000000; // 3122 :   0 - 0x0
      13'hC33: dout  = 8'b00000000; // 3123 :   0 - 0x0
      13'hC34: dout  = 8'b00000000; // 3124 :   0 - 0x0
      13'hC35: dout  = 8'b00000000; // 3125 :   0 - 0x0
      13'hC36: dout  = 8'b00000000; // 3126 :   0 - 0x0
      13'hC37: dout  = 8'b00000000; // 3127 :   0 - 0x0
      13'hC38: dout  = 8'b00000000; // 3128 :   0 - 0x0
      13'hC39: dout  = 8'b00000000; // 3129 :   0 - 0x0
      13'hC3A: dout  = 8'b00000000; // 3130 :   0 - 0x0
      13'hC3B: dout  = 8'b00000000; // 3131 :   0 - 0x0
      13'hC3C: dout  = 8'b00000000; // 3132 :   0 - 0x0
      13'hC3D: dout  = 8'b00000000; // 3133 :   0 - 0x0
      13'hC3E: dout  = 8'b00000000; // 3134 :   0 - 0x0
      13'hC3F: dout  = 8'b00000000; // 3135 :   0 - 0x0
      13'hC40: dout  = 8'b00000000; // 3136 :   0 - 0x0 -- Sprite 0xc4
      13'hC41: dout  = 8'b00000000; // 3137 :   0 - 0x0
      13'hC42: dout  = 8'b00000000; // 3138 :   0 - 0x0
      13'hC43: dout  = 8'b00000000; // 3139 :   0 - 0x0
      13'hC44: dout  = 8'b00000000; // 3140 :   0 - 0x0
      13'hC45: dout  = 8'b00000000; // 3141 :   0 - 0x0
      13'hC46: dout  = 8'b00000000; // 3142 :   0 - 0x0
      13'hC47: dout  = 8'b00000000; // 3143 :   0 - 0x0
      13'hC48: dout  = 8'b00000000; // 3144 :   0 - 0x0
      13'hC49: dout  = 8'b00000000; // 3145 :   0 - 0x0
      13'hC4A: dout  = 8'b00000000; // 3146 :   0 - 0x0
      13'hC4B: dout  = 8'b00000000; // 3147 :   0 - 0x0
      13'hC4C: dout  = 8'b00000000; // 3148 :   0 - 0x0
      13'hC4D: dout  = 8'b00000000; // 3149 :   0 - 0x0
      13'hC4E: dout  = 8'b00000000; // 3150 :   0 - 0x0
      13'hC4F: dout  = 8'b00000000; // 3151 :   0 - 0x0
      13'hC50: dout  = 8'b00000000; // 3152 :   0 - 0x0 -- Sprite 0xc5
      13'hC51: dout  = 8'b00000000; // 3153 :   0 - 0x0
      13'hC52: dout  = 8'b00000000; // 3154 :   0 - 0x0
      13'hC53: dout  = 8'b00000000; // 3155 :   0 - 0x0
      13'hC54: dout  = 8'b00000000; // 3156 :   0 - 0x0
      13'hC55: dout  = 8'b00000000; // 3157 :   0 - 0x0
      13'hC56: dout  = 8'b00000000; // 3158 :   0 - 0x0
      13'hC57: dout  = 8'b00000000; // 3159 :   0 - 0x0
      13'hC58: dout  = 8'b00000000; // 3160 :   0 - 0x0
      13'hC59: dout  = 8'b00000000; // 3161 :   0 - 0x0
      13'hC5A: dout  = 8'b00000000; // 3162 :   0 - 0x0
      13'hC5B: dout  = 8'b00000000; // 3163 :   0 - 0x0
      13'hC5C: dout  = 8'b00000000; // 3164 :   0 - 0x0
      13'hC5D: dout  = 8'b00000000; // 3165 :   0 - 0x0
      13'hC5E: dout  = 8'b00000000; // 3166 :   0 - 0x0
      13'hC5F: dout  = 8'b00000000; // 3167 :   0 - 0x0
      13'hC60: dout  = 8'b00000000; // 3168 :   0 - 0x0 -- Sprite 0xc6
      13'hC61: dout  = 8'b00000000; // 3169 :   0 - 0x0
      13'hC62: dout  = 8'b00000000; // 3170 :   0 - 0x0
      13'hC63: dout  = 8'b00000000; // 3171 :   0 - 0x0
      13'hC64: dout  = 8'b00000000; // 3172 :   0 - 0x0
      13'hC65: dout  = 8'b00000000; // 3173 :   0 - 0x0
      13'hC66: dout  = 8'b00000000; // 3174 :   0 - 0x0
      13'hC67: dout  = 8'b00000000; // 3175 :   0 - 0x0
      13'hC68: dout  = 8'b00000000; // 3176 :   0 - 0x0
      13'hC69: dout  = 8'b00000000; // 3177 :   0 - 0x0
      13'hC6A: dout  = 8'b00000000; // 3178 :   0 - 0x0
      13'hC6B: dout  = 8'b00000000; // 3179 :   0 - 0x0
      13'hC6C: dout  = 8'b00000000; // 3180 :   0 - 0x0
      13'hC6D: dout  = 8'b00000000; // 3181 :   0 - 0x0
      13'hC6E: dout  = 8'b00000000; // 3182 :   0 - 0x0
      13'hC6F: dout  = 8'b00000000; // 3183 :   0 - 0x0
      13'hC70: dout  = 8'b00000000; // 3184 :   0 - 0x0 -- Sprite 0xc7
      13'hC71: dout  = 8'b00000000; // 3185 :   0 - 0x0
      13'hC72: dout  = 8'b00000000; // 3186 :   0 - 0x0
      13'hC73: dout  = 8'b00000000; // 3187 :   0 - 0x0
      13'hC74: dout  = 8'b00000000; // 3188 :   0 - 0x0
      13'hC75: dout  = 8'b00000000; // 3189 :   0 - 0x0
      13'hC76: dout  = 8'b00000000; // 3190 :   0 - 0x0
      13'hC77: dout  = 8'b00000000; // 3191 :   0 - 0x0
      13'hC78: dout  = 8'b00000000; // 3192 :   0 - 0x0
      13'hC79: dout  = 8'b00000000; // 3193 :   0 - 0x0
      13'hC7A: dout  = 8'b00000000; // 3194 :   0 - 0x0
      13'hC7B: dout  = 8'b00000000; // 3195 :   0 - 0x0
      13'hC7C: dout  = 8'b00000000; // 3196 :   0 - 0x0
      13'hC7D: dout  = 8'b00000000; // 3197 :   0 - 0x0
      13'hC7E: dout  = 8'b00000000; // 3198 :   0 - 0x0
      13'hC7F: dout  = 8'b00000000; // 3199 :   0 - 0x0
      13'hC80: dout  = 8'b00000000; // 3200 :   0 - 0x0 -- Sprite 0xc8
      13'hC81: dout  = 8'b00000000; // 3201 :   0 - 0x0
      13'hC82: dout  = 8'b00000000; // 3202 :   0 - 0x0
      13'hC83: dout  = 8'b00000000; // 3203 :   0 - 0x0
      13'hC84: dout  = 8'b00000000; // 3204 :   0 - 0x0
      13'hC85: dout  = 8'b00000000; // 3205 :   0 - 0x0
      13'hC86: dout  = 8'b00000000; // 3206 :   0 - 0x0
      13'hC87: dout  = 8'b00000000; // 3207 :   0 - 0x0
      13'hC88: dout  = 8'b00000000; // 3208 :   0 - 0x0
      13'hC89: dout  = 8'b00000000; // 3209 :   0 - 0x0
      13'hC8A: dout  = 8'b00000000; // 3210 :   0 - 0x0
      13'hC8B: dout  = 8'b00000000; // 3211 :   0 - 0x0
      13'hC8C: dout  = 8'b00000000; // 3212 :   0 - 0x0
      13'hC8D: dout  = 8'b00000000; // 3213 :   0 - 0x0
      13'hC8E: dout  = 8'b00000000; // 3214 :   0 - 0x0
      13'hC8F: dout  = 8'b00000000; // 3215 :   0 - 0x0
      13'hC90: dout  = 8'b00000000; // 3216 :   0 - 0x0 -- Sprite 0xc9
      13'hC91: dout  = 8'b00000000; // 3217 :   0 - 0x0
      13'hC92: dout  = 8'b00000000; // 3218 :   0 - 0x0
      13'hC93: dout  = 8'b00000000; // 3219 :   0 - 0x0
      13'hC94: dout  = 8'b00000000; // 3220 :   0 - 0x0
      13'hC95: dout  = 8'b00000000; // 3221 :   0 - 0x0
      13'hC96: dout  = 8'b00000000; // 3222 :   0 - 0x0
      13'hC97: dout  = 8'b00000000; // 3223 :   0 - 0x0
      13'hC98: dout  = 8'b00000000; // 3224 :   0 - 0x0
      13'hC99: dout  = 8'b00000000; // 3225 :   0 - 0x0
      13'hC9A: dout  = 8'b00000000; // 3226 :   0 - 0x0
      13'hC9B: dout  = 8'b00000000; // 3227 :   0 - 0x0
      13'hC9C: dout  = 8'b00000000; // 3228 :   0 - 0x0
      13'hC9D: dout  = 8'b00000000; // 3229 :   0 - 0x0
      13'hC9E: dout  = 8'b00000000; // 3230 :   0 - 0x0
      13'hC9F: dout  = 8'b00000000; // 3231 :   0 - 0x0
      13'hCA0: dout  = 8'b00000000; // 3232 :   0 - 0x0 -- Sprite 0xca
      13'hCA1: dout  = 8'b00000000; // 3233 :   0 - 0x0
      13'hCA2: dout  = 8'b00000000; // 3234 :   0 - 0x0
      13'hCA3: dout  = 8'b00000000; // 3235 :   0 - 0x0
      13'hCA4: dout  = 8'b00000000; // 3236 :   0 - 0x0
      13'hCA5: dout  = 8'b00000000; // 3237 :   0 - 0x0
      13'hCA6: dout  = 8'b00000000; // 3238 :   0 - 0x0
      13'hCA7: dout  = 8'b00000000; // 3239 :   0 - 0x0
      13'hCA8: dout  = 8'b00000000; // 3240 :   0 - 0x0
      13'hCA9: dout  = 8'b00000000; // 3241 :   0 - 0x0
      13'hCAA: dout  = 8'b00000000; // 3242 :   0 - 0x0
      13'hCAB: dout  = 8'b00000000; // 3243 :   0 - 0x0
      13'hCAC: dout  = 8'b00000000; // 3244 :   0 - 0x0
      13'hCAD: dout  = 8'b00000000; // 3245 :   0 - 0x0
      13'hCAE: dout  = 8'b00000000; // 3246 :   0 - 0x0
      13'hCAF: dout  = 8'b00000000; // 3247 :   0 - 0x0
      13'hCB0: dout  = 8'b00000000; // 3248 :   0 - 0x0 -- Sprite 0xcb
      13'hCB1: dout  = 8'b00000000; // 3249 :   0 - 0x0
      13'hCB2: dout  = 8'b00000000; // 3250 :   0 - 0x0
      13'hCB3: dout  = 8'b00000000; // 3251 :   0 - 0x0
      13'hCB4: dout  = 8'b00000000; // 3252 :   0 - 0x0
      13'hCB5: dout  = 8'b00000000; // 3253 :   0 - 0x0
      13'hCB6: dout  = 8'b00000000; // 3254 :   0 - 0x0
      13'hCB7: dout  = 8'b00000000; // 3255 :   0 - 0x0
      13'hCB8: dout  = 8'b00000000; // 3256 :   0 - 0x0
      13'hCB9: dout  = 8'b00000000; // 3257 :   0 - 0x0
      13'hCBA: dout  = 8'b00000000; // 3258 :   0 - 0x0
      13'hCBB: dout  = 8'b00000000; // 3259 :   0 - 0x0
      13'hCBC: dout  = 8'b00000000; // 3260 :   0 - 0x0
      13'hCBD: dout  = 8'b00000000; // 3261 :   0 - 0x0
      13'hCBE: dout  = 8'b00000000; // 3262 :   0 - 0x0
      13'hCBF: dout  = 8'b00000000; // 3263 :   0 - 0x0
      13'hCC0: dout  = 8'b00000000; // 3264 :   0 - 0x0 -- Sprite 0xcc
      13'hCC1: dout  = 8'b00000000; // 3265 :   0 - 0x0
      13'hCC2: dout  = 8'b00000000; // 3266 :   0 - 0x0
      13'hCC3: dout  = 8'b00000000; // 3267 :   0 - 0x0
      13'hCC4: dout  = 8'b00000000; // 3268 :   0 - 0x0
      13'hCC5: dout  = 8'b00000000; // 3269 :   0 - 0x0
      13'hCC6: dout  = 8'b00000000; // 3270 :   0 - 0x0
      13'hCC7: dout  = 8'b00000000; // 3271 :   0 - 0x0
      13'hCC8: dout  = 8'b00000000; // 3272 :   0 - 0x0
      13'hCC9: dout  = 8'b00000000; // 3273 :   0 - 0x0
      13'hCCA: dout  = 8'b00000000; // 3274 :   0 - 0x0
      13'hCCB: dout  = 8'b00000000; // 3275 :   0 - 0x0
      13'hCCC: dout  = 8'b00000000; // 3276 :   0 - 0x0
      13'hCCD: dout  = 8'b00000000; // 3277 :   0 - 0x0
      13'hCCE: dout  = 8'b00000000; // 3278 :   0 - 0x0
      13'hCCF: dout  = 8'b00000000; // 3279 :   0 - 0x0
      13'hCD0: dout  = 8'b00000000; // 3280 :   0 - 0x0 -- Sprite 0xcd
      13'hCD1: dout  = 8'b00000000; // 3281 :   0 - 0x0
      13'hCD2: dout  = 8'b00000000; // 3282 :   0 - 0x0
      13'hCD3: dout  = 8'b00000000; // 3283 :   0 - 0x0
      13'hCD4: dout  = 8'b00000000; // 3284 :   0 - 0x0
      13'hCD5: dout  = 8'b00000000; // 3285 :   0 - 0x0
      13'hCD6: dout  = 8'b00000000; // 3286 :   0 - 0x0
      13'hCD7: dout  = 8'b00000000; // 3287 :   0 - 0x0
      13'hCD8: dout  = 8'b00000000; // 3288 :   0 - 0x0
      13'hCD9: dout  = 8'b00000000; // 3289 :   0 - 0x0
      13'hCDA: dout  = 8'b00000000; // 3290 :   0 - 0x0
      13'hCDB: dout  = 8'b00000000; // 3291 :   0 - 0x0
      13'hCDC: dout  = 8'b00000000; // 3292 :   0 - 0x0
      13'hCDD: dout  = 8'b00000000; // 3293 :   0 - 0x0
      13'hCDE: dout  = 8'b00000000; // 3294 :   0 - 0x0
      13'hCDF: dout  = 8'b00000000; // 3295 :   0 - 0x0
      13'hCE0: dout  = 8'b00000000; // 3296 :   0 - 0x0 -- Sprite 0xce
      13'hCE1: dout  = 8'b00000000; // 3297 :   0 - 0x0
      13'hCE2: dout  = 8'b00000000; // 3298 :   0 - 0x0
      13'hCE3: dout  = 8'b00000000; // 3299 :   0 - 0x0
      13'hCE4: dout  = 8'b00000000; // 3300 :   0 - 0x0
      13'hCE5: dout  = 8'b00000000; // 3301 :   0 - 0x0
      13'hCE6: dout  = 8'b00000000; // 3302 :   0 - 0x0
      13'hCE7: dout  = 8'b00000000; // 3303 :   0 - 0x0
      13'hCE8: dout  = 8'b00000000; // 3304 :   0 - 0x0
      13'hCE9: dout  = 8'b00000000; // 3305 :   0 - 0x0
      13'hCEA: dout  = 8'b00000000; // 3306 :   0 - 0x0
      13'hCEB: dout  = 8'b00000000; // 3307 :   0 - 0x0
      13'hCEC: dout  = 8'b00000000; // 3308 :   0 - 0x0
      13'hCED: dout  = 8'b00000000; // 3309 :   0 - 0x0
      13'hCEE: dout  = 8'b00000000; // 3310 :   0 - 0x0
      13'hCEF: dout  = 8'b00000000; // 3311 :   0 - 0x0
      13'hCF0: dout  = 8'b00000000; // 3312 :   0 - 0x0 -- Sprite 0xcf
      13'hCF1: dout  = 8'b00000000; // 3313 :   0 - 0x0
      13'hCF2: dout  = 8'b00000000; // 3314 :   0 - 0x0
      13'hCF3: dout  = 8'b00000000; // 3315 :   0 - 0x0
      13'hCF4: dout  = 8'b00000000; // 3316 :   0 - 0x0
      13'hCF5: dout  = 8'b00000000; // 3317 :   0 - 0x0
      13'hCF6: dout  = 8'b00000000; // 3318 :   0 - 0x0
      13'hCF7: dout  = 8'b00000000; // 3319 :   0 - 0x0
      13'hCF8: dout  = 8'b00000000; // 3320 :   0 - 0x0
      13'hCF9: dout  = 8'b00000000; // 3321 :   0 - 0x0
      13'hCFA: dout  = 8'b00000000; // 3322 :   0 - 0x0
      13'hCFB: dout  = 8'b00000000; // 3323 :   0 - 0x0
      13'hCFC: dout  = 8'b00000000; // 3324 :   0 - 0x0
      13'hCFD: dout  = 8'b00000000; // 3325 :   0 - 0x0
      13'hCFE: dout  = 8'b00000000; // 3326 :   0 - 0x0
      13'hCFF: dout  = 8'b00000000; // 3327 :   0 - 0x0
      13'hD00: dout  = 8'b00000000; // 3328 :   0 - 0x0 -- Sprite 0xd0
      13'hD01: dout  = 8'b00000000; // 3329 :   0 - 0x0
      13'hD02: dout  = 8'b00000000; // 3330 :   0 - 0x0
      13'hD03: dout  = 8'b00000000; // 3331 :   0 - 0x0
      13'hD04: dout  = 8'b00000000; // 3332 :   0 - 0x0
      13'hD05: dout  = 8'b00000000; // 3333 :   0 - 0x0
      13'hD06: dout  = 8'b00000000; // 3334 :   0 - 0x0
      13'hD07: dout  = 8'b00000000; // 3335 :   0 - 0x0
      13'hD08: dout  = 8'b00000000; // 3336 :   0 - 0x0
      13'hD09: dout  = 8'b00000000; // 3337 :   0 - 0x0
      13'hD0A: dout  = 8'b00000000; // 3338 :   0 - 0x0
      13'hD0B: dout  = 8'b00000000; // 3339 :   0 - 0x0
      13'hD0C: dout  = 8'b00000000; // 3340 :   0 - 0x0
      13'hD0D: dout  = 8'b00000000; // 3341 :   0 - 0x0
      13'hD0E: dout  = 8'b00000000; // 3342 :   0 - 0x0
      13'hD0F: dout  = 8'b00000000; // 3343 :   0 - 0x0
      13'hD10: dout  = 8'b00000000; // 3344 :   0 - 0x0 -- Sprite 0xd1
      13'hD11: dout  = 8'b00000000; // 3345 :   0 - 0x0
      13'hD12: dout  = 8'b00000000; // 3346 :   0 - 0x0
      13'hD13: dout  = 8'b00000000; // 3347 :   0 - 0x0
      13'hD14: dout  = 8'b00000000; // 3348 :   0 - 0x0
      13'hD15: dout  = 8'b00000000; // 3349 :   0 - 0x0
      13'hD16: dout  = 8'b00000000; // 3350 :   0 - 0x0
      13'hD17: dout  = 8'b00000000; // 3351 :   0 - 0x0
      13'hD18: dout  = 8'b00000000; // 3352 :   0 - 0x0
      13'hD19: dout  = 8'b00000000; // 3353 :   0 - 0x0
      13'hD1A: dout  = 8'b00000000; // 3354 :   0 - 0x0
      13'hD1B: dout  = 8'b00000000; // 3355 :   0 - 0x0
      13'hD1C: dout  = 8'b00000000; // 3356 :   0 - 0x0
      13'hD1D: dout  = 8'b00000000; // 3357 :   0 - 0x0
      13'hD1E: dout  = 8'b00000000; // 3358 :   0 - 0x0
      13'hD1F: dout  = 8'b00000000; // 3359 :   0 - 0x0
      13'hD20: dout  = 8'b00000000; // 3360 :   0 - 0x0 -- Sprite 0xd2
      13'hD21: dout  = 8'b00000000; // 3361 :   0 - 0x0
      13'hD22: dout  = 8'b00000000; // 3362 :   0 - 0x0
      13'hD23: dout  = 8'b00000000; // 3363 :   0 - 0x0
      13'hD24: dout  = 8'b00000000; // 3364 :   0 - 0x0
      13'hD25: dout  = 8'b00000000; // 3365 :   0 - 0x0
      13'hD26: dout  = 8'b00000000; // 3366 :   0 - 0x0
      13'hD27: dout  = 8'b00000000; // 3367 :   0 - 0x0
      13'hD28: dout  = 8'b00000000; // 3368 :   0 - 0x0
      13'hD29: dout  = 8'b00000000; // 3369 :   0 - 0x0
      13'hD2A: dout  = 8'b00000000; // 3370 :   0 - 0x0
      13'hD2B: dout  = 8'b00000000; // 3371 :   0 - 0x0
      13'hD2C: dout  = 8'b00000000; // 3372 :   0 - 0x0
      13'hD2D: dout  = 8'b00000000; // 3373 :   0 - 0x0
      13'hD2E: dout  = 8'b00000000; // 3374 :   0 - 0x0
      13'hD2F: dout  = 8'b00000000; // 3375 :   0 - 0x0
      13'hD30: dout  = 8'b00000000; // 3376 :   0 - 0x0 -- Sprite 0xd3
      13'hD31: dout  = 8'b00000000; // 3377 :   0 - 0x0
      13'hD32: dout  = 8'b00000000; // 3378 :   0 - 0x0
      13'hD33: dout  = 8'b00000000; // 3379 :   0 - 0x0
      13'hD34: dout  = 8'b00000000; // 3380 :   0 - 0x0
      13'hD35: dout  = 8'b00000000; // 3381 :   0 - 0x0
      13'hD36: dout  = 8'b00000000; // 3382 :   0 - 0x0
      13'hD37: dout  = 8'b00000000; // 3383 :   0 - 0x0
      13'hD38: dout  = 8'b00000000; // 3384 :   0 - 0x0
      13'hD39: dout  = 8'b00000000; // 3385 :   0 - 0x0
      13'hD3A: dout  = 8'b00000000; // 3386 :   0 - 0x0
      13'hD3B: dout  = 8'b00000000; // 3387 :   0 - 0x0
      13'hD3C: dout  = 8'b00000000; // 3388 :   0 - 0x0
      13'hD3D: dout  = 8'b00000000; // 3389 :   0 - 0x0
      13'hD3E: dout  = 8'b00000000; // 3390 :   0 - 0x0
      13'hD3F: dout  = 8'b00000000; // 3391 :   0 - 0x0
      13'hD40: dout  = 8'b00000000; // 3392 :   0 - 0x0 -- Sprite 0xd4
      13'hD41: dout  = 8'b00000000; // 3393 :   0 - 0x0
      13'hD42: dout  = 8'b00000000; // 3394 :   0 - 0x0
      13'hD43: dout  = 8'b00000000; // 3395 :   0 - 0x0
      13'hD44: dout  = 8'b00000000; // 3396 :   0 - 0x0
      13'hD45: dout  = 8'b00000000; // 3397 :   0 - 0x0
      13'hD46: dout  = 8'b00000000; // 3398 :   0 - 0x0
      13'hD47: dout  = 8'b00000000; // 3399 :   0 - 0x0
      13'hD48: dout  = 8'b00000000; // 3400 :   0 - 0x0
      13'hD49: dout  = 8'b00000000; // 3401 :   0 - 0x0
      13'hD4A: dout  = 8'b00000000; // 3402 :   0 - 0x0
      13'hD4B: dout  = 8'b00000000; // 3403 :   0 - 0x0
      13'hD4C: dout  = 8'b00000000; // 3404 :   0 - 0x0
      13'hD4D: dout  = 8'b00000000; // 3405 :   0 - 0x0
      13'hD4E: dout  = 8'b00000000; // 3406 :   0 - 0x0
      13'hD4F: dout  = 8'b00000000; // 3407 :   0 - 0x0
      13'hD50: dout  = 8'b00000000; // 3408 :   0 - 0x0 -- Sprite 0xd5
      13'hD51: dout  = 8'b00000000; // 3409 :   0 - 0x0
      13'hD52: dout  = 8'b00000000; // 3410 :   0 - 0x0
      13'hD53: dout  = 8'b00000000; // 3411 :   0 - 0x0
      13'hD54: dout  = 8'b00000000; // 3412 :   0 - 0x0
      13'hD55: dout  = 8'b00000000; // 3413 :   0 - 0x0
      13'hD56: dout  = 8'b00000000; // 3414 :   0 - 0x0
      13'hD57: dout  = 8'b00000000; // 3415 :   0 - 0x0
      13'hD58: dout  = 8'b00000000; // 3416 :   0 - 0x0
      13'hD59: dout  = 8'b00000000; // 3417 :   0 - 0x0
      13'hD5A: dout  = 8'b00000000; // 3418 :   0 - 0x0
      13'hD5B: dout  = 8'b00000000; // 3419 :   0 - 0x0
      13'hD5C: dout  = 8'b00000000; // 3420 :   0 - 0x0
      13'hD5D: dout  = 8'b00000000; // 3421 :   0 - 0x0
      13'hD5E: dout  = 8'b00000000; // 3422 :   0 - 0x0
      13'hD5F: dout  = 8'b00000000; // 3423 :   0 - 0x0
      13'hD60: dout  = 8'b00000000; // 3424 :   0 - 0x0 -- Sprite 0xd6
      13'hD61: dout  = 8'b00000000; // 3425 :   0 - 0x0
      13'hD62: dout  = 8'b00000000; // 3426 :   0 - 0x0
      13'hD63: dout  = 8'b00000000; // 3427 :   0 - 0x0
      13'hD64: dout  = 8'b00000000; // 3428 :   0 - 0x0
      13'hD65: dout  = 8'b00000000; // 3429 :   0 - 0x0
      13'hD66: dout  = 8'b00000000; // 3430 :   0 - 0x0
      13'hD67: dout  = 8'b00000000; // 3431 :   0 - 0x0
      13'hD68: dout  = 8'b00000000; // 3432 :   0 - 0x0
      13'hD69: dout  = 8'b00000000; // 3433 :   0 - 0x0
      13'hD6A: dout  = 8'b00000000; // 3434 :   0 - 0x0
      13'hD6B: dout  = 8'b00000000; // 3435 :   0 - 0x0
      13'hD6C: dout  = 8'b00000000; // 3436 :   0 - 0x0
      13'hD6D: dout  = 8'b00000000; // 3437 :   0 - 0x0
      13'hD6E: dout  = 8'b00000000; // 3438 :   0 - 0x0
      13'hD6F: dout  = 8'b00000000; // 3439 :   0 - 0x0
      13'hD70: dout  = 8'b00000000; // 3440 :   0 - 0x0 -- Sprite 0xd7
      13'hD71: dout  = 8'b00000000; // 3441 :   0 - 0x0
      13'hD72: dout  = 8'b00000000; // 3442 :   0 - 0x0
      13'hD73: dout  = 8'b00000000; // 3443 :   0 - 0x0
      13'hD74: dout  = 8'b00000000; // 3444 :   0 - 0x0
      13'hD75: dout  = 8'b00000000; // 3445 :   0 - 0x0
      13'hD76: dout  = 8'b00000000; // 3446 :   0 - 0x0
      13'hD77: dout  = 8'b00000000; // 3447 :   0 - 0x0
      13'hD78: dout  = 8'b00000000; // 3448 :   0 - 0x0
      13'hD79: dout  = 8'b00000000; // 3449 :   0 - 0x0
      13'hD7A: dout  = 8'b00000000; // 3450 :   0 - 0x0
      13'hD7B: dout  = 8'b00000000; // 3451 :   0 - 0x0
      13'hD7C: dout  = 8'b00000000; // 3452 :   0 - 0x0
      13'hD7D: dout  = 8'b00000000; // 3453 :   0 - 0x0
      13'hD7E: dout  = 8'b00000000; // 3454 :   0 - 0x0
      13'hD7F: dout  = 8'b00000000; // 3455 :   0 - 0x0
      13'hD80: dout  = 8'b00000000; // 3456 :   0 - 0x0 -- Sprite 0xd8
      13'hD81: dout  = 8'b00000000; // 3457 :   0 - 0x0
      13'hD82: dout  = 8'b00000000; // 3458 :   0 - 0x0
      13'hD83: dout  = 8'b00000000; // 3459 :   0 - 0x0
      13'hD84: dout  = 8'b00000000; // 3460 :   0 - 0x0
      13'hD85: dout  = 8'b00000000; // 3461 :   0 - 0x0
      13'hD86: dout  = 8'b00000000; // 3462 :   0 - 0x0
      13'hD87: dout  = 8'b00000000; // 3463 :   0 - 0x0
      13'hD88: dout  = 8'b00000000; // 3464 :   0 - 0x0
      13'hD89: dout  = 8'b00000000; // 3465 :   0 - 0x0
      13'hD8A: dout  = 8'b00000000; // 3466 :   0 - 0x0
      13'hD8B: dout  = 8'b00000000; // 3467 :   0 - 0x0
      13'hD8C: dout  = 8'b00000000; // 3468 :   0 - 0x0
      13'hD8D: dout  = 8'b00000000; // 3469 :   0 - 0x0
      13'hD8E: dout  = 8'b00000000; // 3470 :   0 - 0x0
      13'hD8F: dout  = 8'b00000000; // 3471 :   0 - 0x0
      13'hD90: dout  = 8'b00000000; // 3472 :   0 - 0x0 -- Sprite 0xd9
      13'hD91: dout  = 8'b00000000; // 3473 :   0 - 0x0
      13'hD92: dout  = 8'b00000000; // 3474 :   0 - 0x0
      13'hD93: dout  = 8'b00000000; // 3475 :   0 - 0x0
      13'hD94: dout  = 8'b00000000; // 3476 :   0 - 0x0
      13'hD95: dout  = 8'b00000000; // 3477 :   0 - 0x0
      13'hD96: dout  = 8'b00000000; // 3478 :   0 - 0x0
      13'hD97: dout  = 8'b00000000; // 3479 :   0 - 0x0
      13'hD98: dout  = 8'b00000000; // 3480 :   0 - 0x0
      13'hD99: dout  = 8'b00000000; // 3481 :   0 - 0x0
      13'hD9A: dout  = 8'b00000000; // 3482 :   0 - 0x0
      13'hD9B: dout  = 8'b00000000; // 3483 :   0 - 0x0
      13'hD9C: dout  = 8'b00000000; // 3484 :   0 - 0x0
      13'hD9D: dout  = 8'b00000000; // 3485 :   0 - 0x0
      13'hD9E: dout  = 8'b00000000; // 3486 :   0 - 0x0
      13'hD9F: dout  = 8'b00000000; // 3487 :   0 - 0x0
      13'hDA0: dout  = 8'b00000000; // 3488 :   0 - 0x0 -- Sprite 0xda
      13'hDA1: dout  = 8'b00000000; // 3489 :   0 - 0x0
      13'hDA2: dout  = 8'b00000000; // 3490 :   0 - 0x0
      13'hDA3: dout  = 8'b00000000; // 3491 :   0 - 0x0
      13'hDA4: dout  = 8'b00000000; // 3492 :   0 - 0x0
      13'hDA5: dout  = 8'b00000000; // 3493 :   0 - 0x0
      13'hDA6: dout  = 8'b00000000; // 3494 :   0 - 0x0
      13'hDA7: dout  = 8'b00000000; // 3495 :   0 - 0x0
      13'hDA8: dout  = 8'b00000000; // 3496 :   0 - 0x0
      13'hDA9: dout  = 8'b00000000; // 3497 :   0 - 0x0
      13'hDAA: dout  = 8'b00000000; // 3498 :   0 - 0x0
      13'hDAB: dout  = 8'b00000000; // 3499 :   0 - 0x0
      13'hDAC: dout  = 8'b00000000; // 3500 :   0 - 0x0
      13'hDAD: dout  = 8'b00000000; // 3501 :   0 - 0x0
      13'hDAE: dout  = 8'b00000000; // 3502 :   0 - 0x0
      13'hDAF: dout  = 8'b00000000; // 3503 :   0 - 0x0
      13'hDB0: dout  = 8'b00000000; // 3504 :   0 - 0x0 -- Sprite 0xdb
      13'hDB1: dout  = 8'b00000000; // 3505 :   0 - 0x0
      13'hDB2: dout  = 8'b00000000; // 3506 :   0 - 0x0
      13'hDB3: dout  = 8'b00000000; // 3507 :   0 - 0x0
      13'hDB4: dout  = 8'b00000000; // 3508 :   0 - 0x0
      13'hDB5: dout  = 8'b00000000; // 3509 :   0 - 0x0
      13'hDB6: dout  = 8'b00000000; // 3510 :   0 - 0x0
      13'hDB7: dout  = 8'b00000000; // 3511 :   0 - 0x0
      13'hDB8: dout  = 8'b00000000; // 3512 :   0 - 0x0
      13'hDB9: dout  = 8'b00000000; // 3513 :   0 - 0x0
      13'hDBA: dout  = 8'b00000000; // 3514 :   0 - 0x0
      13'hDBB: dout  = 8'b00000000; // 3515 :   0 - 0x0
      13'hDBC: dout  = 8'b00000000; // 3516 :   0 - 0x0
      13'hDBD: dout  = 8'b00000000; // 3517 :   0 - 0x0
      13'hDBE: dout  = 8'b00000000; // 3518 :   0 - 0x0
      13'hDBF: dout  = 8'b00000000; // 3519 :   0 - 0x0
      13'hDC0: dout  = 8'b00000000; // 3520 :   0 - 0x0 -- Sprite 0xdc
      13'hDC1: dout  = 8'b00000000; // 3521 :   0 - 0x0
      13'hDC2: dout  = 8'b00000000; // 3522 :   0 - 0x0
      13'hDC3: dout  = 8'b00000000; // 3523 :   0 - 0x0
      13'hDC4: dout  = 8'b00000000; // 3524 :   0 - 0x0
      13'hDC5: dout  = 8'b00000000; // 3525 :   0 - 0x0
      13'hDC6: dout  = 8'b00000000; // 3526 :   0 - 0x0
      13'hDC7: dout  = 8'b00000000; // 3527 :   0 - 0x0
      13'hDC8: dout  = 8'b00000000; // 3528 :   0 - 0x0
      13'hDC9: dout  = 8'b00000000; // 3529 :   0 - 0x0
      13'hDCA: dout  = 8'b00000000; // 3530 :   0 - 0x0
      13'hDCB: dout  = 8'b00000000; // 3531 :   0 - 0x0
      13'hDCC: dout  = 8'b00000000; // 3532 :   0 - 0x0
      13'hDCD: dout  = 8'b00000000; // 3533 :   0 - 0x0
      13'hDCE: dout  = 8'b00000000; // 3534 :   0 - 0x0
      13'hDCF: dout  = 8'b00000000; // 3535 :   0 - 0x0
      13'hDD0: dout  = 8'b00000000; // 3536 :   0 - 0x0 -- Sprite 0xdd
      13'hDD1: dout  = 8'b00000000; // 3537 :   0 - 0x0
      13'hDD2: dout  = 8'b00000000; // 3538 :   0 - 0x0
      13'hDD3: dout  = 8'b00000000; // 3539 :   0 - 0x0
      13'hDD4: dout  = 8'b00000000; // 3540 :   0 - 0x0
      13'hDD5: dout  = 8'b00000000; // 3541 :   0 - 0x0
      13'hDD6: dout  = 8'b00000000; // 3542 :   0 - 0x0
      13'hDD7: dout  = 8'b00000000; // 3543 :   0 - 0x0
      13'hDD8: dout  = 8'b00000000; // 3544 :   0 - 0x0
      13'hDD9: dout  = 8'b00000000; // 3545 :   0 - 0x0
      13'hDDA: dout  = 8'b00000000; // 3546 :   0 - 0x0
      13'hDDB: dout  = 8'b00000000; // 3547 :   0 - 0x0
      13'hDDC: dout  = 8'b00000000; // 3548 :   0 - 0x0
      13'hDDD: dout  = 8'b00000000; // 3549 :   0 - 0x0
      13'hDDE: dout  = 8'b00000000; // 3550 :   0 - 0x0
      13'hDDF: dout  = 8'b00000000; // 3551 :   0 - 0x0
      13'hDE0: dout  = 8'b00000000; // 3552 :   0 - 0x0 -- Sprite 0xde
      13'hDE1: dout  = 8'b00000000; // 3553 :   0 - 0x0
      13'hDE2: dout  = 8'b00000000; // 3554 :   0 - 0x0
      13'hDE3: dout  = 8'b00000000; // 3555 :   0 - 0x0
      13'hDE4: dout  = 8'b00000000; // 3556 :   0 - 0x0
      13'hDE5: dout  = 8'b00000000; // 3557 :   0 - 0x0
      13'hDE6: dout  = 8'b00000000; // 3558 :   0 - 0x0
      13'hDE7: dout  = 8'b00000000; // 3559 :   0 - 0x0
      13'hDE8: dout  = 8'b00000000; // 3560 :   0 - 0x0
      13'hDE9: dout  = 8'b00000000; // 3561 :   0 - 0x0
      13'hDEA: dout  = 8'b00000000; // 3562 :   0 - 0x0
      13'hDEB: dout  = 8'b00000000; // 3563 :   0 - 0x0
      13'hDEC: dout  = 8'b00000000; // 3564 :   0 - 0x0
      13'hDED: dout  = 8'b00000000; // 3565 :   0 - 0x0
      13'hDEE: dout  = 8'b00000000; // 3566 :   0 - 0x0
      13'hDEF: dout  = 8'b00000000; // 3567 :   0 - 0x0
      13'hDF0: dout  = 8'b00000000; // 3568 :   0 - 0x0 -- Sprite 0xdf
      13'hDF1: dout  = 8'b00000000; // 3569 :   0 - 0x0
      13'hDF2: dout  = 8'b00000000; // 3570 :   0 - 0x0
      13'hDF3: dout  = 8'b00000000; // 3571 :   0 - 0x0
      13'hDF4: dout  = 8'b00000000; // 3572 :   0 - 0x0
      13'hDF5: dout  = 8'b00000000; // 3573 :   0 - 0x0
      13'hDF6: dout  = 8'b00000000; // 3574 :   0 - 0x0
      13'hDF7: dout  = 8'b00000000; // 3575 :   0 - 0x0
      13'hDF8: dout  = 8'b00000000; // 3576 :   0 - 0x0
      13'hDF9: dout  = 8'b00000000; // 3577 :   0 - 0x0
      13'hDFA: dout  = 8'b00000000; // 3578 :   0 - 0x0
      13'hDFB: dout  = 8'b00000000; // 3579 :   0 - 0x0
      13'hDFC: dout  = 8'b00000000; // 3580 :   0 - 0x0
      13'hDFD: dout  = 8'b00000000; // 3581 :   0 - 0x0
      13'hDFE: dout  = 8'b00000000; // 3582 :   0 - 0x0
      13'hDFF: dout  = 8'b00000000; // 3583 :   0 - 0x0
      13'hE00: dout  = 8'b00000000; // 3584 :   0 - 0x0 -- Sprite 0xe0
      13'hE01: dout  = 8'b00000000; // 3585 :   0 - 0x0
      13'hE02: dout  = 8'b00000000; // 3586 :   0 - 0x0
      13'hE03: dout  = 8'b00000000; // 3587 :   0 - 0x0
      13'hE04: dout  = 8'b00000000; // 3588 :   0 - 0x0
      13'hE05: dout  = 8'b00000000; // 3589 :   0 - 0x0
      13'hE06: dout  = 8'b00000000; // 3590 :   0 - 0x0
      13'hE07: dout  = 8'b00000000; // 3591 :   0 - 0x0
      13'hE08: dout  = 8'b00000000; // 3592 :   0 - 0x0
      13'hE09: dout  = 8'b00000000; // 3593 :   0 - 0x0
      13'hE0A: dout  = 8'b00000000; // 3594 :   0 - 0x0
      13'hE0B: dout  = 8'b00000000; // 3595 :   0 - 0x0
      13'hE0C: dout  = 8'b00000000; // 3596 :   0 - 0x0
      13'hE0D: dout  = 8'b00000000; // 3597 :   0 - 0x0
      13'hE0E: dout  = 8'b00000000; // 3598 :   0 - 0x0
      13'hE0F: dout  = 8'b00000000; // 3599 :   0 - 0x0
      13'hE10: dout  = 8'b00000000; // 3600 :   0 - 0x0 -- Sprite 0xe1
      13'hE11: dout  = 8'b00000000; // 3601 :   0 - 0x0
      13'hE12: dout  = 8'b00000000; // 3602 :   0 - 0x0
      13'hE13: dout  = 8'b00000000; // 3603 :   0 - 0x0
      13'hE14: dout  = 8'b00000000; // 3604 :   0 - 0x0
      13'hE15: dout  = 8'b00000000; // 3605 :   0 - 0x0
      13'hE16: dout  = 8'b00000000; // 3606 :   0 - 0x0
      13'hE17: dout  = 8'b00000000; // 3607 :   0 - 0x0
      13'hE18: dout  = 8'b00000000; // 3608 :   0 - 0x0
      13'hE19: dout  = 8'b00000000; // 3609 :   0 - 0x0
      13'hE1A: dout  = 8'b00000000; // 3610 :   0 - 0x0
      13'hE1B: dout  = 8'b00000000; // 3611 :   0 - 0x0
      13'hE1C: dout  = 8'b00000000; // 3612 :   0 - 0x0
      13'hE1D: dout  = 8'b00000000; // 3613 :   0 - 0x0
      13'hE1E: dout  = 8'b00000000; // 3614 :   0 - 0x0
      13'hE1F: dout  = 8'b00000000; // 3615 :   0 - 0x0
      13'hE20: dout  = 8'b00000000; // 3616 :   0 - 0x0 -- Sprite 0xe2
      13'hE21: dout  = 8'b00000000; // 3617 :   0 - 0x0
      13'hE22: dout  = 8'b00000000; // 3618 :   0 - 0x0
      13'hE23: dout  = 8'b00000000; // 3619 :   0 - 0x0
      13'hE24: dout  = 8'b00000000; // 3620 :   0 - 0x0
      13'hE25: dout  = 8'b00000000; // 3621 :   0 - 0x0
      13'hE26: dout  = 8'b00000000; // 3622 :   0 - 0x0
      13'hE27: dout  = 8'b00000000; // 3623 :   0 - 0x0
      13'hE28: dout  = 8'b00000000; // 3624 :   0 - 0x0
      13'hE29: dout  = 8'b00000000; // 3625 :   0 - 0x0
      13'hE2A: dout  = 8'b00000000; // 3626 :   0 - 0x0
      13'hE2B: dout  = 8'b00000000; // 3627 :   0 - 0x0
      13'hE2C: dout  = 8'b00000000; // 3628 :   0 - 0x0
      13'hE2D: dout  = 8'b00000000; // 3629 :   0 - 0x0
      13'hE2E: dout  = 8'b00000000; // 3630 :   0 - 0x0
      13'hE2F: dout  = 8'b00000000; // 3631 :   0 - 0x0
      13'hE30: dout  = 8'b00000000; // 3632 :   0 - 0x0 -- Sprite 0xe3
      13'hE31: dout  = 8'b00000000; // 3633 :   0 - 0x0
      13'hE32: dout  = 8'b00000000; // 3634 :   0 - 0x0
      13'hE33: dout  = 8'b00000000; // 3635 :   0 - 0x0
      13'hE34: dout  = 8'b00000000; // 3636 :   0 - 0x0
      13'hE35: dout  = 8'b00000000; // 3637 :   0 - 0x0
      13'hE36: dout  = 8'b00000000; // 3638 :   0 - 0x0
      13'hE37: dout  = 8'b00000000; // 3639 :   0 - 0x0
      13'hE38: dout  = 8'b00000000; // 3640 :   0 - 0x0
      13'hE39: dout  = 8'b00000000; // 3641 :   0 - 0x0
      13'hE3A: dout  = 8'b00000000; // 3642 :   0 - 0x0
      13'hE3B: dout  = 8'b00000000; // 3643 :   0 - 0x0
      13'hE3C: dout  = 8'b00000000; // 3644 :   0 - 0x0
      13'hE3D: dout  = 8'b00000000; // 3645 :   0 - 0x0
      13'hE3E: dout  = 8'b00000000; // 3646 :   0 - 0x0
      13'hE3F: dout  = 8'b00000000; // 3647 :   0 - 0x0
      13'hE40: dout  = 8'b00000000; // 3648 :   0 - 0x0 -- Sprite 0xe4
      13'hE41: dout  = 8'b00000000; // 3649 :   0 - 0x0
      13'hE42: dout  = 8'b00000000; // 3650 :   0 - 0x0
      13'hE43: dout  = 8'b00000000; // 3651 :   0 - 0x0
      13'hE44: dout  = 8'b00000000; // 3652 :   0 - 0x0
      13'hE45: dout  = 8'b00000000; // 3653 :   0 - 0x0
      13'hE46: dout  = 8'b00000000; // 3654 :   0 - 0x0
      13'hE47: dout  = 8'b00000000; // 3655 :   0 - 0x0
      13'hE48: dout  = 8'b00000000; // 3656 :   0 - 0x0
      13'hE49: dout  = 8'b00000000; // 3657 :   0 - 0x0
      13'hE4A: dout  = 8'b00000000; // 3658 :   0 - 0x0
      13'hE4B: dout  = 8'b00000000; // 3659 :   0 - 0x0
      13'hE4C: dout  = 8'b00000000; // 3660 :   0 - 0x0
      13'hE4D: dout  = 8'b00000000; // 3661 :   0 - 0x0
      13'hE4E: dout  = 8'b00000000; // 3662 :   0 - 0x0
      13'hE4F: dout  = 8'b00000000; // 3663 :   0 - 0x0
      13'hE50: dout  = 8'b00000000; // 3664 :   0 - 0x0 -- Sprite 0xe5
      13'hE51: dout  = 8'b00000000; // 3665 :   0 - 0x0
      13'hE52: dout  = 8'b00000000; // 3666 :   0 - 0x0
      13'hE53: dout  = 8'b00000000; // 3667 :   0 - 0x0
      13'hE54: dout  = 8'b00000000; // 3668 :   0 - 0x0
      13'hE55: dout  = 8'b00000000; // 3669 :   0 - 0x0
      13'hE56: dout  = 8'b00000000; // 3670 :   0 - 0x0
      13'hE57: dout  = 8'b00000000; // 3671 :   0 - 0x0
      13'hE58: dout  = 8'b00000000; // 3672 :   0 - 0x0
      13'hE59: dout  = 8'b00000000; // 3673 :   0 - 0x0
      13'hE5A: dout  = 8'b00000000; // 3674 :   0 - 0x0
      13'hE5B: dout  = 8'b00000000; // 3675 :   0 - 0x0
      13'hE5C: dout  = 8'b00000000; // 3676 :   0 - 0x0
      13'hE5D: dout  = 8'b00000000; // 3677 :   0 - 0x0
      13'hE5E: dout  = 8'b00000000; // 3678 :   0 - 0x0
      13'hE5F: dout  = 8'b00000000; // 3679 :   0 - 0x0
      13'hE60: dout  = 8'b00000000; // 3680 :   0 - 0x0 -- Sprite 0xe6
      13'hE61: dout  = 8'b00000000; // 3681 :   0 - 0x0
      13'hE62: dout  = 8'b00000000; // 3682 :   0 - 0x0
      13'hE63: dout  = 8'b00000000; // 3683 :   0 - 0x0
      13'hE64: dout  = 8'b00000000; // 3684 :   0 - 0x0
      13'hE65: dout  = 8'b00000000; // 3685 :   0 - 0x0
      13'hE66: dout  = 8'b00000000; // 3686 :   0 - 0x0
      13'hE67: dout  = 8'b00000000; // 3687 :   0 - 0x0
      13'hE68: dout  = 8'b00000000; // 3688 :   0 - 0x0
      13'hE69: dout  = 8'b00000000; // 3689 :   0 - 0x0
      13'hE6A: dout  = 8'b00000000; // 3690 :   0 - 0x0
      13'hE6B: dout  = 8'b00000000; // 3691 :   0 - 0x0
      13'hE6C: dout  = 8'b00000000; // 3692 :   0 - 0x0
      13'hE6D: dout  = 8'b00000000; // 3693 :   0 - 0x0
      13'hE6E: dout  = 8'b00000000; // 3694 :   0 - 0x0
      13'hE6F: dout  = 8'b00000000; // 3695 :   0 - 0x0
      13'hE70: dout  = 8'b00000000; // 3696 :   0 - 0x0 -- Sprite 0xe7
      13'hE71: dout  = 8'b00000000; // 3697 :   0 - 0x0
      13'hE72: dout  = 8'b00000000; // 3698 :   0 - 0x0
      13'hE73: dout  = 8'b00000000; // 3699 :   0 - 0x0
      13'hE74: dout  = 8'b00000000; // 3700 :   0 - 0x0
      13'hE75: dout  = 8'b00000000; // 3701 :   0 - 0x0
      13'hE76: dout  = 8'b00000000; // 3702 :   0 - 0x0
      13'hE77: dout  = 8'b00000000; // 3703 :   0 - 0x0
      13'hE78: dout  = 8'b00000000; // 3704 :   0 - 0x0
      13'hE79: dout  = 8'b00000000; // 3705 :   0 - 0x0
      13'hE7A: dout  = 8'b00000000; // 3706 :   0 - 0x0
      13'hE7B: dout  = 8'b00000000; // 3707 :   0 - 0x0
      13'hE7C: dout  = 8'b00000000; // 3708 :   0 - 0x0
      13'hE7D: dout  = 8'b00000000; // 3709 :   0 - 0x0
      13'hE7E: dout  = 8'b00000000; // 3710 :   0 - 0x0
      13'hE7F: dout  = 8'b00000000; // 3711 :   0 - 0x0
      13'hE80: dout  = 8'b00000000; // 3712 :   0 - 0x0 -- Sprite 0xe8
      13'hE81: dout  = 8'b00000000; // 3713 :   0 - 0x0
      13'hE82: dout  = 8'b00000000; // 3714 :   0 - 0x0
      13'hE83: dout  = 8'b00000000; // 3715 :   0 - 0x0
      13'hE84: dout  = 8'b00000000; // 3716 :   0 - 0x0
      13'hE85: dout  = 8'b00000000; // 3717 :   0 - 0x0
      13'hE86: dout  = 8'b00000000; // 3718 :   0 - 0x0
      13'hE87: dout  = 8'b00000000; // 3719 :   0 - 0x0
      13'hE88: dout  = 8'b00000000; // 3720 :   0 - 0x0
      13'hE89: dout  = 8'b00000000; // 3721 :   0 - 0x0
      13'hE8A: dout  = 8'b00000000; // 3722 :   0 - 0x0
      13'hE8B: dout  = 8'b00000000; // 3723 :   0 - 0x0
      13'hE8C: dout  = 8'b00000000; // 3724 :   0 - 0x0
      13'hE8D: dout  = 8'b00000000; // 3725 :   0 - 0x0
      13'hE8E: dout  = 8'b00000000; // 3726 :   0 - 0x0
      13'hE8F: dout  = 8'b00000000; // 3727 :   0 - 0x0
      13'hE90: dout  = 8'b00000000; // 3728 :   0 - 0x0 -- Sprite 0xe9
      13'hE91: dout  = 8'b00000000; // 3729 :   0 - 0x0
      13'hE92: dout  = 8'b00000000; // 3730 :   0 - 0x0
      13'hE93: dout  = 8'b00000000; // 3731 :   0 - 0x0
      13'hE94: dout  = 8'b00000000; // 3732 :   0 - 0x0
      13'hE95: dout  = 8'b00000000; // 3733 :   0 - 0x0
      13'hE96: dout  = 8'b00000000; // 3734 :   0 - 0x0
      13'hE97: dout  = 8'b00000000; // 3735 :   0 - 0x0
      13'hE98: dout  = 8'b00000000; // 3736 :   0 - 0x0
      13'hE99: dout  = 8'b00000000; // 3737 :   0 - 0x0
      13'hE9A: dout  = 8'b00000000; // 3738 :   0 - 0x0
      13'hE9B: dout  = 8'b00000000; // 3739 :   0 - 0x0
      13'hE9C: dout  = 8'b00000000; // 3740 :   0 - 0x0
      13'hE9D: dout  = 8'b00000000; // 3741 :   0 - 0x0
      13'hE9E: dout  = 8'b00000000; // 3742 :   0 - 0x0
      13'hE9F: dout  = 8'b00000000; // 3743 :   0 - 0x0
      13'hEA0: dout  = 8'b00000000; // 3744 :   0 - 0x0 -- Sprite 0xea
      13'hEA1: dout  = 8'b00000000; // 3745 :   0 - 0x0
      13'hEA2: dout  = 8'b00000000; // 3746 :   0 - 0x0
      13'hEA3: dout  = 8'b00000000; // 3747 :   0 - 0x0
      13'hEA4: dout  = 8'b00000000; // 3748 :   0 - 0x0
      13'hEA5: dout  = 8'b00000000; // 3749 :   0 - 0x0
      13'hEA6: dout  = 8'b00000000; // 3750 :   0 - 0x0
      13'hEA7: dout  = 8'b00000000; // 3751 :   0 - 0x0
      13'hEA8: dout  = 8'b00000000; // 3752 :   0 - 0x0
      13'hEA9: dout  = 8'b00000000; // 3753 :   0 - 0x0
      13'hEAA: dout  = 8'b00000000; // 3754 :   0 - 0x0
      13'hEAB: dout  = 8'b00000000; // 3755 :   0 - 0x0
      13'hEAC: dout  = 8'b00000000; // 3756 :   0 - 0x0
      13'hEAD: dout  = 8'b00000000; // 3757 :   0 - 0x0
      13'hEAE: dout  = 8'b00000000; // 3758 :   0 - 0x0
      13'hEAF: dout  = 8'b00000000; // 3759 :   0 - 0x0
      13'hEB0: dout  = 8'b00000000; // 3760 :   0 - 0x0 -- Sprite 0xeb
      13'hEB1: dout  = 8'b00000000; // 3761 :   0 - 0x0
      13'hEB2: dout  = 8'b00000000; // 3762 :   0 - 0x0
      13'hEB3: dout  = 8'b00000000; // 3763 :   0 - 0x0
      13'hEB4: dout  = 8'b00000000; // 3764 :   0 - 0x0
      13'hEB5: dout  = 8'b00000000; // 3765 :   0 - 0x0
      13'hEB6: dout  = 8'b00000000; // 3766 :   0 - 0x0
      13'hEB7: dout  = 8'b00000000; // 3767 :   0 - 0x0
      13'hEB8: dout  = 8'b00000000; // 3768 :   0 - 0x0
      13'hEB9: dout  = 8'b00000000; // 3769 :   0 - 0x0
      13'hEBA: dout  = 8'b00000000; // 3770 :   0 - 0x0
      13'hEBB: dout  = 8'b00000000; // 3771 :   0 - 0x0
      13'hEBC: dout  = 8'b00000000; // 3772 :   0 - 0x0
      13'hEBD: dout  = 8'b00000000; // 3773 :   0 - 0x0
      13'hEBE: dout  = 8'b00000000; // 3774 :   0 - 0x0
      13'hEBF: dout  = 8'b00000000; // 3775 :   0 - 0x0
      13'hEC0: dout  = 8'b00000000; // 3776 :   0 - 0x0 -- Sprite 0xec
      13'hEC1: dout  = 8'b00000000; // 3777 :   0 - 0x0
      13'hEC2: dout  = 8'b00000000; // 3778 :   0 - 0x0
      13'hEC3: dout  = 8'b00000000; // 3779 :   0 - 0x0
      13'hEC4: dout  = 8'b00000000; // 3780 :   0 - 0x0
      13'hEC5: dout  = 8'b00000000; // 3781 :   0 - 0x0
      13'hEC6: dout  = 8'b00000000; // 3782 :   0 - 0x0
      13'hEC7: dout  = 8'b00000000; // 3783 :   0 - 0x0
      13'hEC8: dout  = 8'b00000000; // 3784 :   0 - 0x0
      13'hEC9: dout  = 8'b00000000; // 3785 :   0 - 0x0
      13'hECA: dout  = 8'b00000000; // 3786 :   0 - 0x0
      13'hECB: dout  = 8'b00000000; // 3787 :   0 - 0x0
      13'hECC: dout  = 8'b00000000; // 3788 :   0 - 0x0
      13'hECD: dout  = 8'b00000000; // 3789 :   0 - 0x0
      13'hECE: dout  = 8'b00000000; // 3790 :   0 - 0x0
      13'hECF: dout  = 8'b00000000; // 3791 :   0 - 0x0
      13'hED0: dout  = 8'b00000000; // 3792 :   0 - 0x0 -- Sprite 0xed
      13'hED1: dout  = 8'b00000000; // 3793 :   0 - 0x0
      13'hED2: dout  = 8'b00000000; // 3794 :   0 - 0x0
      13'hED3: dout  = 8'b00000000; // 3795 :   0 - 0x0
      13'hED4: dout  = 8'b00000000; // 3796 :   0 - 0x0
      13'hED5: dout  = 8'b00000000; // 3797 :   0 - 0x0
      13'hED6: dout  = 8'b00000000; // 3798 :   0 - 0x0
      13'hED7: dout  = 8'b00000000; // 3799 :   0 - 0x0
      13'hED8: dout  = 8'b00000000; // 3800 :   0 - 0x0
      13'hED9: dout  = 8'b00000000; // 3801 :   0 - 0x0
      13'hEDA: dout  = 8'b00000000; // 3802 :   0 - 0x0
      13'hEDB: dout  = 8'b00000000; // 3803 :   0 - 0x0
      13'hEDC: dout  = 8'b00000000; // 3804 :   0 - 0x0
      13'hEDD: dout  = 8'b00000000; // 3805 :   0 - 0x0
      13'hEDE: dout  = 8'b00000000; // 3806 :   0 - 0x0
      13'hEDF: dout  = 8'b00000000; // 3807 :   0 - 0x0
      13'hEE0: dout  = 8'b00000000; // 3808 :   0 - 0x0 -- Sprite 0xee
      13'hEE1: dout  = 8'b00000000; // 3809 :   0 - 0x0
      13'hEE2: dout  = 8'b00000000; // 3810 :   0 - 0x0
      13'hEE3: dout  = 8'b00000000; // 3811 :   0 - 0x0
      13'hEE4: dout  = 8'b00000000; // 3812 :   0 - 0x0
      13'hEE5: dout  = 8'b00000000; // 3813 :   0 - 0x0
      13'hEE6: dout  = 8'b00000000; // 3814 :   0 - 0x0
      13'hEE7: dout  = 8'b00000000; // 3815 :   0 - 0x0
      13'hEE8: dout  = 8'b00000000; // 3816 :   0 - 0x0
      13'hEE9: dout  = 8'b00000000; // 3817 :   0 - 0x0
      13'hEEA: dout  = 8'b00000000; // 3818 :   0 - 0x0
      13'hEEB: dout  = 8'b00000000; // 3819 :   0 - 0x0
      13'hEEC: dout  = 8'b00000000; // 3820 :   0 - 0x0
      13'hEED: dout  = 8'b00000000; // 3821 :   0 - 0x0
      13'hEEE: dout  = 8'b00000000; // 3822 :   0 - 0x0
      13'hEEF: dout  = 8'b00000000; // 3823 :   0 - 0x0
      13'hEF0: dout  = 8'b00000000; // 3824 :   0 - 0x0 -- Sprite 0xef
      13'hEF1: dout  = 8'b00000000; // 3825 :   0 - 0x0
      13'hEF2: dout  = 8'b00000000; // 3826 :   0 - 0x0
      13'hEF3: dout  = 8'b00000000; // 3827 :   0 - 0x0
      13'hEF4: dout  = 8'b00000000; // 3828 :   0 - 0x0
      13'hEF5: dout  = 8'b00000000; // 3829 :   0 - 0x0
      13'hEF6: dout  = 8'b00000000; // 3830 :   0 - 0x0
      13'hEF7: dout  = 8'b00000000; // 3831 :   0 - 0x0
      13'hEF8: dout  = 8'b00000000; // 3832 :   0 - 0x0
      13'hEF9: dout  = 8'b00000000; // 3833 :   0 - 0x0
      13'hEFA: dout  = 8'b00000000; // 3834 :   0 - 0x0
      13'hEFB: dout  = 8'b00000000; // 3835 :   0 - 0x0
      13'hEFC: dout  = 8'b00000000; // 3836 :   0 - 0x0
      13'hEFD: dout  = 8'b00000000; // 3837 :   0 - 0x0
      13'hEFE: dout  = 8'b00000000; // 3838 :   0 - 0x0
      13'hEFF: dout  = 8'b00000000; // 3839 :   0 - 0x0
      13'hF00: dout  = 8'b00000000; // 3840 :   0 - 0x0 -- Sprite 0xf0
      13'hF01: dout  = 8'b00000000; // 3841 :   0 - 0x0
      13'hF02: dout  = 8'b00000000; // 3842 :   0 - 0x0
      13'hF03: dout  = 8'b00000000; // 3843 :   0 - 0x0
      13'hF04: dout  = 8'b00000000; // 3844 :   0 - 0x0
      13'hF05: dout  = 8'b00000000; // 3845 :   0 - 0x0
      13'hF06: dout  = 8'b00000000; // 3846 :   0 - 0x0
      13'hF07: dout  = 8'b00000000; // 3847 :   0 - 0x0
      13'hF08: dout  = 8'b00000000; // 3848 :   0 - 0x0
      13'hF09: dout  = 8'b00000000; // 3849 :   0 - 0x0
      13'hF0A: dout  = 8'b00000000; // 3850 :   0 - 0x0
      13'hF0B: dout  = 8'b00000000; // 3851 :   0 - 0x0
      13'hF0C: dout  = 8'b00000000; // 3852 :   0 - 0x0
      13'hF0D: dout  = 8'b00000000; // 3853 :   0 - 0x0
      13'hF0E: dout  = 8'b00000000; // 3854 :   0 - 0x0
      13'hF0F: dout  = 8'b00000000; // 3855 :   0 - 0x0
      13'hF10: dout  = 8'b00000000; // 3856 :   0 - 0x0 -- Sprite 0xf1
      13'hF11: dout  = 8'b00000000; // 3857 :   0 - 0x0
      13'hF12: dout  = 8'b00000000; // 3858 :   0 - 0x0
      13'hF13: dout  = 8'b00000000; // 3859 :   0 - 0x0
      13'hF14: dout  = 8'b00000000; // 3860 :   0 - 0x0
      13'hF15: dout  = 8'b00000000; // 3861 :   0 - 0x0
      13'hF16: dout  = 8'b00000000; // 3862 :   0 - 0x0
      13'hF17: dout  = 8'b00000000; // 3863 :   0 - 0x0
      13'hF18: dout  = 8'b00000000; // 3864 :   0 - 0x0
      13'hF19: dout  = 8'b00000000; // 3865 :   0 - 0x0
      13'hF1A: dout  = 8'b00000000; // 3866 :   0 - 0x0
      13'hF1B: dout  = 8'b00000000; // 3867 :   0 - 0x0
      13'hF1C: dout  = 8'b00000000; // 3868 :   0 - 0x0
      13'hF1D: dout  = 8'b00000000; // 3869 :   0 - 0x0
      13'hF1E: dout  = 8'b00000000; // 3870 :   0 - 0x0
      13'hF1F: dout  = 8'b00000000; // 3871 :   0 - 0x0
      13'hF20: dout  = 8'b00000000; // 3872 :   0 - 0x0 -- Sprite 0xf2
      13'hF21: dout  = 8'b00000000; // 3873 :   0 - 0x0
      13'hF22: dout  = 8'b00000000; // 3874 :   0 - 0x0
      13'hF23: dout  = 8'b00000000; // 3875 :   0 - 0x0
      13'hF24: dout  = 8'b00000000; // 3876 :   0 - 0x0
      13'hF25: dout  = 8'b00000000; // 3877 :   0 - 0x0
      13'hF26: dout  = 8'b00000000; // 3878 :   0 - 0x0
      13'hF27: dout  = 8'b00000000; // 3879 :   0 - 0x0
      13'hF28: dout  = 8'b00000000; // 3880 :   0 - 0x0
      13'hF29: dout  = 8'b00000000; // 3881 :   0 - 0x0
      13'hF2A: dout  = 8'b00000000; // 3882 :   0 - 0x0
      13'hF2B: dout  = 8'b00000000; // 3883 :   0 - 0x0
      13'hF2C: dout  = 8'b00000000; // 3884 :   0 - 0x0
      13'hF2D: dout  = 8'b00000000; // 3885 :   0 - 0x0
      13'hF2E: dout  = 8'b00000000; // 3886 :   0 - 0x0
      13'hF2F: dout  = 8'b00000000; // 3887 :   0 - 0x0
      13'hF30: dout  = 8'b00000000; // 3888 :   0 - 0x0 -- Sprite 0xf3
      13'hF31: dout  = 8'b00000000; // 3889 :   0 - 0x0
      13'hF32: dout  = 8'b00000000; // 3890 :   0 - 0x0
      13'hF33: dout  = 8'b00000000; // 3891 :   0 - 0x0
      13'hF34: dout  = 8'b00000000; // 3892 :   0 - 0x0
      13'hF35: dout  = 8'b00000000; // 3893 :   0 - 0x0
      13'hF36: dout  = 8'b00000000; // 3894 :   0 - 0x0
      13'hF37: dout  = 8'b00000000; // 3895 :   0 - 0x0
      13'hF38: dout  = 8'b00000000; // 3896 :   0 - 0x0
      13'hF39: dout  = 8'b00000000; // 3897 :   0 - 0x0
      13'hF3A: dout  = 8'b00000000; // 3898 :   0 - 0x0
      13'hF3B: dout  = 8'b00000000; // 3899 :   0 - 0x0
      13'hF3C: dout  = 8'b00000000; // 3900 :   0 - 0x0
      13'hF3D: dout  = 8'b00000000; // 3901 :   0 - 0x0
      13'hF3E: dout  = 8'b00000000; // 3902 :   0 - 0x0
      13'hF3F: dout  = 8'b00000000; // 3903 :   0 - 0x0
      13'hF40: dout  = 8'b00000000; // 3904 :   0 - 0x0 -- Sprite 0xf4
      13'hF41: dout  = 8'b00000000; // 3905 :   0 - 0x0
      13'hF42: dout  = 8'b00000000; // 3906 :   0 - 0x0
      13'hF43: dout  = 8'b00000000; // 3907 :   0 - 0x0
      13'hF44: dout  = 8'b00000000; // 3908 :   0 - 0x0
      13'hF45: dout  = 8'b00000000; // 3909 :   0 - 0x0
      13'hF46: dout  = 8'b00000000; // 3910 :   0 - 0x0
      13'hF47: dout  = 8'b00000000; // 3911 :   0 - 0x0
      13'hF48: dout  = 8'b00000000; // 3912 :   0 - 0x0
      13'hF49: dout  = 8'b00000000; // 3913 :   0 - 0x0
      13'hF4A: dout  = 8'b00000000; // 3914 :   0 - 0x0
      13'hF4B: dout  = 8'b00000000; // 3915 :   0 - 0x0
      13'hF4C: dout  = 8'b00000000; // 3916 :   0 - 0x0
      13'hF4D: dout  = 8'b00000000; // 3917 :   0 - 0x0
      13'hF4E: dout  = 8'b00000000; // 3918 :   0 - 0x0
      13'hF4F: dout  = 8'b00000000; // 3919 :   0 - 0x0
      13'hF50: dout  = 8'b00000000; // 3920 :   0 - 0x0 -- Sprite 0xf5
      13'hF51: dout  = 8'b00000000; // 3921 :   0 - 0x0
      13'hF52: dout  = 8'b00000000; // 3922 :   0 - 0x0
      13'hF53: dout  = 8'b00000000; // 3923 :   0 - 0x0
      13'hF54: dout  = 8'b00000000; // 3924 :   0 - 0x0
      13'hF55: dout  = 8'b00000000; // 3925 :   0 - 0x0
      13'hF56: dout  = 8'b00000000; // 3926 :   0 - 0x0
      13'hF57: dout  = 8'b00000000; // 3927 :   0 - 0x0
      13'hF58: dout  = 8'b00000000; // 3928 :   0 - 0x0
      13'hF59: dout  = 8'b00000000; // 3929 :   0 - 0x0
      13'hF5A: dout  = 8'b00000000; // 3930 :   0 - 0x0
      13'hF5B: dout  = 8'b00000000; // 3931 :   0 - 0x0
      13'hF5C: dout  = 8'b00000000; // 3932 :   0 - 0x0
      13'hF5D: dout  = 8'b00000000; // 3933 :   0 - 0x0
      13'hF5E: dout  = 8'b00000000; // 3934 :   0 - 0x0
      13'hF5F: dout  = 8'b00000000; // 3935 :   0 - 0x0
      13'hF60: dout  = 8'b00000000; // 3936 :   0 - 0x0 -- Sprite 0xf6
      13'hF61: dout  = 8'b00000000; // 3937 :   0 - 0x0
      13'hF62: dout  = 8'b00000000; // 3938 :   0 - 0x0
      13'hF63: dout  = 8'b00000000; // 3939 :   0 - 0x0
      13'hF64: dout  = 8'b00000000; // 3940 :   0 - 0x0
      13'hF65: dout  = 8'b00000000; // 3941 :   0 - 0x0
      13'hF66: dout  = 8'b00000000; // 3942 :   0 - 0x0
      13'hF67: dout  = 8'b00000000; // 3943 :   0 - 0x0
      13'hF68: dout  = 8'b00000000; // 3944 :   0 - 0x0
      13'hF69: dout  = 8'b00000000; // 3945 :   0 - 0x0
      13'hF6A: dout  = 8'b00000000; // 3946 :   0 - 0x0
      13'hF6B: dout  = 8'b00000000; // 3947 :   0 - 0x0
      13'hF6C: dout  = 8'b00000000; // 3948 :   0 - 0x0
      13'hF6D: dout  = 8'b00000000; // 3949 :   0 - 0x0
      13'hF6E: dout  = 8'b00000000; // 3950 :   0 - 0x0
      13'hF6F: dout  = 8'b00000000; // 3951 :   0 - 0x0
      13'hF70: dout  = 8'b00000000; // 3952 :   0 - 0x0 -- Sprite 0xf7
      13'hF71: dout  = 8'b00000000; // 3953 :   0 - 0x0
      13'hF72: dout  = 8'b00000000; // 3954 :   0 - 0x0
      13'hF73: dout  = 8'b00000000; // 3955 :   0 - 0x0
      13'hF74: dout  = 8'b00000000; // 3956 :   0 - 0x0
      13'hF75: dout  = 8'b00000000; // 3957 :   0 - 0x0
      13'hF76: dout  = 8'b00000000; // 3958 :   0 - 0x0
      13'hF77: dout  = 8'b00000000; // 3959 :   0 - 0x0
      13'hF78: dout  = 8'b00000000; // 3960 :   0 - 0x0
      13'hF79: dout  = 8'b00000000; // 3961 :   0 - 0x0
      13'hF7A: dout  = 8'b00000000; // 3962 :   0 - 0x0
      13'hF7B: dout  = 8'b00000000; // 3963 :   0 - 0x0
      13'hF7C: dout  = 8'b00000000; // 3964 :   0 - 0x0
      13'hF7D: dout  = 8'b00000000; // 3965 :   0 - 0x0
      13'hF7E: dout  = 8'b00000000; // 3966 :   0 - 0x0
      13'hF7F: dout  = 8'b00000000; // 3967 :   0 - 0x0
      13'hF80: dout  = 8'b00000000; // 3968 :   0 - 0x0 -- Sprite 0xf8
      13'hF81: dout  = 8'b00000000; // 3969 :   0 - 0x0
      13'hF82: dout  = 8'b00000000; // 3970 :   0 - 0x0
      13'hF83: dout  = 8'b00000000; // 3971 :   0 - 0x0
      13'hF84: dout  = 8'b00000000; // 3972 :   0 - 0x0
      13'hF85: dout  = 8'b00000000; // 3973 :   0 - 0x0
      13'hF86: dout  = 8'b00000000; // 3974 :   0 - 0x0
      13'hF87: dout  = 8'b00000000; // 3975 :   0 - 0x0
      13'hF88: dout  = 8'b00000000; // 3976 :   0 - 0x0
      13'hF89: dout  = 8'b00000000; // 3977 :   0 - 0x0
      13'hF8A: dout  = 8'b00000000; // 3978 :   0 - 0x0
      13'hF8B: dout  = 8'b00000000; // 3979 :   0 - 0x0
      13'hF8C: dout  = 8'b00000000; // 3980 :   0 - 0x0
      13'hF8D: dout  = 8'b00000000; // 3981 :   0 - 0x0
      13'hF8E: dout  = 8'b00000000; // 3982 :   0 - 0x0
      13'hF8F: dout  = 8'b00000000; // 3983 :   0 - 0x0
      13'hF90: dout  = 8'b00000000; // 3984 :   0 - 0x0 -- Sprite 0xf9
      13'hF91: dout  = 8'b00000000; // 3985 :   0 - 0x0
      13'hF92: dout  = 8'b00000000; // 3986 :   0 - 0x0
      13'hF93: dout  = 8'b00000000; // 3987 :   0 - 0x0
      13'hF94: dout  = 8'b00000000; // 3988 :   0 - 0x0
      13'hF95: dout  = 8'b00000000; // 3989 :   0 - 0x0
      13'hF96: dout  = 8'b00000000; // 3990 :   0 - 0x0
      13'hF97: dout  = 8'b00000000; // 3991 :   0 - 0x0
      13'hF98: dout  = 8'b00000000; // 3992 :   0 - 0x0
      13'hF99: dout  = 8'b00000000; // 3993 :   0 - 0x0
      13'hF9A: dout  = 8'b00000000; // 3994 :   0 - 0x0
      13'hF9B: dout  = 8'b00000000; // 3995 :   0 - 0x0
      13'hF9C: dout  = 8'b00000000; // 3996 :   0 - 0x0
      13'hF9D: dout  = 8'b00000000; // 3997 :   0 - 0x0
      13'hF9E: dout  = 8'b00000000; // 3998 :   0 - 0x0
      13'hF9F: dout  = 8'b00000000; // 3999 :   0 - 0x0
      13'hFA0: dout  = 8'b00000000; // 4000 :   0 - 0x0 -- Sprite 0xfa
      13'hFA1: dout  = 8'b00000000; // 4001 :   0 - 0x0
      13'hFA2: dout  = 8'b00000000; // 4002 :   0 - 0x0
      13'hFA3: dout  = 8'b00000000; // 4003 :   0 - 0x0
      13'hFA4: dout  = 8'b00000000; // 4004 :   0 - 0x0
      13'hFA5: dout  = 8'b00000000; // 4005 :   0 - 0x0
      13'hFA6: dout  = 8'b00000000; // 4006 :   0 - 0x0
      13'hFA7: dout  = 8'b00000000; // 4007 :   0 - 0x0
      13'hFA8: dout  = 8'b00000000; // 4008 :   0 - 0x0
      13'hFA9: dout  = 8'b00000000; // 4009 :   0 - 0x0
      13'hFAA: dout  = 8'b00000000; // 4010 :   0 - 0x0
      13'hFAB: dout  = 8'b00000000; // 4011 :   0 - 0x0
      13'hFAC: dout  = 8'b00000000; // 4012 :   0 - 0x0
      13'hFAD: dout  = 8'b00000000; // 4013 :   0 - 0x0
      13'hFAE: dout  = 8'b00000000; // 4014 :   0 - 0x0
      13'hFAF: dout  = 8'b00000000; // 4015 :   0 - 0x0
      13'hFB0: dout  = 8'b00000000; // 4016 :   0 - 0x0 -- Sprite 0xfb
      13'hFB1: dout  = 8'b00000000; // 4017 :   0 - 0x0
      13'hFB2: dout  = 8'b00000000; // 4018 :   0 - 0x0
      13'hFB3: dout  = 8'b00000000; // 4019 :   0 - 0x0
      13'hFB4: dout  = 8'b00000000; // 4020 :   0 - 0x0
      13'hFB5: dout  = 8'b00000000; // 4021 :   0 - 0x0
      13'hFB6: dout  = 8'b00000000; // 4022 :   0 - 0x0
      13'hFB7: dout  = 8'b00000000; // 4023 :   0 - 0x0
      13'hFB8: dout  = 8'b00000000; // 4024 :   0 - 0x0
      13'hFB9: dout  = 8'b00000000; // 4025 :   0 - 0x0
      13'hFBA: dout  = 8'b00000000; // 4026 :   0 - 0x0
      13'hFBB: dout  = 8'b00000000; // 4027 :   0 - 0x0
      13'hFBC: dout  = 8'b00000000; // 4028 :   0 - 0x0
      13'hFBD: dout  = 8'b00000000; // 4029 :   0 - 0x0
      13'hFBE: dout  = 8'b00000000; // 4030 :   0 - 0x0
      13'hFBF: dout  = 8'b00000000; // 4031 :   0 - 0x0
      13'hFC0: dout  = 8'b00000000; // 4032 :   0 - 0x0 -- Sprite 0xfc
      13'hFC1: dout  = 8'b00000000; // 4033 :   0 - 0x0
      13'hFC2: dout  = 8'b00000000; // 4034 :   0 - 0x0
      13'hFC3: dout  = 8'b00000000; // 4035 :   0 - 0x0
      13'hFC4: dout  = 8'b00000000; // 4036 :   0 - 0x0
      13'hFC5: dout  = 8'b00000000; // 4037 :   0 - 0x0
      13'hFC6: dout  = 8'b00000000; // 4038 :   0 - 0x0
      13'hFC7: dout  = 8'b00000000; // 4039 :   0 - 0x0
      13'hFC8: dout  = 8'b00000000; // 4040 :   0 - 0x0
      13'hFC9: dout  = 8'b00000000; // 4041 :   0 - 0x0
      13'hFCA: dout  = 8'b00000000; // 4042 :   0 - 0x0
      13'hFCB: dout  = 8'b00000000; // 4043 :   0 - 0x0
      13'hFCC: dout  = 8'b00000000; // 4044 :   0 - 0x0
      13'hFCD: dout  = 8'b00000000; // 4045 :   0 - 0x0
      13'hFCE: dout  = 8'b00000000; // 4046 :   0 - 0x0
      13'hFCF: dout  = 8'b00000000; // 4047 :   0 - 0x0
      13'hFD0: dout  = 8'b00000000; // 4048 :   0 - 0x0 -- Sprite 0xfd
      13'hFD1: dout  = 8'b00000000; // 4049 :   0 - 0x0
      13'hFD2: dout  = 8'b00000000; // 4050 :   0 - 0x0
      13'hFD3: dout  = 8'b00000000; // 4051 :   0 - 0x0
      13'hFD4: dout  = 8'b00000000; // 4052 :   0 - 0x0
      13'hFD5: dout  = 8'b00000000; // 4053 :   0 - 0x0
      13'hFD6: dout  = 8'b00000000; // 4054 :   0 - 0x0
      13'hFD7: dout  = 8'b00000000; // 4055 :   0 - 0x0
      13'hFD8: dout  = 8'b00000000; // 4056 :   0 - 0x0
      13'hFD9: dout  = 8'b00000000; // 4057 :   0 - 0x0
      13'hFDA: dout  = 8'b00000000; // 4058 :   0 - 0x0
      13'hFDB: dout  = 8'b00000000; // 4059 :   0 - 0x0
      13'hFDC: dout  = 8'b00000000; // 4060 :   0 - 0x0
      13'hFDD: dout  = 8'b00000000; // 4061 :   0 - 0x0
      13'hFDE: dout  = 8'b00000000; // 4062 :   0 - 0x0
      13'hFDF: dout  = 8'b00000000; // 4063 :   0 - 0x0
      13'hFE0: dout  = 8'b00000000; // 4064 :   0 - 0x0 -- Sprite 0xfe
      13'hFE1: dout  = 8'b00000000; // 4065 :   0 - 0x0
      13'hFE2: dout  = 8'b00000000; // 4066 :   0 - 0x0
      13'hFE3: dout  = 8'b00000000; // 4067 :   0 - 0x0
      13'hFE4: dout  = 8'b00000000; // 4068 :   0 - 0x0
      13'hFE5: dout  = 8'b00000000; // 4069 :   0 - 0x0
      13'hFE6: dout  = 8'b00000000; // 4070 :   0 - 0x0
      13'hFE7: dout  = 8'b00000000; // 4071 :   0 - 0x0
      13'hFE8: dout  = 8'b00000000; // 4072 :   0 - 0x0
      13'hFE9: dout  = 8'b00000000; // 4073 :   0 - 0x0
      13'hFEA: dout  = 8'b00000000; // 4074 :   0 - 0x0
      13'hFEB: dout  = 8'b00000000; // 4075 :   0 - 0x0
      13'hFEC: dout  = 8'b00000000; // 4076 :   0 - 0x0
      13'hFED: dout  = 8'b00000000; // 4077 :   0 - 0x0
      13'hFEE: dout  = 8'b00000000; // 4078 :   0 - 0x0
      13'hFEF: dout  = 8'b00000000; // 4079 :   0 - 0x0
      13'hFF0: dout  = 8'b00000000; // 4080 :   0 - 0x0 -- Sprite 0xff
      13'hFF1: dout  = 8'b00000000; // 4081 :   0 - 0x0
      13'hFF2: dout  = 8'b00000000; // 4082 :   0 - 0x0
      13'hFF3: dout  = 8'b00000000; // 4083 :   0 - 0x0
      13'hFF4: dout  = 8'b00000000; // 4084 :   0 - 0x0
      13'hFF5: dout  = 8'b00000000; // 4085 :   0 - 0x0
      13'hFF6: dout  = 8'b00000000; // 4086 :   0 - 0x0
      13'hFF7: dout  = 8'b00000000; // 4087 :   0 - 0x0
      13'hFF8: dout  = 8'b00000000; // 4088 :   0 - 0x0
      13'hFF9: dout  = 8'b00000000; // 4089 :   0 - 0x0
      13'hFFA: dout  = 8'b00000000; // 4090 :   0 - 0x0
      13'hFFB: dout  = 8'b00000000; // 4091 :   0 - 0x0
      13'hFFC: dout  = 8'b00000000; // 4092 :   0 - 0x0
      13'hFFD: dout  = 8'b00000000; // 4093 :   0 - 0x0
      13'hFFE: dout  = 8'b00000000; // 4094 :   0 - 0x0
      13'hFFF: dout  = 8'b00000000; // 4095 :   0 - 0x0
          // Pattern Table 1---------
      13'h1000: dout  = 8'b00111110; // 4096 :  62 - 0x3e -- Background 0x0
      13'h1001: dout  = 8'b01111111; // 4097 : 127 - 0x7f
      13'h1002: dout  = 8'b01110111; // 4098 : 119 - 0x77
      13'h1003: dout  = 8'b01111111; // 4099 : 127 - 0x7f
      13'h1004: dout  = 8'b01111111; // 4100 : 127 - 0x7f
      13'h1005: dout  = 8'b01110111; // 4101 : 119 - 0x77
      13'h1006: dout  = 8'b01111111; // 4102 : 127 - 0x7f
      13'h1007: dout  = 8'b00111110; // 4103 :  62 - 0x3e
      13'h1008: dout  = 8'b11000011; // 4104 : 195 - 0xc3
      13'h1009: dout  = 8'b10000001; // 4105 : 129 - 0x81
      13'h100A: dout  = 8'b10011001; // 4106 : 153 - 0x99
      13'h100B: dout  = 8'b10010001; // 4107 : 145 - 0x91
      13'h100C: dout  = 8'b10001001; // 4108 : 137 - 0x89
      13'h100D: dout  = 8'b10011001; // 4109 : 153 - 0x99
      13'h100E: dout  = 8'b10000001; // 4110 : 129 - 0x81
      13'h100F: dout  = 8'b11000011; // 4111 : 195 - 0xc3
      13'h1010: dout  = 8'b00011100; // 4112 :  28 - 0x1c -- Background 0x1
      13'h1011: dout  = 8'b00111100; // 4113 :  60 - 0x3c
      13'h1012: dout  = 8'b01111100; // 4114 : 124 - 0x7c
      13'h1013: dout  = 8'b00011100; // 4115 :  28 - 0x1c
      13'h1014: dout  = 8'b00011100; // 4116 :  28 - 0x1c
      13'h1015: dout  = 8'b00011100; // 4117 :  28 - 0x1c
      13'h1016: dout  = 8'b01111111; // 4118 : 127 - 0x7f
      13'h1017: dout  = 8'b01111111; // 4119 : 127 - 0x7f
      13'h1018: dout  = 8'b11100111; // 4120 : 231 - 0xe7
      13'h1019: dout  = 8'b11000111; // 4121 : 199 - 0xc7
      13'h101A: dout  = 8'b10000111; // 4122 : 135 - 0x87
      13'h101B: dout  = 8'b11100111; // 4123 : 231 - 0xe7
      13'h101C: dout  = 8'b11100111; // 4124 : 231 - 0xe7
      13'h101D: dout  = 8'b11100111; // 4125 : 231 - 0xe7
      13'h101E: dout  = 8'b10000001; // 4126 : 129 - 0x81
      13'h101F: dout  = 8'b10000001; // 4127 : 129 - 0x81
      13'h1020: dout  = 8'b00111110; // 4128 :  62 - 0x3e -- Background 0x2
      13'h1021: dout  = 8'b01111111; // 4129 : 127 - 0x7f
      13'h1022: dout  = 8'b00000111; // 4130 :   7 - 0x7
      13'h1023: dout  = 8'b00111111; // 4131 :  63 - 0x3f
      13'h1024: dout  = 8'b01111111; // 4132 : 127 - 0x7f
      13'h1025: dout  = 8'b01110000; // 4133 : 112 - 0x70
      13'h1026: dout  = 8'b01111111; // 4134 : 127 - 0x7f
      13'h1027: dout  = 8'b01111111; // 4135 : 127 - 0x7f
      13'h1028: dout  = 8'b11000011; // 4136 : 195 - 0xc3
      13'h1029: dout  = 8'b10000001; // 4137 : 129 - 0x81
      13'h102A: dout  = 8'b11111001; // 4138 : 249 - 0xf9
      13'h102B: dout  = 8'b11000001; // 4139 : 193 - 0xc1
      13'h102C: dout  = 8'b10000001; // 4140 : 129 - 0x81
      13'h102D: dout  = 8'b10011111; // 4141 : 159 - 0x9f
      13'h102E: dout  = 8'b10000001; // 4142 : 129 - 0x81
      13'h102F: dout  = 8'b10000001; // 4143 : 129 - 0x81
      13'h1030: dout  = 8'b00111110; // 4144 :  62 - 0x3e -- Background 0x3
      13'h1031: dout  = 8'b01111111; // 4145 : 127 - 0x7f
      13'h1032: dout  = 8'b00000111; // 4146 :   7 - 0x7
      13'h1033: dout  = 8'b00011111; // 4147 :  31 - 0x1f
      13'h1034: dout  = 8'b00011111; // 4148 :  31 - 0x1f
      13'h1035: dout  = 8'b00000111; // 4149 :   7 - 0x7
      13'h1036: dout  = 8'b01111111; // 4150 : 127 - 0x7f
      13'h1037: dout  = 8'b00111110; // 4151 :  62 - 0x3e
      13'h1038: dout  = 8'b11000011; // 4152 : 195 - 0xc3
      13'h1039: dout  = 8'b10000001; // 4153 : 129 - 0x81
      13'h103A: dout  = 8'b11111001; // 4154 : 249 - 0xf9
      13'h103B: dout  = 8'b11100001; // 4155 : 225 - 0xe1
      13'h103C: dout  = 8'b11100001; // 4156 : 225 - 0xe1
      13'h103D: dout  = 8'b11111001; // 4157 : 249 - 0xf9
      13'h103E: dout  = 8'b10000001; // 4158 : 129 - 0x81
      13'h103F: dout  = 8'b11000011; // 4159 : 195 - 0xc3
      13'h1040: dout  = 8'b00110000; // 4160 :  48 - 0x30 -- Background 0x4
      13'h1041: dout  = 8'b01110000; // 4161 : 112 - 0x70
      13'h1042: dout  = 8'b01110111; // 4162 : 119 - 0x77
      13'h1043: dout  = 8'b01110111; // 4163 : 119 - 0x77
      13'h1044: dout  = 8'b01111111; // 4164 : 127 - 0x7f
      13'h1045: dout  = 8'b01111111; // 4165 : 127 - 0x7f
      13'h1046: dout  = 8'b00000111; // 4166 :   7 - 0x7
      13'h1047: dout  = 8'b00000111; // 4167 :   7 - 0x7
      13'h1048: dout  = 8'b11011111; // 4168 : 223 - 0xdf
      13'h1049: dout  = 8'b10011111; // 4169 : 159 - 0x9f
      13'h104A: dout  = 8'b10011001; // 4170 : 153 - 0x99
      13'h104B: dout  = 8'b10011001; // 4171 : 153 - 0x99
      13'h104C: dout  = 8'b10000000; // 4172 : 128 - 0x80
      13'h104D: dout  = 8'b10000000; // 4173 : 128 - 0x80
      13'h104E: dout  = 8'b11111001; // 4174 : 249 - 0xf9
      13'h104F: dout  = 8'b11111001; // 4175 : 249 - 0xf9
      13'h1050: dout  = 8'b01111111; // 4176 : 127 - 0x7f -- Background 0x5
      13'h1051: dout  = 8'b01111111; // 4177 : 127 - 0x7f
      13'h1052: dout  = 8'b01110000; // 4178 : 112 - 0x70
      13'h1053: dout  = 8'b01111110; // 4179 : 126 - 0x7e
      13'h1054: dout  = 8'b01111111; // 4180 : 127 - 0x7f
      13'h1055: dout  = 8'b00000111; // 4181 :   7 - 0x7
      13'h1056: dout  = 8'b01111111; // 4182 : 127 - 0x7f
      13'h1057: dout  = 8'b00111110; // 4183 :  62 - 0x3e
      13'h1058: dout  = 8'b10000001; // 4184 : 129 - 0x81
      13'h1059: dout  = 8'b10000001; // 4185 : 129 - 0x81
      13'h105A: dout  = 8'b10011111; // 4186 : 159 - 0x9f
      13'h105B: dout  = 8'b10000011; // 4187 : 131 - 0x83
      13'h105C: dout  = 8'b10000001; // 4188 : 129 - 0x81
      13'h105D: dout  = 8'b11111001; // 4189 : 249 - 0xf9
      13'h105E: dout  = 8'b10000001; // 4190 : 129 - 0x81
      13'h105F: dout  = 8'b11000011; // 4191 : 195 - 0xc3
      13'h1060: dout  = 8'b00111110; // 4192 :  62 - 0x3e -- Background 0x6
      13'h1061: dout  = 8'b01111111; // 4193 : 127 - 0x7f
      13'h1062: dout  = 8'b01110000; // 4194 : 112 - 0x70
      13'h1063: dout  = 8'b01111110; // 4195 : 126 - 0x7e
      13'h1064: dout  = 8'b01111111; // 4196 : 127 - 0x7f
      13'h1065: dout  = 8'b01110111; // 4197 : 119 - 0x77
      13'h1066: dout  = 8'b01111111; // 4198 : 127 - 0x7f
      13'h1067: dout  = 8'b00111110; // 4199 :  62 - 0x3e
      13'h1068: dout  = 8'b11000011; // 4200 : 195 - 0xc3
      13'h1069: dout  = 8'b10000001; // 4201 : 129 - 0x81
      13'h106A: dout  = 8'b10011111; // 4202 : 159 - 0x9f
      13'h106B: dout  = 8'b10000011; // 4203 : 131 - 0x83
      13'h106C: dout  = 8'b10000001; // 4204 : 129 - 0x81
      13'h106D: dout  = 8'b10011001; // 4205 : 153 - 0x99
      13'h106E: dout  = 8'b10000001; // 4206 : 129 - 0x81
      13'h106F: dout  = 8'b11000011; // 4207 : 195 - 0xc3
      13'h1070: dout  = 8'b01111111; // 4208 : 127 - 0x7f -- Background 0x7
      13'h1071: dout  = 8'b01111111; // 4209 : 127 - 0x7f
      13'h1072: dout  = 8'b00000111; // 4210 :   7 - 0x7
      13'h1073: dout  = 8'b00001110; // 4211 :  14 - 0xe
      13'h1074: dout  = 8'b00001110; // 4212 :  14 - 0xe
      13'h1075: dout  = 8'b00011100; // 4213 :  28 - 0x1c
      13'h1076: dout  = 8'b00011100; // 4214 :  28 - 0x1c
      13'h1077: dout  = 8'b00011100; // 4215 :  28 - 0x1c
      13'h1078: dout  = 8'b10000001; // 4216 : 129 - 0x81
      13'h1079: dout  = 8'b10000001; // 4217 : 129 - 0x81
      13'h107A: dout  = 8'b11111001; // 4218 : 249 - 0xf9
      13'h107B: dout  = 8'b11110011; // 4219 : 243 - 0xf3
      13'h107C: dout  = 8'b11110011; // 4220 : 243 - 0xf3
      13'h107D: dout  = 8'b11100111; // 4221 : 231 - 0xe7
      13'h107E: dout  = 8'b11100111; // 4222 : 231 - 0xe7
      13'h107F: dout  = 8'b11100111; // 4223 : 231 - 0xe7
      13'h1080: dout  = 8'b00111110; // 4224 :  62 - 0x3e -- Background 0x8
      13'h1081: dout  = 8'b01111111; // 4225 : 127 - 0x7f
      13'h1082: dout  = 8'b01110111; // 4226 : 119 - 0x77
      13'h1083: dout  = 8'b00111110; // 4227 :  62 - 0x3e
      13'h1084: dout  = 8'b01111111; // 4228 : 127 - 0x7f
      13'h1085: dout  = 8'b01110111; // 4229 : 119 - 0x77
      13'h1086: dout  = 8'b01111111; // 4230 : 127 - 0x7f
      13'h1087: dout  = 8'b00111110; // 4231 :  62 - 0x3e
      13'h1088: dout  = 8'b11000011; // 4232 : 195 - 0xc3
      13'h1089: dout  = 8'b10000001; // 4233 : 129 - 0x81
      13'h108A: dout  = 8'b10011001; // 4234 : 153 - 0x99
      13'h108B: dout  = 8'b11000011; // 4235 : 195 - 0xc3
      13'h108C: dout  = 8'b10000001; // 4236 : 129 - 0x81
      13'h108D: dout  = 8'b10011001; // 4237 : 153 - 0x99
      13'h108E: dout  = 8'b10000001; // 4238 : 129 - 0x81
      13'h108F: dout  = 8'b11000011; // 4239 : 195 - 0xc3
      13'h1090: dout  = 8'b00111110; // 4240 :  62 - 0x3e -- Background 0x9
      13'h1091: dout  = 8'b01111111; // 4241 : 127 - 0x7f
      13'h1092: dout  = 8'b01110111; // 4242 : 119 - 0x77
      13'h1093: dout  = 8'b01111111; // 4243 : 127 - 0x7f
      13'h1094: dout  = 8'b00111111; // 4244 :  63 - 0x3f
      13'h1095: dout  = 8'b00000111; // 4245 :   7 - 0x7
      13'h1096: dout  = 8'b01111111; // 4246 : 127 - 0x7f
      13'h1097: dout  = 8'b00111110; // 4247 :  62 - 0x3e
      13'h1098: dout  = 8'b11000011; // 4248 : 195 - 0xc3
      13'h1099: dout  = 8'b10000001; // 4249 : 129 - 0x81
      13'h109A: dout  = 8'b10011001; // 4250 : 153 - 0x99
      13'h109B: dout  = 8'b10000001; // 4251 : 129 - 0x81
      13'h109C: dout  = 8'b11000001; // 4252 : 193 - 0xc1
      13'h109D: dout  = 8'b11111001; // 4253 : 249 - 0xf9
      13'h109E: dout  = 8'b10000001; // 4254 : 129 - 0x81
      13'h109F: dout  = 8'b11000011; // 4255 : 195 - 0xc3
      13'h10A0: dout  = 8'b00000000; // 4256 :   0 - 0x0 -- Background 0xa
      13'h10A1: dout  = 8'b00000000; // 4257 :   0 - 0x0
      13'h10A2: dout  = 8'b00000000; // 4258 :   0 - 0x0
      13'h10A3: dout  = 8'b00000000; // 4259 :   0 - 0x0
      13'h10A4: dout  = 8'b00000000; // 4260 :   0 - 0x0
      13'h10A5: dout  = 8'b00110000; // 4261 :  48 - 0x30
      13'h10A6: dout  = 8'b01111000; // 4262 : 120 - 0x78
      13'h10A7: dout  = 8'b00110000; // 4263 :  48 - 0x30
      13'h10A8: dout  = 8'b11111111; // 4264 : 255 - 0xff
      13'h10A9: dout  = 8'b11111111; // 4265 : 255 - 0xff
      13'h10AA: dout  = 8'b11111111; // 4266 : 255 - 0xff
      13'h10AB: dout  = 8'b11111111; // 4267 : 255 - 0xff
      13'h10AC: dout  = 8'b11111111; // 4268 : 255 - 0xff
      13'h10AD: dout  = 8'b11011111; // 4269 : 223 - 0xdf
      13'h10AE: dout  = 8'b10001111; // 4270 : 143 - 0x8f
      13'h10AF: dout  = 8'b11011111; // 4271 : 223 - 0xdf
      13'h10B0: dout  = 8'b01110000; // 4272 : 112 - 0x70 -- Background 0xb
      13'h10B1: dout  = 8'b11111000; // 4273 : 248 - 0xf8
      13'h10B2: dout  = 8'b11111000; // 4274 : 248 - 0xf8
      13'h10B3: dout  = 8'b11111000; // 4275 : 248 - 0xf8
      13'h10B4: dout  = 8'b01110000; // 4276 : 112 - 0x70
      13'h10B5: dout  = 8'b00000000; // 4277 :   0 - 0x0
      13'h10B6: dout  = 8'b01110000; // 4278 : 112 - 0x70
      13'h10B7: dout  = 8'b01110000; // 4279 : 112 - 0x70
      13'h10B8: dout  = 8'b10011111; // 4280 : 159 - 0x9f
      13'h10B9: dout  = 8'b00001111; // 4281 :  15 - 0xf
      13'h10BA: dout  = 8'b00001111; // 4282 :  15 - 0xf
      13'h10BB: dout  = 8'b00001111; // 4283 :  15 - 0xf
      13'h10BC: dout  = 8'b10011111; // 4284 : 159 - 0x9f
      13'h10BD: dout  = 8'b11111111; // 4285 : 255 - 0xff
      13'h10BE: dout  = 8'b10011111; // 4286 : 159 - 0x9f
      13'h10BF: dout  = 8'b10011111; // 4287 : 159 - 0x9f
      13'h10C0: dout  = 8'b01111000; // 4288 : 120 - 0x78 -- Background 0xc
      13'h10C1: dout  = 8'b11111100; // 4289 : 252 - 0xfc
      13'h10C2: dout  = 8'b00011100; // 4290 :  28 - 0x1c
      13'h10C3: dout  = 8'b00111000; // 4291 :  56 - 0x38
      13'h10C4: dout  = 8'b00110000; // 4292 :  48 - 0x30
      13'h10C5: dout  = 8'b00000000; // 4293 :   0 - 0x0
      13'h10C6: dout  = 8'b01110000; // 4294 : 112 - 0x70
      13'h10C7: dout  = 8'b01110000; // 4295 : 112 - 0x70
      13'h10C8: dout  = 8'b10001111; // 4296 : 143 - 0x8f
      13'h10C9: dout  = 8'b00100111; // 4297 :  39 - 0x27
      13'h10CA: dout  = 8'b11100111; // 4298 : 231 - 0xe7
      13'h10CB: dout  = 8'b11001111; // 4299 : 207 - 0xcf
      13'h10CC: dout  = 8'b11011111; // 4300 : 223 - 0xdf
      13'h10CD: dout  = 8'b11111111; // 4301 : 255 - 0xff
      13'h10CE: dout  = 8'b10011111; // 4302 : 159 - 0x9f
      13'h10CF: dout  = 8'b10011111; // 4303 : 159 - 0x9f
      13'h10D0: dout  = 8'b00111100; // 4304 :  60 - 0x3c -- Background 0xd
      13'h10D1: dout  = 8'b01111110; // 4305 : 126 - 0x7e
      13'h10D2: dout  = 8'b11011011; // 4306 : 219 - 0xdb
      13'h10D3: dout  = 8'b11011111; // 4307 : 223 - 0xdf
      13'h10D4: dout  = 8'b11000011; // 4308 : 195 - 0xc3
      13'h10D5: dout  = 8'b01100110; // 4309 : 102 - 0x66
      13'h10D6: dout  = 8'b00111100; // 4310 :  60 - 0x3c
      13'h10D7: dout  = 8'b00000000; // 4311 :   0 - 0x0
      13'h10D8: dout  = 8'b11000111; // 4312 : 199 - 0xc7
      13'h10D9: dout  = 8'b10101011; // 4313 : 171 - 0xab
      13'h10DA: dout  = 8'b01101101; // 4314 : 109 - 0x6d
      13'h10DB: dout  = 8'b01100101; // 4315 : 101 - 0x65
      13'h10DC: dout  = 8'b01111101; // 4316 : 125 - 0x7d
      13'h10DD: dout  = 8'b10111011; // 4317 : 187 - 0xbb
      13'h10DE: dout  = 8'b11000111; // 4318 : 199 - 0xc7
      13'h10DF: dout  = 8'b11111111; // 4319 : 255 - 0xff
      13'h10E0: dout  = 8'b00000000; // 4320 :   0 - 0x0 -- Background 0xe
      13'h10E1: dout  = 8'b00000000; // 4321 :   0 - 0x0
      13'h10E2: dout  = 8'b00000000; // 4322 :   0 - 0x0
      13'h10E3: dout  = 8'b00111100; // 4323 :  60 - 0x3c
      13'h10E4: dout  = 8'b00111110; // 4324 :  62 - 0x3e
      13'h10E5: dout  = 8'b00011110; // 4325 :  30 - 0x1e
      13'h10E6: dout  = 8'b00000000; // 4326 :   0 - 0x0
      13'h10E7: dout  = 8'b00000000; // 4327 :   0 - 0x0
      13'h10E8: dout  = 8'b11111111; // 4328 : 255 - 0xff
      13'h10E9: dout  = 8'b11111111; // 4329 : 255 - 0xff
      13'h10EA: dout  = 8'b11111111; // 4330 : 255 - 0xff
      13'h10EB: dout  = 8'b11000011; // 4331 : 195 - 0xc3
      13'h10EC: dout  = 8'b11000011; // 4332 : 195 - 0xc3
      13'h10ED: dout  = 8'b11111111; // 4333 : 255 - 0xff
      13'h10EE: dout  = 8'b11111111; // 4334 : 255 - 0xff
      13'h10EF: dout  = 8'b11111111; // 4335 : 255 - 0xff
      13'h10F0: dout  = 8'b11111111; // 4336 : 255 - 0xff -- Background 0xf
      13'h10F1: dout  = 8'b11111111; // 4337 : 255 - 0xff
      13'h10F2: dout  = 8'b11111111; // 4338 : 255 - 0xff
      13'h10F3: dout  = 8'b11111111; // 4339 : 255 - 0xff
      13'h10F4: dout  = 8'b11111111; // 4340 : 255 - 0xff
      13'h10F5: dout  = 8'b11111111; // 4341 : 255 - 0xff
      13'h10F6: dout  = 8'b11100000; // 4342 : 224 - 0xe0
      13'h10F7: dout  = 8'b11100000; // 4343 : 224 - 0xe0
      13'h10F8: dout  = 8'b00000001; // 4344 :   1 - 0x1
      13'h10F9: dout  = 8'b00101001; // 4345 :  41 - 0x29
      13'h10FA: dout  = 8'b01010101; // 4346 :  85 - 0x55
      13'h10FB: dout  = 8'b00101001; // 4347 :  41 - 0x29
      13'h10FC: dout  = 8'b01010101; // 4348 :  85 - 0x55
      13'h10FD: dout  = 8'b00000001; // 4349 :   1 - 0x1
      13'h10FE: dout  = 8'b00111111; // 4350 :  63 - 0x3f
      13'h10FF: dout  = 8'b00111111; // 4351 :  63 - 0x3f
      13'h1100: dout  = 8'b00001110; // 4352 :  14 - 0xe -- Background 0x10
      13'h1101: dout  = 8'b00001110; // 4353 :  14 - 0xe
      13'h1102: dout  = 8'b00011100; // 4354 :  28 - 0x1c
      13'h1103: dout  = 8'b00011100; // 4355 :  28 - 0x1c
      13'h1104: dout  = 8'b00011100; // 4356 :  28 - 0x1c
      13'h1105: dout  = 8'b00011100; // 4357 :  28 - 0x1c
      13'h1106: dout  = 8'b00111000; // 4358 :  56 - 0x38
      13'h1107: dout  = 8'b00111000; // 4359 :  56 - 0x38
      13'h1108: dout  = 8'b11110011; // 4360 : 243 - 0xf3
      13'h1109: dout  = 8'b11110011; // 4361 : 243 - 0xf3
      13'h110A: dout  = 8'b11100111; // 4362 : 231 - 0xe7
      13'h110B: dout  = 8'b11100111; // 4363 : 231 - 0xe7
      13'h110C: dout  = 8'b11100111; // 4364 : 231 - 0xe7
      13'h110D: dout  = 8'b11100111; // 4365 : 231 - 0xe7
      13'h110E: dout  = 8'b11001111; // 4366 : 207 - 0xcf
      13'h110F: dout  = 8'b11001111; // 4367 : 207 - 0xcf
      13'h1110: dout  = 8'b00011100; // 4368 :  28 - 0x1c -- Background 0x11
      13'h1111: dout  = 8'b00111110; // 4369 :  62 - 0x3e
      13'h1112: dout  = 8'b01110111; // 4370 : 119 - 0x77
      13'h1113: dout  = 8'b01110111; // 4371 : 119 - 0x77
      13'h1114: dout  = 8'b01111111; // 4372 : 127 - 0x7f
      13'h1115: dout  = 8'b01111111; // 4373 : 127 - 0x7f
      13'h1116: dout  = 8'b01110111; // 4374 : 119 - 0x77
      13'h1117: dout  = 8'b01110111; // 4375 : 119 - 0x77
      13'h1118: dout  = 8'b11100111; // 4376 : 231 - 0xe7
      13'h1119: dout  = 8'b11000011; // 4377 : 195 - 0xc3
      13'h111A: dout  = 8'b10011001; // 4378 : 153 - 0x99
      13'h111B: dout  = 8'b10011001; // 4379 : 153 - 0x99
      13'h111C: dout  = 8'b10000001; // 4380 : 129 - 0x81
      13'h111D: dout  = 8'b10000001; // 4381 : 129 - 0x81
      13'h111E: dout  = 8'b10011001; // 4382 : 153 - 0x99
      13'h111F: dout  = 8'b10011001; // 4383 : 153 - 0x99
      13'h1120: dout  = 8'b01111110; // 4384 : 126 - 0x7e -- Background 0x12
      13'h1121: dout  = 8'b01110111; // 4385 : 119 - 0x77
      13'h1122: dout  = 8'b01110111; // 4386 : 119 - 0x77
      13'h1123: dout  = 8'b01111110; // 4387 : 126 - 0x7e
      13'h1124: dout  = 8'b01111110; // 4388 : 126 - 0x7e
      13'h1125: dout  = 8'b01110111; // 4389 : 119 - 0x77
      13'h1126: dout  = 8'b01110111; // 4390 : 119 - 0x77
      13'h1127: dout  = 8'b01111110; // 4391 : 126 - 0x7e
      13'h1128: dout  = 8'b10000011; // 4392 : 131 - 0x83
      13'h1129: dout  = 8'b10011001; // 4393 : 153 - 0x99
      13'h112A: dout  = 8'b10011001; // 4394 : 153 - 0x99
      13'h112B: dout  = 8'b10000011; // 4395 : 131 - 0x83
      13'h112C: dout  = 8'b10000011; // 4396 : 131 - 0x83
      13'h112D: dout  = 8'b10011001; // 4397 : 153 - 0x99
      13'h112E: dout  = 8'b10011001; // 4398 : 153 - 0x99
      13'h112F: dout  = 8'b10000011; // 4399 : 131 - 0x83
      13'h1130: dout  = 8'b00111110; // 4400 :  62 - 0x3e -- Background 0x13
      13'h1131: dout  = 8'b01111111; // 4401 : 127 - 0x7f
      13'h1132: dout  = 8'b01110111; // 4402 : 119 - 0x77
      13'h1133: dout  = 8'b01110000; // 4403 : 112 - 0x70
      13'h1134: dout  = 8'b01110000; // 4404 : 112 - 0x70
      13'h1135: dout  = 8'b01110111; // 4405 : 119 - 0x77
      13'h1136: dout  = 8'b01111111; // 4406 : 127 - 0x7f
      13'h1137: dout  = 8'b00111110; // 4407 :  62 - 0x3e
      13'h1138: dout  = 8'b11000011; // 4408 : 195 - 0xc3
      13'h1139: dout  = 8'b10000001; // 4409 : 129 - 0x81
      13'h113A: dout  = 8'b10011001; // 4410 : 153 - 0x99
      13'h113B: dout  = 8'b10011111; // 4411 : 159 - 0x9f
      13'h113C: dout  = 8'b10011111; // 4412 : 159 - 0x9f
      13'h113D: dout  = 8'b10011001; // 4413 : 153 - 0x99
      13'h113E: dout  = 8'b10000001; // 4414 : 129 - 0x81
      13'h113F: dout  = 8'b11000011; // 4415 : 195 - 0xc3
      13'h1140: dout  = 8'b01111110; // 4416 : 126 - 0x7e -- Background 0x14
      13'h1141: dout  = 8'b01111111; // 4417 : 127 - 0x7f
      13'h1142: dout  = 8'b01110111; // 4418 : 119 - 0x77
      13'h1143: dout  = 8'b01110111; // 4419 : 119 - 0x77
      13'h1144: dout  = 8'b01110111; // 4420 : 119 - 0x77
      13'h1145: dout  = 8'b01110111; // 4421 : 119 - 0x77
      13'h1146: dout  = 8'b01111111; // 4422 : 127 - 0x7f
      13'h1147: dout  = 8'b01111110; // 4423 : 126 - 0x7e
      13'h1148: dout  = 8'b10000011; // 4424 : 131 - 0x83
      13'h1149: dout  = 8'b10000001; // 4425 : 129 - 0x81
      13'h114A: dout  = 8'b10011001; // 4426 : 153 - 0x99
      13'h114B: dout  = 8'b10011001; // 4427 : 153 - 0x99
      13'h114C: dout  = 8'b10011001; // 4428 : 153 - 0x99
      13'h114D: dout  = 8'b10011001; // 4429 : 153 - 0x99
      13'h114E: dout  = 8'b10000001; // 4430 : 129 - 0x81
      13'h114F: dout  = 8'b10000011; // 4431 : 131 - 0x83
      13'h1150: dout  = 8'b01111111; // 4432 : 127 - 0x7f -- Background 0x15
      13'h1151: dout  = 8'b01111111; // 4433 : 127 - 0x7f
      13'h1152: dout  = 8'b01110000; // 4434 : 112 - 0x70
      13'h1153: dout  = 8'b01111100; // 4435 : 124 - 0x7c
      13'h1154: dout  = 8'b01111100; // 4436 : 124 - 0x7c
      13'h1155: dout  = 8'b01110000; // 4437 : 112 - 0x70
      13'h1156: dout  = 8'b01111111; // 4438 : 127 - 0x7f
      13'h1157: dout  = 8'b01111111; // 4439 : 127 - 0x7f
      13'h1158: dout  = 8'b10000001; // 4440 : 129 - 0x81
      13'h1159: dout  = 8'b10000001; // 4441 : 129 - 0x81
      13'h115A: dout  = 8'b10011111; // 4442 : 159 - 0x9f
      13'h115B: dout  = 8'b10000111; // 4443 : 135 - 0x87
      13'h115C: dout  = 8'b10000111; // 4444 : 135 - 0x87
      13'h115D: dout  = 8'b10011111; // 4445 : 159 - 0x9f
      13'h115E: dout  = 8'b10000001; // 4446 : 129 - 0x81
      13'h115F: dout  = 8'b10000001; // 4447 : 129 - 0x81
      13'h1160: dout  = 8'b01111111; // 4448 : 127 - 0x7f -- Background 0x16
      13'h1161: dout  = 8'b01111111; // 4449 : 127 - 0x7f
      13'h1162: dout  = 8'b01110000; // 4450 : 112 - 0x70
      13'h1163: dout  = 8'b01111100; // 4451 : 124 - 0x7c
      13'h1164: dout  = 8'b01111100; // 4452 : 124 - 0x7c
      13'h1165: dout  = 8'b01110000; // 4453 : 112 - 0x70
      13'h1166: dout  = 8'b01110000; // 4454 : 112 - 0x70
      13'h1167: dout  = 8'b01110000; // 4455 : 112 - 0x70
      13'h1168: dout  = 8'b10000001; // 4456 : 129 - 0x81
      13'h1169: dout  = 8'b10000001; // 4457 : 129 - 0x81
      13'h116A: dout  = 8'b10011111; // 4458 : 159 - 0x9f
      13'h116B: dout  = 8'b10000111; // 4459 : 135 - 0x87
      13'h116C: dout  = 8'b10000111; // 4460 : 135 - 0x87
      13'h116D: dout  = 8'b10011111; // 4461 : 159 - 0x9f
      13'h116E: dout  = 8'b10011111; // 4462 : 159 - 0x9f
      13'h116F: dout  = 8'b10011111; // 4463 : 159 - 0x9f
      13'h1170: dout  = 8'b00111110; // 4464 :  62 - 0x3e -- Background 0x17
      13'h1171: dout  = 8'b01111111; // 4465 : 127 - 0x7f
      13'h1172: dout  = 8'b01110111; // 4466 : 119 - 0x77
      13'h1173: dout  = 8'b01110000; // 4467 : 112 - 0x70
      13'h1174: dout  = 8'b01111111; // 4468 : 127 - 0x7f
      13'h1175: dout  = 8'b01110111; // 4469 : 119 - 0x77
      13'h1176: dout  = 8'b01111111; // 4470 : 127 - 0x7f
      13'h1177: dout  = 8'b00111110; // 4471 :  62 - 0x3e
      13'h1178: dout  = 8'b11000011; // 4472 : 195 - 0xc3
      13'h1179: dout  = 8'b10000001; // 4473 : 129 - 0x81
      13'h117A: dout  = 8'b10011001; // 4474 : 153 - 0x99
      13'h117B: dout  = 8'b10011111; // 4475 : 159 - 0x9f
      13'h117C: dout  = 8'b10010001; // 4476 : 145 - 0x91
      13'h117D: dout  = 8'b10011001; // 4477 : 153 - 0x99
      13'h117E: dout  = 8'b10000001; // 4478 : 129 - 0x81
      13'h117F: dout  = 8'b11000011; // 4479 : 195 - 0xc3
      13'h1180: dout  = 8'b01110111; // 4480 : 119 - 0x77 -- Background 0x18
      13'h1181: dout  = 8'b01110111; // 4481 : 119 - 0x77
      13'h1182: dout  = 8'b01110111; // 4482 : 119 - 0x77
      13'h1183: dout  = 8'b01111111; // 4483 : 127 - 0x7f
      13'h1184: dout  = 8'b01111111; // 4484 : 127 - 0x7f
      13'h1185: dout  = 8'b01110111; // 4485 : 119 - 0x77
      13'h1186: dout  = 8'b01110111; // 4486 : 119 - 0x77
      13'h1187: dout  = 8'b01110111; // 4487 : 119 - 0x77
      13'h1188: dout  = 8'b10011001; // 4488 : 153 - 0x99
      13'h1189: dout  = 8'b10011001; // 4489 : 153 - 0x99
      13'h118A: dout  = 8'b10011001; // 4490 : 153 - 0x99
      13'h118B: dout  = 8'b10000001; // 4491 : 129 - 0x81
      13'h118C: dout  = 8'b10000001; // 4492 : 129 - 0x81
      13'h118D: dout  = 8'b10011001; // 4493 : 153 - 0x99
      13'h118E: dout  = 8'b10011001; // 4494 : 153 - 0x99
      13'h118F: dout  = 8'b10011001; // 4495 : 153 - 0x99
      13'h1190: dout  = 8'b00111110; // 4496 :  62 - 0x3e -- Background 0x19
      13'h1191: dout  = 8'b00111110; // 4497 :  62 - 0x3e
      13'h1192: dout  = 8'b00011100; // 4498 :  28 - 0x1c
      13'h1193: dout  = 8'b00011100; // 4499 :  28 - 0x1c
      13'h1194: dout  = 8'b00011100; // 4500 :  28 - 0x1c
      13'h1195: dout  = 8'b00011100; // 4501 :  28 - 0x1c
      13'h1196: dout  = 8'b00111110; // 4502 :  62 - 0x3e
      13'h1197: dout  = 8'b00111110; // 4503 :  62 - 0x3e
      13'h1198: dout  = 8'b11000011; // 4504 : 195 - 0xc3
      13'h1199: dout  = 8'b11000011; // 4505 : 195 - 0xc3
      13'h119A: dout  = 8'b11100111; // 4506 : 231 - 0xe7
      13'h119B: dout  = 8'b11100111; // 4507 : 231 - 0xe7
      13'h119C: dout  = 8'b11100111; // 4508 : 231 - 0xe7
      13'h119D: dout  = 8'b11100111; // 4509 : 231 - 0xe7
      13'h119E: dout  = 8'b11000011; // 4510 : 195 - 0xc3
      13'h119F: dout  = 8'b11000011; // 4511 : 195 - 0xc3
      13'h11A0: dout  = 8'b00000111; // 4512 :   7 - 0x7 -- Background 0x1a
      13'h11A1: dout  = 8'b00000111; // 4513 :   7 - 0x7
      13'h11A2: dout  = 8'b00000111; // 4514 :   7 - 0x7
      13'h11A3: dout  = 8'b00000111; // 4515 :   7 - 0x7
      13'h11A4: dout  = 8'b00000111; // 4516 :   7 - 0x7
      13'h11A5: dout  = 8'b01110111; // 4517 : 119 - 0x77
      13'h11A6: dout  = 8'b01111111; // 4518 : 127 - 0x7f
      13'h11A7: dout  = 8'b00111110; // 4519 :  62 - 0x3e
      13'h11A8: dout  = 8'b11111001; // 4520 : 249 - 0xf9
      13'h11A9: dout  = 8'b11111001; // 4521 : 249 - 0xf9
      13'h11AA: dout  = 8'b11111001; // 4522 : 249 - 0xf9
      13'h11AB: dout  = 8'b11111001; // 4523 : 249 - 0xf9
      13'h11AC: dout  = 8'b11111001; // 4524 : 249 - 0xf9
      13'h11AD: dout  = 8'b10011001; // 4525 : 153 - 0x99
      13'h11AE: dout  = 8'b10000001; // 4526 : 129 - 0x81
      13'h11AF: dout  = 8'b11000011; // 4527 : 195 - 0xc3
      13'h11B0: dout  = 8'b01110011; // 4528 : 115 - 0x73 -- Background 0x1b
      13'h11B1: dout  = 8'b01110111; // 4529 : 119 - 0x77
      13'h11B2: dout  = 8'b01111110; // 4530 : 126 - 0x7e
      13'h11B3: dout  = 8'b01111100; // 4531 : 124 - 0x7c
      13'h11B4: dout  = 8'b01111110; // 4532 : 126 - 0x7e
      13'h11B5: dout  = 8'b01110111; // 4533 : 119 - 0x77
      13'h11B6: dout  = 8'b01110111; // 4534 : 119 - 0x77
      13'h11B7: dout  = 8'b01110111; // 4535 : 119 - 0x77
      13'h11B8: dout  = 8'b10011101; // 4536 : 157 - 0x9d
      13'h11B9: dout  = 8'b10011001; // 4537 : 153 - 0x99
      13'h11BA: dout  = 8'b10010011; // 4538 : 147 - 0x93
      13'h11BB: dout  = 8'b10000111; // 4539 : 135 - 0x87
      13'h11BC: dout  = 8'b10000011; // 4540 : 131 - 0x83
      13'h11BD: dout  = 8'b10011001; // 4541 : 153 - 0x99
      13'h11BE: dout  = 8'b10011001; // 4542 : 153 - 0x99
      13'h11BF: dout  = 8'b10011001; // 4543 : 153 - 0x99
      13'h11C0: dout  = 8'b01110000; // 4544 : 112 - 0x70 -- Background 0x1c
      13'h11C1: dout  = 8'b01110000; // 4545 : 112 - 0x70
      13'h11C2: dout  = 8'b01110000; // 4546 : 112 - 0x70
      13'h11C3: dout  = 8'b01110000; // 4547 : 112 - 0x70
      13'h11C4: dout  = 8'b01110000; // 4548 : 112 - 0x70
      13'h11C5: dout  = 8'b01110000; // 4549 : 112 - 0x70
      13'h11C6: dout  = 8'b01111111; // 4550 : 127 - 0x7f
      13'h11C7: dout  = 8'b01111111; // 4551 : 127 - 0x7f
      13'h11C8: dout  = 8'b10011111; // 4552 : 159 - 0x9f
      13'h11C9: dout  = 8'b10011111; // 4553 : 159 - 0x9f
      13'h11CA: dout  = 8'b10011111; // 4554 : 159 - 0x9f
      13'h11CB: dout  = 8'b10011111; // 4555 : 159 - 0x9f
      13'h11CC: dout  = 8'b10011111; // 4556 : 159 - 0x9f
      13'h11CD: dout  = 8'b10011111; // 4557 : 159 - 0x9f
      13'h11CE: dout  = 8'b10000001; // 4558 : 129 - 0x81
      13'h11CF: dout  = 8'b10000001; // 4559 : 129 - 0x81
      13'h11D0: dout  = 8'b11100111; // 4560 : 231 - 0xe7 -- Background 0x1d
      13'h11D1: dout  = 8'b11111111; // 4561 : 255 - 0xff
      13'h11D2: dout  = 8'b11111111; // 4562 : 255 - 0xff
      13'h11D3: dout  = 8'b11111111; // 4563 : 255 - 0xff
      13'h11D4: dout  = 8'b11111111; // 4564 : 255 - 0xff
      13'h11D5: dout  = 8'b11100111; // 4565 : 231 - 0xe7
      13'h11D6: dout  = 8'b11100111; // 4566 : 231 - 0xe7
      13'h11D7: dout  = 8'b11100111; // 4567 : 231 - 0xe7
      13'h11D8: dout  = 8'b00111001; // 4568 :  57 - 0x39
      13'h11D9: dout  = 8'b00010001; // 4569 :  17 - 0x11
      13'h11DA: dout  = 8'b00000001; // 4570 :   1 - 0x1
      13'h11DB: dout  = 8'b00000001; // 4571 :   1 - 0x1
      13'h11DC: dout  = 8'b00101001; // 4572 :  41 - 0x29
      13'h11DD: dout  = 8'b00111001; // 4573 :  57 - 0x39
      13'h11DE: dout  = 8'b00111001; // 4574 :  57 - 0x39
      13'h11DF: dout  = 8'b00111001; // 4575 :  57 - 0x39
      13'h11E0: dout  = 8'b01110111; // 4576 : 119 - 0x77 -- Background 0x1e
      13'h11E1: dout  = 8'b01110111; // 4577 : 119 - 0x77
      13'h11E2: dout  = 8'b01111111; // 4578 : 127 - 0x7f
      13'h11E3: dout  = 8'b01111111; // 4579 : 127 - 0x7f
      13'h11E4: dout  = 8'b01111111; // 4580 : 127 - 0x7f
      13'h11E5: dout  = 8'b01111111; // 4581 : 127 - 0x7f
      13'h11E6: dout  = 8'b01110111; // 4582 : 119 - 0x77
      13'h11E7: dout  = 8'b01110111; // 4583 : 119 - 0x77
      13'h11E8: dout  = 8'b10011001; // 4584 : 153 - 0x99
      13'h11E9: dout  = 8'b10011001; // 4585 : 153 - 0x99
      13'h11EA: dout  = 8'b10001001; // 4586 : 137 - 0x89
      13'h11EB: dout  = 8'b10000001; // 4587 : 129 - 0x81
      13'h11EC: dout  = 8'b10000001; // 4588 : 129 - 0x81
      13'h11ED: dout  = 8'b10010001; // 4589 : 145 - 0x91
      13'h11EE: dout  = 8'b10011001; // 4590 : 153 - 0x99
      13'h11EF: dout  = 8'b10011001; // 4591 : 153 - 0x99
      13'h11F0: dout  = 8'b00111100; // 4592 :  60 - 0x3c -- Background 0x1f
      13'h11F1: dout  = 8'b01111110; // 4593 : 126 - 0x7e
      13'h11F2: dout  = 8'b11100111; // 4594 : 231 - 0xe7
      13'h11F3: dout  = 8'b11100111; // 4595 : 231 - 0xe7
      13'h11F4: dout  = 8'b11100111; // 4596 : 231 - 0xe7
      13'h11F5: dout  = 8'b11100111; // 4597 : 231 - 0xe7
      13'h11F6: dout  = 8'b01111110; // 4598 : 126 - 0x7e
      13'h11F7: dout  = 8'b00111100; // 4599 :  60 - 0x3c
      13'h11F8: dout  = 8'b11000111; // 4600 : 199 - 0xc7
      13'h11F9: dout  = 8'b10000011; // 4601 : 131 - 0x83
      13'h11FA: dout  = 8'b00111001; // 4602 :  57 - 0x39
      13'h11FB: dout  = 8'b00111001; // 4603 :  57 - 0x39
      13'h11FC: dout  = 8'b00111001; // 4604 :  57 - 0x39
      13'h11FD: dout  = 8'b00111001; // 4605 :  57 - 0x39
      13'h11FE: dout  = 8'b10000011; // 4606 : 131 - 0x83
      13'h11FF: dout  = 8'b11000111; // 4607 : 199 - 0xc7
      13'h1200: dout  = 8'b01111110; // 4608 : 126 - 0x7e -- Background 0x20
      13'h1201: dout  = 8'b01111111; // 4609 : 127 - 0x7f
      13'h1202: dout  = 8'b01110111; // 4610 : 119 - 0x77
      13'h1203: dout  = 8'b01110111; // 4611 : 119 - 0x77
      13'h1204: dout  = 8'b01111111; // 4612 : 127 - 0x7f
      13'h1205: dout  = 8'b01111110; // 4613 : 126 - 0x7e
      13'h1206: dout  = 8'b01110000; // 4614 : 112 - 0x70
      13'h1207: dout  = 8'b01110000; // 4615 : 112 - 0x70
      13'h1208: dout  = 8'b10000011; // 4616 : 131 - 0x83
      13'h1209: dout  = 8'b10000001; // 4617 : 129 - 0x81
      13'h120A: dout  = 8'b10011001; // 4618 : 153 - 0x99
      13'h120B: dout  = 8'b10011001; // 4619 : 153 - 0x99
      13'h120C: dout  = 8'b10000001; // 4620 : 129 - 0x81
      13'h120D: dout  = 8'b10000011; // 4621 : 131 - 0x83
      13'h120E: dout  = 8'b10011111; // 4622 : 159 - 0x9f
      13'h120F: dout  = 8'b10011111; // 4623 : 159 - 0x9f
      13'h1210: dout  = 8'b00111100; // 4624 :  60 - 0x3c -- Background 0x21
      13'h1211: dout  = 8'b01111110; // 4625 : 126 - 0x7e
      13'h1212: dout  = 8'b11100111; // 4626 : 231 - 0xe7
      13'h1213: dout  = 8'b11100111; // 4627 : 231 - 0xe7
      13'h1214: dout  = 8'b11100111; // 4628 : 231 - 0xe7
      13'h1215: dout  = 8'b11101110; // 4629 : 238 - 0xee
      13'h1216: dout  = 8'b01111111; // 4630 : 127 - 0x7f
      13'h1217: dout  = 8'b00111111; // 4631 :  63 - 0x3f
      13'h1218: dout  = 8'b11000111; // 4632 : 199 - 0xc7
      13'h1219: dout  = 8'b10000011; // 4633 : 131 - 0x83
      13'h121A: dout  = 8'b00111001; // 4634 :  57 - 0x39
      13'h121B: dout  = 8'b00111001; // 4635 :  57 - 0x39
      13'h121C: dout  = 8'b00111001; // 4636 :  57 - 0x39
      13'h121D: dout  = 8'b00110011; // 4637 :  51 - 0x33
      13'h121E: dout  = 8'b10000001; // 4638 : 129 - 0x81
      13'h121F: dout  = 8'b11001001; // 4639 : 201 - 0xc9
      13'h1220: dout  = 8'b01111110; // 4640 : 126 - 0x7e -- Background 0x22
      13'h1221: dout  = 8'b01111111; // 4641 : 127 - 0x7f
      13'h1222: dout  = 8'b01110111; // 4642 : 119 - 0x77
      13'h1223: dout  = 8'b01110111; // 4643 : 119 - 0x77
      13'h1224: dout  = 8'b01111111; // 4644 : 127 - 0x7f
      13'h1225: dout  = 8'b01111110; // 4645 : 126 - 0x7e
      13'h1226: dout  = 8'b01110111; // 4646 : 119 - 0x77
      13'h1227: dout  = 8'b01110111; // 4647 : 119 - 0x77
      13'h1228: dout  = 8'b10000011; // 4648 : 131 - 0x83
      13'h1229: dout  = 8'b10000001; // 4649 : 129 - 0x81
      13'h122A: dout  = 8'b10011001; // 4650 : 153 - 0x99
      13'h122B: dout  = 8'b10011001; // 4651 : 153 - 0x99
      13'h122C: dout  = 8'b10000001; // 4652 : 129 - 0x81
      13'h122D: dout  = 8'b10000011; // 4653 : 131 - 0x83
      13'h122E: dout  = 8'b10011001; // 4654 : 153 - 0x99
      13'h122F: dout  = 8'b10011001; // 4655 : 153 - 0x99
      13'h1230: dout  = 8'b00111110; // 4656 :  62 - 0x3e -- Background 0x23
      13'h1231: dout  = 8'b01111111; // 4657 : 127 - 0x7f
      13'h1232: dout  = 8'b01110000; // 4658 : 112 - 0x70
      13'h1233: dout  = 8'b01111110; // 4659 : 126 - 0x7e
      13'h1234: dout  = 8'b00111111; // 4660 :  63 - 0x3f
      13'h1235: dout  = 8'b00000111; // 4661 :   7 - 0x7
      13'h1236: dout  = 8'b01111111; // 4662 : 127 - 0x7f
      13'h1237: dout  = 8'b00111110; // 4663 :  62 - 0x3e
      13'h1238: dout  = 8'b11000011; // 4664 : 195 - 0xc3
      13'h1239: dout  = 8'b10000001; // 4665 : 129 - 0x81
      13'h123A: dout  = 8'b10011111; // 4666 : 159 - 0x9f
      13'h123B: dout  = 8'b10000011; // 4667 : 131 - 0x83
      13'h123C: dout  = 8'b11000001; // 4668 : 193 - 0xc1
      13'h123D: dout  = 8'b11111001; // 4669 : 249 - 0xf9
      13'h123E: dout  = 8'b10000001; // 4670 : 129 - 0x81
      13'h123F: dout  = 8'b11000011; // 4671 : 195 - 0xc3
      13'h1240: dout  = 8'b01111111; // 4672 : 127 - 0x7f -- Background 0x24
      13'h1241: dout  = 8'b01111111; // 4673 : 127 - 0x7f
      13'h1242: dout  = 8'b00011100; // 4674 :  28 - 0x1c
      13'h1243: dout  = 8'b00011100; // 4675 :  28 - 0x1c
      13'h1244: dout  = 8'b00011100; // 4676 :  28 - 0x1c
      13'h1245: dout  = 8'b00011100; // 4677 :  28 - 0x1c
      13'h1246: dout  = 8'b00011100; // 4678 :  28 - 0x1c
      13'h1247: dout  = 8'b00011100; // 4679 :  28 - 0x1c
      13'h1248: dout  = 8'b10000001; // 4680 : 129 - 0x81
      13'h1249: dout  = 8'b10000001; // 4681 : 129 - 0x81
      13'h124A: dout  = 8'b11100111; // 4682 : 231 - 0xe7
      13'h124B: dout  = 8'b11100111; // 4683 : 231 - 0xe7
      13'h124C: dout  = 8'b11100111; // 4684 : 231 - 0xe7
      13'h124D: dout  = 8'b11100111; // 4685 : 231 - 0xe7
      13'h124E: dout  = 8'b11100111; // 4686 : 231 - 0xe7
      13'h124F: dout  = 8'b11100111; // 4687 : 231 - 0xe7
      13'h1250: dout  = 8'b01110111; // 4688 : 119 - 0x77 -- Background 0x25
      13'h1251: dout  = 8'b01110111; // 4689 : 119 - 0x77
      13'h1252: dout  = 8'b01110111; // 4690 : 119 - 0x77
      13'h1253: dout  = 8'b01110111; // 4691 : 119 - 0x77
      13'h1254: dout  = 8'b01110111; // 4692 : 119 - 0x77
      13'h1255: dout  = 8'b01110111; // 4693 : 119 - 0x77
      13'h1256: dout  = 8'b01111111; // 4694 : 127 - 0x7f
      13'h1257: dout  = 8'b00111110; // 4695 :  62 - 0x3e
      13'h1258: dout  = 8'b10011001; // 4696 : 153 - 0x99
      13'h1259: dout  = 8'b10011001; // 4697 : 153 - 0x99
      13'h125A: dout  = 8'b10011001; // 4698 : 153 - 0x99
      13'h125B: dout  = 8'b10011001; // 4699 : 153 - 0x99
      13'h125C: dout  = 8'b10011001; // 4700 : 153 - 0x99
      13'h125D: dout  = 8'b10011001; // 4701 : 153 - 0x99
      13'h125E: dout  = 8'b10000001; // 4702 : 129 - 0x81
      13'h125F: dout  = 8'b11000011; // 4703 : 195 - 0xc3
      13'h1260: dout  = 8'b01110111; // 4704 : 119 - 0x77 -- Background 0x26
      13'h1261: dout  = 8'b01110111; // 4705 : 119 - 0x77
      13'h1262: dout  = 8'b01110111; // 4706 : 119 - 0x77
      13'h1263: dout  = 8'b01110111; // 4707 : 119 - 0x77
      13'h1264: dout  = 8'b01110111; // 4708 : 119 - 0x77
      13'h1265: dout  = 8'b01110111; // 4709 : 119 - 0x77
      13'h1266: dout  = 8'b00111110; // 4710 :  62 - 0x3e
      13'h1267: dout  = 8'b00011100; // 4711 :  28 - 0x1c
      13'h1268: dout  = 8'b10011001; // 4712 : 153 - 0x99
      13'h1269: dout  = 8'b10011001; // 4713 : 153 - 0x99
      13'h126A: dout  = 8'b10011001; // 4714 : 153 - 0x99
      13'h126B: dout  = 8'b10011001; // 4715 : 153 - 0x99
      13'h126C: dout  = 8'b10011001; // 4716 : 153 - 0x99
      13'h126D: dout  = 8'b10011001; // 4717 : 153 - 0x99
      13'h126E: dout  = 8'b11000011; // 4718 : 195 - 0xc3
      13'h126F: dout  = 8'b11100111; // 4719 : 231 - 0xe7
      13'h1270: dout  = 8'b11100111; // 4720 : 231 - 0xe7 -- Background 0x27
      13'h1271: dout  = 8'b11100111; // 4721 : 231 - 0xe7
      13'h1272: dout  = 8'b11100111; // 4722 : 231 - 0xe7
      13'h1273: dout  = 8'b11100111; // 4723 : 231 - 0xe7
      13'h1274: dout  = 8'b11110111; // 4724 : 247 - 0xf7
      13'h1275: dout  = 8'b11111111; // 4725 : 255 - 0xff
      13'h1276: dout  = 8'b11111111; // 4726 : 255 - 0xff
      13'h1277: dout  = 8'b01111110; // 4727 : 126 - 0x7e
      13'h1278: dout  = 8'b00111001; // 4728 :  57 - 0x39
      13'h1279: dout  = 8'b00111001; // 4729 :  57 - 0x39
      13'h127A: dout  = 8'b00111001; // 4730 :  57 - 0x39
      13'h127B: dout  = 8'b00111001; // 4731 :  57 - 0x39
      13'h127C: dout  = 8'b00101001; // 4732 :  41 - 0x29
      13'h127D: dout  = 8'b00000001; // 4733 :   1 - 0x1
      13'h127E: dout  = 8'b00000001; // 4734 :   1 - 0x1
      13'h127F: dout  = 8'b10010011; // 4735 : 147 - 0x93
      13'h1280: dout  = 8'b01110111; // 4736 : 119 - 0x77 -- Background 0x28
      13'h1281: dout  = 8'b01110111; // 4737 : 119 - 0x77
      13'h1282: dout  = 8'b01110111; // 4738 : 119 - 0x77
      13'h1283: dout  = 8'b00111110; // 4739 :  62 - 0x3e
      13'h1284: dout  = 8'b00111110; // 4740 :  62 - 0x3e
      13'h1285: dout  = 8'b01110111; // 4741 : 119 - 0x77
      13'h1286: dout  = 8'b01110111; // 4742 : 119 - 0x77
      13'h1287: dout  = 8'b01110111; // 4743 : 119 - 0x77
      13'h1288: dout  = 8'b10011001; // 4744 : 153 - 0x99
      13'h1289: dout  = 8'b10011001; // 4745 : 153 - 0x99
      13'h128A: dout  = 8'b10011001; // 4746 : 153 - 0x99
      13'h128B: dout  = 8'b11000011; // 4747 : 195 - 0xc3
      13'h128C: dout  = 8'b11000011; // 4748 : 195 - 0xc3
      13'h128D: dout  = 8'b10011001; // 4749 : 153 - 0x99
      13'h128E: dout  = 8'b10011001; // 4750 : 153 - 0x99
      13'h128F: dout  = 8'b10011001; // 4751 : 153 - 0x99
      13'h1290: dout  = 8'b01110111; // 4752 : 119 - 0x77 -- Background 0x29
      13'h1291: dout  = 8'b01110111; // 4753 : 119 - 0x77
      13'h1292: dout  = 8'b01110111; // 4754 : 119 - 0x77
      13'h1293: dout  = 8'b01111111; // 4755 : 127 - 0x7f
      13'h1294: dout  = 8'b00111110; // 4756 :  62 - 0x3e
      13'h1295: dout  = 8'b00011100; // 4757 :  28 - 0x1c
      13'h1296: dout  = 8'b00011100; // 4758 :  28 - 0x1c
      13'h1297: dout  = 8'b00011100; // 4759 :  28 - 0x1c
      13'h1298: dout  = 8'b10011001; // 4760 : 153 - 0x99
      13'h1299: dout  = 8'b10011001; // 4761 : 153 - 0x99
      13'h129A: dout  = 8'b10011001; // 4762 : 153 - 0x99
      13'h129B: dout  = 8'b10000001; // 4763 : 129 - 0x81
      13'h129C: dout  = 8'b11000011; // 4764 : 195 - 0xc3
      13'h129D: dout  = 8'b11100111; // 4765 : 231 - 0xe7
      13'h129E: dout  = 8'b11100111; // 4766 : 231 - 0xe7
      13'h129F: dout  = 8'b11100111; // 4767 : 231 - 0xe7
      13'h12A0: dout  = 8'b01111111; // 4768 : 127 - 0x7f -- Background 0x2a
      13'h12A1: dout  = 8'b01111111; // 4769 : 127 - 0x7f
      13'h12A2: dout  = 8'b00001110; // 4770 :  14 - 0xe
      13'h12A3: dout  = 8'b00011100; // 4771 :  28 - 0x1c
      13'h12A4: dout  = 8'b00011100; // 4772 :  28 - 0x1c
      13'h12A5: dout  = 8'b00111000; // 4773 :  56 - 0x38
      13'h12A6: dout  = 8'b01111111; // 4774 : 127 - 0x7f
      13'h12A7: dout  = 8'b01111111; // 4775 : 127 - 0x7f
      13'h12A8: dout  = 8'b10000001; // 4776 : 129 - 0x81
      13'h12A9: dout  = 8'b10000001; // 4777 : 129 - 0x81
      13'h12AA: dout  = 8'b11110011; // 4778 : 243 - 0xf3
      13'h12AB: dout  = 8'b11100111; // 4779 : 231 - 0xe7
      13'h12AC: dout  = 8'b11100111; // 4780 : 231 - 0xe7
      13'h12AD: dout  = 8'b11001111; // 4781 : 207 - 0xcf
      13'h12AE: dout  = 8'b10000001; // 4782 : 129 - 0x81
      13'h12AF: dout  = 8'b10000001; // 4783 : 129 - 0x81
      13'h12B0: dout  = 8'b00111110; // 4784 :  62 - 0x3e -- Background 0x2b
      13'h12B1: dout  = 8'b01100011; // 4785 :  99 - 0x63
      13'h12B2: dout  = 8'b01101111; // 4786 : 111 - 0x6f
      13'h12B3: dout  = 8'b01111111; // 4787 : 127 - 0x7f
      13'h12B4: dout  = 8'b01111111; // 4788 : 127 - 0x7f
      13'h12B5: dout  = 8'b01111110; // 4789 : 126 - 0x7e
      13'h12B6: dout  = 8'b01100000; // 4790 :  96 - 0x60
      13'h12B7: dout  = 8'b00111111; // 4791 :  63 - 0x3f
      13'h12B8: dout  = 8'b11000011; // 4792 : 195 - 0xc3
      13'h12B9: dout  = 8'b10111101; // 4793 : 189 - 0xbd
      13'h12BA: dout  = 8'b10110101; // 4794 : 181 - 0xb5
      13'h12BB: dout  = 8'b10101001; // 4795 : 169 - 0xa9
      13'h12BC: dout  = 8'b10101001; // 4796 : 169 - 0xa9
      13'h12BD: dout  = 8'b10100011; // 4797 : 163 - 0xa3
      13'h12BE: dout  = 8'b10111111; // 4798 : 191 - 0xbf
      13'h12BF: dout  = 8'b11000001; // 4799 : 193 - 0xc1
      13'h12C0: dout  = 8'b00000000; // 4800 :   0 - 0x0 -- Background 0x2c
      13'h12C1: dout  = 8'b01110000; // 4801 : 112 - 0x70
      13'h12C2: dout  = 8'b01111100; // 4802 : 124 - 0x7c
      13'h12C3: dout  = 8'b01111111; // 4803 : 127 - 0x7f
      13'h12C4: dout  = 8'b01111111; // 4804 : 127 - 0x7f
      13'h12C5: dout  = 8'b01111100; // 4805 : 124 - 0x7c
      13'h12C6: dout  = 8'b01110000; // 4806 : 112 - 0x70
      13'h12C7: dout  = 8'b00000000; // 4807 :   0 - 0x0
      13'h12C8: dout  = 8'b11111111; // 4808 : 255 - 0xff
      13'h12C9: dout  = 8'b10011111; // 4809 : 159 - 0x9f
      13'h12CA: dout  = 8'b10000111; // 4810 : 135 - 0x87
      13'h12CB: dout  = 8'b10000001; // 4811 : 129 - 0x81
      13'h12CC: dout  = 8'b10000001; // 4812 : 129 - 0x81
      13'h12CD: dout  = 8'b10000111; // 4813 : 135 - 0x87
      13'h12CE: dout  = 8'b10011111; // 4814 : 159 - 0x9f
      13'h12CF: dout  = 8'b11111111; // 4815 : 255 - 0xff
      13'h12D0: dout  = 8'b00000000; // 4816 :   0 - 0x0 -- Background 0x2d
      13'h12D1: dout  = 8'b01110000; // 4817 : 112 - 0x70
      13'h12D2: dout  = 8'b01110000; // 4818 : 112 - 0x70
      13'h12D3: dout  = 8'b00000000; // 4819 :   0 - 0x0
      13'h12D4: dout  = 8'b00000000; // 4820 :   0 - 0x0
      13'h12D5: dout  = 8'b01110000; // 4821 : 112 - 0x70
      13'h12D6: dout  = 8'b01110000; // 4822 : 112 - 0x70
      13'h12D7: dout  = 8'b00000000; // 4823 :   0 - 0x0
      13'h12D8: dout  = 8'b11111111; // 4824 : 255 - 0xff
      13'h12D9: dout  = 8'b10011111; // 4825 : 159 - 0x9f
      13'h12DA: dout  = 8'b10011111; // 4826 : 159 - 0x9f
      13'h12DB: dout  = 8'b11111111; // 4827 : 255 - 0xff
      13'h12DC: dout  = 8'b11111111; // 4828 : 255 - 0xff
      13'h12DD: dout  = 8'b10011111; // 4829 : 159 - 0x9f
      13'h12DE: dout  = 8'b10011111; // 4830 : 159 - 0x9f
      13'h12DF: dout  = 8'b11111111; // 4831 : 255 - 0xff
      13'h12E0: dout  = 8'b00000000; // 4832 :   0 - 0x0 -- Background 0x2e
      13'h12E1: dout  = 8'b00000000; // 4833 :   0 - 0x0
      13'h12E2: dout  = 8'b00000000; // 4834 :   0 - 0x0
      13'h12E3: dout  = 8'b00000000; // 4835 :   0 - 0x0
      13'h12E4: dout  = 8'b00000000; // 4836 :   0 - 0x0
      13'h12E5: dout  = 8'b00000000; // 4837 :   0 - 0x0
      13'h12E6: dout  = 8'b00000000; // 4838 :   0 - 0x0
      13'h12E7: dout  = 8'b00000000; // 4839 :   0 - 0x0
      13'h12E8: dout  = 8'b00000000; // 4840 :   0 - 0x0
      13'h12E9: dout  = 8'b00000000; // 4841 :   0 - 0x0
      13'h12EA: dout  = 8'b00000000; // 4842 :   0 - 0x0
      13'h12EB: dout  = 8'b00000000; // 4843 :   0 - 0x0
      13'h12EC: dout  = 8'b00000000; // 4844 :   0 - 0x0
      13'h12ED: dout  = 8'b00000000; // 4845 :   0 - 0x0
      13'h12EE: dout  = 8'b00000000; // 4846 :   0 - 0x0
      13'h12EF: dout  = 8'b00000000; // 4847 :   0 - 0x0
      13'h12F0: dout  = 8'b00000000; // 4848 :   0 - 0x0 -- Background 0x2f
      13'h12F1: dout  = 8'b00000000; // 4849 :   0 - 0x0
      13'h12F2: dout  = 8'b00000000; // 4850 :   0 - 0x0
      13'h12F3: dout  = 8'b00000000; // 4851 :   0 - 0x0
      13'h12F4: dout  = 8'b00000000; // 4852 :   0 - 0x0
      13'h12F5: dout  = 8'b00000000; // 4853 :   0 - 0x0
      13'h12F6: dout  = 8'b00000000; // 4854 :   0 - 0x0
      13'h12F7: dout  = 8'b00000000; // 4855 :   0 - 0x0
      13'h12F8: dout  = 8'b00000000; // 4856 :   0 - 0x0
      13'h12F9: dout  = 8'b00000000; // 4857 :   0 - 0x0
      13'h12FA: dout  = 8'b00000000; // 4858 :   0 - 0x0
      13'h12FB: dout  = 8'b00000000; // 4859 :   0 - 0x0
      13'h12FC: dout  = 8'b00000000; // 4860 :   0 - 0x0
      13'h12FD: dout  = 8'b00000000; // 4861 :   0 - 0x0
      13'h12FE: dout  = 8'b00000000; // 4862 :   0 - 0x0
      13'h12FF: dout  = 8'b00000000; // 4863 :   0 - 0x0
      13'h1300: dout  = 8'b00000000; // 4864 :   0 - 0x0 -- Background 0x30
      13'h1301: dout  = 8'b00000000; // 4865 :   0 - 0x0
      13'h1302: dout  = 8'b00000000; // 4866 :   0 - 0x0
      13'h1303: dout  = 8'b00000000; // 4867 :   0 - 0x0
      13'h1304: dout  = 8'b00000000; // 4868 :   0 - 0x0
      13'h1305: dout  = 8'b00000000; // 4869 :   0 - 0x0
      13'h1306: dout  = 8'b00000000; // 4870 :   0 - 0x0
      13'h1307: dout  = 8'b00000000; // 4871 :   0 - 0x0
      13'h1308: dout  = 8'b00000000; // 4872 :   0 - 0x0
      13'h1309: dout  = 8'b00000000; // 4873 :   0 - 0x0
      13'h130A: dout  = 8'b00000000; // 4874 :   0 - 0x0
      13'h130B: dout  = 8'b00000000; // 4875 :   0 - 0x0
      13'h130C: dout  = 8'b00000000; // 4876 :   0 - 0x0
      13'h130D: dout  = 8'b00000000; // 4877 :   0 - 0x0
      13'h130E: dout  = 8'b00000000; // 4878 :   0 - 0x0
      13'h130F: dout  = 8'b00000000; // 4879 :   0 - 0x0
      13'h1310: dout  = 8'b00000000; // 4880 :   0 - 0x0 -- Background 0x31
      13'h1311: dout  = 8'b00000000; // 4881 :   0 - 0x0
      13'h1312: dout  = 8'b00000000; // 4882 :   0 - 0x0
      13'h1313: dout  = 8'b00000000; // 4883 :   0 - 0x0
      13'h1314: dout  = 8'b00000000; // 4884 :   0 - 0x0
      13'h1315: dout  = 8'b00000000; // 4885 :   0 - 0x0
      13'h1316: dout  = 8'b00000000; // 4886 :   0 - 0x0
      13'h1317: dout  = 8'b00000000; // 4887 :   0 - 0x0
      13'h1318: dout  = 8'b00000000; // 4888 :   0 - 0x0
      13'h1319: dout  = 8'b00000000; // 4889 :   0 - 0x0
      13'h131A: dout  = 8'b00000000; // 4890 :   0 - 0x0
      13'h131B: dout  = 8'b00000000; // 4891 :   0 - 0x0
      13'h131C: dout  = 8'b00000000; // 4892 :   0 - 0x0
      13'h131D: dout  = 8'b00000000; // 4893 :   0 - 0x0
      13'h131E: dout  = 8'b00000000; // 4894 :   0 - 0x0
      13'h131F: dout  = 8'b00000000; // 4895 :   0 - 0x0
      13'h1320: dout  = 8'b00000000; // 4896 :   0 - 0x0 -- Background 0x32
      13'h1321: dout  = 8'b00000000; // 4897 :   0 - 0x0
      13'h1322: dout  = 8'b00000000; // 4898 :   0 - 0x0
      13'h1323: dout  = 8'b00000000; // 4899 :   0 - 0x0
      13'h1324: dout  = 8'b00000000; // 4900 :   0 - 0x0
      13'h1325: dout  = 8'b00000000; // 4901 :   0 - 0x0
      13'h1326: dout  = 8'b00000000; // 4902 :   0 - 0x0
      13'h1327: dout  = 8'b00000000; // 4903 :   0 - 0x0
      13'h1328: dout  = 8'b00000000; // 4904 :   0 - 0x0
      13'h1329: dout  = 8'b00000000; // 4905 :   0 - 0x0
      13'h132A: dout  = 8'b00000000; // 4906 :   0 - 0x0
      13'h132B: dout  = 8'b00000000; // 4907 :   0 - 0x0
      13'h132C: dout  = 8'b00000000; // 4908 :   0 - 0x0
      13'h132D: dout  = 8'b00000000; // 4909 :   0 - 0x0
      13'h132E: dout  = 8'b00000000; // 4910 :   0 - 0x0
      13'h132F: dout  = 8'b00000000; // 4911 :   0 - 0x0
      13'h1330: dout  = 8'b00000000; // 4912 :   0 - 0x0 -- Background 0x33
      13'h1331: dout  = 8'b00000000; // 4913 :   0 - 0x0
      13'h1332: dout  = 8'b00000000; // 4914 :   0 - 0x0
      13'h1333: dout  = 8'b00000000; // 4915 :   0 - 0x0
      13'h1334: dout  = 8'b00000000; // 4916 :   0 - 0x0
      13'h1335: dout  = 8'b00000000; // 4917 :   0 - 0x0
      13'h1336: dout  = 8'b00000000; // 4918 :   0 - 0x0
      13'h1337: dout  = 8'b00000000; // 4919 :   0 - 0x0
      13'h1338: dout  = 8'b00000000; // 4920 :   0 - 0x0
      13'h1339: dout  = 8'b00000000; // 4921 :   0 - 0x0
      13'h133A: dout  = 8'b00000000; // 4922 :   0 - 0x0
      13'h133B: dout  = 8'b00000000; // 4923 :   0 - 0x0
      13'h133C: dout  = 8'b00000000; // 4924 :   0 - 0x0
      13'h133D: dout  = 8'b00000000; // 4925 :   0 - 0x0
      13'h133E: dout  = 8'b00000000; // 4926 :   0 - 0x0
      13'h133F: dout  = 8'b00000000; // 4927 :   0 - 0x0
      13'h1340: dout  = 8'b00000000; // 4928 :   0 - 0x0 -- Background 0x34
      13'h1341: dout  = 8'b00000000; // 4929 :   0 - 0x0
      13'h1342: dout  = 8'b00000000; // 4930 :   0 - 0x0
      13'h1343: dout  = 8'b00000000; // 4931 :   0 - 0x0
      13'h1344: dout  = 8'b00000000; // 4932 :   0 - 0x0
      13'h1345: dout  = 8'b00000000; // 4933 :   0 - 0x0
      13'h1346: dout  = 8'b00000000; // 4934 :   0 - 0x0
      13'h1347: dout  = 8'b00000000; // 4935 :   0 - 0x0
      13'h1348: dout  = 8'b00000000; // 4936 :   0 - 0x0
      13'h1349: dout  = 8'b00000000; // 4937 :   0 - 0x0
      13'h134A: dout  = 8'b00000000; // 4938 :   0 - 0x0
      13'h134B: dout  = 8'b00000000; // 4939 :   0 - 0x0
      13'h134C: dout  = 8'b00000000; // 4940 :   0 - 0x0
      13'h134D: dout  = 8'b00000000; // 4941 :   0 - 0x0
      13'h134E: dout  = 8'b00000000; // 4942 :   0 - 0x0
      13'h134F: dout  = 8'b00000000; // 4943 :   0 - 0x0
      13'h1350: dout  = 8'b00000000; // 4944 :   0 - 0x0 -- Background 0x35
      13'h1351: dout  = 8'b00000000; // 4945 :   0 - 0x0
      13'h1352: dout  = 8'b00000000; // 4946 :   0 - 0x0
      13'h1353: dout  = 8'b00000000; // 4947 :   0 - 0x0
      13'h1354: dout  = 8'b00000000; // 4948 :   0 - 0x0
      13'h1355: dout  = 8'b00000000; // 4949 :   0 - 0x0
      13'h1356: dout  = 8'b00000000; // 4950 :   0 - 0x0
      13'h1357: dout  = 8'b00000000; // 4951 :   0 - 0x0
      13'h1358: dout  = 8'b00000000; // 4952 :   0 - 0x0
      13'h1359: dout  = 8'b00000000; // 4953 :   0 - 0x0
      13'h135A: dout  = 8'b00000000; // 4954 :   0 - 0x0
      13'h135B: dout  = 8'b00000000; // 4955 :   0 - 0x0
      13'h135C: dout  = 8'b00000000; // 4956 :   0 - 0x0
      13'h135D: dout  = 8'b00000000; // 4957 :   0 - 0x0
      13'h135E: dout  = 8'b00000000; // 4958 :   0 - 0x0
      13'h135F: dout  = 8'b00000000; // 4959 :   0 - 0x0
      13'h1360: dout  = 8'b00000000; // 4960 :   0 - 0x0 -- Background 0x36
      13'h1361: dout  = 8'b00000000; // 4961 :   0 - 0x0
      13'h1362: dout  = 8'b00000000; // 4962 :   0 - 0x0
      13'h1363: dout  = 8'b00000000; // 4963 :   0 - 0x0
      13'h1364: dout  = 8'b00000000; // 4964 :   0 - 0x0
      13'h1365: dout  = 8'b00000000; // 4965 :   0 - 0x0
      13'h1366: dout  = 8'b00000000; // 4966 :   0 - 0x0
      13'h1367: dout  = 8'b00000000; // 4967 :   0 - 0x0
      13'h1368: dout  = 8'b00000000; // 4968 :   0 - 0x0
      13'h1369: dout  = 8'b00000000; // 4969 :   0 - 0x0
      13'h136A: dout  = 8'b00000000; // 4970 :   0 - 0x0
      13'h136B: dout  = 8'b00000000; // 4971 :   0 - 0x0
      13'h136C: dout  = 8'b00000000; // 4972 :   0 - 0x0
      13'h136D: dout  = 8'b00000000; // 4973 :   0 - 0x0
      13'h136E: dout  = 8'b00000000; // 4974 :   0 - 0x0
      13'h136F: dout  = 8'b00000000; // 4975 :   0 - 0x0
      13'h1370: dout  = 8'b00000000; // 4976 :   0 - 0x0 -- Background 0x37
      13'h1371: dout  = 8'b00000000; // 4977 :   0 - 0x0
      13'h1372: dout  = 8'b00000000; // 4978 :   0 - 0x0
      13'h1373: dout  = 8'b00000000; // 4979 :   0 - 0x0
      13'h1374: dout  = 8'b00000000; // 4980 :   0 - 0x0
      13'h1375: dout  = 8'b00000000; // 4981 :   0 - 0x0
      13'h1376: dout  = 8'b00000000; // 4982 :   0 - 0x0
      13'h1377: dout  = 8'b00000000; // 4983 :   0 - 0x0
      13'h1378: dout  = 8'b00000000; // 4984 :   0 - 0x0
      13'h1379: dout  = 8'b00000000; // 4985 :   0 - 0x0
      13'h137A: dout  = 8'b00000000; // 4986 :   0 - 0x0
      13'h137B: dout  = 8'b00000000; // 4987 :   0 - 0x0
      13'h137C: dout  = 8'b00000000; // 4988 :   0 - 0x0
      13'h137D: dout  = 8'b00000000; // 4989 :   0 - 0x0
      13'h137E: dout  = 8'b00000000; // 4990 :   0 - 0x0
      13'h137F: dout  = 8'b00000000; // 4991 :   0 - 0x0
      13'h1380: dout  = 8'b00000000; // 4992 :   0 - 0x0 -- Background 0x38
      13'h1381: dout  = 8'b00000000; // 4993 :   0 - 0x0
      13'h1382: dout  = 8'b00000000; // 4994 :   0 - 0x0
      13'h1383: dout  = 8'b00000000; // 4995 :   0 - 0x0
      13'h1384: dout  = 8'b00000000; // 4996 :   0 - 0x0
      13'h1385: dout  = 8'b00000000; // 4997 :   0 - 0x0
      13'h1386: dout  = 8'b00000000; // 4998 :   0 - 0x0
      13'h1387: dout  = 8'b00000000; // 4999 :   0 - 0x0
      13'h1388: dout  = 8'b00000000; // 5000 :   0 - 0x0
      13'h1389: dout  = 8'b00000000; // 5001 :   0 - 0x0
      13'h138A: dout  = 8'b00000000; // 5002 :   0 - 0x0
      13'h138B: dout  = 8'b00000000; // 5003 :   0 - 0x0
      13'h138C: dout  = 8'b00000000; // 5004 :   0 - 0x0
      13'h138D: dout  = 8'b00000000; // 5005 :   0 - 0x0
      13'h138E: dout  = 8'b00000000; // 5006 :   0 - 0x0
      13'h138F: dout  = 8'b00000000; // 5007 :   0 - 0x0
      13'h1390: dout  = 8'b00000000; // 5008 :   0 - 0x0 -- Background 0x39
      13'h1391: dout  = 8'b00000000; // 5009 :   0 - 0x0
      13'h1392: dout  = 8'b00000000; // 5010 :   0 - 0x0
      13'h1393: dout  = 8'b00000000; // 5011 :   0 - 0x0
      13'h1394: dout  = 8'b00000000; // 5012 :   0 - 0x0
      13'h1395: dout  = 8'b00000000; // 5013 :   0 - 0x0
      13'h1396: dout  = 8'b00000000; // 5014 :   0 - 0x0
      13'h1397: dout  = 8'b00000000; // 5015 :   0 - 0x0
      13'h1398: dout  = 8'b00000000; // 5016 :   0 - 0x0
      13'h1399: dout  = 8'b00000000; // 5017 :   0 - 0x0
      13'h139A: dout  = 8'b00000000; // 5018 :   0 - 0x0
      13'h139B: dout  = 8'b00000000; // 5019 :   0 - 0x0
      13'h139C: dout  = 8'b00000000; // 5020 :   0 - 0x0
      13'h139D: dout  = 8'b00000000; // 5021 :   0 - 0x0
      13'h139E: dout  = 8'b00000000; // 5022 :   0 - 0x0
      13'h139F: dout  = 8'b00000000; // 5023 :   0 - 0x0
      13'h13A0: dout  = 8'b00000000; // 5024 :   0 - 0x0 -- Background 0x3a
      13'h13A1: dout  = 8'b00000000; // 5025 :   0 - 0x0
      13'h13A2: dout  = 8'b00000000; // 5026 :   0 - 0x0
      13'h13A3: dout  = 8'b00000000; // 5027 :   0 - 0x0
      13'h13A4: dout  = 8'b00000000; // 5028 :   0 - 0x0
      13'h13A5: dout  = 8'b00000000; // 5029 :   0 - 0x0
      13'h13A6: dout  = 8'b00000000; // 5030 :   0 - 0x0
      13'h13A7: dout  = 8'b00000000; // 5031 :   0 - 0x0
      13'h13A8: dout  = 8'b00000000; // 5032 :   0 - 0x0
      13'h13A9: dout  = 8'b00000000; // 5033 :   0 - 0x0
      13'h13AA: dout  = 8'b00000000; // 5034 :   0 - 0x0
      13'h13AB: dout  = 8'b00000000; // 5035 :   0 - 0x0
      13'h13AC: dout  = 8'b00000000; // 5036 :   0 - 0x0
      13'h13AD: dout  = 8'b00000000; // 5037 :   0 - 0x0
      13'h13AE: dout  = 8'b00000000; // 5038 :   0 - 0x0
      13'h13AF: dout  = 8'b00000000; // 5039 :   0 - 0x0
      13'h13B0: dout  = 8'b00000000; // 5040 :   0 - 0x0 -- Background 0x3b
      13'h13B1: dout  = 8'b00000000; // 5041 :   0 - 0x0
      13'h13B2: dout  = 8'b00000000; // 5042 :   0 - 0x0
      13'h13B3: dout  = 8'b00000000; // 5043 :   0 - 0x0
      13'h13B4: dout  = 8'b00000000; // 5044 :   0 - 0x0
      13'h13B5: dout  = 8'b00000000; // 5045 :   0 - 0x0
      13'h13B6: dout  = 8'b00000000; // 5046 :   0 - 0x0
      13'h13B7: dout  = 8'b00000000; // 5047 :   0 - 0x0
      13'h13B8: dout  = 8'b00000000; // 5048 :   0 - 0x0
      13'h13B9: dout  = 8'b00000000; // 5049 :   0 - 0x0
      13'h13BA: dout  = 8'b00000000; // 5050 :   0 - 0x0
      13'h13BB: dout  = 8'b00000000; // 5051 :   0 - 0x0
      13'h13BC: dout  = 8'b00000000; // 5052 :   0 - 0x0
      13'h13BD: dout  = 8'b00000000; // 5053 :   0 - 0x0
      13'h13BE: dout  = 8'b00000000; // 5054 :   0 - 0x0
      13'h13BF: dout  = 8'b00000000; // 5055 :   0 - 0x0
      13'h13C0: dout  = 8'b00000000; // 5056 :   0 - 0x0 -- Background 0x3c
      13'h13C1: dout  = 8'b00000000; // 5057 :   0 - 0x0
      13'h13C2: dout  = 8'b00000000; // 5058 :   0 - 0x0
      13'h13C3: dout  = 8'b00000000; // 5059 :   0 - 0x0
      13'h13C4: dout  = 8'b00000000; // 5060 :   0 - 0x0
      13'h13C5: dout  = 8'b00000000; // 5061 :   0 - 0x0
      13'h13C6: dout  = 8'b00000000; // 5062 :   0 - 0x0
      13'h13C7: dout  = 8'b00000000; // 5063 :   0 - 0x0
      13'h13C8: dout  = 8'b00000000; // 5064 :   0 - 0x0
      13'h13C9: dout  = 8'b00000000; // 5065 :   0 - 0x0
      13'h13CA: dout  = 8'b00000000; // 5066 :   0 - 0x0
      13'h13CB: dout  = 8'b00000000; // 5067 :   0 - 0x0
      13'h13CC: dout  = 8'b00000000; // 5068 :   0 - 0x0
      13'h13CD: dout  = 8'b00000000; // 5069 :   0 - 0x0
      13'h13CE: dout  = 8'b00000000; // 5070 :   0 - 0x0
      13'h13CF: dout  = 8'b00000000; // 5071 :   0 - 0x0
      13'h13D0: dout  = 8'b00000000; // 5072 :   0 - 0x0 -- Background 0x3d
      13'h13D1: dout  = 8'b00000000; // 5073 :   0 - 0x0
      13'h13D2: dout  = 8'b00000000; // 5074 :   0 - 0x0
      13'h13D3: dout  = 8'b00000000; // 5075 :   0 - 0x0
      13'h13D4: dout  = 8'b00000000; // 5076 :   0 - 0x0
      13'h13D5: dout  = 8'b00000000; // 5077 :   0 - 0x0
      13'h13D6: dout  = 8'b00000000; // 5078 :   0 - 0x0
      13'h13D7: dout  = 8'b00000000; // 5079 :   0 - 0x0
      13'h13D8: dout  = 8'b00000000; // 5080 :   0 - 0x0
      13'h13D9: dout  = 8'b00000000; // 5081 :   0 - 0x0
      13'h13DA: dout  = 8'b00000000; // 5082 :   0 - 0x0
      13'h13DB: dout  = 8'b00000000; // 5083 :   0 - 0x0
      13'h13DC: dout  = 8'b00000000; // 5084 :   0 - 0x0
      13'h13DD: dout  = 8'b00000000; // 5085 :   0 - 0x0
      13'h13DE: dout  = 8'b00000000; // 5086 :   0 - 0x0
      13'h13DF: dout  = 8'b00000000; // 5087 :   0 - 0x0
      13'h13E0: dout  = 8'b00000000; // 5088 :   0 - 0x0 -- Background 0x3e
      13'h13E1: dout  = 8'b00000000; // 5089 :   0 - 0x0
      13'h13E2: dout  = 8'b00000000; // 5090 :   0 - 0x0
      13'h13E3: dout  = 8'b00000000; // 5091 :   0 - 0x0
      13'h13E4: dout  = 8'b00000000; // 5092 :   0 - 0x0
      13'h13E5: dout  = 8'b00000000; // 5093 :   0 - 0x0
      13'h13E6: dout  = 8'b00000000; // 5094 :   0 - 0x0
      13'h13E7: dout  = 8'b00000000; // 5095 :   0 - 0x0
      13'h13E8: dout  = 8'b00000000; // 5096 :   0 - 0x0
      13'h13E9: dout  = 8'b00000000; // 5097 :   0 - 0x0
      13'h13EA: dout  = 8'b00000000; // 5098 :   0 - 0x0
      13'h13EB: dout  = 8'b00000000; // 5099 :   0 - 0x0
      13'h13EC: dout  = 8'b00000000; // 5100 :   0 - 0x0
      13'h13ED: dout  = 8'b00000000; // 5101 :   0 - 0x0
      13'h13EE: dout  = 8'b00000000; // 5102 :   0 - 0x0
      13'h13EF: dout  = 8'b00000000; // 5103 :   0 - 0x0
      13'h13F0: dout  = 8'b00000000; // 5104 :   0 - 0x0 -- Background 0x3f
      13'h13F1: dout  = 8'b00000000; // 5105 :   0 - 0x0
      13'h13F2: dout  = 8'b00000000; // 5106 :   0 - 0x0
      13'h13F3: dout  = 8'b00000000; // 5107 :   0 - 0x0
      13'h13F4: dout  = 8'b00000000; // 5108 :   0 - 0x0
      13'h13F5: dout  = 8'b00000000; // 5109 :   0 - 0x0
      13'h13F6: dout  = 8'b00000000; // 5110 :   0 - 0x0
      13'h13F7: dout  = 8'b00000000; // 5111 :   0 - 0x0
      13'h13F8: dout  = 8'b00000000; // 5112 :   0 - 0x0
      13'h13F9: dout  = 8'b00000000; // 5113 :   0 - 0x0
      13'h13FA: dout  = 8'b00000000; // 5114 :   0 - 0x0
      13'h13FB: dout  = 8'b00000000; // 5115 :   0 - 0x0
      13'h13FC: dout  = 8'b00000000; // 5116 :   0 - 0x0
      13'h13FD: dout  = 8'b00000000; // 5117 :   0 - 0x0
      13'h13FE: dout  = 8'b00000000; // 5118 :   0 - 0x0
      13'h13FF: dout  = 8'b00000000; // 5119 :   0 - 0x0
      13'h1400: dout  = 8'b00000000; // 5120 :   0 - 0x0 -- Background 0x40
      13'h1401: dout  = 8'b00000000; // 5121 :   0 - 0x0
      13'h1402: dout  = 8'b00000000; // 5122 :   0 - 0x0
      13'h1403: dout  = 8'b00000000; // 5123 :   0 - 0x0
      13'h1404: dout  = 8'b00000000; // 5124 :   0 - 0x0
      13'h1405: dout  = 8'b00000000; // 5125 :   0 - 0x0
      13'h1406: dout  = 8'b00000000; // 5126 :   0 - 0x0
      13'h1407: dout  = 8'b00000000; // 5127 :   0 - 0x0
      13'h1408: dout  = 8'b00000000; // 5128 :   0 - 0x0
      13'h1409: dout  = 8'b00000000; // 5129 :   0 - 0x0
      13'h140A: dout  = 8'b00000000; // 5130 :   0 - 0x0
      13'h140B: dout  = 8'b00000000; // 5131 :   0 - 0x0
      13'h140C: dout  = 8'b00000000; // 5132 :   0 - 0x0
      13'h140D: dout  = 8'b00000000; // 5133 :   0 - 0x0
      13'h140E: dout  = 8'b00000000; // 5134 :   0 - 0x0
      13'h140F: dout  = 8'b00000000; // 5135 :   0 - 0x0
      13'h1410: dout  = 8'b00000000; // 5136 :   0 - 0x0 -- Background 0x41
      13'h1411: dout  = 8'b00000000; // 5137 :   0 - 0x0
      13'h1412: dout  = 8'b00000000; // 5138 :   0 - 0x0
      13'h1413: dout  = 8'b00000000; // 5139 :   0 - 0x0
      13'h1414: dout  = 8'b00000000; // 5140 :   0 - 0x0
      13'h1415: dout  = 8'b00000000; // 5141 :   0 - 0x0
      13'h1416: dout  = 8'b00000000; // 5142 :   0 - 0x0
      13'h1417: dout  = 8'b00000000; // 5143 :   0 - 0x0
      13'h1418: dout  = 8'b00000000; // 5144 :   0 - 0x0
      13'h1419: dout  = 8'b00000000; // 5145 :   0 - 0x0
      13'h141A: dout  = 8'b00000000; // 5146 :   0 - 0x0
      13'h141B: dout  = 8'b00000000; // 5147 :   0 - 0x0
      13'h141C: dout  = 8'b00000000; // 5148 :   0 - 0x0
      13'h141D: dout  = 8'b00000000; // 5149 :   0 - 0x0
      13'h141E: dout  = 8'b00000000; // 5150 :   0 - 0x0
      13'h141F: dout  = 8'b00000000; // 5151 :   0 - 0x0
      13'h1420: dout  = 8'b00000000; // 5152 :   0 - 0x0 -- Background 0x42
      13'h1421: dout  = 8'b00000000; // 5153 :   0 - 0x0
      13'h1422: dout  = 8'b00000000; // 5154 :   0 - 0x0
      13'h1423: dout  = 8'b00000000; // 5155 :   0 - 0x0
      13'h1424: dout  = 8'b00000000; // 5156 :   0 - 0x0
      13'h1425: dout  = 8'b00000000; // 5157 :   0 - 0x0
      13'h1426: dout  = 8'b00000000; // 5158 :   0 - 0x0
      13'h1427: dout  = 8'b00000000; // 5159 :   0 - 0x0
      13'h1428: dout  = 8'b00000000; // 5160 :   0 - 0x0
      13'h1429: dout  = 8'b00000000; // 5161 :   0 - 0x0
      13'h142A: dout  = 8'b00000000; // 5162 :   0 - 0x0
      13'h142B: dout  = 8'b00000000; // 5163 :   0 - 0x0
      13'h142C: dout  = 8'b00000000; // 5164 :   0 - 0x0
      13'h142D: dout  = 8'b00000000; // 5165 :   0 - 0x0
      13'h142E: dout  = 8'b00000000; // 5166 :   0 - 0x0
      13'h142F: dout  = 8'b00000000; // 5167 :   0 - 0x0
      13'h1430: dout  = 8'b00000000; // 5168 :   0 - 0x0 -- Background 0x43
      13'h1431: dout  = 8'b00000000; // 5169 :   0 - 0x0
      13'h1432: dout  = 8'b00000000; // 5170 :   0 - 0x0
      13'h1433: dout  = 8'b00000000; // 5171 :   0 - 0x0
      13'h1434: dout  = 8'b00000000; // 5172 :   0 - 0x0
      13'h1435: dout  = 8'b00000000; // 5173 :   0 - 0x0
      13'h1436: dout  = 8'b00000000; // 5174 :   0 - 0x0
      13'h1437: dout  = 8'b00000000; // 5175 :   0 - 0x0
      13'h1438: dout  = 8'b00000000; // 5176 :   0 - 0x0
      13'h1439: dout  = 8'b00000000; // 5177 :   0 - 0x0
      13'h143A: dout  = 8'b00000000; // 5178 :   0 - 0x0
      13'h143B: dout  = 8'b00000000; // 5179 :   0 - 0x0
      13'h143C: dout  = 8'b00000000; // 5180 :   0 - 0x0
      13'h143D: dout  = 8'b00000000; // 5181 :   0 - 0x0
      13'h143E: dout  = 8'b00000000; // 5182 :   0 - 0x0
      13'h143F: dout  = 8'b00000000; // 5183 :   0 - 0x0
      13'h1440: dout  = 8'b00000000; // 5184 :   0 - 0x0 -- Background 0x44
      13'h1441: dout  = 8'b00000000; // 5185 :   0 - 0x0
      13'h1442: dout  = 8'b00000000; // 5186 :   0 - 0x0
      13'h1443: dout  = 8'b00000000; // 5187 :   0 - 0x0
      13'h1444: dout  = 8'b00000000; // 5188 :   0 - 0x0
      13'h1445: dout  = 8'b00000000; // 5189 :   0 - 0x0
      13'h1446: dout  = 8'b00000000; // 5190 :   0 - 0x0
      13'h1447: dout  = 8'b00000000; // 5191 :   0 - 0x0
      13'h1448: dout  = 8'b00000000; // 5192 :   0 - 0x0
      13'h1449: dout  = 8'b00000000; // 5193 :   0 - 0x0
      13'h144A: dout  = 8'b00000000; // 5194 :   0 - 0x0
      13'h144B: dout  = 8'b00000000; // 5195 :   0 - 0x0
      13'h144C: dout  = 8'b00000000; // 5196 :   0 - 0x0
      13'h144D: dout  = 8'b00000000; // 5197 :   0 - 0x0
      13'h144E: dout  = 8'b00000000; // 5198 :   0 - 0x0
      13'h144F: dout  = 8'b00000000; // 5199 :   0 - 0x0
      13'h1450: dout  = 8'b00000000; // 5200 :   0 - 0x0 -- Background 0x45
      13'h1451: dout  = 8'b00000000; // 5201 :   0 - 0x0
      13'h1452: dout  = 8'b00000000; // 5202 :   0 - 0x0
      13'h1453: dout  = 8'b00000000; // 5203 :   0 - 0x0
      13'h1454: dout  = 8'b00000000; // 5204 :   0 - 0x0
      13'h1455: dout  = 8'b00000000; // 5205 :   0 - 0x0
      13'h1456: dout  = 8'b00000000; // 5206 :   0 - 0x0
      13'h1457: dout  = 8'b00000000; // 5207 :   0 - 0x0
      13'h1458: dout  = 8'b00000000; // 5208 :   0 - 0x0
      13'h1459: dout  = 8'b00000000; // 5209 :   0 - 0x0
      13'h145A: dout  = 8'b00000000; // 5210 :   0 - 0x0
      13'h145B: dout  = 8'b00000000; // 5211 :   0 - 0x0
      13'h145C: dout  = 8'b00000000; // 5212 :   0 - 0x0
      13'h145D: dout  = 8'b00000000; // 5213 :   0 - 0x0
      13'h145E: dout  = 8'b00000000; // 5214 :   0 - 0x0
      13'h145F: dout  = 8'b00000000; // 5215 :   0 - 0x0
      13'h1460: dout  = 8'b00000000; // 5216 :   0 - 0x0 -- Background 0x46
      13'h1461: dout  = 8'b00000000; // 5217 :   0 - 0x0
      13'h1462: dout  = 8'b00000000; // 5218 :   0 - 0x0
      13'h1463: dout  = 8'b00000000; // 5219 :   0 - 0x0
      13'h1464: dout  = 8'b00000000; // 5220 :   0 - 0x0
      13'h1465: dout  = 8'b00000000; // 5221 :   0 - 0x0
      13'h1466: dout  = 8'b00000000; // 5222 :   0 - 0x0
      13'h1467: dout  = 8'b00000000; // 5223 :   0 - 0x0
      13'h1468: dout  = 8'b00000000; // 5224 :   0 - 0x0
      13'h1469: dout  = 8'b00000000; // 5225 :   0 - 0x0
      13'h146A: dout  = 8'b00000000; // 5226 :   0 - 0x0
      13'h146B: dout  = 8'b00000000; // 5227 :   0 - 0x0
      13'h146C: dout  = 8'b00000000; // 5228 :   0 - 0x0
      13'h146D: dout  = 8'b00000000; // 5229 :   0 - 0x0
      13'h146E: dout  = 8'b00000000; // 5230 :   0 - 0x0
      13'h146F: dout  = 8'b00000000; // 5231 :   0 - 0x0
      13'h1470: dout  = 8'b00000000; // 5232 :   0 - 0x0 -- Background 0x47
      13'h1471: dout  = 8'b00000000; // 5233 :   0 - 0x0
      13'h1472: dout  = 8'b00000000; // 5234 :   0 - 0x0
      13'h1473: dout  = 8'b00000000; // 5235 :   0 - 0x0
      13'h1474: dout  = 8'b00000000; // 5236 :   0 - 0x0
      13'h1475: dout  = 8'b00000000; // 5237 :   0 - 0x0
      13'h1476: dout  = 8'b00000000; // 5238 :   0 - 0x0
      13'h1477: dout  = 8'b00000000; // 5239 :   0 - 0x0
      13'h1478: dout  = 8'b00000000; // 5240 :   0 - 0x0
      13'h1479: dout  = 8'b00000000; // 5241 :   0 - 0x0
      13'h147A: dout  = 8'b00000000; // 5242 :   0 - 0x0
      13'h147B: dout  = 8'b00000000; // 5243 :   0 - 0x0
      13'h147C: dout  = 8'b00000000; // 5244 :   0 - 0x0
      13'h147D: dout  = 8'b00000000; // 5245 :   0 - 0x0
      13'h147E: dout  = 8'b00000000; // 5246 :   0 - 0x0
      13'h147F: dout  = 8'b00000000; // 5247 :   0 - 0x0
      13'h1480: dout  = 8'b00000000; // 5248 :   0 - 0x0 -- Background 0x48
      13'h1481: dout  = 8'b00000000; // 5249 :   0 - 0x0
      13'h1482: dout  = 8'b00000000; // 5250 :   0 - 0x0
      13'h1483: dout  = 8'b00000000; // 5251 :   0 - 0x0
      13'h1484: dout  = 8'b00000000; // 5252 :   0 - 0x0
      13'h1485: dout  = 8'b00000000; // 5253 :   0 - 0x0
      13'h1486: dout  = 8'b00000000; // 5254 :   0 - 0x0
      13'h1487: dout  = 8'b00000000; // 5255 :   0 - 0x0
      13'h1488: dout  = 8'b00000000; // 5256 :   0 - 0x0
      13'h1489: dout  = 8'b00000000; // 5257 :   0 - 0x0
      13'h148A: dout  = 8'b00000000; // 5258 :   0 - 0x0
      13'h148B: dout  = 8'b00000000; // 5259 :   0 - 0x0
      13'h148C: dout  = 8'b00000000; // 5260 :   0 - 0x0
      13'h148D: dout  = 8'b00000000; // 5261 :   0 - 0x0
      13'h148E: dout  = 8'b00000000; // 5262 :   0 - 0x0
      13'h148F: dout  = 8'b00000000; // 5263 :   0 - 0x0
      13'h1490: dout  = 8'b00000000; // 5264 :   0 - 0x0 -- Background 0x49
      13'h1491: dout  = 8'b00000000; // 5265 :   0 - 0x0
      13'h1492: dout  = 8'b00000000; // 5266 :   0 - 0x0
      13'h1493: dout  = 8'b00000000; // 5267 :   0 - 0x0
      13'h1494: dout  = 8'b00000000; // 5268 :   0 - 0x0
      13'h1495: dout  = 8'b00000000; // 5269 :   0 - 0x0
      13'h1496: dout  = 8'b00000000; // 5270 :   0 - 0x0
      13'h1497: dout  = 8'b00000000; // 5271 :   0 - 0x0
      13'h1498: dout  = 8'b00000000; // 5272 :   0 - 0x0
      13'h1499: dout  = 8'b00000000; // 5273 :   0 - 0x0
      13'h149A: dout  = 8'b00000000; // 5274 :   0 - 0x0
      13'h149B: dout  = 8'b00000000; // 5275 :   0 - 0x0
      13'h149C: dout  = 8'b00000000; // 5276 :   0 - 0x0
      13'h149D: dout  = 8'b00000000; // 5277 :   0 - 0x0
      13'h149E: dout  = 8'b00000000; // 5278 :   0 - 0x0
      13'h149F: dout  = 8'b00000000; // 5279 :   0 - 0x0
      13'h14A0: dout  = 8'b00000000; // 5280 :   0 - 0x0 -- Background 0x4a
      13'h14A1: dout  = 8'b00000000; // 5281 :   0 - 0x0
      13'h14A2: dout  = 8'b00000000; // 5282 :   0 - 0x0
      13'h14A3: dout  = 8'b00000000; // 5283 :   0 - 0x0
      13'h14A4: dout  = 8'b00000000; // 5284 :   0 - 0x0
      13'h14A5: dout  = 8'b00000000; // 5285 :   0 - 0x0
      13'h14A6: dout  = 8'b00000000; // 5286 :   0 - 0x0
      13'h14A7: dout  = 8'b00000000; // 5287 :   0 - 0x0
      13'h14A8: dout  = 8'b00000000; // 5288 :   0 - 0x0
      13'h14A9: dout  = 8'b00000000; // 5289 :   0 - 0x0
      13'h14AA: dout  = 8'b00000000; // 5290 :   0 - 0x0
      13'h14AB: dout  = 8'b00000000; // 5291 :   0 - 0x0
      13'h14AC: dout  = 8'b00000000; // 5292 :   0 - 0x0
      13'h14AD: dout  = 8'b00000000; // 5293 :   0 - 0x0
      13'h14AE: dout  = 8'b00000000; // 5294 :   0 - 0x0
      13'h14AF: dout  = 8'b00000000; // 5295 :   0 - 0x0
      13'h14B0: dout  = 8'b00000000; // 5296 :   0 - 0x0 -- Background 0x4b
      13'h14B1: dout  = 8'b00000000; // 5297 :   0 - 0x0
      13'h14B2: dout  = 8'b00000000; // 5298 :   0 - 0x0
      13'h14B3: dout  = 8'b00000000; // 5299 :   0 - 0x0
      13'h14B4: dout  = 8'b00000000; // 5300 :   0 - 0x0
      13'h14B5: dout  = 8'b00000000; // 5301 :   0 - 0x0
      13'h14B6: dout  = 8'b00000000; // 5302 :   0 - 0x0
      13'h14B7: dout  = 8'b00000000; // 5303 :   0 - 0x0
      13'h14B8: dout  = 8'b00000000; // 5304 :   0 - 0x0
      13'h14B9: dout  = 8'b00000000; // 5305 :   0 - 0x0
      13'h14BA: dout  = 8'b00000000; // 5306 :   0 - 0x0
      13'h14BB: dout  = 8'b00000000; // 5307 :   0 - 0x0
      13'h14BC: dout  = 8'b00000000; // 5308 :   0 - 0x0
      13'h14BD: dout  = 8'b00000000; // 5309 :   0 - 0x0
      13'h14BE: dout  = 8'b00000000; // 5310 :   0 - 0x0
      13'h14BF: dout  = 8'b00000000; // 5311 :   0 - 0x0
      13'h14C0: dout  = 8'b00000000; // 5312 :   0 - 0x0 -- Background 0x4c
      13'h14C1: dout  = 8'b00000000; // 5313 :   0 - 0x0
      13'h14C2: dout  = 8'b00000000; // 5314 :   0 - 0x0
      13'h14C3: dout  = 8'b00000000; // 5315 :   0 - 0x0
      13'h14C4: dout  = 8'b00000000; // 5316 :   0 - 0x0
      13'h14C5: dout  = 8'b00000000; // 5317 :   0 - 0x0
      13'h14C6: dout  = 8'b00000000; // 5318 :   0 - 0x0
      13'h14C7: dout  = 8'b00000000; // 5319 :   0 - 0x0
      13'h14C8: dout  = 8'b00000000; // 5320 :   0 - 0x0
      13'h14C9: dout  = 8'b00000000; // 5321 :   0 - 0x0
      13'h14CA: dout  = 8'b00000000; // 5322 :   0 - 0x0
      13'h14CB: dout  = 8'b00000000; // 5323 :   0 - 0x0
      13'h14CC: dout  = 8'b00000000; // 5324 :   0 - 0x0
      13'h14CD: dout  = 8'b00000000; // 5325 :   0 - 0x0
      13'h14CE: dout  = 8'b00000000; // 5326 :   0 - 0x0
      13'h14CF: dout  = 8'b00000000; // 5327 :   0 - 0x0
      13'h14D0: dout  = 8'b00000000; // 5328 :   0 - 0x0 -- Background 0x4d
      13'h14D1: dout  = 8'b00000000; // 5329 :   0 - 0x0
      13'h14D2: dout  = 8'b00000000; // 5330 :   0 - 0x0
      13'h14D3: dout  = 8'b00000000; // 5331 :   0 - 0x0
      13'h14D4: dout  = 8'b00000000; // 5332 :   0 - 0x0
      13'h14D5: dout  = 8'b00000000; // 5333 :   0 - 0x0
      13'h14D6: dout  = 8'b00000000; // 5334 :   0 - 0x0
      13'h14D7: dout  = 8'b00000000; // 5335 :   0 - 0x0
      13'h14D8: dout  = 8'b00000000; // 5336 :   0 - 0x0
      13'h14D9: dout  = 8'b00000000; // 5337 :   0 - 0x0
      13'h14DA: dout  = 8'b00000000; // 5338 :   0 - 0x0
      13'h14DB: dout  = 8'b00000000; // 5339 :   0 - 0x0
      13'h14DC: dout  = 8'b00000000; // 5340 :   0 - 0x0
      13'h14DD: dout  = 8'b00000000; // 5341 :   0 - 0x0
      13'h14DE: dout  = 8'b00000000; // 5342 :   0 - 0x0
      13'h14DF: dout  = 8'b00000000; // 5343 :   0 - 0x0
      13'h14E0: dout  = 8'b00000000; // 5344 :   0 - 0x0 -- Background 0x4e
      13'h14E1: dout  = 8'b00000000; // 5345 :   0 - 0x0
      13'h14E2: dout  = 8'b00000000; // 5346 :   0 - 0x0
      13'h14E3: dout  = 8'b00000000; // 5347 :   0 - 0x0
      13'h14E4: dout  = 8'b00000000; // 5348 :   0 - 0x0
      13'h14E5: dout  = 8'b00000000; // 5349 :   0 - 0x0
      13'h14E6: dout  = 8'b00000000; // 5350 :   0 - 0x0
      13'h14E7: dout  = 8'b00000000; // 5351 :   0 - 0x0
      13'h14E8: dout  = 8'b00000000; // 5352 :   0 - 0x0
      13'h14E9: dout  = 8'b00000000; // 5353 :   0 - 0x0
      13'h14EA: dout  = 8'b00000000; // 5354 :   0 - 0x0
      13'h14EB: dout  = 8'b00000000; // 5355 :   0 - 0x0
      13'h14EC: dout  = 8'b00000000; // 5356 :   0 - 0x0
      13'h14ED: dout  = 8'b00000000; // 5357 :   0 - 0x0
      13'h14EE: dout  = 8'b00000000; // 5358 :   0 - 0x0
      13'h14EF: dout  = 8'b00000000; // 5359 :   0 - 0x0
      13'h14F0: dout  = 8'b00000000; // 5360 :   0 - 0x0 -- Background 0x4f
      13'h14F1: dout  = 8'b00000000; // 5361 :   0 - 0x0
      13'h14F2: dout  = 8'b00000000; // 5362 :   0 - 0x0
      13'h14F3: dout  = 8'b00000000; // 5363 :   0 - 0x0
      13'h14F4: dout  = 8'b00000000; // 5364 :   0 - 0x0
      13'h14F5: dout  = 8'b00000000; // 5365 :   0 - 0x0
      13'h14F6: dout  = 8'b00000000; // 5366 :   0 - 0x0
      13'h14F7: dout  = 8'b00000000; // 5367 :   0 - 0x0
      13'h14F8: dout  = 8'b00000000; // 5368 :   0 - 0x0
      13'h14F9: dout  = 8'b00000000; // 5369 :   0 - 0x0
      13'h14FA: dout  = 8'b00000000; // 5370 :   0 - 0x0
      13'h14FB: dout  = 8'b00000000; // 5371 :   0 - 0x0
      13'h14FC: dout  = 8'b00000000; // 5372 :   0 - 0x0
      13'h14FD: dout  = 8'b00000000; // 5373 :   0 - 0x0
      13'h14FE: dout  = 8'b00000000; // 5374 :   0 - 0x0
      13'h14FF: dout  = 8'b00000000; // 5375 :   0 - 0x0
      13'h1500: dout  = 8'b00000000; // 5376 :   0 - 0x0 -- Background 0x50
      13'h1501: dout  = 8'b00000000; // 5377 :   0 - 0x0
      13'h1502: dout  = 8'b00000000; // 5378 :   0 - 0x0
      13'h1503: dout  = 8'b00000000; // 5379 :   0 - 0x0
      13'h1504: dout  = 8'b00000000; // 5380 :   0 - 0x0
      13'h1505: dout  = 8'b00000000; // 5381 :   0 - 0x0
      13'h1506: dout  = 8'b00000000; // 5382 :   0 - 0x0
      13'h1507: dout  = 8'b00000000; // 5383 :   0 - 0x0
      13'h1508: dout  = 8'b00000000; // 5384 :   0 - 0x0
      13'h1509: dout  = 8'b00000000; // 5385 :   0 - 0x0
      13'h150A: dout  = 8'b00000000; // 5386 :   0 - 0x0
      13'h150B: dout  = 8'b00000000; // 5387 :   0 - 0x0
      13'h150C: dout  = 8'b00000000; // 5388 :   0 - 0x0
      13'h150D: dout  = 8'b00000000; // 5389 :   0 - 0x0
      13'h150E: dout  = 8'b00000000; // 5390 :   0 - 0x0
      13'h150F: dout  = 8'b00000000; // 5391 :   0 - 0x0
      13'h1510: dout  = 8'b00000000; // 5392 :   0 - 0x0 -- Background 0x51
      13'h1511: dout  = 8'b00000000; // 5393 :   0 - 0x0
      13'h1512: dout  = 8'b00000000; // 5394 :   0 - 0x0
      13'h1513: dout  = 8'b00000000; // 5395 :   0 - 0x0
      13'h1514: dout  = 8'b00000000; // 5396 :   0 - 0x0
      13'h1515: dout  = 8'b00000000; // 5397 :   0 - 0x0
      13'h1516: dout  = 8'b00000000; // 5398 :   0 - 0x0
      13'h1517: dout  = 8'b00000000; // 5399 :   0 - 0x0
      13'h1518: dout  = 8'b00000000; // 5400 :   0 - 0x0
      13'h1519: dout  = 8'b00000000; // 5401 :   0 - 0x0
      13'h151A: dout  = 8'b00000000; // 5402 :   0 - 0x0
      13'h151B: dout  = 8'b00000000; // 5403 :   0 - 0x0
      13'h151C: dout  = 8'b00000000; // 5404 :   0 - 0x0
      13'h151D: dout  = 8'b00000000; // 5405 :   0 - 0x0
      13'h151E: dout  = 8'b00000000; // 5406 :   0 - 0x0
      13'h151F: dout  = 8'b00000000; // 5407 :   0 - 0x0
      13'h1520: dout  = 8'b00000000; // 5408 :   0 - 0x0 -- Background 0x52
      13'h1521: dout  = 8'b00000000; // 5409 :   0 - 0x0
      13'h1522: dout  = 8'b00000000; // 5410 :   0 - 0x0
      13'h1523: dout  = 8'b00000000; // 5411 :   0 - 0x0
      13'h1524: dout  = 8'b00000000; // 5412 :   0 - 0x0
      13'h1525: dout  = 8'b00000000; // 5413 :   0 - 0x0
      13'h1526: dout  = 8'b00000000; // 5414 :   0 - 0x0
      13'h1527: dout  = 8'b00000000; // 5415 :   0 - 0x0
      13'h1528: dout  = 8'b00000000; // 5416 :   0 - 0x0
      13'h1529: dout  = 8'b00000000; // 5417 :   0 - 0x0
      13'h152A: dout  = 8'b00000000; // 5418 :   0 - 0x0
      13'h152B: dout  = 8'b00000000; // 5419 :   0 - 0x0
      13'h152C: dout  = 8'b00000000; // 5420 :   0 - 0x0
      13'h152D: dout  = 8'b00000000; // 5421 :   0 - 0x0
      13'h152E: dout  = 8'b00000000; // 5422 :   0 - 0x0
      13'h152F: dout  = 8'b00000000; // 5423 :   0 - 0x0
      13'h1530: dout  = 8'b00000000; // 5424 :   0 - 0x0 -- Background 0x53
      13'h1531: dout  = 8'b00000000; // 5425 :   0 - 0x0
      13'h1532: dout  = 8'b00000000; // 5426 :   0 - 0x0
      13'h1533: dout  = 8'b00000000; // 5427 :   0 - 0x0
      13'h1534: dout  = 8'b00000000; // 5428 :   0 - 0x0
      13'h1535: dout  = 8'b00000000; // 5429 :   0 - 0x0
      13'h1536: dout  = 8'b00000000; // 5430 :   0 - 0x0
      13'h1537: dout  = 8'b00000000; // 5431 :   0 - 0x0
      13'h1538: dout  = 8'b00000000; // 5432 :   0 - 0x0
      13'h1539: dout  = 8'b00000000; // 5433 :   0 - 0x0
      13'h153A: dout  = 8'b00000000; // 5434 :   0 - 0x0
      13'h153B: dout  = 8'b00000000; // 5435 :   0 - 0x0
      13'h153C: dout  = 8'b00000000; // 5436 :   0 - 0x0
      13'h153D: dout  = 8'b00000000; // 5437 :   0 - 0x0
      13'h153E: dout  = 8'b00000000; // 5438 :   0 - 0x0
      13'h153F: dout  = 8'b00000000; // 5439 :   0 - 0x0
      13'h1540: dout  = 8'b00000000; // 5440 :   0 - 0x0 -- Background 0x54
      13'h1541: dout  = 8'b00000000; // 5441 :   0 - 0x0
      13'h1542: dout  = 8'b00000000; // 5442 :   0 - 0x0
      13'h1543: dout  = 8'b00000000; // 5443 :   0 - 0x0
      13'h1544: dout  = 8'b00000000; // 5444 :   0 - 0x0
      13'h1545: dout  = 8'b00000000; // 5445 :   0 - 0x0
      13'h1546: dout  = 8'b00000000; // 5446 :   0 - 0x0
      13'h1547: dout  = 8'b00000000; // 5447 :   0 - 0x0
      13'h1548: dout  = 8'b00000000; // 5448 :   0 - 0x0
      13'h1549: dout  = 8'b00000000; // 5449 :   0 - 0x0
      13'h154A: dout  = 8'b00000000; // 5450 :   0 - 0x0
      13'h154B: dout  = 8'b00000000; // 5451 :   0 - 0x0
      13'h154C: dout  = 8'b00000000; // 5452 :   0 - 0x0
      13'h154D: dout  = 8'b00000000; // 5453 :   0 - 0x0
      13'h154E: dout  = 8'b00000000; // 5454 :   0 - 0x0
      13'h154F: dout  = 8'b00000000; // 5455 :   0 - 0x0
      13'h1550: dout  = 8'b00000000; // 5456 :   0 - 0x0 -- Background 0x55
      13'h1551: dout  = 8'b00000000; // 5457 :   0 - 0x0
      13'h1552: dout  = 8'b00000000; // 5458 :   0 - 0x0
      13'h1553: dout  = 8'b00000000; // 5459 :   0 - 0x0
      13'h1554: dout  = 8'b00000000; // 5460 :   0 - 0x0
      13'h1555: dout  = 8'b00000000; // 5461 :   0 - 0x0
      13'h1556: dout  = 8'b00000000; // 5462 :   0 - 0x0
      13'h1557: dout  = 8'b00000000; // 5463 :   0 - 0x0
      13'h1558: dout  = 8'b00000000; // 5464 :   0 - 0x0
      13'h1559: dout  = 8'b00000000; // 5465 :   0 - 0x0
      13'h155A: dout  = 8'b00000000; // 5466 :   0 - 0x0
      13'h155B: dout  = 8'b00000000; // 5467 :   0 - 0x0
      13'h155C: dout  = 8'b00000000; // 5468 :   0 - 0x0
      13'h155D: dout  = 8'b00000000; // 5469 :   0 - 0x0
      13'h155E: dout  = 8'b00000000; // 5470 :   0 - 0x0
      13'h155F: dout  = 8'b00000000; // 5471 :   0 - 0x0
      13'h1560: dout  = 8'b00000000; // 5472 :   0 - 0x0 -- Background 0x56
      13'h1561: dout  = 8'b00000000; // 5473 :   0 - 0x0
      13'h1562: dout  = 8'b00000000; // 5474 :   0 - 0x0
      13'h1563: dout  = 8'b00000000; // 5475 :   0 - 0x0
      13'h1564: dout  = 8'b00000000; // 5476 :   0 - 0x0
      13'h1565: dout  = 8'b00000000; // 5477 :   0 - 0x0
      13'h1566: dout  = 8'b00000000; // 5478 :   0 - 0x0
      13'h1567: dout  = 8'b00000000; // 5479 :   0 - 0x0
      13'h1568: dout  = 8'b00000000; // 5480 :   0 - 0x0
      13'h1569: dout  = 8'b00000000; // 5481 :   0 - 0x0
      13'h156A: dout  = 8'b00000000; // 5482 :   0 - 0x0
      13'h156B: dout  = 8'b00000000; // 5483 :   0 - 0x0
      13'h156C: dout  = 8'b00000000; // 5484 :   0 - 0x0
      13'h156D: dout  = 8'b00000000; // 5485 :   0 - 0x0
      13'h156E: dout  = 8'b00000000; // 5486 :   0 - 0x0
      13'h156F: dout  = 8'b00000000; // 5487 :   0 - 0x0
      13'h1570: dout  = 8'b00000000; // 5488 :   0 - 0x0 -- Background 0x57
      13'h1571: dout  = 8'b00000000; // 5489 :   0 - 0x0
      13'h1572: dout  = 8'b00000000; // 5490 :   0 - 0x0
      13'h1573: dout  = 8'b00000000; // 5491 :   0 - 0x0
      13'h1574: dout  = 8'b00000000; // 5492 :   0 - 0x0
      13'h1575: dout  = 8'b00000000; // 5493 :   0 - 0x0
      13'h1576: dout  = 8'b00000000; // 5494 :   0 - 0x0
      13'h1577: dout  = 8'b00000000; // 5495 :   0 - 0x0
      13'h1578: dout  = 8'b00000000; // 5496 :   0 - 0x0
      13'h1579: dout  = 8'b00000000; // 5497 :   0 - 0x0
      13'h157A: dout  = 8'b00000000; // 5498 :   0 - 0x0
      13'h157B: dout  = 8'b00000000; // 5499 :   0 - 0x0
      13'h157C: dout  = 8'b00000000; // 5500 :   0 - 0x0
      13'h157D: dout  = 8'b00000000; // 5501 :   0 - 0x0
      13'h157E: dout  = 8'b00000000; // 5502 :   0 - 0x0
      13'h157F: dout  = 8'b00000000; // 5503 :   0 - 0x0
      13'h1580: dout  = 8'b00000000; // 5504 :   0 - 0x0 -- Background 0x58
      13'h1581: dout  = 8'b00000000; // 5505 :   0 - 0x0
      13'h1582: dout  = 8'b00000000; // 5506 :   0 - 0x0
      13'h1583: dout  = 8'b00000000; // 5507 :   0 - 0x0
      13'h1584: dout  = 8'b00000000; // 5508 :   0 - 0x0
      13'h1585: dout  = 8'b00000000; // 5509 :   0 - 0x0
      13'h1586: dout  = 8'b00000000; // 5510 :   0 - 0x0
      13'h1587: dout  = 8'b00000000; // 5511 :   0 - 0x0
      13'h1588: dout  = 8'b00000000; // 5512 :   0 - 0x0
      13'h1589: dout  = 8'b00000000; // 5513 :   0 - 0x0
      13'h158A: dout  = 8'b00000000; // 5514 :   0 - 0x0
      13'h158B: dout  = 8'b00000000; // 5515 :   0 - 0x0
      13'h158C: dout  = 8'b00000000; // 5516 :   0 - 0x0
      13'h158D: dout  = 8'b00000000; // 5517 :   0 - 0x0
      13'h158E: dout  = 8'b00000000; // 5518 :   0 - 0x0
      13'h158F: dout  = 8'b00000000; // 5519 :   0 - 0x0
      13'h1590: dout  = 8'b00000000; // 5520 :   0 - 0x0 -- Background 0x59
      13'h1591: dout  = 8'b00000000; // 5521 :   0 - 0x0
      13'h1592: dout  = 8'b00000000; // 5522 :   0 - 0x0
      13'h1593: dout  = 8'b00000000; // 5523 :   0 - 0x0
      13'h1594: dout  = 8'b00000000; // 5524 :   0 - 0x0
      13'h1595: dout  = 8'b00000000; // 5525 :   0 - 0x0
      13'h1596: dout  = 8'b00000000; // 5526 :   0 - 0x0
      13'h1597: dout  = 8'b00000000; // 5527 :   0 - 0x0
      13'h1598: dout  = 8'b00000000; // 5528 :   0 - 0x0
      13'h1599: dout  = 8'b00000000; // 5529 :   0 - 0x0
      13'h159A: dout  = 8'b00000000; // 5530 :   0 - 0x0
      13'h159B: dout  = 8'b00000000; // 5531 :   0 - 0x0
      13'h159C: dout  = 8'b00000000; // 5532 :   0 - 0x0
      13'h159D: dout  = 8'b00000000; // 5533 :   0 - 0x0
      13'h159E: dout  = 8'b00000000; // 5534 :   0 - 0x0
      13'h159F: dout  = 8'b00000000; // 5535 :   0 - 0x0
      13'h15A0: dout  = 8'b00000000; // 5536 :   0 - 0x0 -- Background 0x5a
      13'h15A1: dout  = 8'b00000000; // 5537 :   0 - 0x0
      13'h15A2: dout  = 8'b00000000; // 5538 :   0 - 0x0
      13'h15A3: dout  = 8'b00000000; // 5539 :   0 - 0x0
      13'h15A4: dout  = 8'b00000000; // 5540 :   0 - 0x0
      13'h15A5: dout  = 8'b00000000; // 5541 :   0 - 0x0
      13'h15A6: dout  = 8'b00000000; // 5542 :   0 - 0x0
      13'h15A7: dout  = 8'b00000000; // 5543 :   0 - 0x0
      13'h15A8: dout  = 8'b00000000; // 5544 :   0 - 0x0
      13'h15A9: dout  = 8'b00000000; // 5545 :   0 - 0x0
      13'h15AA: dout  = 8'b00000000; // 5546 :   0 - 0x0
      13'h15AB: dout  = 8'b00000000; // 5547 :   0 - 0x0
      13'h15AC: dout  = 8'b00000000; // 5548 :   0 - 0x0
      13'h15AD: dout  = 8'b00000000; // 5549 :   0 - 0x0
      13'h15AE: dout  = 8'b00000000; // 5550 :   0 - 0x0
      13'h15AF: dout  = 8'b00000000; // 5551 :   0 - 0x0
      13'h15B0: dout  = 8'b00000000; // 5552 :   0 - 0x0 -- Background 0x5b
      13'h15B1: dout  = 8'b00000000; // 5553 :   0 - 0x0
      13'h15B2: dout  = 8'b00000000; // 5554 :   0 - 0x0
      13'h15B3: dout  = 8'b00000000; // 5555 :   0 - 0x0
      13'h15B4: dout  = 8'b00000000; // 5556 :   0 - 0x0
      13'h15B5: dout  = 8'b00000000; // 5557 :   0 - 0x0
      13'h15B6: dout  = 8'b00000000; // 5558 :   0 - 0x0
      13'h15B7: dout  = 8'b00000000; // 5559 :   0 - 0x0
      13'h15B8: dout  = 8'b00000000; // 5560 :   0 - 0x0
      13'h15B9: dout  = 8'b00000000; // 5561 :   0 - 0x0
      13'h15BA: dout  = 8'b00000000; // 5562 :   0 - 0x0
      13'h15BB: dout  = 8'b00000000; // 5563 :   0 - 0x0
      13'h15BC: dout  = 8'b00000000; // 5564 :   0 - 0x0
      13'h15BD: dout  = 8'b00000000; // 5565 :   0 - 0x0
      13'h15BE: dout  = 8'b00000000; // 5566 :   0 - 0x0
      13'h15BF: dout  = 8'b00000000; // 5567 :   0 - 0x0
      13'h15C0: dout  = 8'b00000000; // 5568 :   0 - 0x0 -- Background 0x5c
      13'h15C1: dout  = 8'b00000000; // 5569 :   0 - 0x0
      13'h15C2: dout  = 8'b00000000; // 5570 :   0 - 0x0
      13'h15C3: dout  = 8'b00000000; // 5571 :   0 - 0x0
      13'h15C4: dout  = 8'b00000000; // 5572 :   0 - 0x0
      13'h15C5: dout  = 8'b00000000; // 5573 :   0 - 0x0
      13'h15C6: dout  = 8'b00000000; // 5574 :   0 - 0x0
      13'h15C7: dout  = 8'b00000000; // 5575 :   0 - 0x0
      13'h15C8: dout  = 8'b00000000; // 5576 :   0 - 0x0
      13'h15C9: dout  = 8'b00000000; // 5577 :   0 - 0x0
      13'h15CA: dout  = 8'b00000000; // 5578 :   0 - 0x0
      13'h15CB: dout  = 8'b00000000; // 5579 :   0 - 0x0
      13'h15CC: dout  = 8'b00000000; // 5580 :   0 - 0x0
      13'h15CD: dout  = 8'b00000000; // 5581 :   0 - 0x0
      13'h15CE: dout  = 8'b00000000; // 5582 :   0 - 0x0
      13'h15CF: dout  = 8'b00000000; // 5583 :   0 - 0x0
      13'h15D0: dout  = 8'b00000000; // 5584 :   0 - 0x0 -- Background 0x5d
      13'h15D1: dout  = 8'b00000000; // 5585 :   0 - 0x0
      13'h15D2: dout  = 8'b00000000; // 5586 :   0 - 0x0
      13'h15D3: dout  = 8'b00000000; // 5587 :   0 - 0x0
      13'h15D4: dout  = 8'b00000000; // 5588 :   0 - 0x0
      13'h15D5: dout  = 8'b00000000; // 5589 :   0 - 0x0
      13'h15D6: dout  = 8'b00000000; // 5590 :   0 - 0x0
      13'h15D7: dout  = 8'b00000000; // 5591 :   0 - 0x0
      13'h15D8: dout  = 8'b00000000; // 5592 :   0 - 0x0
      13'h15D9: dout  = 8'b00000000; // 5593 :   0 - 0x0
      13'h15DA: dout  = 8'b00000000; // 5594 :   0 - 0x0
      13'h15DB: dout  = 8'b00000000; // 5595 :   0 - 0x0
      13'h15DC: dout  = 8'b00000000; // 5596 :   0 - 0x0
      13'h15DD: dout  = 8'b00000000; // 5597 :   0 - 0x0
      13'h15DE: dout  = 8'b00000000; // 5598 :   0 - 0x0
      13'h15DF: dout  = 8'b00000000; // 5599 :   0 - 0x0
      13'h15E0: dout  = 8'b00000000; // 5600 :   0 - 0x0 -- Background 0x5e
      13'h15E1: dout  = 8'b00000000; // 5601 :   0 - 0x0
      13'h15E2: dout  = 8'b00000000; // 5602 :   0 - 0x0
      13'h15E3: dout  = 8'b00000000; // 5603 :   0 - 0x0
      13'h15E4: dout  = 8'b00000000; // 5604 :   0 - 0x0
      13'h15E5: dout  = 8'b00000000; // 5605 :   0 - 0x0
      13'h15E6: dout  = 8'b00000000; // 5606 :   0 - 0x0
      13'h15E7: dout  = 8'b00000000; // 5607 :   0 - 0x0
      13'h15E8: dout  = 8'b00000000; // 5608 :   0 - 0x0
      13'h15E9: dout  = 8'b00000000; // 5609 :   0 - 0x0
      13'h15EA: dout  = 8'b00000000; // 5610 :   0 - 0x0
      13'h15EB: dout  = 8'b00000000; // 5611 :   0 - 0x0
      13'h15EC: dout  = 8'b00000000; // 5612 :   0 - 0x0
      13'h15ED: dout  = 8'b00000000; // 5613 :   0 - 0x0
      13'h15EE: dout  = 8'b00000000; // 5614 :   0 - 0x0
      13'h15EF: dout  = 8'b00000000; // 5615 :   0 - 0x0
      13'h15F0: dout  = 8'b00000000; // 5616 :   0 - 0x0 -- Background 0x5f
      13'h15F1: dout  = 8'b00000000; // 5617 :   0 - 0x0
      13'h15F2: dout  = 8'b00000000; // 5618 :   0 - 0x0
      13'h15F3: dout  = 8'b00000000; // 5619 :   0 - 0x0
      13'h15F4: dout  = 8'b00000000; // 5620 :   0 - 0x0
      13'h15F5: dout  = 8'b00000000; // 5621 :   0 - 0x0
      13'h15F6: dout  = 8'b00000000; // 5622 :   0 - 0x0
      13'h15F7: dout  = 8'b00000000; // 5623 :   0 - 0x0
      13'h15F8: dout  = 8'b00000000; // 5624 :   0 - 0x0
      13'h15F9: dout  = 8'b00000000; // 5625 :   0 - 0x0
      13'h15FA: dout  = 8'b00000000; // 5626 :   0 - 0x0
      13'h15FB: dout  = 8'b00000000; // 5627 :   0 - 0x0
      13'h15FC: dout  = 8'b00000000; // 5628 :   0 - 0x0
      13'h15FD: dout  = 8'b00000000; // 5629 :   0 - 0x0
      13'h15FE: dout  = 8'b00000000; // 5630 :   0 - 0x0
      13'h15FF: dout  = 8'b00000000; // 5631 :   0 - 0x0
      13'h1600: dout  = 8'b00000000; // 5632 :   0 - 0x0 -- Background 0x60
      13'h1601: dout  = 8'b00000000; // 5633 :   0 - 0x0
      13'h1602: dout  = 8'b00000000; // 5634 :   0 - 0x0
      13'h1603: dout  = 8'b00000000; // 5635 :   0 - 0x0
      13'h1604: dout  = 8'b00000000; // 5636 :   0 - 0x0
      13'h1605: dout  = 8'b00000000; // 5637 :   0 - 0x0
      13'h1606: dout  = 8'b00000000; // 5638 :   0 - 0x0
      13'h1607: dout  = 8'b00000000; // 5639 :   0 - 0x0
      13'h1608: dout  = 8'b00000000; // 5640 :   0 - 0x0
      13'h1609: dout  = 8'b00000000; // 5641 :   0 - 0x0
      13'h160A: dout  = 8'b00000000; // 5642 :   0 - 0x0
      13'h160B: dout  = 8'b00000000; // 5643 :   0 - 0x0
      13'h160C: dout  = 8'b00000000; // 5644 :   0 - 0x0
      13'h160D: dout  = 8'b00000000; // 5645 :   0 - 0x0
      13'h160E: dout  = 8'b00000000; // 5646 :   0 - 0x0
      13'h160F: dout  = 8'b00000000; // 5647 :   0 - 0x0
      13'h1610: dout  = 8'b00000000; // 5648 :   0 - 0x0 -- Background 0x61
      13'h1611: dout  = 8'b00000000; // 5649 :   0 - 0x0
      13'h1612: dout  = 8'b00000000; // 5650 :   0 - 0x0
      13'h1613: dout  = 8'b00000000; // 5651 :   0 - 0x0
      13'h1614: dout  = 8'b00000000; // 5652 :   0 - 0x0
      13'h1615: dout  = 8'b00000000; // 5653 :   0 - 0x0
      13'h1616: dout  = 8'b00000000; // 5654 :   0 - 0x0
      13'h1617: dout  = 8'b00000000; // 5655 :   0 - 0x0
      13'h1618: dout  = 8'b00000000; // 5656 :   0 - 0x0
      13'h1619: dout  = 8'b00000000; // 5657 :   0 - 0x0
      13'h161A: dout  = 8'b00000000; // 5658 :   0 - 0x0
      13'h161B: dout  = 8'b00000000; // 5659 :   0 - 0x0
      13'h161C: dout  = 8'b00000000; // 5660 :   0 - 0x0
      13'h161D: dout  = 8'b00000000; // 5661 :   0 - 0x0
      13'h161E: dout  = 8'b00000000; // 5662 :   0 - 0x0
      13'h161F: dout  = 8'b00000000; // 5663 :   0 - 0x0
      13'h1620: dout  = 8'b00000000; // 5664 :   0 - 0x0 -- Background 0x62
      13'h1621: dout  = 8'b00000000; // 5665 :   0 - 0x0
      13'h1622: dout  = 8'b00000000; // 5666 :   0 - 0x0
      13'h1623: dout  = 8'b00000000; // 5667 :   0 - 0x0
      13'h1624: dout  = 8'b00000000; // 5668 :   0 - 0x0
      13'h1625: dout  = 8'b00000000; // 5669 :   0 - 0x0
      13'h1626: dout  = 8'b00000000; // 5670 :   0 - 0x0
      13'h1627: dout  = 8'b00000000; // 5671 :   0 - 0x0
      13'h1628: dout  = 8'b00000000; // 5672 :   0 - 0x0
      13'h1629: dout  = 8'b00000000; // 5673 :   0 - 0x0
      13'h162A: dout  = 8'b00000000; // 5674 :   0 - 0x0
      13'h162B: dout  = 8'b00000000; // 5675 :   0 - 0x0
      13'h162C: dout  = 8'b00000000; // 5676 :   0 - 0x0
      13'h162D: dout  = 8'b00000000; // 5677 :   0 - 0x0
      13'h162E: dout  = 8'b00000000; // 5678 :   0 - 0x0
      13'h162F: dout  = 8'b00000000; // 5679 :   0 - 0x0
      13'h1630: dout  = 8'b00000000; // 5680 :   0 - 0x0 -- Background 0x63
      13'h1631: dout  = 8'b00000000; // 5681 :   0 - 0x0
      13'h1632: dout  = 8'b00000000; // 5682 :   0 - 0x0
      13'h1633: dout  = 8'b00000000; // 5683 :   0 - 0x0
      13'h1634: dout  = 8'b00000000; // 5684 :   0 - 0x0
      13'h1635: dout  = 8'b00000000; // 5685 :   0 - 0x0
      13'h1636: dout  = 8'b00000000; // 5686 :   0 - 0x0
      13'h1637: dout  = 8'b00000000; // 5687 :   0 - 0x0
      13'h1638: dout  = 8'b00000000; // 5688 :   0 - 0x0
      13'h1639: dout  = 8'b00000000; // 5689 :   0 - 0x0
      13'h163A: dout  = 8'b00000000; // 5690 :   0 - 0x0
      13'h163B: dout  = 8'b00000000; // 5691 :   0 - 0x0
      13'h163C: dout  = 8'b00000000; // 5692 :   0 - 0x0
      13'h163D: dout  = 8'b00000000; // 5693 :   0 - 0x0
      13'h163E: dout  = 8'b00000000; // 5694 :   0 - 0x0
      13'h163F: dout  = 8'b00000000; // 5695 :   0 - 0x0
      13'h1640: dout  = 8'b00000000; // 5696 :   0 - 0x0 -- Background 0x64
      13'h1641: dout  = 8'b00000000; // 5697 :   0 - 0x0
      13'h1642: dout  = 8'b00000000; // 5698 :   0 - 0x0
      13'h1643: dout  = 8'b00000000; // 5699 :   0 - 0x0
      13'h1644: dout  = 8'b00000000; // 5700 :   0 - 0x0
      13'h1645: dout  = 8'b00000000; // 5701 :   0 - 0x0
      13'h1646: dout  = 8'b00000000; // 5702 :   0 - 0x0
      13'h1647: dout  = 8'b00000000; // 5703 :   0 - 0x0
      13'h1648: dout  = 8'b00000000; // 5704 :   0 - 0x0
      13'h1649: dout  = 8'b00000000; // 5705 :   0 - 0x0
      13'h164A: dout  = 8'b00000000; // 5706 :   0 - 0x0
      13'h164B: dout  = 8'b00000000; // 5707 :   0 - 0x0
      13'h164C: dout  = 8'b00000000; // 5708 :   0 - 0x0
      13'h164D: dout  = 8'b00000000; // 5709 :   0 - 0x0
      13'h164E: dout  = 8'b00000000; // 5710 :   0 - 0x0
      13'h164F: dout  = 8'b00000000; // 5711 :   0 - 0x0
      13'h1650: dout  = 8'b00000000; // 5712 :   0 - 0x0 -- Background 0x65
      13'h1651: dout  = 8'b00000000; // 5713 :   0 - 0x0
      13'h1652: dout  = 8'b00000000; // 5714 :   0 - 0x0
      13'h1653: dout  = 8'b00000000; // 5715 :   0 - 0x0
      13'h1654: dout  = 8'b00000000; // 5716 :   0 - 0x0
      13'h1655: dout  = 8'b00000000; // 5717 :   0 - 0x0
      13'h1656: dout  = 8'b00000000; // 5718 :   0 - 0x0
      13'h1657: dout  = 8'b00000000; // 5719 :   0 - 0x0
      13'h1658: dout  = 8'b00000000; // 5720 :   0 - 0x0
      13'h1659: dout  = 8'b00000000; // 5721 :   0 - 0x0
      13'h165A: dout  = 8'b00000000; // 5722 :   0 - 0x0
      13'h165B: dout  = 8'b00000000; // 5723 :   0 - 0x0
      13'h165C: dout  = 8'b00000000; // 5724 :   0 - 0x0
      13'h165D: dout  = 8'b00000000; // 5725 :   0 - 0x0
      13'h165E: dout  = 8'b00000000; // 5726 :   0 - 0x0
      13'h165F: dout  = 8'b00000000; // 5727 :   0 - 0x0
      13'h1660: dout  = 8'b00000000; // 5728 :   0 - 0x0 -- Background 0x66
      13'h1661: dout  = 8'b00000000; // 5729 :   0 - 0x0
      13'h1662: dout  = 8'b00000000; // 5730 :   0 - 0x0
      13'h1663: dout  = 8'b00000000; // 5731 :   0 - 0x0
      13'h1664: dout  = 8'b00000000; // 5732 :   0 - 0x0
      13'h1665: dout  = 8'b00000000; // 5733 :   0 - 0x0
      13'h1666: dout  = 8'b00000000; // 5734 :   0 - 0x0
      13'h1667: dout  = 8'b00000000; // 5735 :   0 - 0x0
      13'h1668: dout  = 8'b00000000; // 5736 :   0 - 0x0
      13'h1669: dout  = 8'b00000000; // 5737 :   0 - 0x0
      13'h166A: dout  = 8'b00000000; // 5738 :   0 - 0x0
      13'h166B: dout  = 8'b00000000; // 5739 :   0 - 0x0
      13'h166C: dout  = 8'b00000000; // 5740 :   0 - 0x0
      13'h166D: dout  = 8'b00000000; // 5741 :   0 - 0x0
      13'h166E: dout  = 8'b00000000; // 5742 :   0 - 0x0
      13'h166F: dout  = 8'b00000000; // 5743 :   0 - 0x0
      13'h1670: dout  = 8'b00000000; // 5744 :   0 - 0x0 -- Background 0x67
      13'h1671: dout  = 8'b00000000; // 5745 :   0 - 0x0
      13'h1672: dout  = 8'b00000000; // 5746 :   0 - 0x0
      13'h1673: dout  = 8'b00000000; // 5747 :   0 - 0x0
      13'h1674: dout  = 8'b00000000; // 5748 :   0 - 0x0
      13'h1675: dout  = 8'b00000000; // 5749 :   0 - 0x0
      13'h1676: dout  = 8'b00000000; // 5750 :   0 - 0x0
      13'h1677: dout  = 8'b00000000; // 5751 :   0 - 0x0
      13'h1678: dout  = 8'b00000000; // 5752 :   0 - 0x0
      13'h1679: dout  = 8'b00000000; // 5753 :   0 - 0x0
      13'h167A: dout  = 8'b00000000; // 5754 :   0 - 0x0
      13'h167B: dout  = 8'b00000000; // 5755 :   0 - 0x0
      13'h167C: dout  = 8'b00000000; // 5756 :   0 - 0x0
      13'h167D: dout  = 8'b00000000; // 5757 :   0 - 0x0
      13'h167E: dout  = 8'b00000000; // 5758 :   0 - 0x0
      13'h167F: dout  = 8'b00000000; // 5759 :   0 - 0x0
      13'h1680: dout  = 8'b00000000; // 5760 :   0 - 0x0 -- Background 0x68
      13'h1681: dout  = 8'b00000000; // 5761 :   0 - 0x0
      13'h1682: dout  = 8'b00000000; // 5762 :   0 - 0x0
      13'h1683: dout  = 8'b00000000; // 5763 :   0 - 0x0
      13'h1684: dout  = 8'b00000000; // 5764 :   0 - 0x0
      13'h1685: dout  = 8'b00000000; // 5765 :   0 - 0x0
      13'h1686: dout  = 8'b00000000; // 5766 :   0 - 0x0
      13'h1687: dout  = 8'b00000000; // 5767 :   0 - 0x0
      13'h1688: dout  = 8'b00000000; // 5768 :   0 - 0x0
      13'h1689: dout  = 8'b00000000; // 5769 :   0 - 0x0
      13'h168A: dout  = 8'b00000000; // 5770 :   0 - 0x0
      13'h168B: dout  = 8'b00000000; // 5771 :   0 - 0x0
      13'h168C: dout  = 8'b00000000; // 5772 :   0 - 0x0
      13'h168D: dout  = 8'b00000000; // 5773 :   0 - 0x0
      13'h168E: dout  = 8'b00000000; // 5774 :   0 - 0x0
      13'h168F: dout  = 8'b00000000; // 5775 :   0 - 0x0
      13'h1690: dout  = 8'b00000000; // 5776 :   0 - 0x0 -- Background 0x69
      13'h1691: dout  = 8'b00000000; // 5777 :   0 - 0x0
      13'h1692: dout  = 8'b00000000; // 5778 :   0 - 0x0
      13'h1693: dout  = 8'b00000000; // 5779 :   0 - 0x0
      13'h1694: dout  = 8'b00000000; // 5780 :   0 - 0x0
      13'h1695: dout  = 8'b00000000; // 5781 :   0 - 0x0
      13'h1696: dout  = 8'b00000000; // 5782 :   0 - 0x0
      13'h1697: dout  = 8'b00000000; // 5783 :   0 - 0x0
      13'h1698: dout  = 8'b00000000; // 5784 :   0 - 0x0
      13'h1699: dout  = 8'b00000000; // 5785 :   0 - 0x0
      13'h169A: dout  = 8'b00000000; // 5786 :   0 - 0x0
      13'h169B: dout  = 8'b00000000; // 5787 :   0 - 0x0
      13'h169C: dout  = 8'b00000000; // 5788 :   0 - 0x0
      13'h169D: dout  = 8'b00000000; // 5789 :   0 - 0x0
      13'h169E: dout  = 8'b00000000; // 5790 :   0 - 0x0
      13'h169F: dout  = 8'b00000000; // 5791 :   0 - 0x0
      13'h16A0: dout  = 8'b00000000; // 5792 :   0 - 0x0 -- Background 0x6a
      13'h16A1: dout  = 8'b00000000; // 5793 :   0 - 0x0
      13'h16A2: dout  = 8'b00000000; // 5794 :   0 - 0x0
      13'h16A3: dout  = 8'b00000000; // 5795 :   0 - 0x0
      13'h16A4: dout  = 8'b00000000; // 5796 :   0 - 0x0
      13'h16A5: dout  = 8'b00000000; // 5797 :   0 - 0x0
      13'h16A6: dout  = 8'b00000000; // 5798 :   0 - 0x0
      13'h16A7: dout  = 8'b00000000; // 5799 :   0 - 0x0
      13'h16A8: dout  = 8'b00000000; // 5800 :   0 - 0x0
      13'h16A9: dout  = 8'b00000000; // 5801 :   0 - 0x0
      13'h16AA: dout  = 8'b00000000; // 5802 :   0 - 0x0
      13'h16AB: dout  = 8'b00000000; // 5803 :   0 - 0x0
      13'h16AC: dout  = 8'b00000000; // 5804 :   0 - 0x0
      13'h16AD: dout  = 8'b00000000; // 5805 :   0 - 0x0
      13'h16AE: dout  = 8'b00000000; // 5806 :   0 - 0x0
      13'h16AF: dout  = 8'b00000000; // 5807 :   0 - 0x0
      13'h16B0: dout  = 8'b00000000; // 5808 :   0 - 0x0 -- Background 0x6b
      13'h16B1: dout  = 8'b00000000; // 5809 :   0 - 0x0
      13'h16B2: dout  = 8'b00000000; // 5810 :   0 - 0x0
      13'h16B3: dout  = 8'b00000000; // 5811 :   0 - 0x0
      13'h16B4: dout  = 8'b00000000; // 5812 :   0 - 0x0
      13'h16B5: dout  = 8'b00000000; // 5813 :   0 - 0x0
      13'h16B6: dout  = 8'b00000000; // 5814 :   0 - 0x0
      13'h16B7: dout  = 8'b00000000; // 5815 :   0 - 0x0
      13'h16B8: dout  = 8'b00000000; // 5816 :   0 - 0x0
      13'h16B9: dout  = 8'b00000000; // 5817 :   0 - 0x0
      13'h16BA: dout  = 8'b00000000; // 5818 :   0 - 0x0
      13'h16BB: dout  = 8'b00000000; // 5819 :   0 - 0x0
      13'h16BC: dout  = 8'b00000000; // 5820 :   0 - 0x0
      13'h16BD: dout  = 8'b00000000; // 5821 :   0 - 0x0
      13'h16BE: dout  = 8'b00000000; // 5822 :   0 - 0x0
      13'h16BF: dout  = 8'b00000000; // 5823 :   0 - 0x0
      13'h16C0: dout  = 8'b00000000; // 5824 :   0 - 0x0 -- Background 0x6c
      13'h16C1: dout  = 8'b00000000; // 5825 :   0 - 0x0
      13'h16C2: dout  = 8'b00000000; // 5826 :   0 - 0x0
      13'h16C3: dout  = 8'b00000000; // 5827 :   0 - 0x0
      13'h16C4: dout  = 8'b00000000; // 5828 :   0 - 0x0
      13'h16C5: dout  = 8'b00000000; // 5829 :   0 - 0x0
      13'h16C6: dout  = 8'b00000000; // 5830 :   0 - 0x0
      13'h16C7: dout  = 8'b00000000; // 5831 :   0 - 0x0
      13'h16C8: dout  = 8'b00000000; // 5832 :   0 - 0x0
      13'h16C9: dout  = 8'b00000000; // 5833 :   0 - 0x0
      13'h16CA: dout  = 8'b00000000; // 5834 :   0 - 0x0
      13'h16CB: dout  = 8'b00000000; // 5835 :   0 - 0x0
      13'h16CC: dout  = 8'b00000000; // 5836 :   0 - 0x0
      13'h16CD: dout  = 8'b00000000; // 5837 :   0 - 0x0
      13'h16CE: dout  = 8'b00000000; // 5838 :   0 - 0x0
      13'h16CF: dout  = 8'b00000000; // 5839 :   0 - 0x0
      13'h16D0: dout  = 8'b00000000; // 5840 :   0 - 0x0 -- Background 0x6d
      13'h16D1: dout  = 8'b00000000; // 5841 :   0 - 0x0
      13'h16D2: dout  = 8'b00000000; // 5842 :   0 - 0x0
      13'h16D3: dout  = 8'b00000000; // 5843 :   0 - 0x0
      13'h16D4: dout  = 8'b00000000; // 5844 :   0 - 0x0
      13'h16D5: dout  = 8'b00000000; // 5845 :   0 - 0x0
      13'h16D6: dout  = 8'b00000000; // 5846 :   0 - 0x0
      13'h16D7: dout  = 8'b00000000; // 5847 :   0 - 0x0
      13'h16D8: dout  = 8'b00000000; // 5848 :   0 - 0x0
      13'h16D9: dout  = 8'b00000000; // 5849 :   0 - 0x0
      13'h16DA: dout  = 8'b00000000; // 5850 :   0 - 0x0
      13'h16DB: dout  = 8'b00000000; // 5851 :   0 - 0x0
      13'h16DC: dout  = 8'b00000000; // 5852 :   0 - 0x0
      13'h16DD: dout  = 8'b00000000; // 5853 :   0 - 0x0
      13'h16DE: dout  = 8'b00000000; // 5854 :   0 - 0x0
      13'h16DF: dout  = 8'b00000000; // 5855 :   0 - 0x0
      13'h16E0: dout  = 8'b00000000; // 5856 :   0 - 0x0 -- Background 0x6e
      13'h16E1: dout  = 8'b00000000; // 5857 :   0 - 0x0
      13'h16E2: dout  = 8'b00000000; // 5858 :   0 - 0x0
      13'h16E3: dout  = 8'b00000000; // 5859 :   0 - 0x0
      13'h16E4: dout  = 8'b00000000; // 5860 :   0 - 0x0
      13'h16E5: dout  = 8'b00000000; // 5861 :   0 - 0x0
      13'h16E6: dout  = 8'b00000000; // 5862 :   0 - 0x0
      13'h16E7: dout  = 8'b00000000; // 5863 :   0 - 0x0
      13'h16E8: dout  = 8'b00000000; // 5864 :   0 - 0x0
      13'h16E9: dout  = 8'b00000000; // 5865 :   0 - 0x0
      13'h16EA: dout  = 8'b00000000; // 5866 :   0 - 0x0
      13'h16EB: dout  = 8'b00000000; // 5867 :   0 - 0x0
      13'h16EC: dout  = 8'b00000000; // 5868 :   0 - 0x0
      13'h16ED: dout  = 8'b00000000; // 5869 :   0 - 0x0
      13'h16EE: dout  = 8'b00000000; // 5870 :   0 - 0x0
      13'h16EF: dout  = 8'b00000000; // 5871 :   0 - 0x0
      13'h16F0: dout  = 8'b00000000; // 5872 :   0 - 0x0 -- Background 0x6f
      13'h16F1: dout  = 8'b00000000; // 5873 :   0 - 0x0
      13'h16F2: dout  = 8'b00000000; // 5874 :   0 - 0x0
      13'h16F3: dout  = 8'b00000000; // 5875 :   0 - 0x0
      13'h16F4: dout  = 8'b00000000; // 5876 :   0 - 0x0
      13'h16F5: dout  = 8'b00000000; // 5877 :   0 - 0x0
      13'h16F6: dout  = 8'b00000000; // 5878 :   0 - 0x0
      13'h16F7: dout  = 8'b00000000; // 5879 :   0 - 0x0
      13'h16F8: dout  = 8'b00000000; // 5880 :   0 - 0x0
      13'h16F9: dout  = 8'b00000000; // 5881 :   0 - 0x0
      13'h16FA: dout  = 8'b00000000; // 5882 :   0 - 0x0
      13'h16FB: dout  = 8'b00000000; // 5883 :   0 - 0x0
      13'h16FC: dout  = 8'b00000000; // 5884 :   0 - 0x0
      13'h16FD: dout  = 8'b00000000; // 5885 :   0 - 0x0
      13'h16FE: dout  = 8'b00000000; // 5886 :   0 - 0x0
      13'h16FF: dout  = 8'b00000000; // 5887 :   0 - 0x0
      13'h1700: dout  = 8'b00000000; // 5888 :   0 - 0x0 -- Background 0x70
      13'h1701: dout  = 8'b00000000; // 5889 :   0 - 0x0
      13'h1702: dout  = 8'b00000000; // 5890 :   0 - 0x0
      13'h1703: dout  = 8'b00000000; // 5891 :   0 - 0x0
      13'h1704: dout  = 8'b00000000; // 5892 :   0 - 0x0
      13'h1705: dout  = 8'b00000000; // 5893 :   0 - 0x0
      13'h1706: dout  = 8'b00000000; // 5894 :   0 - 0x0
      13'h1707: dout  = 8'b00000000; // 5895 :   0 - 0x0
      13'h1708: dout  = 8'b00000000; // 5896 :   0 - 0x0
      13'h1709: dout  = 8'b00000000; // 5897 :   0 - 0x0
      13'h170A: dout  = 8'b00000000; // 5898 :   0 - 0x0
      13'h170B: dout  = 8'b00000000; // 5899 :   0 - 0x0
      13'h170C: dout  = 8'b00000000; // 5900 :   0 - 0x0
      13'h170D: dout  = 8'b00000000; // 5901 :   0 - 0x0
      13'h170E: dout  = 8'b00000000; // 5902 :   0 - 0x0
      13'h170F: dout  = 8'b00000000; // 5903 :   0 - 0x0
      13'h1710: dout  = 8'b00000000; // 5904 :   0 - 0x0 -- Background 0x71
      13'h1711: dout  = 8'b00000000; // 5905 :   0 - 0x0
      13'h1712: dout  = 8'b00000000; // 5906 :   0 - 0x0
      13'h1713: dout  = 8'b00000000; // 5907 :   0 - 0x0
      13'h1714: dout  = 8'b00000000; // 5908 :   0 - 0x0
      13'h1715: dout  = 8'b00000000; // 5909 :   0 - 0x0
      13'h1716: dout  = 8'b00000000; // 5910 :   0 - 0x0
      13'h1717: dout  = 8'b00000000; // 5911 :   0 - 0x0
      13'h1718: dout  = 8'b00000000; // 5912 :   0 - 0x0
      13'h1719: dout  = 8'b00000000; // 5913 :   0 - 0x0
      13'h171A: dout  = 8'b00000000; // 5914 :   0 - 0x0
      13'h171B: dout  = 8'b00000000; // 5915 :   0 - 0x0
      13'h171C: dout  = 8'b00000000; // 5916 :   0 - 0x0
      13'h171D: dout  = 8'b00000000; // 5917 :   0 - 0x0
      13'h171E: dout  = 8'b00000000; // 5918 :   0 - 0x0
      13'h171F: dout  = 8'b00000000; // 5919 :   0 - 0x0
      13'h1720: dout  = 8'b00000000; // 5920 :   0 - 0x0 -- Background 0x72
      13'h1721: dout  = 8'b00000000; // 5921 :   0 - 0x0
      13'h1722: dout  = 8'b00000000; // 5922 :   0 - 0x0
      13'h1723: dout  = 8'b00000000; // 5923 :   0 - 0x0
      13'h1724: dout  = 8'b00000000; // 5924 :   0 - 0x0
      13'h1725: dout  = 8'b00000000; // 5925 :   0 - 0x0
      13'h1726: dout  = 8'b00000000; // 5926 :   0 - 0x0
      13'h1727: dout  = 8'b00000000; // 5927 :   0 - 0x0
      13'h1728: dout  = 8'b00000000; // 5928 :   0 - 0x0
      13'h1729: dout  = 8'b00000000; // 5929 :   0 - 0x0
      13'h172A: dout  = 8'b00000000; // 5930 :   0 - 0x0
      13'h172B: dout  = 8'b00000000; // 5931 :   0 - 0x0
      13'h172C: dout  = 8'b00000000; // 5932 :   0 - 0x0
      13'h172D: dout  = 8'b00000000; // 5933 :   0 - 0x0
      13'h172E: dout  = 8'b00000000; // 5934 :   0 - 0x0
      13'h172F: dout  = 8'b00000000; // 5935 :   0 - 0x0
      13'h1730: dout  = 8'b00000000; // 5936 :   0 - 0x0 -- Background 0x73
      13'h1731: dout  = 8'b00000000; // 5937 :   0 - 0x0
      13'h1732: dout  = 8'b00000000; // 5938 :   0 - 0x0
      13'h1733: dout  = 8'b00000000; // 5939 :   0 - 0x0
      13'h1734: dout  = 8'b00000000; // 5940 :   0 - 0x0
      13'h1735: dout  = 8'b00000000; // 5941 :   0 - 0x0
      13'h1736: dout  = 8'b00000000; // 5942 :   0 - 0x0
      13'h1737: dout  = 8'b00000000; // 5943 :   0 - 0x0
      13'h1738: dout  = 8'b00000000; // 5944 :   0 - 0x0
      13'h1739: dout  = 8'b00000000; // 5945 :   0 - 0x0
      13'h173A: dout  = 8'b00000000; // 5946 :   0 - 0x0
      13'h173B: dout  = 8'b00000000; // 5947 :   0 - 0x0
      13'h173C: dout  = 8'b00000000; // 5948 :   0 - 0x0
      13'h173D: dout  = 8'b00000000; // 5949 :   0 - 0x0
      13'h173E: dout  = 8'b00000000; // 5950 :   0 - 0x0
      13'h173F: dout  = 8'b00000000; // 5951 :   0 - 0x0
      13'h1740: dout  = 8'b00000000; // 5952 :   0 - 0x0 -- Background 0x74
      13'h1741: dout  = 8'b00000000; // 5953 :   0 - 0x0
      13'h1742: dout  = 8'b00000000; // 5954 :   0 - 0x0
      13'h1743: dout  = 8'b00000000; // 5955 :   0 - 0x0
      13'h1744: dout  = 8'b00000000; // 5956 :   0 - 0x0
      13'h1745: dout  = 8'b00000000; // 5957 :   0 - 0x0
      13'h1746: dout  = 8'b00000000; // 5958 :   0 - 0x0
      13'h1747: dout  = 8'b00000000; // 5959 :   0 - 0x0
      13'h1748: dout  = 8'b00000000; // 5960 :   0 - 0x0
      13'h1749: dout  = 8'b00000000; // 5961 :   0 - 0x0
      13'h174A: dout  = 8'b00000000; // 5962 :   0 - 0x0
      13'h174B: dout  = 8'b00000000; // 5963 :   0 - 0x0
      13'h174C: dout  = 8'b00000000; // 5964 :   0 - 0x0
      13'h174D: dout  = 8'b00000000; // 5965 :   0 - 0x0
      13'h174E: dout  = 8'b00000000; // 5966 :   0 - 0x0
      13'h174F: dout  = 8'b00000000; // 5967 :   0 - 0x0
      13'h1750: dout  = 8'b00000000; // 5968 :   0 - 0x0 -- Background 0x75
      13'h1751: dout  = 8'b00000000; // 5969 :   0 - 0x0
      13'h1752: dout  = 8'b00000000; // 5970 :   0 - 0x0
      13'h1753: dout  = 8'b00000000; // 5971 :   0 - 0x0
      13'h1754: dout  = 8'b00000000; // 5972 :   0 - 0x0
      13'h1755: dout  = 8'b00000000; // 5973 :   0 - 0x0
      13'h1756: dout  = 8'b00000000; // 5974 :   0 - 0x0
      13'h1757: dout  = 8'b00000000; // 5975 :   0 - 0x0
      13'h1758: dout  = 8'b00000000; // 5976 :   0 - 0x0
      13'h1759: dout  = 8'b00000000; // 5977 :   0 - 0x0
      13'h175A: dout  = 8'b00000000; // 5978 :   0 - 0x0
      13'h175B: dout  = 8'b00000000; // 5979 :   0 - 0x0
      13'h175C: dout  = 8'b00000000; // 5980 :   0 - 0x0
      13'h175D: dout  = 8'b00000000; // 5981 :   0 - 0x0
      13'h175E: dout  = 8'b00000000; // 5982 :   0 - 0x0
      13'h175F: dout  = 8'b00000000; // 5983 :   0 - 0x0
      13'h1760: dout  = 8'b00000000; // 5984 :   0 - 0x0 -- Background 0x76
      13'h1761: dout  = 8'b00000000; // 5985 :   0 - 0x0
      13'h1762: dout  = 8'b00000000; // 5986 :   0 - 0x0
      13'h1763: dout  = 8'b00000000; // 5987 :   0 - 0x0
      13'h1764: dout  = 8'b00000000; // 5988 :   0 - 0x0
      13'h1765: dout  = 8'b00000000; // 5989 :   0 - 0x0
      13'h1766: dout  = 8'b00000000; // 5990 :   0 - 0x0
      13'h1767: dout  = 8'b00000000; // 5991 :   0 - 0x0
      13'h1768: dout  = 8'b00000000; // 5992 :   0 - 0x0
      13'h1769: dout  = 8'b00000000; // 5993 :   0 - 0x0
      13'h176A: dout  = 8'b00000000; // 5994 :   0 - 0x0
      13'h176B: dout  = 8'b00000000; // 5995 :   0 - 0x0
      13'h176C: dout  = 8'b00000000; // 5996 :   0 - 0x0
      13'h176D: dout  = 8'b00000000; // 5997 :   0 - 0x0
      13'h176E: dout  = 8'b00000000; // 5998 :   0 - 0x0
      13'h176F: dout  = 8'b00000000; // 5999 :   0 - 0x0
      13'h1770: dout  = 8'b00000000; // 6000 :   0 - 0x0 -- Background 0x77
      13'h1771: dout  = 8'b00000000; // 6001 :   0 - 0x0
      13'h1772: dout  = 8'b00000000; // 6002 :   0 - 0x0
      13'h1773: dout  = 8'b00000000; // 6003 :   0 - 0x0
      13'h1774: dout  = 8'b00000000; // 6004 :   0 - 0x0
      13'h1775: dout  = 8'b00000000; // 6005 :   0 - 0x0
      13'h1776: dout  = 8'b00000000; // 6006 :   0 - 0x0
      13'h1777: dout  = 8'b00000000; // 6007 :   0 - 0x0
      13'h1778: dout  = 8'b00000000; // 6008 :   0 - 0x0
      13'h1779: dout  = 8'b00000000; // 6009 :   0 - 0x0
      13'h177A: dout  = 8'b00000000; // 6010 :   0 - 0x0
      13'h177B: dout  = 8'b00000000; // 6011 :   0 - 0x0
      13'h177C: dout  = 8'b00000000; // 6012 :   0 - 0x0
      13'h177D: dout  = 8'b00000000; // 6013 :   0 - 0x0
      13'h177E: dout  = 8'b00000000; // 6014 :   0 - 0x0
      13'h177F: dout  = 8'b00000000; // 6015 :   0 - 0x0
      13'h1780: dout  = 8'b00000000; // 6016 :   0 - 0x0 -- Background 0x78
      13'h1781: dout  = 8'b00000000; // 6017 :   0 - 0x0
      13'h1782: dout  = 8'b00000000; // 6018 :   0 - 0x0
      13'h1783: dout  = 8'b00000000; // 6019 :   0 - 0x0
      13'h1784: dout  = 8'b00000000; // 6020 :   0 - 0x0
      13'h1785: dout  = 8'b00000000; // 6021 :   0 - 0x0
      13'h1786: dout  = 8'b00000000; // 6022 :   0 - 0x0
      13'h1787: dout  = 8'b00000000; // 6023 :   0 - 0x0
      13'h1788: dout  = 8'b00000000; // 6024 :   0 - 0x0
      13'h1789: dout  = 8'b00000000; // 6025 :   0 - 0x0
      13'h178A: dout  = 8'b00000000; // 6026 :   0 - 0x0
      13'h178B: dout  = 8'b00000000; // 6027 :   0 - 0x0
      13'h178C: dout  = 8'b00000000; // 6028 :   0 - 0x0
      13'h178D: dout  = 8'b00000000; // 6029 :   0 - 0x0
      13'h178E: dout  = 8'b00000000; // 6030 :   0 - 0x0
      13'h178F: dout  = 8'b00000000; // 6031 :   0 - 0x0
      13'h1790: dout  = 8'b00000000; // 6032 :   0 - 0x0 -- Background 0x79
      13'h1791: dout  = 8'b00000000; // 6033 :   0 - 0x0
      13'h1792: dout  = 8'b00000000; // 6034 :   0 - 0x0
      13'h1793: dout  = 8'b00000000; // 6035 :   0 - 0x0
      13'h1794: dout  = 8'b00000000; // 6036 :   0 - 0x0
      13'h1795: dout  = 8'b00000000; // 6037 :   0 - 0x0
      13'h1796: dout  = 8'b00000000; // 6038 :   0 - 0x0
      13'h1797: dout  = 8'b00000000; // 6039 :   0 - 0x0
      13'h1798: dout  = 8'b00000000; // 6040 :   0 - 0x0
      13'h1799: dout  = 8'b00000000; // 6041 :   0 - 0x0
      13'h179A: dout  = 8'b00000000; // 6042 :   0 - 0x0
      13'h179B: dout  = 8'b00000000; // 6043 :   0 - 0x0
      13'h179C: dout  = 8'b00000000; // 6044 :   0 - 0x0
      13'h179D: dout  = 8'b00000000; // 6045 :   0 - 0x0
      13'h179E: dout  = 8'b00000000; // 6046 :   0 - 0x0
      13'h179F: dout  = 8'b00000000; // 6047 :   0 - 0x0
      13'h17A0: dout  = 8'b00000000; // 6048 :   0 - 0x0 -- Background 0x7a
      13'h17A1: dout  = 8'b00000000; // 6049 :   0 - 0x0
      13'h17A2: dout  = 8'b00000000; // 6050 :   0 - 0x0
      13'h17A3: dout  = 8'b00000000; // 6051 :   0 - 0x0
      13'h17A4: dout  = 8'b00000000; // 6052 :   0 - 0x0
      13'h17A5: dout  = 8'b00000000; // 6053 :   0 - 0x0
      13'h17A6: dout  = 8'b00000000; // 6054 :   0 - 0x0
      13'h17A7: dout  = 8'b00000000; // 6055 :   0 - 0x0
      13'h17A8: dout  = 8'b00000000; // 6056 :   0 - 0x0
      13'h17A9: dout  = 8'b00000000; // 6057 :   0 - 0x0
      13'h17AA: dout  = 8'b00000000; // 6058 :   0 - 0x0
      13'h17AB: dout  = 8'b00000000; // 6059 :   0 - 0x0
      13'h17AC: dout  = 8'b00000000; // 6060 :   0 - 0x0
      13'h17AD: dout  = 8'b00000000; // 6061 :   0 - 0x0
      13'h17AE: dout  = 8'b00000000; // 6062 :   0 - 0x0
      13'h17AF: dout  = 8'b00000000; // 6063 :   0 - 0x0
      13'h17B0: dout  = 8'b00000000; // 6064 :   0 - 0x0 -- Background 0x7b
      13'h17B1: dout  = 8'b00000000; // 6065 :   0 - 0x0
      13'h17B2: dout  = 8'b00000000; // 6066 :   0 - 0x0
      13'h17B3: dout  = 8'b00000000; // 6067 :   0 - 0x0
      13'h17B4: dout  = 8'b00000000; // 6068 :   0 - 0x0
      13'h17B5: dout  = 8'b00000000; // 6069 :   0 - 0x0
      13'h17B6: dout  = 8'b00000000; // 6070 :   0 - 0x0
      13'h17B7: dout  = 8'b00000000; // 6071 :   0 - 0x0
      13'h17B8: dout  = 8'b00000000; // 6072 :   0 - 0x0
      13'h17B9: dout  = 8'b00000000; // 6073 :   0 - 0x0
      13'h17BA: dout  = 8'b00000000; // 6074 :   0 - 0x0
      13'h17BB: dout  = 8'b00000000; // 6075 :   0 - 0x0
      13'h17BC: dout  = 8'b00000000; // 6076 :   0 - 0x0
      13'h17BD: dout  = 8'b00000000; // 6077 :   0 - 0x0
      13'h17BE: dout  = 8'b00000000; // 6078 :   0 - 0x0
      13'h17BF: dout  = 8'b00000000; // 6079 :   0 - 0x0
      13'h17C0: dout  = 8'b00000000; // 6080 :   0 - 0x0 -- Background 0x7c
      13'h17C1: dout  = 8'b00000000; // 6081 :   0 - 0x0
      13'h17C2: dout  = 8'b00000000; // 6082 :   0 - 0x0
      13'h17C3: dout  = 8'b00000000; // 6083 :   0 - 0x0
      13'h17C4: dout  = 8'b00000000; // 6084 :   0 - 0x0
      13'h17C5: dout  = 8'b00000000; // 6085 :   0 - 0x0
      13'h17C6: dout  = 8'b00000000; // 6086 :   0 - 0x0
      13'h17C7: dout  = 8'b00000000; // 6087 :   0 - 0x0
      13'h17C8: dout  = 8'b00000000; // 6088 :   0 - 0x0
      13'h17C9: dout  = 8'b00000000; // 6089 :   0 - 0x0
      13'h17CA: dout  = 8'b00000000; // 6090 :   0 - 0x0
      13'h17CB: dout  = 8'b00000000; // 6091 :   0 - 0x0
      13'h17CC: dout  = 8'b00000000; // 6092 :   0 - 0x0
      13'h17CD: dout  = 8'b00000000; // 6093 :   0 - 0x0
      13'h17CE: dout  = 8'b00000000; // 6094 :   0 - 0x0
      13'h17CF: dout  = 8'b00000000; // 6095 :   0 - 0x0
      13'h17D0: dout  = 8'b00000000; // 6096 :   0 - 0x0 -- Background 0x7d
      13'h17D1: dout  = 8'b00000000; // 6097 :   0 - 0x0
      13'h17D2: dout  = 8'b00000000; // 6098 :   0 - 0x0
      13'h17D3: dout  = 8'b00000000; // 6099 :   0 - 0x0
      13'h17D4: dout  = 8'b00000000; // 6100 :   0 - 0x0
      13'h17D5: dout  = 8'b00000000; // 6101 :   0 - 0x0
      13'h17D6: dout  = 8'b00000000; // 6102 :   0 - 0x0
      13'h17D7: dout  = 8'b00000000; // 6103 :   0 - 0x0
      13'h17D8: dout  = 8'b00000000; // 6104 :   0 - 0x0
      13'h17D9: dout  = 8'b00000000; // 6105 :   0 - 0x0
      13'h17DA: dout  = 8'b00000000; // 6106 :   0 - 0x0
      13'h17DB: dout  = 8'b00000000; // 6107 :   0 - 0x0
      13'h17DC: dout  = 8'b00000000; // 6108 :   0 - 0x0
      13'h17DD: dout  = 8'b00000000; // 6109 :   0 - 0x0
      13'h17DE: dout  = 8'b00000000; // 6110 :   0 - 0x0
      13'h17DF: dout  = 8'b00000000; // 6111 :   0 - 0x0
      13'h17E0: dout  = 8'b00000000; // 6112 :   0 - 0x0 -- Background 0x7e
      13'h17E1: dout  = 8'b00000000; // 6113 :   0 - 0x0
      13'h17E2: dout  = 8'b00000000; // 6114 :   0 - 0x0
      13'h17E3: dout  = 8'b00000000; // 6115 :   0 - 0x0
      13'h17E4: dout  = 8'b00000000; // 6116 :   0 - 0x0
      13'h17E5: dout  = 8'b00000000; // 6117 :   0 - 0x0
      13'h17E6: dout  = 8'b00000000; // 6118 :   0 - 0x0
      13'h17E7: dout  = 8'b00000000; // 6119 :   0 - 0x0
      13'h17E8: dout  = 8'b00000000; // 6120 :   0 - 0x0
      13'h17E9: dout  = 8'b00000000; // 6121 :   0 - 0x0
      13'h17EA: dout  = 8'b00000000; // 6122 :   0 - 0x0
      13'h17EB: dout  = 8'b00000000; // 6123 :   0 - 0x0
      13'h17EC: dout  = 8'b00000000; // 6124 :   0 - 0x0
      13'h17ED: dout  = 8'b00000000; // 6125 :   0 - 0x0
      13'h17EE: dout  = 8'b00000000; // 6126 :   0 - 0x0
      13'h17EF: dout  = 8'b00000000; // 6127 :   0 - 0x0
      13'h17F0: dout  = 8'b00000000; // 6128 :   0 - 0x0 -- Background 0x7f
      13'h17F1: dout  = 8'b00000000; // 6129 :   0 - 0x0
      13'h17F2: dout  = 8'b00000000; // 6130 :   0 - 0x0
      13'h17F3: dout  = 8'b00000000; // 6131 :   0 - 0x0
      13'h17F4: dout  = 8'b00000000; // 6132 :   0 - 0x0
      13'h17F5: dout  = 8'b00000000; // 6133 :   0 - 0x0
      13'h17F6: dout  = 8'b00000000; // 6134 :   0 - 0x0
      13'h17F7: dout  = 8'b00000000; // 6135 :   0 - 0x0
      13'h17F8: dout  = 8'b00000000; // 6136 :   0 - 0x0
      13'h17F9: dout  = 8'b00000000; // 6137 :   0 - 0x0
      13'h17FA: dout  = 8'b00000000; // 6138 :   0 - 0x0
      13'h17FB: dout  = 8'b00000000; // 6139 :   0 - 0x0
      13'h17FC: dout  = 8'b00000000; // 6140 :   0 - 0x0
      13'h17FD: dout  = 8'b00000000; // 6141 :   0 - 0x0
      13'h17FE: dout  = 8'b00000000; // 6142 :   0 - 0x0
      13'h17FF: dout  = 8'b00000000; // 6143 :   0 - 0x0
      13'h1800: dout  = 8'b00000000; // 6144 :   0 - 0x0 -- Background 0x80
      13'h1801: dout  = 8'b00000000; // 6145 :   0 - 0x0
      13'h1802: dout  = 8'b00000000; // 6146 :   0 - 0x0
      13'h1803: dout  = 8'b00000000; // 6147 :   0 - 0x0
      13'h1804: dout  = 8'b00000000; // 6148 :   0 - 0x0
      13'h1805: dout  = 8'b00000000; // 6149 :   0 - 0x0
      13'h1806: dout  = 8'b00000000; // 6150 :   0 - 0x0
      13'h1807: dout  = 8'b00000000; // 6151 :   0 - 0x0
      13'h1808: dout  = 8'b00000000; // 6152 :   0 - 0x0
      13'h1809: dout  = 8'b00000000; // 6153 :   0 - 0x0
      13'h180A: dout  = 8'b00000000; // 6154 :   0 - 0x0
      13'h180B: dout  = 8'b00000000; // 6155 :   0 - 0x0
      13'h180C: dout  = 8'b00000000; // 6156 :   0 - 0x0
      13'h180D: dout  = 8'b00000000; // 6157 :   0 - 0x0
      13'h180E: dout  = 8'b00000000; // 6158 :   0 - 0x0
      13'h180F: dout  = 8'b00000000; // 6159 :   0 - 0x0
      13'h1810: dout  = 8'b00000000; // 6160 :   0 - 0x0 -- Background 0x81
      13'h1811: dout  = 8'b00000000; // 6161 :   0 - 0x0
      13'h1812: dout  = 8'b00000000; // 6162 :   0 - 0x0
      13'h1813: dout  = 8'b00000000; // 6163 :   0 - 0x0
      13'h1814: dout  = 8'b00000000; // 6164 :   0 - 0x0
      13'h1815: dout  = 8'b00000000; // 6165 :   0 - 0x0
      13'h1816: dout  = 8'b00000000; // 6166 :   0 - 0x0
      13'h1817: dout  = 8'b00000000; // 6167 :   0 - 0x0
      13'h1818: dout  = 8'b00000000; // 6168 :   0 - 0x0
      13'h1819: dout  = 8'b00000000; // 6169 :   0 - 0x0
      13'h181A: dout  = 8'b00000000; // 6170 :   0 - 0x0
      13'h181B: dout  = 8'b00000000; // 6171 :   0 - 0x0
      13'h181C: dout  = 8'b00000000; // 6172 :   0 - 0x0
      13'h181D: dout  = 8'b00000000; // 6173 :   0 - 0x0
      13'h181E: dout  = 8'b00000000; // 6174 :   0 - 0x0
      13'h181F: dout  = 8'b00000000; // 6175 :   0 - 0x0
      13'h1820: dout  = 8'b00000000; // 6176 :   0 - 0x0 -- Background 0x82
      13'h1821: dout  = 8'b00000000; // 6177 :   0 - 0x0
      13'h1822: dout  = 8'b00000000; // 6178 :   0 - 0x0
      13'h1823: dout  = 8'b00000000; // 6179 :   0 - 0x0
      13'h1824: dout  = 8'b00000000; // 6180 :   0 - 0x0
      13'h1825: dout  = 8'b00000000; // 6181 :   0 - 0x0
      13'h1826: dout  = 8'b00000000; // 6182 :   0 - 0x0
      13'h1827: dout  = 8'b00000000; // 6183 :   0 - 0x0
      13'h1828: dout  = 8'b00000000; // 6184 :   0 - 0x0
      13'h1829: dout  = 8'b00000000; // 6185 :   0 - 0x0
      13'h182A: dout  = 8'b00000000; // 6186 :   0 - 0x0
      13'h182B: dout  = 8'b00000000; // 6187 :   0 - 0x0
      13'h182C: dout  = 8'b00000000; // 6188 :   0 - 0x0
      13'h182D: dout  = 8'b00000000; // 6189 :   0 - 0x0
      13'h182E: dout  = 8'b00000000; // 6190 :   0 - 0x0
      13'h182F: dout  = 8'b00000000; // 6191 :   0 - 0x0
      13'h1830: dout  = 8'b00000000; // 6192 :   0 - 0x0 -- Background 0x83
      13'h1831: dout  = 8'b00000000; // 6193 :   0 - 0x0
      13'h1832: dout  = 8'b00000000; // 6194 :   0 - 0x0
      13'h1833: dout  = 8'b00000000; // 6195 :   0 - 0x0
      13'h1834: dout  = 8'b00000000; // 6196 :   0 - 0x0
      13'h1835: dout  = 8'b00000000; // 6197 :   0 - 0x0
      13'h1836: dout  = 8'b00000000; // 6198 :   0 - 0x0
      13'h1837: dout  = 8'b00000000; // 6199 :   0 - 0x0
      13'h1838: dout  = 8'b00000000; // 6200 :   0 - 0x0
      13'h1839: dout  = 8'b00000000; // 6201 :   0 - 0x0
      13'h183A: dout  = 8'b00000000; // 6202 :   0 - 0x0
      13'h183B: dout  = 8'b00000000; // 6203 :   0 - 0x0
      13'h183C: dout  = 8'b00000000; // 6204 :   0 - 0x0
      13'h183D: dout  = 8'b00000000; // 6205 :   0 - 0x0
      13'h183E: dout  = 8'b00000000; // 6206 :   0 - 0x0
      13'h183F: dout  = 8'b00000000; // 6207 :   0 - 0x0
      13'h1840: dout  = 8'b00000000; // 6208 :   0 - 0x0 -- Background 0x84
      13'h1841: dout  = 8'b00000000; // 6209 :   0 - 0x0
      13'h1842: dout  = 8'b00000000; // 6210 :   0 - 0x0
      13'h1843: dout  = 8'b00000000; // 6211 :   0 - 0x0
      13'h1844: dout  = 8'b00000000; // 6212 :   0 - 0x0
      13'h1845: dout  = 8'b00000000; // 6213 :   0 - 0x0
      13'h1846: dout  = 8'b00000000; // 6214 :   0 - 0x0
      13'h1847: dout  = 8'b00000000; // 6215 :   0 - 0x0
      13'h1848: dout  = 8'b00000000; // 6216 :   0 - 0x0
      13'h1849: dout  = 8'b00000000; // 6217 :   0 - 0x0
      13'h184A: dout  = 8'b00000000; // 6218 :   0 - 0x0
      13'h184B: dout  = 8'b00000000; // 6219 :   0 - 0x0
      13'h184C: dout  = 8'b00000000; // 6220 :   0 - 0x0
      13'h184D: dout  = 8'b00000000; // 6221 :   0 - 0x0
      13'h184E: dout  = 8'b00000000; // 6222 :   0 - 0x0
      13'h184F: dout  = 8'b00000000; // 6223 :   0 - 0x0
      13'h1850: dout  = 8'b00000000; // 6224 :   0 - 0x0 -- Background 0x85
      13'h1851: dout  = 8'b00000000; // 6225 :   0 - 0x0
      13'h1852: dout  = 8'b00000000; // 6226 :   0 - 0x0
      13'h1853: dout  = 8'b00000000; // 6227 :   0 - 0x0
      13'h1854: dout  = 8'b00000000; // 6228 :   0 - 0x0
      13'h1855: dout  = 8'b00000000; // 6229 :   0 - 0x0
      13'h1856: dout  = 8'b00000000; // 6230 :   0 - 0x0
      13'h1857: dout  = 8'b00000000; // 6231 :   0 - 0x0
      13'h1858: dout  = 8'b00000000; // 6232 :   0 - 0x0
      13'h1859: dout  = 8'b00000000; // 6233 :   0 - 0x0
      13'h185A: dout  = 8'b00000000; // 6234 :   0 - 0x0
      13'h185B: dout  = 8'b00000000; // 6235 :   0 - 0x0
      13'h185C: dout  = 8'b00000000; // 6236 :   0 - 0x0
      13'h185D: dout  = 8'b00000000; // 6237 :   0 - 0x0
      13'h185E: dout  = 8'b00000000; // 6238 :   0 - 0x0
      13'h185F: dout  = 8'b00000000; // 6239 :   0 - 0x0
      13'h1860: dout  = 8'b00000000; // 6240 :   0 - 0x0 -- Background 0x86
      13'h1861: dout  = 8'b00000000; // 6241 :   0 - 0x0
      13'h1862: dout  = 8'b00000000; // 6242 :   0 - 0x0
      13'h1863: dout  = 8'b00000000; // 6243 :   0 - 0x0
      13'h1864: dout  = 8'b00000000; // 6244 :   0 - 0x0
      13'h1865: dout  = 8'b00000000; // 6245 :   0 - 0x0
      13'h1866: dout  = 8'b00000000; // 6246 :   0 - 0x0
      13'h1867: dout  = 8'b00000000; // 6247 :   0 - 0x0
      13'h1868: dout  = 8'b00000000; // 6248 :   0 - 0x0
      13'h1869: dout  = 8'b00000000; // 6249 :   0 - 0x0
      13'h186A: dout  = 8'b00000000; // 6250 :   0 - 0x0
      13'h186B: dout  = 8'b00000000; // 6251 :   0 - 0x0
      13'h186C: dout  = 8'b00000000; // 6252 :   0 - 0x0
      13'h186D: dout  = 8'b00000000; // 6253 :   0 - 0x0
      13'h186E: dout  = 8'b00000000; // 6254 :   0 - 0x0
      13'h186F: dout  = 8'b00000000; // 6255 :   0 - 0x0
      13'h1870: dout  = 8'b00000000; // 6256 :   0 - 0x0 -- Background 0x87
      13'h1871: dout  = 8'b00000000; // 6257 :   0 - 0x0
      13'h1872: dout  = 8'b00000000; // 6258 :   0 - 0x0
      13'h1873: dout  = 8'b00000000; // 6259 :   0 - 0x0
      13'h1874: dout  = 8'b00000000; // 6260 :   0 - 0x0
      13'h1875: dout  = 8'b00000000; // 6261 :   0 - 0x0
      13'h1876: dout  = 8'b00000000; // 6262 :   0 - 0x0
      13'h1877: dout  = 8'b00000000; // 6263 :   0 - 0x0
      13'h1878: dout  = 8'b00000000; // 6264 :   0 - 0x0
      13'h1879: dout  = 8'b00000000; // 6265 :   0 - 0x0
      13'h187A: dout  = 8'b00000000; // 6266 :   0 - 0x0
      13'h187B: dout  = 8'b00000000; // 6267 :   0 - 0x0
      13'h187C: dout  = 8'b00000000; // 6268 :   0 - 0x0
      13'h187D: dout  = 8'b00000000; // 6269 :   0 - 0x0
      13'h187E: dout  = 8'b00000000; // 6270 :   0 - 0x0
      13'h187F: dout  = 8'b00000000; // 6271 :   0 - 0x0
      13'h1880: dout  = 8'b00000000; // 6272 :   0 - 0x0 -- Background 0x88
      13'h1881: dout  = 8'b00000000; // 6273 :   0 - 0x0
      13'h1882: dout  = 8'b00000000; // 6274 :   0 - 0x0
      13'h1883: dout  = 8'b00000000; // 6275 :   0 - 0x0
      13'h1884: dout  = 8'b00000000; // 6276 :   0 - 0x0
      13'h1885: dout  = 8'b00000000; // 6277 :   0 - 0x0
      13'h1886: dout  = 8'b00000000; // 6278 :   0 - 0x0
      13'h1887: dout  = 8'b00000000; // 6279 :   0 - 0x0
      13'h1888: dout  = 8'b00000000; // 6280 :   0 - 0x0
      13'h1889: dout  = 8'b00000000; // 6281 :   0 - 0x0
      13'h188A: dout  = 8'b00000000; // 6282 :   0 - 0x0
      13'h188B: dout  = 8'b00000000; // 6283 :   0 - 0x0
      13'h188C: dout  = 8'b00000000; // 6284 :   0 - 0x0
      13'h188D: dout  = 8'b00000000; // 6285 :   0 - 0x0
      13'h188E: dout  = 8'b00000000; // 6286 :   0 - 0x0
      13'h188F: dout  = 8'b00000000; // 6287 :   0 - 0x0
      13'h1890: dout  = 8'b00000000; // 6288 :   0 - 0x0 -- Background 0x89
      13'h1891: dout  = 8'b00000000; // 6289 :   0 - 0x0
      13'h1892: dout  = 8'b00000000; // 6290 :   0 - 0x0
      13'h1893: dout  = 8'b00000000; // 6291 :   0 - 0x0
      13'h1894: dout  = 8'b00000000; // 6292 :   0 - 0x0
      13'h1895: dout  = 8'b00000000; // 6293 :   0 - 0x0
      13'h1896: dout  = 8'b00000000; // 6294 :   0 - 0x0
      13'h1897: dout  = 8'b00000000; // 6295 :   0 - 0x0
      13'h1898: dout  = 8'b00000000; // 6296 :   0 - 0x0
      13'h1899: dout  = 8'b00000000; // 6297 :   0 - 0x0
      13'h189A: dout  = 8'b00000000; // 6298 :   0 - 0x0
      13'h189B: dout  = 8'b00000000; // 6299 :   0 - 0x0
      13'h189C: dout  = 8'b00000000; // 6300 :   0 - 0x0
      13'h189D: dout  = 8'b00000000; // 6301 :   0 - 0x0
      13'h189E: dout  = 8'b00000000; // 6302 :   0 - 0x0
      13'h189F: dout  = 8'b00000000; // 6303 :   0 - 0x0
      13'h18A0: dout  = 8'b00000000; // 6304 :   0 - 0x0 -- Background 0x8a
      13'h18A1: dout  = 8'b00000000; // 6305 :   0 - 0x0
      13'h18A2: dout  = 8'b00000000; // 6306 :   0 - 0x0
      13'h18A3: dout  = 8'b00000000; // 6307 :   0 - 0x0
      13'h18A4: dout  = 8'b00000000; // 6308 :   0 - 0x0
      13'h18A5: dout  = 8'b00000000; // 6309 :   0 - 0x0
      13'h18A6: dout  = 8'b00000000; // 6310 :   0 - 0x0
      13'h18A7: dout  = 8'b00000000; // 6311 :   0 - 0x0
      13'h18A8: dout  = 8'b00000000; // 6312 :   0 - 0x0
      13'h18A9: dout  = 8'b00000000; // 6313 :   0 - 0x0
      13'h18AA: dout  = 8'b00000000; // 6314 :   0 - 0x0
      13'h18AB: dout  = 8'b00000000; // 6315 :   0 - 0x0
      13'h18AC: dout  = 8'b00000000; // 6316 :   0 - 0x0
      13'h18AD: dout  = 8'b00000000; // 6317 :   0 - 0x0
      13'h18AE: dout  = 8'b00000000; // 6318 :   0 - 0x0
      13'h18AF: dout  = 8'b00000000; // 6319 :   0 - 0x0
      13'h18B0: dout  = 8'b00000000; // 6320 :   0 - 0x0 -- Background 0x8b
      13'h18B1: dout  = 8'b00000000; // 6321 :   0 - 0x0
      13'h18B2: dout  = 8'b00000000; // 6322 :   0 - 0x0
      13'h18B3: dout  = 8'b00000000; // 6323 :   0 - 0x0
      13'h18B4: dout  = 8'b00000000; // 6324 :   0 - 0x0
      13'h18B5: dout  = 8'b00000000; // 6325 :   0 - 0x0
      13'h18B6: dout  = 8'b00000000; // 6326 :   0 - 0x0
      13'h18B7: dout  = 8'b00000000; // 6327 :   0 - 0x0
      13'h18B8: dout  = 8'b00000000; // 6328 :   0 - 0x0
      13'h18B9: dout  = 8'b00000000; // 6329 :   0 - 0x0
      13'h18BA: dout  = 8'b00000000; // 6330 :   0 - 0x0
      13'h18BB: dout  = 8'b00000000; // 6331 :   0 - 0x0
      13'h18BC: dout  = 8'b00000000; // 6332 :   0 - 0x0
      13'h18BD: dout  = 8'b00000000; // 6333 :   0 - 0x0
      13'h18BE: dout  = 8'b00000000; // 6334 :   0 - 0x0
      13'h18BF: dout  = 8'b00000000; // 6335 :   0 - 0x0
      13'h18C0: dout  = 8'b00000000; // 6336 :   0 - 0x0 -- Background 0x8c
      13'h18C1: dout  = 8'b00000000; // 6337 :   0 - 0x0
      13'h18C2: dout  = 8'b00000000; // 6338 :   0 - 0x0
      13'h18C3: dout  = 8'b00000000; // 6339 :   0 - 0x0
      13'h18C4: dout  = 8'b00000000; // 6340 :   0 - 0x0
      13'h18C5: dout  = 8'b00000000; // 6341 :   0 - 0x0
      13'h18C6: dout  = 8'b00000000; // 6342 :   0 - 0x0
      13'h18C7: dout  = 8'b00000000; // 6343 :   0 - 0x0
      13'h18C8: dout  = 8'b00000000; // 6344 :   0 - 0x0
      13'h18C9: dout  = 8'b00000000; // 6345 :   0 - 0x0
      13'h18CA: dout  = 8'b00000000; // 6346 :   0 - 0x0
      13'h18CB: dout  = 8'b00000000; // 6347 :   0 - 0x0
      13'h18CC: dout  = 8'b00000000; // 6348 :   0 - 0x0
      13'h18CD: dout  = 8'b00000000; // 6349 :   0 - 0x0
      13'h18CE: dout  = 8'b00000000; // 6350 :   0 - 0x0
      13'h18CF: dout  = 8'b00000000; // 6351 :   0 - 0x0
      13'h18D0: dout  = 8'b00000000; // 6352 :   0 - 0x0 -- Background 0x8d
      13'h18D1: dout  = 8'b00000000; // 6353 :   0 - 0x0
      13'h18D2: dout  = 8'b00000000; // 6354 :   0 - 0x0
      13'h18D3: dout  = 8'b00000000; // 6355 :   0 - 0x0
      13'h18D4: dout  = 8'b00000000; // 6356 :   0 - 0x0
      13'h18D5: dout  = 8'b00000000; // 6357 :   0 - 0x0
      13'h18D6: dout  = 8'b00000000; // 6358 :   0 - 0x0
      13'h18D7: dout  = 8'b00000000; // 6359 :   0 - 0x0
      13'h18D8: dout  = 8'b00000000; // 6360 :   0 - 0x0
      13'h18D9: dout  = 8'b00000000; // 6361 :   0 - 0x0
      13'h18DA: dout  = 8'b00000000; // 6362 :   0 - 0x0
      13'h18DB: dout  = 8'b00000000; // 6363 :   0 - 0x0
      13'h18DC: dout  = 8'b00000000; // 6364 :   0 - 0x0
      13'h18DD: dout  = 8'b00000000; // 6365 :   0 - 0x0
      13'h18DE: dout  = 8'b00000000; // 6366 :   0 - 0x0
      13'h18DF: dout  = 8'b00000000; // 6367 :   0 - 0x0
      13'h18E0: dout  = 8'b00000000; // 6368 :   0 - 0x0 -- Background 0x8e
      13'h18E1: dout  = 8'b00000000; // 6369 :   0 - 0x0
      13'h18E2: dout  = 8'b00000000; // 6370 :   0 - 0x0
      13'h18E3: dout  = 8'b00000000; // 6371 :   0 - 0x0
      13'h18E4: dout  = 8'b00000000; // 6372 :   0 - 0x0
      13'h18E5: dout  = 8'b00000000; // 6373 :   0 - 0x0
      13'h18E6: dout  = 8'b00000000; // 6374 :   0 - 0x0
      13'h18E7: dout  = 8'b00000000; // 6375 :   0 - 0x0
      13'h18E8: dout  = 8'b00000000; // 6376 :   0 - 0x0
      13'h18E9: dout  = 8'b00000000; // 6377 :   0 - 0x0
      13'h18EA: dout  = 8'b00000000; // 6378 :   0 - 0x0
      13'h18EB: dout  = 8'b00000000; // 6379 :   0 - 0x0
      13'h18EC: dout  = 8'b00000000; // 6380 :   0 - 0x0
      13'h18ED: dout  = 8'b00000000; // 6381 :   0 - 0x0
      13'h18EE: dout  = 8'b00000000; // 6382 :   0 - 0x0
      13'h18EF: dout  = 8'b00000000; // 6383 :   0 - 0x0
      13'h18F0: dout  = 8'b00000000; // 6384 :   0 - 0x0 -- Background 0x8f
      13'h18F1: dout  = 8'b00000000; // 6385 :   0 - 0x0
      13'h18F2: dout  = 8'b00000000; // 6386 :   0 - 0x0
      13'h18F3: dout  = 8'b00000000; // 6387 :   0 - 0x0
      13'h18F4: dout  = 8'b00000000; // 6388 :   0 - 0x0
      13'h18F5: dout  = 8'b00000000; // 6389 :   0 - 0x0
      13'h18F6: dout  = 8'b00000000; // 6390 :   0 - 0x0
      13'h18F7: dout  = 8'b00000000; // 6391 :   0 - 0x0
      13'h18F8: dout  = 8'b00000000; // 6392 :   0 - 0x0
      13'h18F9: dout  = 8'b00000000; // 6393 :   0 - 0x0
      13'h18FA: dout  = 8'b00000000; // 6394 :   0 - 0x0
      13'h18FB: dout  = 8'b00000000; // 6395 :   0 - 0x0
      13'h18FC: dout  = 8'b00000000; // 6396 :   0 - 0x0
      13'h18FD: dout  = 8'b00000000; // 6397 :   0 - 0x0
      13'h18FE: dout  = 8'b00000000; // 6398 :   0 - 0x0
      13'h18FF: dout  = 8'b00000000; // 6399 :   0 - 0x0
      13'h1900: dout  = 8'b00000000; // 6400 :   0 - 0x0 -- Background 0x90
      13'h1901: dout  = 8'b00000000; // 6401 :   0 - 0x0
      13'h1902: dout  = 8'b00000000; // 6402 :   0 - 0x0
      13'h1903: dout  = 8'b00000000; // 6403 :   0 - 0x0
      13'h1904: dout  = 8'b00000000; // 6404 :   0 - 0x0
      13'h1905: dout  = 8'b00000000; // 6405 :   0 - 0x0
      13'h1906: dout  = 8'b00000000; // 6406 :   0 - 0x0
      13'h1907: dout  = 8'b00000000; // 6407 :   0 - 0x0
      13'h1908: dout  = 8'b00000000; // 6408 :   0 - 0x0
      13'h1909: dout  = 8'b00000000; // 6409 :   0 - 0x0
      13'h190A: dout  = 8'b00000000; // 6410 :   0 - 0x0
      13'h190B: dout  = 8'b00000000; // 6411 :   0 - 0x0
      13'h190C: dout  = 8'b00000000; // 6412 :   0 - 0x0
      13'h190D: dout  = 8'b00000000; // 6413 :   0 - 0x0
      13'h190E: dout  = 8'b00000000; // 6414 :   0 - 0x0
      13'h190F: dout  = 8'b00000000; // 6415 :   0 - 0x0
      13'h1910: dout  = 8'b00000000; // 6416 :   0 - 0x0 -- Background 0x91
      13'h1911: dout  = 8'b00000000; // 6417 :   0 - 0x0
      13'h1912: dout  = 8'b00000000; // 6418 :   0 - 0x0
      13'h1913: dout  = 8'b00000000; // 6419 :   0 - 0x0
      13'h1914: dout  = 8'b00000000; // 6420 :   0 - 0x0
      13'h1915: dout  = 8'b00000000; // 6421 :   0 - 0x0
      13'h1916: dout  = 8'b00000000; // 6422 :   0 - 0x0
      13'h1917: dout  = 8'b00000000; // 6423 :   0 - 0x0
      13'h1918: dout  = 8'b00000000; // 6424 :   0 - 0x0
      13'h1919: dout  = 8'b00000000; // 6425 :   0 - 0x0
      13'h191A: dout  = 8'b00000000; // 6426 :   0 - 0x0
      13'h191B: dout  = 8'b00000000; // 6427 :   0 - 0x0
      13'h191C: dout  = 8'b00000000; // 6428 :   0 - 0x0
      13'h191D: dout  = 8'b00000000; // 6429 :   0 - 0x0
      13'h191E: dout  = 8'b00000000; // 6430 :   0 - 0x0
      13'h191F: dout  = 8'b00000000; // 6431 :   0 - 0x0
      13'h1920: dout  = 8'b00000000; // 6432 :   0 - 0x0 -- Background 0x92
      13'h1921: dout  = 8'b00000000; // 6433 :   0 - 0x0
      13'h1922: dout  = 8'b00000000; // 6434 :   0 - 0x0
      13'h1923: dout  = 8'b00000000; // 6435 :   0 - 0x0
      13'h1924: dout  = 8'b00000000; // 6436 :   0 - 0x0
      13'h1925: dout  = 8'b00000000; // 6437 :   0 - 0x0
      13'h1926: dout  = 8'b00000000; // 6438 :   0 - 0x0
      13'h1927: dout  = 8'b00000000; // 6439 :   0 - 0x0
      13'h1928: dout  = 8'b00000000; // 6440 :   0 - 0x0
      13'h1929: dout  = 8'b00000000; // 6441 :   0 - 0x0
      13'h192A: dout  = 8'b00000000; // 6442 :   0 - 0x0
      13'h192B: dout  = 8'b00000000; // 6443 :   0 - 0x0
      13'h192C: dout  = 8'b00000000; // 6444 :   0 - 0x0
      13'h192D: dout  = 8'b00000000; // 6445 :   0 - 0x0
      13'h192E: dout  = 8'b00000000; // 6446 :   0 - 0x0
      13'h192F: dout  = 8'b00000000; // 6447 :   0 - 0x0
      13'h1930: dout  = 8'b00000000; // 6448 :   0 - 0x0 -- Background 0x93
      13'h1931: dout  = 8'b00000000; // 6449 :   0 - 0x0
      13'h1932: dout  = 8'b00000000; // 6450 :   0 - 0x0
      13'h1933: dout  = 8'b00000000; // 6451 :   0 - 0x0
      13'h1934: dout  = 8'b00000000; // 6452 :   0 - 0x0
      13'h1935: dout  = 8'b00000000; // 6453 :   0 - 0x0
      13'h1936: dout  = 8'b00000000; // 6454 :   0 - 0x0
      13'h1937: dout  = 8'b00000000; // 6455 :   0 - 0x0
      13'h1938: dout  = 8'b00000000; // 6456 :   0 - 0x0
      13'h1939: dout  = 8'b00000000; // 6457 :   0 - 0x0
      13'h193A: dout  = 8'b00000000; // 6458 :   0 - 0x0
      13'h193B: dout  = 8'b00000000; // 6459 :   0 - 0x0
      13'h193C: dout  = 8'b00000000; // 6460 :   0 - 0x0
      13'h193D: dout  = 8'b00000000; // 6461 :   0 - 0x0
      13'h193E: dout  = 8'b00000000; // 6462 :   0 - 0x0
      13'h193F: dout  = 8'b00000000; // 6463 :   0 - 0x0
      13'h1940: dout  = 8'b00000000; // 6464 :   0 - 0x0 -- Background 0x94
      13'h1941: dout  = 8'b00000000; // 6465 :   0 - 0x0
      13'h1942: dout  = 8'b00000000; // 6466 :   0 - 0x0
      13'h1943: dout  = 8'b00000000; // 6467 :   0 - 0x0
      13'h1944: dout  = 8'b00000000; // 6468 :   0 - 0x0
      13'h1945: dout  = 8'b00000000; // 6469 :   0 - 0x0
      13'h1946: dout  = 8'b00000000; // 6470 :   0 - 0x0
      13'h1947: dout  = 8'b00000000; // 6471 :   0 - 0x0
      13'h1948: dout  = 8'b00000000; // 6472 :   0 - 0x0
      13'h1949: dout  = 8'b00000000; // 6473 :   0 - 0x0
      13'h194A: dout  = 8'b00000000; // 6474 :   0 - 0x0
      13'h194B: dout  = 8'b00000000; // 6475 :   0 - 0x0
      13'h194C: dout  = 8'b00000000; // 6476 :   0 - 0x0
      13'h194D: dout  = 8'b00000000; // 6477 :   0 - 0x0
      13'h194E: dout  = 8'b00000000; // 6478 :   0 - 0x0
      13'h194F: dout  = 8'b00000000; // 6479 :   0 - 0x0
      13'h1950: dout  = 8'b00000000; // 6480 :   0 - 0x0 -- Background 0x95
      13'h1951: dout  = 8'b00000000; // 6481 :   0 - 0x0
      13'h1952: dout  = 8'b00000000; // 6482 :   0 - 0x0
      13'h1953: dout  = 8'b00000000; // 6483 :   0 - 0x0
      13'h1954: dout  = 8'b00000000; // 6484 :   0 - 0x0
      13'h1955: dout  = 8'b00000000; // 6485 :   0 - 0x0
      13'h1956: dout  = 8'b00000000; // 6486 :   0 - 0x0
      13'h1957: dout  = 8'b00000000; // 6487 :   0 - 0x0
      13'h1958: dout  = 8'b00000000; // 6488 :   0 - 0x0
      13'h1959: dout  = 8'b00000000; // 6489 :   0 - 0x0
      13'h195A: dout  = 8'b00000000; // 6490 :   0 - 0x0
      13'h195B: dout  = 8'b00000000; // 6491 :   0 - 0x0
      13'h195C: dout  = 8'b00000000; // 6492 :   0 - 0x0
      13'h195D: dout  = 8'b00000000; // 6493 :   0 - 0x0
      13'h195E: dout  = 8'b00000000; // 6494 :   0 - 0x0
      13'h195F: dout  = 8'b00000000; // 6495 :   0 - 0x0
      13'h1960: dout  = 8'b00000000; // 6496 :   0 - 0x0 -- Background 0x96
      13'h1961: dout  = 8'b00000000; // 6497 :   0 - 0x0
      13'h1962: dout  = 8'b00000000; // 6498 :   0 - 0x0
      13'h1963: dout  = 8'b00000000; // 6499 :   0 - 0x0
      13'h1964: dout  = 8'b00000000; // 6500 :   0 - 0x0
      13'h1965: dout  = 8'b00000000; // 6501 :   0 - 0x0
      13'h1966: dout  = 8'b00000000; // 6502 :   0 - 0x0
      13'h1967: dout  = 8'b00000000; // 6503 :   0 - 0x0
      13'h1968: dout  = 8'b00000000; // 6504 :   0 - 0x0
      13'h1969: dout  = 8'b00000000; // 6505 :   0 - 0x0
      13'h196A: dout  = 8'b00000000; // 6506 :   0 - 0x0
      13'h196B: dout  = 8'b00000000; // 6507 :   0 - 0x0
      13'h196C: dout  = 8'b00000000; // 6508 :   0 - 0x0
      13'h196D: dout  = 8'b00000000; // 6509 :   0 - 0x0
      13'h196E: dout  = 8'b00000000; // 6510 :   0 - 0x0
      13'h196F: dout  = 8'b00000000; // 6511 :   0 - 0x0
      13'h1970: dout  = 8'b00000000; // 6512 :   0 - 0x0 -- Background 0x97
      13'h1971: dout  = 8'b00000000; // 6513 :   0 - 0x0
      13'h1972: dout  = 8'b00000000; // 6514 :   0 - 0x0
      13'h1973: dout  = 8'b00000000; // 6515 :   0 - 0x0
      13'h1974: dout  = 8'b00000000; // 6516 :   0 - 0x0
      13'h1975: dout  = 8'b00000000; // 6517 :   0 - 0x0
      13'h1976: dout  = 8'b00000000; // 6518 :   0 - 0x0
      13'h1977: dout  = 8'b00000000; // 6519 :   0 - 0x0
      13'h1978: dout  = 8'b00000000; // 6520 :   0 - 0x0
      13'h1979: dout  = 8'b00000000; // 6521 :   0 - 0x0
      13'h197A: dout  = 8'b00000000; // 6522 :   0 - 0x0
      13'h197B: dout  = 8'b00000000; // 6523 :   0 - 0x0
      13'h197C: dout  = 8'b00000000; // 6524 :   0 - 0x0
      13'h197D: dout  = 8'b00000000; // 6525 :   0 - 0x0
      13'h197E: dout  = 8'b00000000; // 6526 :   0 - 0x0
      13'h197F: dout  = 8'b00000000; // 6527 :   0 - 0x0
      13'h1980: dout  = 8'b00000000; // 6528 :   0 - 0x0 -- Background 0x98
      13'h1981: dout  = 8'b00000000; // 6529 :   0 - 0x0
      13'h1982: dout  = 8'b00000000; // 6530 :   0 - 0x0
      13'h1983: dout  = 8'b00000000; // 6531 :   0 - 0x0
      13'h1984: dout  = 8'b00000000; // 6532 :   0 - 0x0
      13'h1985: dout  = 8'b00000000; // 6533 :   0 - 0x0
      13'h1986: dout  = 8'b00000000; // 6534 :   0 - 0x0
      13'h1987: dout  = 8'b00000000; // 6535 :   0 - 0x0
      13'h1988: dout  = 8'b00000000; // 6536 :   0 - 0x0
      13'h1989: dout  = 8'b00000000; // 6537 :   0 - 0x0
      13'h198A: dout  = 8'b00000000; // 6538 :   0 - 0x0
      13'h198B: dout  = 8'b00000000; // 6539 :   0 - 0x0
      13'h198C: dout  = 8'b00000000; // 6540 :   0 - 0x0
      13'h198D: dout  = 8'b00000000; // 6541 :   0 - 0x0
      13'h198E: dout  = 8'b00000000; // 6542 :   0 - 0x0
      13'h198F: dout  = 8'b00000000; // 6543 :   0 - 0x0
      13'h1990: dout  = 8'b00000000; // 6544 :   0 - 0x0 -- Background 0x99
      13'h1991: dout  = 8'b00000000; // 6545 :   0 - 0x0
      13'h1992: dout  = 8'b00000000; // 6546 :   0 - 0x0
      13'h1993: dout  = 8'b00000000; // 6547 :   0 - 0x0
      13'h1994: dout  = 8'b00000000; // 6548 :   0 - 0x0
      13'h1995: dout  = 8'b00000000; // 6549 :   0 - 0x0
      13'h1996: dout  = 8'b00000000; // 6550 :   0 - 0x0
      13'h1997: dout  = 8'b00000000; // 6551 :   0 - 0x0
      13'h1998: dout  = 8'b00000000; // 6552 :   0 - 0x0
      13'h1999: dout  = 8'b00000000; // 6553 :   0 - 0x0
      13'h199A: dout  = 8'b00000000; // 6554 :   0 - 0x0
      13'h199B: dout  = 8'b00000000; // 6555 :   0 - 0x0
      13'h199C: dout  = 8'b00000000; // 6556 :   0 - 0x0
      13'h199D: dout  = 8'b00000000; // 6557 :   0 - 0x0
      13'h199E: dout  = 8'b00000000; // 6558 :   0 - 0x0
      13'h199F: dout  = 8'b00000000; // 6559 :   0 - 0x0
      13'h19A0: dout  = 8'b00000000; // 6560 :   0 - 0x0 -- Background 0x9a
      13'h19A1: dout  = 8'b00000000; // 6561 :   0 - 0x0
      13'h19A2: dout  = 8'b00000000; // 6562 :   0 - 0x0
      13'h19A3: dout  = 8'b00000000; // 6563 :   0 - 0x0
      13'h19A4: dout  = 8'b00000000; // 6564 :   0 - 0x0
      13'h19A5: dout  = 8'b00000000; // 6565 :   0 - 0x0
      13'h19A6: dout  = 8'b00000000; // 6566 :   0 - 0x0
      13'h19A7: dout  = 8'b00000000; // 6567 :   0 - 0x0
      13'h19A8: dout  = 8'b00000000; // 6568 :   0 - 0x0
      13'h19A9: dout  = 8'b00000000; // 6569 :   0 - 0x0
      13'h19AA: dout  = 8'b00000000; // 6570 :   0 - 0x0
      13'h19AB: dout  = 8'b00000000; // 6571 :   0 - 0x0
      13'h19AC: dout  = 8'b00000000; // 6572 :   0 - 0x0
      13'h19AD: dout  = 8'b00000000; // 6573 :   0 - 0x0
      13'h19AE: dout  = 8'b00000000; // 6574 :   0 - 0x0
      13'h19AF: dout  = 8'b00000000; // 6575 :   0 - 0x0
      13'h19B0: dout  = 8'b00000000; // 6576 :   0 - 0x0 -- Background 0x9b
      13'h19B1: dout  = 8'b00000000; // 6577 :   0 - 0x0
      13'h19B2: dout  = 8'b00000000; // 6578 :   0 - 0x0
      13'h19B3: dout  = 8'b00000000; // 6579 :   0 - 0x0
      13'h19B4: dout  = 8'b00000000; // 6580 :   0 - 0x0
      13'h19B5: dout  = 8'b00000000; // 6581 :   0 - 0x0
      13'h19B6: dout  = 8'b00000000; // 6582 :   0 - 0x0
      13'h19B7: dout  = 8'b00000000; // 6583 :   0 - 0x0
      13'h19B8: dout  = 8'b00000000; // 6584 :   0 - 0x0
      13'h19B9: dout  = 8'b00000000; // 6585 :   0 - 0x0
      13'h19BA: dout  = 8'b00000000; // 6586 :   0 - 0x0
      13'h19BB: dout  = 8'b00000000; // 6587 :   0 - 0x0
      13'h19BC: dout  = 8'b00000000; // 6588 :   0 - 0x0
      13'h19BD: dout  = 8'b00000000; // 6589 :   0 - 0x0
      13'h19BE: dout  = 8'b00000000; // 6590 :   0 - 0x0
      13'h19BF: dout  = 8'b00000000; // 6591 :   0 - 0x0
      13'h19C0: dout  = 8'b00000000; // 6592 :   0 - 0x0 -- Background 0x9c
      13'h19C1: dout  = 8'b00000000; // 6593 :   0 - 0x0
      13'h19C2: dout  = 8'b00000000; // 6594 :   0 - 0x0
      13'h19C3: dout  = 8'b00000000; // 6595 :   0 - 0x0
      13'h19C4: dout  = 8'b00000000; // 6596 :   0 - 0x0
      13'h19C5: dout  = 8'b00000000; // 6597 :   0 - 0x0
      13'h19C6: dout  = 8'b00000000; // 6598 :   0 - 0x0
      13'h19C7: dout  = 8'b00000000; // 6599 :   0 - 0x0
      13'h19C8: dout  = 8'b00000000; // 6600 :   0 - 0x0
      13'h19C9: dout  = 8'b00000000; // 6601 :   0 - 0x0
      13'h19CA: dout  = 8'b00000000; // 6602 :   0 - 0x0
      13'h19CB: dout  = 8'b00000000; // 6603 :   0 - 0x0
      13'h19CC: dout  = 8'b00000000; // 6604 :   0 - 0x0
      13'h19CD: dout  = 8'b00000000; // 6605 :   0 - 0x0
      13'h19CE: dout  = 8'b00000000; // 6606 :   0 - 0x0
      13'h19CF: dout  = 8'b00000000; // 6607 :   0 - 0x0
      13'h19D0: dout  = 8'b00000000; // 6608 :   0 - 0x0 -- Background 0x9d
      13'h19D1: dout  = 8'b00000000; // 6609 :   0 - 0x0
      13'h19D2: dout  = 8'b00000000; // 6610 :   0 - 0x0
      13'h19D3: dout  = 8'b00000000; // 6611 :   0 - 0x0
      13'h19D4: dout  = 8'b00000000; // 6612 :   0 - 0x0
      13'h19D5: dout  = 8'b00000000; // 6613 :   0 - 0x0
      13'h19D6: dout  = 8'b00000000; // 6614 :   0 - 0x0
      13'h19D7: dout  = 8'b00000000; // 6615 :   0 - 0x0
      13'h19D8: dout  = 8'b00000000; // 6616 :   0 - 0x0
      13'h19D9: dout  = 8'b00000000; // 6617 :   0 - 0x0
      13'h19DA: dout  = 8'b00000000; // 6618 :   0 - 0x0
      13'h19DB: dout  = 8'b00000000; // 6619 :   0 - 0x0
      13'h19DC: dout  = 8'b00000000; // 6620 :   0 - 0x0
      13'h19DD: dout  = 8'b00000000; // 6621 :   0 - 0x0
      13'h19DE: dout  = 8'b00000000; // 6622 :   0 - 0x0
      13'h19DF: dout  = 8'b00000000; // 6623 :   0 - 0x0
      13'h19E0: dout  = 8'b00000000; // 6624 :   0 - 0x0 -- Background 0x9e
      13'h19E1: dout  = 8'b00000000; // 6625 :   0 - 0x0
      13'h19E2: dout  = 8'b00000000; // 6626 :   0 - 0x0
      13'h19E3: dout  = 8'b00000000; // 6627 :   0 - 0x0
      13'h19E4: dout  = 8'b00000000; // 6628 :   0 - 0x0
      13'h19E5: dout  = 8'b00000000; // 6629 :   0 - 0x0
      13'h19E6: dout  = 8'b00000000; // 6630 :   0 - 0x0
      13'h19E7: dout  = 8'b00000000; // 6631 :   0 - 0x0
      13'h19E8: dout  = 8'b00000000; // 6632 :   0 - 0x0
      13'h19E9: dout  = 8'b00000000; // 6633 :   0 - 0x0
      13'h19EA: dout  = 8'b00000000; // 6634 :   0 - 0x0
      13'h19EB: dout  = 8'b00000000; // 6635 :   0 - 0x0
      13'h19EC: dout  = 8'b00000000; // 6636 :   0 - 0x0
      13'h19ED: dout  = 8'b00000000; // 6637 :   0 - 0x0
      13'h19EE: dout  = 8'b00000000; // 6638 :   0 - 0x0
      13'h19EF: dout  = 8'b00000000; // 6639 :   0 - 0x0
      13'h19F0: dout  = 8'b00000000; // 6640 :   0 - 0x0 -- Background 0x9f
      13'h19F1: dout  = 8'b00000000; // 6641 :   0 - 0x0
      13'h19F2: dout  = 8'b00000000; // 6642 :   0 - 0x0
      13'h19F3: dout  = 8'b00000000; // 6643 :   0 - 0x0
      13'h19F4: dout  = 8'b00000000; // 6644 :   0 - 0x0
      13'h19F5: dout  = 8'b00000000; // 6645 :   0 - 0x0
      13'h19F6: dout  = 8'b00000000; // 6646 :   0 - 0x0
      13'h19F7: dout  = 8'b00000000; // 6647 :   0 - 0x0
      13'h19F8: dout  = 8'b00000000; // 6648 :   0 - 0x0
      13'h19F9: dout  = 8'b00000000; // 6649 :   0 - 0x0
      13'h19FA: dout  = 8'b00000000; // 6650 :   0 - 0x0
      13'h19FB: dout  = 8'b00000000; // 6651 :   0 - 0x0
      13'h19FC: dout  = 8'b00000000; // 6652 :   0 - 0x0
      13'h19FD: dout  = 8'b00000000; // 6653 :   0 - 0x0
      13'h19FE: dout  = 8'b00000000; // 6654 :   0 - 0x0
      13'h19FF: dout  = 8'b00000000; // 6655 :   0 - 0x0
      13'h1A00: dout  = 8'b00000000; // 6656 :   0 - 0x0 -- Background 0xa0
      13'h1A01: dout  = 8'b00000000; // 6657 :   0 - 0x0
      13'h1A02: dout  = 8'b00000000; // 6658 :   0 - 0x0
      13'h1A03: dout  = 8'b00000000; // 6659 :   0 - 0x0
      13'h1A04: dout  = 8'b00000000; // 6660 :   0 - 0x0
      13'h1A05: dout  = 8'b00000000; // 6661 :   0 - 0x0
      13'h1A06: dout  = 8'b00000000; // 6662 :   0 - 0x0
      13'h1A07: dout  = 8'b00000000; // 6663 :   0 - 0x0
      13'h1A08: dout  = 8'b00000000; // 6664 :   0 - 0x0
      13'h1A09: dout  = 8'b00000000; // 6665 :   0 - 0x0
      13'h1A0A: dout  = 8'b00000000; // 6666 :   0 - 0x0
      13'h1A0B: dout  = 8'b00000000; // 6667 :   0 - 0x0
      13'h1A0C: dout  = 8'b00000000; // 6668 :   0 - 0x0
      13'h1A0D: dout  = 8'b00000000; // 6669 :   0 - 0x0
      13'h1A0E: dout  = 8'b00000000; // 6670 :   0 - 0x0
      13'h1A0F: dout  = 8'b00000000; // 6671 :   0 - 0x0
      13'h1A10: dout  = 8'b00000000; // 6672 :   0 - 0x0 -- Background 0xa1
      13'h1A11: dout  = 8'b00000000; // 6673 :   0 - 0x0
      13'h1A12: dout  = 8'b00000000; // 6674 :   0 - 0x0
      13'h1A13: dout  = 8'b00000000; // 6675 :   0 - 0x0
      13'h1A14: dout  = 8'b00000000; // 6676 :   0 - 0x0
      13'h1A15: dout  = 8'b00000000; // 6677 :   0 - 0x0
      13'h1A16: dout  = 8'b00000000; // 6678 :   0 - 0x0
      13'h1A17: dout  = 8'b00000000; // 6679 :   0 - 0x0
      13'h1A18: dout  = 8'b00000000; // 6680 :   0 - 0x0
      13'h1A19: dout  = 8'b00000000; // 6681 :   0 - 0x0
      13'h1A1A: dout  = 8'b00000000; // 6682 :   0 - 0x0
      13'h1A1B: dout  = 8'b00000000; // 6683 :   0 - 0x0
      13'h1A1C: dout  = 8'b00000000; // 6684 :   0 - 0x0
      13'h1A1D: dout  = 8'b00000000; // 6685 :   0 - 0x0
      13'h1A1E: dout  = 8'b00000000; // 6686 :   0 - 0x0
      13'h1A1F: dout  = 8'b00000000; // 6687 :   0 - 0x0
      13'h1A20: dout  = 8'b00000000; // 6688 :   0 - 0x0 -- Background 0xa2
      13'h1A21: dout  = 8'b00000000; // 6689 :   0 - 0x0
      13'h1A22: dout  = 8'b00000000; // 6690 :   0 - 0x0
      13'h1A23: dout  = 8'b00000000; // 6691 :   0 - 0x0
      13'h1A24: dout  = 8'b00000000; // 6692 :   0 - 0x0
      13'h1A25: dout  = 8'b00000000; // 6693 :   0 - 0x0
      13'h1A26: dout  = 8'b00000000; // 6694 :   0 - 0x0
      13'h1A27: dout  = 8'b00000000; // 6695 :   0 - 0x0
      13'h1A28: dout  = 8'b00000000; // 6696 :   0 - 0x0
      13'h1A29: dout  = 8'b00000000; // 6697 :   0 - 0x0
      13'h1A2A: dout  = 8'b00000000; // 6698 :   0 - 0x0
      13'h1A2B: dout  = 8'b00000000; // 6699 :   0 - 0x0
      13'h1A2C: dout  = 8'b00000000; // 6700 :   0 - 0x0
      13'h1A2D: dout  = 8'b00000000; // 6701 :   0 - 0x0
      13'h1A2E: dout  = 8'b00000000; // 6702 :   0 - 0x0
      13'h1A2F: dout  = 8'b00000000; // 6703 :   0 - 0x0
      13'h1A30: dout  = 8'b00000000; // 6704 :   0 - 0x0 -- Background 0xa3
      13'h1A31: dout  = 8'b00000000; // 6705 :   0 - 0x0
      13'h1A32: dout  = 8'b00000000; // 6706 :   0 - 0x0
      13'h1A33: dout  = 8'b00000000; // 6707 :   0 - 0x0
      13'h1A34: dout  = 8'b00000000; // 6708 :   0 - 0x0
      13'h1A35: dout  = 8'b00000000; // 6709 :   0 - 0x0
      13'h1A36: dout  = 8'b00000000; // 6710 :   0 - 0x0
      13'h1A37: dout  = 8'b00000000; // 6711 :   0 - 0x0
      13'h1A38: dout  = 8'b00000000; // 6712 :   0 - 0x0
      13'h1A39: dout  = 8'b00000000; // 6713 :   0 - 0x0
      13'h1A3A: dout  = 8'b00000000; // 6714 :   0 - 0x0
      13'h1A3B: dout  = 8'b00000000; // 6715 :   0 - 0x0
      13'h1A3C: dout  = 8'b00000000; // 6716 :   0 - 0x0
      13'h1A3D: dout  = 8'b00000000; // 6717 :   0 - 0x0
      13'h1A3E: dout  = 8'b00000000; // 6718 :   0 - 0x0
      13'h1A3F: dout  = 8'b00000000; // 6719 :   0 - 0x0
      13'h1A40: dout  = 8'b00000000; // 6720 :   0 - 0x0 -- Background 0xa4
      13'h1A41: dout  = 8'b00000000; // 6721 :   0 - 0x0
      13'h1A42: dout  = 8'b00000000; // 6722 :   0 - 0x0
      13'h1A43: dout  = 8'b00000000; // 6723 :   0 - 0x0
      13'h1A44: dout  = 8'b00000000; // 6724 :   0 - 0x0
      13'h1A45: dout  = 8'b00000000; // 6725 :   0 - 0x0
      13'h1A46: dout  = 8'b00000000; // 6726 :   0 - 0x0
      13'h1A47: dout  = 8'b00000000; // 6727 :   0 - 0x0
      13'h1A48: dout  = 8'b00000000; // 6728 :   0 - 0x0
      13'h1A49: dout  = 8'b00000000; // 6729 :   0 - 0x0
      13'h1A4A: dout  = 8'b00000000; // 6730 :   0 - 0x0
      13'h1A4B: dout  = 8'b00000000; // 6731 :   0 - 0x0
      13'h1A4C: dout  = 8'b00000000; // 6732 :   0 - 0x0
      13'h1A4D: dout  = 8'b00000000; // 6733 :   0 - 0x0
      13'h1A4E: dout  = 8'b00000000; // 6734 :   0 - 0x0
      13'h1A4F: dout  = 8'b00000000; // 6735 :   0 - 0x0
      13'h1A50: dout  = 8'b00000000; // 6736 :   0 - 0x0 -- Background 0xa5
      13'h1A51: dout  = 8'b00000000; // 6737 :   0 - 0x0
      13'h1A52: dout  = 8'b00000000; // 6738 :   0 - 0x0
      13'h1A53: dout  = 8'b00000000; // 6739 :   0 - 0x0
      13'h1A54: dout  = 8'b00000000; // 6740 :   0 - 0x0
      13'h1A55: dout  = 8'b00000000; // 6741 :   0 - 0x0
      13'h1A56: dout  = 8'b00000000; // 6742 :   0 - 0x0
      13'h1A57: dout  = 8'b00000000; // 6743 :   0 - 0x0
      13'h1A58: dout  = 8'b00000000; // 6744 :   0 - 0x0
      13'h1A59: dout  = 8'b00000000; // 6745 :   0 - 0x0
      13'h1A5A: dout  = 8'b00000000; // 6746 :   0 - 0x0
      13'h1A5B: dout  = 8'b00000000; // 6747 :   0 - 0x0
      13'h1A5C: dout  = 8'b00000000; // 6748 :   0 - 0x0
      13'h1A5D: dout  = 8'b00000000; // 6749 :   0 - 0x0
      13'h1A5E: dout  = 8'b00000000; // 6750 :   0 - 0x0
      13'h1A5F: dout  = 8'b00000000; // 6751 :   0 - 0x0
      13'h1A60: dout  = 8'b00000000; // 6752 :   0 - 0x0 -- Background 0xa6
      13'h1A61: dout  = 8'b00000000; // 6753 :   0 - 0x0
      13'h1A62: dout  = 8'b00000000; // 6754 :   0 - 0x0
      13'h1A63: dout  = 8'b00000000; // 6755 :   0 - 0x0
      13'h1A64: dout  = 8'b00000000; // 6756 :   0 - 0x0
      13'h1A65: dout  = 8'b00000000; // 6757 :   0 - 0x0
      13'h1A66: dout  = 8'b00000000; // 6758 :   0 - 0x0
      13'h1A67: dout  = 8'b00000000; // 6759 :   0 - 0x0
      13'h1A68: dout  = 8'b00000000; // 6760 :   0 - 0x0
      13'h1A69: dout  = 8'b00000000; // 6761 :   0 - 0x0
      13'h1A6A: dout  = 8'b00000000; // 6762 :   0 - 0x0
      13'h1A6B: dout  = 8'b00000000; // 6763 :   0 - 0x0
      13'h1A6C: dout  = 8'b00000000; // 6764 :   0 - 0x0
      13'h1A6D: dout  = 8'b00000000; // 6765 :   0 - 0x0
      13'h1A6E: dout  = 8'b00000000; // 6766 :   0 - 0x0
      13'h1A6F: dout  = 8'b00000000; // 6767 :   0 - 0x0
      13'h1A70: dout  = 8'b00000000; // 6768 :   0 - 0x0 -- Background 0xa7
      13'h1A71: dout  = 8'b00000000; // 6769 :   0 - 0x0
      13'h1A72: dout  = 8'b00000000; // 6770 :   0 - 0x0
      13'h1A73: dout  = 8'b00000000; // 6771 :   0 - 0x0
      13'h1A74: dout  = 8'b00000000; // 6772 :   0 - 0x0
      13'h1A75: dout  = 8'b00000000; // 6773 :   0 - 0x0
      13'h1A76: dout  = 8'b00000000; // 6774 :   0 - 0x0
      13'h1A77: dout  = 8'b00000000; // 6775 :   0 - 0x0
      13'h1A78: dout  = 8'b00000000; // 6776 :   0 - 0x0
      13'h1A79: dout  = 8'b00000000; // 6777 :   0 - 0x0
      13'h1A7A: dout  = 8'b00000000; // 6778 :   0 - 0x0
      13'h1A7B: dout  = 8'b00000000; // 6779 :   0 - 0x0
      13'h1A7C: dout  = 8'b00000000; // 6780 :   0 - 0x0
      13'h1A7D: dout  = 8'b00000000; // 6781 :   0 - 0x0
      13'h1A7E: dout  = 8'b00000000; // 6782 :   0 - 0x0
      13'h1A7F: dout  = 8'b00000000; // 6783 :   0 - 0x0
      13'h1A80: dout  = 8'b00000000; // 6784 :   0 - 0x0 -- Background 0xa8
      13'h1A81: dout  = 8'b00000000; // 6785 :   0 - 0x0
      13'h1A82: dout  = 8'b00000000; // 6786 :   0 - 0x0
      13'h1A83: dout  = 8'b00000000; // 6787 :   0 - 0x0
      13'h1A84: dout  = 8'b00000000; // 6788 :   0 - 0x0
      13'h1A85: dout  = 8'b00000000; // 6789 :   0 - 0x0
      13'h1A86: dout  = 8'b00000000; // 6790 :   0 - 0x0
      13'h1A87: dout  = 8'b00000000; // 6791 :   0 - 0x0
      13'h1A88: dout  = 8'b00000000; // 6792 :   0 - 0x0
      13'h1A89: dout  = 8'b00000000; // 6793 :   0 - 0x0
      13'h1A8A: dout  = 8'b00000000; // 6794 :   0 - 0x0
      13'h1A8B: dout  = 8'b00000000; // 6795 :   0 - 0x0
      13'h1A8C: dout  = 8'b00000000; // 6796 :   0 - 0x0
      13'h1A8D: dout  = 8'b00000000; // 6797 :   0 - 0x0
      13'h1A8E: dout  = 8'b00000000; // 6798 :   0 - 0x0
      13'h1A8F: dout  = 8'b00000000; // 6799 :   0 - 0x0
      13'h1A90: dout  = 8'b00000000; // 6800 :   0 - 0x0 -- Background 0xa9
      13'h1A91: dout  = 8'b00000000; // 6801 :   0 - 0x0
      13'h1A92: dout  = 8'b00000000; // 6802 :   0 - 0x0
      13'h1A93: dout  = 8'b00000000; // 6803 :   0 - 0x0
      13'h1A94: dout  = 8'b00000000; // 6804 :   0 - 0x0
      13'h1A95: dout  = 8'b00000000; // 6805 :   0 - 0x0
      13'h1A96: dout  = 8'b00000000; // 6806 :   0 - 0x0
      13'h1A97: dout  = 8'b00000000; // 6807 :   0 - 0x0
      13'h1A98: dout  = 8'b00000000; // 6808 :   0 - 0x0
      13'h1A99: dout  = 8'b00000000; // 6809 :   0 - 0x0
      13'h1A9A: dout  = 8'b00000000; // 6810 :   0 - 0x0
      13'h1A9B: dout  = 8'b00000000; // 6811 :   0 - 0x0
      13'h1A9C: dout  = 8'b00000000; // 6812 :   0 - 0x0
      13'h1A9D: dout  = 8'b00000000; // 6813 :   0 - 0x0
      13'h1A9E: dout  = 8'b00000000; // 6814 :   0 - 0x0
      13'h1A9F: dout  = 8'b00000000; // 6815 :   0 - 0x0
      13'h1AA0: dout  = 8'b00000000; // 6816 :   0 - 0x0 -- Background 0xaa
      13'h1AA1: dout  = 8'b00000000; // 6817 :   0 - 0x0
      13'h1AA2: dout  = 8'b00000000; // 6818 :   0 - 0x0
      13'h1AA3: dout  = 8'b00000000; // 6819 :   0 - 0x0
      13'h1AA4: dout  = 8'b00000000; // 6820 :   0 - 0x0
      13'h1AA5: dout  = 8'b00000000; // 6821 :   0 - 0x0
      13'h1AA6: dout  = 8'b00000000; // 6822 :   0 - 0x0
      13'h1AA7: dout  = 8'b00000000; // 6823 :   0 - 0x0
      13'h1AA8: dout  = 8'b00000000; // 6824 :   0 - 0x0
      13'h1AA9: dout  = 8'b00000000; // 6825 :   0 - 0x0
      13'h1AAA: dout  = 8'b00000000; // 6826 :   0 - 0x0
      13'h1AAB: dout  = 8'b00000000; // 6827 :   0 - 0x0
      13'h1AAC: dout  = 8'b00000000; // 6828 :   0 - 0x0
      13'h1AAD: dout  = 8'b00000000; // 6829 :   0 - 0x0
      13'h1AAE: dout  = 8'b00000000; // 6830 :   0 - 0x0
      13'h1AAF: dout  = 8'b00000000; // 6831 :   0 - 0x0
      13'h1AB0: dout  = 8'b00000000; // 6832 :   0 - 0x0 -- Background 0xab
      13'h1AB1: dout  = 8'b00000000; // 6833 :   0 - 0x0
      13'h1AB2: dout  = 8'b00000000; // 6834 :   0 - 0x0
      13'h1AB3: dout  = 8'b00000000; // 6835 :   0 - 0x0
      13'h1AB4: dout  = 8'b00000000; // 6836 :   0 - 0x0
      13'h1AB5: dout  = 8'b00000000; // 6837 :   0 - 0x0
      13'h1AB6: dout  = 8'b00000000; // 6838 :   0 - 0x0
      13'h1AB7: dout  = 8'b00000000; // 6839 :   0 - 0x0
      13'h1AB8: dout  = 8'b00000000; // 6840 :   0 - 0x0
      13'h1AB9: dout  = 8'b00000000; // 6841 :   0 - 0x0
      13'h1ABA: dout  = 8'b00000000; // 6842 :   0 - 0x0
      13'h1ABB: dout  = 8'b00000000; // 6843 :   0 - 0x0
      13'h1ABC: dout  = 8'b00000000; // 6844 :   0 - 0x0
      13'h1ABD: dout  = 8'b00000000; // 6845 :   0 - 0x0
      13'h1ABE: dout  = 8'b00000000; // 6846 :   0 - 0x0
      13'h1ABF: dout  = 8'b00000000; // 6847 :   0 - 0x0
      13'h1AC0: dout  = 8'b00000000; // 6848 :   0 - 0x0 -- Background 0xac
      13'h1AC1: dout  = 8'b00000000; // 6849 :   0 - 0x0
      13'h1AC2: dout  = 8'b00000000; // 6850 :   0 - 0x0
      13'h1AC3: dout  = 8'b00000000; // 6851 :   0 - 0x0
      13'h1AC4: dout  = 8'b00000000; // 6852 :   0 - 0x0
      13'h1AC5: dout  = 8'b00000000; // 6853 :   0 - 0x0
      13'h1AC6: dout  = 8'b00000000; // 6854 :   0 - 0x0
      13'h1AC7: dout  = 8'b00000000; // 6855 :   0 - 0x0
      13'h1AC8: dout  = 8'b00000000; // 6856 :   0 - 0x0
      13'h1AC9: dout  = 8'b00000000; // 6857 :   0 - 0x0
      13'h1ACA: dout  = 8'b00000000; // 6858 :   0 - 0x0
      13'h1ACB: dout  = 8'b00000000; // 6859 :   0 - 0x0
      13'h1ACC: dout  = 8'b00000000; // 6860 :   0 - 0x0
      13'h1ACD: dout  = 8'b00000000; // 6861 :   0 - 0x0
      13'h1ACE: dout  = 8'b00000000; // 6862 :   0 - 0x0
      13'h1ACF: dout  = 8'b00000000; // 6863 :   0 - 0x0
      13'h1AD0: dout  = 8'b00000000; // 6864 :   0 - 0x0 -- Background 0xad
      13'h1AD1: dout  = 8'b00000000; // 6865 :   0 - 0x0
      13'h1AD2: dout  = 8'b00000000; // 6866 :   0 - 0x0
      13'h1AD3: dout  = 8'b00000000; // 6867 :   0 - 0x0
      13'h1AD4: dout  = 8'b00000000; // 6868 :   0 - 0x0
      13'h1AD5: dout  = 8'b00000000; // 6869 :   0 - 0x0
      13'h1AD6: dout  = 8'b00000000; // 6870 :   0 - 0x0
      13'h1AD7: dout  = 8'b00000000; // 6871 :   0 - 0x0
      13'h1AD8: dout  = 8'b00000000; // 6872 :   0 - 0x0
      13'h1AD9: dout  = 8'b00000000; // 6873 :   0 - 0x0
      13'h1ADA: dout  = 8'b00000000; // 6874 :   0 - 0x0
      13'h1ADB: dout  = 8'b00000000; // 6875 :   0 - 0x0
      13'h1ADC: dout  = 8'b00000000; // 6876 :   0 - 0x0
      13'h1ADD: dout  = 8'b00000000; // 6877 :   0 - 0x0
      13'h1ADE: dout  = 8'b00000000; // 6878 :   0 - 0x0
      13'h1ADF: dout  = 8'b00000000; // 6879 :   0 - 0x0
      13'h1AE0: dout  = 8'b00000000; // 6880 :   0 - 0x0 -- Background 0xae
      13'h1AE1: dout  = 8'b00000000; // 6881 :   0 - 0x0
      13'h1AE2: dout  = 8'b00000000; // 6882 :   0 - 0x0
      13'h1AE3: dout  = 8'b00000000; // 6883 :   0 - 0x0
      13'h1AE4: dout  = 8'b00000000; // 6884 :   0 - 0x0
      13'h1AE5: dout  = 8'b00000000; // 6885 :   0 - 0x0
      13'h1AE6: dout  = 8'b00000000; // 6886 :   0 - 0x0
      13'h1AE7: dout  = 8'b00000000; // 6887 :   0 - 0x0
      13'h1AE8: dout  = 8'b00000000; // 6888 :   0 - 0x0
      13'h1AE9: dout  = 8'b00000000; // 6889 :   0 - 0x0
      13'h1AEA: dout  = 8'b00000000; // 6890 :   0 - 0x0
      13'h1AEB: dout  = 8'b00000000; // 6891 :   0 - 0x0
      13'h1AEC: dout  = 8'b00000000; // 6892 :   0 - 0x0
      13'h1AED: dout  = 8'b00000000; // 6893 :   0 - 0x0
      13'h1AEE: dout  = 8'b00000000; // 6894 :   0 - 0x0
      13'h1AEF: dout  = 8'b00000000; // 6895 :   0 - 0x0
      13'h1AF0: dout  = 8'b00000000; // 6896 :   0 - 0x0 -- Background 0xaf
      13'h1AF1: dout  = 8'b00000000; // 6897 :   0 - 0x0
      13'h1AF2: dout  = 8'b00000000; // 6898 :   0 - 0x0
      13'h1AF3: dout  = 8'b00000000; // 6899 :   0 - 0x0
      13'h1AF4: dout  = 8'b00000000; // 6900 :   0 - 0x0
      13'h1AF5: dout  = 8'b00000000; // 6901 :   0 - 0x0
      13'h1AF6: dout  = 8'b00000000; // 6902 :   0 - 0x0
      13'h1AF7: dout  = 8'b00000000; // 6903 :   0 - 0x0
      13'h1AF8: dout  = 8'b00000000; // 6904 :   0 - 0x0
      13'h1AF9: dout  = 8'b00000000; // 6905 :   0 - 0x0
      13'h1AFA: dout  = 8'b00000000; // 6906 :   0 - 0x0
      13'h1AFB: dout  = 8'b00000000; // 6907 :   0 - 0x0
      13'h1AFC: dout  = 8'b00000000; // 6908 :   0 - 0x0
      13'h1AFD: dout  = 8'b00000000; // 6909 :   0 - 0x0
      13'h1AFE: dout  = 8'b00000000; // 6910 :   0 - 0x0
      13'h1AFF: dout  = 8'b00000000; // 6911 :   0 - 0x0
      13'h1B00: dout  = 8'b00000000; // 6912 :   0 - 0x0 -- Background 0xb0
      13'h1B01: dout  = 8'b00000000; // 6913 :   0 - 0x0
      13'h1B02: dout  = 8'b00000000; // 6914 :   0 - 0x0
      13'h1B03: dout  = 8'b00000000; // 6915 :   0 - 0x0
      13'h1B04: dout  = 8'b00000000; // 6916 :   0 - 0x0
      13'h1B05: dout  = 8'b00000000; // 6917 :   0 - 0x0
      13'h1B06: dout  = 8'b00000000; // 6918 :   0 - 0x0
      13'h1B07: dout  = 8'b00000000; // 6919 :   0 - 0x0
      13'h1B08: dout  = 8'b00000000; // 6920 :   0 - 0x0
      13'h1B09: dout  = 8'b00000000; // 6921 :   0 - 0x0
      13'h1B0A: dout  = 8'b00000000; // 6922 :   0 - 0x0
      13'h1B0B: dout  = 8'b00000000; // 6923 :   0 - 0x0
      13'h1B0C: dout  = 8'b00000000; // 6924 :   0 - 0x0
      13'h1B0D: dout  = 8'b00000000; // 6925 :   0 - 0x0
      13'h1B0E: dout  = 8'b00000000; // 6926 :   0 - 0x0
      13'h1B0F: dout  = 8'b00000000; // 6927 :   0 - 0x0
      13'h1B10: dout  = 8'b00000000; // 6928 :   0 - 0x0 -- Background 0xb1
      13'h1B11: dout  = 8'b00000000; // 6929 :   0 - 0x0
      13'h1B12: dout  = 8'b00000000; // 6930 :   0 - 0x0
      13'h1B13: dout  = 8'b00000000; // 6931 :   0 - 0x0
      13'h1B14: dout  = 8'b00000000; // 6932 :   0 - 0x0
      13'h1B15: dout  = 8'b00000000; // 6933 :   0 - 0x0
      13'h1B16: dout  = 8'b00000000; // 6934 :   0 - 0x0
      13'h1B17: dout  = 8'b00000000; // 6935 :   0 - 0x0
      13'h1B18: dout  = 8'b00000000; // 6936 :   0 - 0x0
      13'h1B19: dout  = 8'b00000000; // 6937 :   0 - 0x0
      13'h1B1A: dout  = 8'b00000000; // 6938 :   0 - 0x0
      13'h1B1B: dout  = 8'b00000000; // 6939 :   0 - 0x0
      13'h1B1C: dout  = 8'b00000000; // 6940 :   0 - 0x0
      13'h1B1D: dout  = 8'b00000000; // 6941 :   0 - 0x0
      13'h1B1E: dout  = 8'b00000000; // 6942 :   0 - 0x0
      13'h1B1F: dout  = 8'b00000000; // 6943 :   0 - 0x0
      13'h1B20: dout  = 8'b00000000; // 6944 :   0 - 0x0 -- Background 0xb2
      13'h1B21: dout  = 8'b00000000; // 6945 :   0 - 0x0
      13'h1B22: dout  = 8'b00000000; // 6946 :   0 - 0x0
      13'h1B23: dout  = 8'b00000000; // 6947 :   0 - 0x0
      13'h1B24: dout  = 8'b00000000; // 6948 :   0 - 0x0
      13'h1B25: dout  = 8'b00000000; // 6949 :   0 - 0x0
      13'h1B26: dout  = 8'b00000000; // 6950 :   0 - 0x0
      13'h1B27: dout  = 8'b00000000; // 6951 :   0 - 0x0
      13'h1B28: dout  = 8'b00000000; // 6952 :   0 - 0x0
      13'h1B29: dout  = 8'b00000000; // 6953 :   0 - 0x0
      13'h1B2A: dout  = 8'b00000000; // 6954 :   0 - 0x0
      13'h1B2B: dout  = 8'b00000000; // 6955 :   0 - 0x0
      13'h1B2C: dout  = 8'b00000000; // 6956 :   0 - 0x0
      13'h1B2D: dout  = 8'b00000000; // 6957 :   0 - 0x0
      13'h1B2E: dout  = 8'b00000000; // 6958 :   0 - 0x0
      13'h1B2F: dout  = 8'b00000000; // 6959 :   0 - 0x0
      13'h1B30: dout  = 8'b00000000; // 6960 :   0 - 0x0 -- Background 0xb3
      13'h1B31: dout  = 8'b00000000; // 6961 :   0 - 0x0
      13'h1B32: dout  = 8'b00000000; // 6962 :   0 - 0x0
      13'h1B33: dout  = 8'b00000000; // 6963 :   0 - 0x0
      13'h1B34: dout  = 8'b00000000; // 6964 :   0 - 0x0
      13'h1B35: dout  = 8'b00000000; // 6965 :   0 - 0x0
      13'h1B36: dout  = 8'b00000000; // 6966 :   0 - 0x0
      13'h1B37: dout  = 8'b00000000; // 6967 :   0 - 0x0
      13'h1B38: dout  = 8'b00000000; // 6968 :   0 - 0x0
      13'h1B39: dout  = 8'b00000000; // 6969 :   0 - 0x0
      13'h1B3A: dout  = 8'b00000000; // 6970 :   0 - 0x0
      13'h1B3B: dout  = 8'b00000000; // 6971 :   0 - 0x0
      13'h1B3C: dout  = 8'b00000000; // 6972 :   0 - 0x0
      13'h1B3D: dout  = 8'b00000000; // 6973 :   0 - 0x0
      13'h1B3E: dout  = 8'b00000000; // 6974 :   0 - 0x0
      13'h1B3F: dout  = 8'b00000000; // 6975 :   0 - 0x0
      13'h1B40: dout  = 8'b00000000; // 6976 :   0 - 0x0 -- Background 0xb4
      13'h1B41: dout  = 8'b00000000; // 6977 :   0 - 0x0
      13'h1B42: dout  = 8'b00000000; // 6978 :   0 - 0x0
      13'h1B43: dout  = 8'b00000000; // 6979 :   0 - 0x0
      13'h1B44: dout  = 8'b00000000; // 6980 :   0 - 0x0
      13'h1B45: dout  = 8'b00000000; // 6981 :   0 - 0x0
      13'h1B46: dout  = 8'b00000000; // 6982 :   0 - 0x0
      13'h1B47: dout  = 8'b00000000; // 6983 :   0 - 0x0
      13'h1B48: dout  = 8'b00000000; // 6984 :   0 - 0x0
      13'h1B49: dout  = 8'b00000000; // 6985 :   0 - 0x0
      13'h1B4A: dout  = 8'b00000000; // 6986 :   0 - 0x0
      13'h1B4B: dout  = 8'b00000000; // 6987 :   0 - 0x0
      13'h1B4C: dout  = 8'b00000000; // 6988 :   0 - 0x0
      13'h1B4D: dout  = 8'b00000000; // 6989 :   0 - 0x0
      13'h1B4E: dout  = 8'b00000000; // 6990 :   0 - 0x0
      13'h1B4F: dout  = 8'b00000000; // 6991 :   0 - 0x0
      13'h1B50: dout  = 8'b00000000; // 6992 :   0 - 0x0 -- Background 0xb5
      13'h1B51: dout  = 8'b00000000; // 6993 :   0 - 0x0
      13'h1B52: dout  = 8'b00000000; // 6994 :   0 - 0x0
      13'h1B53: dout  = 8'b00000000; // 6995 :   0 - 0x0
      13'h1B54: dout  = 8'b00000000; // 6996 :   0 - 0x0
      13'h1B55: dout  = 8'b00000000; // 6997 :   0 - 0x0
      13'h1B56: dout  = 8'b00000000; // 6998 :   0 - 0x0
      13'h1B57: dout  = 8'b00000000; // 6999 :   0 - 0x0
      13'h1B58: dout  = 8'b00000000; // 7000 :   0 - 0x0
      13'h1B59: dout  = 8'b00000000; // 7001 :   0 - 0x0
      13'h1B5A: dout  = 8'b00000000; // 7002 :   0 - 0x0
      13'h1B5B: dout  = 8'b00000000; // 7003 :   0 - 0x0
      13'h1B5C: dout  = 8'b00000000; // 7004 :   0 - 0x0
      13'h1B5D: dout  = 8'b00000000; // 7005 :   0 - 0x0
      13'h1B5E: dout  = 8'b00000000; // 7006 :   0 - 0x0
      13'h1B5F: dout  = 8'b00000000; // 7007 :   0 - 0x0
      13'h1B60: dout  = 8'b00000000; // 7008 :   0 - 0x0 -- Background 0xb6
      13'h1B61: dout  = 8'b00000000; // 7009 :   0 - 0x0
      13'h1B62: dout  = 8'b00000000; // 7010 :   0 - 0x0
      13'h1B63: dout  = 8'b00000000; // 7011 :   0 - 0x0
      13'h1B64: dout  = 8'b00000000; // 7012 :   0 - 0x0
      13'h1B65: dout  = 8'b00000000; // 7013 :   0 - 0x0
      13'h1B66: dout  = 8'b00000000; // 7014 :   0 - 0x0
      13'h1B67: dout  = 8'b00000000; // 7015 :   0 - 0x0
      13'h1B68: dout  = 8'b00000000; // 7016 :   0 - 0x0
      13'h1B69: dout  = 8'b00000000; // 7017 :   0 - 0x0
      13'h1B6A: dout  = 8'b00000000; // 7018 :   0 - 0x0
      13'h1B6B: dout  = 8'b00000000; // 7019 :   0 - 0x0
      13'h1B6C: dout  = 8'b00000000; // 7020 :   0 - 0x0
      13'h1B6D: dout  = 8'b00000000; // 7021 :   0 - 0x0
      13'h1B6E: dout  = 8'b00000000; // 7022 :   0 - 0x0
      13'h1B6F: dout  = 8'b00000000; // 7023 :   0 - 0x0
      13'h1B70: dout  = 8'b00000000; // 7024 :   0 - 0x0 -- Background 0xb7
      13'h1B71: dout  = 8'b00000000; // 7025 :   0 - 0x0
      13'h1B72: dout  = 8'b00000000; // 7026 :   0 - 0x0
      13'h1B73: dout  = 8'b00000000; // 7027 :   0 - 0x0
      13'h1B74: dout  = 8'b00000000; // 7028 :   0 - 0x0
      13'h1B75: dout  = 8'b00000000; // 7029 :   0 - 0x0
      13'h1B76: dout  = 8'b00000000; // 7030 :   0 - 0x0
      13'h1B77: dout  = 8'b00000000; // 7031 :   0 - 0x0
      13'h1B78: dout  = 8'b00000000; // 7032 :   0 - 0x0
      13'h1B79: dout  = 8'b00000000; // 7033 :   0 - 0x0
      13'h1B7A: dout  = 8'b00000000; // 7034 :   0 - 0x0
      13'h1B7B: dout  = 8'b00000000; // 7035 :   0 - 0x0
      13'h1B7C: dout  = 8'b00000000; // 7036 :   0 - 0x0
      13'h1B7D: dout  = 8'b00000000; // 7037 :   0 - 0x0
      13'h1B7E: dout  = 8'b00000000; // 7038 :   0 - 0x0
      13'h1B7F: dout  = 8'b00000000; // 7039 :   0 - 0x0
      13'h1B80: dout  = 8'b00000000; // 7040 :   0 - 0x0 -- Background 0xb8
      13'h1B81: dout  = 8'b00000000; // 7041 :   0 - 0x0
      13'h1B82: dout  = 8'b00000000; // 7042 :   0 - 0x0
      13'h1B83: dout  = 8'b00000000; // 7043 :   0 - 0x0
      13'h1B84: dout  = 8'b00000000; // 7044 :   0 - 0x0
      13'h1B85: dout  = 8'b00000000; // 7045 :   0 - 0x0
      13'h1B86: dout  = 8'b00000000; // 7046 :   0 - 0x0
      13'h1B87: dout  = 8'b00000000; // 7047 :   0 - 0x0
      13'h1B88: dout  = 8'b00000000; // 7048 :   0 - 0x0
      13'h1B89: dout  = 8'b00000000; // 7049 :   0 - 0x0
      13'h1B8A: dout  = 8'b00000000; // 7050 :   0 - 0x0
      13'h1B8B: dout  = 8'b00000000; // 7051 :   0 - 0x0
      13'h1B8C: dout  = 8'b00000000; // 7052 :   0 - 0x0
      13'h1B8D: dout  = 8'b00000000; // 7053 :   0 - 0x0
      13'h1B8E: dout  = 8'b00000000; // 7054 :   0 - 0x0
      13'h1B8F: dout  = 8'b00000000; // 7055 :   0 - 0x0
      13'h1B90: dout  = 8'b00000000; // 7056 :   0 - 0x0 -- Background 0xb9
      13'h1B91: dout  = 8'b00000000; // 7057 :   0 - 0x0
      13'h1B92: dout  = 8'b00000000; // 7058 :   0 - 0x0
      13'h1B93: dout  = 8'b00000000; // 7059 :   0 - 0x0
      13'h1B94: dout  = 8'b00000000; // 7060 :   0 - 0x0
      13'h1B95: dout  = 8'b00000000; // 7061 :   0 - 0x0
      13'h1B96: dout  = 8'b00000000; // 7062 :   0 - 0x0
      13'h1B97: dout  = 8'b00000000; // 7063 :   0 - 0x0
      13'h1B98: dout  = 8'b00000000; // 7064 :   0 - 0x0
      13'h1B99: dout  = 8'b00000000; // 7065 :   0 - 0x0
      13'h1B9A: dout  = 8'b00000000; // 7066 :   0 - 0x0
      13'h1B9B: dout  = 8'b00000000; // 7067 :   0 - 0x0
      13'h1B9C: dout  = 8'b00000000; // 7068 :   0 - 0x0
      13'h1B9D: dout  = 8'b00000000; // 7069 :   0 - 0x0
      13'h1B9E: dout  = 8'b00000000; // 7070 :   0 - 0x0
      13'h1B9F: dout  = 8'b00000000; // 7071 :   0 - 0x0
      13'h1BA0: dout  = 8'b00000000; // 7072 :   0 - 0x0 -- Background 0xba
      13'h1BA1: dout  = 8'b00000000; // 7073 :   0 - 0x0
      13'h1BA2: dout  = 8'b00000000; // 7074 :   0 - 0x0
      13'h1BA3: dout  = 8'b00000000; // 7075 :   0 - 0x0
      13'h1BA4: dout  = 8'b00000000; // 7076 :   0 - 0x0
      13'h1BA5: dout  = 8'b00000000; // 7077 :   0 - 0x0
      13'h1BA6: dout  = 8'b00000000; // 7078 :   0 - 0x0
      13'h1BA7: dout  = 8'b00000000; // 7079 :   0 - 0x0
      13'h1BA8: dout  = 8'b00000000; // 7080 :   0 - 0x0
      13'h1BA9: dout  = 8'b00000000; // 7081 :   0 - 0x0
      13'h1BAA: dout  = 8'b00000000; // 7082 :   0 - 0x0
      13'h1BAB: dout  = 8'b00000000; // 7083 :   0 - 0x0
      13'h1BAC: dout  = 8'b00000000; // 7084 :   0 - 0x0
      13'h1BAD: dout  = 8'b00000000; // 7085 :   0 - 0x0
      13'h1BAE: dout  = 8'b00000000; // 7086 :   0 - 0x0
      13'h1BAF: dout  = 8'b00000000; // 7087 :   0 - 0x0
      13'h1BB0: dout  = 8'b00000000; // 7088 :   0 - 0x0 -- Background 0xbb
      13'h1BB1: dout  = 8'b00000000; // 7089 :   0 - 0x0
      13'h1BB2: dout  = 8'b00000000; // 7090 :   0 - 0x0
      13'h1BB3: dout  = 8'b00000000; // 7091 :   0 - 0x0
      13'h1BB4: dout  = 8'b00000000; // 7092 :   0 - 0x0
      13'h1BB5: dout  = 8'b00000000; // 7093 :   0 - 0x0
      13'h1BB6: dout  = 8'b00000000; // 7094 :   0 - 0x0
      13'h1BB7: dout  = 8'b00000000; // 7095 :   0 - 0x0
      13'h1BB8: dout  = 8'b00000000; // 7096 :   0 - 0x0
      13'h1BB9: dout  = 8'b00000000; // 7097 :   0 - 0x0
      13'h1BBA: dout  = 8'b00000000; // 7098 :   0 - 0x0
      13'h1BBB: dout  = 8'b00000000; // 7099 :   0 - 0x0
      13'h1BBC: dout  = 8'b00000000; // 7100 :   0 - 0x0
      13'h1BBD: dout  = 8'b00000000; // 7101 :   0 - 0x0
      13'h1BBE: dout  = 8'b00000000; // 7102 :   0 - 0x0
      13'h1BBF: dout  = 8'b00000000; // 7103 :   0 - 0x0
      13'h1BC0: dout  = 8'b00000000; // 7104 :   0 - 0x0 -- Background 0xbc
      13'h1BC1: dout  = 8'b00000000; // 7105 :   0 - 0x0
      13'h1BC2: dout  = 8'b00000000; // 7106 :   0 - 0x0
      13'h1BC3: dout  = 8'b00000000; // 7107 :   0 - 0x0
      13'h1BC4: dout  = 8'b00000000; // 7108 :   0 - 0x0
      13'h1BC5: dout  = 8'b00000000; // 7109 :   0 - 0x0
      13'h1BC6: dout  = 8'b00000000; // 7110 :   0 - 0x0
      13'h1BC7: dout  = 8'b00000000; // 7111 :   0 - 0x0
      13'h1BC8: dout  = 8'b00000000; // 7112 :   0 - 0x0
      13'h1BC9: dout  = 8'b00000000; // 7113 :   0 - 0x0
      13'h1BCA: dout  = 8'b00000000; // 7114 :   0 - 0x0
      13'h1BCB: dout  = 8'b00000000; // 7115 :   0 - 0x0
      13'h1BCC: dout  = 8'b00000000; // 7116 :   0 - 0x0
      13'h1BCD: dout  = 8'b00000000; // 7117 :   0 - 0x0
      13'h1BCE: dout  = 8'b00000000; // 7118 :   0 - 0x0
      13'h1BCF: dout  = 8'b00000000; // 7119 :   0 - 0x0
      13'h1BD0: dout  = 8'b00000000; // 7120 :   0 - 0x0 -- Background 0xbd
      13'h1BD1: dout  = 8'b00000000; // 7121 :   0 - 0x0
      13'h1BD2: dout  = 8'b00000000; // 7122 :   0 - 0x0
      13'h1BD3: dout  = 8'b00000000; // 7123 :   0 - 0x0
      13'h1BD4: dout  = 8'b00000000; // 7124 :   0 - 0x0
      13'h1BD5: dout  = 8'b00000000; // 7125 :   0 - 0x0
      13'h1BD6: dout  = 8'b00000000; // 7126 :   0 - 0x0
      13'h1BD7: dout  = 8'b00000000; // 7127 :   0 - 0x0
      13'h1BD8: dout  = 8'b00000000; // 7128 :   0 - 0x0
      13'h1BD9: dout  = 8'b00000000; // 7129 :   0 - 0x0
      13'h1BDA: dout  = 8'b00000000; // 7130 :   0 - 0x0
      13'h1BDB: dout  = 8'b00000000; // 7131 :   0 - 0x0
      13'h1BDC: dout  = 8'b00000000; // 7132 :   0 - 0x0
      13'h1BDD: dout  = 8'b00000000; // 7133 :   0 - 0x0
      13'h1BDE: dout  = 8'b00000000; // 7134 :   0 - 0x0
      13'h1BDF: dout  = 8'b00000000; // 7135 :   0 - 0x0
      13'h1BE0: dout  = 8'b00000000; // 7136 :   0 - 0x0 -- Background 0xbe
      13'h1BE1: dout  = 8'b00000000; // 7137 :   0 - 0x0
      13'h1BE2: dout  = 8'b00000000; // 7138 :   0 - 0x0
      13'h1BE3: dout  = 8'b00000000; // 7139 :   0 - 0x0
      13'h1BE4: dout  = 8'b00000000; // 7140 :   0 - 0x0
      13'h1BE5: dout  = 8'b00000000; // 7141 :   0 - 0x0
      13'h1BE6: dout  = 8'b00000000; // 7142 :   0 - 0x0
      13'h1BE7: dout  = 8'b00000000; // 7143 :   0 - 0x0
      13'h1BE8: dout  = 8'b00000000; // 7144 :   0 - 0x0
      13'h1BE9: dout  = 8'b00000000; // 7145 :   0 - 0x0
      13'h1BEA: dout  = 8'b00000000; // 7146 :   0 - 0x0
      13'h1BEB: dout  = 8'b00000000; // 7147 :   0 - 0x0
      13'h1BEC: dout  = 8'b00000000; // 7148 :   0 - 0x0
      13'h1BED: dout  = 8'b00000000; // 7149 :   0 - 0x0
      13'h1BEE: dout  = 8'b00000000; // 7150 :   0 - 0x0
      13'h1BEF: dout  = 8'b00000000; // 7151 :   0 - 0x0
      13'h1BF0: dout  = 8'b00000000; // 7152 :   0 - 0x0 -- Background 0xbf
      13'h1BF1: dout  = 8'b00000000; // 7153 :   0 - 0x0
      13'h1BF2: dout  = 8'b00000000; // 7154 :   0 - 0x0
      13'h1BF3: dout  = 8'b00000000; // 7155 :   0 - 0x0
      13'h1BF4: dout  = 8'b00000000; // 7156 :   0 - 0x0
      13'h1BF5: dout  = 8'b00000000; // 7157 :   0 - 0x0
      13'h1BF6: dout  = 8'b00000000; // 7158 :   0 - 0x0
      13'h1BF7: dout  = 8'b00000000; // 7159 :   0 - 0x0
      13'h1BF8: dout  = 8'b00000000; // 7160 :   0 - 0x0
      13'h1BF9: dout  = 8'b00000000; // 7161 :   0 - 0x0
      13'h1BFA: dout  = 8'b00000000; // 7162 :   0 - 0x0
      13'h1BFB: dout  = 8'b00000000; // 7163 :   0 - 0x0
      13'h1BFC: dout  = 8'b00000000; // 7164 :   0 - 0x0
      13'h1BFD: dout  = 8'b00000000; // 7165 :   0 - 0x0
      13'h1BFE: dout  = 8'b00000000; // 7166 :   0 - 0x0
      13'h1BFF: dout  = 8'b00000000; // 7167 :   0 - 0x0
      13'h1C00: dout  = 8'b00000000; // 7168 :   0 - 0x0 -- Background 0xc0
      13'h1C01: dout  = 8'b00000000; // 7169 :   0 - 0x0
      13'h1C02: dout  = 8'b00000000; // 7170 :   0 - 0x0
      13'h1C03: dout  = 8'b00000000; // 7171 :   0 - 0x0
      13'h1C04: dout  = 8'b00000000; // 7172 :   0 - 0x0
      13'h1C05: dout  = 8'b00000000; // 7173 :   0 - 0x0
      13'h1C06: dout  = 8'b00000000; // 7174 :   0 - 0x0
      13'h1C07: dout  = 8'b00000000; // 7175 :   0 - 0x0
      13'h1C08: dout  = 8'b00000000; // 7176 :   0 - 0x0
      13'h1C09: dout  = 8'b00000000; // 7177 :   0 - 0x0
      13'h1C0A: dout  = 8'b00000000; // 7178 :   0 - 0x0
      13'h1C0B: dout  = 8'b00000000; // 7179 :   0 - 0x0
      13'h1C0C: dout  = 8'b00000000; // 7180 :   0 - 0x0
      13'h1C0D: dout  = 8'b00000000; // 7181 :   0 - 0x0
      13'h1C0E: dout  = 8'b00000000; // 7182 :   0 - 0x0
      13'h1C0F: dout  = 8'b00000000; // 7183 :   0 - 0x0
      13'h1C10: dout  = 8'b00000000; // 7184 :   0 - 0x0 -- Background 0xc1
      13'h1C11: dout  = 8'b00000000; // 7185 :   0 - 0x0
      13'h1C12: dout  = 8'b00000000; // 7186 :   0 - 0x0
      13'h1C13: dout  = 8'b00000000; // 7187 :   0 - 0x0
      13'h1C14: dout  = 8'b00000000; // 7188 :   0 - 0x0
      13'h1C15: dout  = 8'b00000000; // 7189 :   0 - 0x0
      13'h1C16: dout  = 8'b00000000; // 7190 :   0 - 0x0
      13'h1C17: dout  = 8'b00000000; // 7191 :   0 - 0x0
      13'h1C18: dout  = 8'b00000000; // 7192 :   0 - 0x0
      13'h1C19: dout  = 8'b00000000; // 7193 :   0 - 0x0
      13'h1C1A: dout  = 8'b00000000; // 7194 :   0 - 0x0
      13'h1C1B: dout  = 8'b00000000; // 7195 :   0 - 0x0
      13'h1C1C: dout  = 8'b00000000; // 7196 :   0 - 0x0
      13'h1C1D: dout  = 8'b00000000; // 7197 :   0 - 0x0
      13'h1C1E: dout  = 8'b00000000; // 7198 :   0 - 0x0
      13'h1C1F: dout  = 8'b00000000; // 7199 :   0 - 0x0
      13'h1C20: dout  = 8'b00000000; // 7200 :   0 - 0x0 -- Background 0xc2
      13'h1C21: dout  = 8'b00000000; // 7201 :   0 - 0x0
      13'h1C22: dout  = 8'b00000000; // 7202 :   0 - 0x0
      13'h1C23: dout  = 8'b00000000; // 7203 :   0 - 0x0
      13'h1C24: dout  = 8'b00000000; // 7204 :   0 - 0x0
      13'h1C25: dout  = 8'b00000000; // 7205 :   0 - 0x0
      13'h1C26: dout  = 8'b00000000; // 7206 :   0 - 0x0
      13'h1C27: dout  = 8'b00000000; // 7207 :   0 - 0x0
      13'h1C28: dout  = 8'b00000000; // 7208 :   0 - 0x0
      13'h1C29: dout  = 8'b00000000; // 7209 :   0 - 0x0
      13'h1C2A: dout  = 8'b00000000; // 7210 :   0 - 0x0
      13'h1C2B: dout  = 8'b00000000; // 7211 :   0 - 0x0
      13'h1C2C: dout  = 8'b00000000; // 7212 :   0 - 0x0
      13'h1C2D: dout  = 8'b00000000; // 7213 :   0 - 0x0
      13'h1C2E: dout  = 8'b00000000; // 7214 :   0 - 0x0
      13'h1C2F: dout  = 8'b00000000; // 7215 :   0 - 0x0
      13'h1C30: dout  = 8'b00000000; // 7216 :   0 - 0x0 -- Background 0xc3
      13'h1C31: dout  = 8'b00000000; // 7217 :   0 - 0x0
      13'h1C32: dout  = 8'b00000000; // 7218 :   0 - 0x0
      13'h1C33: dout  = 8'b00000000; // 7219 :   0 - 0x0
      13'h1C34: dout  = 8'b00000000; // 7220 :   0 - 0x0
      13'h1C35: dout  = 8'b00000000; // 7221 :   0 - 0x0
      13'h1C36: dout  = 8'b00000000; // 7222 :   0 - 0x0
      13'h1C37: dout  = 8'b00000000; // 7223 :   0 - 0x0
      13'h1C38: dout  = 8'b00000000; // 7224 :   0 - 0x0
      13'h1C39: dout  = 8'b00000000; // 7225 :   0 - 0x0
      13'h1C3A: dout  = 8'b00000000; // 7226 :   0 - 0x0
      13'h1C3B: dout  = 8'b00000000; // 7227 :   0 - 0x0
      13'h1C3C: dout  = 8'b00000000; // 7228 :   0 - 0x0
      13'h1C3D: dout  = 8'b00000000; // 7229 :   0 - 0x0
      13'h1C3E: dout  = 8'b00000000; // 7230 :   0 - 0x0
      13'h1C3F: dout  = 8'b00000000; // 7231 :   0 - 0x0
      13'h1C40: dout  = 8'b00000000; // 7232 :   0 - 0x0 -- Background 0xc4
      13'h1C41: dout  = 8'b00000000; // 7233 :   0 - 0x0
      13'h1C42: dout  = 8'b00000000; // 7234 :   0 - 0x0
      13'h1C43: dout  = 8'b00000000; // 7235 :   0 - 0x0
      13'h1C44: dout  = 8'b00000000; // 7236 :   0 - 0x0
      13'h1C45: dout  = 8'b00000000; // 7237 :   0 - 0x0
      13'h1C46: dout  = 8'b00000000; // 7238 :   0 - 0x0
      13'h1C47: dout  = 8'b00000000; // 7239 :   0 - 0x0
      13'h1C48: dout  = 8'b00000000; // 7240 :   0 - 0x0
      13'h1C49: dout  = 8'b00000000; // 7241 :   0 - 0x0
      13'h1C4A: dout  = 8'b00000000; // 7242 :   0 - 0x0
      13'h1C4B: dout  = 8'b00000000; // 7243 :   0 - 0x0
      13'h1C4C: dout  = 8'b00000000; // 7244 :   0 - 0x0
      13'h1C4D: dout  = 8'b00000000; // 7245 :   0 - 0x0
      13'h1C4E: dout  = 8'b00000000; // 7246 :   0 - 0x0
      13'h1C4F: dout  = 8'b00000000; // 7247 :   0 - 0x0
      13'h1C50: dout  = 8'b00000000; // 7248 :   0 - 0x0 -- Background 0xc5
      13'h1C51: dout  = 8'b00000000; // 7249 :   0 - 0x0
      13'h1C52: dout  = 8'b00000000; // 7250 :   0 - 0x0
      13'h1C53: dout  = 8'b00000000; // 7251 :   0 - 0x0
      13'h1C54: dout  = 8'b00000000; // 7252 :   0 - 0x0
      13'h1C55: dout  = 8'b00000000; // 7253 :   0 - 0x0
      13'h1C56: dout  = 8'b00000000; // 7254 :   0 - 0x0
      13'h1C57: dout  = 8'b00000000; // 7255 :   0 - 0x0
      13'h1C58: dout  = 8'b00000000; // 7256 :   0 - 0x0
      13'h1C59: dout  = 8'b00000000; // 7257 :   0 - 0x0
      13'h1C5A: dout  = 8'b00000000; // 7258 :   0 - 0x0
      13'h1C5B: dout  = 8'b00000000; // 7259 :   0 - 0x0
      13'h1C5C: dout  = 8'b00000000; // 7260 :   0 - 0x0
      13'h1C5D: dout  = 8'b00000000; // 7261 :   0 - 0x0
      13'h1C5E: dout  = 8'b00000000; // 7262 :   0 - 0x0
      13'h1C5F: dout  = 8'b00000000; // 7263 :   0 - 0x0
      13'h1C60: dout  = 8'b00000000; // 7264 :   0 - 0x0 -- Background 0xc6
      13'h1C61: dout  = 8'b00000000; // 7265 :   0 - 0x0
      13'h1C62: dout  = 8'b00000000; // 7266 :   0 - 0x0
      13'h1C63: dout  = 8'b00000000; // 7267 :   0 - 0x0
      13'h1C64: dout  = 8'b00000000; // 7268 :   0 - 0x0
      13'h1C65: dout  = 8'b00000000; // 7269 :   0 - 0x0
      13'h1C66: dout  = 8'b00000000; // 7270 :   0 - 0x0
      13'h1C67: dout  = 8'b00000000; // 7271 :   0 - 0x0
      13'h1C68: dout  = 8'b00000000; // 7272 :   0 - 0x0
      13'h1C69: dout  = 8'b00000000; // 7273 :   0 - 0x0
      13'h1C6A: dout  = 8'b00000000; // 7274 :   0 - 0x0
      13'h1C6B: dout  = 8'b00000000; // 7275 :   0 - 0x0
      13'h1C6C: dout  = 8'b00000000; // 7276 :   0 - 0x0
      13'h1C6D: dout  = 8'b00000000; // 7277 :   0 - 0x0
      13'h1C6E: dout  = 8'b00000000; // 7278 :   0 - 0x0
      13'h1C6F: dout  = 8'b00000000; // 7279 :   0 - 0x0
      13'h1C70: dout  = 8'b00000000; // 7280 :   0 - 0x0 -- Background 0xc7
      13'h1C71: dout  = 8'b00000000; // 7281 :   0 - 0x0
      13'h1C72: dout  = 8'b00000000; // 7282 :   0 - 0x0
      13'h1C73: dout  = 8'b00000000; // 7283 :   0 - 0x0
      13'h1C74: dout  = 8'b00000000; // 7284 :   0 - 0x0
      13'h1C75: dout  = 8'b00000000; // 7285 :   0 - 0x0
      13'h1C76: dout  = 8'b00000000; // 7286 :   0 - 0x0
      13'h1C77: dout  = 8'b00000000; // 7287 :   0 - 0x0
      13'h1C78: dout  = 8'b00000000; // 7288 :   0 - 0x0
      13'h1C79: dout  = 8'b00000000; // 7289 :   0 - 0x0
      13'h1C7A: dout  = 8'b00000000; // 7290 :   0 - 0x0
      13'h1C7B: dout  = 8'b00000000; // 7291 :   0 - 0x0
      13'h1C7C: dout  = 8'b00000000; // 7292 :   0 - 0x0
      13'h1C7D: dout  = 8'b00000000; // 7293 :   0 - 0x0
      13'h1C7E: dout  = 8'b00000000; // 7294 :   0 - 0x0
      13'h1C7F: dout  = 8'b00000000; // 7295 :   0 - 0x0
      13'h1C80: dout  = 8'b00000000; // 7296 :   0 - 0x0 -- Background 0xc8
      13'h1C81: dout  = 8'b00000000; // 7297 :   0 - 0x0
      13'h1C82: dout  = 8'b00000000; // 7298 :   0 - 0x0
      13'h1C83: dout  = 8'b00000000; // 7299 :   0 - 0x0
      13'h1C84: dout  = 8'b00000000; // 7300 :   0 - 0x0
      13'h1C85: dout  = 8'b00000000; // 7301 :   0 - 0x0
      13'h1C86: dout  = 8'b00000000; // 7302 :   0 - 0x0
      13'h1C87: dout  = 8'b00000000; // 7303 :   0 - 0x0
      13'h1C88: dout  = 8'b00000000; // 7304 :   0 - 0x0
      13'h1C89: dout  = 8'b00000000; // 7305 :   0 - 0x0
      13'h1C8A: dout  = 8'b00000000; // 7306 :   0 - 0x0
      13'h1C8B: dout  = 8'b00000000; // 7307 :   0 - 0x0
      13'h1C8C: dout  = 8'b00000000; // 7308 :   0 - 0x0
      13'h1C8D: dout  = 8'b00000000; // 7309 :   0 - 0x0
      13'h1C8E: dout  = 8'b00000000; // 7310 :   0 - 0x0
      13'h1C8F: dout  = 8'b00000000; // 7311 :   0 - 0x0
      13'h1C90: dout  = 8'b00000000; // 7312 :   0 - 0x0 -- Background 0xc9
      13'h1C91: dout  = 8'b00000000; // 7313 :   0 - 0x0
      13'h1C92: dout  = 8'b00000000; // 7314 :   0 - 0x0
      13'h1C93: dout  = 8'b00000000; // 7315 :   0 - 0x0
      13'h1C94: dout  = 8'b00000000; // 7316 :   0 - 0x0
      13'h1C95: dout  = 8'b00000000; // 7317 :   0 - 0x0
      13'h1C96: dout  = 8'b00000000; // 7318 :   0 - 0x0
      13'h1C97: dout  = 8'b00000000; // 7319 :   0 - 0x0
      13'h1C98: dout  = 8'b00000000; // 7320 :   0 - 0x0
      13'h1C99: dout  = 8'b00000000; // 7321 :   0 - 0x0
      13'h1C9A: dout  = 8'b00000000; // 7322 :   0 - 0x0
      13'h1C9B: dout  = 8'b00000000; // 7323 :   0 - 0x0
      13'h1C9C: dout  = 8'b00000000; // 7324 :   0 - 0x0
      13'h1C9D: dout  = 8'b00000000; // 7325 :   0 - 0x0
      13'h1C9E: dout  = 8'b00000000; // 7326 :   0 - 0x0
      13'h1C9F: dout  = 8'b00000000; // 7327 :   0 - 0x0
      13'h1CA0: dout  = 8'b00000000; // 7328 :   0 - 0x0 -- Background 0xca
      13'h1CA1: dout  = 8'b00000000; // 7329 :   0 - 0x0
      13'h1CA2: dout  = 8'b00000000; // 7330 :   0 - 0x0
      13'h1CA3: dout  = 8'b00000000; // 7331 :   0 - 0x0
      13'h1CA4: dout  = 8'b00000000; // 7332 :   0 - 0x0
      13'h1CA5: dout  = 8'b00000000; // 7333 :   0 - 0x0
      13'h1CA6: dout  = 8'b00000000; // 7334 :   0 - 0x0
      13'h1CA7: dout  = 8'b00000000; // 7335 :   0 - 0x0
      13'h1CA8: dout  = 8'b00000000; // 7336 :   0 - 0x0
      13'h1CA9: dout  = 8'b00000000; // 7337 :   0 - 0x0
      13'h1CAA: dout  = 8'b00000000; // 7338 :   0 - 0x0
      13'h1CAB: dout  = 8'b00000000; // 7339 :   0 - 0x0
      13'h1CAC: dout  = 8'b00000000; // 7340 :   0 - 0x0
      13'h1CAD: dout  = 8'b00000000; // 7341 :   0 - 0x0
      13'h1CAE: dout  = 8'b00000000; // 7342 :   0 - 0x0
      13'h1CAF: dout  = 8'b00000000; // 7343 :   0 - 0x0
      13'h1CB0: dout  = 8'b00000000; // 7344 :   0 - 0x0 -- Background 0xcb
      13'h1CB1: dout  = 8'b00000000; // 7345 :   0 - 0x0
      13'h1CB2: dout  = 8'b00000000; // 7346 :   0 - 0x0
      13'h1CB3: dout  = 8'b00000000; // 7347 :   0 - 0x0
      13'h1CB4: dout  = 8'b00000000; // 7348 :   0 - 0x0
      13'h1CB5: dout  = 8'b00000000; // 7349 :   0 - 0x0
      13'h1CB6: dout  = 8'b00000000; // 7350 :   0 - 0x0
      13'h1CB7: dout  = 8'b00000000; // 7351 :   0 - 0x0
      13'h1CB8: dout  = 8'b00000000; // 7352 :   0 - 0x0
      13'h1CB9: dout  = 8'b00000000; // 7353 :   0 - 0x0
      13'h1CBA: dout  = 8'b00000000; // 7354 :   0 - 0x0
      13'h1CBB: dout  = 8'b00000000; // 7355 :   0 - 0x0
      13'h1CBC: dout  = 8'b00000000; // 7356 :   0 - 0x0
      13'h1CBD: dout  = 8'b00000000; // 7357 :   0 - 0x0
      13'h1CBE: dout  = 8'b00000000; // 7358 :   0 - 0x0
      13'h1CBF: dout  = 8'b00000000; // 7359 :   0 - 0x0
      13'h1CC0: dout  = 8'b00000000; // 7360 :   0 - 0x0 -- Background 0xcc
      13'h1CC1: dout  = 8'b00000000; // 7361 :   0 - 0x0
      13'h1CC2: dout  = 8'b00000000; // 7362 :   0 - 0x0
      13'h1CC3: dout  = 8'b00000000; // 7363 :   0 - 0x0
      13'h1CC4: dout  = 8'b00000000; // 7364 :   0 - 0x0
      13'h1CC5: dout  = 8'b00000000; // 7365 :   0 - 0x0
      13'h1CC6: dout  = 8'b00000000; // 7366 :   0 - 0x0
      13'h1CC7: dout  = 8'b00000000; // 7367 :   0 - 0x0
      13'h1CC8: dout  = 8'b00000000; // 7368 :   0 - 0x0
      13'h1CC9: dout  = 8'b00000000; // 7369 :   0 - 0x0
      13'h1CCA: dout  = 8'b00000000; // 7370 :   0 - 0x0
      13'h1CCB: dout  = 8'b00000000; // 7371 :   0 - 0x0
      13'h1CCC: dout  = 8'b00000000; // 7372 :   0 - 0x0
      13'h1CCD: dout  = 8'b00000000; // 7373 :   0 - 0x0
      13'h1CCE: dout  = 8'b00000000; // 7374 :   0 - 0x0
      13'h1CCF: dout  = 8'b00000000; // 7375 :   0 - 0x0
      13'h1CD0: dout  = 8'b00111111; // 7376 :  63 - 0x3f -- Background 0xcd
      13'h1CD1: dout  = 8'b01111111; // 7377 : 127 - 0x7f
      13'h1CD2: dout  = 8'b11111111; // 7378 : 255 - 0xff
      13'h1CD3: dout  = 8'b11110000; // 7379 : 240 - 0xf0
      13'h1CD4: dout  = 8'b11100000; // 7380 : 224 - 0xe0
      13'h1CD5: dout  = 8'b11100011; // 7381 : 227 - 0xe3
      13'h1CD6: dout  = 8'b11100111; // 7382 : 231 - 0xe7
      13'h1CD7: dout  = 8'b11100111; // 7383 : 231 - 0xe7
      13'h1CD8: dout  = 8'b11000000; // 7384 : 192 - 0xc0
      13'h1CD9: dout  = 8'b10000000; // 7385 : 128 - 0x80
      13'h1CDA: dout  = 8'b00000000; // 7386 :   0 - 0x0
      13'h1CDB: dout  = 8'b00001111; // 7387 :  15 - 0xf
      13'h1CDC: dout  = 8'b00011111; // 7388 :  31 - 0x1f
      13'h1CDD: dout  = 8'b00011100; // 7389 :  28 - 0x1c
      13'h1CDE: dout  = 8'b00011000; // 7390 :  24 - 0x18
      13'h1CDF: dout  = 8'b00011000; // 7391 :  24 - 0x18
      13'h1CE0: dout  = 8'b11111100; // 7392 : 252 - 0xfc -- Background 0xce
      13'h1CE1: dout  = 8'b11111110; // 7393 : 254 - 0xfe
      13'h1CE2: dout  = 8'b11111111; // 7394 : 255 - 0xff
      13'h1CE3: dout  = 8'b00001111; // 7395 :  15 - 0xf
      13'h1CE4: dout  = 8'b00000111; // 7396 :   7 - 0x7
      13'h1CE5: dout  = 8'b11000111; // 7397 : 199 - 0xc7
      13'h1CE6: dout  = 8'b11100111; // 7398 : 231 - 0xe7
      13'h1CE7: dout  = 8'b11100111; // 7399 : 231 - 0xe7
      13'h1CE8: dout  = 8'b00000011; // 7400 :   3 - 0x3
      13'h1CE9: dout  = 8'b00000001; // 7401 :   1 - 0x1
      13'h1CEA: dout  = 8'b00000000; // 7402 :   0 - 0x0
      13'h1CEB: dout  = 8'b11110000; // 7403 : 240 - 0xf0
      13'h1CEC: dout  = 8'b11111000; // 7404 : 248 - 0xf8
      13'h1CED: dout  = 8'b00111000; // 7405 :  56 - 0x38
      13'h1CEE: dout  = 8'b00011000; // 7406 :  24 - 0x18
      13'h1CEF: dout  = 8'b00011000; // 7407 :  24 - 0x18
      13'h1CF0: dout  = 8'b00000000; // 7408 :   0 - 0x0 -- Background 0xcf
      13'h1CF1: dout  = 8'b00000000; // 7409 :   0 - 0x0
      13'h1CF2: dout  = 8'b00000000; // 7410 :   0 - 0x0
      13'h1CF3: dout  = 8'b00000000; // 7411 :   0 - 0x0
      13'h1CF4: dout  = 8'b00000000; // 7412 :   0 - 0x0
      13'h1CF5: dout  = 8'b00000000; // 7413 :   0 - 0x0
      13'h1CF6: dout  = 8'b00000000; // 7414 :   0 - 0x0
      13'h1CF7: dout  = 8'b00000000; // 7415 :   0 - 0x0
      13'h1CF8: dout  = 8'b00000000; // 7416 :   0 - 0x0
      13'h1CF9: dout  = 8'b00000000; // 7417 :   0 - 0x0
      13'h1CFA: dout  = 8'b00000000; // 7418 :   0 - 0x0
      13'h1CFB: dout  = 8'b00000000; // 7419 :   0 - 0x0
      13'h1CFC: dout  = 8'b00000000; // 7420 :   0 - 0x0
      13'h1CFD: dout  = 8'b00000000; // 7421 :   0 - 0x0
      13'h1CFE: dout  = 8'b00000000; // 7422 :   0 - 0x0
      13'h1CFF: dout  = 8'b00000000; // 7423 :   0 - 0x0
      13'h1D00: dout  = 8'b00000000; // 7424 :   0 - 0x0 -- Background 0xd0
      13'h1D01: dout  = 8'b00000000; // 7425 :   0 - 0x0
      13'h1D02: dout  = 8'b00000000; // 7426 :   0 - 0x0
      13'h1D03: dout  = 8'b00000000; // 7427 :   0 - 0x0
      13'h1D04: dout  = 8'b00000000; // 7428 :   0 - 0x0
      13'h1D05: dout  = 8'b00000000; // 7429 :   0 - 0x0
      13'h1D06: dout  = 8'b00000000; // 7430 :   0 - 0x0
      13'h1D07: dout  = 8'b00000000; // 7431 :   0 - 0x0
      13'h1D08: dout  = 8'b00000000; // 7432 :   0 - 0x0
      13'h1D09: dout  = 8'b00000000; // 7433 :   0 - 0x0
      13'h1D0A: dout  = 8'b00000000; // 7434 :   0 - 0x0
      13'h1D0B: dout  = 8'b00000000; // 7435 :   0 - 0x0
      13'h1D0C: dout  = 8'b00000000; // 7436 :   0 - 0x0
      13'h1D0D: dout  = 8'b00000000; // 7437 :   0 - 0x0
      13'h1D0E: dout  = 8'b00000000; // 7438 :   0 - 0x0
      13'h1D0F: dout  = 8'b00000000; // 7439 :   0 - 0x0
      13'h1D10: dout  = 8'b00000000; // 7440 :   0 - 0x0 -- Background 0xd1
      13'h1D11: dout  = 8'b00000000; // 7441 :   0 - 0x0
      13'h1D12: dout  = 8'b00000000; // 7442 :   0 - 0x0
      13'h1D13: dout  = 8'b00000000; // 7443 :   0 - 0x0
      13'h1D14: dout  = 8'b00000000; // 7444 :   0 - 0x0
      13'h1D15: dout  = 8'b00000000; // 7445 :   0 - 0x0
      13'h1D16: dout  = 8'b00000000; // 7446 :   0 - 0x0
      13'h1D17: dout  = 8'b00000000; // 7447 :   0 - 0x0
      13'h1D18: dout  = 8'b00000000; // 7448 :   0 - 0x0
      13'h1D19: dout  = 8'b00000000; // 7449 :   0 - 0x0
      13'h1D1A: dout  = 8'b00000000; // 7450 :   0 - 0x0
      13'h1D1B: dout  = 8'b00000000; // 7451 :   0 - 0x0
      13'h1D1C: dout  = 8'b00000000; // 7452 :   0 - 0x0
      13'h1D1D: dout  = 8'b00000000; // 7453 :   0 - 0x0
      13'h1D1E: dout  = 8'b00000000; // 7454 :   0 - 0x0
      13'h1D1F: dout  = 8'b00000000; // 7455 :   0 - 0x0
      13'h1D20: dout  = 8'b00000000; // 7456 :   0 - 0x0 -- Background 0xd2
      13'h1D21: dout  = 8'b00000000; // 7457 :   0 - 0x0
      13'h1D22: dout  = 8'b00000000; // 7458 :   0 - 0x0
      13'h1D23: dout  = 8'b00000000; // 7459 :   0 - 0x0
      13'h1D24: dout  = 8'b00000000; // 7460 :   0 - 0x0
      13'h1D25: dout  = 8'b00000000; // 7461 :   0 - 0x0
      13'h1D26: dout  = 8'b00000000; // 7462 :   0 - 0x0
      13'h1D27: dout  = 8'b00000000; // 7463 :   0 - 0x0
      13'h1D28: dout  = 8'b00000000; // 7464 :   0 - 0x0
      13'h1D29: dout  = 8'b00000000; // 7465 :   0 - 0x0
      13'h1D2A: dout  = 8'b00000000; // 7466 :   0 - 0x0
      13'h1D2B: dout  = 8'b00000000; // 7467 :   0 - 0x0
      13'h1D2C: dout  = 8'b00000000; // 7468 :   0 - 0x0
      13'h1D2D: dout  = 8'b00000000; // 7469 :   0 - 0x0
      13'h1D2E: dout  = 8'b00000000; // 7470 :   0 - 0x0
      13'h1D2F: dout  = 8'b00000000; // 7471 :   0 - 0x0
      13'h1D30: dout  = 8'b00000000; // 7472 :   0 - 0x0 -- Background 0xd3
      13'h1D31: dout  = 8'b00000000; // 7473 :   0 - 0x0
      13'h1D32: dout  = 8'b00000000; // 7474 :   0 - 0x0
      13'h1D33: dout  = 8'b00000000; // 7475 :   0 - 0x0
      13'h1D34: dout  = 8'b00000000; // 7476 :   0 - 0x0
      13'h1D35: dout  = 8'b00000000; // 7477 :   0 - 0x0
      13'h1D36: dout  = 8'b00000000; // 7478 :   0 - 0x0
      13'h1D37: dout  = 8'b00000000; // 7479 :   0 - 0x0
      13'h1D38: dout  = 8'b00000000; // 7480 :   0 - 0x0
      13'h1D39: dout  = 8'b00000000; // 7481 :   0 - 0x0
      13'h1D3A: dout  = 8'b00000000; // 7482 :   0 - 0x0
      13'h1D3B: dout  = 8'b00000000; // 7483 :   0 - 0x0
      13'h1D3C: dout  = 8'b00000000; // 7484 :   0 - 0x0
      13'h1D3D: dout  = 8'b00000000; // 7485 :   0 - 0x0
      13'h1D3E: dout  = 8'b00000000; // 7486 :   0 - 0x0
      13'h1D3F: dout  = 8'b00000000; // 7487 :   0 - 0x0
      13'h1D40: dout  = 8'b00000000; // 7488 :   0 - 0x0 -- Background 0xd4
      13'h1D41: dout  = 8'b00000000; // 7489 :   0 - 0x0
      13'h1D42: dout  = 8'b00000000; // 7490 :   0 - 0x0
      13'h1D43: dout  = 8'b00000000; // 7491 :   0 - 0x0
      13'h1D44: dout  = 8'b00000000; // 7492 :   0 - 0x0
      13'h1D45: dout  = 8'b00000000; // 7493 :   0 - 0x0
      13'h1D46: dout  = 8'b00000000; // 7494 :   0 - 0x0
      13'h1D47: dout  = 8'b00000000; // 7495 :   0 - 0x0
      13'h1D48: dout  = 8'b00000000; // 7496 :   0 - 0x0
      13'h1D49: dout  = 8'b00000000; // 7497 :   0 - 0x0
      13'h1D4A: dout  = 8'b00000000; // 7498 :   0 - 0x0
      13'h1D4B: dout  = 8'b00000000; // 7499 :   0 - 0x0
      13'h1D4C: dout  = 8'b00000000; // 7500 :   0 - 0x0
      13'h1D4D: dout  = 8'b00000000; // 7501 :   0 - 0x0
      13'h1D4E: dout  = 8'b00000000; // 7502 :   0 - 0x0
      13'h1D4F: dout  = 8'b00000000; // 7503 :   0 - 0x0
      13'h1D50: dout  = 8'b00000000; // 7504 :   0 - 0x0 -- Background 0xd5
      13'h1D51: dout  = 8'b00000000; // 7505 :   0 - 0x0
      13'h1D52: dout  = 8'b00000000; // 7506 :   0 - 0x0
      13'h1D53: dout  = 8'b00000000; // 7507 :   0 - 0x0
      13'h1D54: dout  = 8'b00000000; // 7508 :   0 - 0x0
      13'h1D55: dout  = 8'b00000000; // 7509 :   0 - 0x0
      13'h1D56: dout  = 8'b00000000; // 7510 :   0 - 0x0
      13'h1D57: dout  = 8'b00000000; // 7511 :   0 - 0x0
      13'h1D58: dout  = 8'b00000000; // 7512 :   0 - 0x0
      13'h1D59: dout  = 8'b00000000; // 7513 :   0 - 0x0
      13'h1D5A: dout  = 8'b00000000; // 7514 :   0 - 0x0
      13'h1D5B: dout  = 8'b00000000; // 7515 :   0 - 0x0
      13'h1D5C: dout  = 8'b00000000; // 7516 :   0 - 0x0
      13'h1D5D: dout  = 8'b00000000; // 7517 :   0 - 0x0
      13'h1D5E: dout  = 8'b00000000; // 7518 :   0 - 0x0
      13'h1D5F: dout  = 8'b00000000; // 7519 :   0 - 0x0
      13'h1D60: dout  = 8'b00000000; // 7520 :   0 - 0x0 -- Background 0xd6
      13'h1D61: dout  = 8'b00000000; // 7521 :   0 - 0x0
      13'h1D62: dout  = 8'b00000000; // 7522 :   0 - 0x0
      13'h1D63: dout  = 8'b00000000; // 7523 :   0 - 0x0
      13'h1D64: dout  = 8'b00000000; // 7524 :   0 - 0x0
      13'h1D65: dout  = 8'b00000000; // 7525 :   0 - 0x0
      13'h1D66: dout  = 8'b00000000; // 7526 :   0 - 0x0
      13'h1D67: dout  = 8'b00000000; // 7527 :   0 - 0x0
      13'h1D68: dout  = 8'b00000000; // 7528 :   0 - 0x0
      13'h1D69: dout  = 8'b00000000; // 7529 :   0 - 0x0
      13'h1D6A: dout  = 8'b00000000; // 7530 :   0 - 0x0
      13'h1D6B: dout  = 8'b00000000; // 7531 :   0 - 0x0
      13'h1D6C: dout  = 8'b00000000; // 7532 :   0 - 0x0
      13'h1D6D: dout  = 8'b00000000; // 7533 :   0 - 0x0
      13'h1D6E: dout  = 8'b00000000; // 7534 :   0 - 0x0
      13'h1D6F: dout  = 8'b00000000; // 7535 :   0 - 0x0
      13'h1D70: dout  = 8'b00000000; // 7536 :   0 - 0x0 -- Background 0xd7
      13'h1D71: dout  = 8'b00000000; // 7537 :   0 - 0x0
      13'h1D72: dout  = 8'b00000000; // 7538 :   0 - 0x0
      13'h1D73: dout  = 8'b00000000; // 7539 :   0 - 0x0
      13'h1D74: dout  = 8'b00000000; // 7540 :   0 - 0x0
      13'h1D75: dout  = 8'b00000000; // 7541 :   0 - 0x0
      13'h1D76: dout  = 8'b00000000; // 7542 :   0 - 0x0
      13'h1D77: dout  = 8'b00000000; // 7543 :   0 - 0x0
      13'h1D78: dout  = 8'b00000000; // 7544 :   0 - 0x0
      13'h1D79: dout  = 8'b00000000; // 7545 :   0 - 0x0
      13'h1D7A: dout  = 8'b00000000; // 7546 :   0 - 0x0
      13'h1D7B: dout  = 8'b00000000; // 7547 :   0 - 0x0
      13'h1D7C: dout  = 8'b00000000; // 7548 :   0 - 0x0
      13'h1D7D: dout  = 8'b00000000; // 7549 :   0 - 0x0
      13'h1D7E: dout  = 8'b00000000; // 7550 :   0 - 0x0
      13'h1D7F: dout  = 8'b00000000; // 7551 :   0 - 0x0
      13'h1D80: dout  = 8'b00000000; // 7552 :   0 - 0x0 -- Background 0xd8
      13'h1D81: dout  = 8'b00000000; // 7553 :   0 - 0x0
      13'h1D82: dout  = 8'b00000000; // 7554 :   0 - 0x0
      13'h1D83: dout  = 8'b00000000; // 7555 :   0 - 0x0
      13'h1D84: dout  = 8'b00000000; // 7556 :   0 - 0x0
      13'h1D85: dout  = 8'b00000000; // 7557 :   0 - 0x0
      13'h1D86: dout  = 8'b00000000; // 7558 :   0 - 0x0
      13'h1D87: dout  = 8'b00000000; // 7559 :   0 - 0x0
      13'h1D88: dout  = 8'b00000000; // 7560 :   0 - 0x0
      13'h1D89: dout  = 8'b00000000; // 7561 :   0 - 0x0
      13'h1D8A: dout  = 8'b00000000; // 7562 :   0 - 0x0
      13'h1D8B: dout  = 8'b00000000; // 7563 :   0 - 0x0
      13'h1D8C: dout  = 8'b00000000; // 7564 :   0 - 0x0
      13'h1D8D: dout  = 8'b00000000; // 7565 :   0 - 0x0
      13'h1D8E: dout  = 8'b00000000; // 7566 :   0 - 0x0
      13'h1D8F: dout  = 8'b00000000; // 7567 :   0 - 0x0
      13'h1D90: dout  = 8'b00000000; // 7568 :   0 - 0x0 -- Background 0xd9
      13'h1D91: dout  = 8'b00000000; // 7569 :   0 - 0x0
      13'h1D92: dout  = 8'b00000000; // 7570 :   0 - 0x0
      13'h1D93: dout  = 8'b00000000; // 7571 :   0 - 0x0
      13'h1D94: dout  = 8'b00000000; // 7572 :   0 - 0x0
      13'h1D95: dout  = 8'b00000000; // 7573 :   0 - 0x0
      13'h1D96: dout  = 8'b00000000; // 7574 :   0 - 0x0
      13'h1D97: dout  = 8'b00000000; // 7575 :   0 - 0x0
      13'h1D98: dout  = 8'b00000000; // 7576 :   0 - 0x0
      13'h1D99: dout  = 8'b00000000; // 7577 :   0 - 0x0
      13'h1D9A: dout  = 8'b00000000; // 7578 :   0 - 0x0
      13'h1D9B: dout  = 8'b00000000; // 7579 :   0 - 0x0
      13'h1D9C: dout  = 8'b00000000; // 7580 :   0 - 0x0
      13'h1D9D: dout  = 8'b00000000; // 7581 :   0 - 0x0
      13'h1D9E: dout  = 8'b00000000; // 7582 :   0 - 0x0
      13'h1D9F: dout  = 8'b00000000; // 7583 :   0 - 0x0
      13'h1DA0: dout  = 8'b00000000; // 7584 :   0 - 0x0 -- Background 0xda
      13'h1DA1: dout  = 8'b00000000; // 7585 :   0 - 0x0
      13'h1DA2: dout  = 8'b00000000; // 7586 :   0 - 0x0
      13'h1DA3: dout  = 8'b00000000; // 7587 :   0 - 0x0
      13'h1DA4: dout  = 8'b00000000; // 7588 :   0 - 0x0
      13'h1DA5: dout  = 8'b00000000; // 7589 :   0 - 0x0
      13'h1DA6: dout  = 8'b00000000; // 7590 :   0 - 0x0
      13'h1DA7: dout  = 8'b00000000; // 7591 :   0 - 0x0
      13'h1DA8: dout  = 8'b00000000; // 7592 :   0 - 0x0
      13'h1DA9: dout  = 8'b00000000; // 7593 :   0 - 0x0
      13'h1DAA: dout  = 8'b00000000; // 7594 :   0 - 0x0
      13'h1DAB: dout  = 8'b00000000; // 7595 :   0 - 0x0
      13'h1DAC: dout  = 8'b00000000; // 7596 :   0 - 0x0
      13'h1DAD: dout  = 8'b00000000; // 7597 :   0 - 0x0
      13'h1DAE: dout  = 8'b00000000; // 7598 :   0 - 0x0
      13'h1DAF: dout  = 8'b00000000; // 7599 :   0 - 0x0
      13'h1DB0: dout  = 8'b00000000; // 7600 :   0 - 0x0 -- Background 0xdb
      13'h1DB1: dout  = 8'b00000000; // 7601 :   0 - 0x0
      13'h1DB2: dout  = 8'b00000000; // 7602 :   0 - 0x0
      13'h1DB3: dout  = 8'b00000000; // 7603 :   0 - 0x0
      13'h1DB4: dout  = 8'b00000000; // 7604 :   0 - 0x0
      13'h1DB5: dout  = 8'b00000000; // 7605 :   0 - 0x0
      13'h1DB6: dout  = 8'b00000000; // 7606 :   0 - 0x0
      13'h1DB7: dout  = 8'b00000000; // 7607 :   0 - 0x0
      13'h1DB8: dout  = 8'b00000000; // 7608 :   0 - 0x0
      13'h1DB9: dout  = 8'b00000000; // 7609 :   0 - 0x0
      13'h1DBA: dout  = 8'b00000000; // 7610 :   0 - 0x0
      13'h1DBB: dout  = 8'b00000000; // 7611 :   0 - 0x0
      13'h1DBC: dout  = 8'b00000000; // 7612 :   0 - 0x0
      13'h1DBD: dout  = 8'b00000000; // 7613 :   0 - 0x0
      13'h1DBE: dout  = 8'b00000000; // 7614 :   0 - 0x0
      13'h1DBF: dout  = 8'b00000000; // 7615 :   0 - 0x0
      13'h1DC0: dout  = 8'b00000000; // 7616 :   0 - 0x0 -- Background 0xdc
      13'h1DC1: dout  = 8'b00000000; // 7617 :   0 - 0x0
      13'h1DC2: dout  = 8'b00000000; // 7618 :   0 - 0x0
      13'h1DC3: dout  = 8'b00000000; // 7619 :   0 - 0x0
      13'h1DC4: dout  = 8'b00000000; // 7620 :   0 - 0x0
      13'h1DC5: dout  = 8'b00000000; // 7621 :   0 - 0x0
      13'h1DC6: dout  = 8'b00000000; // 7622 :   0 - 0x0
      13'h1DC7: dout  = 8'b00000000; // 7623 :   0 - 0x0
      13'h1DC8: dout  = 8'b00000000; // 7624 :   0 - 0x0
      13'h1DC9: dout  = 8'b00000000; // 7625 :   0 - 0x0
      13'h1DCA: dout  = 8'b00000000; // 7626 :   0 - 0x0
      13'h1DCB: dout  = 8'b00000000; // 7627 :   0 - 0x0
      13'h1DCC: dout  = 8'b00000000; // 7628 :   0 - 0x0
      13'h1DCD: dout  = 8'b00000000; // 7629 :   0 - 0x0
      13'h1DCE: dout  = 8'b00000000; // 7630 :   0 - 0x0
      13'h1DCF: dout  = 8'b00000000; // 7631 :   0 - 0x0
      13'h1DD0: dout  = 8'b11100111; // 7632 : 231 - 0xe7 -- Background 0xdd
      13'h1DD1: dout  = 8'b11100111; // 7633 : 231 - 0xe7
      13'h1DD2: dout  = 8'b11100011; // 7634 : 227 - 0xe3
      13'h1DD3: dout  = 8'b11100000; // 7635 : 224 - 0xe0
      13'h1DD4: dout  = 8'b11110000; // 7636 : 240 - 0xf0
      13'h1DD5: dout  = 8'b11111111; // 7637 : 255 - 0xff
      13'h1DD6: dout  = 8'b01111111; // 7638 : 127 - 0x7f
      13'h1DD7: dout  = 8'b00111111; // 7639 :  63 - 0x3f
      13'h1DD8: dout  = 8'b00011000; // 7640 :  24 - 0x18
      13'h1DD9: dout  = 8'b00011000; // 7641 :  24 - 0x18
      13'h1DDA: dout  = 8'b00011100; // 7642 :  28 - 0x1c
      13'h1DDB: dout  = 8'b00011111; // 7643 :  31 - 0x1f
      13'h1DDC: dout  = 8'b00001111; // 7644 :  15 - 0xf
      13'h1DDD: dout  = 8'b00000000; // 7645 :   0 - 0x0
      13'h1DDE: dout  = 8'b10000000; // 7646 : 128 - 0x80
      13'h1DDF: dout  = 8'b11000000; // 7647 : 192 - 0xc0
      13'h1DE0: dout  = 8'b11100111; // 7648 : 231 - 0xe7 -- Background 0xde
      13'h1DE1: dout  = 8'b11100111; // 7649 : 231 - 0xe7
      13'h1DE2: dout  = 8'b11000111; // 7650 : 199 - 0xc7
      13'h1DE3: dout  = 8'b00000111; // 7651 :   7 - 0x7
      13'h1DE4: dout  = 8'b00001111; // 7652 :  15 - 0xf
      13'h1DE5: dout  = 8'b11111111; // 7653 : 255 - 0xff
      13'h1DE6: dout  = 8'b11111110; // 7654 : 254 - 0xfe
      13'h1DE7: dout  = 8'b11111100; // 7655 : 252 - 0xfc
      13'h1DE8: dout  = 8'b00011000; // 7656 :  24 - 0x18
      13'h1DE9: dout  = 8'b00011000; // 7657 :  24 - 0x18
      13'h1DEA: dout  = 8'b00111000; // 7658 :  56 - 0x38
      13'h1DEB: dout  = 8'b11111000; // 7659 : 248 - 0xf8
      13'h1DEC: dout  = 8'b11110000; // 7660 : 240 - 0xf0
      13'h1DED: dout  = 8'b00000000; // 7661 :   0 - 0x0
      13'h1DEE: dout  = 8'b00000001; // 7662 :   1 - 0x1
      13'h1DEF: dout  = 8'b00000011; // 7663 :   3 - 0x3
      13'h1DF0: dout  = 8'b00000000; // 7664 :   0 - 0x0 -- Background 0xdf
      13'h1DF1: dout  = 8'b00000000; // 7665 :   0 - 0x0
      13'h1DF2: dout  = 8'b00000000; // 7666 :   0 - 0x0
      13'h1DF3: dout  = 8'b00000000; // 7667 :   0 - 0x0
      13'h1DF4: dout  = 8'b00000000; // 7668 :   0 - 0x0
      13'h1DF5: dout  = 8'b00000000; // 7669 :   0 - 0x0
      13'h1DF6: dout  = 8'b00000000; // 7670 :   0 - 0x0
      13'h1DF7: dout  = 8'b00000000; // 7671 :   0 - 0x0
      13'h1DF8: dout  = 8'b00000000; // 7672 :   0 - 0x0
      13'h1DF9: dout  = 8'b00000000; // 7673 :   0 - 0x0
      13'h1DFA: dout  = 8'b00000000; // 7674 :   0 - 0x0
      13'h1DFB: dout  = 8'b00000000; // 7675 :   0 - 0x0
      13'h1DFC: dout  = 8'b00000000; // 7676 :   0 - 0x0
      13'h1DFD: dout  = 8'b00000000; // 7677 :   0 - 0x0
      13'h1DFE: dout  = 8'b00000000; // 7678 :   0 - 0x0
      13'h1DFF: dout  = 8'b00000000; // 7679 :   0 - 0x0
      13'h1E00: dout  = 8'b00000000; // 7680 :   0 - 0x0 -- Background 0xe0
      13'h1E01: dout  = 8'b00000000; // 7681 :   0 - 0x0
      13'h1E02: dout  = 8'b00000000; // 7682 :   0 - 0x0
      13'h1E03: dout  = 8'b00000000; // 7683 :   0 - 0x0
      13'h1E04: dout  = 8'b00000000; // 7684 :   0 - 0x0
      13'h1E05: dout  = 8'b00000000; // 7685 :   0 - 0x0
      13'h1E06: dout  = 8'b00000000; // 7686 :   0 - 0x0
      13'h1E07: dout  = 8'b00000000; // 7687 :   0 - 0x0
      13'h1E08: dout  = 8'b00000000; // 7688 :   0 - 0x0
      13'h1E09: dout  = 8'b00000000; // 7689 :   0 - 0x0
      13'h1E0A: dout  = 8'b00000000; // 7690 :   0 - 0x0
      13'h1E0B: dout  = 8'b00000000; // 7691 :   0 - 0x0
      13'h1E0C: dout  = 8'b00000000; // 7692 :   0 - 0x0
      13'h1E0D: dout  = 8'b00000000; // 7693 :   0 - 0x0
      13'h1E0E: dout  = 8'b00000000; // 7694 :   0 - 0x0
      13'h1E0F: dout  = 8'b00000000; // 7695 :   0 - 0x0
      13'h1E10: dout  = 8'b00000000; // 7696 :   0 - 0x0 -- Background 0xe1
      13'h1E11: dout  = 8'b00000000; // 7697 :   0 - 0x0
      13'h1E12: dout  = 8'b00000000; // 7698 :   0 - 0x0
      13'h1E13: dout  = 8'b00000000; // 7699 :   0 - 0x0
      13'h1E14: dout  = 8'b00000000; // 7700 :   0 - 0x0
      13'h1E15: dout  = 8'b00000000; // 7701 :   0 - 0x0
      13'h1E16: dout  = 8'b00000000; // 7702 :   0 - 0x0
      13'h1E17: dout  = 8'b00000000; // 7703 :   0 - 0x0
      13'h1E18: dout  = 8'b00000000; // 7704 :   0 - 0x0
      13'h1E19: dout  = 8'b00000000; // 7705 :   0 - 0x0
      13'h1E1A: dout  = 8'b00000000; // 7706 :   0 - 0x0
      13'h1E1B: dout  = 8'b00000000; // 7707 :   0 - 0x0
      13'h1E1C: dout  = 8'b00000000; // 7708 :   0 - 0x0
      13'h1E1D: dout  = 8'b00000000; // 7709 :   0 - 0x0
      13'h1E1E: dout  = 8'b00000000; // 7710 :   0 - 0x0
      13'h1E1F: dout  = 8'b00000000; // 7711 :   0 - 0x0
      13'h1E20: dout  = 8'b00000000; // 7712 :   0 - 0x0 -- Background 0xe2
      13'h1E21: dout  = 8'b00000000; // 7713 :   0 - 0x0
      13'h1E22: dout  = 8'b00000000; // 7714 :   0 - 0x0
      13'h1E23: dout  = 8'b00000000; // 7715 :   0 - 0x0
      13'h1E24: dout  = 8'b00000000; // 7716 :   0 - 0x0
      13'h1E25: dout  = 8'b00000000; // 7717 :   0 - 0x0
      13'h1E26: dout  = 8'b00000000; // 7718 :   0 - 0x0
      13'h1E27: dout  = 8'b00000000; // 7719 :   0 - 0x0
      13'h1E28: dout  = 8'b00000000; // 7720 :   0 - 0x0
      13'h1E29: dout  = 8'b00000000; // 7721 :   0 - 0x0
      13'h1E2A: dout  = 8'b00000000; // 7722 :   0 - 0x0
      13'h1E2B: dout  = 8'b00000000; // 7723 :   0 - 0x0
      13'h1E2C: dout  = 8'b00000000; // 7724 :   0 - 0x0
      13'h1E2D: dout  = 8'b00000000; // 7725 :   0 - 0x0
      13'h1E2E: dout  = 8'b00000000; // 7726 :   0 - 0x0
      13'h1E2F: dout  = 8'b00000000; // 7727 :   0 - 0x0
      13'h1E30: dout  = 8'b00000000; // 7728 :   0 - 0x0 -- Background 0xe3
      13'h1E31: dout  = 8'b00000000; // 7729 :   0 - 0x0
      13'h1E32: dout  = 8'b00000000; // 7730 :   0 - 0x0
      13'h1E33: dout  = 8'b00000000; // 7731 :   0 - 0x0
      13'h1E34: dout  = 8'b00000000; // 7732 :   0 - 0x0
      13'h1E35: dout  = 8'b00000000; // 7733 :   0 - 0x0
      13'h1E36: dout  = 8'b00000000; // 7734 :   0 - 0x0
      13'h1E37: dout  = 8'b00000000; // 7735 :   0 - 0x0
      13'h1E38: dout  = 8'b00000000; // 7736 :   0 - 0x0
      13'h1E39: dout  = 8'b00000000; // 7737 :   0 - 0x0
      13'h1E3A: dout  = 8'b00000000; // 7738 :   0 - 0x0
      13'h1E3B: dout  = 8'b00000000; // 7739 :   0 - 0x0
      13'h1E3C: dout  = 8'b00000000; // 7740 :   0 - 0x0
      13'h1E3D: dout  = 8'b00000000; // 7741 :   0 - 0x0
      13'h1E3E: dout  = 8'b00000000; // 7742 :   0 - 0x0
      13'h1E3F: dout  = 8'b00000000; // 7743 :   0 - 0x0
      13'h1E40: dout  = 8'b00000000; // 7744 :   0 - 0x0 -- Background 0xe4
      13'h1E41: dout  = 8'b00000000; // 7745 :   0 - 0x0
      13'h1E42: dout  = 8'b00000000; // 7746 :   0 - 0x0
      13'h1E43: dout  = 8'b00000000; // 7747 :   0 - 0x0
      13'h1E44: dout  = 8'b00000000; // 7748 :   0 - 0x0
      13'h1E45: dout  = 8'b00000000; // 7749 :   0 - 0x0
      13'h1E46: dout  = 8'b00000000; // 7750 :   0 - 0x0
      13'h1E47: dout  = 8'b00000000; // 7751 :   0 - 0x0
      13'h1E48: dout  = 8'b00000000; // 7752 :   0 - 0x0
      13'h1E49: dout  = 8'b00000000; // 7753 :   0 - 0x0
      13'h1E4A: dout  = 8'b00000000; // 7754 :   0 - 0x0
      13'h1E4B: dout  = 8'b00000000; // 7755 :   0 - 0x0
      13'h1E4C: dout  = 8'b00000000; // 7756 :   0 - 0x0
      13'h1E4D: dout  = 8'b00000000; // 7757 :   0 - 0x0
      13'h1E4E: dout  = 8'b00000000; // 7758 :   0 - 0x0
      13'h1E4F: dout  = 8'b00000000; // 7759 :   0 - 0x0
      13'h1E50: dout  = 8'b01111111; // 7760 : 127 - 0x7f -- Background 0xe5
      13'h1E51: dout  = 8'b11111111; // 7761 : 255 - 0xff
      13'h1E52: dout  = 8'b11111111; // 7762 : 255 - 0xff
      13'h1E53: dout  = 8'b11100000; // 7763 : 224 - 0xe0
      13'h1E54: dout  = 8'b11100000; // 7764 : 224 - 0xe0
      13'h1E55: dout  = 8'b11100000; // 7765 : 224 - 0xe0
      13'h1E56: dout  = 8'b11100000; // 7766 : 224 - 0xe0
      13'h1E57: dout  = 8'b11100001; // 7767 : 225 - 0xe1
      13'h1E58: dout  = 8'b00000000; // 7768 :   0 - 0x0
      13'h1E59: dout  = 8'b00000000; // 7769 :   0 - 0x0
      13'h1E5A: dout  = 8'b00000000; // 7770 :   0 - 0x0
      13'h1E5B: dout  = 8'b00000000; // 7771 :   0 - 0x0
      13'h1E5C: dout  = 8'b00000000; // 7772 :   0 - 0x0
      13'h1E5D: dout  = 8'b00000000; // 7773 :   0 - 0x0
      13'h1E5E: dout  = 8'b00000000; // 7774 :   0 - 0x0
      13'h1E5F: dout  = 8'b00000000; // 7775 :   0 - 0x0
      13'h1E60: dout  = 8'b11111110; // 7776 : 254 - 0xfe -- Background 0xe6
      13'h1E61: dout  = 8'b11111111; // 7777 : 255 - 0xff
      13'h1E62: dout  = 8'b11111111; // 7778 : 255 - 0xff
      13'h1E63: dout  = 8'b00000111; // 7779 :   7 - 0x7
      13'h1E64: dout  = 8'b00000111; // 7780 :   7 - 0x7
      13'h1E65: dout  = 8'b00000111; // 7781 :   7 - 0x7
      13'h1E66: dout  = 8'b00000111; // 7782 :   7 - 0x7
      13'h1E67: dout  = 8'b10000111; // 7783 : 135 - 0x87
      13'h1E68: dout  = 8'b00000000; // 7784 :   0 - 0x0
      13'h1E69: dout  = 8'b00000000; // 7785 :   0 - 0x0
      13'h1E6A: dout  = 8'b00000000; // 7786 :   0 - 0x0
      13'h1E6B: dout  = 8'b00000000; // 7787 :   0 - 0x0
      13'h1E6C: dout  = 8'b00000000; // 7788 :   0 - 0x0
      13'h1E6D: dout  = 8'b00000000; // 7789 :   0 - 0x0
      13'h1E6E: dout  = 8'b00000000; // 7790 :   0 - 0x0
      13'h1E6F: dout  = 8'b00000000; // 7791 :   0 - 0x0
      13'h1E70: dout  = 8'b00011111; // 7792 :  31 - 0x1f -- Background 0xe7
      13'h1E71: dout  = 8'b00100000; // 7793 :  32 - 0x20
      13'h1E72: dout  = 8'b01000000; // 7794 :  64 - 0x40
      13'h1E73: dout  = 8'b10000000; // 7795 : 128 - 0x80
      13'h1E74: dout  = 8'b10000000; // 7796 : 128 - 0x80
      13'h1E75: dout  = 8'b10000011; // 7797 : 131 - 0x83
      13'h1E76: dout  = 8'b10000111; // 7798 : 135 - 0x87
      13'h1E77: dout  = 8'b10000111; // 7799 : 135 - 0x87
      13'h1E78: dout  = 8'b11100000; // 7800 : 224 - 0xe0
      13'h1E79: dout  = 8'b11000000; // 7801 : 192 - 0xc0
      13'h1E7A: dout  = 8'b10000000; // 7802 : 128 - 0x80
      13'h1E7B: dout  = 8'b00000000; // 7803 :   0 - 0x0
      13'h1E7C: dout  = 8'b00000000; // 7804 :   0 - 0x0
      13'h1E7D: dout  = 8'b00000000; // 7805 :   0 - 0x0
      13'h1E7E: dout  = 8'b00000000; // 7806 :   0 - 0x0
      13'h1E7F: dout  = 8'b00000000; // 7807 :   0 - 0x0
      13'h1E80: dout  = 8'b11111000; // 7808 : 248 - 0xf8 -- Background 0xe8
      13'h1E81: dout  = 8'b00000100; // 7809 :   4 - 0x4
      13'h1E82: dout  = 8'b00000010; // 7810 :   2 - 0x2
      13'h1E83: dout  = 8'b00000001; // 7811 :   1 - 0x1
      13'h1E84: dout  = 8'b00000001; // 7812 :   1 - 0x1
      13'h1E85: dout  = 8'b11000001; // 7813 : 193 - 0xc1
      13'h1E86: dout  = 8'b11100001; // 7814 : 225 - 0xe1
      13'h1E87: dout  = 8'b11100001; // 7815 : 225 - 0xe1
      13'h1E88: dout  = 8'b00000111; // 7816 :   7 - 0x7
      13'h1E89: dout  = 8'b00000011; // 7817 :   3 - 0x3
      13'h1E8A: dout  = 8'b00000001; // 7818 :   1 - 0x1
      13'h1E8B: dout  = 8'b00000000; // 7819 :   0 - 0x0
      13'h1E8C: dout  = 8'b00000000; // 7820 :   0 - 0x0
      13'h1E8D: dout  = 8'b00000000; // 7821 :   0 - 0x0
      13'h1E8E: dout  = 8'b00000000; // 7822 :   0 - 0x0
      13'h1E8F: dout  = 8'b00000000; // 7823 :   0 - 0x0
      13'h1E90: dout  = 8'b00000000; // 7824 :   0 - 0x0 -- Background 0xe9
      13'h1E91: dout  = 8'b00000000; // 7825 :   0 - 0x0
      13'h1E92: dout  = 8'b00001000; // 7826 :   8 - 0x8
      13'h1E93: dout  = 8'b00010100; // 7827 :  20 - 0x14
      13'h1E94: dout  = 8'b00000000; // 7828 :   0 - 0x0
      13'h1E95: dout  = 8'b00000000; // 7829 :   0 - 0x0
      13'h1E96: dout  = 8'b01000000; // 7830 :  64 - 0x40
      13'h1E97: dout  = 8'b10100000; // 7831 : 160 - 0xa0
      13'h1E98: dout  = 8'b11111111; // 7832 : 255 - 0xff
      13'h1E99: dout  = 8'b11111111; // 7833 : 255 - 0xff
      13'h1E9A: dout  = 8'b11111111; // 7834 : 255 - 0xff
      13'h1E9B: dout  = 8'b11111111; // 7835 : 255 - 0xff
      13'h1E9C: dout  = 8'b11111111; // 7836 : 255 - 0xff
      13'h1E9D: dout  = 8'b11111111; // 7837 : 255 - 0xff
      13'h1E9E: dout  = 8'b11111111; // 7838 : 255 - 0xff
      13'h1E9F: dout  = 8'b11111111; // 7839 : 255 - 0xff
      13'h1EA0: dout  = 8'b01000000; // 7840 :  64 - 0x40 -- Background 0xea
      13'h1EA1: dout  = 8'b10100010; // 7841 : 162 - 0xa2
      13'h1EA2: dout  = 8'b00000101; // 7842 :   5 - 0x5
      13'h1EA3: dout  = 8'b00000000; // 7843 :   0 - 0x0
      13'h1EA4: dout  = 8'b00000000; // 7844 :   0 - 0x0
      13'h1EA5: dout  = 8'b00010000; // 7845 :  16 - 0x10
      13'h1EA6: dout  = 8'b00101000; // 7846 :  40 - 0x28
      13'h1EA7: dout  = 8'b00000000; // 7847 :   0 - 0x0
      13'h1EA8: dout  = 8'b11111111; // 7848 : 255 - 0xff
      13'h1EA9: dout  = 8'b11111111; // 7849 : 255 - 0xff
      13'h1EAA: dout  = 8'b11111111; // 7850 : 255 - 0xff
      13'h1EAB: dout  = 8'b11111111; // 7851 : 255 - 0xff
      13'h1EAC: dout  = 8'b11111111; // 7852 : 255 - 0xff
      13'h1EAD: dout  = 8'b11111111; // 7853 : 255 - 0xff
      13'h1EAE: dout  = 8'b11111111; // 7854 : 255 - 0xff
      13'h1EAF: dout  = 8'b11111111; // 7855 : 255 - 0xff
      13'h1EB0: dout  = 8'b11111111; // 7856 : 255 - 0xff -- Background 0xeb
      13'h1EB1: dout  = 8'b11111111; // 7857 : 255 - 0xff
      13'h1EB2: dout  = 8'b11111111; // 7858 : 255 - 0xff
      13'h1EB3: dout  = 8'b00000000; // 7859 :   0 - 0x0
      13'h1EB4: dout  = 8'b00000000; // 7860 :   0 - 0x0
      13'h1EB5: dout  = 8'b00000000; // 7861 :   0 - 0x0
      13'h1EB6: dout  = 8'b00000000; // 7862 :   0 - 0x0
      13'h1EB7: dout  = 8'b11111111; // 7863 : 255 - 0xff
      13'h1EB8: dout  = 8'b00000000; // 7864 :   0 - 0x0
      13'h1EB9: dout  = 8'b00000000; // 7865 :   0 - 0x0
      13'h1EBA: dout  = 8'b00000000; // 7866 :   0 - 0x0
      13'h1EBB: dout  = 8'b00000000; // 7867 :   0 - 0x0
      13'h1EBC: dout  = 8'b00000000; // 7868 :   0 - 0x0
      13'h1EBD: dout  = 8'b00000000; // 7869 :   0 - 0x0
      13'h1EBE: dout  = 8'b00000000; // 7870 :   0 - 0x0
      13'h1EBF: dout  = 8'b00000000; // 7871 :   0 - 0x0
      13'h1EC0: dout  = 8'b11100001; // 7872 : 225 - 0xe1 -- Background 0xec
      13'h1EC1: dout  = 8'b11100001; // 7873 : 225 - 0xe1
      13'h1EC2: dout  = 8'b11100001; // 7874 : 225 - 0xe1
      13'h1EC3: dout  = 8'b11100001; // 7875 : 225 - 0xe1
      13'h1EC4: dout  = 8'b11100001; // 7876 : 225 - 0xe1
      13'h1EC5: dout  = 8'b11100001; // 7877 : 225 - 0xe1
      13'h1EC6: dout  = 8'b11100001; // 7878 : 225 - 0xe1
      13'h1EC7: dout  = 8'b11100001; // 7879 : 225 - 0xe1
      13'h1EC8: dout  = 8'b00000000; // 7880 :   0 - 0x0
      13'h1EC9: dout  = 8'b00000000; // 7881 :   0 - 0x0
      13'h1ECA: dout  = 8'b00000000; // 7882 :   0 - 0x0
      13'h1ECB: dout  = 8'b00000000; // 7883 :   0 - 0x0
      13'h1ECC: dout  = 8'b00000000; // 7884 :   0 - 0x0
      13'h1ECD: dout  = 8'b00000000; // 7885 :   0 - 0x0
      13'h1ECE: dout  = 8'b00000000; // 7886 :   0 - 0x0
      13'h1ECF: dout  = 8'b00000000; // 7887 :   0 - 0x0
      13'h1ED0: dout  = 8'b11111111; // 7888 : 255 - 0xff -- Background 0xed
      13'h1ED1: dout  = 8'b11111111; // 7889 : 255 - 0xff
      13'h1ED2: dout  = 8'b11111111; // 7890 : 255 - 0xff
      13'h1ED3: dout  = 8'b00000000; // 7891 :   0 - 0x0
      13'h1ED4: dout  = 8'b00000000; // 7892 :   0 - 0x0
      13'h1ED5: dout  = 8'b11111111; // 7893 : 255 - 0xff
      13'h1ED6: dout  = 8'b11111111; // 7894 : 255 - 0xff
      13'h1ED7: dout  = 8'b11111111; // 7895 : 255 - 0xff
      13'h1ED8: dout  = 8'b00000000; // 7896 :   0 - 0x0
      13'h1ED9: dout  = 8'b00000000; // 7897 :   0 - 0x0
      13'h1EDA: dout  = 8'b00000000; // 7898 :   0 - 0x0
      13'h1EDB: dout  = 8'b11111111; // 7899 : 255 - 0xff
      13'h1EDC: dout  = 8'b11111111; // 7900 : 255 - 0xff
      13'h1EDD: dout  = 8'b00000000; // 7901 :   0 - 0x0
      13'h1EDE: dout  = 8'b00000000; // 7902 :   0 - 0x0
      13'h1EDF: dout  = 8'b00000000; // 7903 :   0 - 0x0
      13'h1EE0: dout  = 8'b11100111; // 7904 : 231 - 0xe7 -- Background 0xee
      13'h1EE1: dout  = 8'b11100111; // 7905 : 231 - 0xe7
      13'h1EE2: dout  = 8'b11100111; // 7906 : 231 - 0xe7
      13'h1EE3: dout  = 8'b11100111; // 7907 : 231 - 0xe7
      13'h1EE4: dout  = 8'b11100111; // 7908 : 231 - 0xe7
      13'h1EE5: dout  = 8'b11100111; // 7909 : 231 - 0xe7
      13'h1EE6: dout  = 8'b11100111; // 7910 : 231 - 0xe7
      13'h1EE7: dout  = 8'b11100111; // 7911 : 231 - 0xe7
      13'h1EE8: dout  = 8'b00011000; // 7912 :  24 - 0x18
      13'h1EE9: dout  = 8'b00011000; // 7913 :  24 - 0x18
      13'h1EEA: dout  = 8'b00011000; // 7914 :  24 - 0x18
      13'h1EEB: dout  = 8'b00011000; // 7915 :  24 - 0x18
      13'h1EEC: dout  = 8'b00011000; // 7916 :  24 - 0x18
      13'h1EED: dout  = 8'b00011000; // 7917 :  24 - 0x18
      13'h1EEE: dout  = 8'b00011000; // 7918 :  24 - 0x18
      13'h1EEF: dout  = 8'b00011000; // 7919 :  24 - 0x18
      13'h1EF0: dout  = 8'b11111111; // 7920 : 255 - 0xff -- Background 0xef
      13'h1EF1: dout  = 8'b11111111; // 7921 : 255 - 0xff
      13'h1EF2: dout  = 8'b11111111; // 7922 : 255 - 0xff
      13'h1EF3: dout  = 8'b11111111; // 7923 : 255 - 0xff
      13'h1EF4: dout  = 8'b11111111; // 7924 : 255 - 0xff
      13'h1EF5: dout  = 8'b11111111; // 7925 : 255 - 0xff
      13'h1EF6: dout  = 8'b11111111; // 7926 : 255 - 0xff
      13'h1EF7: dout  = 8'b11111111; // 7927 : 255 - 0xff
      13'h1EF8: dout  = 8'b00110011; // 7928 :  51 - 0x33
      13'h1EF9: dout  = 8'b00110011; // 7929 :  51 - 0x33
      13'h1EFA: dout  = 8'b11001100; // 7930 : 204 - 0xcc
      13'h1EFB: dout  = 8'b11001100; // 7931 : 204 - 0xcc
      13'h1EFC: dout  = 8'b00110011; // 7932 :  51 - 0x33
      13'h1EFD: dout  = 8'b00110011; // 7933 :  51 - 0x33
      13'h1EFE: dout  = 8'b11001100; // 7934 : 204 - 0xcc
      13'h1EFF: dout  = 8'b11001100; // 7935 : 204 - 0xcc
      13'h1F00: dout  = 8'b00000000; // 7936 :   0 - 0x0 -- Background 0xf0
      13'h1F01: dout  = 8'b00000000; // 7937 :   0 - 0x0
      13'h1F02: dout  = 8'b00000000; // 7938 :   0 - 0x0
      13'h1F03: dout  = 8'b00000000; // 7939 :   0 - 0x0
      13'h1F04: dout  = 8'b00000000; // 7940 :   0 - 0x0
      13'h1F05: dout  = 8'b00000000; // 7941 :   0 - 0x0
      13'h1F06: dout  = 8'b00000000; // 7942 :   0 - 0x0
      13'h1F07: dout  = 8'b00000000; // 7943 :   0 - 0x0
      13'h1F08: dout  = 8'b00000000; // 7944 :   0 - 0x0
      13'h1F09: dout  = 8'b00000000; // 7945 :   0 - 0x0
      13'h1F0A: dout  = 8'b00000000; // 7946 :   0 - 0x0
      13'h1F0B: dout  = 8'b00000000; // 7947 :   0 - 0x0
      13'h1F0C: dout  = 8'b00000000; // 7948 :   0 - 0x0
      13'h1F0D: dout  = 8'b00000000; // 7949 :   0 - 0x0
      13'h1F0E: dout  = 8'b00000000; // 7950 :   0 - 0x0
      13'h1F0F: dout  = 8'b00000000; // 7951 :   0 - 0x0
      13'h1F10: dout  = 8'b00000000; // 7952 :   0 - 0x0 -- Background 0xf1
      13'h1F11: dout  = 8'b00000000; // 7953 :   0 - 0x0
      13'h1F12: dout  = 8'b00000000; // 7954 :   0 - 0x0
      13'h1F13: dout  = 8'b00000000; // 7955 :   0 - 0x0
      13'h1F14: dout  = 8'b00000000; // 7956 :   0 - 0x0
      13'h1F15: dout  = 8'b00000000; // 7957 :   0 - 0x0
      13'h1F16: dout  = 8'b00000000; // 7958 :   0 - 0x0
      13'h1F17: dout  = 8'b00000000; // 7959 :   0 - 0x0
      13'h1F18: dout  = 8'b00000000; // 7960 :   0 - 0x0
      13'h1F19: dout  = 8'b00000000; // 7961 :   0 - 0x0
      13'h1F1A: dout  = 8'b00000000; // 7962 :   0 - 0x0
      13'h1F1B: dout  = 8'b00000000; // 7963 :   0 - 0x0
      13'h1F1C: dout  = 8'b00000000; // 7964 :   0 - 0x0
      13'h1F1D: dout  = 8'b00000000; // 7965 :   0 - 0x0
      13'h1F1E: dout  = 8'b00000000; // 7966 :   0 - 0x0
      13'h1F1F: dout  = 8'b00000000; // 7967 :   0 - 0x0
      13'h1F20: dout  = 8'b00000000; // 7968 :   0 - 0x0 -- Background 0xf2
      13'h1F21: dout  = 8'b00000000; // 7969 :   0 - 0x0
      13'h1F22: dout  = 8'b00000000; // 7970 :   0 - 0x0
      13'h1F23: dout  = 8'b00000000; // 7971 :   0 - 0x0
      13'h1F24: dout  = 8'b00000000; // 7972 :   0 - 0x0
      13'h1F25: dout  = 8'b00000000; // 7973 :   0 - 0x0
      13'h1F26: dout  = 8'b00000000; // 7974 :   0 - 0x0
      13'h1F27: dout  = 8'b00000000; // 7975 :   0 - 0x0
      13'h1F28: dout  = 8'b00000000; // 7976 :   0 - 0x0
      13'h1F29: dout  = 8'b00000000; // 7977 :   0 - 0x0
      13'h1F2A: dout  = 8'b00000000; // 7978 :   0 - 0x0
      13'h1F2B: dout  = 8'b00000000; // 7979 :   0 - 0x0
      13'h1F2C: dout  = 8'b00000000; // 7980 :   0 - 0x0
      13'h1F2D: dout  = 8'b00000000; // 7981 :   0 - 0x0
      13'h1F2E: dout  = 8'b00000000; // 7982 :   0 - 0x0
      13'h1F2F: dout  = 8'b00000000; // 7983 :   0 - 0x0
      13'h1F30: dout  = 8'b00000000; // 7984 :   0 - 0x0 -- Background 0xf3
      13'h1F31: dout  = 8'b00000000; // 7985 :   0 - 0x0
      13'h1F32: dout  = 8'b00000000; // 7986 :   0 - 0x0
      13'h1F33: dout  = 8'b00000000; // 7987 :   0 - 0x0
      13'h1F34: dout  = 8'b00000000; // 7988 :   0 - 0x0
      13'h1F35: dout  = 8'b00000000; // 7989 :   0 - 0x0
      13'h1F36: dout  = 8'b00000000; // 7990 :   0 - 0x0
      13'h1F37: dout  = 8'b00000000; // 7991 :   0 - 0x0
      13'h1F38: dout  = 8'b00000000; // 7992 :   0 - 0x0
      13'h1F39: dout  = 8'b00000000; // 7993 :   0 - 0x0
      13'h1F3A: dout  = 8'b00000000; // 7994 :   0 - 0x0
      13'h1F3B: dout  = 8'b00000000; // 7995 :   0 - 0x0
      13'h1F3C: dout  = 8'b00000000; // 7996 :   0 - 0x0
      13'h1F3D: dout  = 8'b00000000; // 7997 :   0 - 0x0
      13'h1F3E: dout  = 8'b00000000; // 7998 :   0 - 0x0
      13'h1F3F: dout  = 8'b00000000; // 7999 :   0 - 0x0
      13'h1F40: dout  = 8'b11100111; // 8000 : 231 - 0xe7 -- Background 0xf4
      13'h1F41: dout  = 8'b10011001; // 8001 : 153 - 0x99
      13'h1F42: dout  = 8'b10000001; // 8002 : 129 - 0x81
      13'h1F43: dout  = 8'b11000011; // 8003 : 195 - 0xc3
      13'h1F44: dout  = 8'b11111111; // 8004 : 255 - 0xff
      13'h1F45: dout  = 8'b10111101; // 8005 : 189 - 0xbd
      13'h1F46: dout  = 8'b10000001; // 8006 : 129 - 0x81
      13'h1F47: dout  = 8'b11000011; // 8007 : 195 - 0xc3
      13'h1F48: dout  = 8'b00100100; // 8008 :  36 - 0x24
      13'h1F49: dout  = 8'b00011000; // 8009 :  24 - 0x18
      13'h1F4A: dout  = 8'b00000000; // 8010 :   0 - 0x0
      13'h1F4B: dout  = 8'b01000010; // 8011 :  66 - 0x42
      13'h1F4C: dout  = 8'b01111110; // 8012 : 126 - 0x7e
      13'h1F4D: dout  = 8'b00111100; // 8013 :  60 - 0x3c
      13'h1F4E: dout  = 8'b00000000; // 8014 :   0 - 0x0
      13'h1F4F: dout  = 8'b00000000; // 8015 :   0 - 0x0
      13'h1F50: dout  = 8'b11100001; // 8016 : 225 - 0xe1 -- Background 0xf5
      13'h1F51: dout  = 8'b11100000; // 8017 : 224 - 0xe0
      13'h1F52: dout  = 8'b11100000; // 8018 : 224 - 0xe0
      13'h1F53: dout  = 8'b11100000; // 8019 : 224 - 0xe0
      13'h1F54: dout  = 8'b11100000; // 8020 : 224 - 0xe0
      13'h1F55: dout  = 8'b11111111; // 8021 : 255 - 0xff
      13'h1F56: dout  = 8'b11111111; // 8022 : 255 - 0xff
      13'h1F57: dout  = 8'b01111111; // 8023 : 127 - 0x7f
      13'h1F58: dout  = 8'b00000000; // 8024 :   0 - 0x0
      13'h1F59: dout  = 8'b00000000; // 8025 :   0 - 0x0
      13'h1F5A: dout  = 8'b00000000; // 8026 :   0 - 0x0
      13'h1F5B: dout  = 8'b00000000; // 8027 :   0 - 0x0
      13'h1F5C: dout  = 8'b00000000; // 8028 :   0 - 0x0
      13'h1F5D: dout  = 8'b00000000; // 8029 :   0 - 0x0
      13'h1F5E: dout  = 8'b00000000; // 8030 :   0 - 0x0
      13'h1F5F: dout  = 8'b00000000; // 8031 :   0 - 0x0
      13'h1F60: dout  = 8'b10000111; // 8032 : 135 - 0x87 -- Background 0xf6
      13'h1F61: dout  = 8'b00000111; // 8033 :   7 - 0x7
      13'h1F62: dout  = 8'b00000111; // 8034 :   7 - 0x7
      13'h1F63: dout  = 8'b00000111; // 8035 :   7 - 0x7
      13'h1F64: dout  = 8'b00000111; // 8036 :   7 - 0x7
      13'h1F65: dout  = 8'b11111111; // 8037 : 255 - 0xff
      13'h1F66: dout  = 8'b11111111; // 8038 : 255 - 0xff
      13'h1F67: dout  = 8'b11111110; // 8039 : 254 - 0xfe
      13'h1F68: dout  = 8'b00000000; // 8040 :   0 - 0x0
      13'h1F69: dout  = 8'b00000000; // 8041 :   0 - 0x0
      13'h1F6A: dout  = 8'b00000000; // 8042 :   0 - 0x0
      13'h1F6B: dout  = 8'b00000000; // 8043 :   0 - 0x0
      13'h1F6C: dout  = 8'b00000000; // 8044 :   0 - 0x0
      13'h1F6D: dout  = 8'b00000000; // 8045 :   0 - 0x0
      13'h1F6E: dout  = 8'b00000000; // 8046 :   0 - 0x0
      13'h1F6F: dout  = 8'b00000000; // 8047 :   0 - 0x0
      13'h1F70: dout  = 8'b10000111; // 8048 : 135 - 0x87 -- Background 0xf7
      13'h1F71: dout  = 8'b10000111; // 8049 : 135 - 0x87
      13'h1F72: dout  = 8'b10000011; // 8050 : 131 - 0x83
      13'h1F73: dout  = 8'b10000000; // 8051 : 128 - 0x80
      13'h1F74: dout  = 8'b10000000; // 8052 : 128 - 0x80
      13'h1F75: dout  = 8'b01000000; // 8053 :  64 - 0x40
      13'h1F76: dout  = 8'b00100000; // 8054 :  32 - 0x20
      13'h1F77: dout  = 8'b00011111; // 8055 :  31 - 0x1f
      13'h1F78: dout  = 8'b00000000; // 8056 :   0 - 0x0
      13'h1F79: dout  = 8'b00000000; // 8057 :   0 - 0x0
      13'h1F7A: dout  = 8'b00000000; // 8058 :   0 - 0x0
      13'h1F7B: dout  = 8'b00000000; // 8059 :   0 - 0x0
      13'h1F7C: dout  = 8'b00000000; // 8060 :   0 - 0x0
      13'h1F7D: dout  = 8'b10000000; // 8061 : 128 - 0x80
      13'h1F7E: dout  = 8'b11000000; // 8062 : 192 - 0xc0
      13'h1F7F: dout  = 8'b11100000; // 8063 : 224 - 0xe0
      13'h1F80: dout  = 8'b11100001; // 8064 : 225 - 0xe1 -- Background 0xf8
      13'h1F81: dout  = 8'b11100001; // 8065 : 225 - 0xe1
      13'h1F82: dout  = 8'b11000001; // 8066 : 193 - 0xc1
      13'h1F83: dout  = 8'b00000001; // 8067 :   1 - 0x1
      13'h1F84: dout  = 8'b00000001; // 8068 :   1 - 0x1
      13'h1F85: dout  = 8'b00000010; // 8069 :   2 - 0x2
      13'h1F86: dout  = 8'b00000100; // 8070 :   4 - 0x4
      13'h1F87: dout  = 8'b11111000; // 8071 : 248 - 0xf8
      13'h1F88: dout  = 8'b00000000; // 8072 :   0 - 0x0
      13'h1F89: dout  = 8'b00000000; // 8073 :   0 - 0x0
      13'h1F8A: dout  = 8'b00000000; // 8074 :   0 - 0x0
      13'h1F8B: dout  = 8'b00000000; // 8075 :   0 - 0x0
      13'h1F8C: dout  = 8'b00000000; // 8076 :   0 - 0x0
      13'h1F8D: dout  = 8'b00000001; // 8077 :   1 - 0x1
      13'h1F8E: dout  = 8'b00000011; // 8078 :   3 - 0x3
      13'h1F8F: dout  = 8'b00000111; // 8079 :   7 - 0x7
      13'h1F90: dout  = 8'b00000000; // 8080 :   0 - 0x0 -- Background 0xf9
      13'h1F91: dout  = 8'b00000010; // 8081 :   2 - 0x2
      13'h1F92: dout  = 8'b00000101; // 8082 :   5 - 0x5
      13'h1F93: dout  = 8'b00000000; // 8083 :   0 - 0x0
      13'h1F94: dout  = 8'b00100000; // 8084 :  32 - 0x20
      13'h1F95: dout  = 8'b01010000; // 8085 :  80 - 0x50
      13'h1F96: dout  = 8'b00000000; // 8086 :   0 - 0x0
      13'h1F97: dout  = 8'b00000000; // 8087 :   0 - 0x0
      13'h1F98: dout  = 8'b11111111; // 8088 : 255 - 0xff
      13'h1F99: dout  = 8'b11111111; // 8089 : 255 - 0xff
      13'h1F9A: dout  = 8'b11111111; // 8090 : 255 - 0xff
      13'h1F9B: dout  = 8'b11111111; // 8091 : 255 - 0xff
      13'h1F9C: dout  = 8'b11111111; // 8092 : 255 - 0xff
      13'h1F9D: dout  = 8'b11111111; // 8093 : 255 - 0xff
      13'h1F9E: dout  = 8'b11111111; // 8094 : 255 - 0xff
      13'h1F9F: dout  = 8'b11111111; // 8095 : 255 - 0xff
      13'h1FA0: dout  = 8'b00000000; // 8096 :   0 - 0x0 -- Background 0xfa
      13'h1FA1: dout  = 8'b00000000; // 8097 :   0 - 0x0
      13'h1FA2: dout  = 8'b00000000; // 8098 :   0 - 0x0
      13'h1FA3: dout  = 8'b00000000; // 8099 :   0 - 0x0
      13'h1FA4: dout  = 8'b00000000; // 8100 :   0 - 0x0
      13'h1FA5: dout  = 8'b00000000; // 8101 :   0 - 0x0
      13'h1FA6: dout  = 8'b00000000; // 8102 :   0 - 0x0
      13'h1FA7: dout  = 8'b00000000; // 8103 :   0 - 0x0
      13'h1FA8: dout  = 8'b11111111; // 8104 : 255 - 0xff
      13'h1FA9: dout  = 8'b11111111; // 8105 : 255 - 0xff
      13'h1FAA: dout  = 8'b11111111; // 8106 : 255 - 0xff
      13'h1FAB: dout  = 8'b11111111; // 8107 : 255 - 0xff
      13'h1FAC: dout  = 8'b11111111; // 8108 : 255 - 0xff
      13'h1FAD: dout  = 8'b11111111; // 8109 : 255 - 0xff
      13'h1FAE: dout  = 8'b11111111; // 8110 : 255 - 0xff
      13'h1FAF: dout  = 8'b11111111; // 8111 : 255 - 0xff
      13'h1FB0: dout  = 8'b11111111; // 8112 : 255 - 0xff -- Background 0xfb
      13'h1FB1: dout  = 8'b00000000; // 8113 :   0 - 0x0
      13'h1FB2: dout  = 8'b00000000; // 8114 :   0 - 0x0
      13'h1FB3: dout  = 8'b00000000; // 8115 :   0 - 0x0
      13'h1FB4: dout  = 8'b00000000; // 8116 :   0 - 0x0
      13'h1FB5: dout  = 8'b11111111; // 8117 : 255 - 0xff
      13'h1FB6: dout  = 8'b11111111; // 8118 : 255 - 0xff
      13'h1FB7: dout  = 8'b11111111; // 8119 : 255 - 0xff
      13'h1FB8: dout  = 8'b00000000; // 8120 :   0 - 0x0
      13'h1FB9: dout  = 8'b00000000; // 8121 :   0 - 0x0
      13'h1FBA: dout  = 8'b00000000; // 8122 :   0 - 0x0
      13'h1FBB: dout  = 8'b00000000; // 8123 :   0 - 0x0
      13'h1FBC: dout  = 8'b00000000; // 8124 :   0 - 0x0
      13'h1FBD: dout  = 8'b00000000; // 8125 :   0 - 0x0
      13'h1FBE: dout  = 8'b00000000; // 8126 :   0 - 0x0
      13'h1FBF: dout  = 8'b00000000; // 8127 :   0 - 0x0
      13'h1FC0: dout  = 8'b10000111; // 8128 : 135 - 0x87 -- Background 0xfc
      13'h1FC1: dout  = 8'b10000111; // 8129 : 135 - 0x87
      13'h1FC2: dout  = 8'b10000111; // 8130 : 135 - 0x87
      13'h1FC3: dout  = 8'b10000111; // 8131 : 135 - 0x87
      13'h1FC4: dout  = 8'b10000111; // 8132 : 135 - 0x87
      13'h1FC5: dout  = 8'b10000111; // 8133 : 135 - 0x87
      13'h1FC6: dout  = 8'b10000111; // 8134 : 135 - 0x87
      13'h1FC7: dout  = 8'b10000111; // 8135 : 135 - 0x87
      13'h1FC8: dout  = 8'b00000000; // 8136 :   0 - 0x0
      13'h1FC9: dout  = 8'b00000000; // 8137 :   0 - 0x0
      13'h1FCA: dout  = 8'b00000000; // 8138 :   0 - 0x0
      13'h1FCB: dout  = 8'b00000000; // 8139 :   0 - 0x0
      13'h1FCC: dout  = 8'b00000000; // 8140 :   0 - 0x0
      13'h1FCD: dout  = 8'b00000000; // 8141 :   0 - 0x0
      13'h1FCE: dout  = 8'b00000000; // 8142 :   0 - 0x0
      13'h1FCF: dout  = 8'b00000000; // 8143 :   0 - 0x0
      13'h1FD0: dout  = 8'b11111111; // 8144 : 255 - 0xff -- Background 0xfd
      13'h1FD1: dout  = 8'b11111111; // 8145 : 255 - 0xff
      13'h1FD2: dout  = 8'b11111111; // 8146 : 255 - 0xff
      13'h1FD3: dout  = 8'b11000011; // 8147 : 195 - 0xc3
      13'h1FD4: dout  = 8'b11000011; // 8148 : 195 - 0xc3
      13'h1FD5: dout  = 8'b11111111; // 8149 : 255 - 0xff
      13'h1FD6: dout  = 8'b11111111; // 8150 : 255 - 0xff
      13'h1FD7: dout  = 8'b11111111; // 8151 : 255 - 0xff
      13'h1FD8: dout  = 8'b00000000; // 8152 :   0 - 0x0
      13'h1FD9: dout  = 8'b00000000; // 8153 :   0 - 0x0
      13'h1FDA: dout  = 8'b00000000; // 8154 :   0 - 0x0
      13'h1FDB: dout  = 8'b00111100; // 8155 :  60 - 0x3c
      13'h1FDC: dout  = 8'b00111100; // 8156 :  60 - 0x3c
      13'h1FDD: dout  = 8'b00000000; // 8157 :   0 - 0x0
      13'h1FDE: dout  = 8'b00000000; // 8158 :   0 - 0x0
      13'h1FDF: dout  = 8'b00000000; // 8159 :   0 - 0x0
      13'h1FE0: dout  = 8'b11111111; // 8160 : 255 - 0xff -- Background 0xfe
      13'h1FE1: dout  = 8'b11111111; // 8161 : 255 - 0xff
      13'h1FE2: dout  = 8'b11100111; // 8162 : 231 - 0xe7
      13'h1FE3: dout  = 8'b11100111; // 8163 : 231 - 0xe7
      13'h1FE4: dout  = 8'b11100111; // 8164 : 231 - 0xe7
      13'h1FE5: dout  = 8'b11100111; // 8165 : 231 - 0xe7
      13'h1FE6: dout  = 8'b11111111; // 8166 : 255 - 0xff
      13'h1FE7: dout  = 8'b11111111; // 8167 : 255 - 0xff
      13'h1FE8: dout  = 8'b00000000; // 8168 :   0 - 0x0
      13'h1FE9: dout  = 8'b00000000; // 8169 :   0 - 0x0
      13'h1FEA: dout  = 8'b00011000; // 8170 :  24 - 0x18
      13'h1FEB: dout  = 8'b00011000; // 8171 :  24 - 0x18
      13'h1FEC: dout  = 8'b00011000; // 8172 :  24 - 0x18
      13'h1FED: dout  = 8'b00011000; // 8173 :  24 - 0x18
      13'h1FEE: dout  = 8'b00000000; // 8174 :   0 - 0x0
      13'h1FEF: dout  = 8'b00000000; // 8175 :   0 - 0x0
      13'h1FF0: dout  = 8'b11111111; // 8176 : 255 - 0xff -- Background 0xff
      13'h1FF1: dout  = 8'b11111111; // 8177 : 255 - 0xff
      13'h1FF2: dout  = 8'b11111111; // 8178 : 255 - 0xff
      13'h1FF3: dout  = 8'b11111111; // 8179 : 255 - 0xff
      13'h1FF4: dout  = 8'b11111111; // 8180 : 255 - 0xff
      13'h1FF5: dout  = 8'b11111111; // 8181 : 255 - 0xff
      13'h1FF6: dout  = 8'b11111111; // 8182 : 255 - 0xff
      13'h1FF7: dout  = 8'b11111111; // 8183 : 255 - 0xff
      13'h1FF8: dout  = 8'b00000000; // 8184 :   0 - 0x0
      13'h1FF9: dout  = 8'b00000000; // 8185 :   0 - 0x0
      13'h1FFA: dout  = 8'b00000000; // 8186 :   0 - 0x0
      13'h1FFB: dout  = 8'b00000000; // 8187 :   0 - 0x0
      13'h1FFC: dout  = 8'b00000000; // 8188 :   0 - 0x0
      13'h1FFD: dout  = 8'b00000000; // 8189 :   0 - 0x0
      13'h1FFE: dout  = 8'b00000000; // 8190 :   0 - 0x0
      13'h1FFF: dout  = 8'b00000000; // 8191 :   0 - 0x0
    endcase
  end

endmodule
