//- Autcmatically generated verilog ROM from a NES memory file----
//-   PATTERN TABLE WITH ONLY ONE COLOR PLANE
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


//-  Original memory dump file name: pacman_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_PTABLE_PACMAN_color1
  (
     //input     clk,   // clock
     input      [12-1:0] addr,  //4096 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                              //  address:   value 
                              //    dec  : dec - hex
          // Sprite pattern Table
      12'h0: dout  = 8'b00000000; //    0 :   0 - 0x0 -- Sprite 0x0
      12'h1: dout  = 8'b00000000; //    1 :   0 - 0x0
      12'h2: dout  = 8'b00000000; //    2 :   0 - 0x0
      12'h3: dout  = 8'b00000000; //    3 :   0 - 0x0
      12'h4: dout  = 8'b00000000; //    4 :   0 - 0x0
      12'h5: dout  = 8'b00000000; //    5 :   0 - 0x0
      12'h6: dout  = 8'b00000000; //    6 :   0 - 0x0
      12'h7: dout  = 8'b00000000; //    7 :   0 - 0x0
      12'h8: dout  = 8'b00000000; //    8 :   0 - 0x0 -- Sprite 0x1
      12'h9: dout  = 8'b00000000; //    9 :   0 - 0x0
      12'hA: dout  = 8'b00000000; //   10 :   0 - 0x0
      12'hB: dout  = 8'b00000000; //   11 :   0 - 0x0
      12'hC: dout  = 8'b00000000; //   12 :   0 - 0x0
      12'hD: dout  = 8'b00000000; //   13 :   0 - 0x0
      12'hE: dout  = 8'b00000000; //   14 :   0 - 0x0
      12'hF: dout  = 8'b00000000; //   15 :   0 - 0x0
      12'h10: dout  = 8'b00000000; //   16 :   0 - 0x0 -- Sprite 0x2
      12'h11: dout  = 8'b00000000; //   17 :   0 - 0x0
      12'h12: dout  = 8'b00000000; //   18 :   0 - 0x0
      12'h13: dout  = 8'b00000000; //   19 :   0 - 0x0
      12'h14: dout  = 8'b00000000; //   20 :   0 - 0x0
      12'h15: dout  = 8'b00000000; //   21 :   0 - 0x0
      12'h16: dout  = 8'b00000000; //   22 :   0 - 0x0
      12'h17: dout  = 8'b00000000; //   23 :   0 - 0x0
      12'h18: dout  = 8'b00000000; //   24 :   0 - 0x0 -- Sprite 0x3
      12'h19: dout  = 8'b00000000; //   25 :   0 - 0x0
      12'h1A: dout  = 8'b00000000; //   26 :   0 - 0x0
      12'h1B: dout  = 8'b00000000; //   27 :   0 - 0x0
      12'h1C: dout  = 8'b00000000; //   28 :   0 - 0x0
      12'h1D: dout  = 8'b00000000; //   29 :   0 - 0x0
      12'h1E: dout  = 8'b00000000; //   30 :   0 - 0x0
      12'h1F: dout  = 8'b00000000; //   31 :   0 - 0x0
      12'h20: dout  = 8'b00000000; //   32 :   0 - 0x0 -- Sprite 0x4
      12'h21: dout  = 8'b00000000; //   33 :   0 - 0x0
      12'h22: dout  = 8'b00000000; //   34 :   0 - 0x0
      12'h23: dout  = 8'b00000000; //   35 :   0 - 0x0
      12'h24: dout  = 8'b00000000; //   36 :   0 - 0x0
      12'h25: dout  = 8'b00000000; //   37 :   0 - 0x0
      12'h26: dout  = 8'b00000000; //   38 :   0 - 0x0
      12'h27: dout  = 8'b00000000; //   39 :   0 - 0x0
      12'h28: dout  = 8'b00000000; //   40 :   0 - 0x0 -- Sprite 0x5
      12'h29: dout  = 8'b00000000; //   41 :   0 - 0x0
      12'h2A: dout  = 8'b00000000; //   42 :   0 - 0x0
      12'h2B: dout  = 8'b00000000; //   43 :   0 - 0x0
      12'h2C: dout  = 8'b00000000; //   44 :   0 - 0x0
      12'h2D: dout  = 8'b00000000; //   45 :   0 - 0x0
      12'h2E: dout  = 8'b00000000; //   46 :   0 - 0x0
      12'h2F: dout  = 8'b00000000; //   47 :   0 - 0x0
      12'h30: dout  = 8'b00000000; //   48 :   0 - 0x0 -- Sprite 0x6
      12'h31: dout  = 8'b00000000; //   49 :   0 - 0x0
      12'h32: dout  = 8'b00000000; //   50 :   0 - 0x0
      12'h33: dout  = 8'b00000000; //   51 :   0 - 0x0
      12'h34: dout  = 8'b00000000; //   52 :   0 - 0x0
      12'h35: dout  = 8'b00000000; //   53 :   0 - 0x0
      12'h36: dout  = 8'b00000000; //   54 :   0 - 0x0
      12'h37: dout  = 8'b00000000; //   55 :   0 - 0x0
      12'h38: dout  = 8'b00000000; //   56 :   0 - 0x0 -- Sprite 0x7
      12'h39: dout  = 8'b00000000; //   57 :   0 - 0x0
      12'h3A: dout  = 8'b00000000; //   58 :   0 - 0x0
      12'h3B: dout  = 8'b00000000; //   59 :   0 - 0x0
      12'h3C: dout  = 8'b00000000; //   60 :   0 - 0x0
      12'h3D: dout  = 8'b00000000; //   61 :   0 - 0x0
      12'h3E: dout  = 8'b00000000; //   62 :   0 - 0x0
      12'h3F: dout  = 8'b00000000; //   63 :   0 - 0x0
      12'h40: dout  = 8'b00000000; //   64 :   0 - 0x0 -- Sprite 0x8
      12'h41: dout  = 8'b00000000; //   65 :   0 - 0x0
      12'h42: dout  = 8'b00000000; //   66 :   0 - 0x0
      12'h43: dout  = 8'b00000000; //   67 :   0 - 0x0
      12'h44: dout  = 8'b00000000; //   68 :   0 - 0x0
      12'h45: dout  = 8'b00000000; //   69 :   0 - 0x0
      12'h46: dout  = 8'b00000000; //   70 :   0 - 0x0
      12'h47: dout  = 8'b00000000; //   71 :   0 - 0x0
      12'h48: dout  = 8'b00000000; //   72 :   0 - 0x0 -- Sprite 0x9
      12'h49: dout  = 8'b00000000; //   73 :   0 - 0x0
      12'h4A: dout  = 8'b00000000; //   74 :   0 - 0x0
      12'h4B: dout  = 8'b00000000; //   75 :   0 - 0x0
      12'h4C: dout  = 8'b00000000; //   76 :   0 - 0x0
      12'h4D: dout  = 8'b00000000; //   77 :   0 - 0x0
      12'h4E: dout  = 8'b00000000; //   78 :   0 - 0x0
      12'h4F: dout  = 8'b00000000; //   79 :   0 - 0x0
      12'h50: dout  = 8'b00000000; //   80 :   0 - 0x0 -- Sprite 0xa
      12'h51: dout  = 8'b00000000; //   81 :   0 - 0x0
      12'h52: dout  = 8'b00000000; //   82 :   0 - 0x0
      12'h53: dout  = 8'b00000000; //   83 :   0 - 0x0
      12'h54: dout  = 8'b00000000; //   84 :   0 - 0x0
      12'h55: dout  = 8'b00000000; //   85 :   0 - 0x0
      12'h56: dout  = 8'b00000000; //   86 :   0 - 0x0
      12'h57: dout  = 8'b00000000; //   87 :   0 - 0x0
      12'h58: dout  = 8'b00000000; //   88 :   0 - 0x0 -- Sprite 0xb
      12'h59: dout  = 8'b00000000; //   89 :   0 - 0x0
      12'h5A: dout  = 8'b00000000; //   90 :   0 - 0x0
      12'h5B: dout  = 8'b00000000; //   91 :   0 - 0x0
      12'h5C: dout  = 8'b00000000; //   92 :   0 - 0x0
      12'h5D: dout  = 8'b00000000; //   93 :   0 - 0x0
      12'h5E: dout  = 8'b00000000; //   94 :   0 - 0x0
      12'h5F: dout  = 8'b00000000; //   95 :   0 - 0x0
      12'h60: dout  = 8'b00000000; //   96 :   0 - 0x0 -- Sprite 0xc
      12'h61: dout  = 8'b00000000; //   97 :   0 - 0x0
      12'h62: dout  = 8'b00000000; //   98 :   0 - 0x0
      12'h63: dout  = 8'b00000000; //   99 :   0 - 0x0
      12'h64: dout  = 8'b00000000; //  100 :   0 - 0x0
      12'h65: dout  = 8'b00000000; //  101 :   0 - 0x0
      12'h66: dout  = 8'b00000000; //  102 :   0 - 0x0
      12'h67: dout  = 8'b00000000; //  103 :   0 - 0x0
      12'h68: dout  = 8'b00000000; //  104 :   0 - 0x0 -- Sprite 0xd
      12'h69: dout  = 8'b00000000; //  105 :   0 - 0x0
      12'h6A: dout  = 8'b00000000; //  106 :   0 - 0x0
      12'h6B: dout  = 8'b00000000; //  107 :   0 - 0x0
      12'h6C: dout  = 8'b00000000; //  108 :   0 - 0x0
      12'h6D: dout  = 8'b00000000; //  109 :   0 - 0x0
      12'h6E: dout  = 8'b00000000; //  110 :   0 - 0x0
      12'h6F: dout  = 8'b00000000; //  111 :   0 - 0x0
      12'h70: dout  = 8'b00000000; //  112 :   0 - 0x0 -- Sprite 0xe
      12'h71: dout  = 8'b00000000; //  113 :   0 - 0x0
      12'h72: dout  = 8'b00000000; //  114 :   0 - 0x0
      12'h73: dout  = 8'b00000000; //  115 :   0 - 0x0
      12'h74: dout  = 8'b00000000; //  116 :   0 - 0x0
      12'h75: dout  = 8'b00000000; //  117 :   0 - 0x0
      12'h76: dout  = 8'b00000000; //  118 :   0 - 0x0
      12'h77: dout  = 8'b00000000; //  119 :   0 - 0x0
      12'h78: dout  = 8'b00000000; //  120 :   0 - 0x0 -- Sprite 0xf
      12'h79: dout  = 8'b00000000; //  121 :   0 - 0x0
      12'h7A: dout  = 8'b00000000; //  122 :   0 - 0x0
      12'h7B: dout  = 8'b00000000; //  123 :   0 - 0x0
      12'h7C: dout  = 8'b00000000; //  124 :   0 - 0x0
      12'h7D: dout  = 8'b00000000; //  125 :   0 - 0x0
      12'h7E: dout  = 8'b00000000; //  126 :   0 - 0x0
      12'h7F: dout  = 8'b00000000; //  127 :   0 - 0x0
      12'h80: dout  = 8'b00000000; //  128 :   0 - 0x0 -- Sprite 0x10
      12'h81: dout  = 8'b00000000; //  129 :   0 - 0x0
      12'h82: dout  = 8'b00000000; //  130 :   0 - 0x0
      12'h83: dout  = 8'b00000000; //  131 :   0 - 0x0
      12'h84: dout  = 8'b00000000; //  132 :   0 - 0x0
      12'h85: dout  = 8'b00000000; //  133 :   0 - 0x0
      12'h86: dout  = 8'b00000000; //  134 :   0 - 0x0
      12'h87: dout  = 8'b00000000; //  135 :   0 - 0x0
      12'h88: dout  = 8'b00000000; //  136 :   0 - 0x0 -- Sprite 0x11
      12'h89: dout  = 8'b00000000; //  137 :   0 - 0x0
      12'h8A: dout  = 8'b00000000; //  138 :   0 - 0x0
      12'h8B: dout  = 8'b00000000; //  139 :   0 - 0x0
      12'h8C: dout  = 8'b00000000; //  140 :   0 - 0x0
      12'h8D: dout  = 8'b00000000; //  141 :   0 - 0x0
      12'h8E: dout  = 8'b00000000; //  142 :   0 - 0x0
      12'h8F: dout  = 8'b00000000; //  143 :   0 - 0x0
      12'h90: dout  = 8'b00000000; //  144 :   0 - 0x0 -- Sprite 0x12
      12'h91: dout  = 8'b00000000; //  145 :   0 - 0x0
      12'h92: dout  = 8'b00000000; //  146 :   0 - 0x0
      12'h93: dout  = 8'b00000000; //  147 :   0 - 0x0
      12'h94: dout  = 8'b00000000; //  148 :   0 - 0x0
      12'h95: dout  = 8'b00000000; //  149 :   0 - 0x0
      12'h96: dout  = 8'b00000000; //  150 :   0 - 0x0
      12'h97: dout  = 8'b00000000; //  151 :   0 - 0x0
      12'h98: dout  = 8'b00000000; //  152 :   0 - 0x0 -- Sprite 0x13
      12'h99: dout  = 8'b00000000; //  153 :   0 - 0x0
      12'h9A: dout  = 8'b00000000; //  154 :   0 - 0x0
      12'h9B: dout  = 8'b00000000; //  155 :   0 - 0x0
      12'h9C: dout  = 8'b00000000; //  156 :   0 - 0x0
      12'h9D: dout  = 8'b00000000; //  157 :   0 - 0x0
      12'h9E: dout  = 8'b00000000; //  158 :   0 - 0x0
      12'h9F: dout  = 8'b00000000; //  159 :   0 - 0x0
      12'hA0: dout  = 8'b00000000; //  160 :   0 - 0x0 -- Sprite 0x14
      12'hA1: dout  = 8'b00000000; //  161 :   0 - 0x0
      12'hA2: dout  = 8'b00000000; //  162 :   0 - 0x0
      12'hA3: dout  = 8'b00000000; //  163 :   0 - 0x0
      12'hA4: dout  = 8'b00000000; //  164 :   0 - 0x0
      12'hA5: dout  = 8'b00000000; //  165 :   0 - 0x0
      12'hA6: dout  = 8'b00000000; //  166 :   0 - 0x0
      12'hA7: dout  = 8'b00000000; //  167 :   0 - 0x0
      12'hA8: dout  = 8'b00000000; //  168 :   0 - 0x0 -- Sprite 0x15
      12'hA9: dout  = 8'b00000000; //  169 :   0 - 0x0
      12'hAA: dout  = 8'b00000000; //  170 :   0 - 0x0
      12'hAB: dout  = 8'b00000000; //  171 :   0 - 0x0
      12'hAC: dout  = 8'b00000000; //  172 :   0 - 0x0
      12'hAD: dout  = 8'b00000000; //  173 :   0 - 0x0
      12'hAE: dout  = 8'b00000000; //  174 :   0 - 0x0
      12'hAF: dout  = 8'b00000000; //  175 :   0 - 0x0
      12'hB0: dout  = 8'b00000000; //  176 :   0 - 0x0 -- Sprite 0x16
      12'hB1: dout  = 8'b00000000; //  177 :   0 - 0x0
      12'hB2: dout  = 8'b00000000; //  178 :   0 - 0x0
      12'hB3: dout  = 8'b00000000; //  179 :   0 - 0x0
      12'hB4: dout  = 8'b00000000; //  180 :   0 - 0x0
      12'hB5: dout  = 8'b00000000; //  181 :   0 - 0x0
      12'hB6: dout  = 8'b00000000; //  182 :   0 - 0x0
      12'hB7: dout  = 8'b00000000; //  183 :   0 - 0x0
      12'hB8: dout  = 8'b00000000; //  184 :   0 - 0x0 -- Sprite 0x17
      12'hB9: dout  = 8'b00000000; //  185 :   0 - 0x0
      12'hBA: dout  = 8'b00000000; //  186 :   0 - 0x0
      12'hBB: dout  = 8'b00000000; //  187 :   0 - 0x0
      12'hBC: dout  = 8'b00000000; //  188 :   0 - 0x0
      12'hBD: dout  = 8'b00000000; //  189 :   0 - 0x0
      12'hBE: dout  = 8'b00000000; //  190 :   0 - 0x0
      12'hBF: dout  = 8'b00000000; //  191 :   0 - 0x0
      12'hC0: dout  = 8'b00000000; //  192 :   0 - 0x0 -- Sprite 0x18
      12'hC1: dout  = 8'b00000000; //  193 :   0 - 0x0
      12'hC2: dout  = 8'b00000011; //  194 :   3 - 0x3
      12'hC3: dout  = 8'b00000011; //  195 :   3 - 0x3
      12'hC4: dout  = 8'b00010011; //  196 :  19 - 0x13
      12'hC5: dout  = 8'b00111111; //  197 :  63 - 0x3f
      12'hC6: dout  = 8'b00111111; //  198 :  63 - 0x3f
      12'hC7: dout  = 8'b01111111; //  199 : 127 - 0x7f
      12'hC8: dout  = 8'b01111111; //  200 : 127 - 0x7f -- Sprite 0x19
      12'hC9: dout  = 8'b01111111; //  201 : 127 - 0x7f
      12'hCA: dout  = 8'b01111111; //  202 : 127 - 0x7f
      12'hCB: dout  = 8'b01111111; //  203 : 127 - 0x7f
      12'hCC: dout  = 8'b01101110; //  204 : 110 - 0x6e
      12'hCD: dout  = 8'b01000110; //  205 :  70 - 0x46
      12'hCE: dout  = 8'b00000000; //  206 :   0 - 0x0
      12'hCF: dout  = 8'b00000000; //  207 :   0 - 0x0
      12'hD0: dout  = 8'b01111111; //  208 : 127 - 0x7f -- Sprite 0x1a
      12'hD1: dout  = 8'b01111111; //  209 : 127 - 0x7f
      12'hD2: dout  = 8'b01111111; //  210 : 127 - 0x7f
      12'hD3: dout  = 8'b01111111; //  211 : 127 - 0x7f
      12'hD4: dout  = 8'b01111011; //  212 : 123 - 0x7b
      12'hD5: dout  = 8'b00110001; //  213 :  49 - 0x31
      12'hD6: dout  = 8'b00000000; //  214 :   0 - 0x0
      12'hD7: dout  = 8'b00000000; //  215 :   0 - 0x0
      12'hD8: dout  = 8'b00000000; //  216 :   0 - 0x0 -- Sprite 0x1b
      12'hD9: dout  = 8'b00000011; //  217 :   3 - 0x3
      12'hDA: dout  = 8'b00001111; //  218 :  15 - 0xf
      12'hDB: dout  = 8'b00011111; //  219 :  31 - 0x1f
      12'hDC: dout  = 8'b00111111; //  220 :  63 - 0x3f
      12'hDD: dout  = 8'b00111111; //  221 :  63 - 0x3f
      12'hDE: dout  = 8'b00001111; //  222 :  15 - 0xf
      12'hDF: dout  = 8'b01001111; //  223 :  79 - 0x4f
      12'hE0: dout  = 8'b00000000; //  224 :   0 - 0x0 -- Sprite 0x1c
      12'hE1: dout  = 8'b11000000; //  225 : 192 - 0xc0
      12'hE2: dout  = 8'b11110000; //  226 : 240 - 0xf0
      12'hE3: dout  = 8'b11111000; //  227 : 248 - 0xf8
      12'hE4: dout  = 8'b11111100; //  228 : 252 - 0xfc
      12'hE5: dout  = 8'b11111100; //  229 : 252 - 0xfc
      12'hE6: dout  = 8'b00111100; //  230 :  60 - 0x3c
      12'hE7: dout  = 8'b00111110; //  231 :  62 - 0x3e
      12'hE8: dout  = 8'b01111111; //  232 : 127 - 0x7f -- Sprite 0x1d
      12'hE9: dout  = 8'b01111111; //  233 : 127 - 0x7f
      12'hEA: dout  = 8'b01111111; //  234 : 127 - 0x7f
      12'hEB: dout  = 8'b01111111; //  235 : 127 - 0x7f
      12'hEC: dout  = 8'b01101110; //  236 : 110 - 0x6e
      12'hED: dout  = 8'b01000110; //  237 :  70 - 0x46
      12'hEE: dout  = 8'b00000000; //  238 :   0 - 0x0
      12'hEF: dout  = 8'b00000000; //  239 :   0 - 0x0
      12'hF0: dout  = 8'b01111111; //  240 : 127 - 0x7f -- Sprite 0x1e
      12'hF1: dout  = 8'b01111111; //  241 : 127 - 0x7f
      12'hF2: dout  = 8'b01111111; //  242 : 127 - 0x7f
      12'hF3: dout  = 8'b01111111; //  243 : 127 - 0x7f
      12'hF4: dout  = 8'b01111011; //  244 : 123 - 0x7b
      12'hF5: dout  = 8'b00110001; //  245 :  49 - 0x31
      12'hF6: dout  = 8'b00000000; //  246 :   0 - 0x0
      12'hF7: dout  = 8'b00000000; //  247 :   0 - 0x0
      12'hF8: dout  = 8'b11111110; //  248 : 254 - 0xfe -- Sprite 0x1f
      12'hF9: dout  = 8'b11111110; //  249 : 254 - 0xfe
      12'hFA: dout  = 8'b11111110; //  250 : 254 - 0xfe
      12'hFB: dout  = 8'b11111110; //  251 : 254 - 0xfe
      12'hFC: dout  = 8'b01110110; //  252 : 118 - 0x76
      12'hFD: dout  = 8'b01100010; //  253 :  98 - 0x62
      12'hFE: dout  = 8'b00000000; //  254 :   0 - 0x0
      12'hFF: dout  = 8'b00000000; //  255 :   0 - 0x0
      12'h100: dout  = 8'b11111110; //  256 : 254 - 0xfe -- Sprite 0x20
      12'h101: dout  = 8'b11111110; //  257 : 254 - 0xfe
      12'h102: dout  = 8'b11111110; //  258 : 254 - 0xfe
      12'h103: dout  = 8'b11111110; //  259 : 254 - 0xfe
      12'h104: dout  = 8'b11011110; //  260 : 222 - 0xde
      12'h105: dout  = 8'b10001100; //  261 : 140 - 0x8c
      12'h106: dout  = 8'b00000000; //  262 :   0 - 0x0
      12'h107: dout  = 8'b00000000; //  263 :   0 - 0x0
      12'h108: dout  = 8'b00000000; //  264 :   0 - 0x0 -- Sprite 0x21
      12'h109: dout  = 8'b00000011; //  265 :   3 - 0x3
      12'h10A: dout  = 8'b00001111; //  266 :  15 - 0xf
      12'h10B: dout  = 8'b00011111; //  267 :  31 - 0x1f
      12'h10C: dout  = 8'b00111111; //  268 :  63 - 0x3f
      12'h10D: dout  = 8'b00111111; //  269 :  63 - 0x3f
      12'h10E: dout  = 8'b00111111; //  270 :  63 - 0x3f
      12'h10F: dout  = 8'b01111111; //  271 : 127 - 0x7f
      12'h110: dout  = 8'b01110011; //  272 : 115 - 0x73 -- Sprite 0x22
      12'h111: dout  = 8'b01110011; //  273 : 115 - 0x73
      12'h112: dout  = 8'b01111111; //  274 : 127 - 0x7f
      12'h113: dout  = 8'b01111111; //  275 : 127 - 0x7f
      12'h114: dout  = 8'b01101110; //  276 : 110 - 0x6e
      12'h115: dout  = 8'b01000110; //  277 :  70 - 0x46
      12'h116: dout  = 8'b00000000; //  278 :   0 - 0x0
      12'h117: dout  = 8'b00000000; //  279 :   0 - 0x0
      12'h118: dout  = 8'b01110011; //  280 : 115 - 0x73 -- Sprite 0x23
      12'h119: dout  = 8'b01110011; //  281 : 115 - 0x73
      12'h11A: dout  = 8'b01111111; //  282 : 127 - 0x7f
      12'h11B: dout  = 8'b01111111; //  283 : 127 - 0x7f
      12'h11C: dout  = 8'b01110111; //  284 : 119 - 0x77
      12'h11D: dout  = 8'b00100011; //  285 :  35 - 0x23
      12'h11E: dout  = 8'b00000000; //  286 :   0 - 0x0
      12'h11F: dout  = 8'b00000000; //  287 :   0 - 0x0
      12'h120: dout  = 8'b00000000; //  288 :   0 - 0x0 -- Sprite 0x24
      12'h121: dout  = 8'b00000000; //  289 :   0 - 0x0
      12'h122: dout  = 8'b00000000; //  290 :   0 - 0x0
      12'h123: dout  = 8'b00000000; //  291 :   0 - 0x0
      12'h124: dout  = 8'b00000000; //  292 :   0 - 0x0
      12'h125: dout  = 8'b00000110; //  293 :   6 - 0x6
      12'h126: dout  = 8'b00000110; //  294 :   6 - 0x6
      12'h127: dout  = 8'b00000000; //  295 :   0 - 0x0
      12'h128: dout  = 8'b00000000; //  296 :   0 - 0x0 -- Sprite 0x25
      12'h129: dout  = 8'b00011001; //  297 :  25 - 0x19
      12'h12A: dout  = 8'b00100110; //  298 :  38 - 0x26
      12'h12B: dout  = 8'b00000000; //  299 :   0 - 0x0
      12'h12C: dout  = 8'b00000000; //  300 :   0 - 0x0
      12'h12D: dout  = 8'b00000000; //  301 :   0 - 0x0
      12'h12E: dout  = 8'b00000000; //  302 :   0 - 0x0
      12'h12F: dout  = 8'b00000000; //  303 :   0 - 0x0
      12'h130: dout  = 8'b00000000; //  304 :   0 - 0x0 -- Sprite 0x26
      12'h131: dout  = 8'b00011001; //  305 :  25 - 0x19
      12'h132: dout  = 8'b00100110; //  306 :  38 - 0x26
      12'h133: dout  = 8'b00000000; //  307 :   0 - 0x0
      12'h134: dout  = 8'b00000000; //  308 :   0 - 0x0
      12'h135: dout  = 8'b00000000; //  309 :   0 - 0x0
      12'h136: dout  = 8'b00000000; //  310 :   0 - 0x0
      12'h137: dout  = 8'b00000000; //  311 :   0 - 0x0
      12'h138: dout  = 8'b00000000; //  312 :   0 - 0x0 -- Sprite 0x27
      12'h139: dout  = 8'b00001100; //  313 :  12 - 0xc
      12'h13A: dout  = 8'b00010010; //  314 :  18 - 0x12
      12'h13B: dout  = 8'b00010010; //  315 :  18 - 0x12
      12'h13C: dout  = 8'b00011110; //  316 :  30 - 0x1e
      12'h13D: dout  = 8'b00001100; //  317 :  12 - 0xc
      12'h13E: dout  = 8'b00000000; //  318 :   0 - 0x0
      12'h13F: dout  = 8'b00000000; //  319 :   0 - 0x0
      12'h140: dout  = 8'b00000000; //  320 :   0 - 0x0 -- Sprite 0x28
      12'h141: dout  = 8'b00000000; //  321 :   0 - 0x0
      12'h142: dout  = 8'b00000000; //  322 :   0 - 0x0
      12'h143: dout  = 8'b00000000; //  323 :   0 - 0x0
      12'h144: dout  = 8'b00000000; //  324 :   0 - 0x0
      12'h145: dout  = 8'b00111000; //  325 :  56 - 0x38
      12'h146: dout  = 8'b01001101; //  326 :  77 - 0x4d
      12'h147: dout  = 8'b01001101; //  327 :  77 - 0x4d
      12'h148: dout  = 8'b00000000; //  328 :   0 - 0x0 -- Sprite 0x29
      12'h149: dout  = 8'b00000000; //  329 :   0 - 0x0
      12'h14A: dout  = 8'b00000000; //  330 :   0 - 0x0
      12'h14B: dout  = 8'b00000000; //  331 :   0 - 0x0
      12'h14C: dout  = 8'b00000000; //  332 :   0 - 0x0
      12'h14D: dout  = 8'b11100000; //  333 : 224 - 0xe0
      12'h14E: dout  = 8'b00110000; //  334 :  48 - 0x30
      12'h14F: dout  = 8'b00110000; //  335 :  48 - 0x30
      12'h150: dout  = 8'b00111000; //  336 :  56 - 0x38 -- Sprite 0x2a
      12'h151: dout  = 8'b00000000; //  337 :   0 - 0x0
      12'h152: dout  = 8'b00000000; //  338 :   0 - 0x0
      12'h153: dout  = 8'b00000000; //  339 :   0 - 0x0
      12'h154: dout  = 8'b00000000; //  340 :   0 - 0x0
      12'h155: dout  = 8'b00000000; //  341 :   0 - 0x0
      12'h156: dout  = 8'b00000000; //  342 :   0 - 0x0
      12'h157: dout  = 8'b00000000; //  343 :   0 - 0x0
      12'h158: dout  = 8'b11100000; //  344 : 224 - 0xe0 -- Sprite 0x2b
      12'h159: dout  = 8'b00000000; //  345 :   0 - 0x0
      12'h15A: dout  = 8'b00000000; //  346 :   0 - 0x0
      12'h15B: dout  = 8'b00000000; //  347 :   0 - 0x0
      12'h15C: dout  = 8'b00000000; //  348 :   0 - 0x0
      12'h15D: dout  = 8'b00000000; //  349 :   0 - 0x0
      12'h15E: dout  = 8'b00000000; //  350 :   0 - 0x0
      12'h15F: dout  = 8'b00000000; //  351 :   0 - 0x0
      12'h160: dout  = 8'b00000000; //  352 :   0 - 0x0 -- Sprite 0x2c
      12'h161: dout  = 8'b00000000; //  353 :   0 - 0x0
      12'h162: dout  = 8'b00000000; //  354 :   0 - 0x0
      12'h163: dout  = 8'b00000000; //  355 :   0 - 0x0
      12'h164: dout  = 8'b00000000; //  356 :   0 - 0x0
      12'h165: dout  = 8'b00000000; //  357 :   0 - 0x0
      12'h166: dout  = 8'b00001100; //  358 :  12 - 0xc
      12'h167: dout  = 8'b00011110; //  359 :  30 - 0x1e
      12'h168: dout  = 8'b00010010; //  360 :  18 - 0x12 -- Sprite 0x2d
      12'h169: dout  = 8'b00010010; //  361 :  18 - 0x12
      12'h16A: dout  = 8'b00001100; //  362 :  12 - 0xc
      12'h16B: dout  = 8'b00000000; //  363 :   0 - 0x0
      12'h16C: dout  = 8'b00000000; //  364 :   0 - 0x0
      12'h16D: dout  = 8'b00000000; //  365 :   0 - 0x0
      12'h16E: dout  = 8'b00000000; //  366 :   0 - 0x0
      12'h16F: dout  = 8'b00000000; //  367 :   0 - 0x0
      12'h170: dout  = 8'b00000000; //  368 :   0 - 0x0 -- Sprite 0x2e
      12'h171: dout  = 8'b00000000; //  369 :   0 - 0x0
      12'h172: dout  = 8'b00000000; //  370 :   0 - 0x0
      12'h173: dout  = 8'b00010001; //  371 :  17 - 0x11
      12'h174: dout  = 8'b00110010; //  372 :  50 - 0x32
      12'h175: dout  = 8'b00010010; //  373 :  18 - 0x12
      12'h176: dout  = 8'b00010010; //  374 :  18 - 0x12
      12'h177: dout  = 8'b00010010; //  375 :  18 - 0x12
      12'h178: dout  = 8'b00000000; //  376 :   0 - 0x0 -- Sprite 0x2f
      12'h179: dout  = 8'b00000000; //  377 :   0 - 0x0
      12'h17A: dout  = 8'b00000000; //  378 :   0 - 0x0
      12'h17B: dout  = 8'b10001100; //  379 : 140 - 0x8c
      12'h17C: dout  = 8'b01010010; //  380 :  82 - 0x52
      12'h17D: dout  = 8'b01010010; //  381 :  82 - 0x52
      12'h17E: dout  = 8'b01010010; //  382 :  82 - 0x52
      12'h17F: dout  = 8'b01010010; //  383 :  82 - 0x52
      12'h180: dout  = 8'b00010010; //  384 :  18 - 0x12 -- Sprite 0x30
      12'h181: dout  = 8'b00111001; //  385 :  57 - 0x39
      12'h182: dout  = 8'b00000000; //  386 :   0 - 0x0
      12'h183: dout  = 8'b00000000; //  387 :   0 - 0x0
      12'h184: dout  = 8'b00000000; //  388 :   0 - 0x0
      12'h185: dout  = 8'b00000000; //  389 :   0 - 0x0
      12'h186: dout  = 8'b00000000; //  390 :   0 - 0x0
      12'h187: dout  = 8'b00000000; //  391 :   0 - 0x0
      12'h188: dout  = 8'b01010010; //  392 :  82 - 0x52 -- Sprite 0x31
      12'h189: dout  = 8'b10001100; //  393 : 140 - 0x8c
      12'h18A: dout  = 8'b00000000; //  394 :   0 - 0x0
      12'h18B: dout  = 8'b00000000; //  395 :   0 - 0x0
      12'h18C: dout  = 8'b00000000; //  396 :   0 - 0x0
      12'h18D: dout  = 8'b00000000; //  397 :   0 - 0x0
      12'h18E: dout  = 8'b00000000; //  398 :   0 - 0x0
      12'h18F: dout  = 8'b00000000; //  399 :   0 - 0x0
      12'h190: dout  = 8'b00000000; //  400 :   0 - 0x0 -- Sprite 0x32
      12'h191: dout  = 8'b00000000; //  401 :   0 - 0x0
      12'h192: dout  = 8'b00000000; //  402 :   0 - 0x0
      12'h193: dout  = 8'b01110001; //  403 : 113 - 0x71
      12'h194: dout  = 8'b10001010; //  404 : 138 - 0x8a
      12'h195: dout  = 8'b00001010; //  405 :  10 - 0xa
      12'h196: dout  = 8'b00010010; //  406 :  18 - 0x12
      12'h197: dout  = 8'b00100010; //  407 :  34 - 0x22
      12'h198: dout  = 8'b01000010; //  408 :  66 - 0x42 -- Sprite 0x33
      12'h199: dout  = 8'b11111001; //  409 : 249 - 0xf9
      12'h19A: dout  = 8'b00000000; //  410 :   0 - 0x0
      12'h19B: dout  = 8'b00000000; //  411 :   0 - 0x0
      12'h19C: dout  = 8'b00000000; //  412 :   0 - 0x0
      12'h19D: dout  = 8'b00000000; //  413 :   0 - 0x0
      12'h19E: dout  = 8'b00000000; //  414 :   0 - 0x0
      12'h19F: dout  = 8'b00000000; //  415 :   0 - 0x0
      12'h1A0: dout  = 8'b00000000; //  416 :   0 - 0x0 -- Sprite 0x34
      12'h1A1: dout  = 8'b00000000; //  417 :   0 - 0x0
      12'h1A2: dout  = 8'b00000000; //  418 :   0 - 0x0
      12'h1A3: dout  = 8'b00110001; //  419 :  49 - 0x31
      12'h1A4: dout  = 8'b01001010; //  420 :  74 - 0x4a
      12'h1A5: dout  = 8'b00001010; //  421 :  10 - 0xa
      12'h1A6: dout  = 8'b00110010; //  422 :  50 - 0x32
      12'h1A7: dout  = 8'b00001010; //  423 :  10 - 0xa
      12'h1A8: dout  = 8'b01001010; //  424 :  74 - 0x4a -- Sprite 0x35
      12'h1A9: dout  = 8'b00110001; //  425 :  49 - 0x31
      12'h1AA: dout  = 8'b00000000; //  426 :   0 - 0x0
      12'h1AB: dout  = 8'b00000000; //  427 :   0 - 0x0
      12'h1AC: dout  = 8'b00000000; //  428 :   0 - 0x0
      12'h1AD: dout  = 8'b00000000; //  429 :   0 - 0x0
      12'h1AE: dout  = 8'b00000000; //  430 :   0 - 0x0
      12'h1AF: dout  = 8'b00000000; //  431 :   0 - 0x0
      12'h1B0: dout  = 8'b00000000; //  432 :   0 - 0x0 -- Sprite 0x36
      12'h1B1: dout  = 8'b00000000; //  433 :   0 - 0x0
      12'h1B2: dout  = 8'b00000000; //  434 :   0 - 0x0
      12'h1B3: dout  = 8'b00010001; //  435 :  17 - 0x11
      12'h1B4: dout  = 8'b00110010; //  436 :  50 - 0x32
      12'h1B5: dout  = 8'b01010010; //  437 :  82 - 0x52
      12'h1B6: dout  = 8'b10010010; //  438 : 146 - 0x92
      12'h1B7: dout  = 8'b11111010; //  439 : 250 - 0xfa
      12'h1B8: dout  = 8'b00010010; //  440 :  18 - 0x12 -- Sprite 0x37
      12'h1B9: dout  = 8'b00010001; //  441 :  17 - 0x11
      12'h1BA: dout  = 8'b00000000; //  442 :   0 - 0x0
      12'h1BB: dout  = 8'b00000000; //  443 :   0 - 0x0
      12'h1BC: dout  = 8'b00000000; //  444 :   0 - 0x0
      12'h1BD: dout  = 8'b00000000; //  445 :   0 - 0x0
      12'h1BE: dout  = 8'b00000000; //  446 :   0 - 0x0
      12'h1BF: dout  = 8'b00000000; //  447 :   0 - 0x0
      12'h1C0: dout  = 8'b00000000; //  448 :   0 - 0x0 -- Sprite 0x38
      12'h1C1: dout  = 8'b00000000; //  449 :   0 - 0x0
      12'h1C2: dout  = 8'b00000000; //  450 :   0 - 0x0
      12'h1C3: dout  = 8'b01110001; //  451 : 113 - 0x71
      12'h1C4: dout  = 8'b01000010; //  452 :  66 - 0x42
      12'h1C5: dout  = 8'b01000010; //  453 :  66 - 0x42
      12'h1C6: dout  = 8'b01110010; //  454 : 114 - 0x72
      12'h1C7: dout  = 8'b00001010; //  455 :  10 - 0xa
      12'h1C8: dout  = 8'b00001010; //  456 :  10 - 0xa -- Sprite 0x39
      12'h1C9: dout  = 8'b01110001; //  457 : 113 - 0x71
      12'h1CA: dout  = 8'b00000000; //  458 :   0 - 0x0
      12'h1CB: dout  = 8'b00000000; //  459 :   0 - 0x0
      12'h1CC: dout  = 8'b00000000; //  460 :   0 - 0x0
      12'h1CD: dout  = 8'b00000000; //  461 :   0 - 0x0
      12'h1CE: dout  = 8'b00000000; //  462 :   0 - 0x0
      12'h1CF: dout  = 8'b00000000; //  463 :   0 - 0x0
      12'h1D0: dout  = 8'b00000000; //  464 :   0 - 0x0 -- Sprite 0x3a
      12'h1D1: dout  = 8'b00000000; //  465 :   0 - 0x0
      12'h1D2: dout  = 8'b00000000; //  466 :   0 - 0x0
      12'h1D3: dout  = 8'b01110001; //  467 : 113 - 0x71
      12'h1D4: dout  = 8'b00001010; //  468 :  10 - 0xa
      12'h1D5: dout  = 8'b00010010; //  469 :  18 - 0x12
      12'h1D6: dout  = 8'b00010010; //  470 :  18 - 0x12
      12'h1D7: dout  = 8'b00100010; //  471 :  34 - 0x22
      12'h1D8: dout  = 8'b00100010; //  472 :  34 - 0x22 -- Sprite 0x3b
      12'h1D9: dout  = 8'b00100001; //  473 :  33 - 0x21
      12'h1DA: dout  = 8'b00000000; //  474 :   0 - 0x0
      12'h1DB: dout  = 8'b00000000; //  475 :   0 - 0x0
      12'h1DC: dout  = 8'b00000000; //  476 :   0 - 0x0
      12'h1DD: dout  = 8'b00000000; //  477 :   0 - 0x0
      12'h1DE: dout  = 8'b00000000; //  478 :   0 - 0x0
      12'h1DF: dout  = 8'b00000000; //  479 :   0 - 0x0
      12'h1E0: dout  = 8'b00000000; //  480 :   0 - 0x0 -- Sprite 0x3c
      12'h1E1: dout  = 8'b00000000; //  481 :   0 - 0x0
      12'h1E2: dout  = 8'b00000000; //  482 :   0 - 0x0
      12'h1E3: dout  = 8'b01110001; //  483 : 113 - 0x71
      12'h1E4: dout  = 8'b10001010; //  484 : 138 - 0x8a
      12'h1E5: dout  = 8'b10001010; //  485 : 138 - 0x8a
      12'h1E6: dout  = 8'b01110010; //  486 : 114 - 0x72
      12'h1E7: dout  = 8'b10001010; //  487 : 138 - 0x8a
      12'h1E8: dout  = 8'b10001010; //  488 : 138 - 0x8a -- Sprite 0x3d
      12'h1E9: dout  = 8'b01110001; //  489 : 113 - 0x71
      12'h1EA: dout  = 8'b00000000; //  490 :   0 - 0x0
      12'h1EB: dout  = 8'b00000000; //  491 :   0 - 0x0
      12'h1EC: dout  = 8'b00000000; //  492 :   0 - 0x0
      12'h1ED: dout  = 8'b00000000; //  493 :   0 - 0x0
      12'h1EE: dout  = 8'b00000000; //  494 :   0 - 0x0
      12'h1EF: dout  = 8'b00000000; //  495 :   0 - 0x0
      12'h1F0: dout  = 8'b00000000; //  496 :   0 - 0x0 -- Sprite 0x3e
      12'h1F1: dout  = 8'b00000000; //  497 :   0 - 0x0
      12'h1F2: dout  = 8'b00000000; //  498 :   0 - 0x0
      12'h1F3: dout  = 8'b10011000; //  499 : 152 - 0x98
      12'h1F4: dout  = 8'b10100101; //  500 : 165 - 0xa5
      12'h1F5: dout  = 8'b10100101; //  501 : 165 - 0xa5
      12'h1F6: dout  = 8'b10100101; //  502 : 165 - 0xa5
      12'h1F7: dout  = 8'b10100101; //  503 : 165 - 0xa5
      12'h1F8: dout  = 8'b00000000; //  504 :   0 - 0x0 -- Sprite 0x3f
      12'h1F9: dout  = 8'b00000000; //  505 :   0 - 0x0
      12'h1FA: dout  = 8'b00000000; //  506 :   0 - 0x0
      12'h1FB: dout  = 8'b11000110; //  507 : 198 - 0xc6
      12'h1FC: dout  = 8'b00101001; //  508 :  41 - 0x29
      12'h1FD: dout  = 8'b00101001; //  509 :  41 - 0x29
      12'h1FE: dout  = 8'b00101001; //  510 :  41 - 0x29
      12'h1FF: dout  = 8'b00101001; //  511 :  41 - 0x29
      12'h200: dout  = 8'b10100101; //  512 : 165 - 0xa5 -- Sprite 0x40
      12'h201: dout  = 8'b10011000; //  513 : 152 - 0x98
      12'h202: dout  = 8'b00000000; //  514 :   0 - 0x0
      12'h203: dout  = 8'b00000000; //  515 :   0 - 0x0
      12'h204: dout  = 8'b00000000; //  516 :   0 - 0x0
      12'h205: dout  = 8'b00000000; //  517 :   0 - 0x0
      12'h206: dout  = 8'b00000000; //  518 :   0 - 0x0
      12'h207: dout  = 8'b00000000; //  519 :   0 - 0x0
      12'h208: dout  = 8'b00101001; //  520 :  41 - 0x29 -- Sprite 0x41
      12'h209: dout  = 8'b11000110; //  521 : 198 - 0xc6
      12'h20A: dout  = 8'b00000000; //  522 :   0 - 0x0
      12'h20B: dout  = 8'b00000000; //  523 :   0 - 0x0
      12'h20C: dout  = 8'b00000000; //  524 :   0 - 0x0
      12'h20D: dout  = 8'b00000000; //  525 :   0 - 0x0
      12'h20E: dout  = 8'b00000000; //  526 :   0 - 0x0
      12'h20F: dout  = 8'b00000000; //  527 :   0 - 0x0
      12'h210: dout  = 8'b00000000; //  528 :   0 - 0x0 -- Sprite 0x42
      12'h211: dout  = 8'b00000000; //  529 :   0 - 0x0
      12'h212: dout  = 8'b00000000; //  530 :   0 - 0x0
      12'h213: dout  = 8'b10011100; //  531 : 156 - 0x9c
      12'h214: dout  = 8'b10100001; //  532 : 161 - 0xa1
      12'h215: dout  = 8'b10100001; //  533 : 161 - 0xa1
      12'h216: dout  = 8'b10111101; //  534 : 189 - 0xbd
      12'h217: dout  = 8'b10100101; //  535 : 165 - 0xa5
      12'h218: dout  = 8'b10100101; //  536 : 165 - 0xa5 -- Sprite 0x43
      12'h219: dout  = 8'b10011000; //  537 : 152 - 0x98
      12'h21A: dout  = 8'b00000000; //  538 :   0 - 0x0
      12'h21B: dout  = 8'b00000000; //  539 :   0 - 0x0
      12'h21C: dout  = 8'b00000000; //  540 :   0 - 0x0
      12'h21D: dout  = 8'b00000000; //  541 :   0 - 0x0
      12'h21E: dout  = 8'b00000000; //  542 :   0 - 0x0
      12'h21F: dout  = 8'b00000000; //  543 :   0 - 0x0
      12'h220: dout  = 8'b00000000; //  544 :   0 - 0x0 -- Sprite 0x44
      12'h221: dout  = 8'b00000000; //  545 :   0 - 0x0
      12'h222: dout  = 8'b00000000; //  546 :   0 - 0x0
      12'h223: dout  = 8'b01100010; //  547 :  98 - 0x62
      12'h224: dout  = 8'b10010101; //  548 : 149 - 0x95
      12'h225: dout  = 8'b00010101; //  549 :  21 - 0x15
      12'h226: dout  = 8'b00100101; //  550 :  37 - 0x25
      12'h227: dout  = 8'b01000101; //  551 :  69 - 0x45
      12'h228: dout  = 8'b00000000; //  552 :   0 - 0x0 -- Sprite 0x45
      12'h229: dout  = 8'b00000000; //  553 :   0 - 0x0
      12'h22A: dout  = 8'b00000000; //  554 :   0 - 0x0
      12'h22B: dout  = 8'b00100010; //  555 :  34 - 0x22
      12'h22C: dout  = 8'b01010101; //  556 :  85 - 0x55
      12'h22D: dout  = 8'b01010101; //  557 :  85 - 0x55
      12'h22E: dout  = 8'b01010101; //  558 :  85 - 0x55
      12'h22F: dout  = 8'b01010101; //  559 :  85 - 0x55
      12'h230: dout  = 8'b10000101; //  560 : 133 - 0x85 -- Sprite 0x46
      12'h231: dout  = 8'b11110010; //  561 : 242 - 0xf2
      12'h232: dout  = 8'b00000000; //  562 :   0 - 0x0
      12'h233: dout  = 8'b00000000; //  563 :   0 - 0x0
      12'h234: dout  = 8'b00000000; //  564 :   0 - 0x0
      12'h235: dout  = 8'b00000000; //  565 :   0 - 0x0
      12'h236: dout  = 8'b00000000; //  566 :   0 - 0x0
      12'h237: dout  = 8'b00000000; //  567 :   0 - 0x0
      12'h238: dout  = 8'b01010101; //  568 :  85 - 0x55 -- Sprite 0x47
      12'h239: dout  = 8'b00100010; //  569 :  34 - 0x22
      12'h23A: dout  = 8'b00000000; //  570 :   0 - 0x0
      12'h23B: dout  = 8'b00000000; //  571 :   0 - 0x0
      12'h23C: dout  = 8'b00000000; //  572 :   0 - 0x0
      12'h23D: dout  = 8'b00000000; //  573 :   0 - 0x0
      12'h23E: dout  = 8'b00000000; //  574 :   0 - 0x0
      12'h23F: dout  = 8'b00000000; //  575 :   0 - 0x0
      12'h240: dout  = 8'b00000000; //  576 :   0 - 0x0 -- Sprite 0x48
      12'h241: dout  = 8'b00000000; //  577 :   0 - 0x0
      12'h242: dout  = 8'b00000000; //  578 :   0 - 0x0
      12'h243: dout  = 8'b01100010; //  579 :  98 - 0x62
      12'h244: dout  = 8'b10010101; //  580 : 149 - 0x95
      12'h245: dout  = 8'b00010101; //  581 :  21 - 0x15
      12'h246: dout  = 8'b01100101; //  582 : 101 - 0x65
      12'h247: dout  = 8'b00010101; //  583 :  21 - 0x15
      12'h248: dout  = 8'b10010101; //  584 : 149 - 0x95 -- Sprite 0x49
      12'h249: dout  = 8'b01100010; //  585 :  98 - 0x62
      12'h24A: dout  = 8'b00000000; //  586 :   0 - 0x0
      12'h24B: dout  = 8'b00000000; //  587 :   0 - 0x0
      12'h24C: dout  = 8'b00000000; //  588 :   0 - 0x0
      12'h24D: dout  = 8'b00000000; //  589 :   0 - 0x0
      12'h24E: dout  = 8'b00000000; //  590 :   0 - 0x0
      12'h24F: dout  = 8'b00000000; //  591 :   0 - 0x0
      12'h250: dout  = 8'b00000000; //  592 :   0 - 0x0 -- Sprite 0x4a
      12'h251: dout  = 8'b00000000; //  593 :   0 - 0x0
      12'h252: dout  = 8'b00000000; //  594 :   0 - 0x0
      12'h253: dout  = 8'b11100010; //  595 : 226 - 0xe2
      12'h254: dout  = 8'b10000101; //  596 : 133 - 0x85
      12'h255: dout  = 8'b10000101; //  597 : 133 - 0x85
      12'h256: dout  = 8'b11100101; //  598 : 229 - 0xe5
      12'h257: dout  = 8'b00010101; //  599 :  21 - 0x15
      12'h258: dout  = 8'b00010101; //  600 :  21 - 0x15 -- Sprite 0x4b
      12'h259: dout  = 8'b11100010; //  601 : 226 - 0xe2
      12'h25A: dout  = 8'b00000000; //  602 :   0 - 0x0
      12'h25B: dout  = 8'b00000000; //  603 :   0 - 0x0
      12'h25C: dout  = 8'b00000000; //  604 :   0 - 0x0
      12'h25D: dout  = 8'b00000000; //  605 :   0 - 0x0
      12'h25E: dout  = 8'b00000000; //  606 :   0 - 0x0
      12'h25F: dout  = 8'b00000000; //  607 :   0 - 0x0
      12'h260: dout  = 8'b00000000; //  608 :   0 - 0x0 -- Sprite 0x4c
      12'h261: dout  = 8'b00000000; //  609 :   0 - 0x0
      12'h262: dout  = 8'b00000000; //  610 :   0 - 0x0
      12'h263: dout  = 8'b00000000; //  611 :   0 - 0x0
      12'h264: dout  = 8'b00000000; //  612 :   0 - 0x0
      12'h265: dout  = 8'b00000000; //  613 :   0 - 0x0
      12'h266: dout  = 8'b00000000; //  614 :   0 - 0x0
      12'h267: dout  = 8'b00000000; //  615 :   0 - 0x0
      12'h268: dout  = 8'b00000000; //  616 :   0 - 0x0 -- Sprite 0x4d
      12'h269: dout  = 8'b00000000; //  617 :   0 - 0x0
      12'h26A: dout  = 8'b00000000; //  618 :   0 - 0x0
      12'h26B: dout  = 8'b00000000; //  619 :   0 - 0x0
      12'h26C: dout  = 8'b00000000; //  620 :   0 - 0x0
      12'h26D: dout  = 8'b00000000; //  621 :   0 - 0x0
      12'h26E: dout  = 8'b00000000; //  622 :   0 - 0x0
      12'h26F: dout  = 8'b00000000; //  623 :   0 - 0x0
      12'h270: dout  = 8'b00000000; //  624 :   0 - 0x0 -- Sprite 0x4e
      12'h271: dout  = 8'b00000000; //  625 :   0 - 0x0
      12'h272: dout  = 8'b00000000; //  626 :   0 - 0x0
      12'h273: dout  = 8'b00000000; //  627 :   0 - 0x0
      12'h274: dout  = 8'b00000000; //  628 :   0 - 0x0
      12'h275: dout  = 8'b00000000; //  629 :   0 - 0x0
      12'h276: dout  = 8'b00000000; //  630 :   0 - 0x0
      12'h277: dout  = 8'b00000000; //  631 :   0 - 0x0
      12'h278: dout  = 8'b00000000; //  632 :   0 - 0x0 -- Sprite 0x4f
      12'h279: dout  = 8'b00000000; //  633 :   0 - 0x0
      12'h27A: dout  = 8'b00000000; //  634 :   0 - 0x0
      12'h27B: dout  = 8'b00000000; //  635 :   0 - 0x0
      12'h27C: dout  = 8'b00000000; //  636 :   0 - 0x0
      12'h27D: dout  = 8'b00000000; //  637 :   0 - 0x0
      12'h27E: dout  = 8'b00000000; //  638 :   0 - 0x0
      12'h27F: dout  = 8'b00000000; //  639 :   0 - 0x0
      12'h280: dout  = 8'b00000000; //  640 :   0 - 0x0 -- Sprite 0x50
      12'h281: dout  = 8'b00000000; //  641 :   0 - 0x0
      12'h282: dout  = 8'b00000000; //  642 :   0 - 0x0
      12'h283: dout  = 8'b00000000; //  643 :   0 - 0x0
      12'h284: dout  = 8'b00000000; //  644 :   0 - 0x0
      12'h285: dout  = 8'b00000000; //  645 :   0 - 0x0
      12'h286: dout  = 8'b00000000; //  646 :   0 - 0x0
      12'h287: dout  = 8'b00000000; //  647 :   0 - 0x0
      12'h288: dout  = 8'b00000000; //  648 :   0 - 0x0 -- Sprite 0x51
      12'h289: dout  = 8'b00000000; //  649 :   0 - 0x0
      12'h28A: dout  = 8'b00000000; //  650 :   0 - 0x0
      12'h28B: dout  = 8'b00000000; //  651 :   0 - 0x0
      12'h28C: dout  = 8'b00000000; //  652 :   0 - 0x0
      12'h28D: dout  = 8'b00000000; //  653 :   0 - 0x0
      12'h28E: dout  = 8'b00000000; //  654 :   0 - 0x0
      12'h28F: dout  = 8'b00000000; //  655 :   0 - 0x0
      12'h290: dout  = 8'b00000000; //  656 :   0 - 0x0 -- Sprite 0x52
      12'h291: dout  = 8'b00000000; //  657 :   0 - 0x0
      12'h292: dout  = 8'b00000000; //  658 :   0 - 0x0
      12'h293: dout  = 8'b00000000; //  659 :   0 - 0x0
      12'h294: dout  = 8'b00000000; //  660 :   0 - 0x0
      12'h295: dout  = 8'b00000000; //  661 :   0 - 0x0
      12'h296: dout  = 8'b00000000; //  662 :   0 - 0x0
      12'h297: dout  = 8'b00000000; //  663 :   0 - 0x0
      12'h298: dout  = 8'b00000000; //  664 :   0 - 0x0 -- Sprite 0x53
      12'h299: dout  = 8'b00000000; //  665 :   0 - 0x0
      12'h29A: dout  = 8'b00000000; //  666 :   0 - 0x0
      12'h29B: dout  = 8'b00000000; //  667 :   0 - 0x0
      12'h29C: dout  = 8'b00000000; //  668 :   0 - 0x0
      12'h29D: dout  = 8'b00000000; //  669 :   0 - 0x0
      12'h29E: dout  = 8'b00000000; //  670 :   0 - 0x0
      12'h29F: dout  = 8'b00000000; //  671 :   0 - 0x0
      12'h2A0: dout  = 8'b00000000; //  672 :   0 - 0x0 -- Sprite 0x54
      12'h2A1: dout  = 8'b00000000; //  673 :   0 - 0x0
      12'h2A2: dout  = 8'b00000000; //  674 :   0 - 0x0
      12'h2A3: dout  = 8'b00000000; //  675 :   0 - 0x0
      12'h2A4: dout  = 8'b00000000; //  676 :   0 - 0x0
      12'h2A5: dout  = 8'b00000000; //  677 :   0 - 0x0
      12'h2A6: dout  = 8'b00000000; //  678 :   0 - 0x0
      12'h2A7: dout  = 8'b00000000; //  679 :   0 - 0x0
      12'h2A8: dout  = 8'b00000000; //  680 :   0 - 0x0 -- Sprite 0x55
      12'h2A9: dout  = 8'b00000000; //  681 :   0 - 0x0
      12'h2AA: dout  = 8'b00000000; //  682 :   0 - 0x0
      12'h2AB: dout  = 8'b00000000; //  683 :   0 - 0x0
      12'h2AC: dout  = 8'b00000000; //  684 :   0 - 0x0
      12'h2AD: dout  = 8'b00000000; //  685 :   0 - 0x0
      12'h2AE: dout  = 8'b00000000; //  686 :   0 - 0x0
      12'h2AF: dout  = 8'b00000000; //  687 :   0 - 0x0
      12'h2B0: dout  = 8'b00000000; //  688 :   0 - 0x0 -- Sprite 0x56
      12'h2B1: dout  = 8'b00000000; //  689 :   0 - 0x0
      12'h2B2: dout  = 8'b00000000; //  690 :   0 - 0x0
      12'h2B3: dout  = 8'b00000000; //  691 :   0 - 0x0
      12'h2B4: dout  = 8'b00000000; //  692 :   0 - 0x0
      12'h2B5: dout  = 8'b00000000; //  693 :   0 - 0x0
      12'h2B6: dout  = 8'b00000000; //  694 :   0 - 0x0
      12'h2B7: dout  = 8'b00000000; //  695 :   0 - 0x0
      12'h2B8: dout  = 8'b00000000; //  696 :   0 - 0x0 -- Sprite 0x57
      12'h2B9: dout  = 8'b00000000; //  697 :   0 - 0x0
      12'h2BA: dout  = 8'b00000000; //  698 :   0 - 0x0
      12'h2BB: dout  = 8'b00000000; //  699 :   0 - 0x0
      12'h2BC: dout  = 8'b00000000; //  700 :   0 - 0x0
      12'h2BD: dout  = 8'b00000000; //  701 :   0 - 0x0
      12'h2BE: dout  = 8'b00000000; //  702 :   0 - 0x0
      12'h2BF: dout  = 8'b00000100; //  703 :   4 - 0x4
      12'h2C0: dout  = 8'b00000110; //  704 :   6 - 0x6 -- Sprite 0x58
      12'h2C1: dout  = 8'b00000110; //  705 :   6 - 0x6
      12'h2C2: dout  = 8'b00000111; //  706 :   7 - 0x7
      12'h2C3: dout  = 8'b00000111; //  707 :   7 - 0x7
      12'h2C4: dout  = 8'b00000111; //  708 :   7 - 0x7
      12'h2C5: dout  = 8'b00000111; //  709 :   7 - 0x7
      12'h2C6: dout  = 8'b00000000; //  710 :   0 - 0x0
      12'h2C7: dout  = 8'b00000000; //  711 :   0 - 0x0
      12'h2C8: dout  = 8'b00000000; //  712 :   0 - 0x0 -- Sprite 0x59
      12'h2C9: dout  = 8'b00000000; //  713 :   0 - 0x0
      12'h2CA: dout  = 8'b00000000; //  714 :   0 - 0x0
      12'h2CB: dout  = 8'b00000000; //  715 :   0 - 0x0
      12'h2CC: dout  = 8'b00000000; //  716 :   0 - 0x0
      12'h2CD: dout  = 8'b00000000; //  717 :   0 - 0x0
      12'h2CE: dout  = 8'b00000000; //  718 :   0 - 0x0
      12'h2CF: dout  = 8'b00010000; //  719 :  16 - 0x10
      12'h2D0: dout  = 8'b00011100; //  720 :  28 - 0x1c -- Sprite 0x5a
      12'h2D1: dout  = 8'b00011110; //  721 :  30 - 0x1e
      12'h2D2: dout  = 8'b00011111; //  722 :  31 - 0x1f
      12'h2D3: dout  = 8'b00011111; //  723 :  31 - 0x1f
      12'h2D4: dout  = 8'b00011111; //  724 :  31 - 0x1f
      12'h2D5: dout  = 8'b00011111; //  725 :  31 - 0x1f
      12'h2D6: dout  = 8'b00000000; //  726 :   0 - 0x0
      12'h2D7: dout  = 8'b00000000; //  727 :   0 - 0x0
      12'h2D8: dout  = 8'b00000000; //  728 :   0 - 0x0 -- Sprite 0x5b
      12'h2D9: dout  = 8'b00000000; //  729 :   0 - 0x0
      12'h2DA: dout  = 8'b00000000; //  730 :   0 - 0x0
      12'h2DB: dout  = 8'b00000000; //  731 :   0 - 0x0
      12'h2DC: dout  = 8'b00000000; //  732 :   0 - 0x0
      12'h2DD: dout  = 8'b00000000; //  733 :   0 - 0x0
      12'h2DE: dout  = 8'b00000000; //  734 :   0 - 0x0
      12'h2DF: dout  = 8'b11000000; //  735 : 192 - 0xc0
      12'h2E0: dout  = 8'b11110000; //  736 : 240 - 0xf0 -- Sprite 0x5c
      12'h2E1: dout  = 8'b11111100; //  737 : 252 - 0xfc
      12'h2E2: dout  = 8'b11111111; //  738 : 255 - 0xff
      12'h2E3: dout  = 8'b11111111; //  739 : 255 - 0xff
      12'h2E4: dout  = 8'b11111111; //  740 : 255 - 0xff
      12'h2E5: dout  = 8'b11111111; //  741 : 255 - 0xff
      12'h2E6: dout  = 8'b00000000; //  742 :   0 - 0x0
      12'h2E7: dout  = 8'b00000000; //  743 :   0 - 0x0
      12'h2E8: dout  = 8'b00000000; //  744 :   0 - 0x0 -- Sprite 0x5d
      12'h2E9: dout  = 8'b00000000; //  745 :   0 - 0x0
      12'h2EA: dout  = 8'b00000001; //  746 :   1 - 0x1
      12'h2EB: dout  = 8'b00000011; //  747 :   3 - 0x3
      12'h2EC: dout  = 8'b00001111; //  748 :  15 - 0xf
      12'h2ED: dout  = 8'b00001111; //  749 :  15 - 0xf
      12'h2EE: dout  = 8'b00000000; //  750 :   0 - 0x0
      12'h2EF: dout  = 8'b00000000; //  751 :   0 - 0x0
      12'h2F0: dout  = 8'b11111000; //  752 : 248 - 0xf8 -- Sprite 0x5e
      12'h2F1: dout  = 8'b11110000; //  753 : 240 - 0xf0
      12'h2F2: dout  = 8'b11100000; //  754 : 224 - 0xe0
      12'h2F3: dout  = 8'b11110000; //  755 : 240 - 0xf0
      12'h2F4: dout  = 8'b11100000; //  756 : 224 - 0xe0
      12'h2F5: dout  = 8'b11000000; //  757 : 192 - 0xc0
      12'h2F6: dout  = 8'b00000000; //  758 :   0 - 0x0
      12'h2F7: dout  = 8'b00000000; //  759 :   0 - 0x0
      12'h2F8: dout  = 8'b00000000; //  760 :   0 - 0x0 -- Sprite 0x5f
      12'h2F9: dout  = 8'b00000000; //  761 :   0 - 0x0
      12'h2FA: dout  = 8'b00000000; //  762 :   0 - 0x0
      12'h2FB: dout  = 8'b00000000; //  763 :   0 - 0x0
      12'h2FC: dout  = 8'b00000000; //  764 :   0 - 0x0
      12'h2FD: dout  = 8'b00000000; //  765 :   0 - 0x0
      12'h2FE: dout  = 8'b00000000; //  766 :   0 - 0x0
      12'h2FF: dout  = 8'b00000000; //  767 :   0 - 0x0
      12'h300: dout  = 8'b00000000; //  768 :   0 - 0x0 -- Sprite 0x60
      12'h301: dout  = 8'b00000011; //  769 :   3 - 0x3
      12'h302: dout  = 8'b00001111; //  770 :  15 - 0xf
      12'h303: dout  = 8'b00011111; //  771 :  31 - 0x1f
      12'h304: dout  = 8'b00111111; //  772 :  63 - 0x3f
      12'h305: dout  = 8'b00111111; //  773 :  63 - 0x3f
      12'h306: dout  = 8'b00111001; //  774 :  57 - 0x39
      12'h307: dout  = 8'b01111011; //  775 : 123 - 0x7b
      12'h308: dout  = 8'b00000000; //  776 :   0 - 0x0 -- Sprite 0x61
      12'h309: dout  = 8'b11000000; //  777 : 192 - 0xc0
      12'h30A: dout  = 8'b11110000; //  778 : 240 - 0xf0
      12'h30B: dout  = 8'b11111000; //  779 : 248 - 0xf8
      12'h30C: dout  = 8'b11111100; //  780 : 252 - 0xfc
      12'h30D: dout  = 8'b11111100; //  781 : 252 - 0xfc
      12'h30E: dout  = 8'b11100100; //  782 : 228 - 0xe4
      12'h30F: dout  = 8'b11101110; //  783 : 238 - 0xee
      12'h310: dout  = 8'b11111110; //  784 : 254 - 0xfe -- Sprite 0x62
      12'h311: dout  = 8'b11111110; //  785 : 254 - 0xfe
      12'h312: dout  = 8'b11111110; //  786 : 254 - 0xfe
      12'h313: dout  = 8'b11111110; //  787 : 254 - 0xfe
      12'h314: dout  = 8'b11111110; //  788 : 254 - 0xfe
      12'h315: dout  = 8'b01100110; //  789 : 102 - 0x66
      12'h316: dout  = 8'b01000010; //  790 :  66 - 0x42
      12'h317: dout  = 8'b00000000; //  791 :   0 - 0x0
      12'h318: dout  = 8'b11111110; //  792 : 254 - 0xfe -- Sprite 0x63
      12'h319: dout  = 8'b11111110; //  793 : 254 - 0xfe
      12'h31A: dout  = 8'b11111110; //  794 : 254 - 0xfe
      12'h31B: dout  = 8'b11111110; //  795 : 254 - 0xfe
      12'h31C: dout  = 8'b11111110; //  796 : 254 - 0xfe
      12'h31D: dout  = 8'b11011110; //  797 : 222 - 0xde
      12'h31E: dout  = 8'b10001100; //  798 : 140 - 0x8c
      12'h31F: dout  = 8'b00000000; //  799 :   0 - 0x0
      12'h320: dout  = 8'b00000000; //  800 :   0 - 0x0 -- Sprite 0x64
      12'h321: dout  = 8'b00000000; //  801 :   0 - 0x0
      12'h322: dout  = 8'b00000000; //  802 :   0 - 0x0
      12'h323: dout  = 8'b00000000; //  803 :   0 - 0x0
      12'h324: dout  = 8'b00000000; //  804 :   0 - 0x0
      12'h325: dout  = 8'b00000000; //  805 :   0 - 0x0
      12'h326: dout  = 8'b00000000; //  806 :   0 - 0x0
      12'h327: dout  = 8'b00000000; //  807 :   0 - 0x0
      12'h328: dout  = 8'b00000000; //  808 :   0 - 0x0 -- Sprite 0x65
      12'h329: dout  = 8'b00000000; //  809 :   0 - 0x0
      12'h32A: dout  = 8'b00000000; //  810 :   0 - 0x0
      12'h32B: dout  = 8'b00000000; //  811 :   0 - 0x0
      12'h32C: dout  = 8'b01101100; //  812 : 108 - 0x6c
      12'h32D: dout  = 8'b11111110; //  813 : 254 - 0xfe
      12'h32E: dout  = 8'b11111110; //  814 : 254 - 0xfe
      12'h32F: dout  = 8'b11111100; //  815 : 252 - 0xfc
      12'h330: dout  = 8'b00000000; //  816 :   0 - 0x0 -- Sprite 0x66
      12'h331: dout  = 8'b00000000; //  817 :   0 - 0x0
      12'h332: dout  = 8'b00000000; //  818 :   0 - 0x0
      12'h333: dout  = 8'b00000000; //  819 :   0 - 0x0
      12'h334: dout  = 8'b00000000; //  820 :   0 - 0x0
      12'h335: dout  = 8'b00000000; //  821 :   0 - 0x0
      12'h336: dout  = 8'b00000000; //  822 :   0 - 0x0
      12'h337: dout  = 8'b00000000; //  823 :   0 - 0x0
      12'h338: dout  = 8'b00000000; //  824 :   0 - 0x0 -- Sprite 0x67
      12'h339: dout  = 8'b00000000; //  825 :   0 - 0x0
      12'h33A: dout  = 8'b00000000; //  826 :   0 - 0x0
      12'h33B: dout  = 8'b00000000; //  827 :   0 - 0x0
      12'h33C: dout  = 8'b00000000; //  828 :   0 - 0x0
      12'h33D: dout  = 8'b00000000; //  829 :   0 - 0x0
      12'h33E: dout  = 8'b00000000; //  830 :   0 - 0x0
      12'h33F: dout  = 8'b00000000; //  831 :   0 - 0x0
      12'h340: dout  = 8'b00000000; //  832 :   0 - 0x0 -- Sprite 0x68
      12'h341: dout  = 8'b00000000; //  833 :   0 - 0x0
      12'h342: dout  = 8'b00000000; //  834 :   0 - 0x0
      12'h343: dout  = 8'b00000000; //  835 :   0 - 0x0
      12'h344: dout  = 8'b00000000; //  836 :   0 - 0x0
      12'h345: dout  = 8'b00000000; //  837 :   0 - 0x0
      12'h346: dout  = 8'b00000000; //  838 :   0 - 0x0
      12'h347: dout  = 8'b00000000; //  839 :   0 - 0x0
      12'h348: dout  = 8'b00000000; //  840 :   0 - 0x0 -- Sprite 0x69
      12'h349: dout  = 8'b00000000; //  841 :   0 - 0x0
      12'h34A: dout  = 8'b00000000; //  842 :   0 - 0x0
      12'h34B: dout  = 8'b00000000; //  843 :   0 - 0x0
      12'h34C: dout  = 8'b00000000; //  844 :   0 - 0x0
      12'h34D: dout  = 8'b00000000; //  845 :   0 - 0x0
      12'h34E: dout  = 8'b00000000; //  846 :   0 - 0x0
      12'h34F: dout  = 8'b00000000; //  847 :   0 - 0x0
      12'h350: dout  = 8'b00000000; //  848 :   0 - 0x0 -- Sprite 0x6a
      12'h351: dout  = 8'b00011111; //  849 :  31 - 0x1f
      12'h352: dout  = 8'b01111111; //  850 : 127 - 0x7f
      12'h353: dout  = 8'b00111111; //  851 :  63 - 0x3f
      12'h354: dout  = 8'b00001111; //  852 :  15 - 0xf
      12'h355: dout  = 8'b00000111; //  853 :   7 - 0x7
      12'h356: dout  = 8'b00000000; //  854 :   0 - 0x0
      12'h357: dout  = 8'b00000000; //  855 :   0 - 0x0
      12'h358: dout  = 8'b00000000; //  856 :   0 - 0x0 -- Sprite 0x6b
      12'h359: dout  = 8'b00000000; //  857 :   0 - 0x0
      12'h35A: dout  = 8'b11000000; //  858 : 192 - 0xc0
      12'h35B: dout  = 8'b11110000; //  859 : 240 - 0xf0
      12'h35C: dout  = 8'b11111000; //  860 : 248 - 0xf8
      12'h35D: dout  = 8'b11111000; //  861 : 248 - 0xf8
      12'h35E: dout  = 8'b11100000; //  862 : 224 - 0xe0
      12'h35F: dout  = 8'b00000000; //  863 :   0 - 0x0
      12'h360: dout  = 8'b00000000; //  864 :   0 - 0x0 -- Sprite 0x6c
      12'h361: dout  = 8'b00000000; //  865 :   0 - 0x0
      12'h362: dout  = 8'b00000000; //  866 :   0 - 0x0
      12'h363: dout  = 8'b00000000; //  867 :   0 - 0x0
      12'h364: dout  = 8'b00000000; //  868 :   0 - 0x0
      12'h365: dout  = 8'b00000000; //  869 :   0 - 0x0
      12'h366: dout  = 8'b00000000; //  870 :   0 - 0x0
      12'h367: dout  = 8'b00000000; //  871 :   0 - 0x0
      12'h368: dout  = 8'b00000000; //  872 :   0 - 0x0 -- Sprite 0x6d
      12'h369: dout  = 8'b00000000; //  873 :   0 - 0x0
      12'h36A: dout  = 8'b00000000; //  874 :   0 - 0x0
      12'h36B: dout  = 8'b00000000; //  875 :   0 - 0x0
      12'h36C: dout  = 8'b00000000; //  876 :   0 - 0x0
      12'h36D: dout  = 8'b00000000; //  877 :   0 - 0x0
      12'h36E: dout  = 8'b00000000; //  878 :   0 - 0x0
      12'h36F: dout  = 8'b00000000; //  879 :   0 - 0x0
      12'h370: dout  = 8'b00000000; //  880 :   0 - 0x0 -- Sprite 0x6e
      12'h371: dout  = 8'b00000000; //  881 :   0 - 0x0
      12'h372: dout  = 8'b00000000; //  882 :   0 - 0x0
      12'h373: dout  = 8'b00000000; //  883 :   0 - 0x0
      12'h374: dout  = 8'b00000000; //  884 :   0 - 0x0
      12'h375: dout  = 8'b00000000; //  885 :   0 - 0x0
      12'h376: dout  = 8'b00000000; //  886 :   0 - 0x0
      12'h377: dout  = 8'b00000000; //  887 :   0 - 0x0
      12'h378: dout  = 8'b00000000; //  888 :   0 - 0x0 -- Sprite 0x6f
      12'h379: dout  = 8'b00000000; //  889 :   0 - 0x0
      12'h37A: dout  = 8'b00000000; //  890 :   0 - 0x0
      12'h37B: dout  = 8'b00000000; //  891 :   0 - 0x0
      12'h37C: dout  = 8'b00000000; //  892 :   0 - 0x0
      12'h37D: dout  = 8'b00000000; //  893 :   0 - 0x0
      12'h37E: dout  = 8'b00000000; //  894 :   0 - 0x0
      12'h37F: dout  = 8'b00000000; //  895 :   0 - 0x0
      12'h380: dout  = 8'b11111111; //  896 : 255 - 0xff -- Sprite 0x70
      12'h381: dout  = 8'b11111111; //  897 : 255 - 0xff
      12'h382: dout  = 8'b11111111; //  898 : 255 - 0xff
      12'h383: dout  = 8'b11111111; //  899 : 255 - 0xff
      12'h384: dout  = 8'b11111111; //  900 : 255 - 0xff
      12'h385: dout  = 8'b11111111; //  901 : 255 - 0xff
      12'h386: dout  = 8'b11111111; //  902 : 255 - 0xff
      12'h387: dout  = 8'b11111111; //  903 : 255 - 0xff
      12'h388: dout  = 8'b11111111; //  904 : 255 - 0xff -- Sprite 0x71
      12'h389: dout  = 8'b11111111; //  905 : 255 - 0xff
      12'h38A: dout  = 8'b11111111; //  906 : 255 - 0xff
      12'h38B: dout  = 8'b11111111; //  907 : 255 - 0xff
      12'h38C: dout  = 8'b11111111; //  908 : 255 - 0xff
      12'h38D: dout  = 8'b11111111; //  909 : 255 - 0xff
      12'h38E: dout  = 8'b11111111; //  910 : 255 - 0xff
      12'h38F: dout  = 8'b11111111; //  911 : 255 - 0xff
      12'h390: dout  = 8'b11111111; //  912 : 255 - 0xff -- Sprite 0x72
      12'h391: dout  = 8'b11111111; //  913 : 255 - 0xff
      12'h392: dout  = 8'b11111111; //  914 : 255 - 0xff
      12'h393: dout  = 8'b11111111; //  915 : 255 - 0xff
      12'h394: dout  = 8'b11111111; //  916 : 255 - 0xff
      12'h395: dout  = 8'b11111111; //  917 : 255 - 0xff
      12'h396: dout  = 8'b11111111; //  918 : 255 - 0xff
      12'h397: dout  = 8'b11111111; //  919 : 255 - 0xff
      12'h398: dout  = 8'b11111111; //  920 : 255 - 0xff -- Sprite 0x73
      12'h399: dout  = 8'b11111111; //  921 : 255 - 0xff
      12'h39A: dout  = 8'b11111111; //  922 : 255 - 0xff
      12'h39B: dout  = 8'b11111111; //  923 : 255 - 0xff
      12'h39C: dout  = 8'b11111111; //  924 : 255 - 0xff
      12'h39D: dout  = 8'b11111111; //  925 : 255 - 0xff
      12'h39E: dout  = 8'b11111111; //  926 : 255 - 0xff
      12'h39F: dout  = 8'b11111111; //  927 : 255 - 0xff
      12'h3A0: dout  = 8'b11111111; //  928 : 255 - 0xff -- Sprite 0x74
      12'h3A1: dout  = 8'b11111111; //  929 : 255 - 0xff
      12'h3A2: dout  = 8'b11111111; //  930 : 255 - 0xff
      12'h3A3: dout  = 8'b11111111; //  931 : 255 - 0xff
      12'h3A4: dout  = 8'b11111111; //  932 : 255 - 0xff
      12'h3A5: dout  = 8'b11111111; //  933 : 255 - 0xff
      12'h3A6: dout  = 8'b11111111; //  934 : 255 - 0xff
      12'h3A7: dout  = 8'b11111111; //  935 : 255 - 0xff
      12'h3A8: dout  = 8'b11111111; //  936 : 255 - 0xff -- Sprite 0x75
      12'h3A9: dout  = 8'b11111111; //  937 : 255 - 0xff
      12'h3AA: dout  = 8'b11111111; //  938 : 255 - 0xff
      12'h3AB: dout  = 8'b11111111; //  939 : 255 - 0xff
      12'h3AC: dout  = 8'b11111111; //  940 : 255 - 0xff
      12'h3AD: dout  = 8'b11111111; //  941 : 255 - 0xff
      12'h3AE: dout  = 8'b11111111; //  942 : 255 - 0xff
      12'h3AF: dout  = 8'b11111111; //  943 : 255 - 0xff
      12'h3B0: dout  = 8'b11111111; //  944 : 255 - 0xff -- Sprite 0x76
      12'h3B1: dout  = 8'b11111111; //  945 : 255 - 0xff
      12'h3B2: dout  = 8'b11111111; //  946 : 255 - 0xff
      12'h3B3: dout  = 8'b11111111; //  947 : 255 - 0xff
      12'h3B4: dout  = 8'b11111111; //  948 : 255 - 0xff
      12'h3B5: dout  = 8'b11111111; //  949 : 255 - 0xff
      12'h3B6: dout  = 8'b11111111; //  950 : 255 - 0xff
      12'h3B7: dout  = 8'b11111111; //  951 : 255 - 0xff
      12'h3B8: dout  = 8'b11111111; //  952 : 255 - 0xff -- Sprite 0x77
      12'h3B9: dout  = 8'b11111111; //  953 : 255 - 0xff
      12'h3BA: dout  = 8'b11111111; //  954 : 255 - 0xff
      12'h3BB: dout  = 8'b11111111; //  955 : 255 - 0xff
      12'h3BC: dout  = 8'b11111111; //  956 : 255 - 0xff
      12'h3BD: dout  = 8'b11111111; //  957 : 255 - 0xff
      12'h3BE: dout  = 8'b11111111; //  958 : 255 - 0xff
      12'h3BF: dout  = 8'b11111111; //  959 : 255 - 0xff
      12'h3C0: dout  = 8'b11111111; //  960 : 255 - 0xff -- Sprite 0x78
      12'h3C1: dout  = 8'b11111111; //  961 : 255 - 0xff
      12'h3C2: dout  = 8'b11111111; //  962 : 255 - 0xff
      12'h3C3: dout  = 8'b11111111; //  963 : 255 - 0xff
      12'h3C4: dout  = 8'b11111111; //  964 : 255 - 0xff
      12'h3C5: dout  = 8'b11111111; //  965 : 255 - 0xff
      12'h3C6: dout  = 8'b11111111; //  966 : 255 - 0xff
      12'h3C7: dout  = 8'b11111111; //  967 : 255 - 0xff
      12'h3C8: dout  = 8'b11111111; //  968 : 255 - 0xff -- Sprite 0x79
      12'h3C9: dout  = 8'b11111111; //  969 : 255 - 0xff
      12'h3CA: dout  = 8'b11111111; //  970 : 255 - 0xff
      12'h3CB: dout  = 8'b11111111; //  971 : 255 - 0xff
      12'h3CC: dout  = 8'b11111111; //  972 : 255 - 0xff
      12'h3CD: dout  = 8'b11111111; //  973 : 255 - 0xff
      12'h3CE: dout  = 8'b11111111; //  974 : 255 - 0xff
      12'h3CF: dout  = 8'b11111111; //  975 : 255 - 0xff
      12'h3D0: dout  = 8'b11111111; //  976 : 255 - 0xff -- Sprite 0x7a
      12'h3D1: dout  = 8'b11111111; //  977 : 255 - 0xff
      12'h3D2: dout  = 8'b11111111; //  978 : 255 - 0xff
      12'h3D3: dout  = 8'b11111111; //  979 : 255 - 0xff
      12'h3D4: dout  = 8'b11111111; //  980 : 255 - 0xff
      12'h3D5: dout  = 8'b11111111; //  981 : 255 - 0xff
      12'h3D6: dout  = 8'b11111111; //  982 : 255 - 0xff
      12'h3D7: dout  = 8'b11111111; //  983 : 255 - 0xff
      12'h3D8: dout  = 8'b11111111; //  984 : 255 - 0xff -- Sprite 0x7b
      12'h3D9: dout  = 8'b11111111; //  985 : 255 - 0xff
      12'h3DA: dout  = 8'b11111111; //  986 : 255 - 0xff
      12'h3DB: dout  = 8'b11111111; //  987 : 255 - 0xff
      12'h3DC: dout  = 8'b11111111; //  988 : 255 - 0xff
      12'h3DD: dout  = 8'b11111111; //  989 : 255 - 0xff
      12'h3DE: dout  = 8'b11111111; //  990 : 255 - 0xff
      12'h3DF: dout  = 8'b11111111; //  991 : 255 - 0xff
      12'h3E0: dout  = 8'b11111111; //  992 : 255 - 0xff -- Sprite 0x7c
      12'h3E1: dout  = 8'b11111111; //  993 : 255 - 0xff
      12'h3E2: dout  = 8'b11111111; //  994 : 255 - 0xff
      12'h3E3: dout  = 8'b11111111; //  995 : 255 - 0xff
      12'h3E4: dout  = 8'b11111111; //  996 : 255 - 0xff
      12'h3E5: dout  = 8'b11111111; //  997 : 255 - 0xff
      12'h3E6: dout  = 8'b11111111; //  998 : 255 - 0xff
      12'h3E7: dout  = 8'b11111111; //  999 : 255 - 0xff
      12'h3E8: dout  = 8'b11111111; // 1000 : 255 - 0xff -- Sprite 0x7d
      12'h3E9: dout  = 8'b11111111; // 1001 : 255 - 0xff
      12'h3EA: dout  = 8'b11111111; // 1002 : 255 - 0xff
      12'h3EB: dout  = 8'b11111111; // 1003 : 255 - 0xff
      12'h3EC: dout  = 8'b11111111; // 1004 : 255 - 0xff
      12'h3ED: dout  = 8'b11111111; // 1005 : 255 - 0xff
      12'h3EE: dout  = 8'b11111111; // 1006 : 255 - 0xff
      12'h3EF: dout  = 8'b11111111; // 1007 : 255 - 0xff
      12'h3F0: dout  = 8'b11111111; // 1008 : 255 - 0xff -- Sprite 0x7e
      12'h3F1: dout  = 8'b11111111; // 1009 : 255 - 0xff
      12'h3F2: dout  = 8'b11111111; // 1010 : 255 - 0xff
      12'h3F3: dout  = 8'b11111111; // 1011 : 255 - 0xff
      12'h3F4: dout  = 8'b11111111; // 1012 : 255 - 0xff
      12'h3F5: dout  = 8'b11111111; // 1013 : 255 - 0xff
      12'h3F6: dout  = 8'b11111111; // 1014 : 255 - 0xff
      12'h3F7: dout  = 8'b11111111; // 1015 : 255 - 0xff
      12'h3F8: dout  = 8'b11111111; // 1016 : 255 - 0xff -- Sprite 0x7f
      12'h3F9: dout  = 8'b11111111; // 1017 : 255 - 0xff
      12'h3FA: dout  = 8'b11111111; // 1018 : 255 - 0xff
      12'h3FB: dout  = 8'b11111111; // 1019 : 255 - 0xff
      12'h3FC: dout  = 8'b11111111; // 1020 : 255 - 0xff
      12'h3FD: dout  = 8'b11111111; // 1021 : 255 - 0xff
      12'h3FE: dout  = 8'b11111111; // 1022 : 255 - 0xff
      12'h3FF: dout  = 8'b11111111; // 1023 : 255 - 0xff
      12'h400: dout  = 8'b11111111; // 1024 : 255 - 0xff -- Sprite 0x80
      12'h401: dout  = 8'b11111111; // 1025 : 255 - 0xff
      12'h402: dout  = 8'b11111111; // 1026 : 255 - 0xff
      12'h403: dout  = 8'b11111111; // 1027 : 255 - 0xff
      12'h404: dout  = 8'b11111111; // 1028 : 255 - 0xff
      12'h405: dout  = 8'b11111111; // 1029 : 255 - 0xff
      12'h406: dout  = 8'b11111111; // 1030 : 255 - 0xff
      12'h407: dout  = 8'b11111111; // 1031 : 255 - 0xff
      12'h408: dout  = 8'b11111111; // 1032 : 255 - 0xff -- Sprite 0x81
      12'h409: dout  = 8'b11111111; // 1033 : 255 - 0xff
      12'h40A: dout  = 8'b11111111; // 1034 : 255 - 0xff
      12'h40B: dout  = 8'b11111111; // 1035 : 255 - 0xff
      12'h40C: dout  = 8'b11111111; // 1036 : 255 - 0xff
      12'h40D: dout  = 8'b11111111; // 1037 : 255 - 0xff
      12'h40E: dout  = 8'b11111111; // 1038 : 255 - 0xff
      12'h40F: dout  = 8'b11111111; // 1039 : 255 - 0xff
      12'h410: dout  = 8'b11111111; // 1040 : 255 - 0xff -- Sprite 0x82
      12'h411: dout  = 8'b11111111; // 1041 : 255 - 0xff
      12'h412: dout  = 8'b11111111; // 1042 : 255 - 0xff
      12'h413: dout  = 8'b11111111; // 1043 : 255 - 0xff
      12'h414: dout  = 8'b11111111; // 1044 : 255 - 0xff
      12'h415: dout  = 8'b11111111; // 1045 : 255 - 0xff
      12'h416: dout  = 8'b11111111; // 1046 : 255 - 0xff
      12'h417: dout  = 8'b11111111; // 1047 : 255 - 0xff
      12'h418: dout  = 8'b11111111; // 1048 : 255 - 0xff -- Sprite 0x83
      12'h419: dout  = 8'b11111111; // 1049 : 255 - 0xff
      12'h41A: dout  = 8'b11111111; // 1050 : 255 - 0xff
      12'h41B: dout  = 8'b11111111; // 1051 : 255 - 0xff
      12'h41C: dout  = 8'b11111111; // 1052 : 255 - 0xff
      12'h41D: dout  = 8'b11111111; // 1053 : 255 - 0xff
      12'h41E: dout  = 8'b11111111; // 1054 : 255 - 0xff
      12'h41F: dout  = 8'b11111111; // 1055 : 255 - 0xff
      12'h420: dout  = 8'b11111111; // 1056 : 255 - 0xff -- Sprite 0x84
      12'h421: dout  = 8'b11111111; // 1057 : 255 - 0xff
      12'h422: dout  = 8'b11111111; // 1058 : 255 - 0xff
      12'h423: dout  = 8'b11111111; // 1059 : 255 - 0xff
      12'h424: dout  = 8'b11111111; // 1060 : 255 - 0xff
      12'h425: dout  = 8'b11111111; // 1061 : 255 - 0xff
      12'h426: dout  = 8'b11111111; // 1062 : 255 - 0xff
      12'h427: dout  = 8'b11111111; // 1063 : 255 - 0xff
      12'h428: dout  = 8'b11111111; // 1064 : 255 - 0xff -- Sprite 0x85
      12'h429: dout  = 8'b11111111; // 1065 : 255 - 0xff
      12'h42A: dout  = 8'b11111111; // 1066 : 255 - 0xff
      12'h42B: dout  = 8'b11111111; // 1067 : 255 - 0xff
      12'h42C: dout  = 8'b11111111; // 1068 : 255 - 0xff
      12'h42D: dout  = 8'b11111111; // 1069 : 255 - 0xff
      12'h42E: dout  = 8'b11111111; // 1070 : 255 - 0xff
      12'h42F: dout  = 8'b11111111; // 1071 : 255 - 0xff
      12'h430: dout  = 8'b11111111; // 1072 : 255 - 0xff -- Sprite 0x86
      12'h431: dout  = 8'b11111111; // 1073 : 255 - 0xff
      12'h432: dout  = 8'b11111111; // 1074 : 255 - 0xff
      12'h433: dout  = 8'b11111111; // 1075 : 255 - 0xff
      12'h434: dout  = 8'b11111111; // 1076 : 255 - 0xff
      12'h435: dout  = 8'b11111111; // 1077 : 255 - 0xff
      12'h436: dout  = 8'b11111111; // 1078 : 255 - 0xff
      12'h437: dout  = 8'b11111111; // 1079 : 255 - 0xff
      12'h438: dout  = 8'b11111111; // 1080 : 255 - 0xff -- Sprite 0x87
      12'h439: dout  = 8'b11111111; // 1081 : 255 - 0xff
      12'h43A: dout  = 8'b11111111; // 1082 : 255 - 0xff
      12'h43B: dout  = 8'b11111111; // 1083 : 255 - 0xff
      12'h43C: dout  = 8'b11111111; // 1084 : 255 - 0xff
      12'h43D: dout  = 8'b11111111; // 1085 : 255 - 0xff
      12'h43E: dout  = 8'b11111111; // 1086 : 255 - 0xff
      12'h43F: dout  = 8'b11111111; // 1087 : 255 - 0xff
      12'h440: dout  = 8'b11111111; // 1088 : 255 - 0xff -- Sprite 0x88
      12'h441: dout  = 8'b11111111; // 1089 : 255 - 0xff
      12'h442: dout  = 8'b11111111; // 1090 : 255 - 0xff
      12'h443: dout  = 8'b11111111; // 1091 : 255 - 0xff
      12'h444: dout  = 8'b11111111; // 1092 : 255 - 0xff
      12'h445: dout  = 8'b11111111; // 1093 : 255 - 0xff
      12'h446: dout  = 8'b11111111; // 1094 : 255 - 0xff
      12'h447: dout  = 8'b11111111; // 1095 : 255 - 0xff
      12'h448: dout  = 8'b11111111; // 1096 : 255 - 0xff -- Sprite 0x89
      12'h449: dout  = 8'b11111111; // 1097 : 255 - 0xff
      12'h44A: dout  = 8'b11111111; // 1098 : 255 - 0xff
      12'h44B: dout  = 8'b11111111; // 1099 : 255 - 0xff
      12'h44C: dout  = 8'b11111111; // 1100 : 255 - 0xff
      12'h44D: dout  = 8'b11111111; // 1101 : 255 - 0xff
      12'h44E: dout  = 8'b11111111; // 1102 : 255 - 0xff
      12'h44F: dout  = 8'b11111111; // 1103 : 255 - 0xff
      12'h450: dout  = 8'b11111111; // 1104 : 255 - 0xff -- Sprite 0x8a
      12'h451: dout  = 8'b11111111; // 1105 : 255 - 0xff
      12'h452: dout  = 8'b11111111; // 1106 : 255 - 0xff
      12'h453: dout  = 8'b11111111; // 1107 : 255 - 0xff
      12'h454: dout  = 8'b11111111; // 1108 : 255 - 0xff
      12'h455: dout  = 8'b11111111; // 1109 : 255 - 0xff
      12'h456: dout  = 8'b11111111; // 1110 : 255 - 0xff
      12'h457: dout  = 8'b11111111; // 1111 : 255 - 0xff
      12'h458: dout  = 8'b11111111; // 1112 : 255 - 0xff -- Sprite 0x8b
      12'h459: dout  = 8'b11111111; // 1113 : 255 - 0xff
      12'h45A: dout  = 8'b11111111; // 1114 : 255 - 0xff
      12'h45B: dout  = 8'b11111111; // 1115 : 255 - 0xff
      12'h45C: dout  = 8'b11111111; // 1116 : 255 - 0xff
      12'h45D: dout  = 8'b11111111; // 1117 : 255 - 0xff
      12'h45E: dout  = 8'b11111111; // 1118 : 255 - 0xff
      12'h45F: dout  = 8'b11111111; // 1119 : 255 - 0xff
      12'h460: dout  = 8'b11111111; // 1120 : 255 - 0xff -- Sprite 0x8c
      12'h461: dout  = 8'b11111111; // 1121 : 255 - 0xff
      12'h462: dout  = 8'b11111111; // 1122 : 255 - 0xff
      12'h463: dout  = 8'b11111111; // 1123 : 255 - 0xff
      12'h464: dout  = 8'b11111111; // 1124 : 255 - 0xff
      12'h465: dout  = 8'b11111111; // 1125 : 255 - 0xff
      12'h466: dout  = 8'b11111111; // 1126 : 255 - 0xff
      12'h467: dout  = 8'b11111111; // 1127 : 255 - 0xff
      12'h468: dout  = 8'b11111111; // 1128 : 255 - 0xff -- Sprite 0x8d
      12'h469: dout  = 8'b11111111; // 1129 : 255 - 0xff
      12'h46A: dout  = 8'b11111111; // 1130 : 255 - 0xff
      12'h46B: dout  = 8'b11111111; // 1131 : 255 - 0xff
      12'h46C: dout  = 8'b11111111; // 1132 : 255 - 0xff
      12'h46D: dout  = 8'b11111111; // 1133 : 255 - 0xff
      12'h46E: dout  = 8'b11111111; // 1134 : 255 - 0xff
      12'h46F: dout  = 8'b11111111; // 1135 : 255 - 0xff
      12'h470: dout  = 8'b11111111; // 1136 : 255 - 0xff -- Sprite 0x8e
      12'h471: dout  = 8'b11111111; // 1137 : 255 - 0xff
      12'h472: dout  = 8'b11111111; // 1138 : 255 - 0xff
      12'h473: dout  = 8'b11111111; // 1139 : 255 - 0xff
      12'h474: dout  = 8'b11111111; // 1140 : 255 - 0xff
      12'h475: dout  = 8'b11111111; // 1141 : 255 - 0xff
      12'h476: dout  = 8'b11111111; // 1142 : 255 - 0xff
      12'h477: dout  = 8'b11111111; // 1143 : 255 - 0xff
      12'h478: dout  = 8'b11111111; // 1144 : 255 - 0xff -- Sprite 0x8f
      12'h479: dout  = 8'b11111111; // 1145 : 255 - 0xff
      12'h47A: dout  = 8'b11111111; // 1146 : 255 - 0xff
      12'h47B: dout  = 8'b11111111; // 1147 : 255 - 0xff
      12'h47C: dout  = 8'b11111111; // 1148 : 255 - 0xff
      12'h47D: dout  = 8'b11111111; // 1149 : 255 - 0xff
      12'h47E: dout  = 8'b11111111; // 1150 : 255 - 0xff
      12'h47F: dout  = 8'b11111111; // 1151 : 255 - 0xff
      12'h480: dout  = 8'b00000000; // 1152 :   0 - 0x0 -- Sprite 0x90
      12'h481: dout  = 8'b00000000; // 1153 :   0 - 0x0
      12'h482: dout  = 8'b00000000; // 1154 :   0 - 0x0
      12'h483: dout  = 8'b00000000; // 1155 :   0 - 0x0
      12'h484: dout  = 8'b00000000; // 1156 :   0 - 0x0
      12'h485: dout  = 8'b00000000; // 1157 :   0 - 0x0
      12'h486: dout  = 8'b00000000; // 1158 :   0 - 0x0
      12'h487: dout  = 8'b00000000; // 1159 :   0 - 0x0
      12'h488: dout  = 8'b00000000; // 1160 :   0 - 0x0 -- Sprite 0x91
      12'h489: dout  = 8'b00000000; // 1161 :   0 - 0x0
      12'h48A: dout  = 8'b00000000; // 1162 :   0 - 0x0
      12'h48B: dout  = 8'b00000000; // 1163 :   0 - 0x0
      12'h48C: dout  = 8'b00000000; // 1164 :   0 - 0x0
      12'h48D: dout  = 8'b00000000; // 1165 :   0 - 0x0
      12'h48E: dout  = 8'b00000000; // 1166 :   0 - 0x0
      12'h48F: dout  = 8'b00000000; // 1167 :   0 - 0x0
      12'h490: dout  = 8'b00000000; // 1168 :   0 - 0x0 -- Sprite 0x92
      12'h491: dout  = 8'b00000000; // 1169 :   0 - 0x0
      12'h492: dout  = 8'b00000000; // 1170 :   0 - 0x0
      12'h493: dout  = 8'b00000000; // 1171 :   0 - 0x0
      12'h494: dout  = 8'b00000000; // 1172 :   0 - 0x0
      12'h495: dout  = 8'b00000000; // 1173 :   0 - 0x0
      12'h496: dout  = 8'b00000000; // 1174 :   0 - 0x0
      12'h497: dout  = 8'b00000000; // 1175 :   0 - 0x0
      12'h498: dout  = 8'b00000000; // 1176 :   0 - 0x0 -- Sprite 0x93
      12'h499: dout  = 8'b00000000; // 1177 :   0 - 0x0
      12'h49A: dout  = 8'b00000000; // 1178 :   0 - 0x0
      12'h49B: dout  = 8'b00000000; // 1179 :   0 - 0x0
      12'h49C: dout  = 8'b00000000; // 1180 :   0 - 0x0
      12'h49D: dout  = 8'b00000000; // 1181 :   0 - 0x0
      12'h49E: dout  = 8'b00000000; // 1182 :   0 - 0x0
      12'h49F: dout  = 8'b00000000; // 1183 :   0 - 0x0
      12'h4A0: dout  = 8'b00000000; // 1184 :   0 - 0x0 -- Sprite 0x94
      12'h4A1: dout  = 8'b00000000; // 1185 :   0 - 0x0
      12'h4A2: dout  = 8'b00000000; // 1186 :   0 - 0x0
      12'h4A3: dout  = 8'b00000000; // 1187 :   0 - 0x0
      12'h4A4: dout  = 8'b00000000; // 1188 :   0 - 0x0
      12'h4A5: dout  = 8'b00000000; // 1189 :   0 - 0x0
      12'h4A6: dout  = 8'b00000000; // 1190 :   0 - 0x0
      12'h4A7: dout  = 8'b00000000; // 1191 :   0 - 0x0
      12'h4A8: dout  = 8'b00000000; // 1192 :   0 - 0x0 -- Sprite 0x95
      12'h4A9: dout  = 8'b00000000; // 1193 :   0 - 0x0
      12'h4AA: dout  = 8'b00000000; // 1194 :   0 - 0x0
      12'h4AB: dout  = 8'b00000000; // 1195 :   0 - 0x0
      12'h4AC: dout  = 8'b00000000; // 1196 :   0 - 0x0
      12'h4AD: dout  = 8'b00000000; // 1197 :   0 - 0x0
      12'h4AE: dout  = 8'b00000000; // 1198 :   0 - 0x0
      12'h4AF: dout  = 8'b00000000; // 1199 :   0 - 0x0
      12'h4B0: dout  = 8'b00000000; // 1200 :   0 - 0x0 -- Sprite 0x96
      12'h4B1: dout  = 8'b00000000; // 1201 :   0 - 0x0
      12'h4B2: dout  = 8'b00000000; // 1202 :   0 - 0x0
      12'h4B3: dout  = 8'b00000000; // 1203 :   0 - 0x0
      12'h4B4: dout  = 8'b00000000; // 1204 :   0 - 0x0
      12'h4B5: dout  = 8'b00000000; // 1205 :   0 - 0x0
      12'h4B6: dout  = 8'b00000000; // 1206 :   0 - 0x0
      12'h4B7: dout  = 8'b00000000; // 1207 :   0 - 0x0
      12'h4B8: dout  = 8'b00000000; // 1208 :   0 - 0x0 -- Sprite 0x97
      12'h4B9: dout  = 8'b00000000; // 1209 :   0 - 0x0
      12'h4BA: dout  = 8'b00000000; // 1210 :   0 - 0x0
      12'h4BB: dout  = 8'b00000000; // 1211 :   0 - 0x0
      12'h4BC: dout  = 8'b00000000; // 1212 :   0 - 0x0
      12'h4BD: dout  = 8'b00000000; // 1213 :   0 - 0x0
      12'h4BE: dout  = 8'b00000000; // 1214 :   0 - 0x0
      12'h4BF: dout  = 8'b00000000; // 1215 :   0 - 0x0
      12'h4C0: dout  = 8'b00000000; // 1216 :   0 - 0x0 -- Sprite 0x98
      12'h4C1: dout  = 8'b00000000; // 1217 :   0 - 0x0
      12'h4C2: dout  = 8'b00000000; // 1218 :   0 - 0x0
      12'h4C3: dout  = 8'b00000000; // 1219 :   0 - 0x0
      12'h4C4: dout  = 8'b00000000; // 1220 :   0 - 0x0
      12'h4C5: dout  = 8'b00000000; // 1221 :   0 - 0x0
      12'h4C6: dout  = 8'b00000000; // 1222 :   0 - 0x0
      12'h4C7: dout  = 8'b00000000; // 1223 :   0 - 0x0
      12'h4C8: dout  = 8'b00000000; // 1224 :   0 - 0x0 -- Sprite 0x99
      12'h4C9: dout  = 8'b00000000; // 1225 :   0 - 0x0
      12'h4CA: dout  = 8'b00000000; // 1226 :   0 - 0x0
      12'h4CB: dout  = 8'b00000000; // 1227 :   0 - 0x0
      12'h4CC: dout  = 8'b00000000; // 1228 :   0 - 0x0
      12'h4CD: dout  = 8'b00000000; // 1229 :   0 - 0x0
      12'h4CE: dout  = 8'b00000000; // 1230 :   0 - 0x0
      12'h4CF: dout  = 8'b00000000; // 1231 :   0 - 0x0
      12'h4D0: dout  = 8'b00000000; // 1232 :   0 - 0x0 -- Sprite 0x9a
      12'h4D1: dout  = 8'b00000000; // 1233 :   0 - 0x0
      12'h4D2: dout  = 8'b00000000; // 1234 :   0 - 0x0
      12'h4D3: dout  = 8'b00000000; // 1235 :   0 - 0x0
      12'h4D4: dout  = 8'b00000000; // 1236 :   0 - 0x0
      12'h4D5: dout  = 8'b00000000; // 1237 :   0 - 0x0
      12'h4D6: dout  = 8'b00000000; // 1238 :   0 - 0x0
      12'h4D7: dout  = 8'b00000000; // 1239 :   0 - 0x0
      12'h4D8: dout  = 8'b00000000; // 1240 :   0 - 0x0 -- Sprite 0x9b
      12'h4D9: dout  = 8'b00000000; // 1241 :   0 - 0x0
      12'h4DA: dout  = 8'b00000000; // 1242 :   0 - 0x0
      12'h4DB: dout  = 8'b00000000; // 1243 :   0 - 0x0
      12'h4DC: dout  = 8'b00000000; // 1244 :   0 - 0x0
      12'h4DD: dout  = 8'b00000000; // 1245 :   0 - 0x0
      12'h4DE: dout  = 8'b00000000; // 1246 :   0 - 0x0
      12'h4DF: dout  = 8'b00000000; // 1247 :   0 - 0x0
      12'h4E0: dout  = 8'b00000000; // 1248 :   0 - 0x0 -- Sprite 0x9c
      12'h4E1: dout  = 8'b00000000; // 1249 :   0 - 0x0
      12'h4E2: dout  = 8'b00000000; // 1250 :   0 - 0x0
      12'h4E3: dout  = 8'b00000000; // 1251 :   0 - 0x0
      12'h4E4: dout  = 8'b00000000; // 1252 :   0 - 0x0
      12'h4E5: dout  = 8'b00000000; // 1253 :   0 - 0x0
      12'h4E6: dout  = 8'b00000000; // 1254 :   0 - 0x0
      12'h4E7: dout  = 8'b00000000; // 1255 :   0 - 0x0
      12'h4E8: dout  = 8'b00000000; // 1256 :   0 - 0x0 -- Sprite 0x9d
      12'h4E9: dout  = 8'b00000000; // 1257 :   0 - 0x0
      12'h4EA: dout  = 8'b00000000; // 1258 :   0 - 0x0
      12'h4EB: dout  = 8'b00000000; // 1259 :   0 - 0x0
      12'h4EC: dout  = 8'b00000000; // 1260 :   0 - 0x0
      12'h4ED: dout  = 8'b00000000; // 1261 :   0 - 0x0
      12'h4EE: dout  = 8'b00000000; // 1262 :   0 - 0x0
      12'h4EF: dout  = 8'b00000000; // 1263 :   0 - 0x0
      12'h4F0: dout  = 8'b00000000; // 1264 :   0 - 0x0 -- Sprite 0x9e
      12'h4F1: dout  = 8'b00000000; // 1265 :   0 - 0x0
      12'h4F2: dout  = 8'b00000000; // 1266 :   0 - 0x0
      12'h4F3: dout  = 8'b00000000; // 1267 :   0 - 0x0
      12'h4F4: dout  = 8'b00000000; // 1268 :   0 - 0x0
      12'h4F5: dout  = 8'b00000000; // 1269 :   0 - 0x0
      12'h4F6: dout  = 8'b00000000; // 1270 :   0 - 0x0
      12'h4F7: dout  = 8'b00000000; // 1271 :   0 - 0x0
      12'h4F8: dout  = 8'b00000000; // 1272 :   0 - 0x0 -- Sprite 0x9f
      12'h4F9: dout  = 8'b00000000; // 1273 :   0 - 0x0
      12'h4FA: dout  = 8'b00000000; // 1274 :   0 - 0x0
      12'h4FB: dout  = 8'b00000000; // 1275 :   0 - 0x0
      12'h4FC: dout  = 8'b00000000; // 1276 :   0 - 0x0
      12'h4FD: dout  = 8'b00000000; // 1277 :   0 - 0x0
      12'h4FE: dout  = 8'b00000000; // 1278 :   0 - 0x0
      12'h4FF: dout  = 8'b00000000; // 1279 :   0 - 0x0
      12'h500: dout  = 8'b00000000; // 1280 :   0 - 0x0 -- Sprite 0xa0
      12'h501: dout  = 8'b00000000; // 1281 :   0 - 0x0
      12'h502: dout  = 8'b00000000; // 1282 :   0 - 0x0
      12'h503: dout  = 8'b00000000; // 1283 :   0 - 0x0
      12'h504: dout  = 8'b00000000; // 1284 :   0 - 0x0
      12'h505: dout  = 8'b00000000; // 1285 :   0 - 0x0
      12'h506: dout  = 8'b00000000; // 1286 :   0 - 0x0
      12'h507: dout  = 8'b00000000; // 1287 :   0 - 0x0
      12'h508: dout  = 8'b00000000; // 1288 :   0 - 0x0 -- Sprite 0xa1
      12'h509: dout  = 8'b00000000; // 1289 :   0 - 0x0
      12'h50A: dout  = 8'b00000000; // 1290 :   0 - 0x0
      12'h50B: dout  = 8'b00000000; // 1291 :   0 - 0x0
      12'h50C: dout  = 8'b00000000; // 1292 :   0 - 0x0
      12'h50D: dout  = 8'b00000000; // 1293 :   0 - 0x0
      12'h50E: dout  = 8'b00000000; // 1294 :   0 - 0x0
      12'h50F: dout  = 8'b00000000; // 1295 :   0 - 0x0
      12'h510: dout  = 8'b00000000; // 1296 :   0 - 0x0 -- Sprite 0xa2
      12'h511: dout  = 8'b00000000; // 1297 :   0 - 0x0
      12'h512: dout  = 8'b00000000; // 1298 :   0 - 0x0
      12'h513: dout  = 8'b00000000; // 1299 :   0 - 0x0
      12'h514: dout  = 8'b00000000; // 1300 :   0 - 0x0
      12'h515: dout  = 8'b00000000; // 1301 :   0 - 0x0
      12'h516: dout  = 8'b00000000; // 1302 :   0 - 0x0
      12'h517: dout  = 8'b00000000; // 1303 :   0 - 0x0
      12'h518: dout  = 8'b00000000; // 1304 :   0 - 0x0 -- Sprite 0xa3
      12'h519: dout  = 8'b00000000; // 1305 :   0 - 0x0
      12'h51A: dout  = 8'b00000000; // 1306 :   0 - 0x0
      12'h51B: dout  = 8'b00000000; // 1307 :   0 - 0x0
      12'h51C: dout  = 8'b00000000; // 1308 :   0 - 0x0
      12'h51D: dout  = 8'b00000000; // 1309 :   0 - 0x0
      12'h51E: dout  = 8'b00000000; // 1310 :   0 - 0x0
      12'h51F: dout  = 8'b00000000; // 1311 :   0 - 0x0
      12'h520: dout  = 8'b00000000; // 1312 :   0 - 0x0 -- Sprite 0xa4
      12'h521: dout  = 8'b00000000; // 1313 :   0 - 0x0
      12'h522: dout  = 8'b00000000; // 1314 :   0 - 0x0
      12'h523: dout  = 8'b00000000; // 1315 :   0 - 0x0
      12'h524: dout  = 8'b00000000; // 1316 :   0 - 0x0
      12'h525: dout  = 8'b00000000; // 1317 :   0 - 0x0
      12'h526: dout  = 8'b00000000; // 1318 :   0 - 0x0
      12'h527: dout  = 8'b00000000; // 1319 :   0 - 0x0
      12'h528: dout  = 8'b00000000; // 1320 :   0 - 0x0 -- Sprite 0xa5
      12'h529: dout  = 8'b00000000; // 1321 :   0 - 0x0
      12'h52A: dout  = 8'b00000000; // 1322 :   0 - 0x0
      12'h52B: dout  = 8'b00000000; // 1323 :   0 - 0x0
      12'h52C: dout  = 8'b00000000; // 1324 :   0 - 0x0
      12'h52D: dout  = 8'b00000000; // 1325 :   0 - 0x0
      12'h52E: dout  = 8'b00000000; // 1326 :   0 - 0x0
      12'h52F: dout  = 8'b00000000; // 1327 :   0 - 0x0
      12'h530: dout  = 8'b00000000; // 1328 :   0 - 0x0 -- Sprite 0xa6
      12'h531: dout  = 8'b00000000; // 1329 :   0 - 0x0
      12'h532: dout  = 8'b00000000; // 1330 :   0 - 0x0
      12'h533: dout  = 8'b00000000; // 1331 :   0 - 0x0
      12'h534: dout  = 8'b00000000; // 1332 :   0 - 0x0
      12'h535: dout  = 8'b00000000; // 1333 :   0 - 0x0
      12'h536: dout  = 8'b00000000; // 1334 :   0 - 0x0
      12'h537: dout  = 8'b00000000; // 1335 :   0 - 0x0
      12'h538: dout  = 8'b00000000; // 1336 :   0 - 0x0 -- Sprite 0xa7
      12'h539: dout  = 8'b00000000; // 1337 :   0 - 0x0
      12'h53A: dout  = 8'b00000000; // 1338 :   0 - 0x0
      12'h53B: dout  = 8'b00000000; // 1339 :   0 - 0x0
      12'h53C: dout  = 8'b00000000; // 1340 :   0 - 0x0
      12'h53D: dout  = 8'b00000000; // 1341 :   0 - 0x0
      12'h53E: dout  = 8'b00000000; // 1342 :   0 - 0x0
      12'h53F: dout  = 8'b00000000; // 1343 :   0 - 0x0
      12'h540: dout  = 8'b00000000; // 1344 :   0 - 0x0 -- Sprite 0xa8
      12'h541: dout  = 8'b00000000; // 1345 :   0 - 0x0
      12'h542: dout  = 8'b00000000; // 1346 :   0 - 0x0
      12'h543: dout  = 8'b00000000; // 1347 :   0 - 0x0
      12'h544: dout  = 8'b00000000; // 1348 :   0 - 0x0
      12'h545: dout  = 8'b00000000; // 1349 :   0 - 0x0
      12'h546: dout  = 8'b00000000; // 1350 :   0 - 0x0
      12'h547: dout  = 8'b00000000; // 1351 :   0 - 0x0
      12'h548: dout  = 8'b00000000; // 1352 :   0 - 0x0 -- Sprite 0xa9
      12'h549: dout  = 8'b00000000; // 1353 :   0 - 0x0
      12'h54A: dout  = 8'b00000000; // 1354 :   0 - 0x0
      12'h54B: dout  = 8'b00000000; // 1355 :   0 - 0x0
      12'h54C: dout  = 8'b00000000; // 1356 :   0 - 0x0
      12'h54D: dout  = 8'b00000000; // 1357 :   0 - 0x0
      12'h54E: dout  = 8'b00000000; // 1358 :   0 - 0x0
      12'h54F: dout  = 8'b00000000; // 1359 :   0 - 0x0
      12'h550: dout  = 8'b00000000; // 1360 :   0 - 0x0 -- Sprite 0xaa
      12'h551: dout  = 8'b00000000; // 1361 :   0 - 0x0
      12'h552: dout  = 8'b00000000; // 1362 :   0 - 0x0
      12'h553: dout  = 8'b00000000; // 1363 :   0 - 0x0
      12'h554: dout  = 8'b00000000; // 1364 :   0 - 0x0
      12'h555: dout  = 8'b00000000; // 1365 :   0 - 0x0
      12'h556: dout  = 8'b00000000; // 1366 :   0 - 0x0
      12'h557: dout  = 8'b00000000; // 1367 :   0 - 0x0
      12'h558: dout  = 8'b00000000; // 1368 :   0 - 0x0 -- Sprite 0xab
      12'h559: dout  = 8'b00000000; // 1369 :   0 - 0x0
      12'h55A: dout  = 8'b00000000; // 1370 :   0 - 0x0
      12'h55B: dout  = 8'b00000000; // 1371 :   0 - 0x0
      12'h55C: dout  = 8'b00000000; // 1372 :   0 - 0x0
      12'h55D: dout  = 8'b00000000; // 1373 :   0 - 0x0
      12'h55E: dout  = 8'b00000000; // 1374 :   0 - 0x0
      12'h55F: dout  = 8'b00000000; // 1375 :   0 - 0x0
      12'h560: dout  = 8'b00000000; // 1376 :   0 - 0x0 -- Sprite 0xac
      12'h561: dout  = 8'b00000000; // 1377 :   0 - 0x0
      12'h562: dout  = 8'b00000000; // 1378 :   0 - 0x0
      12'h563: dout  = 8'b00000000; // 1379 :   0 - 0x0
      12'h564: dout  = 8'b00000000; // 1380 :   0 - 0x0
      12'h565: dout  = 8'b00000000; // 1381 :   0 - 0x0
      12'h566: dout  = 8'b00000000; // 1382 :   0 - 0x0
      12'h567: dout  = 8'b00000000; // 1383 :   0 - 0x0
      12'h568: dout  = 8'b00000000; // 1384 :   0 - 0x0 -- Sprite 0xad
      12'h569: dout  = 8'b00000000; // 1385 :   0 - 0x0
      12'h56A: dout  = 8'b00000000; // 1386 :   0 - 0x0
      12'h56B: dout  = 8'b00000000; // 1387 :   0 - 0x0
      12'h56C: dout  = 8'b00000000; // 1388 :   0 - 0x0
      12'h56D: dout  = 8'b00000000; // 1389 :   0 - 0x0
      12'h56E: dout  = 8'b00000000; // 1390 :   0 - 0x0
      12'h56F: dout  = 8'b00000000; // 1391 :   0 - 0x0
      12'h570: dout  = 8'b00000000; // 1392 :   0 - 0x0 -- Sprite 0xae
      12'h571: dout  = 8'b00000000; // 1393 :   0 - 0x0
      12'h572: dout  = 8'b00000000; // 1394 :   0 - 0x0
      12'h573: dout  = 8'b00000000; // 1395 :   0 - 0x0
      12'h574: dout  = 8'b00000000; // 1396 :   0 - 0x0
      12'h575: dout  = 8'b00000000; // 1397 :   0 - 0x0
      12'h576: dout  = 8'b00000000; // 1398 :   0 - 0x0
      12'h577: dout  = 8'b00000000; // 1399 :   0 - 0x0
      12'h578: dout  = 8'b00000000; // 1400 :   0 - 0x0 -- Sprite 0xaf
      12'h579: dout  = 8'b00000000; // 1401 :   0 - 0x0
      12'h57A: dout  = 8'b00000000; // 1402 :   0 - 0x0
      12'h57B: dout  = 8'b00000000; // 1403 :   0 - 0x0
      12'h57C: dout  = 8'b00000000; // 1404 :   0 - 0x0
      12'h57D: dout  = 8'b00000000; // 1405 :   0 - 0x0
      12'h57E: dout  = 8'b00000000; // 1406 :   0 - 0x0
      12'h57F: dout  = 8'b00000000; // 1407 :   0 - 0x0
      12'h580: dout  = 8'b01111110; // 1408 : 126 - 0x7e -- Sprite 0xb0
      12'h581: dout  = 8'b01100011; // 1409 :  99 - 0x63
      12'h582: dout  = 8'b01100011; // 1410 :  99 - 0x63
      12'h583: dout  = 8'b01100011; // 1411 :  99 - 0x63
      12'h584: dout  = 8'b01111110; // 1412 : 126 - 0x7e
      12'h585: dout  = 8'b01100000; // 1413 :  96 - 0x60
      12'h586: dout  = 8'b01100000; // 1414 :  96 - 0x60
      12'h587: dout  = 8'b00000000; // 1415 :   0 - 0x0
      12'h588: dout  = 8'b01100000; // 1416 :  96 - 0x60 -- Sprite 0xb1
      12'h589: dout  = 8'b01100000; // 1417 :  96 - 0x60
      12'h58A: dout  = 8'b01100000; // 1418 :  96 - 0x60
      12'h58B: dout  = 8'b01100000; // 1419 :  96 - 0x60
      12'h58C: dout  = 8'b01100000; // 1420 :  96 - 0x60
      12'h58D: dout  = 8'b01100000; // 1421 :  96 - 0x60
      12'h58E: dout  = 8'b01111111; // 1422 : 127 - 0x7f
      12'h58F: dout  = 8'b00000000; // 1423 :   0 - 0x0
      12'h590: dout  = 8'b00011100; // 1424 :  28 - 0x1c -- Sprite 0xb2
      12'h591: dout  = 8'b00110110; // 1425 :  54 - 0x36
      12'h592: dout  = 8'b01100011; // 1426 :  99 - 0x63
      12'h593: dout  = 8'b01100011; // 1427 :  99 - 0x63
      12'h594: dout  = 8'b01111111; // 1428 : 127 - 0x7f
      12'h595: dout  = 8'b01100011; // 1429 :  99 - 0x63
      12'h596: dout  = 8'b01100011; // 1430 :  99 - 0x63
      12'h597: dout  = 8'b00000000; // 1431 :   0 - 0x0
      12'h598: dout  = 8'b00110011; // 1432 :  51 - 0x33 -- Sprite 0xb3
      12'h599: dout  = 8'b00110011; // 1433 :  51 - 0x33
      12'h59A: dout  = 8'b00110011; // 1434 :  51 - 0x33
      12'h59B: dout  = 8'b00011110; // 1435 :  30 - 0x1e
      12'h59C: dout  = 8'b00001100; // 1436 :  12 - 0xc
      12'h59D: dout  = 8'b00001100; // 1437 :  12 - 0xc
      12'h59E: dout  = 8'b00001100; // 1438 :  12 - 0xc
      12'h59F: dout  = 8'b00000000; // 1439 :   0 - 0x0
      12'h5A0: dout  = 8'b01111111; // 1440 : 127 - 0x7f -- Sprite 0xb4
      12'h5A1: dout  = 8'b01100000; // 1441 :  96 - 0x60
      12'h5A2: dout  = 8'b01100000; // 1442 :  96 - 0x60
      12'h5A3: dout  = 8'b01111110; // 1443 : 126 - 0x7e
      12'h5A4: dout  = 8'b01100000; // 1444 :  96 - 0x60
      12'h5A5: dout  = 8'b01100000; // 1445 :  96 - 0x60
      12'h5A6: dout  = 8'b01111111; // 1446 : 127 - 0x7f
      12'h5A7: dout  = 8'b00000000; // 1447 :   0 - 0x0
      12'h5A8: dout  = 8'b01111110; // 1448 : 126 - 0x7e -- Sprite 0xb5
      12'h5A9: dout  = 8'b01100011; // 1449 :  99 - 0x63
      12'h5AA: dout  = 8'b01100011; // 1450 :  99 - 0x63
      12'h5AB: dout  = 8'b01100111; // 1451 : 103 - 0x67
      12'h5AC: dout  = 8'b01111100; // 1452 : 124 - 0x7c
      12'h5AD: dout  = 8'b01101110; // 1453 : 110 - 0x6e
      12'h5AE: dout  = 8'b01100111; // 1454 : 103 - 0x67
      12'h5AF: dout  = 8'b00000000; // 1455 :   0 - 0x0
      12'h5B0: dout  = 8'b00111110; // 1456 :  62 - 0x3e -- Sprite 0xb6
      12'h5B1: dout  = 8'b01100011; // 1457 :  99 - 0x63
      12'h5B2: dout  = 8'b01100011; // 1458 :  99 - 0x63
      12'h5B3: dout  = 8'b01100011; // 1459 :  99 - 0x63
      12'h5B4: dout  = 8'b01100011; // 1460 :  99 - 0x63
      12'h5B5: dout  = 8'b01100011; // 1461 :  99 - 0x63
      12'h5B6: dout  = 8'b00111110; // 1462 :  62 - 0x3e
      12'h5B7: dout  = 8'b00000000; // 1463 :   0 - 0x0
      12'h5B8: dout  = 8'b01100011; // 1464 :  99 - 0x63 -- Sprite 0xb7
      12'h5B9: dout  = 8'b01110011; // 1465 : 115 - 0x73
      12'h5BA: dout  = 8'b01111011; // 1466 : 123 - 0x7b
      12'h5BB: dout  = 8'b01111111; // 1467 : 127 - 0x7f
      12'h5BC: dout  = 8'b01101111; // 1468 : 111 - 0x6f
      12'h5BD: dout  = 8'b01100111; // 1469 : 103 - 0x67
      12'h5BE: dout  = 8'b01100011; // 1470 :  99 - 0x63
      12'h5BF: dout  = 8'b00000000; // 1471 :   0 - 0x0
      12'h5C0: dout  = 8'b00111111; // 1472 :  63 - 0x3f -- Sprite 0xb8
      12'h5C1: dout  = 8'b00001100; // 1473 :  12 - 0xc
      12'h5C2: dout  = 8'b00001100; // 1474 :  12 - 0xc
      12'h5C3: dout  = 8'b00001100; // 1475 :  12 - 0xc
      12'h5C4: dout  = 8'b00001100; // 1476 :  12 - 0xc
      12'h5C5: dout  = 8'b00001100; // 1477 :  12 - 0xc
      12'h5C6: dout  = 8'b00001100; // 1478 :  12 - 0xc
      12'h5C7: dout  = 8'b00000000; // 1479 :   0 - 0x0
      12'h5C8: dout  = 8'b01100011; // 1480 :  99 - 0x63 -- Sprite 0xb9
      12'h5C9: dout  = 8'b01100011; // 1481 :  99 - 0x63
      12'h5CA: dout  = 8'b01101011; // 1482 : 107 - 0x6b
      12'h5CB: dout  = 8'b01111111; // 1483 : 127 - 0x7f
      12'h5CC: dout  = 8'b01111111; // 1484 : 127 - 0x7f
      12'h5CD: dout  = 8'b01110111; // 1485 : 119 - 0x77
      12'h5CE: dout  = 8'b01100011; // 1486 :  99 - 0x63
      12'h5CF: dout  = 8'b00000000; // 1487 :   0 - 0x0
      12'h5D0: dout  = 8'b00000000; // 1488 :   0 - 0x0 -- Sprite 0xba
      12'h5D1: dout  = 8'b00000000; // 1489 :   0 - 0x0
      12'h5D2: dout  = 8'b00000000; // 1490 :   0 - 0x0
      12'h5D3: dout  = 8'b00000000; // 1491 :   0 - 0x0
      12'h5D4: dout  = 8'b00000000; // 1492 :   0 - 0x0
      12'h5D5: dout  = 8'b00000000; // 1493 :   0 - 0x0
      12'h5D6: dout  = 8'b00000000; // 1494 :   0 - 0x0
      12'h5D7: dout  = 8'b00000000; // 1495 :   0 - 0x0
      12'h5D8: dout  = 8'b00000000; // 1496 :   0 - 0x0 -- Sprite 0xbb
      12'h5D9: dout  = 8'b00000000; // 1497 :   0 - 0x0
      12'h5DA: dout  = 8'b00000000; // 1498 :   0 - 0x0
      12'h5DB: dout  = 8'b00000000; // 1499 :   0 - 0x0
      12'h5DC: dout  = 8'b00000000; // 1500 :   0 - 0x0
      12'h5DD: dout  = 8'b00000000; // 1501 :   0 - 0x0
      12'h5DE: dout  = 8'b00000000; // 1502 :   0 - 0x0
      12'h5DF: dout  = 8'b00000000; // 1503 :   0 - 0x0
      12'h5E0: dout  = 8'b00011111; // 1504 :  31 - 0x1f -- Sprite 0xbc
      12'h5E1: dout  = 8'b00110000; // 1505 :  48 - 0x30
      12'h5E2: dout  = 8'b01100000; // 1506 :  96 - 0x60
      12'h5E3: dout  = 8'b01100111; // 1507 : 103 - 0x67
      12'h5E4: dout  = 8'b01100011; // 1508 :  99 - 0x63
      12'h5E5: dout  = 8'b00110011; // 1509 :  51 - 0x33
      12'h5E6: dout  = 8'b00011111; // 1510 :  31 - 0x1f
      12'h5E7: dout  = 8'b00000000; // 1511 :   0 - 0x0
      12'h5E8: dout  = 8'b01100011; // 1512 :  99 - 0x63 -- Sprite 0xbd
      12'h5E9: dout  = 8'b01110111; // 1513 : 119 - 0x77
      12'h5EA: dout  = 8'b01111111; // 1514 : 127 - 0x7f
      12'h5EB: dout  = 8'b01111111; // 1515 : 127 - 0x7f
      12'h5EC: dout  = 8'b01101011; // 1516 : 107 - 0x6b
      12'h5ED: dout  = 8'b01100011; // 1517 :  99 - 0x63
      12'h5EE: dout  = 8'b01100011; // 1518 :  99 - 0x63
      12'h5EF: dout  = 8'b00000000; // 1519 :   0 - 0x0
      12'h5F0: dout  = 8'b01100011; // 1520 :  99 - 0x63 -- Sprite 0xbe
      12'h5F1: dout  = 8'b01100011; // 1521 :  99 - 0x63
      12'h5F2: dout  = 8'b01100011; // 1522 :  99 - 0x63
      12'h5F3: dout  = 8'b01110111; // 1523 : 119 - 0x77
      12'h5F4: dout  = 8'b00111110; // 1524 :  62 - 0x3e
      12'h5F5: dout  = 8'b00011100; // 1525 :  28 - 0x1c
      12'h5F6: dout  = 8'b00001000; // 1526 :   8 - 0x8
      12'h5F7: dout  = 8'b00000000; // 1527 :   0 - 0x0
      12'h5F8: dout  = 8'b00000000; // 1528 :   0 - 0x0 -- Sprite 0xbf
      12'h5F9: dout  = 8'b00000000; // 1529 :   0 - 0x0
      12'h5FA: dout  = 8'b00000000; // 1530 :   0 - 0x0
      12'h5FB: dout  = 8'b00000000; // 1531 :   0 - 0x0
      12'h5FC: dout  = 8'b00000000; // 1532 :   0 - 0x0
      12'h5FD: dout  = 8'b00000000; // 1533 :   0 - 0x0
      12'h5FE: dout  = 8'b00000000; // 1534 :   0 - 0x0
      12'h5FF: dout  = 8'b00000000; // 1535 :   0 - 0x0
      12'h600: dout  = 8'b00000000; // 1536 :   0 - 0x0 -- Sprite 0xc0
      12'h601: dout  = 8'b00000000; // 1537 :   0 - 0x0
      12'h602: dout  = 8'b00000000; // 1538 :   0 - 0x0
      12'h603: dout  = 8'b00000000; // 1539 :   0 - 0x0
      12'h604: dout  = 8'b00000000; // 1540 :   0 - 0x0
      12'h605: dout  = 8'b00000000; // 1541 :   0 - 0x0
      12'h606: dout  = 8'b00000000; // 1542 :   0 - 0x0
      12'h607: dout  = 8'b00000000; // 1543 :   0 - 0x0
      12'h608: dout  = 8'b00000000; // 1544 :   0 - 0x0 -- Sprite 0xc1
      12'h609: dout  = 8'b00000000; // 1545 :   0 - 0x0
      12'h60A: dout  = 8'b00000000; // 1546 :   0 - 0x0
      12'h60B: dout  = 8'b00000000; // 1547 :   0 - 0x0
      12'h60C: dout  = 8'b00000000; // 1548 :   0 - 0x0
      12'h60D: dout  = 8'b00000000; // 1549 :   0 - 0x0
      12'h60E: dout  = 8'b00000000; // 1550 :   0 - 0x0
      12'h60F: dout  = 8'b00000000; // 1551 :   0 - 0x0
      12'h610: dout  = 8'b00000000; // 1552 :   0 - 0x0 -- Sprite 0xc2
      12'h611: dout  = 8'b00000000; // 1553 :   0 - 0x0
      12'h612: dout  = 8'b00000000; // 1554 :   0 - 0x0
      12'h613: dout  = 8'b00000000; // 1555 :   0 - 0x0
      12'h614: dout  = 8'b00000000; // 1556 :   0 - 0x0
      12'h615: dout  = 8'b00000000; // 1557 :   0 - 0x0
      12'h616: dout  = 8'b00000000; // 1558 :   0 - 0x0
      12'h617: dout  = 8'b00000000; // 1559 :   0 - 0x0
      12'h618: dout  = 8'b00000000; // 1560 :   0 - 0x0 -- Sprite 0xc3
      12'h619: dout  = 8'b00000000; // 1561 :   0 - 0x0
      12'h61A: dout  = 8'b00000000; // 1562 :   0 - 0x0
      12'h61B: dout  = 8'b00000000; // 1563 :   0 - 0x0
      12'h61C: dout  = 8'b00000000; // 1564 :   0 - 0x0
      12'h61D: dout  = 8'b00000000; // 1565 :   0 - 0x0
      12'h61E: dout  = 8'b00000000; // 1566 :   0 - 0x0
      12'h61F: dout  = 8'b00000000; // 1567 :   0 - 0x0
      12'h620: dout  = 8'b00000000; // 1568 :   0 - 0x0 -- Sprite 0xc4
      12'h621: dout  = 8'b00000000; // 1569 :   0 - 0x0
      12'h622: dout  = 8'b00000000; // 1570 :   0 - 0x0
      12'h623: dout  = 8'b00000000; // 1571 :   0 - 0x0
      12'h624: dout  = 8'b00000000; // 1572 :   0 - 0x0
      12'h625: dout  = 8'b00000000; // 1573 :   0 - 0x0
      12'h626: dout  = 8'b00000000; // 1574 :   0 - 0x0
      12'h627: dout  = 8'b00000000; // 1575 :   0 - 0x0
      12'h628: dout  = 8'b00000000; // 1576 :   0 - 0x0 -- Sprite 0xc5
      12'h629: dout  = 8'b00000000; // 1577 :   0 - 0x0
      12'h62A: dout  = 8'b00000000; // 1578 :   0 - 0x0
      12'h62B: dout  = 8'b00000000; // 1579 :   0 - 0x0
      12'h62C: dout  = 8'b00000000; // 1580 :   0 - 0x0
      12'h62D: dout  = 8'b00000000; // 1581 :   0 - 0x0
      12'h62E: dout  = 8'b00000000; // 1582 :   0 - 0x0
      12'h62F: dout  = 8'b00000000; // 1583 :   0 - 0x0
      12'h630: dout  = 8'b00000000; // 1584 :   0 - 0x0 -- Sprite 0xc6
      12'h631: dout  = 8'b00000000; // 1585 :   0 - 0x0
      12'h632: dout  = 8'b00000000; // 1586 :   0 - 0x0
      12'h633: dout  = 8'b00000000; // 1587 :   0 - 0x0
      12'h634: dout  = 8'b00000000; // 1588 :   0 - 0x0
      12'h635: dout  = 8'b00000000; // 1589 :   0 - 0x0
      12'h636: dout  = 8'b00000000; // 1590 :   0 - 0x0
      12'h637: dout  = 8'b00000000; // 1591 :   0 - 0x0
      12'h638: dout  = 8'b00000000; // 1592 :   0 - 0x0 -- Sprite 0xc7
      12'h639: dout  = 8'b00000000; // 1593 :   0 - 0x0
      12'h63A: dout  = 8'b00000000; // 1594 :   0 - 0x0
      12'h63B: dout  = 8'b00000000; // 1595 :   0 - 0x0
      12'h63C: dout  = 8'b00000000; // 1596 :   0 - 0x0
      12'h63D: dout  = 8'b00000000; // 1597 :   0 - 0x0
      12'h63E: dout  = 8'b00000000; // 1598 :   0 - 0x0
      12'h63F: dout  = 8'b00000000; // 1599 :   0 - 0x0
      12'h640: dout  = 8'b00000000; // 1600 :   0 - 0x0 -- Sprite 0xc8
      12'h641: dout  = 8'b00000000; // 1601 :   0 - 0x0
      12'h642: dout  = 8'b00000000; // 1602 :   0 - 0x0
      12'h643: dout  = 8'b00000000; // 1603 :   0 - 0x0
      12'h644: dout  = 8'b00000000; // 1604 :   0 - 0x0
      12'h645: dout  = 8'b00000000; // 1605 :   0 - 0x0
      12'h646: dout  = 8'b00000000; // 1606 :   0 - 0x0
      12'h647: dout  = 8'b00000000; // 1607 :   0 - 0x0
      12'h648: dout  = 8'b00000000; // 1608 :   0 - 0x0 -- Sprite 0xc9
      12'h649: dout  = 8'b00000000; // 1609 :   0 - 0x0
      12'h64A: dout  = 8'b00000000; // 1610 :   0 - 0x0
      12'h64B: dout  = 8'b00000000; // 1611 :   0 - 0x0
      12'h64C: dout  = 8'b00000000; // 1612 :   0 - 0x0
      12'h64D: dout  = 8'b00000000; // 1613 :   0 - 0x0
      12'h64E: dout  = 8'b00000000; // 1614 :   0 - 0x0
      12'h64F: dout  = 8'b00000000; // 1615 :   0 - 0x0
      12'h650: dout  = 8'b00000000; // 1616 :   0 - 0x0 -- Sprite 0xca
      12'h651: dout  = 8'b00000000; // 1617 :   0 - 0x0
      12'h652: dout  = 8'b00000000; // 1618 :   0 - 0x0
      12'h653: dout  = 8'b00000000; // 1619 :   0 - 0x0
      12'h654: dout  = 8'b00000000; // 1620 :   0 - 0x0
      12'h655: dout  = 8'b00000000; // 1621 :   0 - 0x0
      12'h656: dout  = 8'b00000000; // 1622 :   0 - 0x0
      12'h657: dout  = 8'b00000000; // 1623 :   0 - 0x0
      12'h658: dout  = 8'b00000000; // 1624 :   0 - 0x0 -- Sprite 0xcb
      12'h659: dout  = 8'b00000000; // 1625 :   0 - 0x0
      12'h65A: dout  = 8'b00000000; // 1626 :   0 - 0x0
      12'h65B: dout  = 8'b00000000; // 1627 :   0 - 0x0
      12'h65C: dout  = 8'b00000000; // 1628 :   0 - 0x0
      12'h65D: dout  = 8'b00000000; // 1629 :   0 - 0x0
      12'h65E: dout  = 8'b00000000; // 1630 :   0 - 0x0
      12'h65F: dout  = 8'b00000000; // 1631 :   0 - 0x0
      12'h660: dout  = 8'b00000000; // 1632 :   0 - 0x0 -- Sprite 0xcc
      12'h661: dout  = 8'b00000000; // 1633 :   0 - 0x0
      12'h662: dout  = 8'b00000000; // 1634 :   0 - 0x0
      12'h663: dout  = 8'b00000000; // 1635 :   0 - 0x0
      12'h664: dout  = 8'b00000000; // 1636 :   0 - 0x0
      12'h665: dout  = 8'b00000000; // 1637 :   0 - 0x0
      12'h666: dout  = 8'b00000000; // 1638 :   0 - 0x0
      12'h667: dout  = 8'b00000000; // 1639 :   0 - 0x0
      12'h668: dout  = 8'b00000000; // 1640 :   0 - 0x0 -- Sprite 0xcd
      12'h669: dout  = 8'b00000000; // 1641 :   0 - 0x0
      12'h66A: dout  = 8'b00000000; // 1642 :   0 - 0x0
      12'h66B: dout  = 8'b00000000; // 1643 :   0 - 0x0
      12'h66C: dout  = 8'b00000000; // 1644 :   0 - 0x0
      12'h66D: dout  = 8'b00000000; // 1645 :   0 - 0x0
      12'h66E: dout  = 8'b00000000; // 1646 :   0 - 0x0
      12'h66F: dout  = 8'b00000000; // 1647 :   0 - 0x0
      12'h670: dout  = 8'b00000000; // 1648 :   0 - 0x0 -- Sprite 0xce
      12'h671: dout  = 8'b00000000; // 1649 :   0 - 0x0
      12'h672: dout  = 8'b00000000; // 1650 :   0 - 0x0
      12'h673: dout  = 8'b00000000; // 1651 :   0 - 0x0
      12'h674: dout  = 8'b00000000; // 1652 :   0 - 0x0
      12'h675: dout  = 8'b00000000; // 1653 :   0 - 0x0
      12'h676: dout  = 8'b00000000; // 1654 :   0 - 0x0
      12'h677: dout  = 8'b00000000; // 1655 :   0 - 0x0
      12'h678: dout  = 8'b00000000; // 1656 :   0 - 0x0 -- Sprite 0xcf
      12'h679: dout  = 8'b00000000; // 1657 :   0 - 0x0
      12'h67A: dout  = 8'b00000000; // 1658 :   0 - 0x0
      12'h67B: dout  = 8'b00000000; // 1659 :   0 - 0x0
      12'h67C: dout  = 8'b00000000; // 1660 :   0 - 0x0
      12'h67D: dout  = 8'b00000000; // 1661 :   0 - 0x0
      12'h67E: dout  = 8'b00000000; // 1662 :   0 - 0x0
      12'h67F: dout  = 8'b00000000; // 1663 :   0 - 0x0
      12'h680: dout  = 8'b11111111; // 1664 : 255 - 0xff -- Sprite 0xd0
      12'h681: dout  = 8'b11111111; // 1665 : 255 - 0xff
      12'h682: dout  = 8'b11111111; // 1666 : 255 - 0xff
      12'h683: dout  = 8'b11111111; // 1667 : 255 - 0xff
      12'h684: dout  = 8'b11111111; // 1668 : 255 - 0xff
      12'h685: dout  = 8'b11111111; // 1669 : 255 - 0xff
      12'h686: dout  = 8'b11111111; // 1670 : 255 - 0xff
      12'h687: dout  = 8'b11111111; // 1671 : 255 - 0xff
      12'h688: dout  = 8'b11111111; // 1672 : 255 - 0xff -- Sprite 0xd1
      12'h689: dout  = 8'b11111111; // 1673 : 255 - 0xff
      12'h68A: dout  = 8'b11111111; // 1674 : 255 - 0xff
      12'h68B: dout  = 8'b11111111; // 1675 : 255 - 0xff
      12'h68C: dout  = 8'b11111111; // 1676 : 255 - 0xff
      12'h68D: dout  = 8'b11111111; // 1677 : 255 - 0xff
      12'h68E: dout  = 8'b11111111; // 1678 : 255 - 0xff
      12'h68F: dout  = 8'b11111111; // 1679 : 255 - 0xff
      12'h690: dout  = 8'b11111111; // 1680 : 255 - 0xff -- Sprite 0xd2
      12'h691: dout  = 8'b11111111; // 1681 : 255 - 0xff
      12'h692: dout  = 8'b11111111; // 1682 : 255 - 0xff
      12'h693: dout  = 8'b11111111; // 1683 : 255 - 0xff
      12'h694: dout  = 8'b11111111; // 1684 : 255 - 0xff
      12'h695: dout  = 8'b11111111; // 1685 : 255 - 0xff
      12'h696: dout  = 8'b11111111; // 1686 : 255 - 0xff
      12'h697: dout  = 8'b11111111; // 1687 : 255 - 0xff
      12'h698: dout  = 8'b11111111; // 1688 : 255 - 0xff -- Sprite 0xd3
      12'h699: dout  = 8'b11111111; // 1689 : 255 - 0xff
      12'h69A: dout  = 8'b11111111; // 1690 : 255 - 0xff
      12'h69B: dout  = 8'b11111111; // 1691 : 255 - 0xff
      12'h69C: dout  = 8'b11111111; // 1692 : 255 - 0xff
      12'h69D: dout  = 8'b11111111; // 1693 : 255 - 0xff
      12'h69E: dout  = 8'b11111111; // 1694 : 255 - 0xff
      12'h69F: dout  = 8'b11111111; // 1695 : 255 - 0xff
      12'h6A0: dout  = 8'b11111111; // 1696 : 255 - 0xff -- Sprite 0xd4
      12'h6A1: dout  = 8'b11111111; // 1697 : 255 - 0xff
      12'h6A2: dout  = 8'b11111111; // 1698 : 255 - 0xff
      12'h6A3: dout  = 8'b11111111; // 1699 : 255 - 0xff
      12'h6A4: dout  = 8'b11111111; // 1700 : 255 - 0xff
      12'h6A5: dout  = 8'b11111111; // 1701 : 255 - 0xff
      12'h6A6: dout  = 8'b11111111; // 1702 : 255 - 0xff
      12'h6A7: dout  = 8'b11111111; // 1703 : 255 - 0xff
      12'h6A8: dout  = 8'b11111111; // 1704 : 255 - 0xff -- Sprite 0xd5
      12'h6A9: dout  = 8'b11111111; // 1705 : 255 - 0xff
      12'h6AA: dout  = 8'b11111111; // 1706 : 255 - 0xff
      12'h6AB: dout  = 8'b11111111; // 1707 : 255 - 0xff
      12'h6AC: dout  = 8'b11111111; // 1708 : 255 - 0xff
      12'h6AD: dout  = 8'b11111111; // 1709 : 255 - 0xff
      12'h6AE: dout  = 8'b11111111; // 1710 : 255 - 0xff
      12'h6AF: dout  = 8'b11111111; // 1711 : 255 - 0xff
      12'h6B0: dout  = 8'b11111111; // 1712 : 255 - 0xff -- Sprite 0xd6
      12'h6B1: dout  = 8'b11111111; // 1713 : 255 - 0xff
      12'h6B2: dout  = 8'b11111111; // 1714 : 255 - 0xff
      12'h6B3: dout  = 8'b11111111; // 1715 : 255 - 0xff
      12'h6B4: dout  = 8'b11111111; // 1716 : 255 - 0xff
      12'h6B5: dout  = 8'b11111111; // 1717 : 255 - 0xff
      12'h6B6: dout  = 8'b11111111; // 1718 : 255 - 0xff
      12'h6B7: dout  = 8'b11111111; // 1719 : 255 - 0xff
      12'h6B8: dout  = 8'b11111111; // 1720 : 255 - 0xff -- Sprite 0xd7
      12'h6B9: dout  = 8'b11111111; // 1721 : 255 - 0xff
      12'h6BA: dout  = 8'b11111111; // 1722 : 255 - 0xff
      12'h6BB: dout  = 8'b11111111; // 1723 : 255 - 0xff
      12'h6BC: dout  = 8'b11111111; // 1724 : 255 - 0xff
      12'h6BD: dout  = 8'b11111111; // 1725 : 255 - 0xff
      12'h6BE: dout  = 8'b11111111; // 1726 : 255 - 0xff
      12'h6BF: dout  = 8'b11111111; // 1727 : 255 - 0xff
      12'h6C0: dout  = 8'b11111111; // 1728 : 255 - 0xff -- Sprite 0xd8
      12'h6C1: dout  = 8'b11111111; // 1729 : 255 - 0xff
      12'h6C2: dout  = 8'b11111111; // 1730 : 255 - 0xff
      12'h6C3: dout  = 8'b11111111; // 1731 : 255 - 0xff
      12'h6C4: dout  = 8'b11111111; // 1732 : 255 - 0xff
      12'h6C5: dout  = 8'b11111111; // 1733 : 255 - 0xff
      12'h6C6: dout  = 8'b11111111; // 1734 : 255 - 0xff
      12'h6C7: dout  = 8'b11111111; // 1735 : 255 - 0xff
      12'h6C8: dout  = 8'b11111111; // 1736 : 255 - 0xff -- Sprite 0xd9
      12'h6C9: dout  = 8'b11111111; // 1737 : 255 - 0xff
      12'h6CA: dout  = 8'b11111111; // 1738 : 255 - 0xff
      12'h6CB: dout  = 8'b11111111; // 1739 : 255 - 0xff
      12'h6CC: dout  = 8'b11111111; // 1740 : 255 - 0xff
      12'h6CD: dout  = 8'b11111111; // 1741 : 255 - 0xff
      12'h6CE: dout  = 8'b11111111; // 1742 : 255 - 0xff
      12'h6CF: dout  = 8'b11111111; // 1743 : 255 - 0xff
      12'h6D0: dout  = 8'b11111111; // 1744 : 255 - 0xff -- Sprite 0xda
      12'h6D1: dout  = 8'b11111111; // 1745 : 255 - 0xff
      12'h6D2: dout  = 8'b11111111; // 1746 : 255 - 0xff
      12'h6D3: dout  = 8'b11111111; // 1747 : 255 - 0xff
      12'h6D4: dout  = 8'b11111111; // 1748 : 255 - 0xff
      12'h6D5: dout  = 8'b11111111; // 1749 : 255 - 0xff
      12'h6D6: dout  = 8'b11111111; // 1750 : 255 - 0xff
      12'h6D7: dout  = 8'b11111111; // 1751 : 255 - 0xff
      12'h6D8: dout  = 8'b11111111; // 1752 : 255 - 0xff -- Sprite 0xdb
      12'h6D9: dout  = 8'b11111111; // 1753 : 255 - 0xff
      12'h6DA: dout  = 8'b11111111; // 1754 : 255 - 0xff
      12'h6DB: dout  = 8'b11111111; // 1755 : 255 - 0xff
      12'h6DC: dout  = 8'b11111111; // 1756 : 255 - 0xff
      12'h6DD: dout  = 8'b11111111; // 1757 : 255 - 0xff
      12'h6DE: dout  = 8'b11111111; // 1758 : 255 - 0xff
      12'h6DF: dout  = 8'b11111111; // 1759 : 255 - 0xff
      12'h6E0: dout  = 8'b11111111; // 1760 : 255 - 0xff -- Sprite 0xdc
      12'h6E1: dout  = 8'b11111111; // 1761 : 255 - 0xff
      12'h6E2: dout  = 8'b11111111; // 1762 : 255 - 0xff
      12'h6E3: dout  = 8'b11111111; // 1763 : 255 - 0xff
      12'h6E4: dout  = 8'b11111111; // 1764 : 255 - 0xff
      12'h6E5: dout  = 8'b11111111; // 1765 : 255 - 0xff
      12'h6E6: dout  = 8'b11111111; // 1766 : 255 - 0xff
      12'h6E7: dout  = 8'b11111111; // 1767 : 255 - 0xff
      12'h6E8: dout  = 8'b11111111; // 1768 : 255 - 0xff -- Sprite 0xdd
      12'h6E9: dout  = 8'b11111111; // 1769 : 255 - 0xff
      12'h6EA: dout  = 8'b11111111; // 1770 : 255 - 0xff
      12'h6EB: dout  = 8'b11111111; // 1771 : 255 - 0xff
      12'h6EC: dout  = 8'b11111111; // 1772 : 255 - 0xff
      12'h6ED: dout  = 8'b11111111; // 1773 : 255 - 0xff
      12'h6EE: dout  = 8'b11111111; // 1774 : 255 - 0xff
      12'h6EF: dout  = 8'b11111111; // 1775 : 255 - 0xff
      12'h6F0: dout  = 8'b11111111; // 1776 : 255 - 0xff -- Sprite 0xde
      12'h6F1: dout  = 8'b11111111; // 1777 : 255 - 0xff
      12'h6F2: dout  = 8'b11111111; // 1778 : 255 - 0xff
      12'h6F3: dout  = 8'b11111111; // 1779 : 255 - 0xff
      12'h6F4: dout  = 8'b11111111; // 1780 : 255 - 0xff
      12'h6F5: dout  = 8'b11111111; // 1781 : 255 - 0xff
      12'h6F6: dout  = 8'b11111111; // 1782 : 255 - 0xff
      12'h6F7: dout  = 8'b11111111; // 1783 : 255 - 0xff
      12'h6F8: dout  = 8'b11111111; // 1784 : 255 - 0xff -- Sprite 0xdf
      12'h6F9: dout  = 8'b11111111; // 1785 : 255 - 0xff
      12'h6FA: dout  = 8'b11111111; // 1786 : 255 - 0xff
      12'h6FB: dout  = 8'b11111111; // 1787 : 255 - 0xff
      12'h6FC: dout  = 8'b11111111; // 1788 : 255 - 0xff
      12'h6FD: dout  = 8'b11111111; // 1789 : 255 - 0xff
      12'h6FE: dout  = 8'b11111111; // 1790 : 255 - 0xff
      12'h6FF: dout  = 8'b11111111; // 1791 : 255 - 0xff
      12'h700: dout  = 8'b11111111; // 1792 : 255 - 0xff -- Sprite 0xe0
      12'h701: dout  = 8'b11111111; // 1793 : 255 - 0xff
      12'h702: dout  = 8'b11111111; // 1794 : 255 - 0xff
      12'h703: dout  = 8'b11111111; // 1795 : 255 - 0xff
      12'h704: dout  = 8'b11111111; // 1796 : 255 - 0xff
      12'h705: dout  = 8'b11111111; // 1797 : 255 - 0xff
      12'h706: dout  = 8'b11111111; // 1798 : 255 - 0xff
      12'h707: dout  = 8'b11111111; // 1799 : 255 - 0xff
      12'h708: dout  = 8'b11111111; // 1800 : 255 - 0xff -- Sprite 0xe1
      12'h709: dout  = 8'b11111111; // 1801 : 255 - 0xff
      12'h70A: dout  = 8'b11111111; // 1802 : 255 - 0xff
      12'h70B: dout  = 8'b11111111; // 1803 : 255 - 0xff
      12'h70C: dout  = 8'b11111111; // 1804 : 255 - 0xff
      12'h70D: dout  = 8'b11111111; // 1805 : 255 - 0xff
      12'h70E: dout  = 8'b11111111; // 1806 : 255 - 0xff
      12'h70F: dout  = 8'b11111111; // 1807 : 255 - 0xff
      12'h710: dout  = 8'b11111111; // 1808 : 255 - 0xff -- Sprite 0xe2
      12'h711: dout  = 8'b11111111; // 1809 : 255 - 0xff
      12'h712: dout  = 8'b11111111; // 1810 : 255 - 0xff
      12'h713: dout  = 8'b11111111; // 1811 : 255 - 0xff
      12'h714: dout  = 8'b11111111; // 1812 : 255 - 0xff
      12'h715: dout  = 8'b11111111; // 1813 : 255 - 0xff
      12'h716: dout  = 8'b11111111; // 1814 : 255 - 0xff
      12'h717: dout  = 8'b11111111; // 1815 : 255 - 0xff
      12'h718: dout  = 8'b11111111; // 1816 : 255 - 0xff -- Sprite 0xe3
      12'h719: dout  = 8'b11111111; // 1817 : 255 - 0xff
      12'h71A: dout  = 8'b11111111; // 1818 : 255 - 0xff
      12'h71B: dout  = 8'b11111111; // 1819 : 255 - 0xff
      12'h71C: dout  = 8'b11111111; // 1820 : 255 - 0xff
      12'h71D: dout  = 8'b11111111; // 1821 : 255 - 0xff
      12'h71E: dout  = 8'b11111111; // 1822 : 255 - 0xff
      12'h71F: dout  = 8'b11111111; // 1823 : 255 - 0xff
      12'h720: dout  = 8'b11111111; // 1824 : 255 - 0xff -- Sprite 0xe4
      12'h721: dout  = 8'b11111111; // 1825 : 255 - 0xff
      12'h722: dout  = 8'b11111111; // 1826 : 255 - 0xff
      12'h723: dout  = 8'b11111111; // 1827 : 255 - 0xff
      12'h724: dout  = 8'b11111111; // 1828 : 255 - 0xff
      12'h725: dout  = 8'b11111111; // 1829 : 255 - 0xff
      12'h726: dout  = 8'b11111111; // 1830 : 255 - 0xff
      12'h727: dout  = 8'b11111111; // 1831 : 255 - 0xff
      12'h728: dout  = 8'b11111111; // 1832 : 255 - 0xff -- Sprite 0xe5
      12'h729: dout  = 8'b11111111; // 1833 : 255 - 0xff
      12'h72A: dout  = 8'b11111111; // 1834 : 255 - 0xff
      12'h72B: dout  = 8'b11111111; // 1835 : 255 - 0xff
      12'h72C: dout  = 8'b11111111; // 1836 : 255 - 0xff
      12'h72D: dout  = 8'b11111111; // 1837 : 255 - 0xff
      12'h72E: dout  = 8'b11111111; // 1838 : 255 - 0xff
      12'h72F: dout  = 8'b11111111; // 1839 : 255 - 0xff
      12'h730: dout  = 8'b11111111; // 1840 : 255 - 0xff -- Sprite 0xe6
      12'h731: dout  = 8'b11111111; // 1841 : 255 - 0xff
      12'h732: dout  = 8'b11111111; // 1842 : 255 - 0xff
      12'h733: dout  = 8'b11111111; // 1843 : 255 - 0xff
      12'h734: dout  = 8'b11111111; // 1844 : 255 - 0xff
      12'h735: dout  = 8'b11111111; // 1845 : 255 - 0xff
      12'h736: dout  = 8'b11111111; // 1846 : 255 - 0xff
      12'h737: dout  = 8'b11111111; // 1847 : 255 - 0xff
      12'h738: dout  = 8'b11111111; // 1848 : 255 - 0xff -- Sprite 0xe7
      12'h739: dout  = 8'b11111111; // 1849 : 255 - 0xff
      12'h73A: dout  = 8'b11111111; // 1850 : 255 - 0xff
      12'h73B: dout  = 8'b11111111; // 1851 : 255 - 0xff
      12'h73C: dout  = 8'b11111111; // 1852 : 255 - 0xff
      12'h73D: dout  = 8'b11111111; // 1853 : 255 - 0xff
      12'h73E: dout  = 8'b11111111; // 1854 : 255 - 0xff
      12'h73F: dout  = 8'b11111111; // 1855 : 255 - 0xff
      12'h740: dout  = 8'b11111111; // 1856 : 255 - 0xff -- Sprite 0xe8
      12'h741: dout  = 8'b11111111; // 1857 : 255 - 0xff
      12'h742: dout  = 8'b11111111; // 1858 : 255 - 0xff
      12'h743: dout  = 8'b11111111; // 1859 : 255 - 0xff
      12'h744: dout  = 8'b11111111; // 1860 : 255 - 0xff
      12'h745: dout  = 8'b11111111; // 1861 : 255 - 0xff
      12'h746: dout  = 8'b11111111; // 1862 : 255 - 0xff
      12'h747: dout  = 8'b11111111; // 1863 : 255 - 0xff
      12'h748: dout  = 8'b11111111; // 1864 : 255 - 0xff -- Sprite 0xe9
      12'h749: dout  = 8'b11111111; // 1865 : 255 - 0xff
      12'h74A: dout  = 8'b11111111; // 1866 : 255 - 0xff
      12'h74B: dout  = 8'b11111111; // 1867 : 255 - 0xff
      12'h74C: dout  = 8'b11111111; // 1868 : 255 - 0xff
      12'h74D: dout  = 8'b11111111; // 1869 : 255 - 0xff
      12'h74E: dout  = 8'b11111111; // 1870 : 255 - 0xff
      12'h74F: dout  = 8'b11111111; // 1871 : 255 - 0xff
      12'h750: dout  = 8'b11111111; // 1872 : 255 - 0xff -- Sprite 0xea
      12'h751: dout  = 8'b11111111; // 1873 : 255 - 0xff
      12'h752: dout  = 8'b11111111; // 1874 : 255 - 0xff
      12'h753: dout  = 8'b11111111; // 1875 : 255 - 0xff
      12'h754: dout  = 8'b11111111; // 1876 : 255 - 0xff
      12'h755: dout  = 8'b11111111; // 1877 : 255 - 0xff
      12'h756: dout  = 8'b11111111; // 1878 : 255 - 0xff
      12'h757: dout  = 8'b11111111; // 1879 : 255 - 0xff
      12'h758: dout  = 8'b11111111; // 1880 : 255 - 0xff -- Sprite 0xeb
      12'h759: dout  = 8'b11111111; // 1881 : 255 - 0xff
      12'h75A: dout  = 8'b11111111; // 1882 : 255 - 0xff
      12'h75B: dout  = 8'b11111111; // 1883 : 255 - 0xff
      12'h75C: dout  = 8'b11111111; // 1884 : 255 - 0xff
      12'h75D: dout  = 8'b11111111; // 1885 : 255 - 0xff
      12'h75E: dout  = 8'b11111111; // 1886 : 255 - 0xff
      12'h75F: dout  = 8'b11111111; // 1887 : 255 - 0xff
      12'h760: dout  = 8'b11111111; // 1888 : 255 - 0xff -- Sprite 0xec
      12'h761: dout  = 8'b11111111; // 1889 : 255 - 0xff
      12'h762: dout  = 8'b11111111; // 1890 : 255 - 0xff
      12'h763: dout  = 8'b11111111; // 1891 : 255 - 0xff
      12'h764: dout  = 8'b11111111; // 1892 : 255 - 0xff
      12'h765: dout  = 8'b11111111; // 1893 : 255 - 0xff
      12'h766: dout  = 8'b11111111; // 1894 : 255 - 0xff
      12'h767: dout  = 8'b11111111; // 1895 : 255 - 0xff
      12'h768: dout  = 8'b11111111; // 1896 : 255 - 0xff -- Sprite 0xed
      12'h769: dout  = 8'b11111111; // 1897 : 255 - 0xff
      12'h76A: dout  = 8'b11111111; // 1898 : 255 - 0xff
      12'h76B: dout  = 8'b11111111; // 1899 : 255 - 0xff
      12'h76C: dout  = 8'b11111111; // 1900 : 255 - 0xff
      12'h76D: dout  = 8'b11111111; // 1901 : 255 - 0xff
      12'h76E: dout  = 8'b11111111; // 1902 : 255 - 0xff
      12'h76F: dout  = 8'b11111111; // 1903 : 255 - 0xff
      12'h770: dout  = 8'b11111111; // 1904 : 255 - 0xff -- Sprite 0xee
      12'h771: dout  = 8'b11111111; // 1905 : 255 - 0xff
      12'h772: dout  = 8'b11111111; // 1906 : 255 - 0xff
      12'h773: dout  = 8'b11111111; // 1907 : 255 - 0xff
      12'h774: dout  = 8'b11111111; // 1908 : 255 - 0xff
      12'h775: dout  = 8'b11111111; // 1909 : 255 - 0xff
      12'h776: dout  = 8'b11111111; // 1910 : 255 - 0xff
      12'h777: dout  = 8'b11111111; // 1911 : 255 - 0xff
      12'h778: dout  = 8'b11111111; // 1912 : 255 - 0xff -- Sprite 0xef
      12'h779: dout  = 8'b11111111; // 1913 : 255 - 0xff
      12'h77A: dout  = 8'b11111111; // 1914 : 255 - 0xff
      12'h77B: dout  = 8'b11111111; // 1915 : 255 - 0xff
      12'h77C: dout  = 8'b11111111; // 1916 : 255 - 0xff
      12'h77D: dout  = 8'b11111111; // 1917 : 255 - 0xff
      12'h77E: dout  = 8'b11111111; // 1918 : 255 - 0xff
      12'h77F: dout  = 8'b11111111; // 1919 : 255 - 0xff
      12'h780: dout  = 8'b11111111; // 1920 : 255 - 0xff -- Sprite 0xf0
      12'h781: dout  = 8'b11111111; // 1921 : 255 - 0xff
      12'h782: dout  = 8'b11111111; // 1922 : 255 - 0xff
      12'h783: dout  = 8'b11111111; // 1923 : 255 - 0xff
      12'h784: dout  = 8'b11111111; // 1924 : 255 - 0xff
      12'h785: dout  = 8'b11111111; // 1925 : 255 - 0xff
      12'h786: dout  = 8'b11111111; // 1926 : 255 - 0xff
      12'h787: dout  = 8'b11111111; // 1927 : 255 - 0xff
      12'h788: dout  = 8'b11111111; // 1928 : 255 - 0xff -- Sprite 0xf1
      12'h789: dout  = 8'b11111111; // 1929 : 255 - 0xff
      12'h78A: dout  = 8'b11111111; // 1930 : 255 - 0xff
      12'h78B: dout  = 8'b11111111; // 1931 : 255 - 0xff
      12'h78C: dout  = 8'b11111111; // 1932 : 255 - 0xff
      12'h78D: dout  = 8'b11111111; // 1933 : 255 - 0xff
      12'h78E: dout  = 8'b11111111; // 1934 : 255 - 0xff
      12'h78F: dout  = 8'b11111111; // 1935 : 255 - 0xff
      12'h790: dout  = 8'b11111111; // 1936 : 255 - 0xff -- Sprite 0xf2
      12'h791: dout  = 8'b11111111; // 1937 : 255 - 0xff
      12'h792: dout  = 8'b11111111; // 1938 : 255 - 0xff
      12'h793: dout  = 8'b11111111; // 1939 : 255 - 0xff
      12'h794: dout  = 8'b11111111; // 1940 : 255 - 0xff
      12'h795: dout  = 8'b11111111; // 1941 : 255 - 0xff
      12'h796: dout  = 8'b11111111; // 1942 : 255 - 0xff
      12'h797: dout  = 8'b11111111; // 1943 : 255 - 0xff
      12'h798: dout  = 8'b11111111; // 1944 : 255 - 0xff -- Sprite 0xf3
      12'h799: dout  = 8'b11111111; // 1945 : 255 - 0xff
      12'h79A: dout  = 8'b11111111; // 1946 : 255 - 0xff
      12'h79B: dout  = 8'b11111111; // 1947 : 255 - 0xff
      12'h79C: dout  = 8'b11111111; // 1948 : 255 - 0xff
      12'h79D: dout  = 8'b11111111; // 1949 : 255 - 0xff
      12'h79E: dout  = 8'b11111111; // 1950 : 255 - 0xff
      12'h79F: dout  = 8'b11111111; // 1951 : 255 - 0xff
      12'h7A0: dout  = 8'b11111111; // 1952 : 255 - 0xff -- Sprite 0xf4
      12'h7A1: dout  = 8'b11111111; // 1953 : 255 - 0xff
      12'h7A2: dout  = 8'b11111111; // 1954 : 255 - 0xff
      12'h7A3: dout  = 8'b11111111; // 1955 : 255 - 0xff
      12'h7A4: dout  = 8'b11111111; // 1956 : 255 - 0xff
      12'h7A5: dout  = 8'b11111111; // 1957 : 255 - 0xff
      12'h7A6: dout  = 8'b11111111; // 1958 : 255 - 0xff
      12'h7A7: dout  = 8'b11111111; // 1959 : 255 - 0xff
      12'h7A8: dout  = 8'b11111111; // 1960 : 255 - 0xff -- Sprite 0xf5
      12'h7A9: dout  = 8'b11111111; // 1961 : 255 - 0xff
      12'h7AA: dout  = 8'b11111111; // 1962 : 255 - 0xff
      12'h7AB: dout  = 8'b11111111; // 1963 : 255 - 0xff
      12'h7AC: dout  = 8'b11111111; // 1964 : 255 - 0xff
      12'h7AD: dout  = 8'b11111111; // 1965 : 255 - 0xff
      12'h7AE: dout  = 8'b11111111; // 1966 : 255 - 0xff
      12'h7AF: dout  = 8'b11111111; // 1967 : 255 - 0xff
      12'h7B0: dout  = 8'b11111111; // 1968 : 255 - 0xff -- Sprite 0xf6
      12'h7B1: dout  = 8'b11111111; // 1969 : 255 - 0xff
      12'h7B2: dout  = 8'b11111111; // 1970 : 255 - 0xff
      12'h7B3: dout  = 8'b11111111; // 1971 : 255 - 0xff
      12'h7B4: dout  = 8'b11111111; // 1972 : 255 - 0xff
      12'h7B5: dout  = 8'b11111111; // 1973 : 255 - 0xff
      12'h7B6: dout  = 8'b11111111; // 1974 : 255 - 0xff
      12'h7B7: dout  = 8'b11111111; // 1975 : 255 - 0xff
      12'h7B8: dout  = 8'b11111111; // 1976 : 255 - 0xff -- Sprite 0xf7
      12'h7B9: dout  = 8'b11111111; // 1977 : 255 - 0xff
      12'h7BA: dout  = 8'b11111111; // 1978 : 255 - 0xff
      12'h7BB: dout  = 8'b11111111; // 1979 : 255 - 0xff
      12'h7BC: dout  = 8'b11111111; // 1980 : 255 - 0xff
      12'h7BD: dout  = 8'b11111111; // 1981 : 255 - 0xff
      12'h7BE: dout  = 8'b11111111; // 1982 : 255 - 0xff
      12'h7BF: dout  = 8'b11111111; // 1983 : 255 - 0xff
      12'h7C0: dout  = 8'b11111111; // 1984 : 255 - 0xff -- Sprite 0xf8
      12'h7C1: dout  = 8'b11111111; // 1985 : 255 - 0xff
      12'h7C2: dout  = 8'b11111111; // 1986 : 255 - 0xff
      12'h7C3: dout  = 8'b11111111; // 1987 : 255 - 0xff
      12'h7C4: dout  = 8'b11111111; // 1988 : 255 - 0xff
      12'h7C5: dout  = 8'b11111111; // 1989 : 255 - 0xff
      12'h7C6: dout  = 8'b11111111; // 1990 : 255 - 0xff
      12'h7C7: dout  = 8'b11111111; // 1991 : 255 - 0xff
      12'h7C8: dout  = 8'b11111111; // 1992 : 255 - 0xff -- Sprite 0xf9
      12'h7C9: dout  = 8'b11111111; // 1993 : 255 - 0xff
      12'h7CA: dout  = 8'b11111111; // 1994 : 255 - 0xff
      12'h7CB: dout  = 8'b11111111; // 1995 : 255 - 0xff
      12'h7CC: dout  = 8'b11111111; // 1996 : 255 - 0xff
      12'h7CD: dout  = 8'b11111111; // 1997 : 255 - 0xff
      12'h7CE: dout  = 8'b11111111; // 1998 : 255 - 0xff
      12'h7CF: dout  = 8'b11111111; // 1999 : 255 - 0xff
      12'h7D0: dout  = 8'b11111111; // 2000 : 255 - 0xff -- Sprite 0xfa
      12'h7D1: dout  = 8'b11111111; // 2001 : 255 - 0xff
      12'h7D2: dout  = 8'b11111111; // 2002 : 255 - 0xff
      12'h7D3: dout  = 8'b11111111; // 2003 : 255 - 0xff
      12'h7D4: dout  = 8'b11111111; // 2004 : 255 - 0xff
      12'h7D5: dout  = 8'b11111111; // 2005 : 255 - 0xff
      12'h7D6: dout  = 8'b11111111; // 2006 : 255 - 0xff
      12'h7D7: dout  = 8'b11111111; // 2007 : 255 - 0xff
      12'h7D8: dout  = 8'b11111111; // 2008 : 255 - 0xff -- Sprite 0xfb
      12'h7D9: dout  = 8'b11111111; // 2009 : 255 - 0xff
      12'h7DA: dout  = 8'b11111111; // 2010 : 255 - 0xff
      12'h7DB: dout  = 8'b11111111; // 2011 : 255 - 0xff
      12'h7DC: dout  = 8'b11111111; // 2012 : 255 - 0xff
      12'h7DD: dout  = 8'b11111111; // 2013 : 255 - 0xff
      12'h7DE: dout  = 8'b11111111; // 2014 : 255 - 0xff
      12'h7DF: dout  = 8'b11111111; // 2015 : 255 - 0xff
      12'h7E0: dout  = 8'b11111111; // 2016 : 255 - 0xff -- Sprite 0xfc
      12'h7E1: dout  = 8'b11111111; // 2017 : 255 - 0xff
      12'h7E2: dout  = 8'b11111111; // 2018 : 255 - 0xff
      12'h7E3: dout  = 8'b11111111; // 2019 : 255 - 0xff
      12'h7E4: dout  = 8'b11111111; // 2020 : 255 - 0xff
      12'h7E5: dout  = 8'b11111111; // 2021 : 255 - 0xff
      12'h7E6: dout  = 8'b11111111; // 2022 : 255 - 0xff
      12'h7E7: dout  = 8'b11111111; // 2023 : 255 - 0xff
      12'h7E8: dout  = 8'b11111111; // 2024 : 255 - 0xff -- Sprite 0xfd
      12'h7E9: dout  = 8'b11111111; // 2025 : 255 - 0xff
      12'h7EA: dout  = 8'b11111111; // 2026 : 255 - 0xff
      12'h7EB: dout  = 8'b11111111; // 2027 : 255 - 0xff
      12'h7EC: dout  = 8'b11111111; // 2028 : 255 - 0xff
      12'h7ED: dout  = 8'b11111111; // 2029 : 255 - 0xff
      12'h7EE: dout  = 8'b11111111; // 2030 : 255 - 0xff
      12'h7EF: dout  = 8'b11111111; // 2031 : 255 - 0xff
      12'h7F0: dout  = 8'b11111111; // 2032 : 255 - 0xff -- Sprite 0xfe
      12'h7F1: dout  = 8'b11111111; // 2033 : 255 - 0xff
      12'h7F2: dout  = 8'b11111111; // 2034 : 255 - 0xff
      12'h7F3: dout  = 8'b11111111; // 2035 : 255 - 0xff
      12'h7F4: dout  = 8'b11111111; // 2036 : 255 - 0xff
      12'h7F5: dout  = 8'b11111111; // 2037 : 255 - 0xff
      12'h7F6: dout  = 8'b11111111; // 2038 : 255 - 0xff
      12'h7F7: dout  = 8'b11111111; // 2039 : 255 - 0xff
      12'h7F8: dout  = 8'b11111111; // 2040 : 255 - 0xff -- Sprite 0xff
      12'h7F9: dout  = 8'b11111111; // 2041 : 255 - 0xff
      12'h7FA: dout  = 8'b11111111; // 2042 : 255 - 0xff
      12'h7FB: dout  = 8'b11111111; // 2043 : 255 - 0xff
      12'h7FC: dout  = 8'b11111111; // 2044 : 255 - 0xff
      12'h7FD: dout  = 8'b11111111; // 2045 : 255 - 0xff
      12'h7FE: dout  = 8'b11111111; // 2046 : 255 - 0xff
      12'h7FF: dout  = 8'b11111111; // 2047 : 255 - 0xff
          // Background pattern Table
      12'h800: dout  = 8'b00000000; // 2048 :   0 - 0x0 -- Background 0x0
      12'h801: dout  = 8'b00000000; // 2049 :   0 - 0x0
      12'h802: dout  = 8'b00000000; // 2050 :   0 - 0x0
      12'h803: dout  = 8'b00000000; // 2051 :   0 - 0x0
      12'h804: dout  = 8'b00000000; // 2052 :   0 - 0x0
      12'h805: dout  = 8'b00000000; // 2053 :   0 - 0x0
      12'h806: dout  = 8'b00000000; // 2054 :   0 - 0x0
      12'h807: dout  = 8'b00000000; // 2055 :   0 - 0x0
      12'h808: dout  = 8'b00000000; // 2056 :   0 - 0x0 -- Background 0x1
      12'h809: dout  = 8'b00111000; // 2057 :  56 - 0x38
      12'h80A: dout  = 8'b01111100; // 2058 : 124 - 0x7c
      12'h80B: dout  = 8'b11111110; // 2059 : 254 - 0xfe
      12'h80C: dout  = 8'b11111110; // 2060 : 254 - 0xfe
      12'h80D: dout  = 8'b11111110; // 2061 : 254 - 0xfe
      12'h80E: dout  = 8'b01111100; // 2062 : 124 - 0x7c
      12'h80F: dout  = 8'b00111000; // 2063 :  56 - 0x38
      12'h810: dout  = 8'b00000000; // 2064 :   0 - 0x0 -- Background 0x2
      12'h811: dout  = 8'b00000000; // 2065 :   0 - 0x0
      12'h812: dout  = 8'b00000000; // 2066 :   0 - 0x0
      12'h813: dout  = 8'b00000000; // 2067 :   0 - 0x0
      12'h814: dout  = 8'b00000000; // 2068 :   0 - 0x0
      12'h815: dout  = 8'b00000000; // 2069 :   0 - 0x0
      12'h816: dout  = 8'b00000000; // 2070 :   0 - 0x0
      12'h817: dout  = 8'b00000000; // 2071 :   0 - 0x0
      12'h818: dout  = 8'b00000000; // 2072 :   0 - 0x0 -- Background 0x3
      12'h819: dout  = 8'b00000000; // 2073 :   0 - 0x0
      12'h81A: dout  = 8'b00000000; // 2074 :   0 - 0x0
      12'h81B: dout  = 8'b00011000; // 2075 :  24 - 0x18
      12'h81C: dout  = 8'b00011000; // 2076 :  24 - 0x18
      12'h81D: dout  = 8'b00000000; // 2077 :   0 - 0x0
      12'h81E: dout  = 8'b00000000; // 2078 :   0 - 0x0
      12'h81F: dout  = 8'b00000000; // 2079 :   0 - 0x0
      12'h820: dout  = 8'b11111111; // 2080 : 255 - 0xff -- Background 0x4
      12'h821: dout  = 8'b11111111; // 2081 : 255 - 0xff
      12'h822: dout  = 8'b11111111; // 2082 : 255 - 0xff
      12'h823: dout  = 8'b11111111; // 2083 : 255 - 0xff
      12'h824: dout  = 8'b11111111; // 2084 : 255 - 0xff
      12'h825: dout  = 8'b11111111; // 2085 : 255 - 0xff
      12'h826: dout  = 8'b11111111; // 2086 : 255 - 0xff
      12'h827: dout  = 8'b11111111; // 2087 : 255 - 0xff
      12'h828: dout  = 8'b00001111; // 2088 :  15 - 0xf -- Background 0x5
      12'h829: dout  = 8'b00001111; // 2089 :  15 - 0xf
      12'h82A: dout  = 8'b00001111; // 2090 :  15 - 0xf
      12'h82B: dout  = 8'b00001111; // 2091 :  15 - 0xf
      12'h82C: dout  = 8'b00001111; // 2092 :  15 - 0xf
      12'h82D: dout  = 8'b00001111; // 2093 :  15 - 0xf
      12'h82E: dout  = 8'b00001111; // 2094 :  15 - 0xf
      12'h82F: dout  = 8'b00001111; // 2095 :  15 - 0xf
      12'h830: dout  = 8'b11110000; // 2096 : 240 - 0xf0 -- Background 0x6
      12'h831: dout  = 8'b11110000; // 2097 : 240 - 0xf0
      12'h832: dout  = 8'b11110000; // 2098 : 240 - 0xf0
      12'h833: dout  = 8'b11110000; // 2099 : 240 - 0xf0
      12'h834: dout  = 8'b11110000; // 2100 : 240 - 0xf0
      12'h835: dout  = 8'b11110000; // 2101 : 240 - 0xf0
      12'h836: dout  = 8'b11110000; // 2102 : 240 - 0xf0
      12'h837: dout  = 8'b11110000; // 2103 : 240 - 0xf0
      12'h838: dout  = 8'b00000000; // 2104 :   0 - 0x0 -- Background 0x7
      12'h839: dout  = 8'b00000000; // 2105 :   0 - 0x0
      12'h83A: dout  = 8'b00000000; // 2106 :   0 - 0x0
      12'h83B: dout  = 8'b00000000; // 2107 :   0 - 0x0
      12'h83C: dout  = 8'b00000000; // 2108 :   0 - 0x0
      12'h83D: dout  = 8'b00000000; // 2109 :   0 - 0x0
      12'h83E: dout  = 8'b00000000; // 2110 :   0 - 0x0
      12'h83F: dout  = 8'b00000000; // 2111 :   0 - 0x0
      12'h840: dout  = 8'b00000000; // 2112 :   0 - 0x0 -- Background 0x8
      12'h841: dout  = 8'b00000000; // 2113 :   0 - 0x0
      12'h842: dout  = 8'b00000000; // 2114 :   0 - 0x0
      12'h843: dout  = 8'b00000000; // 2115 :   0 - 0x0
      12'h844: dout  = 8'b00000000; // 2116 :   0 - 0x0
      12'h845: dout  = 8'b00000000; // 2117 :   0 - 0x0
      12'h846: dout  = 8'b00000000; // 2118 :   0 - 0x0
      12'h847: dout  = 8'b00000000; // 2119 :   0 - 0x0
      12'h848: dout  = 8'b00000000; // 2120 :   0 - 0x0 -- Background 0x9
      12'h849: dout  = 8'b00000000; // 2121 :   0 - 0x0
      12'h84A: dout  = 8'b00000000; // 2122 :   0 - 0x0
      12'h84B: dout  = 8'b00011000; // 2123 :  24 - 0x18
      12'h84C: dout  = 8'b00011000; // 2124 :  24 - 0x18
      12'h84D: dout  = 8'b00000000; // 2125 :   0 - 0x0
      12'h84E: dout  = 8'b00000000; // 2126 :   0 - 0x0
      12'h84F: dout  = 8'b00000000; // 2127 :   0 - 0x0
      12'h850: dout  = 8'b00000000; // 2128 :   0 - 0x0 -- Background 0xa
      12'h851: dout  = 8'b00000000; // 2129 :   0 - 0x0
      12'h852: dout  = 8'b00000000; // 2130 :   0 - 0x0
      12'h853: dout  = 8'b00000000; // 2131 :   0 - 0x0
      12'h854: dout  = 8'b00000000; // 2132 :   0 - 0x0
      12'h855: dout  = 8'b00000000; // 2133 :   0 - 0x0
      12'h856: dout  = 8'b00000000; // 2134 :   0 - 0x0
      12'h857: dout  = 8'b00000000; // 2135 :   0 - 0x0
      12'h858: dout  = 8'b00000000; // 2136 :   0 - 0x0 -- Background 0xb
      12'h859: dout  = 8'b00000000; // 2137 :   0 - 0x0
      12'h85A: dout  = 8'b00000000; // 2138 :   0 - 0x0
      12'h85B: dout  = 8'b00000000; // 2139 :   0 - 0x0
      12'h85C: dout  = 8'b00000000; // 2140 :   0 - 0x0
      12'h85D: dout  = 8'b00000000; // 2141 :   0 - 0x0
      12'h85E: dout  = 8'b00000000; // 2142 :   0 - 0x0
      12'h85F: dout  = 8'b00000000; // 2143 :   0 - 0x0
      12'h860: dout  = 8'b00000000; // 2144 :   0 - 0x0 -- Background 0xc
      12'h861: dout  = 8'b00000000; // 2145 :   0 - 0x0
      12'h862: dout  = 8'b00000000; // 2146 :   0 - 0x0
      12'h863: dout  = 8'b00000000; // 2147 :   0 - 0x0
      12'h864: dout  = 8'b00000000; // 2148 :   0 - 0x0
      12'h865: dout  = 8'b00000000; // 2149 :   0 - 0x0
      12'h866: dout  = 8'b00000000; // 2150 :   0 - 0x0
      12'h867: dout  = 8'b00000000; // 2151 :   0 - 0x0
      12'h868: dout  = 8'b00000000; // 2152 :   0 - 0x0 -- Background 0xd
      12'h869: dout  = 8'b00000000; // 2153 :   0 - 0x0
      12'h86A: dout  = 8'b00000000; // 2154 :   0 - 0x0
      12'h86B: dout  = 8'b00000000; // 2155 :   0 - 0x0
      12'h86C: dout  = 8'b00000000; // 2156 :   0 - 0x0
      12'h86D: dout  = 8'b00000000; // 2157 :   0 - 0x0
      12'h86E: dout  = 8'b00000000; // 2158 :   0 - 0x0
      12'h86F: dout  = 8'b00000000; // 2159 :   0 - 0x0
      12'h870: dout  = 8'b00000000; // 2160 :   0 - 0x0 -- Background 0xe
      12'h871: dout  = 8'b00000000; // 2161 :   0 - 0x0
      12'h872: dout  = 8'b00000000; // 2162 :   0 - 0x0
      12'h873: dout  = 8'b00000000; // 2163 :   0 - 0x0
      12'h874: dout  = 8'b00000000; // 2164 :   0 - 0x0
      12'h875: dout  = 8'b00000000; // 2165 :   0 - 0x0
      12'h876: dout  = 8'b00000000; // 2166 :   0 - 0x0
      12'h877: dout  = 8'b00000000; // 2167 :   0 - 0x0
      12'h878: dout  = 8'b00000000; // 2168 :   0 - 0x0 -- Background 0xf
      12'h879: dout  = 8'b00000000; // 2169 :   0 - 0x0
      12'h87A: dout  = 8'b00000000; // 2170 :   0 - 0x0
      12'h87B: dout  = 8'b00000000; // 2171 :   0 - 0x0
      12'h87C: dout  = 8'b00000000; // 2172 :   0 - 0x0
      12'h87D: dout  = 8'b00000000; // 2173 :   0 - 0x0
      12'h87E: dout  = 8'b00000000; // 2174 :   0 - 0x0
      12'h87F: dout  = 8'b00000000; // 2175 :   0 - 0x0
      12'h880: dout  = 8'b00000000; // 2176 :   0 - 0x0 -- Background 0x10
      12'h881: dout  = 8'b00000000; // 2177 :   0 - 0x0
      12'h882: dout  = 8'b00000000; // 2178 :   0 - 0x0
      12'h883: dout  = 8'b00000000; // 2179 :   0 - 0x0
      12'h884: dout  = 8'b00000000; // 2180 :   0 - 0x0
      12'h885: dout  = 8'b00000000; // 2181 :   0 - 0x0
      12'h886: dout  = 8'b00000000; // 2182 :   0 - 0x0
      12'h887: dout  = 8'b00000000; // 2183 :   0 - 0x0
      12'h888: dout  = 8'b00000000; // 2184 :   0 - 0x0 -- Background 0x11
      12'h889: dout  = 8'b00000000; // 2185 :   0 - 0x0
      12'h88A: dout  = 8'b00000000; // 2186 :   0 - 0x0
      12'h88B: dout  = 8'b00000000; // 2187 :   0 - 0x0
      12'h88C: dout  = 8'b00000000; // 2188 :   0 - 0x0
      12'h88D: dout  = 8'b00000000; // 2189 :   0 - 0x0
      12'h88E: dout  = 8'b00000000; // 2190 :   0 - 0x0
      12'h88F: dout  = 8'b00000000; // 2191 :   0 - 0x0
      12'h890: dout  = 8'b00000000; // 2192 :   0 - 0x0 -- Background 0x12
      12'h891: dout  = 8'b00000000; // 2193 :   0 - 0x0
      12'h892: dout  = 8'b00000000; // 2194 :   0 - 0x0
      12'h893: dout  = 8'b00000000; // 2195 :   0 - 0x0
      12'h894: dout  = 8'b00000000; // 2196 :   0 - 0x0
      12'h895: dout  = 8'b00000000; // 2197 :   0 - 0x0
      12'h896: dout  = 8'b00000000; // 2198 :   0 - 0x0
      12'h897: dout  = 8'b00000000; // 2199 :   0 - 0x0
      12'h898: dout  = 8'b00000000; // 2200 :   0 - 0x0 -- Background 0x13
      12'h899: dout  = 8'b00000000; // 2201 :   0 - 0x0
      12'h89A: dout  = 8'b00000000; // 2202 :   0 - 0x0
      12'h89B: dout  = 8'b00000000; // 2203 :   0 - 0x0
      12'h89C: dout  = 8'b00000000; // 2204 :   0 - 0x0
      12'h89D: dout  = 8'b00000000; // 2205 :   0 - 0x0
      12'h89E: dout  = 8'b00000000; // 2206 :   0 - 0x0
      12'h89F: dout  = 8'b00000000; // 2207 :   0 - 0x0
      12'h8A0: dout  = 8'b00000000; // 2208 :   0 - 0x0 -- Background 0x14
      12'h8A1: dout  = 8'b00000000; // 2209 :   0 - 0x0
      12'h8A2: dout  = 8'b00000000; // 2210 :   0 - 0x0
      12'h8A3: dout  = 8'b00000000; // 2211 :   0 - 0x0
      12'h8A4: dout  = 8'b00000000; // 2212 :   0 - 0x0
      12'h8A5: dout  = 8'b00000000; // 2213 :   0 - 0x0
      12'h8A6: dout  = 8'b00000000; // 2214 :   0 - 0x0
      12'h8A7: dout  = 8'b00000000; // 2215 :   0 - 0x0
      12'h8A8: dout  = 8'b00000000; // 2216 :   0 - 0x0 -- Background 0x15
      12'h8A9: dout  = 8'b00000000; // 2217 :   0 - 0x0
      12'h8AA: dout  = 8'b00000000; // 2218 :   0 - 0x0
      12'h8AB: dout  = 8'b00000000; // 2219 :   0 - 0x0
      12'h8AC: dout  = 8'b00000000; // 2220 :   0 - 0x0
      12'h8AD: dout  = 8'b00000000; // 2221 :   0 - 0x0
      12'h8AE: dout  = 8'b00000000; // 2222 :   0 - 0x0
      12'h8AF: dout  = 8'b00000000; // 2223 :   0 - 0x0
      12'h8B0: dout  = 8'b00000000; // 2224 :   0 - 0x0 -- Background 0x16
      12'h8B1: dout  = 8'b00000000; // 2225 :   0 - 0x0
      12'h8B2: dout  = 8'b00000000; // 2226 :   0 - 0x0
      12'h8B3: dout  = 8'b00000000; // 2227 :   0 - 0x0
      12'h8B4: dout  = 8'b00000000; // 2228 :   0 - 0x0
      12'h8B5: dout  = 8'b00000000; // 2229 :   0 - 0x0
      12'h8B6: dout  = 8'b00000000; // 2230 :   0 - 0x0
      12'h8B7: dout  = 8'b00000000; // 2231 :   0 - 0x0
      12'h8B8: dout  = 8'b00000000; // 2232 :   0 - 0x0 -- Background 0x17
      12'h8B9: dout  = 8'b00000000; // 2233 :   0 - 0x0
      12'h8BA: dout  = 8'b00000000; // 2234 :   0 - 0x0
      12'h8BB: dout  = 8'b00000000; // 2235 :   0 - 0x0
      12'h8BC: dout  = 8'b00000000; // 2236 :   0 - 0x0
      12'h8BD: dout  = 8'b00000000; // 2237 :   0 - 0x0
      12'h8BE: dout  = 8'b00000000; // 2238 :   0 - 0x0
      12'h8BF: dout  = 8'b00000000; // 2239 :   0 - 0x0
      12'h8C0: dout  = 8'b00000000; // 2240 :   0 - 0x0 -- Background 0x18
      12'h8C1: dout  = 8'b00000000; // 2241 :   0 - 0x0
      12'h8C2: dout  = 8'b00000000; // 2242 :   0 - 0x0
      12'h8C3: dout  = 8'b00000000; // 2243 :   0 - 0x0
      12'h8C4: dout  = 8'b00000000; // 2244 :   0 - 0x0
      12'h8C5: dout  = 8'b00000000; // 2245 :   0 - 0x0
      12'h8C6: dout  = 8'b00000000; // 2246 :   0 - 0x0
      12'h8C7: dout  = 8'b00000000; // 2247 :   0 - 0x0
      12'h8C8: dout  = 8'b00000000; // 2248 :   0 - 0x0 -- Background 0x19
      12'h8C9: dout  = 8'b00000000; // 2249 :   0 - 0x0
      12'h8CA: dout  = 8'b00000000; // 2250 :   0 - 0x0
      12'h8CB: dout  = 8'b00000000; // 2251 :   0 - 0x0
      12'h8CC: dout  = 8'b00000000; // 2252 :   0 - 0x0
      12'h8CD: dout  = 8'b00000000; // 2253 :   0 - 0x0
      12'h8CE: dout  = 8'b00000000; // 2254 :   0 - 0x0
      12'h8CF: dout  = 8'b00000000; // 2255 :   0 - 0x0
      12'h8D0: dout  = 8'b00000000; // 2256 :   0 - 0x0 -- Background 0x1a
      12'h8D1: dout  = 8'b00000000; // 2257 :   0 - 0x0
      12'h8D2: dout  = 8'b00000000; // 2258 :   0 - 0x0
      12'h8D3: dout  = 8'b00000000; // 2259 :   0 - 0x0
      12'h8D4: dout  = 8'b00000000; // 2260 :   0 - 0x0
      12'h8D5: dout  = 8'b00000000; // 2261 :   0 - 0x0
      12'h8D6: dout  = 8'b00000000; // 2262 :   0 - 0x0
      12'h8D7: dout  = 8'b00000000; // 2263 :   0 - 0x0
      12'h8D8: dout  = 8'b00000000; // 2264 :   0 - 0x0 -- Background 0x1b
      12'h8D9: dout  = 8'b00000000; // 2265 :   0 - 0x0
      12'h8DA: dout  = 8'b00000000; // 2266 :   0 - 0x0
      12'h8DB: dout  = 8'b00000000; // 2267 :   0 - 0x0
      12'h8DC: dout  = 8'b00000000; // 2268 :   0 - 0x0
      12'h8DD: dout  = 8'b00000000; // 2269 :   0 - 0x0
      12'h8DE: dout  = 8'b00000000; // 2270 :   0 - 0x0
      12'h8DF: dout  = 8'b00000000; // 2271 :   0 - 0x0
      12'h8E0: dout  = 8'b00000000; // 2272 :   0 - 0x0 -- Background 0x1c
      12'h8E1: dout  = 8'b00000000; // 2273 :   0 - 0x0
      12'h8E2: dout  = 8'b00000000; // 2274 :   0 - 0x0
      12'h8E3: dout  = 8'b00000000; // 2275 :   0 - 0x0
      12'h8E4: dout  = 8'b00000000; // 2276 :   0 - 0x0
      12'h8E5: dout  = 8'b00000000; // 2277 :   0 - 0x0
      12'h8E6: dout  = 8'b00000000; // 2278 :   0 - 0x0
      12'h8E7: dout  = 8'b00000000; // 2279 :   0 - 0x0
      12'h8E8: dout  = 8'b00000000; // 2280 :   0 - 0x0 -- Background 0x1d
      12'h8E9: dout  = 8'b00000000; // 2281 :   0 - 0x0
      12'h8EA: dout  = 8'b00000000; // 2282 :   0 - 0x0
      12'h8EB: dout  = 8'b00000000; // 2283 :   0 - 0x0
      12'h8EC: dout  = 8'b00000000; // 2284 :   0 - 0x0
      12'h8ED: dout  = 8'b00000000; // 2285 :   0 - 0x0
      12'h8EE: dout  = 8'b00000000; // 2286 :   0 - 0x0
      12'h8EF: dout  = 8'b00000000; // 2287 :   0 - 0x0
      12'h8F0: dout  = 8'b00000000; // 2288 :   0 - 0x0 -- Background 0x1e
      12'h8F1: dout  = 8'b00000000; // 2289 :   0 - 0x0
      12'h8F2: dout  = 8'b00000000; // 2290 :   0 - 0x0
      12'h8F3: dout  = 8'b00000000; // 2291 :   0 - 0x0
      12'h8F4: dout  = 8'b00000000; // 2292 :   0 - 0x0
      12'h8F5: dout  = 8'b00000000; // 2293 :   0 - 0x0
      12'h8F6: dout  = 8'b00000000; // 2294 :   0 - 0x0
      12'h8F7: dout  = 8'b00000000; // 2295 :   0 - 0x0
      12'h8F8: dout  = 8'b00000000; // 2296 :   0 - 0x0 -- Background 0x1f
      12'h8F9: dout  = 8'b00000000; // 2297 :   0 - 0x0
      12'h8FA: dout  = 8'b00000000; // 2298 :   0 - 0x0
      12'h8FB: dout  = 8'b00000000; // 2299 :   0 - 0x0
      12'h8FC: dout  = 8'b00000000; // 2300 :   0 - 0x0
      12'h8FD: dout  = 8'b00000000; // 2301 :   0 - 0x0
      12'h8FE: dout  = 8'b00000000; // 2302 :   0 - 0x0
      12'h8FF: dout  = 8'b00000000; // 2303 :   0 - 0x0
      12'h900: dout  = 8'b00000000; // 2304 :   0 - 0x0 -- Background 0x20
      12'h901: dout  = 8'b00000000; // 2305 :   0 - 0x0
      12'h902: dout  = 8'b00000000; // 2306 :   0 - 0x0
      12'h903: dout  = 8'b00000000; // 2307 :   0 - 0x0
      12'h904: dout  = 8'b00000000; // 2308 :   0 - 0x0
      12'h905: dout  = 8'b00000000; // 2309 :   0 - 0x0
      12'h906: dout  = 8'b00000000; // 2310 :   0 - 0x0
      12'h907: dout  = 8'b00000000; // 2311 :   0 - 0x0
      12'h908: dout  = 8'b00001111; // 2312 :  15 - 0xf -- Background 0x21
      12'h909: dout  = 8'b00001111; // 2313 :  15 - 0xf
      12'h90A: dout  = 8'b00001111; // 2314 :  15 - 0xf
      12'h90B: dout  = 8'b00000111; // 2315 :   7 - 0x7
      12'h90C: dout  = 8'b00000111; // 2316 :   7 - 0x7
      12'h90D: dout  = 8'b00001111; // 2317 :  15 - 0xf
      12'h90E: dout  = 8'b00001111; // 2318 :  15 - 0xf
      12'h90F: dout  = 8'b00001111; // 2319 :  15 - 0xf
      12'h910: dout  = 8'b11110000; // 2320 : 240 - 0xf0 -- Background 0x22
      12'h911: dout  = 8'b11110000; // 2321 : 240 - 0xf0
      12'h912: dout  = 8'b11110000; // 2322 : 240 - 0xf0
      12'h913: dout  = 8'b11100000; // 2323 : 224 - 0xe0
      12'h914: dout  = 8'b11100000; // 2324 : 224 - 0xe0
      12'h915: dout  = 8'b11110000; // 2325 : 240 - 0xf0
      12'h916: dout  = 8'b11110000; // 2326 : 240 - 0xf0
      12'h917: dout  = 8'b11110000; // 2327 : 240 - 0xf0
      12'h918: dout  = 8'b11111111; // 2328 : 255 - 0xff -- Background 0x23
      12'h919: dout  = 8'b11111111; // 2329 : 255 - 0xff
      12'h91A: dout  = 8'b11100001; // 2330 : 225 - 0xe1
      12'h91B: dout  = 8'b11100001; // 2331 : 225 - 0xe1
      12'h91C: dout  = 8'b11100001; // 2332 : 225 - 0xe1
      12'h91D: dout  = 8'b11100001; // 2333 : 225 - 0xe1
      12'h91E: dout  = 8'b11100001; // 2334 : 225 - 0xe1
      12'h91F: dout  = 8'b11100001; // 2335 : 225 - 0xe1
      12'h920: dout  = 8'b10000111; // 2336 : 135 - 0x87 -- Background 0x24
      12'h921: dout  = 8'b11000111; // 2337 : 199 - 0xc7
      12'h922: dout  = 8'b11000000; // 2338 : 192 - 0xc0
      12'h923: dout  = 8'b11000111; // 2339 : 199 - 0xc7
      12'h924: dout  = 8'b11001111; // 2340 : 207 - 0xcf
      12'h925: dout  = 8'b11001110; // 2341 : 206 - 0xce
      12'h926: dout  = 8'b11001111; // 2342 : 207 - 0xcf
      12'h927: dout  = 8'b11000111; // 2343 : 199 - 0xc7
      12'h928: dout  = 8'b11111000; // 2344 : 248 - 0xf8 -- Background 0x25
      12'h929: dout  = 8'b11111100; // 2345 : 252 - 0xfc
      12'h92A: dout  = 8'b00011100; // 2346 :  28 - 0x1c
      12'h92B: dout  = 8'b11111100; // 2347 : 252 - 0xfc
      12'h92C: dout  = 8'b11111100; // 2348 : 252 - 0xfc
      12'h92D: dout  = 8'b00011100; // 2349 :  28 - 0x1c
      12'h92E: dout  = 8'b11111100; // 2350 : 252 - 0xfc
      12'h92F: dout  = 8'b11111100; // 2351 : 252 - 0xfc
      12'h930: dout  = 8'b11111111; // 2352 : 255 - 0xff -- Background 0x26
      12'h931: dout  = 8'b11111111; // 2353 : 255 - 0xff
      12'h932: dout  = 8'b11100111; // 2354 : 231 - 0xe7
      12'h933: dout  = 8'b11100111; // 2355 : 231 - 0xe7
      12'h934: dout  = 8'b11100111; // 2356 : 231 - 0xe7
      12'h935: dout  = 8'b11100111; // 2357 : 231 - 0xe7
      12'h936: dout  = 8'b11100111; // 2358 : 231 - 0xe7
      12'h937: dout  = 8'b11100111; // 2359 : 231 - 0xe7
      12'h938: dout  = 8'b11110000; // 2360 : 240 - 0xf0 -- Background 0x27
      12'h939: dout  = 8'b11111001; // 2361 : 249 - 0xf9
      12'h93A: dout  = 8'b00111001; // 2362 :  57 - 0x39
      12'h93B: dout  = 8'b00111001; // 2363 :  57 - 0x39
      12'h93C: dout  = 8'b00111001; // 2364 :  57 - 0x39
      12'h93D: dout  = 8'b00111001; // 2365 :  57 - 0x39
      12'h93E: dout  = 8'b00111001; // 2366 :  57 - 0x39
      12'h93F: dout  = 8'b00111000; // 2367 :  56 - 0x38
      12'h940: dout  = 8'b11111111; // 2368 : 255 - 0xff -- Background 0x28
      12'h941: dout  = 8'b11111111; // 2369 : 255 - 0xff
      12'h942: dout  = 8'b11000000; // 2370 : 192 - 0xc0
      12'h943: dout  = 8'b11000000; // 2371 : 192 - 0xc0
      12'h944: dout  = 8'b11000000; // 2372 : 192 - 0xc0
      12'h945: dout  = 8'b11000000; // 2373 : 192 - 0xc0
      12'h946: dout  = 8'b11111111; // 2374 : 255 - 0xff
      12'h947: dout  = 8'b11111111; // 2375 : 255 - 0xff
      12'h948: dout  = 8'b00011111; // 2376 :  31 - 0x1f -- Background 0x29
      12'h949: dout  = 8'b00111111; // 2377 :  63 - 0x3f
      12'h94A: dout  = 8'b00110000; // 2378 :  48 - 0x30
      12'h94B: dout  = 8'b00110000; // 2379 :  48 - 0x30
      12'h94C: dout  = 8'b00110000; // 2380 :  48 - 0x30
      12'h94D: dout  = 8'b00110000; // 2381 :  48 - 0x30
      12'h94E: dout  = 8'b00111111; // 2382 :  63 - 0x3f
      12'h94F: dout  = 8'b00011111; // 2383 :  31 - 0x1f
      12'h950: dout  = 8'b11100011; // 2384 : 227 - 0xe3 -- Background 0x2a
      12'h951: dout  = 8'b11110011; // 2385 : 243 - 0xf3
      12'h952: dout  = 8'b01110000; // 2386 : 112 - 0x70
      12'h953: dout  = 8'b01110000; // 2387 : 112 - 0x70
      12'h954: dout  = 8'b01110000; // 2388 : 112 - 0x70
      12'h955: dout  = 8'b01110000; // 2389 : 112 - 0x70
      12'h956: dout  = 8'b11110000; // 2390 : 240 - 0xf0
      12'h957: dout  = 8'b11100000; // 2391 : 224 - 0xe0
      12'h958: dout  = 8'b11111110; // 2392 : 254 - 0xfe -- Background 0x2b
      12'h959: dout  = 8'b11111110; // 2393 : 254 - 0xfe
      12'h95A: dout  = 8'b01110000; // 2394 : 112 - 0x70
      12'h95B: dout  = 8'b01110000; // 2395 : 112 - 0x70
      12'h95C: dout  = 8'b01110000; // 2396 : 112 - 0x70
      12'h95D: dout  = 8'b01110000; // 2397 : 112 - 0x70
      12'h95E: dout  = 8'b01110000; // 2398 : 112 - 0x70
      12'h95F: dout  = 8'b01110000; // 2399 : 112 - 0x70
      12'h960: dout  = 8'b00000000; // 2400 :   0 - 0x0 -- Background 0x2c
      12'h961: dout  = 8'b00000000; // 2401 :   0 - 0x0
      12'h962: dout  = 8'b00000000; // 2402 :   0 - 0x0
      12'h963: dout  = 8'b00000000; // 2403 :   0 - 0x0
      12'h964: dout  = 8'b00000000; // 2404 :   0 - 0x0
      12'h965: dout  = 8'b00000000; // 2405 :   0 - 0x0
      12'h966: dout  = 8'b00000000; // 2406 :   0 - 0x0
      12'h967: dout  = 8'b00000000; // 2407 :   0 - 0x0
      12'h968: dout  = 8'b11111111; // 2408 : 255 - 0xff -- Background 0x2d
      12'h969: dout  = 8'b11111111; // 2409 : 255 - 0xff
      12'h96A: dout  = 8'b11111111; // 2410 : 255 - 0xff
      12'h96B: dout  = 8'b11111111; // 2411 : 255 - 0xff
      12'h96C: dout  = 8'b11111111; // 2412 : 255 - 0xff
      12'h96D: dout  = 8'b11111111; // 2413 : 255 - 0xff
      12'h96E: dout  = 8'b11111111; // 2414 : 255 - 0xff
      12'h96F: dout  = 8'b11111111; // 2415 : 255 - 0xff
      12'h970: dout  = 8'b00000000; // 2416 :   0 - 0x0 -- Background 0x2e
      12'h971: dout  = 8'b00000000; // 2417 :   0 - 0x0
      12'h972: dout  = 8'b00000000; // 2418 :   0 - 0x0
      12'h973: dout  = 8'b00000000; // 2419 :   0 - 0x0
      12'h974: dout  = 8'b00000000; // 2420 :   0 - 0x0
      12'h975: dout  = 8'b00000000; // 2421 :   0 - 0x0
      12'h976: dout  = 8'b00000000; // 2422 :   0 - 0x0
      12'h977: dout  = 8'b00000000; // 2423 :   0 - 0x0
      12'h978: dout  = 8'b00000000; // 2424 :   0 - 0x0 -- Background 0x2f
      12'h979: dout  = 8'b00000000; // 2425 :   0 - 0x0
      12'h97A: dout  = 8'b00000000; // 2426 :   0 - 0x0
      12'h97B: dout  = 8'b00011000; // 2427 :  24 - 0x18
      12'h97C: dout  = 8'b00011000; // 2428 :  24 - 0x18
      12'h97D: dout  = 8'b00000000; // 2429 :   0 - 0x0
      12'h97E: dout  = 8'b00000000; // 2430 :   0 - 0x0
      12'h97F: dout  = 8'b00000000; // 2431 :   0 - 0x0
      12'h980: dout  = 8'b00000000; // 2432 :   0 - 0x0 -- Background 0x30
      12'h981: dout  = 8'b00000000; // 2433 :   0 - 0x0
      12'h982: dout  = 8'b00000000; // 2434 :   0 - 0x0
      12'h983: dout  = 8'b00000000; // 2435 :   0 - 0x0
      12'h984: dout  = 8'b00000000; // 2436 :   0 - 0x0
      12'h985: dout  = 8'b00000000; // 2437 :   0 - 0x0
      12'h986: dout  = 8'b00000000; // 2438 :   0 - 0x0
      12'h987: dout  = 8'b00000000; // 2439 :   0 - 0x0
      12'h988: dout  = 8'b00000000; // 2440 :   0 - 0x0 -- Background 0x31
      12'h989: dout  = 8'b00000000; // 2441 :   0 - 0x0
      12'h98A: dout  = 8'b00000000; // 2442 :   0 - 0x0
      12'h98B: dout  = 8'b00000000; // 2443 :   0 - 0x0
      12'h98C: dout  = 8'b00000000; // 2444 :   0 - 0x0
      12'h98D: dout  = 8'b00000000; // 2445 :   0 - 0x0
      12'h98E: dout  = 8'b00000000; // 2446 :   0 - 0x0
      12'h98F: dout  = 8'b00000000; // 2447 :   0 - 0x0
      12'h990: dout  = 8'b00000000; // 2448 :   0 - 0x0 -- Background 0x32
      12'h991: dout  = 8'b00000000; // 2449 :   0 - 0x0
      12'h992: dout  = 8'b00000000; // 2450 :   0 - 0x0
      12'h993: dout  = 8'b00000000; // 2451 :   0 - 0x0
      12'h994: dout  = 8'b00000000; // 2452 :   0 - 0x0
      12'h995: dout  = 8'b00000000; // 2453 :   0 - 0x0
      12'h996: dout  = 8'b00000000; // 2454 :   0 - 0x0
      12'h997: dout  = 8'b00000000; // 2455 :   0 - 0x0
      12'h998: dout  = 8'b00000000; // 2456 :   0 - 0x0 -- Background 0x33
      12'h999: dout  = 8'b00000000; // 2457 :   0 - 0x0
      12'h99A: dout  = 8'b00000000; // 2458 :   0 - 0x0
      12'h99B: dout  = 8'b00000000; // 2459 :   0 - 0x0
      12'h99C: dout  = 8'b00000000; // 2460 :   0 - 0x0
      12'h99D: dout  = 8'b00000000; // 2461 :   0 - 0x0
      12'h99E: dout  = 8'b00000000; // 2462 :   0 - 0x0
      12'h99F: dout  = 8'b00000000; // 2463 :   0 - 0x0
      12'h9A0: dout  = 8'b00000000; // 2464 :   0 - 0x0 -- Background 0x34
      12'h9A1: dout  = 8'b00000000; // 2465 :   0 - 0x0
      12'h9A2: dout  = 8'b00000000; // 2466 :   0 - 0x0
      12'h9A3: dout  = 8'b00000000; // 2467 :   0 - 0x0
      12'h9A4: dout  = 8'b00000000; // 2468 :   0 - 0x0
      12'h9A5: dout  = 8'b00000000; // 2469 :   0 - 0x0
      12'h9A6: dout  = 8'b00000000; // 2470 :   0 - 0x0
      12'h9A7: dout  = 8'b00000000; // 2471 :   0 - 0x0
      12'h9A8: dout  = 8'b00000000; // 2472 :   0 - 0x0 -- Background 0x35
      12'h9A9: dout  = 8'b00000000; // 2473 :   0 - 0x0
      12'h9AA: dout  = 8'b00000000; // 2474 :   0 - 0x0
      12'h9AB: dout  = 8'b00000000; // 2475 :   0 - 0x0
      12'h9AC: dout  = 8'b00000000; // 2476 :   0 - 0x0
      12'h9AD: dout  = 8'b00000000; // 2477 :   0 - 0x0
      12'h9AE: dout  = 8'b00000000; // 2478 :   0 - 0x0
      12'h9AF: dout  = 8'b00000000; // 2479 :   0 - 0x0
      12'h9B0: dout  = 8'b00000000; // 2480 :   0 - 0x0 -- Background 0x36
      12'h9B1: dout  = 8'b00000000; // 2481 :   0 - 0x0
      12'h9B2: dout  = 8'b00000000; // 2482 :   0 - 0x0
      12'h9B3: dout  = 8'b00000000; // 2483 :   0 - 0x0
      12'h9B4: dout  = 8'b00000000; // 2484 :   0 - 0x0
      12'h9B5: dout  = 8'b00000000; // 2485 :   0 - 0x0
      12'h9B6: dout  = 8'b00000000; // 2486 :   0 - 0x0
      12'h9B7: dout  = 8'b00000000; // 2487 :   0 - 0x0
      12'h9B8: dout  = 8'b00000000; // 2488 :   0 - 0x0 -- Background 0x37
      12'h9B9: dout  = 8'b00000000; // 2489 :   0 - 0x0
      12'h9BA: dout  = 8'b00000000; // 2490 :   0 - 0x0
      12'h9BB: dout  = 8'b00000000; // 2491 :   0 - 0x0
      12'h9BC: dout  = 8'b00000000; // 2492 :   0 - 0x0
      12'h9BD: dout  = 8'b00000000; // 2493 :   0 - 0x0
      12'h9BE: dout  = 8'b00000000; // 2494 :   0 - 0x0
      12'h9BF: dout  = 8'b00000000; // 2495 :   0 - 0x0
      12'h9C0: dout  = 8'b00000000; // 2496 :   0 - 0x0 -- Background 0x38
      12'h9C1: dout  = 8'b00000000; // 2497 :   0 - 0x0
      12'h9C2: dout  = 8'b00000000; // 2498 :   0 - 0x0
      12'h9C3: dout  = 8'b00000000; // 2499 :   0 - 0x0
      12'h9C4: dout  = 8'b00000000; // 2500 :   0 - 0x0
      12'h9C5: dout  = 8'b00000000; // 2501 :   0 - 0x0
      12'h9C6: dout  = 8'b00000000; // 2502 :   0 - 0x0
      12'h9C7: dout  = 8'b00000000; // 2503 :   0 - 0x0
      12'h9C8: dout  = 8'b00000000; // 2504 :   0 - 0x0 -- Background 0x39
      12'h9C9: dout  = 8'b00000000; // 2505 :   0 - 0x0
      12'h9CA: dout  = 8'b00000000; // 2506 :   0 - 0x0
      12'h9CB: dout  = 8'b00000000; // 2507 :   0 - 0x0
      12'h9CC: dout  = 8'b00000000; // 2508 :   0 - 0x0
      12'h9CD: dout  = 8'b00000000; // 2509 :   0 - 0x0
      12'h9CE: dout  = 8'b00000000; // 2510 :   0 - 0x0
      12'h9CF: dout  = 8'b00000000; // 2511 :   0 - 0x0
      12'h9D0: dout  = 8'b00000000; // 2512 :   0 - 0x0 -- Background 0x3a
      12'h9D1: dout  = 8'b00000000; // 2513 :   0 - 0x0
      12'h9D2: dout  = 8'b00000000; // 2514 :   0 - 0x0
      12'h9D3: dout  = 8'b00000000; // 2515 :   0 - 0x0
      12'h9D4: dout  = 8'b00000000; // 2516 :   0 - 0x0
      12'h9D5: dout  = 8'b00000000; // 2517 :   0 - 0x0
      12'h9D6: dout  = 8'b00000000; // 2518 :   0 - 0x0
      12'h9D7: dout  = 8'b00000000; // 2519 :   0 - 0x0
      12'h9D8: dout  = 8'b00000000; // 2520 :   0 - 0x0 -- Background 0x3b
      12'h9D9: dout  = 8'b00000000; // 2521 :   0 - 0x0
      12'h9DA: dout  = 8'b00000000; // 2522 :   0 - 0x0
      12'h9DB: dout  = 8'b00000000; // 2523 :   0 - 0x0
      12'h9DC: dout  = 8'b00000000; // 2524 :   0 - 0x0
      12'h9DD: dout  = 8'b00000000; // 2525 :   0 - 0x0
      12'h9DE: dout  = 8'b00000000; // 2526 :   0 - 0x0
      12'h9DF: dout  = 8'b00000000; // 2527 :   0 - 0x0
      12'h9E0: dout  = 8'b00000000; // 2528 :   0 - 0x0 -- Background 0x3c
      12'h9E1: dout  = 8'b00000111; // 2529 :   7 - 0x7
      12'h9E2: dout  = 8'b00011111; // 2530 :  31 - 0x1f
      12'h9E3: dout  = 8'b00111111; // 2531 :  63 - 0x3f
      12'h9E4: dout  = 8'b00111111; // 2532 :  63 - 0x3f
      12'h9E5: dout  = 8'b00001111; // 2533 :  15 - 0xf
      12'h9E6: dout  = 8'b00000011; // 2534 :   3 - 0x3
      12'h9E7: dout  = 8'b00000000; // 2535 :   0 - 0x0
      12'h9E8: dout  = 8'b00000000; // 2536 :   0 - 0x0 -- Background 0x3d
      12'h9E9: dout  = 8'b11000000; // 2537 : 192 - 0xc0
      12'h9EA: dout  = 8'b11110000; // 2538 : 240 - 0xf0
      12'h9EB: dout  = 8'b11111000; // 2539 : 248 - 0xf8
      12'h9EC: dout  = 8'b11111000; // 2540 : 248 - 0xf8
      12'h9ED: dout  = 8'b11111100; // 2541 : 252 - 0xfc
      12'h9EE: dout  = 8'b11111100; // 2542 : 252 - 0xfc
      12'h9EF: dout  = 8'b11111100; // 2543 : 252 - 0xfc
      12'h9F0: dout  = 8'b00000000; // 2544 :   0 - 0x0 -- Background 0x3e
      12'h9F1: dout  = 8'b00000011; // 2545 :   3 - 0x3
      12'h9F2: dout  = 8'b00001111; // 2546 :  15 - 0xf
      12'h9F3: dout  = 8'b00111111; // 2547 :  63 - 0x3f
      12'h9F4: dout  = 8'b00111111; // 2548 :  63 - 0x3f
      12'h9F5: dout  = 8'b00011111; // 2549 :  31 - 0x1f
      12'h9F6: dout  = 8'b00000111; // 2550 :   7 - 0x7
      12'h9F7: dout  = 8'b00000000; // 2551 :   0 - 0x0
      12'h9F8: dout  = 8'b11111100; // 2552 : 252 - 0xfc -- Background 0x3f
      12'h9F9: dout  = 8'b11111100; // 2553 : 252 - 0xfc
      12'h9FA: dout  = 8'b11111100; // 2554 : 252 - 0xfc
      12'h9FB: dout  = 8'b11111000; // 2555 : 248 - 0xf8
      12'h9FC: dout  = 8'b11111000; // 2556 : 248 - 0xf8
      12'h9FD: dout  = 8'b11110000; // 2557 : 240 - 0xf0
      12'h9FE: dout  = 8'b11000000; // 2558 : 192 - 0xc0
      12'h9FF: dout  = 8'b00000000; // 2559 :   0 - 0x0
      12'hA00: dout  = 8'b00000000; // 2560 :   0 - 0x0 -- Background 0x40
      12'hA01: dout  = 8'b00000000; // 2561 :   0 - 0x0
      12'hA02: dout  = 8'b00000000; // 2562 :   0 - 0x0
      12'hA03: dout  = 8'b00000000; // 2563 :   0 - 0x0
      12'hA04: dout  = 8'b00000000; // 2564 :   0 - 0x0
      12'hA05: dout  = 8'b00000000; // 2565 :   0 - 0x0
      12'hA06: dout  = 8'b00000000; // 2566 :   0 - 0x0
      12'hA07: dout  = 8'b00000000; // 2567 :   0 - 0x0
      12'hA08: dout  = 8'b00000000; // 2568 :   0 - 0x0 -- Background 0x41
      12'hA09: dout  = 8'b00000000; // 2569 :   0 - 0x0
      12'hA0A: dout  = 8'b00000000; // 2570 :   0 - 0x0
      12'hA0B: dout  = 8'b00000000; // 2571 :   0 - 0x0
      12'hA0C: dout  = 8'b00000000; // 2572 :   0 - 0x0
      12'hA0D: dout  = 8'b00000000; // 2573 :   0 - 0x0
      12'hA0E: dout  = 8'b00000000; // 2574 :   0 - 0x0
      12'hA0F: dout  = 8'b00000000; // 2575 :   0 - 0x0
      12'hA10: dout  = 8'b00000000; // 2576 :   0 - 0x0 -- Background 0x42
      12'hA11: dout  = 8'b00000000; // 2577 :   0 - 0x0
      12'hA12: dout  = 8'b00000000; // 2578 :   0 - 0x0
      12'hA13: dout  = 8'b00000000; // 2579 :   0 - 0x0
      12'hA14: dout  = 8'b00000000; // 2580 :   0 - 0x0
      12'hA15: dout  = 8'b00000000; // 2581 :   0 - 0x0
      12'hA16: dout  = 8'b00000000; // 2582 :   0 - 0x0
      12'hA17: dout  = 8'b00000000; // 2583 :   0 - 0x0
      12'hA18: dout  = 8'b00000000; // 2584 :   0 - 0x0 -- Background 0x43
      12'hA19: dout  = 8'b00000000; // 2585 :   0 - 0x0
      12'hA1A: dout  = 8'b00000000; // 2586 :   0 - 0x0
      12'hA1B: dout  = 8'b00000000; // 2587 :   0 - 0x0
      12'hA1C: dout  = 8'b00000000; // 2588 :   0 - 0x0
      12'hA1D: dout  = 8'b00000000; // 2589 :   0 - 0x0
      12'hA1E: dout  = 8'b00000000; // 2590 :   0 - 0x0
      12'hA1F: dout  = 8'b00000000; // 2591 :   0 - 0x0
      12'hA20: dout  = 8'b00000000; // 2592 :   0 - 0x0 -- Background 0x44
      12'hA21: dout  = 8'b00000000; // 2593 :   0 - 0x0
      12'hA22: dout  = 8'b00000000; // 2594 :   0 - 0x0
      12'hA23: dout  = 8'b00000000; // 2595 :   0 - 0x0
      12'hA24: dout  = 8'b00000000; // 2596 :   0 - 0x0
      12'hA25: dout  = 8'b00000000; // 2597 :   0 - 0x0
      12'hA26: dout  = 8'b00000000; // 2598 :   0 - 0x0
      12'hA27: dout  = 8'b00000000; // 2599 :   0 - 0x0
      12'hA28: dout  = 8'b00000000; // 2600 :   0 - 0x0 -- Background 0x45
      12'hA29: dout  = 8'b00000000; // 2601 :   0 - 0x0
      12'hA2A: dout  = 8'b00000000; // 2602 :   0 - 0x0
      12'hA2B: dout  = 8'b00000000; // 2603 :   0 - 0x0
      12'hA2C: dout  = 8'b00000000; // 2604 :   0 - 0x0
      12'hA2D: dout  = 8'b00000000; // 2605 :   0 - 0x0
      12'hA2E: dout  = 8'b00000000; // 2606 :   0 - 0x0
      12'hA2F: dout  = 8'b00000000; // 2607 :   0 - 0x0
      12'hA30: dout  = 8'b00000000; // 2608 :   0 - 0x0 -- Background 0x46
      12'hA31: dout  = 8'b00000000; // 2609 :   0 - 0x0
      12'hA32: dout  = 8'b00000000; // 2610 :   0 - 0x0
      12'hA33: dout  = 8'b00000000; // 2611 :   0 - 0x0
      12'hA34: dout  = 8'b00000000; // 2612 :   0 - 0x0
      12'hA35: dout  = 8'b00000000; // 2613 :   0 - 0x0
      12'hA36: dout  = 8'b00000000; // 2614 :   0 - 0x0
      12'hA37: dout  = 8'b00000000; // 2615 :   0 - 0x0
      12'hA38: dout  = 8'b00000000; // 2616 :   0 - 0x0 -- Background 0x47
      12'hA39: dout  = 8'b00000000; // 2617 :   0 - 0x0
      12'hA3A: dout  = 8'b00000000; // 2618 :   0 - 0x0
      12'hA3B: dout  = 8'b00000000; // 2619 :   0 - 0x0
      12'hA3C: dout  = 8'b00000000; // 2620 :   0 - 0x0
      12'hA3D: dout  = 8'b00000000; // 2621 :   0 - 0x0
      12'hA3E: dout  = 8'b00000000; // 2622 :   0 - 0x0
      12'hA3F: dout  = 8'b00000000; // 2623 :   0 - 0x0
      12'hA40: dout  = 8'b00000000; // 2624 :   0 - 0x0 -- Background 0x48
      12'hA41: dout  = 8'b00000000; // 2625 :   0 - 0x0
      12'hA42: dout  = 8'b00000000; // 2626 :   0 - 0x0
      12'hA43: dout  = 8'b00000000; // 2627 :   0 - 0x0
      12'hA44: dout  = 8'b00000000; // 2628 :   0 - 0x0
      12'hA45: dout  = 8'b00000000; // 2629 :   0 - 0x0
      12'hA46: dout  = 8'b00000000; // 2630 :   0 - 0x0
      12'hA47: dout  = 8'b00000000; // 2631 :   0 - 0x0
      12'hA48: dout  = 8'b00000000; // 2632 :   0 - 0x0 -- Background 0x49
      12'hA49: dout  = 8'b00000000; // 2633 :   0 - 0x0
      12'hA4A: dout  = 8'b00000000; // 2634 :   0 - 0x0
      12'hA4B: dout  = 8'b00000000; // 2635 :   0 - 0x0
      12'hA4C: dout  = 8'b00000000; // 2636 :   0 - 0x0
      12'hA4D: dout  = 8'b00000000; // 2637 :   0 - 0x0
      12'hA4E: dout  = 8'b00000000; // 2638 :   0 - 0x0
      12'hA4F: dout  = 8'b00000000; // 2639 :   0 - 0x0
      12'hA50: dout  = 8'b00000000; // 2640 :   0 - 0x0 -- Background 0x4a
      12'hA51: dout  = 8'b00000000; // 2641 :   0 - 0x0
      12'hA52: dout  = 8'b00000000; // 2642 :   0 - 0x0
      12'hA53: dout  = 8'b00000000; // 2643 :   0 - 0x0
      12'hA54: dout  = 8'b00000000; // 2644 :   0 - 0x0
      12'hA55: dout  = 8'b00000000; // 2645 :   0 - 0x0
      12'hA56: dout  = 8'b00000000; // 2646 :   0 - 0x0
      12'hA57: dout  = 8'b00000000; // 2647 :   0 - 0x0
      12'hA58: dout  = 8'b00000000; // 2648 :   0 - 0x0 -- Background 0x4b
      12'hA59: dout  = 8'b00000000; // 2649 :   0 - 0x0
      12'hA5A: dout  = 8'b00000000; // 2650 :   0 - 0x0
      12'hA5B: dout  = 8'b00000000; // 2651 :   0 - 0x0
      12'hA5C: dout  = 8'b00000000; // 2652 :   0 - 0x0
      12'hA5D: dout  = 8'b00000000; // 2653 :   0 - 0x0
      12'hA5E: dout  = 8'b00000000; // 2654 :   0 - 0x0
      12'hA5F: dout  = 8'b00000000; // 2655 :   0 - 0x0
      12'hA60: dout  = 8'b00000000; // 2656 :   0 - 0x0 -- Background 0x4c
      12'hA61: dout  = 8'b00000000; // 2657 :   0 - 0x0
      12'hA62: dout  = 8'b00000000; // 2658 :   0 - 0x0
      12'hA63: dout  = 8'b00000000; // 2659 :   0 - 0x0
      12'hA64: dout  = 8'b00000000; // 2660 :   0 - 0x0
      12'hA65: dout  = 8'b00000000; // 2661 :   0 - 0x0
      12'hA66: dout  = 8'b00000000; // 2662 :   0 - 0x0
      12'hA67: dout  = 8'b00000000; // 2663 :   0 - 0x0
      12'hA68: dout  = 8'b00000000; // 2664 :   0 - 0x0 -- Background 0x4d
      12'hA69: dout  = 8'b00000000; // 2665 :   0 - 0x0
      12'hA6A: dout  = 8'b00000000; // 2666 :   0 - 0x0
      12'hA6B: dout  = 8'b00000000; // 2667 :   0 - 0x0
      12'hA6C: dout  = 8'b00000000; // 2668 :   0 - 0x0
      12'hA6D: dout  = 8'b00000000; // 2669 :   0 - 0x0
      12'hA6E: dout  = 8'b00000000; // 2670 :   0 - 0x0
      12'hA6F: dout  = 8'b00000000; // 2671 :   0 - 0x0
      12'hA70: dout  = 8'b00000000; // 2672 :   0 - 0x0 -- Background 0x4e
      12'hA71: dout  = 8'b00000000; // 2673 :   0 - 0x0
      12'hA72: dout  = 8'b00000000; // 2674 :   0 - 0x0
      12'hA73: dout  = 8'b00000000; // 2675 :   0 - 0x0
      12'hA74: dout  = 8'b00000000; // 2676 :   0 - 0x0
      12'hA75: dout  = 8'b00000000; // 2677 :   0 - 0x0
      12'hA76: dout  = 8'b00000000; // 2678 :   0 - 0x0
      12'hA77: dout  = 8'b00000000; // 2679 :   0 - 0x0
      12'hA78: dout  = 8'b00000000; // 2680 :   0 - 0x0 -- Background 0x4f
      12'hA79: dout  = 8'b00000000; // 2681 :   0 - 0x0
      12'hA7A: dout  = 8'b00000000; // 2682 :   0 - 0x0
      12'hA7B: dout  = 8'b00000000; // 2683 :   0 - 0x0
      12'hA7C: dout  = 8'b00000000; // 2684 :   0 - 0x0
      12'hA7D: dout  = 8'b00000000; // 2685 :   0 - 0x0
      12'hA7E: dout  = 8'b00000000; // 2686 :   0 - 0x0
      12'hA7F: dout  = 8'b00000000; // 2687 :   0 - 0x0
      12'hA80: dout  = 8'b00000000; // 2688 :   0 - 0x0 -- Background 0x50
      12'hA81: dout  = 8'b00000000; // 2689 :   0 - 0x0
      12'hA82: dout  = 8'b00000000; // 2690 :   0 - 0x0
      12'hA83: dout  = 8'b00000000; // 2691 :   0 - 0x0
      12'hA84: dout  = 8'b00000000; // 2692 :   0 - 0x0
      12'hA85: dout  = 8'b00000000; // 2693 :   0 - 0x0
      12'hA86: dout  = 8'b00000000; // 2694 :   0 - 0x0
      12'hA87: dout  = 8'b00000000; // 2695 :   0 - 0x0
      12'hA88: dout  = 8'b00000000; // 2696 :   0 - 0x0 -- Background 0x51
      12'hA89: dout  = 8'b00000000; // 2697 :   0 - 0x0
      12'hA8A: dout  = 8'b00000000; // 2698 :   0 - 0x0
      12'hA8B: dout  = 8'b00000000; // 2699 :   0 - 0x0
      12'hA8C: dout  = 8'b00000000; // 2700 :   0 - 0x0
      12'hA8D: dout  = 8'b00000000; // 2701 :   0 - 0x0
      12'hA8E: dout  = 8'b00000000; // 2702 :   0 - 0x0
      12'hA8F: dout  = 8'b00000000; // 2703 :   0 - 0x0
      12'hA90: dout  = 8'b00000000; // 2704 :   0 - 0x0 -- Background 0x52
      12'hA91: dout  = 8'b00000000; // 2705 :   0 - 0x0
      12'hA92: dout  = 8'b00000000; // 2706 :   0 - 0x0
      12'hA93: dout  = 8'b00000000; // 2707 :   0 - 0x0
      12'hA94: dout  = 8'b00000000; // 2708 :   0 - 0x0
      12'hA95: dout  = 8'b00000000; // 2709 :   0 - 0x0
      12'hA96: dout  = 8'b00000000; // 2710 :   0 - 0x0
      12'hA97: dout  = 8'b00000000; // 2711 :   0 - 0x0
      12'hA98: dout  = 8'b00000000; // 2712 :   0 - 0x0 -- Background 0x53
      12'hA99: dout  = 8'b00000000; // 2713 :   0 - 0x0
      12'hA9A: dout  = 8'b00000000; // 2714 :   0 - 0x0
      12'hA9B: dout  = 8'b00000000; // 2715 :   0 - 0x0
      12'hA9C: dout  = 8'b00000000; // 2716 :   0 - 0x0
      12'hA9D: dout  = 8'b00000000; // 2717 :   0 - 0x0
      12'hA9E: dout  = 8'b00000000; // 2718 :   0 - 0x0
      12'hA9F: dout  = 8'b00000000; // 2719 :   0 - 0x0
      12'hAA0: dout  = 8'b00000000; // 2720 :   0 - 0x0 -- Background 0x54
      12'hAA1: dout  = 8'b00000000; // 2721 :   0 - 0x0
      12'hAA2: dout  = 8'b00000000; // 2722 :   0 - 0x0
      12'hAA3: dout  = 8'b00000000; // 2723 :   0 - 0x0
      12'hAA4: dout  = 8'b00000000; // 2724 :   0 - 0x0
      12'hAA5: dout  = 8'b00000000; // 2725 :   0 - 0x0
      12'hAA6: dout  = 8'b00000000; // 2726 :   0 - 0x0
      12'hAA7: dout  = 8'b00000000; // 2727 :   0 - 0x0
      12'hAA8: dout  = 8'b00000000; // 2728 :   0 - 0x0 -- Background 0x55
      12'hAA9: dout  = 8'b00000000; // 2729 :   0 - 0x0
      12'hAAA: dout  = 8'b00000000; // 2730 :   0 - 0x0
      12'hAAB: dout  = 8'b00000000; // 2731 :   0 - 0x0
      12'hAAC: dout  = 8'b00000000; // 2732 :   0 - 0x0
      12'hAAD: dout  = 8'b00000000; // 2733 :   0 - 0x0
      12'hAAE: dout  = 8'b00000000; // 2734 :   0 - 0x0
      12'hAAF: dout  = 8'b00000000; // 2735 :   0 - 0x0
      12'hAB0: dout  = 8'b00000000; // 2736 :   0 - 0x0 -- Background 0x56
      12'hAB1: dout  = 8'b00000000; // 2737 :   0 - 0x0
      12'hAB2: dout  = 8'b00000000; // 2738 :   0 - 0x0
      12'hAB3: dout  = 8'b00000000; // 2739 :   0 - 0x0
      12'hAB4: dout  = 8'b00000000; // 2740 :   0 - 0x0
      12'hAB5: dout  = 8'b00000000; // 2741 :   0 - 0x0
      12'hAB6: dout  = 8'b00000000; // 2742 :   0 - 0x0
      12'hAB7: dout  = 8'b00000000; // 2743 :   0 - 0x0
      12'hAB8: dout  = 8'b00000000; // 2744 :   0 - 0x0 -- Background 0x57
      12'hAB9: dout  = 8'b00000000; // 2745 :   0 - 0x0
      12'hABA: dout  = 8'b00000000; // 2746 :   0 - 0x0
      12'hABB: dout  = 8'b00000000; // 2747 :   0 - 0x0
      12'hABC: dout  = 8'b00000000; // 2748 :   0 - 0x0
      12'hABD: dout  = 8'b00000000; // 2749 :   0 - 0x0
      12'hABE: dout  = 8'b00000000; // 2750 :   0 - 0x0
      12'hABF: dout  = 8'b00000000; // 2751 :   0 - 0x0
      12'hAC0: dout  = 8'b00000000; // 2752 :   0 - 0x0 -- Background 0x58
      12'hAC1: dout  = 8'b00000000; // 2753 :   0 - 0x0
      12'hAC2: dout  = 8'b00000000; // 2754 :   0 - 0x0
      12'hAC3: dout  = 8'b00000000; // 2755 :   0 - 0x0
      12'hAC4: dout  = 8'b00000000; // 2756 :   0 - 0x0
      12'hAC5: dout  = 8'b00000000; // 2757 :   0 - 0x0
      12'hAC6: dout  = 8'b00000000; // 2758 :   0 - 0x0
      12'hAC7: dout  = 8'b00000000; // 2759 :   0 - 0x0
      12'hAC8: dout  = 8'b00000000; // 2760 :   0 - 0x0 -- Background 0x59
      12'hAC9: dout  = 8'b00000000; // 2761 :   0 - 0x0
      12'hACA: dout  = 8'b00000000; // 2762 :   0 - 0x0
      12'hACB: dout  = 8'b00000000; // 2763 :   0 - 0x0
      12'hACC: dout  = 8'b00000000; // 2764 :   0 - 0x0
      12'hACD: dout  = 8'b00000000; // 2765 :   0 - 0x0
      12'hACE: dout  = 8'b00000000; // 2766 :   0 - 0x0
      12'hACF: dout  = 8'b00000000; // 2767 :   0 - 0x0
      12'hAD0: dout  = 8'b00000000; // 2768 :   0 - 0x0 -- Background 0x5a
      12'hAD1: dout  = 8'b00000000; // 2769 :   0 - 0x0
      12'hAD2: dout  = 8'b00000000; // 2770 :   0 - 0x0
      12'hAD3: dout  = 8'b00000000; // 2771 :   0 - 0x0
      12'hAD4: dout  = 8'b00000000; // 2772 :   0 - 0x0
      12'hAD5: dout  = 8'b00000000; // 2773 :   0 - 0x0
      12'hAD6: dout  = 8'b00000000; // 2774 :   0 - 0x0
      12'hAD7: dout  = 8'b00000000; // 2775 :   0 - 0x0
      12'hAD8: dout  = 8'b00000000; // 2776 :   0 - 0x0 -- Background 0x5b
      12'hAD9: dout  = 8'b00000000; // 2777 :   0 - 0x0
      12'hADA: dout  = 8'b00000000; // 2778 :   0 - 0x0
      12'hADB: dout  = 8'b00000000; // 2779 :   0 - 0x0
      12'hADC: dout  = 8'b00000000; // 2780 :   0 - 0x0
      12'hADD: dout  = 8'b00000000; // 2781 :   0 - 0x0
      12'hADE: dout  = 8'b00000000; // 2782 :   0 - 0x0
      12'hADF: dout  = 8'b00000000; // 2783 :   0 - 0x0
      12'hAE0: dout  = 8'b00000000; // 2784 :   0 - 0x0 -- Background 0x5c
      12'hAE1: dout  = 8'b00000000; // 2785 :   0 - 0x0
      12'hAE2: dout  = 8'b00000000; // 2786 :   0 - 0x0
      12'hAE3: dout  = 8'b00000000; // 2787 :   0 - 0x0
      12'hAE4: dout  = 8'b00000000; // 2788 :   0 - 0x0
      12'hAE5: dout  = 8'b00000000; // 2789 :   0 - 0x0
      12'hAE6: dout  = 8'b00000000; // 2790 :   0 - 0x0
      12'hAE7: dout  = 8'b00000000; // 2791 :   0 - 0x0
      12'hAE8: dout  = 8'b00000000; // 2792 :   0 - 0x0 -- Background 0x5d
      12'hAE9: dout  = 8'b00000000; // 2793 :   0 - 0x0
      12'hAEA: dout  = 8'b00000000; // 2794 :   0 - 0x0
      12'hAEB: dout  = 8'b00000000; // 2795 :   0 - 0x0
      12'hAEC: dout  = 8'b00000000; // 2796 :   0 - 0x0
      12'hAED: dout  = 8'b00000000; // 2797 :   0 - 0x0
      12'hAEE: dout  = 8'b00000000; // 2798 :   0 - 0x0
      12'hAEF: dout  = 8'b00000000; // 2799 :   0 - 0x0
      12'hAF0: dout  = 8'b00000000; // 2800 :   0 - 0x0 -- Background 0x5e
      12'hAF1: dout  = 8'b00000000; // 2801 :   0 - 0x0
      12'hAF2: dout  = 8'b00010000; // 2802 :  16 - 0x10
      12'hAF3: dout  = 8'b00010000; // 2803 :  16 - 0x10
      12'hAF4: dout  = 8'b00010000; // 2804 :  16 - 0x10
      12'hAF5: dout  = 8'b00010000; // 2805 :  16 - 0x10
      12'hAF6: dout  = 8'b00000000; // 2806 :   0 - 0x0
      12'hAF7: dout  = 8'b00000000; // 2807 :   0 - 0x0
      12'hAF8: dout  = 8'b00000000; // 2808 :   0 - 0x0 -- Background 0x5f
      12'hAF9: dout  = 8'b00000000; // 2809 :   0 - 0x0
      12'hAFA: dout  = 8'b00000000; // 2810 :   0 - 0x0
      12'hAFB: dout  = 8'b00000000; // 2811 :   0 - 0x0
      12'hAFC: dout  = 8'b00000000; // 2812 :   0 - 0x0
      12'hAFD: dout  = 8'b00000000; // 2813 :   0 - 0x0
      12'hAFE: dout  = 8'b00000000; // 2814 :   0 - 0x0
      12'hAFF: dout  = 8'b00000000; // 2815 :   0 - 0x0
      12'hB00: dout  = 8'b00000000; // 2816 :   0 - 0x0 -- Background 0x60
      12'hB01: dout  = 8'b00000000; // 2817 :   0 - 0x0
      12'hB02: dout  = 8'b00000000; // 2818 :   0 - 0x0
      12'hB03: dout  = 8'b00000000; // 2819 :   0 - 0x0
      12'hB04: dout  = 8'b00000000; // 2820 :   0 - 0x0
      12'hB05: dout  = 8'b00000000; // 2821 :   0 - 0x0
      12'hB06: dout  = 8'b00000000; // 2822 :   0 - 0x0
      12'hB07: dout  = 8'b00000000; // 2823 :   0 - 0x0
      12'hB08: dout  = 8'b00000000; // 2824 :   0 - 0x0 -- Background 0x61
      12'hB09: dout  = 8'b00000000; // 2825 :   0 - 0x0
      12'hB0A: dout  = 8'b00000000; // 2826 :   0 - 0x0
      12'hB0B: dout  = 8'b00000000; // 2827 :   0 - 0x0
      12'hB0C: dout  = 8'b00000000; // 2828 :   0 - 0x0
      12'hB0D: dout  = 8'b00000000; // 2829 :   0 - 0x0
      12'hB0E: dout  = 8'b00000000; // 2830 :   0 - 0x0
      12'hB0F: dout  = 8'b00000000; // 2831 :   0 - 0x0
      12'hB10: dout  = 8'b00000000; // 2832 :   0 - 0x0 -- Background 0x62
      12'hB11: dout  = 8'b00000000; // 2833 :   0 - 0x0
      12'hB12: dout  = 8'b00000000; // 2834 :   0 - 0x0
      12'hB13: dout  = 8'b00000000; // 2835 :   0 - 0x0
      12'hB14: dout  = 8'b00000000; // 2836 :   0 - 0x0
      12'hB15: dout  = 8'b00000000; // 2837 :   0 - 0x0
      12'hB16: dout  = 8'b00000000; // 2838 :   0 - 0x0
      12'hB17: dout  = 8'b00000000; // 2839 :   0 - 0x0
      12'hB18: dout  = 8'b00000000; // 2840 :   0 - 0x0 -- Background 0x63
      12'hB19: dout  = 8'b00000000; // 2841 :   0 - 0x0
      12'hB1A: dout  = 8'b00000000; // 2842 :   0 - 0x0
      12'hB1B: dout  = 8'b00000000; // 2843 :   0 - 0x0
      12'hB1C: dout  = 8'b00000000; // 2844 :   0 - 0x0
      12'hB1D: dout  = 8'b00000000; // 2845 :   0 - 0x0
      12'hB1E: dout  = 8'b00000000; // 2846 :   0 - 0x0
      12'hB1F: dout  = 8'b00000000; // 2847 :   0 - 0x0
      12'hB20: dout  = 8'b00000000; // 2848 :   0 - 0x0 -- Background 0x64
      12'hB21: dout  = 8'b00000000; // 2849 :   0 - 0x0
      12'hB22: dout  = 8'b00000000; // 2850 :   0 - 0x0
      12'hB23: dout  = 8'b00000000; // 2851 :   0 - 0x0
      12'hB24: dout  = 8'b00000000; // 2852 :   0 - 0x0
      12'hB25: dout  = 8'b00000000; // 2853 :   0 - 0x0
      12'hB26: dout  = 8'b00000000; // 2854 :   0 - 0x0
      12'hB27: dout  = 8'b00000000; // 2855 :   0 - 0x0
      12'hB28: dout  = 8'b00000000; // 2856 :   0 - 0x0 -- Background 0x65
      12'hB29: dout  = 8'b00000000; // 2857 :   0 - 0x0
      12'hB2A: dout  = 8'b00000000; // 2858 :   0 - 0x0
      12'hB2B: dout  = 8'b00000000; // 2859 :   0 - 0x0
      12'hB2C: dout  = 8'b00000000; // 2860 :   0 - 0x0
      12'hB2D: dout  = 8'b00000000; // 2861 :   0 - 0x0
      12'hB2E: dout  = 8'b00000000; // 2862 :   0 - 0x0
      12'hB2F: dout  = 8'b00000000; // 2863 :   0 - 0x0
      12'hB30: dout  = 8'b00000000; // 2864 :   0 - 0x0 -- Background 0x66
      12'hB31: dout  = 8'b00000000; // 2865 :   0 - 0x0
      12'hB32: dout  = 8'b00000000; // 2866 :   0 - 0x0
      12'hB33: dout  = 8'b00000000; // 2867 :   0 - 0x0
      12'hB34: dout  = 8'b00000000; // 2868 :   0 - 0x0
      12'hB35: dout  = 8'b00000000; // 2869 :   0 - 0x0
      12'hB36: dout  = 8'b00000000; // 2870 :   0 - 0x0
      12'hB37: dout  = 8'b00000000; // 2871 :   0 - 0x0
      12'hB38: dout  = 8'b00000000; // 2872 :   0 - 0x0 -- Background 0x67
      12'hB39: dout  = 8'b00000000; // 2873 :   0 - 0x0
      12'hB3A: dout  = 8'b00000000; // 2874 :   0 - 0x0
      12'hB3B: dout  = 8'b00000000; // 2875 :   0 - 0x0
      12'hB3C: dout  = 8'b00000000; // 2876 :   0 - 0x0
      12'hB3D: dout  = 8'b00000000; // 2877 :   0 - 0x0
      12'hB3E: dout  = 8'b00000000; // 2878 :   0 - 0x0
      12'hB3F: dout  = 8'b00000000; // 2879 :   0 - 0x0
      12'hB40: dout  = 8'b00000000; // 2880 :   0 - 0x0 -- Background 0x68
      12'hB41: dout  = 8'b00000000; // 2881 :   0 - 0x0
      12'hB42: dout  = 8'b00000000; // 2882 :   0 - 0x0
      12'hB43: dout  = 8'b00000001; // 2883 :   1 - 0x1
      12'hB44: dout  = 8'b00000001; // 2884 :   1 - 0x1
      12'hB45: dout  = 8'b00001011; // 2885 :  11 - 0xb
      12'hB46: dout  = 8'b00011100; // 2886 :  28 - 0x1c
      12'hB47: dout  = 8'b00111111; // 2887 :  63 - 0x3f
      12'hB48: dout  = 8'b00000000; // 2888 :   0 - 0x0 -- Background 0x69
      12'hB49: dout  = 8'b00000000; // 2889 :   0 - 0x0
      12'hB4A: dout  = 8'b00110000; // 2890 :  48 - 0x30
      12'hB4B: dout  = 8'b01111000; // 2891 : 120 - 0x78
      12'hB4C: dout  = 8'b10000000; // 2892 : 128 - 0x80
      12'hB4D: dout  = 8'b11110000; // 2893 : 240 - 0xf0
      12'hB4E: dout  = 8'b11111000; // 2894 : 248 - 0xf8
      12'hB4F: dout  = 8'b11111100; // 2895 : 252 - 0xfc
      12'hB50: dout  = 8'b00111111; // 2896 :  63 - 0x3f -- Background 0x6a
      12'hB51: dout  = 8'b00111111; // 2897 :  63 - 0x3f
      12'hB52: dout  = 8'b00111111; // 2898 :  63 - 0x3f
      12'hB53: dout  = 8'b00011111; // 2899 :  31 - 0x1f
      12'hB54: dout  = 8'b00011111; // 2900 :  31 - 0x1f
      12'hB55: dout  = 8'b00000111; // 2901 :   7 - 0x7
      12'hB56: dout  = 8'b00000000; // 2902 :   0 - 0x0
      12'hB57: dout  = 8'b00000000; // 2903 :   0 - 0x0
      12'hB58: dout  = 8'b11111100; // 2904 : 252 - 0xfc -- Background 0x6b
      12'hB59: dout  = 8'b11101100; // 2905 : 236 - 0xec
      12'hB5A: dout  = 8'b11101100; // 2906 : 236 - 0xec
      12'hB5B: dout  = 8'b11011000; // 2907 : 216 - 0xd8
      12'hB5C: dout  = 8'b11111000; // 2908 : 248 - 0xf8
      12'hB5D: dout  = 8'b11100000; // 2909 : 224 - 0xe0
      12'hB5E: dout  = 8'b00000000; // 2910 :   0 - 0x0
      12'hB5F: dout  = 8'b00000000; // 2911 :   0 - 0x0
      12'hB60: dout  = 8'b00000000; // 2912 :   0 - 0x0 -- Background 0x6c
      12'hB61: dout  = 8'b00000000; // 2913 :   0 - 0x0
      12'hB62: dout  = 8'b00000001; // 2914 :   1 - 0x1
      12'hB63: dout  = 8'b00011101; // 2915 :  29 - 0x1d
      12'hB64: dout  = 8'b00111110; // 2916 :  62 - 0x3e
      12'hB65: dout  = 8'b00111111; // 2917 :  63 - 0x3f
      12'hB66: dout  = 8'b00111111; // 2918 :  63 - 0x3f
      12'hB67: dout  = 8'b00111111; // 2919 :  63 - 0x3f
      12'hB68: dout  = 8'b00000000; // 2920 :   0 - 0x0 -- Background 0x6d
      12'hB69: dout  = 8'b10000000; // 2921 : 128 - 0x80
      12'hB6A: dout  = 8'b00000000; // 2922 :   0 - 0x0
      12'hB6B: dout  = 8'b01110000; // 2923 : 112 - 0x70
      12'hB6C: dout  = 8'b11111000; // 2924 : 248 - 0xf8
      12'hB6D: dout  = 8'b11111100; // 2925 : 252 - 0xfc
      12'hB6E: dout  = 8'b11111100; // 2926 : 252 - 0xfc
      12'hB6F: dout  = 8'b11111100; // 2927 : 252 - 0xfc
      12'hB70: dout  = 8'b00111111; // 2928 :  63 - 0x3f -- Background 0x6e
      12'hB71: dout  = 8'b00111111; // 2929 :  63 - 0x3f
      12'hB72: dout  = 8'b00011111; // 2930 :  31 - 0x1f
      12'hB73: dout  = 8'b00011111; // 2931 :  31 - 0x1f
      12'hB74: dout  = 8'b00001111; // 2932 :  15 - 0xf
      12'hB75: dout  = 8'b00000110; // 2933 :   6 - 0x6
      12'hB76: dout  = 8'b00000000; // 2934 :   0 - 0x0
      12'hB77: dout  = 8'b00000000; // 2935 :   0 - 0x0
      12'hB78: dout  = 8'b11101100; // 2936 : 236 - 0xec -- Background 0x6f
      12'hB79: dout  = 8'b11101100; // 2937 : 236 - 0xec
      12'hB7A: dout  = 8'b11011000; // 2938 : 216 - 0xd8
      12'hB7B: dout  = 8'b11111000; // 2939 : 248 - 0xf8
      12'hB7C: dout  = 8'b11110000; // 2940 : 240 - 0xf0
      12'hB7D: dout  = 8'b11100000; // 2941 : 224 - 0xe0
      12'hB7E: dout  = 8'b00000000; // 2942 :   0 - 0x0
      12'hB7F: dout  = 8'b00000000; // 2943 :   0 - 0x0
      12'hB80: dout  = 8'b00000000; // 2944 :   0 - 0x0 -- Background 0x70
      12'hB81: dout  = 8'b00000000; // 2945 :   0 - 0x0
      12'hB82: dout  = 8'b00000000; // 2946 :   0 - 0x0
      12'hB83: dout  = 8'b00000000; // 2947 :   0 - 0x0
      12'hB84: dout  = 8'b00000000; // 2948 :   0 - 0x0
      12'hB85: dout  = 8'b00000000; // 2949 :   0 - 0x0
      12'hB86: dout  = 8'b00000000; // 2950 :   0 - 0x0
      12'hB87: dout  = 8'b00000000; // 2951 :   0 - 0x0
      12'hB88: dout  = 8'b00000000; // 2952 :   0 - 0x0 -- Background 0x71
      12'hB89: dout  = 8'b00000000; // 2953 :   0 - 0x0
      12'hB8A: dout  = 8'b00000000; // 2954 :   0 - 0x0
      12'hB8B: dout  = 8'b00000000; // 2955 :   0 - 0x0
      12'hB8C: dout  = 8'b00000000; // 2956 :   0 - 0x0
      12'hB8D: dout  = 8'b00000000; // 2957 :   0 - 0x0
      12'hB8E: dout  = 8'b00000000; // 2958 :   0 - 0x0
      12'hB8F: dout  = 8'b00000000; // 2959 :   0 - 0x0
      12'hB90: dout  = 8'b00000000; // 2960 :   0 - 0x0 -- Background 0x72
      12'hB91: dout  = 8'b00000000; // 2961 :   0 - 0x0
      12'hB92: dout  = 8'b00000000; // 2962 :   0 - 0x0
      12'hB93: dout  = 8'b00000000; // 2963 :   0 - 0x0
      12'hB94: dout  = 8'b00000000; // 2964 :   0 - 0x0
      12'hB95: dout  = 8'b00000000; // 2965 :   0 - 0x0
      12'hB96: dout  = 8'b00000000; // 2966 :   0 - 0x0
      12'hB97: dout  = 8'b00000000; // 2967 :   0 - 0x0
      12'hB98: dout  = 8'b00000000; // 2968 :   0 - 0x0 -- Background 0x73
      12'hB99: dout  = 8'b00000000; // 2969 :   0 - 0x0
      12'hB9A: dout  = 8'b00000000; // 2970 :   0 - 0x0
      12'hB9B: dout  = 8'b00000000; // 2971 :   0 - 0x0
      12'hB9C: dout  = 8'b00000000; // 2972 :   0 - 0x0
      12'hB9D: dout  = 8'b00000000; // 2973 :   0 - 0x0
      12'hB9E: dout  = 8'b00000000; // 2974 :   0 - 0x0
      12'hB9F: dout  = 8'b00000000; // 2975 :   0 - 0x0
      12'hBA0: dout  = 8'b00000000; // 2976 :   0 - 0x0 -- Background 0x74
      12'hBA1: dout  = 8'b00000000; // 2977 :   0 - 0x0
      12'hBA2: dout  = 8'b00000000; // 2978 :   0 - 0x0
      12'hBA3: dout  = 8'b00000000; // 2979 :   0 - 0x0
      12'hBA4: dout  = 8'b00010001; // 2980 :  17 - 0x11
      12'hBA5: dout  = 8'b00010011; // 2981 :  19 - 0x13
      12'hBA6: dout  = 8'b00011111; // 2982 :  31 - 0x1f
      12'hBA7: dout  = 8'b00011111; // 2983 :  31 - 0x1f
      12'hBA8: dout  = 8'b00000000; // 2984 :   0 - 0x0 -- Background 0x75
      12'hBA9: dout  = 8'b00000000; // 2985 :   0 - 0x0
      12'hBAA: dout  = 8'b00000000; // 2986 :   0 - 0x0
      12'hBAB: dout  = 8'b10000000; // 2987 : 128 - 0x80
      12'hBAC: dout  = 8'b11000100; // 2988 : 196 - 0xc4
      12'hBAD: dout  = 8'b11100100; // 2989 : 228 - 0xe4
      12'hBAE: dout  = 8'b11111100; // 2990 : 252 - 0xfc
      12'hBAF: dout  = 8'b11111100; // 2991 : 252 - 0xfc
      12'hBB0: dout  = 8'b00011111; // 2992 :  31 - 0x1f -- Background 0x76
      12'hBB1: dout  = 8'b00001110; // 2993 :  14 - 0xe
      12'hBB2: dout  = 8'b00000110; // 2994 :   6 - 0x6
      12'hBB3: dout  = 8'b00000010; // 2995 :   2 - 0x2
      12'hBB4: dout  = 8'b00000000; // 2996 :   0 - 0x0
      12'hBB5: dout  = 8'b00000000; // 2997 :   0 - 0x0
      12'hBB6: dout  = 8'b00000000; // 2998 :   0 - 0x0
      12'hBB7: dout  = 8'b00000000; // 2999 :   0 - 0x0
      12'hBB8: dout  = 8'b11111100; // 3000 : 252 - 0xfc -- Background 0x77
      12'hBB9: dout  = 8'b10111000; // 3001 : 184 - 0xb8
      12'hBBA: dout  = 8'b10110000; // 3002 : 176 - 0xb0
      12'hBBB: dout  = 8'b10100000; // 3003 : 160 - 0xa0
      12'hBBC: dout  = 8'b10000000; // 3004 : 128 - 0x80
      12'hBBD: dout  = 8'b00000000; // 3005 :   0 - 0x0
      12'hBBE: dout  = 8'b00000000; // 3006 :   0 - 0x0
      12'hBBF: dout  = 8'b00000000; // 3007 :   0 - 0x0
      12'hBC0: dout  = 8'b00000000; // 3008 :   0 - 0x0 -- Background 0x78
      12'hBC1: dout  = 8'b00000000; // 3009 :   0 - 0x0
      12'hBC2: dout  = 8'b00000000; // 3010 :   0 - 0x0
      12'hBC3: dout  = 8'b00000001; // 3011 :   1 - 0x1
      12'hBC4: dout  = 8'b00000011; // 3012 :   3 - 0x3
      12'hBC5: dout  = 8'b00000110; // 3013 :   6 - 0x6
      12'hBC6: dout  = 8'b00000110; // 3014 :   6 - 0x6
      12'hBC7: dout  = 8'b00001111; // 3015 :  15 - 0xf
      12'hBC8: dout  = 8'b00000000; // 3016 :   0 - 0x0 -- Background 0x79
      12'hBC9: dout  = 8'b00011000; // 3017 :  24 - 0x18
      12'hBCA: dout  = 8'b11110100; // 3018 : 244 - 0xf4
      12'hBCB: dout  = 8'b11111000; // 3019 : 248 - 0xf8
      12'hBCC: dout  = 8'b00111000; // 3020 :  56 - 0x38
      12'hBCD: dout  = 8'b01111100; // 3021 : 124 - 0x7c
      12'hBCE: dout  = 8'b11111100; // 3022 : 252 - 0xfc
      12'hBCF: dout  = 8'b11111100; // 3023 : 252 - 0xfc
      12'hBD0: dout  = 8'b00001111; // 3024 :  15 - 0xf -- Background 0x7a
      12'hBD1: dout  = 8'b00011111; // 3025 :  31 - 0x1f
      12'hBD2: dout  = 8'b00110000; // 3026 :  48 - 0x30
      12'hBD3: dout  = 8'b00111000; // 3027 :  56 - 0x38
      12'hBD4: dout  = 8'b00011101; // 3028 :  29 - 0x1d
      12'hBD5: dout  = 8'b00000011; // 3029 :   3 - 0x3
      12'hBD6: dout  = 8'b00000011; // 3030 :   3 - 0x3
      12'hBD7: dout  = 8'b00000000; // 3031 :   0 - 0x0
      12'hBD8: dout  = 8'b11111100; // 3032 : 252 - 0xfc -- Background 0x7b
      12'hBD9: dout  = 8'b11111100; // 3033 : 252 - 0xfc
      12'hBDA: dout  = 8'b01111100; // 3034 : 124 - 0x7c
      12'hBDB: dout  = 8'b10001110; // 3035 : 142 - 0x8e
      12'hBDC: dout  = 8'b10000110; // 3036 : 134 - 0x86
      12'hBDD: dout  = 8'b10011100; // 3037 : 156 - 0x9c
      12'hBDE: dout  = 8'b01111000; // 3038 : 120 - 0x78
      12'hBDF: dout  = 8'b00000000; // 3039 :   0 - 0x0
      12'hBE0: dout  = 8'b00000000; // 3040 :   0 - 0x0 -- Background 0x7c
      12'hBE1: dout  = 8'b00000001; // 3041 :   1 - 0x1
      12'hBE2: dout  = 8'b00000110; // 3042 :   6 - 0x6
      12'hBE3: dout  = 8'b00000111; // 3043 :   7 - 0x7
      12'hBE4: dout  = 8'b00000111; // 3044 :   7 - 0x7
      12'hBE5: dout  = 8'b00000111; // 3045 :   7 - 0x7
      12'hBE6: dout  = 8'b00000001; // 3046 :   1 - 0x1
      12'hBE7: dout  = 8'b00000011; // 3047 :   3 - 0x3
      12'hBE8: dout  = 8'b00000000; // 3048 :   0 - 0x0 -- Background 0x7d
      12'hBE9: dout  = 8'b11000000; // 3049 : 192 - 0xc0
      12'hBEA: dout  = 8'b00110000; // 3050 :  48 - 0x30
      12'hBEB: dout  = 8'b11110000; // 3051 : 240 - 0xf0
      12'hBEC: dout  = 8'b11110000; // 3052 : 240 - 0xf0
      12'hBED: dout  = 8'b11110000; // 3053 : 240 - 0xf0
      12'hBEE: dout  = 8'b01000000; // 3054 :  64 - 0x40
      12'hBEF: dout  = 8'b01000000; // 3055 :  64 - 0x40
      12'hBF0: dout  = 8'b00000001; // 3056 :   1 - 0x1 -- Background 0x7e
      12'hBF1: dout  = 8'b00000000; // 3057 :   0 - 0x0
      12'hBF2: dout  = 8'b00000001; // 3058 :   1 - 0x1
      12'hBF3: dout  = 8'b00000011; // 3059 :   3 - 0x3
      12'hBF4: dout  = 8'b00000001; // 3060 :   1 - 0x1
      12'hBF5: dout  = 8'b00000000; // 3061 :   0 - 0x0
      12'hBF6: dout  = 8'b00000000; // 3062 :   0 - 0x0
      12'hBF7: dout  = 8'b00000000; // 3063 :   0 - 0x0
      12'hBF8: dout  = 8'b01000000; // 3064 :  64 - 0x40 -- Background 0x7f
      12'hBF9: dout  = 8'b01000000; // 3065 :  64 - 0x40
      12'hBFA: dout  = 8'b01000000; // 3066 :  64 - 0x40
      12'hBFB: dout  = 8'b01000000; // 3067 :  64 - 0x40
      12'hBFC: dout  = 8'b01000000; // 3068 :  64 - 0x40
      12'hBFD: dout  = 8'b10000000; // 3069 : 128 - 0x80
      12'hBFE: dout  = 8'b00000000; // 3070 :   0 - 0x0
      12'hBFF: dout  = 8'b00000000; // 3071 :   0 - 0x0
      12'hC00: dout  = 8'b00000000; // 3072 :   0 - 0x0 -- Background 0x80
      12'hC01: dout  = 8'b00000000; // 3073 :   0 - 0x0
      12'hC02: dout  = 8'b00000000; // 3074 :   0 - 0x0
      12'hC03: dout  = 8'b00000000; // 3075 :   0 - 0x0
      12'hC04: dout  = 8'b00000000; // 3076 :   0 - 0x0
      12'hC05: dout  = 8'b00011111; // 3077 :  31 - 0x1f
      12'hC06: dout  = 8'b00010000; // 3078 :  16 - 0x10
      12'hC07: dout  = 8'b00010111; // 3079 :  23 - 0x17
      12'hC08: dout  = 8'b00000000; // 3080 :   0 - 0x0 -- Background 0x81
      12'hC09: dout  = 8'b00000000; // 3081 :   0 - 0x0
      12'hC0A: dout  = 8'b00000000; // 3082 :   0 - 0x0
      12'hC0B: dout  = 8'b00000000; // 3083 :   0 - 0x0
      12'hC0C: dout  = 8'b00000000; // 3084 :   0 - 0x0
      12'hC0D: dout  = 8'b11111111; // 3085 : 255 - 0xff
      12'hC0E: dout  = 8'b00000000; // 3086 :   0 - 0x0
      12'hC0F: dout  = 8'b11111111; // 3087 : 255 - 0xff
      12'hC10: dout  = 8'b00000000; // 3088 :   0 - 0x0 -- Background 0x82
      12'hC11: dout  = 8'b00000000; // 3089 :   0 - 0x0
      12'hC12: dout  = 8'b00000000; // 3090 :   0 - 0x0
      12'hC13: dout  = 8'b00000000; // 3091 :   0 - 0x0
      12'hC14: dout  = 8'b00000000; // 3092 :   0 - 0x0
      12'hC15: dout  = 8'b10000000; // 3093 : 128 - 0x80
      12'hC16: dout  = 8'b00000000; // 3094 :   0 - 0x0
      12'hC17: dout  = 8'b11000000; // 3095 : 192 - 0xc0
      12'hC18: dout  = 8'b00000000; // 3096 :   0 - 0x0 -- Background 0x83
      12'hC19: dout  = 8'b00000000; // 3097 :   0 - 0x0
      12'hC1A: dout  = 8'b00000000; // 3098 :   0 - 0x0
      12'hC1B: dout  = 8'b00000000; // 3099 :   0 - 0x0
      12'hC1C: dout  = 8'b00000000; // 3100 :   0 - 0x0
      12'hC1D: dout  = 8'b00001000; // 3101 :   8 - 0x8
      12'hC1E: dout  = 8'b00001000; // 3102 :   8 - 0x8
      12'hC1F: dout  = 8'b00010110; // 3103 :  22 - 0x16
      12'hC20: dout  = 8'b00000000; // 3104 :   0 - 0x0 -- Background 0x84
      12'hC21: dout  = 8'b00000000; // 3105 :   0 - 0x0
      12'hC22: dout  = 8'b00000000; // 3106 :   0 - 0x0
      12'hC23: dout  = 8'b00000000; // 3107 :   0 - 0x0
      12'hC24: dout  = 8'b00000000; // 3108 :   0 - 0x0
      12'hC25: dout  = 8'b00000000; // 3109 :   0 - 0x0
      12'hC26: dout  = 8'b01000000; // 3110 :  64 - 0x40
      12'hC27: dout  = 8'b11000000; // 3111 : 192 - 0xc0
      12'hC28: dout  = 8'b00000000; // 3112 :   0 - 0x0 -- Background 0x85
      12'hC29: dout  = 8'b00000000; // 3113 :   0 - 0x0
      12'hC2A: dout  = 8'b00000000; // 3114 :   0 - 0x0
      12'hC2B: dout  = 8'b00000000; // 3115 :   0 - 0x0
      12'hC2C: dout  = 8'b00000000; // 3116 :   0 - 0x0
      12'hC2D: dout  = 8'b00000001; // 3117 :   1 - 0x1
      12'hC2E: dout  = 8'b00000111; // 3118 :   7 - 0x7
      12'hC2F: dout  = 8'b00001100; // 3119 :  12 - 0xc
      12'hC30: dout  = 8'b00000000; // 3120 :   0 - 0x0 -- Background 0x86
      12'hC31: dout  = 8'b00000000; // 3121 :   0 - 0x0
      12'hC32: dout  = 8'b00000000; // 3122 :   0 - 0x0
      12'hC33: dout  = 8'b00000000; // 3123 :   0 - 0x0
      12'hC34: dout  = 8'b00000000; // 3124 :   0 - 0x0
      12'hC35: dout  = 8'b11000000; // 3125 : 192 - 0xc0
      12'hC36: dout  = 8'b00111111; // 3126 :  63 - 0x3f
      12'hC37: dout  = 8'b11111111; // 3127 : 255 - 0xff
      12'hC38: dout  = 8'b00000000; // 3128 :   0 - 0x0 -- Background 0x87
      12'hC39: dout  = 8'b00000000; // 3129 :   0 - 0x0
      12'hC3A: dout  = 8'b00000000; // 3130 :   0 - 0x0
      12'hC3B: dout  = 8'b00000000; // 3131 :   0 - 0x0
      12'hC3C: dout  = 8'b00000000; // 3132 :   0 - 0x0
      12'hC3D: dout  = 8'b00000000; // 3133 :   0 - 0x0
      12'hC3E: dout  = 8'b00000000; // 3134 :   0 - 0x0
      12'hC3F: dout  = 8'b11000000; // 3135 : 192 - 0xc0
      12'hC40: dout  = 8'b00000000; // 3136 :   0 - 0x0 -- Background 0x88
      12'hC41: dout  = 8'b00000000; // 3137 :   0 - 0x0
      12'hC42: dout  = 8'b00000000; // 3138 :   0 - 0x0
      12'hC43: dout  = 8'b00000000; // 3139 :   0 - 0x0
      12'hC44: dout  = 8'b00000000; // 3140 :   0 - 0x0
      12'hC45: dout  = 8'b00000000; // 3141 :   0 - 0x0
      12'hC46: dout  = 8'b00000000; // 3142 :   0 - 0x0
      12'hC47: dout  = 8'b00000000; // 3143 :   0 - 0x0
      12'hC48: dout  = 8'b00000000; // 3144 :   0 - 0x0 -- Background 0x89
      12'hC49: dout  = 8'b00000000; // 3145 :   0 - 0x0
      12'hC4A: dout  = 8'b00000000; // 3146 :   0 - 0x0
      12'hC4B: dout  = 8'b00000000; // 3147 :   0 - 0x0
      12'hC4C: dout  = 8'b00000000; // 3148 :   0 - 0x0
      12'hC4D: dout  = 8'b01000100; // 3149 :  68 - 0x44
      12'hC4E: dout  = 8'b01010110; // 3150 :  86 - 0x56
      12'hC4F: dout  = 8'b01011011; // 3151 :  91 - 0x5b
      12'hC50: dout  = 8'b00000000; // 3152 :   0 - 0x0 -- Background 0x8a
      12'hC51: dout  = 8'b00000000; // 3153 :   0 - 0x0
      12'hC52: dout  = 8'b00000000; // 3154 :   0 - 0x0
      12'hC53: dout  = 8'b00000000; // 3155 :   0 - 0x0
      12'hC54: dout  = 8'b00000000; // 3156 :   0 - 0x0
      12'hC55: dout  = 8'b00000000; // 3157 :   0 - 0x0
      12'hC56: dout  = 8'b00000000; // 3158 :   0 - 0x0
      12'hC57: dout  = 8'b00000000; // 3159 :   0 - 0x0
      12'hC58: dout  = 8'b00000000; // 3160 :   0 - 0x0 -- Background 0x8b
      12'hC59: dout  = 8'b00000000; // 3161 :   0 - 0x0
      12'hC5A: dout  = 8'b00000000; // 3162 :   0 - 0x0
      12'hC5B: dout  = 8'b00000000; // 3163 :   0 - 0x0
      12'hC5C: dout  = 8'b00000000; // 3164 :   0 - 0x0
      12'hC5D: dout  = 8'b00010000; // 3165 :  16 - 0x10
      12'hC5E: dout  = 8'b00110100; // 3166 :  52 - 0x34
      12'hC5F: dout  = 8'b01101101; // 3167 : 109 - 0x6d
      12'hC60: dout  = 8'b00000000; // 3168 :   0 - 0x0 -- Background 0x8c
      12'hC61: dout  = 8'b00000000; // 3169 :   0 - 0x0
      12'hC62: dout  = 8'b00000000; // 3170 :   0 - 0x0
      12'hC63: dout  = 8'b00000000; // 3171 :   0 - 0x0
      12'hC64: dout  = 8'b00000000; // 3172 :   0 - 0x0
      12'hC65: dout  = 8'b00000000; // 3173 :   0 - 0x0
      12'hC66: dout  = 8'b00000000; // 3174 :   0 - 0x0
      12'hC67: dout  = 8'b00000000; // 3175 :   0 - 0x0
      12'hC68: dout  = 8'b00000000; // 3176 :   0 - 0x0 -- Background 0x8d
      12'hC69: dout  = 8'b00000000; // 3177 :   0 - 0x0
      12'hC6A: dout  = 8'b00000000; // 3178 :   0 - 0x0
      12'hC6B: dout  = 8'b00000000; // 3179 :   0 - 0x0
      12'hC6C: dout  = 8'b01000000; // 3180 :  64 - 0x40
      12'hC6D: dout  = 8'b01001000; // 3181 :  72 - 0x48
      12'hC6E: dout  = 8'b10101000; // 3182 : 168 - 0xa8
      12'hC6F: dout  = 8'b10101100; // 3183 : 172 - 0xac
      12'hC70: dout  = 8'b00000000; // 3184 :   0 - 0x0 -- Background 0x8e
      12'hC71: dout  = 8'b00000000; // 3185 :   0 - 0x0
      12'hC72: dout  = 8'b00000000; // 3186 :   0 - 0x0
      12'hC73: dout  = 8'b00000000; // 3187 :   0 - 0x0
      12'hC74: dout  = 8'b00000010; // 3188 :   2 - 0x2
      12'hC75: dout  = 8'b00000010; // 3189 :   2 - 0x2
      12'hC76: dout  = 8'b00000010; // 3190 :   2 - 0x2
      12'hC77: dout  = 8'b00000010; // 3191 :   2 - 0x2
      12'hC78: dout  = 8'b00000000; // 3192 :   0 - 0x0 -- Background 0x8f
      12'hC79: dout  = 8'b00000000; // 3193 :   0 - 0x0
      12'hC7A: dout  = 8'b00000000; // 3194 :   0 - 0x0
      12'hC7B: dout  = 8'b00000011; // 3195 :   3 - 0x3
      12'hC7C: dout  = 8'b01000011; // 3196 :  67 - 0x43
      12'hC7D: dout  = 8'b01100010; // 3197 :  98 - 0x62
      12'hC7E: dout  = 8'b10110010; // 3198 : 178 - 0xb2
      12'hC7F: dout  = 8'b11011010; // 3199 : 218 - 0xda
      12'hC80: dout  = 8'b00000000; // 3200 :   0 - 0x0 -- Background 0x90
      12'hC81: dout  = 8'b00000000; // 3201 :   0 - 0x0
      12'hC82: dout  = 8'b00000000; // 3202 :   0 - 0x0
      12'hC83: dout  = 8'b11111100; // 3203 : 252 - 0xfc
      12'hC84: dout  = 8'b11111100; // 3204 : 252 - 0xfc
      12'hC85: dout  = 8'b00000000; // 3205 :   0 - 0x0
      12'hC86: dout  = 8'b11111111; // 3206 : 255 - 0xff
      12'hC87: dout  = 8'b11111111; // 3207 : 255 - 0xff
      12'hC88: dout  = 8'b00000000; // 3208 :   0 - 0x0 -- Background 0x91
      12'hC89: dout  = 8'b00000000; // 3209 :   0 - 0x0
      12'hC8A: dout  = 8'b00000000; // 3210 :   0 - 0x0
      12'hC8B: dout  = 8'b00000000; // 3211 :   0 - 0x0
      12'hC8C: dout  = 8'b00000000; // 3212 :   0 - 0x0
      12'hC8D: dout  = 8'b00000000; // 3213 :   0 - 0x0
      12'hC8E: dout  = 8'b00000000; // 3214 :   0 - 0x0
      12'hC8F: dout  = 8'b00000000; // 3215 :   0 - 0x0
      12'hC90: dout  = 8'b00010111; // 3216 :  23 - 0x17 -- Background 0x92
      12'hC91: dout  = 8'b00010111; // 3217 :  23 - 0x17
      12'hC92: dout  = 8'b00010111; // 3218 :  23 - 0x17
      12'hC93: dout  = 8'b00010111; // 3219 :  23 - 0x17
      12'hC94: dout  = 8'b00010111; // 3220 :  23 - 0x17
      12'hC95: dout  = 8'b00010111; // 3221 :  23 - 0x17
      12'hC96: dout  = 8'b00010111; // 3222 :  23 - 0x17
      12'hC97: dout  = 8'b00010111; // 3223 :  23 - 0x17
      12'hC98: dout  = 8'b11111111; // 3224 : 255 - 0xff -- Background 0x93
      12'hC99: dout  = 8'b11111111; // 3225 : 255 - 0xff
      12'hC9A: dout  = 8'b11111111; // 3226 : 255 - 0xff
      12'hC9B: dout  = 8'b11111111; // 3227 : 255 - 0xff
      12'hC9C: dout  = 8'b11111001; // 3228 : 249 - 0xf9
      12'hC9D: dout  = 8'b11111001; // 3229 : 249 - 0xf9
      12'hC9E: dout  = 8'b11111111; // 3230 : 255 - 0xff
      12'hC9F: dout  = 8'b11111111; // 3231 : 255 - 0xff
      12'hCA0: dout  = 8'b11110000; // 3232 : 240 - 0xf0 -- Background 0x94
      12'hCA1: dout  = 8'b11111000; // 3233 : 248 - 0xf8
      12'hCA2: dout  = 8'b11111000; // 3234 : 248 - 0xf8
      12'hCA3: dout  = 8'b11111100; // 3235 : 252 - 0xfc
      12'hCA4: dout  = 8'b11111100; // 3236 : 252 - 0xfc
      12'hCA5: dout  = 8'b11111100; // 3237 : 252 - 0xfc
      12'hCA6: dout  = 8'b01111100; // 3238 : 124 - 0x7c
      12'hCA7: dout  = 8'b01111100; // 3239 : 124 - 0x7c
      12'hCA8: dout  = 8'b00010111; // 3240 :  23 - 0x17 -- Background 0x95
      12'hCA9: dout  = 8'b00101111; // 3241 :  47 - 0x2f
      12'hCAA: dout  = 8'b00101111; // 3242 :  47 - 0x2f
      12'hCAB: dout  = 8'b01011111; // 3243 :  95 - 0x5f
      12'hCAC: dout  = 8'b01011111; // 3244 :  95 - 0x5f
      12'hCAD: dout  = 8'b10111111; // 3245 : 191 - 0xbf
      12'hCAE: dout  = 8'b10111111; // 3246 : 191 - 0xbf
      12'hCAF: dout  = 8'b01111111; // 3247 : 127 - 0x7f
      12'hCB0: dout  = 8'b01100000; // 3248 :  96 - 0x60 -- Background 0x96
      12'hCB1: dout  = 8'b01100000; // 3249 :  96 - 0x60
      12'hCB2: dout  = 8'b10110000; // 3250 : 176 - 0xb0
      12'hCB3: dout  = 8'b10110000; // 3251 : 176 - 0xb0
      12'hCB4: dout  = 8'b11011000; // 3252 : 216 - 0xd8
      12'hCB5: dout  = 8'b11011000; // 3253 : 216 - 0xd8
      12'hCB6: dout  = 8'b11101100; // 3254 : 236 - 0xec
      12'hCB7: dout  = 8'b11101100; // 3255 : 236 - 0xec
      12'hCB8: dout  = 8'b00110011; // 3256 :  51 - 0x33 -- Background 0x97
      12'hCB9: dout  = 8'b00101111; // 3257 :  47 - 0x2f
      12'hCBA: dout  = 8'b01101111; // 3258 : 111 - 0x6f
      12'hCBB: dout  = 8'b01011111; // 3259 :  95 - 0x5f
      12'hCBC: dout  = 8'b11011111; // 3260 : 223 - 0xdf
      12'hCBD: dout  = 8'b10111111; // 3261 : 191 - 0xbf
      12'hCBE: dout  = 8'b10111111; // 3262 : 191 - 0xbf
      12'hCBF: dout  = 8'b10111111; // 3263 : 191 - 0xbf
      12'hCC0: dout  = 8'b11111111; // 3264 : 255 - 0xff -- Background 0x98
      12'hCC1: dout  = 8'b11111111; // 3265 : 255 - 0xff
      12'hCC2: dout  = 8'b11111111; // 3266 : 255 - 0xff
      12'hCC3: dout  = 8'b11111110; // 3267 : 254 - 0xfe
      12'hCC4: dout  = 8'b11111001; // 3268 : 249 - 0xf9
      12'hCC5: dout  = 8'b11100111; // 3269 : 231 - 0xe7
      12'hCC6: dout  = 8'b11111100; // 3270 : 252 - 0xfc
      12'hCC7: dout  = 8'b11110011; // 3271 : 243 - 0xf3
      12'hCC8: dout  = 8'b11110000; // 3272 : 240 - 0xf0 -- Background 0x99
      12'hCC9: dout  = 8'b11111000; // 3273 : 248 - 0xf8
      12'hCCA: dout  = 8'b11111000; // 3274 : 248 - 0xf8
      12'hCCB: dout  = 8'b01110000; // 3275 : 112 - 0x70
      12'hCCC: dout  = 8'b11001100; // 3276 : 204 - 0xcc
      12'hCCD: dout  = 8'b00110000; // 3277 :  48 - 0x30
      12'hCCE: dout  = 8'b11000000; // 3278 : 192 - 0xc0
      12'hCCF: dout  = 8'b00000000; // 3279 :   0 - 0x0
      12'hCD0: dout  = 8'b00000000; // 3280 :   0 - 0x0 -- Background 0x9a
      12'hCD1: dout  = 8'b00000000; // 3281 :   0 - 0x0
      12'hCD2: dout  = 8'b00000000; // 3282 :   0 - 0x0
      12'hCD3: dout  = 8'b00000000; // 3283 :   0 - 0x0
      12'hCD4: dout  = 8'b00111111; // 3284 :  63 - 0x3f
      12'hCD5: dout  = 8'b00100000; // 3285 :  32 - 0x20
      12'hCD6: dout  = 8'b00101111; // 3286 :  47 - 0x2f
      12'hCD7: dout  = 8'b00101111; // 3287 :  47 - 0x2f
      12'hCD8: dout  = 8'b00000000; // 3288 :   0 - 0x0 -- Background 0x9b
      12'hCD9: dout  = 8'b00000000; // 3289 :   0 - 0x0
      12'hCDA: dout  = 8'b00000000; // 3290 :   0 - 0x0
      12'hCDB: dout  = 8'b00000000; // 3291 :   0 - 0x0
      12'hCDC: dout  = 8'b11100000; // 3292 : 224 - 0xe0
      12'hCDD: dout  = 8'b00000000; // 3293 :   0 - 0x0
      12'hCDE: dout  = 8'b11110000; // 3294 : 240 - 0xf0
      12'hCDF: dout  = 8'b11110000; // 3295 : 240 - 0xf0
      12'hCE0: dout  = 8'b01011101; // 3296 :  93 - 0x5d -- Background 0x9c
      12'hCE1: dout  = 8'b01011110; // 3297 :  94 - 0x5e
      12'hCE2: dout  = 8'b01011111; // 3298 :  95 - 0x5f
      12'hCE3: dout  = 8'b01011111; // 3299 :  95 - 0x5f
      12'hCE4: dout  = 8'b01011111; // 3300 :  95 - 0x5f
      12'hCE5: dout  = 8'b01011111; // 3301 :  95 - 0x5f
      12'hCE6: dout  = 8'b01011111; // 3302 :  95 - 0x5f
      12'hCE7: dout  = 8'b01011111; // 3303 :  95 - 0x5f
      12'hCE8: dout  = 8'b10000000; // 3304 : 128 - 0x80 -- Background 0x9d
      12'hCE9: dout  = 8'b11000001; // 3305 : 193 - 0xc1
      12'hCEA: dout  = 8'b01100011; // 3306 :  99 - 0x63
      12'hCEB: dout  = 8'b10110110; // 3307 : 182 - 0xb6
      12'hCEC: dout  = 8'b11011001; // 3308 : 217 - 0xd9
      12'hCED: dout  = 8'b11101011; // 3309 : 235 - 0xeb
      12'hCEE: dout  = 8'b11110111; // 3310 : 247 - 0xf7
      12'hCEF: dout  = 8'b11111111; // 3311 : 255 - 0xff
      12'hCF0: dout  = 8'b11011101; // 3312 : 221 - 0xdd -- Background 0x9e
      12'hCF1: dout  = 8'b10111101; // 3313 : 189 - 0xbd
      12'hCF2: dout  = 8'b01111101; // 3314 : 125 - 0x7d
      12'hCF3: dout  = 8'b11111101; // 3315 : 253 - 0xfd
      12'hCF4: dout  = 8'b11111101; // 3316 : 253 - 0xfd
      12'hCF5: dout  = 8'b11111101; // 3317 : 253 - 0xfd
      12'hCF6: dout  = 8'b11111101; // 3318 : 253 - 0xfd
      12'hCF7: dout  = 8'b11111101; // 3319 : 253 - 0xfd
      12'hCF8: dout  = 8'b00000001; // 3320 :   1 - 0x1 -- Background 0x9f
      12'hCF9: dout  = 8'b00000001; // 3321 :   1 - 0x1
      12'hCFA: dout  = 8'b00000010; // 3322 :   2 - 0x2
      12'hCFB: dout  = 8'b00000010; // 3323 :   2 - 0x2
      12'hCFC: dout  = 8'b00000101; // 3324 :   5 - 0x5
      12'hCFD: dout  = 8'b00000101; // 3325 :   5 - 0x5
      12'hCFE: dout  = 8'b00001011; // 3326 :  11 - 0xb
      12'hCFF: dout  = 8'b00001011; // 3327 :  11 - 0xb
      12'hD00: dout  = 8'b01110100; // 3328 : 116 - 0x74 -- Background 0xa0
      12'hD01: dout  = 8'b01110110; // 3329 : 118 - 0x76
      12'hD02: dout  = 8'b11111010; // 3330 : 250 - 0xfa
      12'hD03: dout  = 8'b11111011; // 3331 : 251 - 0xfb
      12'hD04: dout  = 8'b11111101; // 3332 : 253 - 0xfd
      12'hD05: dout  = 8'b11111101; // 3333 : 253 - 0xfd
      12'hD06: dout  = 8'b11111110; // 3334 : 254 - 0xfe
      12'hD07: dout  = 8'b11111110; // 3335 : 254 - 0xfe
      12'hD08: dout  = 8'b00000010; // 3336 :   2 - 0x2 -- Background 0xa1
      12'hD09: dout  = 8'b00000010; // 3337 :   2 - 0x2
      12'hD0A: dout  = 8'b00000010; // 3338 :   2 - 0x2
      12'hD0B: dout  = 8'b00000010; // 3339 :   2 - 0x2
      12'hD0C: dout  = 8'b00000010; // 3340 :   2 - 0x2
      12'hD0D: dout  = 8'b10000010; // 3341 : 130 - 0x82
      12'hD0E: dout  = 8'b10000010; // 3342 : 130 - 0x82
      12'hD0F: dout  = 8'b11000010; // 3343 : 194 - 0xc2
      12'hD10: dout  = 8'b11101010; // 3344 : 234 - 0xea -- Background 0xa2
      12'hD11: dout  = 8'b11110110; // 3345 : 246 - 0xf6
      12'hD12: dout  = 8'b11111010; // 3346 : 250 - 0xfa
      12'hD13: dout  = 8'b11111010; // 3347 : 250 - 0xfa
      12'hD14: dout  = 8'b11111100; // 3348 : 252 - 0xfc
      12'hD15: dout  = 8'b11111100; // 3349 : 252 - 0xfc
      12'hD16: dout  = 8'b11111110; // 3350 : 254 - 0xfe
      12'hD17: dout  = 8'b11111111; // 3351 : 255 - 0xff
      12'hD18: dout  = 8'b11111111; // 3352 : 255 - 0xff -- Background 0xa3
      12'hD19: dout  = 8'b11111111; // 3353 : 255 - 0xff
      12'hD1A: dout  = 8'b11111111; // 3354 : 255 - 0xff
      12'hD1B: dout  = 8'b11111111; // 3355 : 255 - 0xff
      12'hD1C: dout  = 8'b11111111; // 3356 : 255 - 0xff
      12'hD1D: dout  = 8'b11111111; // 3357 : 255 - 0xff
      12'hD1E: dout  = 8'b11111111; // 3358 : 255 - 0xff
      12'hD1F: dout  = 8'b11111111; // 3359 : 255 - 0xff
      12'hD20: dout  = 8'b01000000; // 3360 :  64 - 0x40 -- Background 0xa4
      12'hD21: dout  = 8'b01000000; // 3361 :  64 - 0x40
      12'hD22: dout  = 8'b01000000; // 3362 :  64 - 0x40
      12'hD23: dout  = 8'b01000000; // 3363 :  64 - 0x40
      12'hD24: dout  = 8'b01000000; // 3364 :  64 - 0x40
      12'hD25: dout  = 8'b01000000; // 3365 :  64 - 0x40
      12'hD26: dout  = 8'b01000000; // 3366 :  64 - 0x40
      12'hD27: dout  = 8'b01000000; // 3367 :  64 - 0x40
      12'hD28: dout  = 8'b11111000; // 3368 : 248 - 0xf8 -- Background 0xa5
      12'hD29: dout  = 8'b11111111; // 3369 : 255 - 0xff
      12'hD2A: dout  = 8'b11111111; // 3370 : 255 - 0xff
      12'hD2B: dout  = 8'b11111000; // 3371 : 248 - 0xf8
      12'hD2C: dout  = 8'b11111011; // 3372 : 251 - 0xfb
      12'hD2D: dout  = 8'b11111010; // 3373 : 250 - 0xfa
      12'hD2E: dout  = 8'b11111010; // 3374 : 250 - 0xfa
      12'hD2F: dout  = 8'b11111010; // 3375 : 250 - 0xfa
      12'hD30: dout  = 8'b11111100; // 3376 : 252 - 0xfc -- Background 0xa6
      12'hD31: dout  = 8'b11111010; // 3377 : 250 - 0xfa
      12'hD32: dout  = 8'b11110110; // 3378 : 246 - 0xf6
      12'hD33: dout  = 8'b00001101; // 3379 :  13 - 0xd
      12'hD34: dout  = 8'b11111001; // 3380 : 249 - 0xf9
      12'hD35: dout  = 8'b00000011; // 3381 :   3 - 0x3
      12'hD36: dout  = 8'b00010011; // 3382 :  19 - 0x13
      12'hD37: dout  = 8'b00110111; // 3383 :  55 - 0x37
      12'hD38: dout  = 8'b01111111; // 3384 : 127 - 0x7f -- Background 0xa7
      12'hD39: dout  = 8'b11111001; // 3385 : 249 - 0xf9
      12'hD3A: dout  = 8'b11111001; // 3386 : 249 - 0xf9
      12'hD3B: dout  = 8'b11111111; // 3387 : 255 - 0xff
      12'hD3C: dout  = 8'b11111110; // 3388 : 254 - 0xfe
      12'hD3D: dout  = 8'b11111100; // 3389 : 252 - 0xfc
      12'hD3E: dout  = 8'b11111111; // 3390 : 255 - 0xff
      12'hD3F: dout  = 8'b11111111; // 3391 : 255 - 0xff
      12'hD40: dout  = 8'b11110110; // 3392 : 246 - 0xf6 -- Background 0xa8
      12'hD41: dout  = 8'b11110110; // 3393 : 246 - 0xf6
      12'hD42: dout  = 8'b11111011; // 3394 : 251 - 0xfb
      12'hD43: dout  = 8'b01111011; // 3395 : 123 - 0x7b
      12'hD44: dout  = 8'b11111101; // 3396 : 253 - 0xfd
      12'hD45: dout  = 8'b11110101; // 3397 : 245 - 0xf5
      12'hD46: dout  = 8'b11110110; // 3398 : 246 - 0xf6
      12'hD47: dout  = 8'b11111010; // 3399 : 250 - 0xfa
      12'hD48: dout  = 8'b10111111; // 3400 : 191 - 0xbf -- Background 0xa9
      12'hD49: dout  = 8'b10111111; // 3401 : 191 - 0xbf
      12'hD4A: dout  = 8'b00111111; // 3402 :  63 - 0x3f
      12'hD4B: dout  = 8'b00111111; // 3403 :  63 - 0x3f
      12'hD4C: dout  = 8'b10111111; // 3404 : 191 - 0xbf
      12'hD4D: dout  = 8'b10011111; // 3405 : 159 - 0x9f
      12'hD4E: dout  = 8'b11001111; // 3406 : 207 - 0xcf
      12'hD4F: dout  = 8'b11010111; // 3407 : 215 - 0xd7
      12'hD50: dout  = 8'b11100100; // 3408 : 228 - 0xe4 -- Background 0xaa
      12'hD51: dout  = 8'b11111000; // 3409 : 248 - 0xf8
      12'hD52: dout  = 8'b11111111; // 3410 : 255 - 0xff
      12'hD53: dout  = 8'b11110011; // 3411 : 243 - 0xf3
      12'hD54: dout  = 8'b11111100; // 3412 : 252 - 0xfc
      12'hD55: dout  = 8'b11111111; // 3413 : 255 - 0xff
      12'hD56: dout  = 8'b11111111; // 3414 : 255 - 0xff
      12'hD57: dout  = 8'b11111111; // 3415 : 255 - 0xff
      12'hD58: dout  = 8'b00000000; // 3416 :   0 - 0x0 -- Background 0xab
      12'hD59: dout  = 8'b00000000; // 3417 :   0 - 0x0
      12'hD5A: dout  = 8'b00000000; // 3418 :   0 - 0x0
      12'hD5B: dout  = 8'b11000000; // 3419 : 192 - 0xc0
      12'hD5C: dout  = 8'b11110000; // 3420 : 240 - 0xf0
      12'hD5D: dout  = 8'b00111100; // 3421 :  60 - 0x3c
      12'hD5E: dout  = 8'b11011000; // 3422 : 216 - 0xd8
      12'hD5F: dout  = 8'b10110110; // 3423 : 182 - 0xb6
      12'hD60: dout  = 8'b00001111; // 3424 :  15 - 0xf -- Background 0xac
      12'hD61: dout  = 8'b00001111; // 3425 :  15 - 0xf
      12'hD62: dout  = 8'b00000000; // 3426 :   0 - 0x0
      12'hD63: dout  = 8'b00000011; // 3427 :   3 - 0x3
      12'hD64: dout  = 8'b00000000; // 3428 :   0 - 0x0
      12'hD65: dout  = 8'b00000000; // 3429 :   0 - 0x0
      12'hD66: dout  = 8'b00000000; // 3430 :   0 - 0x0
      12'hD67: dout  = 8'b00000000; // 3431 :   0 - 0x0
      12'hD68: dout  = 8'b11110100; // 3432 : 244 - 0xf4 -- Background 0xad
      12'hD69: dout  = 8'b11110100; // 3433 : 244 - 0xf4
      12'hD6A: dout  = 8'b00000100; // 3434 :   4 - 0x4
      12'hD6B: dout  = 8'b11111100; // 3435 : 252 - 0xfc
      12'hD6C: dout  = 8'b00000000; // 3436 :   0 - 0x0
      12'hD6D: dout  = 8'b00000000; // 3437 :   0 - 0x0
      12'hD6E: dout  = 8'b00000000; // 3438 :   0 - 0x0
      12'hD6F: dout  = 8'b00000000; // 3439 :   0 - 0x0
      12'hD70: dout  = 8'b01011111; // 3440 :  95 - 0x5f -- Background 0xae
      12'hD71: dout  = 8'b01011111; // 3441 :  95 - 0x5f
      12'hD72: dout  = 8'b01011111; // 3442 :  95 - 0x5f
      12'hD73: dout  = 8'b01011111; // 3443 :  95 - 0x5f
      12'hD74: dout  = 8'b01011111; // 3444 :  95 - 0x5f
      12'hD75: dout  = 8'b01011111; // 3445 :  95 - 0x5f
      12'hD76: dout  = 8'b01011111; // 3446 :  95 - 0x5f
      12'hD77: dout  = 8'b01011111; // 3447 :  95 - 0x5f
      12'hD78: dout  = 8'b11111101; // 3448 : 253 - 0xfd -- Background 0xaf
      12'hD79: dout  = 8'b11111101; // 3449 : 253 - 0xfd
      12'hD7A: dout  = 8'b11111101; // 3450 : 253 - 0xfd
      12'hD7B: dout  = 8'b11111101; // 3451 : 253 - 0xfd
      12'hD7C: dout  = 8'b11110101; // 3452 : 245 - 0xf5
      12'hD7D: dout  = 8'b11110101; // 3453 : 245 - 0xf5
      12'hD7E: dout  = 8'b11110101; // 3454 : 245 - 0xf5
      12'hD7F: dout  = 8'b11110101; // 3455 : 245 - 0xf5
      12'hD80: dout  = 8'b00001100; // 3456 :  12 - 0xc -- Background 0xb0
      12'hD81: dout  = 8'b00011100; // 3457 :  28 - 0x1c
      12'hD82: dout  = 8'b00001100; // 3458 :  12 - 0xc
      12'hD83: dout  = 8'b00001100; // 3459 :  12 - 0xc
      12'hD84: dout  = 8'b00001100; // 3460 :  12 - 0xc
      12'hD85: dout  = 8'b00001100; // 3461 :  12 - 0xc
      12'hD86: dout  = 8'b00111111; // 3462 :  63 - 0x3f
      12'hD87: dout  = 8'b00000000; // 3463 :   0 - 0x0
      12'hD88: dout  = 8'b00111110; // 3464 :  62 - 0x3e -- Background 0xb1
      12'hD89: dout  = 8'b01100011; // 3465 :  99 - 0x63
      12'hD8A: dout  = 8'b00000111; // 3466 :   7 - 0x7
      12'hD8B: dout  = 8'b00011110; // 3467 :  30 - 0x1e
      12'hD8C: dout  = 8'b00111100; // 3468 :  60 - 0x3c
      12'hD8D: dout  = 8'b01110000; // 3469 : 112 - 0x70
      12'hD8E: dout  = 8'b01111111; // 3470 : 127 - 0x7f
      12'hD8F: dout  = 8'b00000000; // 3471 :   0 - 0x0
      12'hD90: dout  = 8'b01111110; // 3472 : 126 - 0x7e -- Background 0xb2
      12'hD91: dout  = 8'b01100011; // 3473 :  99 - 0x63
      12'hD92: dout  = 8'b01100011; // 3474 :  99 - 0x63
      12'hD93: dout  = 8'b01100011; // 3475 :  99 - 0x63
      12'hD94: dout  = 8'b01111110; // 3476 : 126 - 0x7e
      12'hD95: dout  = 8'b01100000; // 3477 :  96 - 0x60
      12'hD96: dout  = 8'b01100000; // 3478 :  96 - 0x60
      12'hD97: dout  = 8'b00000000; // 3479 :   0 - 0x0
      12'hD98: dout  = 8'b01100011; // 3480 :  99 - 0x63 -- Background 0xb3
      12'hD99: dout  = 8'b01100011; // 3481 :  99 - 0x63
      12'hD9A: dout  = 8'b01100011; // 3482 :  99 - 0x63
      12'hD9B: dout  = 8'b01100011; // 3483 :  99 - 0x63
      12'hD9C: dout  = 8'b01100011; // 3484 :  99 - 0x63
      12'hD9D: dout  = 8'b01100011; // 3485 :  99 - 0x63
      12'hD9E: dout  = 8'b00111110; // 3486 :  62 - 0x3e
      12'hD9F: dout  = 8'b00000000; // 3487 :   0 - 0x0
      12'hDA0: dout  = 8'b01100011; // 3488 :  99 - 0x63 -- Background 0xb4
      12'hDA1: dout  = 8'b01100011; // 3489 :  99 - 0x63
      12'hDA2: dout  = 8'b01100011; // 3490 :  99 - 0x63
      12'hDA3: dout  = 8'b01111111; // 3491 : 127 - 0x7f
      12'hDA4: dout  = 8'b01100011; // 3492 :  99 - 0x63
      12'hDA5: dout  = 8'b01100011; // 3493 :  99 - 0x63
      12'hDA6: dout  = 8'b01100011; // 3494 :  99 - 0x63
      12'hDA7: dout  = 8'b00000000; // 3495 :   0 - 0x0
      12'hDA8: dout  = 8'b00111111; // 3496 :  63 - 0x3f -- Background 0xb5
      12'hDA9: dout  = 8'b00001100; // 3497 :  12 - 0xc
      12'hDAA: dout  = 8'b00001100; // 3498 :  12 - 0xc
      12'hDAB: dout  = 8'b00001100; // 3499 :  12 - 0xc
      12'hDAC: dout  = 8'b00001100; // 3500 :  12 - 0xc
      12'hDAD: dout  = 8'b00001100; // 3501 :  12 - 0xc
      12'hDAE: dout  = 8'b00111111; // 3502 :  63 - 0x3f
      12'hDAF: dout  = 8'b00000000; // 3503 :   0 - 0x0
      12'hDB0: dout  = 8'b00000000; // 3504 :   0 - 0x0 -- Background 0xb6
      12'hDB1: dout  = 8'b00000000; // 3505 :   0 - 0x0
      12'hDB2: dout  = 8'b00000000; // 3506 :   0 - 0x0
      12'hDB3: dout  = 8'b01111110; // 3507 : 126 - 0x7e
      12'hDB4: dout  = 8'b00000000; // 3508 :   0 - 0x0
      12'hDB5: dout  = 8'b00000000; // 3509 :   0 - 0x0
      12'hDB6: dout  = 8'b00000000; // 3510 :   0 - 0x0
      12'hDB7: dout  = 8'b00000000; // 3511 :   0 - 0x0
      12'hDB8: dout  = 8'b00111100; // 3512 :  60 - 0x3c -- Background 0xb7
      12'hDB9: dout  = 8'b01100110; // 3513 : 102 - 0x66
      12'hDBA: dout  = 8'b01100000; // 3514 :  96 - 0x60
      12'hDBB: dout  = 8'b00111110; // 3515 :  62 - 0x3e
      12'hDBC: dout  = 8'b00000011; // 3516 :   3 - 0x3
      12'hDBD: dout  = 8'b01100011; // 3517 :  99 - 0x63
      12'hDBE: dout  = 8'b00111110; // 3518 :  62 - 0x3e
      12'hDBF: dout  = 8'b00000000; // 3519 :   0 - 0x0
      12'hDC0: dout  = 8'b00011110; // 3520 :  30 - 0x1e -- Background 0xb8
      12'hDC1: dout  = 8'b00110011; // 3521 :  51 - 0x33
      12'hDC2: dout  = 8'b01100000; // 3522 :  96 - 0x60
      12'hDC3: dout  = 8'b01100000; // 3523 :  96 - 0x60
      12'hDC4: dout  = 8'b01100000; // 3524 :  96 - 0x60
      12'hDC5: dout  = 8'b00110011; // 3525 :  51 - 0x33
      12'hDC6: dout  = 8'b00011110; // 3526 :  30 - 0x1e
      12'hDC7: dout  = 8'b00000000; // 3527 :   0 - 0x0
      12'hDC8: dout  = 8'b00111110; // 3528 :  62 - 0x3e -- Background 0xb9
      12'hDC9: dout  = 8'b01100011; // 3529 :  99 - 0x63
      12'hDCA: dout  = 8'b01100011; // 3530 :  99 - 0x63
      12'hDCB: dout  = 8'b01100011; // 3531 :  99 - 0x63
      12'hDCC: dout  = 8'b01100011; // 3532 :  99 - 0x63
      12'hDCD: dout  = 8'b01100011; // 3533 :  99 - 0x63
      12'hDCE: dout  = 8'b00111110; // 3534 :  62 - 0x3e
      12'hDCF: dout  = 8'b00000000; // 3535 :   0 - 0x0
      12'hDD0: dout  = 8'b01111110; // 3536 : 126 - 0x7e -- Background 0xba
      12'hDD1: dout  = 8'b01100011; // 3537 :  99 - 0x63
      12'hDD2: dout  = 8'b01100011; // 3538 :  99 - 0x63
      12'hDD3: dout  = 8'b01100111; // 3539 : 103 - 0x67
      12'hDD4: dout  = 8'b01111100; // 3540 : 124 - 0x7c
      12'hDD5: dout  = 8'b01101110; // 3541 : 110 - 0x6e
      12'hDD6: dout  = 8'b01100111; // 3542 : 103 - 0x67
      12'hDD7: dout  = 8'b00000000; // 3543 :   0 - 0x0
      12'hDD8: dout  = 8'b01111111; // 3544 : 127 - 0x7f -- Background 0xbb
      12'hDD9: dout  = 8'b01100000; // 3545 :  96 - 0x60
      12'hDDA: dout  = 8'b01100000; // 3546 :  96 - 0x60
      12'hDDB: dout  = 8'b01111110; // 3547 : 126 - 0x7e
      12'hDDC: dout  = 8'b01100000; // 3548 :  96 - 0x60
      12'hDDD: dout  = 8'b01100000; // 3549 :  96 - 0x60
      12'hDDE: dout  = 8'b01111111; // 3550 : 127 - 0x7f
      12'hDDF: dout  = 8'b00000000; // 3551 :   0 - 0x0
      12'hDE0: dout  = 8'b00000000; // 3552 :   0 - 0x0 -- Background 0xbc
      12'hDE1: dout  = 8'b00000000; // 3553 :   0 - 0x0
      12'hDE2: dout  = 8'b00000000; // 3554 :   0 - 0x0
      12'hDE3: dout  = 8'b00000000; // 3555 :   0 - 0x0
      12'hDE4: dout  = 8'b00000000; // 3556 :   0 - 0x0
      12'hDE5: dout  = 8'b00000000; // 3557 :   0 - 0x0
      12'hDE6: dout  = 8'b00000000; // 3558 :   0 - 0x0
      12'hDE7: dout  = 8'b00000000; // 3559 :   0 - 0x0
      12'hDE8: dout  = 8'b00000000; // 3560 :   0 - 0x0 -- Background 0xbd
      12'hDE9: dout  = 8'b00000000; // 3561 :   0 - 0x0
      12'hDEA: dout  = 8'b00000000; // 3562 :   0 - 0x0
      12'hDEB: dout  = 8'b00000000; // 3563 :   0 - 0x0
      12'hDEC: dout  = 8'b00000000; // 3564 :   0 - 0x0
      12'hDED: dout  = 8'b00000000; // 3565 :   0 - 0x0
      12'hDEE: dout  = 8'b00000000; // 3566 :   0 - 0x0
      12'hDEF: dout  = 8'b00000000; // 3567 :   0 - 0x0
      12'hDF0: dout  = 8'b00000000; // 3568 :   0 - 0x0 -- Background 0xbe
      12'hDF1: dout  = 8'b00000000; // 3569 :   0 - 0x0
      12'hDF2: dout  = 8'b00000000; // 3570 :   0 - 0x0
      12'hDF3: dout  = 8'b00000000; // 3571 :   0 - 0x0
      12'hDF4: dout  = 8'b00000000; // 3572 :   0 - 0x0
      12'hDF5: dout  = 8'b00000000; // 3573 :   0 - 0x0
      12'hDF6: dout  = 8'b00000000; // 3574 :   0 - 0x0
      12'hDF7: dout  = 8'b00000000; // 3575 :   0 - 0x0
      12'hDF8: dout  = 8'b00000000; // 3576 :   0 - 0x0 -- Background 0xbf
      12'hDF9: dout  = 8'b00000000; // 3577 :   0 - 0x0
      12'hDFA: dout  = 8'b00000000; // 3578 :   0 - 0x0
      12'hDFB: dout  = 8'b00000000; // 3579 :   0 - 0x0
      12'hDFC: dout  = 8'b00000000; // 3580 :   0 - 0x0
      12'hDFD: dout  = 8'b00000000; // 3581 :   0 - 0x0
      12'hDFE: dout  = 8'b00000000; // 3582 :   0 - 0x0
      12'hDFF: dout  = 8'b00000000; // 3583 :   0 - 0x0
      12'hE00: dout  = 8'b01100011; // 3584 :  99 - 0x63 -- Background 0xc0
      12'hE01: dout  = 8'b01100110; // 3585 : 102 - 0x66
      12'hE02: dout  = 8'b01101100; // 3586 : 108 - 0x6c
      12'hE03: dout  = 8'b01111000; // 3587 : 120 - 0x78
      12'hE04: dout  = 8'b01111100; // 3588 : 124 - 0x7c
      12'hE05: dout  = 8'b01100110; // 3589 : 102 - 0x66
      12'hE06: dout  = 8'b01100011; // 3590 :  99 - 0x63
      12'hE07: dout  = 8'b00000000; // 3591 :   0 - 0x0
      12'hE08: dout  = 8'b00111111; // 3592 :  63 - 0x3f -- Background 0xc1
      12'hE09: dout  = 8'b00001100; // 3593 :  12 - 0xc
      12'hE0A: dout  = 8'b00001100; // 3594 :  12 - 0xc
      12'hE0B: dout  = 8'b00001100; // 3595 :  12 - 0xc
      12'hE0C: dout  = 8'b00001100; // 3596 :  12 - 0xc
      12'hE0D: dout  = 8'b00001100; // 3597 :  12 - 0xc
      12'hE0E: dout  = 8'b00111111; // 3598 :  63 - 0x3f
      12'hE0F: dout  = 8'b00000000; // 3599 :   0 - 0x0
      12'hE10: dout  = 8'b01100011; // 3600 :  99 - 0x63 -- Background 0xc2
      12'hE11: dout  = 8'b01110111; // 3601 : 119 - 0x77
      12'hE12: dout  = 8'b01111111; // 3602 : 127 - 0x7f
      12'hE13: dout  = 8'b01111111; // 3603 : 127 - 0x7f
      12'hE14: dout  = 8'b01101011; // 3604 : 107 - 0x6b
      12'hE15: dout  = 8'b01100011; // 3605 :  99 - 0x63
      12'hE16: dout  = 8'b01100011; // 3606 :  99 - 0x63
      12'hE17: dout  = 8'b00000000; // 3607 :   0 - 0x0
      12'hE18: dout  = 8'b00011100; // 3608 :  28 - 0x1c -- Background 0xc3
      12'hE19: dout  = 8'b00110110; // 3609 :  54 - 0x36
      12'hE1A: dout  = 8'b01100011; // 3610 :  99 - 0x63
      12'hE1B: dout  = 8'b01100011; // 3611 :  99 - 0x63
      12'hE1C: dout  = 8'b01111111; // 3612 : 127 - 0x7f
      12'hE1D: dout  = 8'b01100011; // 3613 :  99 - 0x63
      12'hE1E: dout  = 8'b01100011; // 3614 :  99 - 0x63
      12'hE1F: dout  = 8'b00000000; // 3615 :   0 - 0x0
      12'hE20: dout  = 8'b00011111; // 3616 :  31 - 0x1f -- Background 0xc4
      12'hE21: dout  = 8'b00110000; // 3617 :  48 - 0x30
      12'hE22: dout  = 8'b01100000; // 3618 :  96 - 0x60
      12'hE23: dout  = 8'b01100111; // 3619 : 103 - 0x67
      12'hE24: dout  = 8'b01100011; // 3620 :  99 - 0x63
      12'hE25: dout  = 8'b00110011; // 3621 :  51 - 0x33
      12'hE26: dout  = 8'b00011111; // 3622 :  31 - 0x1f
      12'hE27: dout  = 8'b00000000; // 3623 :   0 - 0x0
      12'hE28: dout  = 8'b01100011; // 3624 :  99 - 0x63 -- Background 0xc5
      12'hE29: dout  = 8'b01100011; // 3625 :  99 - 0x63
      12'hE2A: dout  = 8'b01100011; // 3626 :  99 - 0x63
      12'hE2B: dout  = 8'b01100011; // 3627 :  99 - 0x63
      12'hE2C: dout  = 8'b01100011; // 3628 :  99 - 0x63
      12'hE2D: dout  = 8'b01100011; // 3629 :  99 - 0x63
      12'hE2E: dout  = 8'b00111110; // 3630 :  62 - 0x3e
      12'hE2F: dout  = 8'b00000000; // 3631 :   0 - 0x0
      12'hE30: dout  = 8'b01111110; // 3632 : 126 - 0x7e -- Background 0xc6
      12'hE31: dout  = 8'b01100011; // 3633 :  99 - 0x63
      12'hE32: dout  = 8'b01100011; // 3634 :  99 - 0x63
      12'hE33: dout  = 8'b01100111; // 3635 : 103 - 0x67
      12'hE34: dout  = 8'b01111100; // 3636 : 124 - 0x7c
      12'hE35: dout  = 8'b01101110; // 3637 : 110 - 0x6e
      12'hE36: dout  = 8'b01100111; // 3638 : 103 - 0x67
      12'hE37: dout  = 8'b00000000; // 3639 :   0 - 0x0
      12'hE38: dout  = 8'b01111111; // 3640 : 127 - 0x7f -- Background 0xc7
      12'hE39: dout  = 8'b01100000; // 3641 :  96 - 0x60
      12'hE3A: dout  = 8'b01100000; // 3642 :  96 - 0x60
      12'hE3B: dout  = 8'b01111110; // 3643 : 126 - 0x7e
      12'hE3C: dout  = 8'b01100000; // 3644 :  96 - 0x60
      12'hE3D: dout  = 8'b01100000; // 3645 :  96 - 0x60
      12'hE3E: dout  = 8'b01111111; // 3646 : 127 - 0x7f
      12'hE3F: dout  = 8'b00000000; // 3647 :   0 - 0x0
      12'hE40: dout  = 8'b00110110; // 3648 :  54 - 0x36 -- Background 0xc8
      12'hE41: dout  = 8'b00110110; // 3649 :  54 - 0x36
      12'hE42: dout  = 8'b00010010; // 3650 :  18 - 0x12
      12'hE43: dout  = 8'b00000000; // 3651 :   0 - 0x0
      12'hE44: dout  = 8'b00000000; // 3652 :   0 - 0x0
      12'hE45: dout  = 8'b00000000; // 3653 :   0 - 0x0
      12'hE46: dout  = 8'b00000000; // 3654 :   0 - 0x0
      12'hE47: dout  = 8'b00000000; // 3655 :   0 - 0x0
      12'hE48: dout  = 8'b00111110; // 3656 :  62 - 0x3e -- Background 0xc9
      12'hE49: dout  = 8'b01100011; // 3657 :  99 - 0x63
      12'hE4A: dout  = 8'b01100011; // 3658 :  99 - 0x63
      12'hE4B: dout  = 8'b01100011; // 3659 :  99 - 0x63
      12'hE4C: dout  = 8'b01100011; // 3660 :  99 - 0x63
      12'hE4D: dout  = 8'b01100011; // 3661 :  99 - 0x63
      12'hE4E: dout  = 8'b00111110; // 3662 :  62 - 0x3e
      12'hE4F: dout  = 8'b00000000; // 3663 :   0 - 0x0
      12'hE50: dout  = 8'b00111100; // 3664 :  60 - 0x3c -- Background 0xca
      12'hE51: dout  = 8'b01100110; // 3665 : 102 - 0x66
      12'hE52: dout  = 8'b01100000; // 3666 :  96 - 0x60
      12'hE53: dout  = 8'b00111110; // 3667 :  62 - 0x3e
      12'hE54: dout  = 8'b00000011; // 3668 :   3 - 0x3
      12'hE55: dout  = 8'b01100011; // 3669 :  99 - 0x63
      12'hE56: dout  = 8'b00111110; // 3670 :  62 - 0x3e
      12'hE57: dout  = 8'b00000000; // 3671 :   0 - 0x0
      12'hE58: dout  = 8'b00000000; // 3672 :   0 - 0x0 -- Background 0xcb
      12'hE59: dout  = 8'b00111000; // 3673 :  56 - 0x38
      12'hE5A: dout  = 8'b01111100; // 3674 : 124 - 0x7c
      12'hE5B: dout  = 8'b11111110; // 3675 : 254 - 0xfe
      12'hE5C: dout  = 8'b11111110; // 3676 : 254 - 0xfe
      12'hE5D: dout  = 8'b11111110; // 3677 : 254 - 0xfe
      12'hE5E: dout  = 8'b01111100; // 3678 : 124 - 0x7c
      12'hE5F: dout  = 8'b00111000; // 3679 :  56 - 0x38
      12'hE60: dout  = 8'b00000000; // 3680 :   0 - 0x0 -- Background 0xcc
      12'hE61: dout  = 8'b00000000; // 3681 :   0 - 0x0
      12'hE62: dout  = 8'b00000000; // 3682 :   0 - 0x0
      12'hE63: dout  = 8'b00000000; // 3683 :   0 - 0x0
      12'hE64: dout  = 8'b00000000; // 3684 :   0 - 0x0
      12'hE65: dout  = 8'b00000000; // 3685 :   0 - 0x0
      12'hE66: dout  = 8'b00000000; // 3686 :   0 - 0x0
      12'hE67: dout  = 8'b00000000; // 3687 :   0 - 0x0
      12'hE68: dout  = 8'b00000000; // 3688 :   0 - 0x0 -- Background 0xcd
      12'hE69: dout  = 8'b00000000; // 3689 :   0 - 0x0
      12'hE6A: dout  = 8'b00000000; // 3690 :   0 - 0x0
      12'hE6B: dout  = 8'b00000000; // 3691 :   0 - 0x0
      12'hE6C: dout  = 8'b00000000; // 3692 :   0 - 0x0
      12'hE6D: dout  = 8'b00000000; // 3693 :   0 - 0x0
      12'hE6E: dout  = 8'b00000000; // 3694 :   0 - 0x0
      12'hE6F: dout  = 8'b00000000; // 3695 :   0 - 0x0
      12'hE70: dout  = 8'b00000000; // 3696 :   0 - 0x0 -- Background 0xce
      12'hE71: dout  = 8'b00000000; // 3697 :   0 - 0x0
      12'hE72: dout  = 8'b00000000; // 3698 :   0 - 0x0
      12'hE73: dout  = 8'b00000000; // 3699 :   0 - 0x0
      12'hE74: dout  = 8'b00000000; // 3700 :   0 - 0x0
      12'hE75: dout  = 8'b00000000; // 3701 :   0 - 0x0
      12'hE76: dout  = 8'b00000000; // 3702 :   0 - 0x0
      12'hE77: dout  = 8'b00000000; // 3703 :   0 - 0x0
      12'hE78: dout  = 8'b00000000; // 3704 :   0 - 0x0 -- Background 0xcf
      12'hE79: dout  = 8'b00000000; // 3705 :   0 - 0x0
      12'hE7A: dout  = 8'b00000000; // 3706 :   0 - 0x0
      12'hE7B: dout  = 8'b00000000; // 3707 :   0 - 0x0
      12'hE7C: dout  = 8'b00000000; // 3708 :   0 - 0x0
      12'hE7D: dout  = 8'b00000000; // 3709 :   0 - 0x0
      12'hE7E: dout  = 8'b00000000; // 3710 :   0 - 0x0
      12'hE7F: dout  = 8'b00000000; // 3711 :   0 - 0x0
      12'hE80: dout  = 8'b00010111; // 3712 :  23 - 0x17 -- Background 0xd0
      12'hE81: dout  = 8'b00010111; // 3713 :  23 - 0x17
      12'hE82: dout  = 8'b00101111; // 3714 :  47 - 0x2f
      12'hE83: dout  = 8'b00101111; // 3715 :  47 - 0x2f
      12'hE84: dout  = 8'b01011111; // 3716 :  95 - 0x5f
      12'hE85: dout  = 8'b01011111; // 3717 :  95 - 0x5f
      12'hE86: dout  = 8'b00111111; // 3718 :  63 - 0x3f
      12'hE87: dout  = 8'b00111111; // 3719 :  63 - 0x3f
      12'hE88: dout  = 8'b11111111; // 3720 : 255 - 0xff -- Background 0xd1
      12'hE89: dout  = 8'b11001111; // 3721 : 207 - 0xcf
      12'hE8A: dout  = 8'b11001111; // 3722 : 207 - 0xcf
      12'hE8B: dout  = 8'b11111011; // 3723 : 251 - 0xfb
      12'hE8C: dout  = 8'b11110111; // 3724 : 247 - 0xf7
      12'hE8D: dout  = 8'b11100111; // 3725 : 231 - 0xe7
      12'hE8E: dout  = 8'b11111111; // 3726 : 255 - 0xff
      12'hE8F: dout  = 8'b11111111; // 3727 : 255 - 0xff
      12'hE90: dout  = 8'b01000010; // 3728 :  66 - 0x42 -- Background 0xd2
      12'hE91: dout  = 8'b01100010; // 3729 :  98 - 0x62
      12'hE92: dout  = 8'b10100010; // 3730 : 162 - 0xa2
      12'hE93: dout  = 8'b10110010; // 3731 : 178 - 0xb2
      12'hE94: dout  = 8'b01010010; // 3732 :  82 - 0x52
      12'hE95: dout  = 8'b01011010; // 3733 :  90 - 0x5a
      12'hE96: dout  = 8'b10101010; // 3734 : 170 - 0xaa
      12'hE97: dout  = 8'b10101100; // 3735 : 172 - 0xac
      12'hE98: dout  = 8'b11111111; // 3736 : 255 - 0xff -- Background 0xd3
      12'hE99: dout  = 8'b11111111; // 3737 : 255 - 0xff
      12'hE9A: dout  = 8'b11111111; // 3738 : 255 - 0xff
      12'hE9B: dout  = 8'b11111111; // 3739 : 255 - 0xff
      12'hE9C: dout  = 8'b11111101; // 3740 : 253 - 0xfd
      12'hE9D: dout  = 8'b11111101; // 3741 : 253 - 0xfd
      12'hE9E: dout  = 8'b11111101; // 3742 : 253 - 0xfd
      12'hE9F: dout  = 8'b11111101; // 3743 : 253 - 0xfd
      12'hEA0: dout  = 8'b00000111; // 3744 :   7 - 0x7 -- Background 0xd4
      12'hEA1: dout  = 8'b00000111; // 3745 :   7 - 0x7
      12'hEA2: dout  = 8'b00000000; // 3746 :   0 - 0x0
      12'hEA3: dout  = 8'b00000011; // 3747 :   3 - 0x3
      12'hEA4: dout  = 8'b00000000; // 3748 :   0 - 0x0
      12'hEA5: dout  = 8'b00000000; // 3749 :   0 - 0x0
      12'hEA6: dout  = 8'b00000000; // 3750 :   0 - 0x0
      12'hEA7: dout  = 8'b00000000; // 3751 :   0 - 0x0
      12'hEA8: dout  = 8'b11111010; // 3752 : 250 - 0xfa -- Background 0xd5
      12'hEA9: dout  = 8'b11111010; // 3753 : 250 - 0xfa
      12'hEAA: dout  = 8'b00000010; // 3754 :   2 - 0x2
      12'hEAB: dout  = 8'b11111110; // 3755 : 254 - 0xfe
      12'hEAC: dout  = 8'b00000000; // 3756 :   0 - 0x0
      12'hEAD: dout  = 8'b00000000; // 3757 :   0 - 0x0
      12'hEAE: dout  = 8'b00000000; // 3758 :   0 - 0x0
      12'hEAF: dout  = 8'b00000000; // 3759 :   0 - 0x0
      12'hEB0: dout  = 8'b00001111; // 3760 :  15 - 0xf -- Background 0xd6
      12'hEB1: dout  = 8'b00001111; // 3761 :  15 - 0xf
      12'hEB2: dout  = 8'b00000000; // 3762 :   0 - 0x0
      12'hEB3: dout  = 8'b00000111; // 3763 :   7 - 0x7
      12'hEB4: dout  = 8'b00000000; // 3764 :   0 - 0x0
      12'hEB5: dout  = 8'b00000000; // 3765 :   0 - 0x0
      12'hEB6: dout  = 8'b00000000; // 3766 :   0 - 0x0
      12'hEB7: dout  = 8'b00000000; // 3767 :   0 - 0x0
      12'hEB8: dout  = 8'b11111111; // 3768 : 255 - 0xff -- Background 0xd7
      12'hEB9: dout  = 8'b11111111; // 3769 : 255 - 0xff
      12'hEBA: dout  = 8'b00000000; // 3770 :   0 - 0x0
      12'hEBB: dout  = 8'b11111111; // 3771 : 255 - 0xff
      12'hEBC: dout  = 8'b00000000; // 3772 :   0 - 0x0
      12'hEBD: dout  = 8'b00000000; // 3773 :   0 - 0x0
      12'hEBE: dout  = 8'b00000000; // 3774 :   0 - 0x0
      12'hEBF: dout  = 8'b00000000; // 3775 :   0 - 0x0
      12'hEC0: dout  = 8'b11000011; // 3776 : 195 - 0xc3 -- Background 0xd8
      12'hEC1: dout  = 8'b11111111; // 3777 : 255 - 0xff
      12'hEC2: dout  = 8'b00000000; // 3778 :   0 - 0x0
      12'hEC3: dout  = 8'b11111111; // 3779 : 255 - 0xff
      12'hEC4: dout  = 8'b00000000; // 3780 :   0 - 0x0
      12'hEC5: dout  = 8'b00000000; // 3781 :   0 - 0x0
      12'hEC6: dout  = 8'b00000000; // 3782 :   0 - 0x0
      12'hEC7: dout  = 8'b00000000; // 3783 :   0 - 0x0
      12'hEC8: dout  = 8'b01101011; // 3784 : 107 - 0x6b -- Background 0xd9
      12'hEC9: dout  = 8'b10110101; // 3785 : 181 - 0xb5
      12'hECA: dout  = 8'b00110110; // 3786 :  54 - 0x36
      12'hECB: dout  = 8'b11111000; // 3787 : 248 - 0xf8
      12'hECC: dout  = 8'b00000000; // 3788 :   0 - 0x0
      12'hECD: dout  = 8'b00000000; // 3789 :   0 - 0x0
      12'hECE: dout  = 8'b00000000; // 3790 :   0 - 0x0
      12'hECF: dout  = 8'b00000000; // 3791 :   0 - 0x0
      12'hED0: dout  = 8'b11111111; // 3792 : 255 - 0xff -- Background 0xda
      12'hED1: dout  = 8'b11111111; // 3793 : 255 - 0xff
      12'hED2: dout  = 8'b01111110; // 3794 : 126 - 0x7e
      12'hED3: dout  = 8'b10000001; // 3795 : 129 - 0x81
      12'hED4: dout  = 8'b00011111; // 3796 :  31 - 0x1f
      12'hED5: dout  = 8'b00000000; // 3797 :   0 - 0x0
      12'hED6: dout  = 8'b00000000; // 3798 :   0 - 0x0
      12'hED7: dout  = 8'b00000000; // 3799 :   0 - 0x0
      12'hED8: dout  = 8'b01101100; // 3800 : 108 - 0x6c -- Background 0xdb
      12'hED9: dout  = 8'b11011000; // 3801 : 216 - 0xd8
      12'hEDA: dout  = 8'b00110000; // 3802 :  48 - 0x30
      12'hEDB: dout  = 8'b11100000; // 3803 : 224 - 0xe0
      12'hEDC: dout  = 8'b10000000; // 3804 : 128 - 0x80
      12'hEDD: dout  = 8'b00000000; // 3805 :   0 - 0x0
      12'hEDE: dout  = 8'b00000000; // 3806 :   0 - 0x0
      12'hEDF: dout  = 8'b00000000; // 3807 :   0 - 0x0
      12'hEE0: dout  = 8'b00011111; // 3808 :  31 - 0x1f -- Background 0xdc
      12'hEE1: dout  = 8'b00011111; // 3809 :  31 - 0x1f
      12'hEE2: dout  = 8'b00000000; // 3810 :   0 - 0x0
      12'hEE3: dout  = 8'b00000111; // 3811 :   7 - 0x7
      12'hEE4: dout  = 8'b00000000; // 3812 :   0 - 0x0
      12'hEE5: dout  = 8'b00000000; // 3813 :   0 - 0x0
      12'hEE6: dout  = 8'b00000000; // 3814 :   0 - 0x0
      12'hEE7: dout  = 8'b00000000; // 3815 :   0 - 0x0
      12'hEE8: dout  = 8'b10000101; // 3816 : 133 - 0x85 -- Background 0xdd
      12'hEE9: dout  = 8'b11111101; // 3817 : 253 - 0xfd
      12'hEEA: dout  = 8'b00000001; // 3818 :   1 - 0x1
      12'hEEB: dout  = 8'b11111111; // 3819 : 255 - 0xff
      12'hEEC: dout  = 8'b00000000; // 3820 :   0 - 0x0
      12'hEED: dout  = 8'b00000000; // 3821 :   0 - 0x0
      12'hEEE: dout  = 8'b00000000; // 3822 :   0 - 0x0
      12'hEEF: dout  = 8'b00000000; // 3823 :   0 - 0x0
      12'hEF0: dout  = 8'b01111111; // 3824 : 127 - 0x7f -- Background 0xde
      12'hEF1: dout  = 8'b01111111; // 3825 : 127 - 0x7f
      12'hEF2: dout  = 8'b00000000; // 3826 :   0 - 0x0
      12'hEF3: dout  = 8'b01011111; // 3827 :  95 - 0x5f
      12'hEF4: dout  = 8'b00000000; // 3828 :   0 - 0x0
      12'hEF5: dout  = 8'b00000000; // 3829 :   0 - 0x0
      12'hEF6: dout  = 8'b00000000; // 3830 :   0 - 0x0
      12'hEF7: dout  = 8'b00000000; // 3831 :   0 - 0x0
      12'hEF8: dout  = 8'b11111100; // 3832 : 252 - 0xfc -- Background 0xdf
      12'hEF9: dout  = 8'b11111111; // 3833 : 255 - 0xff
      12'hEFA: dout  = 8'b00000000; // 3834 :   0 - 0x0
      12'hEFB: dout  = 8'b11111111; // 3835 : 255 - 0xff
      12'hEFC: dout  = 8'b00000000; // 3836 :   0 - 0x0
      12'hEFD: dout  = 8'b00000000; // 3837 :   0 - 0x0
      12'hEFE: dout  = 8'b00000000; // 3838 :   0 - 0x0
      12'hEFF: dout  = 8'b00000000; // 3839 :   0 - 0x0
      12'hF00: dout  = 8'b00110100; // 3840 :  52 - 0x34 -- Background 0xe0
      12'hF01: dout  = 8'b11110110; // 3841 : 246 - 0xf6
      12'hF02: dout  = 8'b00000010; // 3842 :   2 - 0x2
      12'hF03: dout  = 8'b11111111; // 3843 : 255 - 0xff
      12'hF04: dout  = 8'b00000000; // 3844 :   0 - 0x0
      12'hF05: dout  = 8'b00000000; // 3845 :   0 - 0x0
      12'hF06: dout  = 8'b00000000; // 3846 :   0 - 0x0
      12'hF07: dout  = 8'b00000000; // 3847 :   0 - 0x0
      12'hF08: dout  = 8'b11111111; // 3848 : 255 - 0xff -- Background 0xe1
      12'hF09: dout  = 8'b11111111; // 3849 : 255 - 0xff
      12'hF0A: dout  = 8'b00000000; // 3850 :   0 - 0x0
      12'hF0B: dout  = 8'b01111111; // 3851 : 127 - 0x7f
      12'hF0C: dout  = 8'b00000000; // 3852 :   0 - 0x0
      12'hF0D: dout  = 8'b00000000; // 3853 :   0 - 0x0
      12'hF0E: dout  = 8'b00000000; // 3854 :   0 - 0x0
      12'hF0F: dout  = 8'b00000000; // 3855 :   0 - 0x0
      12'hF10: dout  = 8'b11100001; // 3856 : 225 - 0xe1 -- Background 0xe2
      12'hF11: dout  = 8'b11111111; // 3857 : 255 - 0xff
      12'hF12: dout  = 8'b00000000; // 3858 :   0 - 0x0
      12'hF13: dout  = 8'b11111111; // 3859 : 255 - 0xff
      12'hF14: dout  = 8'b00000000; // 3860 :   0 - 0x0
      12'hF15: dout  = 8'b00000000; // 3861 :   0 - 0x0
      12'hF16: dout  = 8'b00000000; // 3862 :   0 - 0x0
      12'hF17: dout  = 8'b00000000; // 3863 :   0 - 0x0
      12'hF18: dout  = 8'b01000000; // 3864 :  64 - 0x40 -- Background 0xe3
      12'hF19: dout  = 8'b01000000; // 3865 :  64 - 0x40
      12'hF1A: dout  = 8'b01000000; // 3866 :  64 - 0x40
      12'hF1B: dout  = 8'b11000000; // 3867 : 192 - 0xc0
      12'hF1C: dout  = 8'b00000000; // 3868 :   0 - 0x0
      12'hF1D: dout  = 8'b00000000; // 3869 :   0 - 0x0
      12'hF1E: dout  = 8'b00000000; // 3870 :   0 - 0x0
      12'hF1F: dout  = 8'b00000000; // 3871 :   0 - 0x0
      12'hF20: dout  = 8'b00000000; // 3872 :   0 - 0x0 -- Background 0xe4
      12'hF21: dout  = 8'b00000000; // 3873 :   0 - 0x0
      12'hF22: dout  = 8'b00000000; // 3874 :   0 - 0x0
      12'hF23: dout  = 8'b00000000; // 3875 :   0 - 0x0
      12'hF24: dout  = 8'b00000111; // 3876 :   7 - 0x7
      12'hF25: dout  = 8'b00001111; // 3877 :  15 - 0xf
      12'hF26: dout  = 8'b00001111; // 3878 :  15 - 0xf
      12'hF27: dout  = 8'b00001111; // 3879 :  15 - 0xf
      12'hF28: dout  = 8'b00000000; // 3880 :   0 - 0x0 -- Background 0xe5
      12'hF29: dout  = 8'b00000000; // 3881 :   0 - 0x0
      12'hF2A: dout  = 8'b00000000; // 3882 :   0 - 0x0
      12'hF2B: dout  = 8'b00000000; // 3883 :   0 - 0x0
      12'hF2C: dout  = 8'b11100000; // 3884 : 224 - 0xe0
      12'hF2D: dout  = 8'b11110000; // 3885 : 240 - 0xf0
      12'hF2E: dout  = 8'b11110000; // 3886 : 240 - 0xf0
      12'hF2F: dout  = 8'b11110000; // 3887 : 240 - 0xf0
      12'hF30: dout  = 8'b11110000; // 3888 : 240 - 0xf0 -- Background 0xe6
      12'hF31: dout  = 8'b11110000; // 3889 : 240 - 0xf0
      12'hF32: dout  = 8'b11110000; // 3890 : 240 - 0xf0
      12'hF33: dout  = 8'b11100000; // 3891 : 224 - 0xe0
      12'hF34: dout  = 8'b00000000; // 3892 :   0 - 0x0
      12'hF35: dout  = 8'b00000000; // 3893 :   0 - 0x0
      12'hF36: dout  = 8'b00000000; // 3894 :   0 - 0x0
      12'hF37: dout  = 8'b00000000; // 3895 :   0 - 0x0
      12'hF38: dout  = 8'b00001111; // 3896 :  15 - 0xf -- Background 0xe7
      12'hF39: dout  = 8'b00001111; // 3897 :  15 - 0xf
      12'hF3A: dout  = 8'b00001111; // 3898 :  15 - 0xf
      12'hF3B: dout  = 8'b00000111; // 3899 :   7 - 0x7
      12'hF3C: dout  = 8'b00000000; // 3900 :   0 - 0x0
      12'hF3D: dout  = 8'b00000000; // 3901 :   0 - 0x0
      12'hF3E: dout  = 8'b00000000; // 3902 :   0 - 0x0
      12'hF3F: dout  = 8'b00000000; // 3903 :   0 - 0x0
      12'hF40: dout  = 8'b00000000; // 3904 :   0 - 0x0 -- Background 0xe8
      12'hF41: dout  = 8'b00000000; // 3905 :   0 - 0x0
      12'hF42: dout  = 8'b00000000; // 3906 :   0 - 0x0
      12'hF43: dout  = 8'b00000000; // 3907 :   0 - 0x0
      12'hF44: dout  = 8'b11111111; // 3908 : 255 - 0xff
      12'hF45: dout  = 8'b11111111; // 3909 : 255 - 0xff
      12'hF46: dout  = 8'b11111111; // 3910 : 255 - 0xff
      12'hF47: dout  = 8'b11111111; // 3911 : 255 - 0xff
      12'hF48: dout  = 8'b11110000; // 3912 : 240 - 0xf0 -- Background 0xe9
      12'hF49: dout  = 8'b11110000; // 3913 : 240 - 0xf0
      12'hF4A: dout  = 8'b11110000; // 3914 : 240 - 0xf0
      12'hF4B: dout  = 8'b11110000; // 3915 : 240 - 0xf0
      12'hF4C: dout  = 8'b11110000; // 3916 : 240 - 0xf0
      12'hF4D: dout  = 8'b11110000; // 3917 : 240 - 0xf0
      12'hF4E: dout  = 8'b11110000; // 3918 : 240 - 0xf0
      12'hF4F: dout  = 8'b11110000; // 3919 : 240 - 0xf0
      12'hF50: dout  = 8'b11111111; // 3920 : 255 - 0xff -- Background 0xea
      12'hF51: dout  = 8'b11111111; // 3921 : 255 - 0xff
      12'hF52: dout  = 8'b11111111; // 3922 : 255 - 0xff
      12'hF53: dout  = 8'b11111111; // 3923 : 255 - 0xff
      12'hF54: dout  = 8'b00000000; // 3924 :   0 - 0x0
      12'hF55: dout  = 8'b00000000; // 3925 :   0 - 0x0
      12'hF56: dout  = 8'b00000000; // 3926 :   0 - 0x0
      12'hF57: dout  = 8'b00000000; // 3927 :   0 - 0x0
      12'hF58: dout  = 8'b00001111; // 3928 :  15 - 0xf -- Background 0xeb
      12'hF59: dout  = 8'b00001111; // 3929 :  15 - 0xf
      12'hF5A: dout  = 8'b00001111; // 3930 :  15 - 0xf
      12'hF5B: dout  = 8'b00001111; // 3931 :  15 - 0xf
      12'hF5C: dout  = 8'b00001111; // 3932 :  15 - 0xf
      12'hF5D: dout  = 8'b00001111; // 3933 :  15 - 0xf
      12'hF5E: dout  = 8'b00001111; // 3934 :  15 - 0xf
      12'hF5F: dout  = 8'b00001111; // 3935 :  15 - 0xf
      12'hF60: dout  = 8'b00000000; // 3936 :   0 - 0x0 -- Background 0xec
      12'hF61: dout  = 8'b00000000; // 3937 :   0 - 0x0
      12'hF62: dout  = 8'b00000000; // 3938 :   0 - 0x0
      12'hF63: dout  = 8'b00000000; // 3939 :   0 - 0x0
      12'hF64: dout  = 8'b00000000; // 3940 :   0 - 0x0
      12'hF65: dout  = 8'b00000000; // 3941 :   0 - 0x0
      12'hF66: dout  = 8'b00000000; // 3942 :   0 - 0x0
      12'hF67: dout  = 8'b00000000; // 3943 :   0 - 0x0
      12'hF68: dout  = 8'b00000000; // 3944 :   0 - 0x0 -- Background 0xed
      12'hF69: dout  = 8'b00000000; // 3945 :   0 - 0x0
      12'hF6A: dout  = 8'b00000000; // 3946 :   0 - 0x0
      12'hF6B: dout  = 8'b00000000; // 3947 :   0 - 0x0
      12'hF6C: dout  = 8'b00000000; // 3948 :   0 - 0x0
      12'hF6D: dout  = 8'b00000000; // 3949 :   0 - 0x0
      12'hF6E: dout  = 8'b00000000; // 3950 :   0 - 0x0
      12'hF6F: dout  = 8'b00000000; // 3951 :   0 - 0x0
      12'hF70: dout  = 8'b00000000; // 3952 :   0 - 0x0 -- Background 0xee
      12'hF71: dout  = 8'b00000000; // 3953 :   0 - 0x0
      12'hF72: dout  = 8'b00000000; // 3954 :   0 - 0x0
      12'hF73: dout  = 8'b00000000; // 3955 :   0 - 0x0
      12'hF74: dout  = 8'b00000000; // 3956 :   0 - 0x0
      12'hF75: dout  = 8'b00000000; // 3957 :   0 - 0x0
      12'hF76: dout  = 8'b00000000; // 3958 :   0 - 0x0
      12'hF77: dout  = 8'b00000000; // 3959 :   0 - 0x0
      12'hF78: dout  = 8'b00000000; // 3960 :   0 - 0x0 -- Background 0xef
      12'hF79: dout  = 8'b00000000; // 3961 :   0 - 0x0
      12'hF7A: dout  = 8'b00000000; // 3962 :   0 - 0x0
      12'hF7B: dout  = 8'b00000000; // 3963 :   0 - 0x0
      12'hF7C: dout  = 8'b00000000; // 3964 :   0 - 0x0
      12'hF7D: dout  = 8'b00000000; // 3965 :   0 - 0x0
      12'hF7E: dout  = 8'b00000000; // 3966 :   0 - 0x0
      12'hF7F: dout  = 8'b00000000; // 3967 :   0 - 0x0
      12'hF80: dout  = 8'b11111111; // 3968 : 255 - 0xff -- Background 0xf0
      12'hF81: dout  = 8'b11111111; // 3969 : 255 - 0xff
      12'hF82: dout  = 8'b11111111; // 3970 : 255 - 0xff
      12'hF83: dout  = 8'b11111111; // 3971 : 255 - 0xff
      12'hF84: dout  = 8'b11111111; // 3972 : 255 - 0xff
      12'hF85: dout  = 8'b11111111; // 3973 : 255 - 0xff
      12'hF86: dout  = 8'b11111111; // 3974 : 255 - 0xff
      12'hF87: dout  = 8'b11111111; // 3975 : 255 - 0xff
      12'hF88: dout  = 8'b11111111; // 3976 : 255 - 0xff -- Background 0xf1
      12'hF89: dout  = 8'b11111111; // 3977 : 255 - 0xff
      12'hF8A: dout  = 8'b11111111; // 3978 : 255 - 0xff
      12'hF8B: dout  = 8'b11111111; // 3979 : 255 - 0xff
      12'hF8C: dout  = 8'b11111111; // 3980 : 255 - 0xff
      12'hF8D: dout  = 8'b11111111; // 3981 : 255 - 0xff
      12'hF8E: dout  = 8'b11111111; // 3982 : 255 - 0xff
      12'hF8F: dout  = 8'b11111111; // 3983 : 255 - 0xff
      12'hF90: dout  = 8'b11111111; // 3984 : 255 - 0xff -- Background 0xf2
      12'hF91: dout  = 8'b11111111; // 3985 : 255 - 0xff
      12'hF92: dout  = 8'b11111111; // 3986 : 255 - 0xff
      12'hF93: dout  = 8'b11111111; // 3987 : 255 - 0xff
      12'hF94: dout  = 8'b11111111; // 3988 : 255 - 0xff
      12'hF95: dout  = 8'b11111111; // 3989 : 255 - 0xff
      12'hF96: dout  = 8'b11111111; // 3990 : 255 - 0xff
      12'hF97: dout  = 8'b11111111; // 3991 : 255 - 0xff
      12'hF98: dout  = 8'b11111111; // 3992 : 255 - 0xff -- Background 0xf3
      12'hF99: dout  = 8'b11111111; // 3993 : 255 - 0xff
      12'hF9A: dout  = 8'b11111111; // 3994 : 255 - 0xff
      12'hF9B: dout  = 8'b11111111; // 3995 : 255 - 0xff
      12'hF9C: dout  = 8'b11111111; // 3996 : 255 - 0xff
      12'hF9D: dout  = 8'b11111111; // 3997 : 255 - 0xff
      12'hF9E: dout  = 8'b11111111; // 3998 : 255 - 0xff
      12'hF9F: dout  = 8'b11111111; // 3999 : 255 - 0xff
      12'hFA0: dout  = 8'b11111111; // 4000 : 255 - 0xff -- Background 0xf4
      12'hFA1: dout  = 8'b11111111; // 4001 : 255 - 0xff
      12'hFA2: dout  = 8'b11111111; // 4002 : 255 - 0xff
      12'hFA3: dout  = 8'b11111111; // 4003 : 255 - 0xff
      12'hFA4: dout  = 8'b11111111; // 4004 : 255 - 0xff
      12'hFA5: dout  = 8'b11111111; // 4005 : 255 - 0xff
      12'hFA6: dout  = 8'b11111111; // 4006 : 255 - 0xff
      12'hFA7: dout  = 8'b11111111; // 4007 : 255 - 0xff
      12'hFA8: dout  = 8'b11111111; // 4008 : 255 - 0xff -- Background 0xf5
      12'hFA9: dout  = 8'b11111111; // 4009 : 255 - 0xff
      12'hFAA: dout  = 8'b11111111; // 4010 : 255 - 0xff
      12'hFAB: dout  = 8'b11111111; // 4011 : 255 - 0xff
      12'hFAC: dout  = 8'b11111111; // 4012 : 255 - 0xff
      12'hFAD: dout  = 8'b11111111; // 4013 : 255 - 0xff
      12'hFAE: dout  = 8'b11111111; // 4014 : 255 - 0xff
      12'hFAF: dout  = 8'b11111111; // 4015 : 255 - 0xff
      12'hFB0: dout  = 8'b11111111; // 4016 : 255 - 0xff -- Background 0xf6
      12'hFB1: dout  = 8'b11111111; // 4017 : 255 - 0xff
      12'hFB2: dout  = 8'b11111111; // 4018 : 255 - 0xff
      12'hFB3: dout  = 8'b11111111; // 4019 : 255 - 0xff
      12'hFB4: dout  = 8'b11111111; // 4020 : 255 - 0xff
      12'hFB5: dout  = 8'b11111111; // 4021 : 255 - 0xff
      12'hFB6: dout  = 8'b11111111; // 4022 : 255 - 0xff
      12'hFB7: dout  = 8'b11111111; // 4023 : 255 - 0xff
      12'hFB8: dout  = 8'b11111111; // 4024 : 255 - 0xff -- Background 0xf7
      12'hFB9: dout  = 8'b11111111; // 4025 : 255 - 0xff
      12'hFBA: dout  = 8'b11111111; // 4026 : 255 - 0xff
      12'hFBB: dout  = 8'b11111111; // 4027 : 255 - 0xff
      12'hFBC: dout  = 8'b11111111; // 4028 : 255 - 0xff
      12'hFBD: dout  = 8'b11111111; // 4029 : 255 - 0xff
      12'hFBE: dout  = 8'b11111111; // 4030 : 255 - 0xff
      12'hFBF: dout  = 8'b11111111; // 4031 : 255 - 0xff
      12'hFC0: dout  = 8'b11111111; // 4032 : 255 - 0xff -- Background 0xf8
      12'hFC1: dout  = 8'b11111111; // 4033 : 255 - 0xff
      12'hFC2: dout  = 8'b11111111; // 4034 : 255 - 0xff
      12'hFC3: dout  = 8'b11111111; // 4035 : 255 - 0xff
      12'hFC4: dout  = 8'b11111111; // 4036 : 255 - 0xff
      12'hFC5: dout  = 8'b11111111; // 4037 : 255 - 0xff
      12'hFC6: dout  = 8'b11111111; // 4038 : 255 - 0xff
      12'hFC7: dout  = 8'b11111111; // 4039 : 255 - 0xff
      12'hFC8: dout  = 8'b11111111; // 4040 : 255 - 0xff -- Background 0xf9
      12'hFC9: dout  = 8'b11111111; // 4041 : 255 - 0xff
      12'hFCA: dout  = 8'b11111111; // 4042 : 255 - 0xff
      12'hFCB: dout  = 8'b11111111; // 4043 : 255 - 0xff
      12'hFCC: dout  = 8'b11111111; // 4044 : 255 - 0xff
      12'hFCD: dout  = 8'b11111111; // 4045 : 255 - 0xff
      12'hFCE: dout  = 8'b11111111; // 4046 : 255 - 0xff
      12'hFCF: dout  = 8'b11111111; // 4047 : 255 - 0xff
      12'hFD0: dout  = 8'b11111111; // 4048 : 255 - 0xff -- Background 0xfa
      12'hFD1: dout  = 8'b11111111; // 4049 : 255 - 0xff
      12'hFD2: dout  = 8'b11111111; // 4050 : 255 - 0xff
      12'hFD3: dout  = 8'b11111111; // 4051 : 255 - 0xff
      12'hFD4: dout  = 8'b11111111; // 4052 : 255 - 0xff
      12'hFD5: dout  = 8'b11111111; // 4053 : 255 - 0xff
      12'hFD6: dout  = 8'b11111111; // 4054 : 255 - 0xff
      12'hFD7: dout  = 8'b11111111; // 4055 : 255 - 0xff
      12'hFD8: dout  = 8'b11111111; // 4056 : 255 - 0xff -- Background 0xfb
      12'hFD9: dout  = 8'b11111111; // 4057 : 255 - 0xff
      12'hFDA: dout  = 8'b11111111; // 4058 : 255 - 0xff
      12'hFDB: dout  = 8'b11111111; // 4059 : 255 - 0xff
      12'hFDC: dout  = 8'b11111111; // 4060 : 255 - 0xff
      12'hFDD: dout  = 8'b11111111; // 4061 : 255 - 0xff
      12'hFDE: dout  = 8'b11111111; // 4062 : 255 - 0xff
      12'hFDF: dout  = 8'b11111111; // 4063 : 255 - 0xff
      12'hFE0: dout  = 8'b11111111; // 4064 : 255 - 0xff -- Background 0xfc
      12'hFE1: dout  = 8'b11111111; // 4065 : 255 - 0xff
      12'hFE2: dout  = 8'b11111111; // 4066 : 255 - 0xff
      12'hFE3: dout  = 8'b11111111; // 4067 : 255 - 0xff
      12'hFE4: dout  = 8'b11111111; // 4068 : 255 - 0xff
      12'hFE5: dout  = 8'b11111111; // 4069 : 255 - 0xff
      12'hFE6: dout  = 8'b11111111; // 4070 : 255 - 0xff
      12'hFE7: dout  = 8'b11111111; // 4071 : 255 - 0xff
      12'hFE8: dout  = 8'b11111111; // 4072 : 255 - 0xff -- Background 0xfd
      12'hFE9: dout  = 8'b11111111; // 4073 : 255 - 0xff
      12'hFEA: dout  = 8'b11111111; // 4074 : 255 - 0xff
      12'hFEB: dout  = 8'b11111111; // 4075 : 255 - 0xff
      12'hFEC: dout  = 8'b11111111; // 4076 : 255 - 0xff
      12'hFED: dout  = 8'b11111111; // 4077 : 255 - 0xff
      12'hFEE: dout  = 8'b11111111; // 4078 : 255 - 0xff
      12'hFEF: dout  = 8'b11111111; // 4079 : 255 - 0xff
      12'hFF0: dout  = 8'b11111111; // 4080 : 255 - 0xff -- Background 0xfe
      12'hFF1: dout  = 8'b11111111; // 4081 : 255 - 0xff
      12'hFF2: dout  = 8'b11111111; // 4082 : 255 - 0xff
      12'hFF3: dout  = 8'b11111111; // 4083 : 255 - 0xff
      12'hFF4: dout  = 8'b11111111; // 4084 : 255 - 0xff
      12'hFF5: dout  = 8'b11111111; // 4085 : 255 - 0xff
      12'hFF6: dout  = 8'b11111111; // 4086 : 255 - 0xff
      12'hFF7: dout  = 8'b11111111; // 4087 : 255 - 0xff
      12'hFF8: dout  = 8'b11111111; // 4088 : 255 - 0xff -- Background 0xff
      12'hFF9: dout  = 8'b11111111; // 4089 : 255 - 0xff
      12'hFFA: dout  = 8'b11111111; // 4090 : 255 - 0xff
      12'hFFB: dout  = 8'b11111111; // 4091 : 255 - 0xff
      12'hFFC: dout  = 8'b11111111; // 4092 : 255 - 0xff
      12'hFFD: dout  = 8'b11111111; // 4093 : 255 - 0xff
      12'hFFE: dout  = 8'b11111111; // 4094 : 255 - 0xff
      12'hFFF: dout  = 8'b11111111; // 4095 : 255 - 0xff
    endcase
  end

endmodule
