//-   Background Pattern table BOTH COLOR PLANES
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
//- Autcmatically generated verilog ROM from a NES memory file----


//-  Original memory dump file name: pacman_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_PTABLE_PACMAN_BG
  (
     input     clk,   // clock
     input      [12-1:0] addr,  //4096 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Background pattern Table both color planes
      12'h0: dout <= 8'b00000000; //    0 :   0 - 0x0 -- Background 0x0
      12'h1: dout <= 8'b00000000; //    1 :   0 - 0x0
      12'h2: dout <= 8'b00000000; //    2 :   0 - 0x0
      12'h3: dout <= 8'b00000000; //    3 :   0 - 0x0
      12'h4: dout <= 8'b00000000; //    4 :   0 - 0x0
      12'h5: dout <= 8'b00000000; //    5 :   0 - 0x0
      12'h6: dout <= 8'b00000000; //    6 :   0 - 0x0
      12'h7: dout <= 8'b00000000; //    7 :   0 - 0x0
      12'h8: dout <= 8'b00000000; //    8 :   0 - 0x0 -- plane 1
      12'h9: dout <= 8'b00000000; //    9 :   0 - 0x0
      12'hA: dout <= 8'b00000000; //   10 :   0 - 0x0
      12'hB: dout <= 8'b00000000; //   11 :   0 - 0x0
      12'hC: dout <= 8'b00000000; //   12 :   0 - 0x0
      12'hD: dout <= 8'b00000000; //   13 :   0 - 0x0
      12'hE: dout <= 8'b00000000; //   14 :   0 - 0x0
      12'hF: dout <= 8'b00000000; //   15 :   0 - 0x0
      12'h10: dout <= 8'b00000000; //   16 :   0 - 0x0 -- Background 0x1
      12'h11: dout <= 8'b00111000; //   17 :  56 - 0x38
      12'h12: dout <= 8'b01111100; //   18 : 124 - 0x7c
      12'h13: dout <= 8'b11111110; //   19 : 254 - 0xfe
      12'h14: dout <= 8'b11111110; //   20 : 254 - 0xfe
      12'h15: dout <= 8'b11111110; //   21 : 254 - 0xfe
      12'h16: dout <= 8'b01111100; //   22 : 124 - 0x7c
      12'h17: dout <= 8'b00111000; //   23 :  56 - 0x38
      12'h18: dout <= 8'b00000000; //   24 :   0 - 0x0 -- plane 1
      12'h19: dout <= 8'b00111000; //   25 :  56 - 0x38
      12'h1A: dout <= 8'b01111100; //   26 : 124 - 0x7c
      12'h1B: dout <= 8'b11111110; //   27 : 254 - 0xfe
      12'h1C: dout <= 8'b11111110; //   28 : 254 - 0xfe
      12'h1D: dout <= 8'b11111110; //   29 : 254 - 0xfe
      12'h1E: dout <= 8'b01111100; //   30 : 124 - 0x7c
      12'h1F: dout <= 8'b00111000; //   31 :  56 - 0x38
      12'h20: dout <= 8'b00000000; //   32 :   0 - 0x0 -- Background 0x2
      12'h21: dout <= 8'b00000000; //   33 :   0 - 0x0
      12'h22: dout <= 8'b00000000; //   34 :   0 - 0x0
      12'h23: dout <= 8'b00000000; //   35 :   0 - 0x0
      12'h24: dout <= 8'b00000000; //   36 :   0 - 0x0
      12'h25: dout <= 8'b00000000; //   37 :   0 - 0x0
      12'h26: dout <= 8'b00000000; //   38 :   0 - 0x0
      12'h27: dout <= 8'b00000000; //   39 :   0 - 0x0
      12'h28: dout <= 8'b00000000; //   40 :   0 - 0x0 -- plane 1
      12'h29: dout <= 8'b00000000; //   41 :   0 - 0x0
      12'h2A: dout <= 8'b00000000; //   42 :   0 - 0x0
      12'h2B: dout <= 8'b00000000; //   43 :   0 - 0x0
      12'h2C: dout <= 8'b00000000; //   44 :   0 - 0x0
      12'h2D: dout <= 8'b00000000; //   45 :   0 - 0x0
      12'h2E: dout <= 8'b00000000; //   46 :   0 - 0x0
      12'h2F: dout <= 8'b00000000; //   47 :   0 - 0x0
      12'h30: dout <= 8'b00000000; //   48 :   0 - 0x0 -- Background 0x3
      12'h31: dout <= 8'b00000000; //   49 :   0 - 0x0
      12'h32: dout <= 8'b00000000; //   50 :   0 - 0x0
      12'h33: dout <= 8'b00011000; //   51 :  24 - 0x18
      12'h34: dout <= 8'b00011000; //   52 :  24 - 0x18
      12'h35: dout <= 8'b00000000; //   53 :   0 - 0x0
      12'h36: dout <= 8'b00000000; //   54 :   0 - 0x0
      12'h37: dout <= 8'b00000000; //   55 :   0 - 0x0
      12'h38: dout <= 8'b00000000; //   56 :   0 - 0x0 -- plane 1
      12'h39: dout <= 8'b00000000; //   57 :   0 - 0x0
      12'h3A: dout <= 8'b00000000; //   58 :   0 - 0x0
      12'h3B: dout <= 8'b00011000; //   59 :  24 - 0x18
      12'h3C: dout <= 8'b00011000; //   60 :  24 - 0x18
      12'h3D: dout <= 8'b00000000; //   61 :   0 - 0x0
      12'h3E: dout <= 8'b00000000; //   62 :   0 - 0x0
      12'h3F: dout <= 8'b00000000; //   63 :   0 - 0x0
      12'h40: dout <= 8'b00000000; //   64 :   0 - 0x0 -- Background 0x4
      12'h41: dout <= 8'b00000000; //   65 :   0 - 0x0
      12'h42: dout <= 8'b00000000; //   66 :   0 - 0x0
      12'h43: dout <= 8'b00000000; //   67 :   0 - 0x0
      12'h44: dout <= 8'b00000000; //   68 :   0 - 0x0
      12'h45: dout <= 8'b00000000; //   69 :   0 - 0x0
      12'h46: dout <= 8'b00000000; //   70 :   0 - 0x0
      12'h47: dout <= 8'b00000000; //   71 :   0 - 0x0
      12'h48: dout <= 8'b11111111; //   72 : 255 - 0xff -- plane 1
      12'h49: dout <= 8'b11111111; //   73 : 255 - 0xff
      12'h4A: dout <= 8'b11111111; //   74 : 255 - 0xff
      12'h4B: dout <= 8'b11111111; //   75 : 255 - 0xff
      12'h4C: dout <= 8'b11111111; //   76 : 255 - 0xff
      12'h4D: dout <= 8'b11111111; //   77 : 255 - 0xff
      12'h4E: dout <= 8'b11111111; //   78 : 255 - 0xff
      12'h4F: dout <= 8'b11111111; //   79 : 255 - 0xff
      12'h50: dout <= 8'b00000000; //   80 :   0 - 0x0 -- Background 0x5
      12'h51: dout <= 8'b00000000; //   81 :   0 - 0x0
      12'h52: dout <= 8'b00000000; //   82 :   0 - 0x0
      12'h53: dout <= 8'b00000000; //   83 :   0 - 0x0
      12'h54: dout <= 8'b00000000; //   84 :   0 - 0x0
      12'h55: dout <= 8'b00000000; //   85 :   0 - 0x0
      12'h56: dout <= 8'b00000000; //   86 :   0 - 0x0
      12'h57: dout <= 8'b00000000; //   87 :   0 - 0x0
      12'h58: dout <= 8'b00001111; //   88 :  15 - 0xf -- plane 1
      12'h59: dout <= 8'b00001111; //   89 :  15 - 0xf
      12'h5A: dout <= 8'b00001111; //   90 :  15 - 0xf
      12'h5B: dout <= 8'b00001111; //   91 :  15 - 0xf
      12'h5C: dout <= 8'b00001111; //   92 :  15 - 0xf
      12'h5D: dout <= 8'b00001111; //   93 :  15 - 0xf
      12'h5E: dout <= 8'b00001111; //   94 :  15 - 0xf
      12'h5F: dout <= 8'b00001111; //   95 :  15 - 0xf
      12'h60: dout <= 8'b00000000; //   96 :   0 - 0x0 -- Background 0x6
      12'h61: dout <= 8'b00000000; //   97 :   0 - 0x0
      12'h62: dout <= 8'b00000000; //   98 :   0 - 0x0
      12'h63: dout <= 8'b00000000; //   99 :   0 - 0x0
      12'h64: dout <= 8'b00000000; //  100 :   0 - 0x0
      12'h65: dout <= 8'b00000000; //  101 :   0 - 0x0
      12'h66: dout <= 8'b00000000; //  102 :   0 - 0x0
      12'h67: dout <= 8'b00000000; //  103 :   0 - 0x0
      12'h68: dout <= 8'b11110000; //  104 : 240 - 0xf0 -- plane 1
      12'h69: dout <= 8'b11110000; //  105 : 240 - 0xf0
      12'h6A: dout <= 8'b11110000; //  106 : 240 - 0xf0
      12'h6B: dout <= 8'b11110000; //  107 : 240 - 0xf0
      12'h6C: dout <= 8'b11110000; //  108 : 240 - 0xf0
      12'h6D: dout <= 8'b11110000; //  109 : 240 - 0xf0
      12'h6E: dout <= 8'b11110000; //  110 : 240 - 0xf0
      12'h6F: dout <= 8'b11110000; //  111 : 240 - 0xf0
      12'h70: dout <= 8'b00000000; //  112 :   0 - 0x0 -- Background 0x7
      12'h71: dout <= 8'b00000000; //  113 :   0 - 0x0
      12'h72: dout <= 8'b00000000; //  114 :   0 - 0x0
      12'h73: dout <= 8'b00000000; //  115 :   0 - 0x0
      12'h74: dout <= 8'b00000000; //  116 :   0 - 0x0
      12'h75: dout <= 8'b00000000; //  117 :   0 - 0x0
      12'h76: dout <= 8'b00000000; //  118 :   0 - 0x0
      12'h77: dout <= 8'b00000000; //  119 :   0 - 0x0
      12'h78: dout <= 8'b00000000; //  120 :   0 - 0x0 -- plane 1
      12'h79: dout <= 8'b00000000; //  121 :   0 - 0x0
      12'h7A: dout <= 8'b00000000; //  122 :   0 - 0x0
      12'h7B: dout <= 8'b00000000; //  123 :   0 - 0x0
      12'h7C: dout <= 8'b00000000; //  124 :   0 - 0x0
      12'h7D: dout <= 8'b00000000; //  125 :   0 - 0x0
      12'h7E: dout <= 8'b00000000; //  126 :   0 - 0x0
      12'h7F: dout <= 8'b00000000; //  127 :   0 - 0x0
      12'h80: dout <= 8'b00000000; //  128 :   0 - 0x0 -- Background 0x8
      12'h81: dout <= 8'b00000000; //  129 :   0 - 0x0
      12'h82: dout <= 8'b00000000; //  130 :   0 - 0x0
      12'h83: dout <= 8'b00000000; //  131 :   0 - 0x0
      12'h84: dout <= 8'b00000000; //  132 :   0 - 0x0
      12'h85: dout <= 8'b00000000; //  133 :   0 - 0x0
      12'h86: dout <= 8'b00000000; //  134 :   0 - 0x0
      12'h87: dout <= 8'b00000000; //  135 :   0 - 0x0
      12'h88: dout <= 8'b00000000; //  136 :   0 - 0x0 -- plane 1
      12'h89: dout <= 8'b00000000; //  137 :   0 - 0x0
      12'h8A: dout <= 8'b00000000; //  138 :   0 - 0x0
      12'h8B: dout <= 8'b00000000; //  139 :   0 - 0x0
      12'h8C: dout <= 8'b00000000; //  140 :   0 - 0x0
      12'h8D: dout <= 8'b00000000; //  141 :   0 - 0x0
      12'h8E: dout <= 8'b00000000; //  142 :   0 - 0x0
      12'h8F: dout <= 8'b00000000; //  143 :   0 - 0x0
      12'h90: dout <= 8'b00000000; //  144 :   0 - 0x0 -- Background 0x9
      12'h91: dout <= 8'b00000000; //  145 :   0 - 0x0
      12'h92: dout <= 8'b00000000; //  146 :   0 - 0x0
      12'h93: dout <= 8'b00011000; //  147 :  24 - 0x18
      12'h94: dout <= 8'b00011000; //  148 :  24 - 0x18
      12'h95: dout <= 8'b00000000; //  149 :   0 - 0x0
      12'h96: dout <= 8'b00000000; //  150 :   0 - 0x0
      12'h97: dout <= 8'b00000000; //  151 :   0 - 0x0
      12'h98: dout <= 8'b00000000; //  152 :   0 - 0x0 -- plane 1
      12'h99: dout <= 8'b00000000; //  153 :   0 - 0x0
      12'h9A: dout <= 8'b00000000; //  154 :   0 - 0x0
      12'h9B: dout <= 8'b00011000; //  155 :  24 - 0x18
      12'h9C: dout <= 8'b00011000; //  156 :  24 - 0x18
      12'h9D: dout <= 8'b00000000; //  157 :   0 - 0x0
      12'h9E: dout <= 8'b00000000; //  158 :   0 - 0x0
      12'h9F: dout <= 8'b00000000; //  159 :   0 - 0x0
      12'hA0: dout <= 8'b00000000; //  160 :   0 - 0x0 -- Background 0xa
      12'hA1: dout <= 8'b00000000; //  161 :   0 - 0x0
      12'hA2: dout <= 8'b00000000; //  162 :   0 - 0x0
      12'hA3: dout <= 8'b00000000; //  163 :   0 - 0x0
      12'hA4: dout <= 8'b00000000; //  164 :   0 - 0x0
      12'hA5: dout <= 8'b00000000; //  165 :   0 - 0x0
      12'hA6: dout <= 8'b00000000; //  166 :   0 - 0x0
      12'hA7: dout <= 8'b00000000; //  167 :   0 - 0x0
      12'hA8: dout <= 8'b00000000; //  168 :   0 - 0x0 -- plane 1
      12'hA9: dout <= 8'b00000000; //  169 :   0 - 0x0
      12'hAA: dout <= 8'b00000000; //  170 :   0 - 0x0
      12'hAB: dout <= 8'b00000000; //  171 :   0 - 0x0
      12'hAC: dout <= 8'b00000000; //  172 :   0 - 0x0
      12'hAD: dout <= 8'b00000000; //  173 :   0 - 0x0
      12'hAE: dout <= 8'b00000000; //  174 :   0 - 0x0
      12'hAF: dout <= 8'b00000000; //  175 :   0 - 0x0
      12'hB0: dout <= 8'b00000000; //  176 :   0 - 0x0 -- Background 0xb
      12'hB1: dout <= 8'b00000000; //  177 :   0 - 0x0
      12'hB2: dout <= 8'b00000000; //  178 :   0 - 0x0
      12'hB3: dout <= 8'b00000000; //  179 :   0 - 0x0
      12'hB4: dout <= 8'b00000000; //  180 :   0 - 0x0
      12'hB5: dout <= 8'b00000000; //  181 :   0 - 0x0
      12'hB6: dout <= 8'b00000000; //  182 :   0 - 0x0
      12'hB7: dout <= 8'b00000000; //  183 :   0 - 0x0
      12'hB8: dout <= 8'b00000000; //  184 :   0 - 0x0 -- plane 1
      12'hB9: dout <= 8'b00000000; //  185 :   0 - 0x0
      12'hBA: dout <= 8'b00000000; //  186 :   0 - 0x0
      12'hBB: dout <= 8'b00000000; //  187 :   0 - 0x0
      12'hBC: dout <= 8'b00000000; //  188 :   0 - 0x0
      12'hBD: dout <= 8'b00000000; //  189 :   0 - 0x0
      12'hBE: dout <= 8'b00000000; //  190 :   0 - 0x0
      12'hBF: dout <= 8'b00000000; //  191 :   0 - 0x0
      12'hC0: dout <= 8'b00000000; //  192 :   0 - 0x0 -- Background 0xc
      12'hC1: dout <= 8'b00000000; //  193 :   0 - 0x0
      12'hC2: dout <= 8'b00000000; //  194 :   0 - 0x0
      12'hC3: dout <= 8'b00000000; //  195 :   0 - 0x0
      12'hC4: dout <= 8'b00000000; //  196 :   0 - 0x0
      12'hC5: dout <= 8'b00000000; //  197 :   0 - 0x0
      12'hC6: dout <= 8'b00000000; //  198 :   0 - 0x0
      12'hC7: dout <= 8'b00000000; //  199 :   0 - 0x0
      12'hC8: dout <= 8'b00000000; //  200 :   0 - 0x0 -- plane 1
      12'hC9: dout <= 8'b00000000; //  201 :   0 - 0x0
      12'hCA: dout <= 8'b00000000; //  202 :   0 - 0x0
      12'hCB: dout <= 8'b00000000; //  203 :   0 - 0x0
      12'hCC: dout <= 8'b00000000; //  204 :   0 - 0x0
      12'hCD: dout <= 8'b00000000; //  205 :   0 - 0x0
      12'hCE: dout <= 8'b00000000; //  206 :   0 - 0x0
      12'hCF: dout <= 8'b00000000; //  207 :   0 - 0x0
      12'hD0: dout <= 8'b00000000; //  208 :   0 - 0x0 -- Background 0xd
      12'hD1: dout <= 8'b00000000; //  209 :   0 - 0x0
      12'hD2: dout <= 8'b00000000; //  210 :   0 - 0x0
      12'hD3: dout <= 8'b00000000; //  211 :   0 - 0x0
      12'hD4: dout <= 8'b00000000; //  212 :   0 - 0x0
      12'hD5: dout <= 8'b00000000; //  213 :   0 - 0x0
      12'hD6: dout <= 8'b00000000; //  214 :   0 - 0x0
      12'hD7: dout <= 8'b00000000; //  215 :   0 - 0x0
      12'hD8: dout <= 8'b00000000; //  216 :   0 - 0x0 -- plane 1
      12'hD9: dout <= 8'b00000000; //  217 :   0 - 0x0
      12'hDA: dout <= 8'b00000000; //  218 :   0 - 0x0
      12'hDB: dout <= 8'b00000000; //  219 :   0 - 0x0
      12'hDC: dout <= 8'b00000000; //  220 :   0 - 0x0
      12'hDD: dout <= 8'b00000000; //  221 :   0 - 0x0
      12'hDE: dout <= 8'b00000000; //  222 :   0 - 0x0
      12'hDF: dout <= 8'b00000000; //  223 :   0 - 0x0
      12'hE0: dout <= 8'b00000000; //  224 :   0 - 0x0 -- Background 0xe
      12'hE1: dout <= 8'b00000000; //  225 :   0 - 0x0
      12'hE2: dout <= 8'b00000000; //  226 :   0 - 0x0
      12'hE3: dout <= 8'b00000000; //  227 :   0 - 0x0
      12'hE4: dout <= 8'b00000000; //  228 :   0 - 0x0
      12'hE5: dout <= 8'b00000000; //  229 :   0 - 0x0
      12'hE6: dout <= 8'b00000000; //  230 :   0 - 0x0
      12'hE7: dout <= 8'b00000000; //  231 :   0 - 0x0
      12'hE8: dout <= 8'b00000000; //  232 :   0 - 0x0 -- plane 1
      12'hE9: dout <= 8'b00000000; //  233 :   0 - 0x0
      12'hEA: dout <= 8'b00000000; //  234 :   0 - 0x0
      12'hEB: dout <= 8'b00000000; //  235 :   0 - 0x0
      12'hEC: dout <= 8'b00000000; //  236 :   0 - 0x0
      12'hED: dout <= 8'b00000000; //  237 :   0 - 0x0
      12'hEE: dout <= 8'b00000000; //  238 :   0 - 0x0
      12'hEF: dout <= 8'b00000000; //  239 :   0 - 0x0
      12'hF0: dout <= 8'b00000000; //  240 :   0 - 0x0 -- Background 0xf
      12'hF1: dout <= 8'b00000000; //  241 :   0 - 0x0
      12'hF2: dout <= 8'b00000000; //  242 :   0 - 0x0
      12'hF3: dout <= 8'b00000000; //  243 :   0 - 0x0
      12'hF4: dout <= 8'b00000000; //  244 :   0 - 0x0
      12'hF5: dout <= 8'b00000000; //  245 :   0 - 0x0
      12'hF6: dout <= 8'b00000000; //  246 :   0 - 0x0
      12'hF7: dout <= 8'b00000000; //  247 :   0 - 0x0
      12'hF8: dout <= 8'b00000000; //  248 :   0 - 0x0 -- plane 1
      12'hF9: dout <= 8'b00000000; //  249 :   0 - 0x0
      12'hFA: dout <= 8'b00000000; //  250 :   0 - 0x0
      12'hFB: dout <= 8'b00000000; //  251 :   0 - 0x0
      12'hFC: dout <= 8'b00000000; //  252 :   0 - 0x0
      12'hFD: dout <= 8'b00000000; //  253 :   0 - 0x0
      12'hFE: dout <= 8'b00000000; //  254 :   0 - 0x0
      12'hFF: dout <= 8'b00000000; //  255 :   0 - 0x0
      12'h100: dout <= 8'b00000000; //  256 :   0 - 0x0 -- Background 0x10
      12'h101: dout <= 8'b00000000; //  257 :   0 - 0x0
      12'h102: dout <= 8'b11111111; //  258 : 255 - 0xff
      12'h103: dout <= 8'b00000000; //  259 :   0 - 0x0
      12'h104: dout <= 8'b00000000; //  260 :   0 - 0x0
      12'h105: dout <= 8'b11111111; //  261 : 255 - 0xff
      12'h106: dout <= 8'b00000000; //  262 :   0 - 0x0
      12'h107: dout <= 8'b00000000; //  263 :   0 - 0x0
      12'h108: dout <= 8'b00000000; //  264 :   0 - 0x0 -- plane 1
      12'h109: dout <= 8'b00000000; //  265 :   0 - 0x0
      12'h10A: dout <= 8'b00000000; //  266 :   0 - 0x0
      12'h10B: dout <= 8'b00000000; //  267 :   0 - 0x0
      12'h10C: dout <= 8'b00000000; //  268 :   0 - 0x0
      12'h10D: dout <= 8'b00000000; //  269 :   0 - 0x0
      12'h10E: dout <= 8'b00000000; //  270 :   0 - 0x0
      12'h10F: dout <= 8'b00000000; //  271 :   0 - 0x0
      12'h110: dout <= 8'b00100100; //  272 :  36 - 0x24 -- Background 0x11
      12'h111: dout <= 8'b00100100; //  273 :  36 - 0x24
      12'h112: dout <= 8'b00100100; //  274 :  36 - 0x24
      12'h113: dout <= 8'b00100100; //  275 :  36 - 0x24
      12'h114: dout <= 8'b00100100; //  276 :  36 - 0x24
      12'h115: dout <= 8'b00100100; //  277 :  36 - 0x24
      12'h116: dout <= 8'b00100100; //  278 :  36 - 0x24
      12'h117: dout <= 8'b00100100; //  279 :  36 - 0x24
      12'h118: dout <= 8'b00000000; //  280 :   0 - 0x0 -- plane 1
      12'h119: dout <= 8'b00000000; //  281 :   0 - 0x0
      12'h11A: dout <= 8'b00000000; //  282 :   0 - 0x0
      12'h11B: dout <= 8'b00000000; //  283 :   0 - 0x0
      12'h11C: dout <= 8'b00000000; //  284 :   0 - 0x0
      12'h11D: dout <= 8'b00000000; //  285 :   0 - 0x0
      12'h11E: dout <= 8'b00000000; //  286 :   0 - 0x0
      12'h11F: dout <= 8'b00000000; //  287 :   0 - 0x0
      12'h120: dout <= 8'b00100100; //  288 :  36 - 0x24 -- Background 0x12
      12'h121: dout <= 8'b00100100; //  289 :  36 - 0x24
      12'h122: dout <= 8'b11000011; //  290 : 195 - 0xc3
      12'h123: dout <= 8'b00000000; //  291 :   0 - 0x0
      12'h124: dout <= 8'b00000000; //  292 :   0 - 0x0
      12'h125: dout <= 8'b11111111; //  293 : 255 - 0xff
      12'h126: dout <= 8'b00000000; //  294 :   0 - 0x0
      12'h127: dout <= 8'b00000000; //  295 :   0 - 0x0
      12'h128: dout <= 8'b00000000; //  296 :   0 - 0x0 -- plane 1
      12'h129: dout <= 8'b00000000; //  297 :   0 - 0x0
      12'h12A: dout <= 8'b00000000; //  298 :   0 - 0x0
      12'h12B: dout <= 8'b00000000; //  299 :   0 - 0x0
      12'h12C: dout <= 8'b00000000; //  300 :   0 - 0x0
      12'h12D: dout <= 8'b00000000; //  301 :   0 - 0x0
      12'h12E: dout <= 8'b00000000; //  302 :   0 - 0x0
      12'h12F: dout <= 8'b00000000; //  303 :   0 - 0x0
      12'h130: dout <= 8'b00000000; //  304 :   0 - 0x0 -- Background 0x13
      12'h131: dout <= 8'b00000000; //  305 :   0 - 0x0
      12'h132: dout <= 8'b11111111; //  306 : 255 - 0xff
      12'h133: dout <= 8'b00000000; //  307 :   0 - 0x0
      12'h134: dout <= 8'b00000000; //  308 :   0 - 0x0
      12'h135: dout <= 8'b11000011; //  309 : 195 - 0xc3
      12'h136: dout <= 8'b00100100; //  310 :  36 - 0x24
      12'h137: dout <= 8'b00100100; //  311 :  36 - 0x24
      12'h138: dout <= 8'b00000000; //  312 :   0 - 0x0 -- plane 1
      12'h139: dout <= 8'b00000000; //  313 :   0 - 0x0
      12'h13A: dout <= 8'b00000000; //  314 :   0 - 0x0
      12'h13B: dout <= 8'b00000000; //  315 :   0 - 0x0
      12'h13C: dout <= 8'b00000000; //  316 :   0 - 0x0
      12'h13D: dout <= 8'b00000000; //  317 :   0 - 0x0
      12'h13E: dout <= 8'b00000000; //  318 :   0 - 0x0
      12'h13F: dout <= 8'b00000000; //  319 :   0 - 0x0
      12'h140: dout <= 8'b00100100; //  320 :  36 - 0x24 -- Background 0x14
      12'h141: dout <= 8'b00100100; //  321 :  36 - 0x24
      12'h142: dout <= 8'b11000100; //  322 : 196 - 0xc4
      12'h143: dout <= 8'b00000100; //  323 :   4 - 0x4
      12'h144: dout <= 8'b00000100; //  324 :   4 - 0x4
      12'h145: dout <= 8'b11000100; //  325 : 196 - 0xc4
      12'h146: dout <= 8'b00100100; //  326 :  36 - 0x24
      12'h147: dout <= 8'b00100100; //  327 :  36 - 0x24
      12'h148: dout <= 8'b00000000; //  328 :   0 - 0x0 -- plane 1
      12'h149: dout <= 8'b00000000; //  329 :   0 - 0x0
      12'h14A: dout <= 8'b00000000; //  330 :   0 - 0x0
      12'h14B: dout <= 8'b00000000; //  331 :   0 - 0x0
      12'h14C: dout <= 8'b00000000; //  332 :   0 - 0x0
      12'h14D: dout <= 8'b00000000; //  333 :   0 - 0x0
      12'h14E: dout <= 8'b00000000; //  334 :   0 - 0x0
      12'h14F: dout <= 8'b00000000; //  335 :   0 - 0x0
      12'h150: dout <= 8'b00100100; //  336 :  36 - 0x24 -- Background 0x15
      12'h151: dout <= 8'b00100100; //  337 :  36 - 0x24
      12'h152: dout <= 8'b00100011; //  338 :  35 - 0x23
      12'h153: dout <= 8'b00100000; //  339 :  32 - 0x20
      12'h154: dout <= 8'b00100000; //  340 :  32 - 0x20
      12'h155: dout <= 8'b00100011; //  341 :  35 - 0x23
      12'h156: dout <= 8'b00100100; //  342 :  36 - 0x24
      12'h157: dout <= 8'b00100100; //  343 :  36 - 0x24
      12'h158: dout <= 8'b00000000; //  344 :   0 - 0x0 -- plane 1
      12'h159: dout <= 8'b00000000; //  345 :   0 - 0x0
      12'h15A: dout <= 8'b00000000; //  346 :   0 - 0x0
      12'h15B: dout <= 8'b00000000; //  347 :   0 - 0x0
      12'h15C: dout <= 8'b00000000; //  348 :   0 - 0x0
      12'h15D: dout <= 8'b00000000; //  349 :   0 - 0x0
      12'h15E: dout <= 8'b00000000; //  350 :   0 - 0x0
      12'h15F: dout <= 8'b00000000; //  351 :   0 - 0x0
      12'h160: dout <= 8'b00000000; //  352 :   0 - 0x0 -- Background 0x16
      12'h161: dout <= 8'b00000000; //  353 :   0 - 0x0
      12'h162: dout <= 8'b00001111; //  354 :  15 - 0xf
      12'h163: dout <= 8'b00010000; //  355 :  16 - 0x10
      12'h164: dout <= 8'b11110000; //  356 : 240 - 0xf0
      12'h165: dout <= 8'b00001111; //  357 :  15 - 0xf
      12'h166: dout <= 8'b00000000; //  358 :   0 - 0x0
      12'h167: dout <= 8'b00000000; //  359 :   0 - 0x0
      12'h168: dout <= 8'b00000000; //  360 :   0 - 0x0 -- plane 1
      12'h169: dout <= 8'b00000000; //  361 :   0 - 0x0
      12'h16A: dout <= 8'b00000000; //  362 :   0 - 0x0
      12'h16B: dout <= 8'b00000000; //  363 :   0 - 0x0
      12'h16C: dout <= 8'b00000000; //  364 :   0 - 0x0
      12'h16D: dout <= 8'b00000000; //  365 :   0 - 0x0
      12'h16E: dout <= 8'b00000000; //  366 :   0 - 0x0
      12'h16F: dout <= 8'b00000000; //  367 :   0 - 0x0
      12'h170: dout <= 8'b00000000; //  368 :   0 - 0x0 -- Background 0x17
      12'h171: dout <= 8'b00000000; //  369 :   0 - 0x0
      12'h172: dout <= 8'b11110000; //  370 : 240 - 0xf0
      12'h173: dout <= 8'b00001000; //  371 :   8 - 0x8
      12'h174: dout <= 8'b00001111; //  372 :  15 - 0xf
      12'h175: dout <= 8'b11110000; //  373 : 240 - 0xf0
      12'h176: dout <= 8'b00000000; //  374 :   0 - 0x0
      12'h177: dout <= 8'b00000000; //  375 :   0 - 0x0
      12'h178: dout <= 8'b00000000; //  376 :   0 - 0x0 -- plane 1
      12'h179: dout <= 8'b00000000; //  377 :   0 - 0x0
      12'h17A: dout <= 8'b00000000; //  378 :   0 - 0x0
      12'h17B: dout <= 8'b00000000; //  379 :   0 - 0x0
      12'h17C: dout <= 8'b00000000; //  380 :   0 - 0x0
      12'h17D: dout <= 8'b00000000; //  381 :   0 - 0x0
      12'h17E: dout <= 8'b00000000; //  382 :   0 - 0x0
      12'h17F: dout <= 8'b00000000; //  383 :   0 - 0x0
      12'h180: dout <= 8'b00000000; //  384 :   0 - 0x0 -- Background 0x18
      12'h181: dout <= 8'b00000000; //  385 :   0 - 0x0
      12'h182: dout <= 8'b11110000; //  386 : 240 - 0xf0
      12'h183: dout <= 8'b00001000; //  387 :   8 - 0x8
      12'h184: dout <= 8'b00001000; //  388 :   8 - 0x8
      12'h185: dout <= 8'b11110000; //  389 : 240 - 0xf0
      12'h186: dout <= 8'b00000000; //  390 :   0 - 0x0
      12'h187: dout <= 8'b00000000; //  391 :   0 - 0x0
      12'h188: dout <= 8'b00000000; //  392 :   0 - 0x0 -- plane 1
      12'h189: dout <= 8'b00000000; //  393 :   0 - 0x0
      12'h18A: dout <= 8'b00000000; //  394 :   0 - 0x0
      12'h18B: dout <= 8'b00000000; //  395 :   0 - 0x0
      12'h18C: dout <= 8'b00000000; //  396 :   0 - 0x0
      12'h18D: dout <= 8'b00000000; //  397 :   0 - 0x0
      12'h18E: dout <= 8'b00000000; //  398 :   0 - 0x0
      12'h18F: dout <= 8'b00000000; //  399 :   0 - 0x0
      12'h190: dout <= 8'b00000000; //  400 :   0 - 0x0 -- Background 0x19
      12'h191: dout <= 8'b00000000; //  401 :   0 - 0x0
      12'h192: dout <= 8'b00001111; //  402 :  15 - 0xf
      12'h193: dout <= 8'b00010000; //  403 :  16 - 0x10
      12'h194: dout <= 8'b00010000; //  404 :  16 - 0x10
      12'h195: dout <= 8'b00001111; //  405 :  15 - 0xf
      12'h196: dout <= 8'b00000000; //  406 :   0 - 0x0
      12'h197: dout <= 8'b00000000; //  407 :   0 - 0x0
      12'h198: dout <= 8'b00000000; //  408 :   0 - 0x0 -- plane 1
      12'h199: dout <= 8'b00000000; //  409 :   0 - 0x0
      12'h19A: dout <= 8'b00000000; //  410 :   0 - 0x0
      12'h19B: dout <= 8'b00000000; //  411 :   0 - 0x0
      12'h19C: dout <= 8'b00000000; //  412 :   0 - 0x0
      12'h19D: dout <= 8'b00000000; //  413 :   0 - 0x0
      12'h19E: dout <= 8'b00000000; //  414 :   0 - 0x0
      12'h19F: dout <= 8'b00000000; //  415 :   0 - 0x0
      12'h1A0: dout <= 8'b00100100; //  416 :  36 - 0x24 -- Background 0x1a
      12'h1A1: dout <= 8'b00100100; //  417 :  36 - 0x24
      12'h1A2: dout <= 8'b00100100; //  418 :  36 - 0x24
      12'h1A3: dout <= 8'b00100100; //  419 :  36 - 0x24
      12'h1A4: dout <= 8'b00011000; //  420 :  24 - 0x18
      12'h1A5: dout <= 8'b00000000; //  421 :   0 - 0x0
      12'h1A6: dout <= 8'b00000000; //  422 :   0 - 0x0
      12'h1A7: dout <= 8'b00000000; //  423 :   0 - 0x0
      12'h1A8: dout <= 8'b00000000; //  424 :   0 - 0x0 -- plane 1
      12'h1A9: dout <= 8'b00000000; //  425 :   0 - 0x0
      12'h1AA: dout <= 8'b00000000; //  426 :   0 - 0x0
      12'h1AB: dout <= 8'b00000000; //  427 :   0 - 0x0
      12'h1AC: dout <= 8'b00000000; //  428 :   0 - 0x0
      12'h1AD: dout <= 8'b00000000; //  429 :   0 - 0x0
      12'h1AE: dout <= 8'b00000000; //  430 :   0 - 0x0
      12'h1AF: dout <= 8'b00000000; //  431 :   0 - 0x0
      12'h1B0: dout <= 8'b00000000; //  432 :   0 - 0x0 -- Background 0x1b
      12'h1B1: dout <= 8'b00000000; //  433 :   0 - 0x0
      12'h1B2: dout <= 8'b00000000; //  434 :   0 - 0x0
      12'h1B3: dout <= 8'b00011000; //  435 :  24 - 0x18
      12'h1B4: dout <= 8'b00100100; //  436 :  36 - 0x24
      12'h1B5: dout <= 8'b00100100; //  437 :  36 - 0x24
      12'h1B6: dout <= 8'b00100100; //  438 :  36 - 0x24
      12'h1B7: dout <= 8'b00100100; //  439 :  36 - 0x24
      12'h1B8: dout <= 8'b00000000; //  440 :   0 - 0x0 -- plane 1
      12'h1B9: dout <= 8'b00000000; //  441 :   0 - 0x0
      12'h1BA: dout <= 8'b00000000; //  442 :   0 - 0x0
      12'h1BB: dout <= 8'b00000000; //  443 :   0 - 0x0
      12'h1BC: dout <= 8'b00000000; //  444 :   0 - 0x0
      12'h1BD: dout <= 8'b00000000; //  445 :   0 - 0x0
      12'h1BE: dout <= 8'b00000000; //  446 :   0 - 0x0
      12'h1BF: dout <= 8'b00000000; //  447 :   0 - 0x0
      12'h1C0: dout <= 8'b00100100; //  448 :  36 - 0x24 -- Background 0x1c
      12'h1C1: dout <= 8'b00100100; //  449 :  36 - 0x24
      12'h1C2: dout <= 8'b11000100; //  450 : 196 - 0xc4
      12'h1C3: dout <= 8'b00000100; //  451 :   4 - 0x4
      12'h1C4: dout <= 8'b00001000; //  452 :   8 - 0x8
      12'h1C5: dout <= 8'b11110000; //  453 : 240 - 0xf0
      12'h1C6: dout <= 8'b00000000; //  454 :   0 - 0x0
      12'h1C7: dout <= 8'b00000000; //  455 :   0 - 0x0
      12'h1C8: dout <= 8'b00000000; //  456 :   0 - 0x0 -- plane 1
      12'h1C9: dout <= 8'b00000000; //  457 :   0 - 0x0
      12'h1CA: dout <= 8'b00000000; //  458 :   0 - 0x0
      12'h1CB: dout <= 8'b00000000; //  459 :   0 - 0x0
      12'h1CC: dout <= 8'b00000000; //  460 :   0 - 0x0
      12'h1CD: dout <= 8'b00000000; //  461 :   0 - 0x0
      12'h1CE: dout <= 8'b00000000; //  462 :   0 - 0x0
      12'h1CF: dout <= 8'b00000000; //  463 :   0 - 0x0
      12'h1D0: dout <= 8'b00000000; //  464 :   0 - 0x0 -- Background 0x1d
      12'h1D1: dout <= 8'b00000000; //  465 :   0 - 0x0
      12'h1D2: dout <= 8'b11110000; //  466 : 240 - 0xf0
      12'h1D3: dout <= 8'b00001000; //  467 :   8 - 0x8
      12'h1D4: dout <= 8'b00000100; //  468 :   4 - 0x4
      12'h1D5: dout <= 8'b11000100; //  469 : 196 - 0xc4
      12'h1D6: dout <= 8'b00100100; //  470 :  36 - 0x24
      12'h1D7: dout <= 8'b00100100; //  471 :  36 - 0x24
      12'h1D8: dout <= 8'b00000000; //  472 :   0 - 0x0 -- plane 1
      12'h1D9: dout <= 8'b00000000; //  473 :   0 - 0x0
      12'h1DA: dout <= 8'b00000000; //  474 :   0 - 0x0
      12'h1DB: dout <= 8'b00000000; //  475 :   0 - 0x0
      12'h1DC: dout <= 8'b00000000; //  476 :   0 - 0x0
      12'h1DD: dout <= 8'b00000000; //  477 :   0 - 0x0
      12'h1DE: dout <= 8'b00000000; //  478 :   0 - 0x0
      12'h1DF: dout <= 8'b00000000; //  479 :   0 - 0x0
      12'h1E0: dout <= 8'b00100100; //  480 :  36 - 0x24 -- Background 0x1e
      12'h1E1: dout <= 8'b00100100; //  481 :  36 - 0x24
      12'h1E2: dout <= 8'b00100011; //  482 :  35 - 0x23
      12'h1E3: dout <= 8'b00100000; //  483 :  32 - 0x20
      12'h1E4: dout <= 8'b00010000; //  484 :  16 - 0x10
      12'h1E5: dout <= 8'b00001111; //  485 :  15 - 0xf
      12'h1E6: dout <= 8'b00000000; //  486 :   0 - 0x0
      12'h1E7: dout <= 8'b00000000; //  487 :   0 - 0x0
      12'h1E8: dout <= 8'b00000000; //  488 :   0 - 0x0 -- plane 1
      12'h1E9: dout <= 8'b00000000; //  489 :   0 - 0x0
      12'h1EA: dout <= 8'b00000000; //  490 :   0 - 0x0
      12'h1EB: dout <= 8'b00000000; //  491 :   0 - 0x0
      12'h1EC: dout <= 8'b00000000; //  492 :   0 - 0x0
      12'h1ED: dout <= 8'b00000000; //  493 :   0 - 0x0
      12'h1EE: dout <= 8'b00000000; //  494 :   0 - 0x0
      12'h1EF: dout <= 8'b00000000; //  495 :   0 - 0x0
      12'h1F0: dout <= 8'b00000000; //  496 :   0 - 0x0 -- Background 0x1f
      12'h1F1: dout <= 8'b00000000; //  497 :   0 - 0x0
      12'h1F2: dout <= 8'b00001111; //  498 :  15 - 0xf
      12'h1F3: dout <= 8'b00010000; //  499 :  16 - 0x10
      12'h1F4: dout <= 8'b00100000; //  500 :  32 - 0x20
      12'h1F5: dout <= 8'b00100011; //  501 :  35 - 0x23
      12'h1F6: dout <= 8'b00100100; //  502 :  36 - 0x24
      12'h1F7: dout <= 8'b00100100; //  503 :  36 - 0x24
      12'h1F8: dout <= 8'b00000000; //  504 :   0 - 0x0 -- plane 1
      12'h1F9: dout <= 8'b00000000; //  505 :   0 - 0x0
      12'h1FA: dout <= 8'b00000000; //  506 :   0 - 0x0
      12'h1FB: dout <= 8'b00000000; //  507 :   0 - 0x0
      12'h1FC: dout <= 8'b00000000; //  508 :   0 - 0x0
      12'h1FD: dout <= 8'b00000000; //  509 :   0 - 0x0
      12'h1FE: dout <= 8'b00000000; //  510 :   0 - 0x0
      12'h1FF: dout <= 8'b00000000; //  511 :   0 - 0x0
      12'h200: dout <= 8'b00000000; //  512 :   0 - 0x0 -- Background 0x20
      12'h201: dout <= 8'b00000000; //  513 :   0 - 0x0
      12'h202: dout <= 8'b00000000; //  514 :   0 - 0x0
      12'h203: dout <= 8'b00000000; //  515 :   0 - 0x0
      12'h204: dout <= 8'b00000000; //  516 :   0 - 0x0
      12'h205: dout <= 8'b00000000; //  517 :   0 - 0x0
      12'h206: dout <= 8'b00000000; //  518 :   0 - 0x0
      12'h207: dout <= 8'b00000000; //  519 :   0 - 0x0
      12'h208: dout <= 8'b00000000; //  520 :   0 - 0x0 -- plane 1
      12'h209: dout <= 8'b00000000; //  521 :   0 - 0x0
      12'h20A: dout <= 8'b00000000; //  522 :   0 - 0x0
      12'h20B: dout <= 8'b00000000; //  523 :   0 - 0x0
      12'h20C: dout <= 8'b00000000; //  524 :   0 - 0x0
      12'h20D: dout <= 8'b00000000; //  525 :   0 - 0x0
      12'h20E: dout <= 8'b00000000; //  526 :   0 - 0x0
      12'h20F: dout <= 8'b00000000; //  527 :   0 - 0x0
      12'h210: dout <= 8'b00000000; //  528 :   0 - 0x0 -- Background 0x21
      12'h211: dout <= 8'b00000000; //  529 :   0 - 0x0
      12'h212: dout <= 8'b11110000; //  530 : 240 - 0xf0
      12'h213: dout <= 8'b00001000; //  531 :   8 - 0x8
      12'h214: dout <= 8'b00001000; //  532 :   8 - 0x8
      12'h215: dout <= 8'b11110000; //  533 : 240 - 0xf0
      12'h216: dout <= 8'b00000000; //  534 :   0 - 0x0
      12'h217: dout <= 8'b00000000; //  535 :   0 - 0x0
      12'h218: dout <= 8'b00001111; //  536 :  15 - 0xf -- plane 1
      12'h219: dout <= 8'b00001111; //  537 :  15 - 0xf
      12'h21A: dout <= 8'b00001111; //  538 :  15 - 0xf
      12'h21B: dout <= 8'b00000111; //  539 :   7 - 0x7
      12'h21C: dout <= 8'b00000111; //  540 :   7 - 0x7
      12'h21D: dout <= 8'b00001111; //  541 :  15 - 0xf
      12'h21E: dout <= 8'b00001111; //  542 :  15 - 0xf
      12'h21F: dout <= 8'b00001111; //  543 :  15 - 0xf
      12'h220: dout <= 8'b00000000; //  544 :   0 - 0x0 -- Background 0x22
      12'h221: dout <= 8'b00000000; //  545 :   0 - 0x0
      12'h222: dout <= 8'b00001111; //  546 :  15 - 0xf
      12'h223: dout <= 8'b00010000; //  547 :  16 - 0x10
      12'h224: dout <= 8'b00010000; //  548 :  16 - 0x10
      12'h225: dout <= 8'b00001111; //  549 :  15 - 0xf
      12'h226: dout <= 8'b00000000; //  550 :   0 - 0x0
      12'h227: dout <= 8'b00000000; //  551 :   0 - 0x0
      12'h228: dout <= 8'b11110000; //  552 : 240 - 0xf0 -- plane 1
      12'h229: dout <= 8'b11110000; //  553 : 240 - 0xf0
      12'h22A: dout <= 8'b11110000; //  554 : 240 - 0xf0
      12'h22B: dout <= 8'b11100000; //  555 : 224 - 0xe0
      12'h22C: dout <= 8'b11100000; //  556 : 224 - 0xe0
      12'h22D: dout <= 8'b11110000; //  557 : 240 - 0xf0
      12'h22E: dout <= 8'b11110000; //  558 : 240 - 0xf0
      12'h22F: dout <= 8'b11110000; //  559 : 240 - 0xf0
      12'h230: dout <= 8'b11111111; //  560 : 255 - 0xff -- Background 0x23
      12'h231: dout <= 8'b11111111; //  561 : 255 - 0xff
      12'h232: dout <= 8'b11100001; //  562 : 225 - 0xe1
      12'h233: dout <= 8'b11100001; //  563 : 225 - 0xe1
      12'h234: dout <= 8'b11100001; //  564 : 225 - 0xe1
      12'h235: dout <= 8'b11100001; //  565 : 225 - 0xe1
      12'h236: dout <= 8'b11100001; //  566 : 225 - 0xe1
      12'h237: dout <= 8'b11100001; //  567 : 225 - 0xe1
      12'h238: dout <= 8'b11111111; //  568 : 255 - 0xff -- plane 1
      12'h239: dout <= 8'b11111111; //  569 : 255 - 0xff
      12'h23A: dout <= 8'b11100001; //  570 : 225 - 0xe1
      12'h23B: dout <= 8'b11100001; //  571 : 225 - 0xe1
      12'h23C: dout <= 8'b11100001; //  572 : 225 - 0xe1
      12'h23D: dout <= 8'b11100001; //  573 : 225 - 0xe1
      12'h23E: dout <= 8'b11100001; //  574 : 225 - 0xe1
      12'h23F: dout <= 8'b11100001; //  575 : 225 - 0xe1
      12'h240: dout <= 8'b10000111; //  576 : 135 - 0x87 -- Background 0x24
      12'h241: dout <= 8'b11000111; //  577 : 199 - 0xc7
      12'h242: dout <= 8'b11000000; //  578 : 192 - 0xc0
      12'h243: dout <= 8'b11000111; //  579 : 199 - 0xc7
      12'h244: dout <= 8'b11001111; //  580 : 207 - 0xcf
      12'h245: dout <= 8'b11001110; //  581 : 206 - 0xce
      12'h246: dout <= 8'b11001111; //  582 : 207 - 0xcf
      12'h247: dout <= 8'b11000111; //  583 : 199 - 0xc7
      12'h248: dout <= 8'b10000111; //  584 : 135 - 0x87 -- plane 1
      12'h249: dout <= 8'b11000111; //  585 : 199 - 0xc7
      12'h24A: dout <= 8'b11000000; //  586 : 192 - 0xc0
      12'h24B: dout <= 8'b11000111; //  587 : 199 - 0xc7
      12'h24C: dout <= 8'b11001111; //  588 : 207 - 0xcf
      12'h24D: dout <= 8'b11001110; //  589 : 206 - 0xce
      12'h24E: dout <= 8'b11001111; //  590 : 207 - 0xcf
      12'h24F: dout <= 8'b11000111; //  591 : 199 - 0xc7
      12'h250: dout <= 8'b11111000; //  592 : 248 - 0xf8 -- Background 0x25
      12'h251: dout <= 8'b11111100; //  593 : 252 - 0xfc
      12'h252: dout <= 8'b00011100; //  594 :  28 - 0x1c
      12'h253: dout <= 8'b11111100; //  595 : 252 - 0xfc
      12'h254: dout <= 8'b11111100; //  596 : 252 - 0xfc
      12'h255: dout <= 8'b00011100; //  597 :  28 - 0x1c
      12'h256: dout <= 8'b11111100; //  598 : 252 - 0xfc
      12'h257: dout <= 8'b11111100; //  599 : 252 - 0xfc
      12'h258: dout <= 8'b11111000; //  600 : 248 - 0xf8 -- plane 1
      12'h259: dout <= 8'b11111100; //  601 : 252 - 0xfc
      12'h25A: dout <= 8'b00011100; //  602 :  28 - 0x1c
      12'h25B: dout <= 8'b11111100; //  603 : 252 - 0xfc
      12'h25C: dout <= 8'b11111100; //  604 : 252 - 0xfc
      12'h25D: dout <= 8'b00011100; //  605 :  28 - 0x1c
      12'h25E: dout <= 8'b11111100; //  606 : 252 - 0xfc
      12'h25F: dout <= 8'b11111100; //  607 : 252 - 0xfc
      12'h260: dout <= 8'b11111111; //  608 : 255 - 0xff -- Background 0x26
      12'h261: dout <= 8'b11111111; //  609 : 255 - 0xff
      12'h262: dout <= 8'b11100111; //  610 : 231 - 0xe7
      12'h263: dout <= 8'b11100111; //  611 : 231 - 0xe7
      12'h264: dout <= 8'b11100111; //  612 : 231 - 0xe7
      12'h265: dout <= 8'b11100111; //  613 : 231 - 0xe7
      12'h266: dout <= 8'b11100111; //  614 : 231 - 0xe7
      12'h267: dout <= 8'b11100111; //  615 : 231 - 0xe7
      12'h268: dout <= 8'b11111111; //  616 : 255 - 0xff -- plane 1
      12'h269: dout <= 8'b11111111; //  617 : 255 - 0xff
      12'h26A: dout <= 8'b11100111; //  618 : 231 - 0xe7
      12'h26B: dout <= 8'b11100111; //  619 : 231 - 0xe7
      12'h26C: dout <= 8'b11100111; //  620 : 231 - 0xe7
      12'h26D: dout <= 8'b11100111; //  621 : 231 - 0xe7
      12'h26E: dout <= 8'b11100111; //  622 : 231 - 0xe7
      12'h26F: dout <= 8'b11100111; //  623 : 231 - 0xe7
      12'h270: dout <= 8'b11110000; //  624 : 240 - 0xf0 -- Background 0x27
      12'h271: dout <= 8'b11111001; //  625 : 249 - 0xf9
      12'h272: dout <= 8'b00111001; //  626 :  57 - 0x39
      12'h273: dout <= 8'b00111001; //  627 :  57 - 0x39
      12'h274: dout <= 8'b00111001; //  628 :  57 - 0x39
      12'h275: dout <= 8'b00111001; //  629 :  57 - 0x39
      12'h276: dout <= 8'b00111001; //  630 :  57 - 0x39
      12'h277: dout <= 8'b00111000; //  631 :  56 - 0x38
      12'h278: dout <= 8'b11110000; //  632 : 240 - 0xf0 -- plane 1
      12'h279: dout <= 8'b11111001; //  633 : 249 - 0xf9
      12'h27A: dout <= 8'b00111001; //  634 :  57 - 0x39
      12'h27B: dout <= 8'b00111001; //  635 :  57 - 0x39
      12'h27C: dout <= 8'b00111001; //  636 :  57 - 0x39
      12'h27D: dout <= 8'b00111001; //  637 :  57 - 0x39
      12'h27E: dout <= 8'b00111001; //  638 :  57 - 0x39
      12'h27F: dout <= 8'b00111000; //  639 :  56 - 0x38
      12'h280: dout <= 8'b11111111; //  640 : 255 - 0xff -- Background 0x28
      12'h281: dout <= 8'b11111111; //  641 : 255 - 0xff
      12'h282: dout <= 8'b11000000; //  642 : 192 - 0xc0
      12'h283: dout <= 8'b11000000; //  643 : 192 - 0xc0
      12'h284: dout <= 8'b11000000; //  644 : 192 - 0xc0
      12'h285: dout <= 8'b11000000; //  645 : 192 - 0xc0
      12'h286: dout <= 8'b11111111; //  646 : 255 - 0xff
      12'h287: dout <= 8'b11111111; //  647 : 255 - 0xff
      12'h288: dout <= 8'b11111111; //  648 : 255 - 0xff -- plane 1
      12'h289: dout <= 8'b11111111; //  649 : 255 - 0xff
      12'h28A: dout <= 8'b11000000; //  650 : 192 - 0xc0
      12'h28B: dout <= 8'b11000000; //  651 : 192 - 0xc0
      12'h28C: dout <= 8'b11000000; //  652 : 192 - 0xc0
      12'h28D: dout <= 8'b11000000; //  653 : 192 - 0xc0
      12'h28E: dout <= 8'b11111111; //  654 : 255 - 0xff
      12'h28F: dout <= 8'b11111111; //  655 : 255 - 0xff
      12'h290: dout <= 8'b00011111; //  656 :  31 - 0x1f -- Background 0x29
      12'h291: dout <= 8'b00111111; //  657 :  63 - 0x3f
      12'h292: dout <= 8'b00110000; //  658 :  48 - 0x30
      12'h293: dout <= 8'b00110000; //  659 :  48 - 0x30
      12'h294: dout <= 8'b00110000; //  660 :  48 - 0x30
      12'h295: dout <= 8'b00110000; //  661 :  48 - 0x30
      12'h296: dout <= 8'b00111111; //  662 :  63 - 0x3f
      12'h297: dout <= 8'b00011111; //  663 :  31 - 0x1f
      12'h298: dout <= 8'b00011111; //  664 :  31 - 0x1f -- plane 1
      12'h299: dout <= 8'b00111111; //  665 :  63 - 0x3f
      12'h29A: dout <= 8'b00110000; //  666 :  48 - 0x30
      12'h29B: dout <= 8'b00110000; //  667 :  48 - 0x30
      12'h29C: dout <= 8'b00110000; //  668 :  48 - 0x30
      12'h29D: dout <= 8'b00110000; //  669 :  48 - 0x30
      12'h29E: dout <= 8'b00111111; //  670 :  63 - 0x3f
      12'h29F: dout <= 8'b00011111; //  671 :  31 - 0x1f
      12'h2A0: dout <= 8'b11100011; //  672 : 227 - 0xe3 -- Background 0x2a
      12'h2A1: dout <= 8'b11110011; //  673 : 243 - 0xf3
      12'h2A2: dout <= 8'b01110000; //  674 : 112 - 0x70
      12'h2A3: dout <= 8'b01110000; //  675 : 112 - 0x70
      12'h2A4: dout <= 8'b01110000; //  676 : 112 - 0x70
      12'h2A5: dout <= 8'b01110000; //  677 : 112 - 0x70
      12'h2A6: dout <= 8'b11110000; //  678 : 240 - 0xf0
      12'h2A7: dout <= 8'b11100000; //  679 : 224 - 0xe0
      12'h2A8: dout <= 8'b11100011; //  680 : 227 - 0xe3 -- plane 1
      12'h2A9: dout <= 8'b11110011; //  681 : 243 - 0xf3
      12'h2AA: dout <= 8'b01110000; //  682 : 112 - 0x70
      12'h2AB: dout <= 8'b01110000; //  683 : 112 - 0x70
      12'h2AC: dout <= 8'b01110000; //  684 : 112 - 0x70
      12'h2AD: dout <= 8'b01110000; //  685 : 112 - 0x70
      12'h2AE: dout <= 8'b11110000; //  686 : 240 - 0xf0
      12'h2AF: dout <= 8'b11100000; //  687 : 224 - 0xe0
      12'h2B0: dout <= 8'b11111110; //  688 : 254 - 0xfe -- Background 0x2b
      12'h2B1: dout <= 8'b11111110; //  689 : 254 - 0xfe
      12'h2B2: dout <= 8'b01110000; //  690 : 112 - 0x70
      12'h2B3: dout <= 8'b01110000; //  691 : 112 - 0x70
      12'h2B4: dout <= 8'b01110000; //  692 : 112 - 0x70
      12'h2B5: dout <= 8'b01110000; //  693 : 112 - 0x70
      12'h2B6: dout <= 8'b01110000; //  694 : 112 - 0x70
      12'h2B7: dout <= 8'b01110000; //  695 : 112 - 0x70
      12'h2B8: dout <= 8'b11111110; //  696 : 254 - 0xfe -- plane 1
      12'h2B9: dout <= 8'b11111110; //  697 : 254 - 0xfe
      12'h2BA: dout <= 8'b01110000; //  698 : 112 - 0x70
      12'h2BB: dout <= 8'b01110000; //  699 : 112 - 0x70
      12'h2BC: dout <= 8'b01110000; //  700 : 112 - 0x70
      12'h2BD: dout <= 8'b01110000; //  701 : 112 - 0x70
      12'h2BE: dout <= 8'b01110000; //  702 : 112 - 0x70
      12'h2BF: dout <= 8'b01110000; //  703 : 112 - 0x70
      12'h2C0: dout <= 8'b00000000; //  704 :   0 - 0x0 -- Background 0x2c
      12'h2C1: dout <= 8'b00000000; //  705 :   0 - 0x0
      12'h2C2: dout <= 8'b00000000; //  706 :   0 - 0x0
      12'h2C3: dout <= 8'b00000000; //  707 :   0 - 0x0
      12'h2C4: dout <= 8'b11111111; //  708 : 255 - 0xff
      12'h2C5: dout <= 8'b00000000; //  709 :   0 - 0x0
      12'h2C6: dout <= 8'b00000000; //  710 :   0 - 0x0
      12'h2C7: dout <= 8'b00000000; //  711 :   0 - 0x0
      12'h2C8: dout <= 8'b00000000; //  712 :   0 - 0x0 -- plane 1
      12'h2C9: dout <= 8'b00000000; //  713 :   0 - 0x0
      12'h2CA: dout <= 8'b00000000; //  714 :   0 - 0x0
      12'h2CB: dout <= 8'b00000000; //  715 :   0 - 0x0
      12'h2CC: dout <= 8'b00000000; //  716 :   0 - 0x0
      12'h2CD: dout <= 8'b00000000; //  717 :   0 - 0x0
      12'h2CE: dout <= 8'b00000000; //  718 :   0 - 0x0
      12'h2CF: dout <= 8'b00000000; //  719 :   0 - 0x0
      12'h2D0: dout <= 8'b00000000; //  720 :   0 - 0x0 -- Background 0x2d
      12'h2D1: dout <= 8'b00000000; //  721 :   0 - 0x0
      12'h2D2: dout <= 8'b00000000; //  722 :   0 - 0x0
      12'h2D3: dout <= 8'b00000000; //  723 :   0 - 0x0
      12'h2D4: dout <= 8'b00000000; //  724 :   0 - 0x0
      12'h2D5: dout <= 8'b00000000; //  725 :   0 - 0x0
      12'h2D6: dout <= 8'b00000000; //  726 :   0 - 0x0
      12'h2D7: dout <= 8'b00000000; //  727 :   0 - 0x0
      12'h2D8: dout <= 8'b11111111; //  728 : 255 - 0xff -- plane 1
      12'h2D9: dout <= 8'b11111111; //  729 : 255 - 0xff
      12'h2DA: dout <= 8'b11111111; //  730 : 255 - 0xff
      12'h2DB: dout <= 8'b11111111; //  731 : 255 - 0xff
      12'h2DC: dout <= 8'b11111111; //  732 : 255 - 0xff
      12'h2DD: dout <= 8'b11111111; //  733 : 255 - 0xff
      12'h2DE: dout <= 8'b11111111; //  734 : 255 - 0xff
      12'h2DF: dout <= 8'b11111111; //  735 : 255 - 0xff
      12'h2E0: dout <= 8'b00000000; //  736 :   0 - 0x0 -- Background 0x2e
      12'h2E1: dout <= 8'b00000000; //  737 :   0 - 0x0
      12'h2E2: dout <= 8'b00000000; //  738 :   0 - 0x0
      12'h2E3: dout <= 8'b00011000; //  739 :  24 - 0x18
      12'h2E4: dout <= 8'b00011000; //  740 :  24 - 0x18
      12'h2E5: dout <= 8'b00000000; //  741 :   0 - 0x0
      12'h2E6: dout <= 8'b00000000; //  742 :   0 - 0x0
      12'h2E7: dout <= 8'b00000000; //  743 :   0 - 0x0
      12'h2E8: dout <= 8'b00000000; //  744 :   0 - 0x0 -- plane 1
      12'h2E9: dout <= 8'b00000000; //  745 :   0 - 0x0
      12'h2EA: dout <= 8'b00000000; //  746 :   0 - 0x0
      12'h2EB: dout <= 8'b00000000; //  747 :   0 - 0x0
      12'h2EC: dout <= 8'b00000000; //  748 :   0 - 0x0
      12'h2ED: dout <= 8'b00000000; //  749 :   0 - 0x0
      12'h2EE: dout <= 8'b00000000; //  750 :   0 - 0x0
      12'h2EF: dout <= 8'b00000000; //  751 :   0 - 0x0
      12'h2F0: dout <= 8'b00000000; //  752 :   0 - 0x0 -- Background 0x2f
      12'h2F1: dout <= 8'b00000000; //  753 :   0 - 0x0
      12'h2F2: dout <= 8'b00000000; //  754 :   0 - 0x0
      12'h2F3: dout <= 8'b00000000; //  755 :   0 - 0x0
      12'h2F4: dout <= 8'b00000000; //  756 :   0 - 0x0
      12'h2F5: dout <= 8'b00000000; //  757 :   0 - 0x0
      12'h2F6: dout <= 8'b00000000; //  758 :   0 - 0x0
      12'h2F7: dout <= 8'b00000000; //  759 :   0 - 0x0
      12'h2F8: dout <= 8'b00000000; //  760 :   0 - 0x0 -- plane 1
      12'h2F9: dout <= 8'b00000000; //  761 :   0 - 0x0
      12'h2FA: dout <= 8'b00000000; //  762 :   0 - 0x0
      12'h2FB: dout <= 8'b00011000; //  763 :  24 - 0x18
      12'h2FC: dout <= 8'b00011000; //  764 :  24 - 0x18
      12'h2FD: dout <= 8'b00000000; //  765 :   0 - 0x0
      12'h2FE: dout <= 8'b00000000; //  766 :   0 - 0x0
      12'h2FF: dout <= 8'b00000000; //  767 :   0 - 0x0
      12'h300: dout <= 8'b00011100; //  768 :  28 - 0x1c -- Background 0x30
      12'h301: dout <= 8'b00100110; //  769 :  38 - 0x26
      12'h302: dout <= 8'b01100011; //  770 :  99 - 0x63
      12'h303: dout <= 8'b01100011; //  771 :  99 - 0x63
      12'h304: dout <= 8'b01100011; //  772 :  99 - 0x63
      12'h305: dout <= 8'b00110010; //  773 :  50 - 0x32
      12'h306: dout <= 8'b00011100; //  774 :  28 - 0x1c
      12'h307: dout <= 8'b00000000; //  775 :   0 - 0x0
      12'h308: dout <= 8'b00000000; //  776 :   0 - 0x0 -- plane 1
      12'h309: dout <= 8'b00000000; //  777 :   0 - 0x0
      12'h30A: dout <= 8'b00000000; //  778 :   0 - 0x0
      12'h30B: dout <= 8'b00000000; //  779 :   0 - 0x0
      12'h30C: dout <= 8'b00000000; //  780 :   0 - 0x0
      12'h30D: dout <= 8'b00000000; //  781 :   0 - 0x0
      12'h30E: dout <= 8'b00000000; //  782 :   0 - 0x0
      12'h30F: dout <= 8'b00000000; //  783 :   0 - 0x0
      12'h310: dout <= 8'b00001100; //  784 :  12 - 0xc -- Background 0x31
      12'h311: dout <= 8'b00011100; //  785 :  28 - 0x1c
      12'h312: dout <= 8'b00001100; //  786 :  12 - 0xc
      12'h313: dout <= 8'b00001100; //  787 :  12 - 0xc
      12'h314: dout <= 8'b00001100; //  788 :  12 - 0xc
      12'h315: dout <= 8'b00001100; //  789 :  12 - 0xc
      12'h316: dout <= 8'b00111111; //  790 :  63 - 0x3f
      12'h317: dout <= 8'b00000000; //  791 :   0 - 0x0
      12'h318: dout <= 8'b00000000; //  792 :   0 - 0x0 -- plane 1
      12'h319: dout <= 8'b00000000; //  793 :   0 - 0x0
      12'h31A: dout <= 8'b00000000; //  794 :   0 - 0x0
      12'h31B: dout <= 8'b00000000; //  795 :   0 - 0x0
      12'h31C: dout <= 8'b00000000; //  796 :   0 - 0x0
      12'h31D: dout <= 8'b00000000; //  797 :   0 - 0x0
      12'h31E: dout <= 8'b00000000; //  798 :   0 - 0x0
      12'h31F: dout <= 8'b00000000; //  799 :   0 - 0x0
      12'h320: dout <= 8'b00111110; //  800 :  62 - 0x3e -- Background 0x32
      12'h321: dout <= 8'b01100011; //  801 :  99 - 0x63
      12'h322: dout <= 8'b00000111; //  802 :   7 - 0x7
      12'h323: dout <= 8'b00011110; //  803 :  30 - 0x1e
      12'h324: dout <= 8'b00111100; //  804 :  60 - 0x3c
      12'h325: dout <= 8'b01110000; //  805 : 112 - 0x70
      12'h326: dout <= 8'b01111111; //  806 : 127 - 0x7f
      12'h327: dout <= 8'b00000000; //  807 :   0 - 0x0
      12'h328: dout <= 8'b00000000; //  808 :   0 - 0x0 -- plane 1
      12'h329: dout <= 8'b00000000; //  809 :   0 - 0x0
      12'h32A: dout <= 8'b00000000; //  810 :   0 - 0x0
      12'h32B: dout <= 8'b00000000; //  811 :   0 - 0x0
      12'h32C: dout <= 8'b00000000; //  812 :   0 - 0x0
      12'h32D: dout <= 8'b00000000; //  813 :   0 - 0x0
      12'h32E: dout <= 8'b00000000; //  814 :   0 - 0x0
      12'h32F: dout <= 8'b00000000; //  815 :   0 - 0x0
      12'h330: dout <= 8'b00111111; //  816 :  63 - 0x3f -- Background 0x33
      12'h331: dout <= 8'b00000110; //  817 :   6 - 0x6
      12'h332: dout <= 8'b00001100; //  818 :  12 - 0xc
      12'h333: dout <= 8'b00011110; //  819 :  30 - 0x1e
      12'h334: dout <= 8'b00000011; //  820 :   3 - 0x3
      12'h335: dout <= 8'b01100011; //  821 :  99 - 0x63
      12'h336: dout <= 8'b00111110; //  822 :  62 - 0x3e
      12'h337: dout <= 8'b00000000; //  823 :   0 - 0x0
      12'h338: dout <= 8'b00000000; //  824 :   0 - 0x0 -- plane 1
      12'h339: dout <= 8'b00000000; //  825 :   0 - 0x0
      12'h33A: dout <= 8'b00000000; //  826 :   0 - 0x0
      12'h33B: dout <= 8'b00000000; //  827 :   0 - 0x0
      12'h33C: dout <= 8'b00000000; //  828 :   0 - 0x0
      12'h33D: dout <= 8'b00000000; //  829 :   0 - 0x0
      12'h33E: dout <= 8'b00000000; //  830 :   0 - 0x0
      12'h33F: dout <= 8'b00000000; //  831 :   0 - 0x0
      12'h340: dout <= 8'b00001110; //  832 :  14 - 0xe -- Background 0x34
      12'h341: dout <= 8'b00011110; //  833 :  30 - 0x1e
      12'h342: dout <= 8'b00110110; //  834 :  54 - 0x36
      12'h343: dout <= 8'b01100110; //  835 : 102 - 0x66
      12'h344: dout <= 8'b01111111; //  836 : 127 - 0x7f
      12'h345: dout <= 8'b00000110; //  837 :   6 - 0x6
      12'h346: dout <= 8'b00000110; //  838 :   6 - 0x6
      12'h347: dout <= 8'b00000000; //  839 :   0 - 0x0
      12'h348: dout <= 8'b00000000; //  840 :   0 - 0x0 -- plane 1
      12'h349: dout <= 8'b00000000; //  841 :   0 - 0x0
      12'h34A: dout <= 8'b00000000; //  842 :   0 - 0x0
      12'h34B: dout <= 8'b00000000; //  843 :   0 - 0x0
      12'h34C: dout <= 8'b00000000; //  844 :   0 - 0x0
      12'h34D: dout <= 8'b00000000; //  845 :   0 - 0x0
      12'h34E: dout <= 8'b00000000; //  846 :   0 - 0x0
      12'h34F: dout <= 8'b00000000; //  847 :   0 - 0x0
      12'h350: dout <= 8'b01111110; //  848 : 126 - 0x7e -- Background 0x35
      12'h351: dout <= 8'b01100000; //  849 :  96 - 0x60
      12'h352: dout <= 8'b01111110; //  850 : 126 - 0x7e
      12'h353: dout <= 8'b00000011; //  851 :   3 - 0x3
      12'h354: dout <= 8'b00000011; //  852 :   3 - 0x3
      12'h355: dout <= 8'b01100011; //  853 :  99 - 0x63
      12'h356: dout <= 8'b00111110; //  854 :  62 - 0x3e
      12'h357: dout <= 8'b00000000; //  855 :   0 - 0x0
      12'h358: dout <= 8'b00000000; //  856 :   0 - 0x0 -- plane 1
      12'h359: dout <= 8'b00000000; //  857 :   0 - 0x0
      12'h35A: dout <= 8'b00000000; //  858 :   0 - 0x0
      12'h35B: dout <= 8'b00000000; //  859 :   0 - 0x0
      12'h35C: dout <= 8'b00000000; //  860 :   0 - 0x0
      12'h35D: dout <= 8'b00000000; //  861 :   0 - 0x0
      12'h35E: dout <= 8'b00000000; //  862 :   0 - 0x0
      12'h35F: dout <= 8'b00000000; //  863 :   0 - 0x0
      12'h360: dout <= 8'b00011110; //  864 :  30 - 0x1e -- Background 0x36
      12'h361: dout <= 8'b00110000; //  865 :  48 - 0x30
      12'h362: dout <= 8'b01100000; //  866 :  96 - 0x60
      12'h363: dout <= 8'b01111110; //  867 : 126 - 0x7e
      12'h364: dout <= 8'b01100011; //  868 :  99 - 0x63
      12'h365: dout <= 8'b01100011; //  869 :  99 - 0x63
      12'h366: dout <= 8'b00111110; //  870 :  62 - 0x3e
      12'h367: dout <= 8'b00000000; //  871 :   0 - 0x0
      12'h368: dout <= 8'b00000000; //  872 :   0 - 0x0 -- plane 1
      12'h369: dout <= 8'b00000000; //  873 :   0 - 0x0
      12'h36A: dout <= 8'b00000000; //  874 :   0 - 0x0
      12'h36B: dout <= 8'b00000000; //  875 :   0 - 0x0
      12'h36C: dout <= 8'b00000000; //  876 :   0 - 0x0
      12'h36D: dout <= 8'b00000000; //  877 :   0 - 0x0
      12'h36E: dout <= 8'b00000000; //  878 :   0 - 0x0
      12'h36F: dout <= 8'b00000000; //  879 :   0 - 0x0
      12'h370: dout <= 8'b01111111; //  880 : 127 - 0x7f -- Background 0x37
      12'h371: dout <= 8'b01100011; //  881 :  99 - 0x63
      12'h372: dout <= 8'b00000110; //  882 :   6 - 0x6
      12'h373: dout <= 8'b00001100; //  883 :  12 - 0xc
      12'h374: dout <= 8'b00011000; //  884 :  24 - 0x18
      12'h375: dout <= 8'b00011000; //  885 :  24 - 0x18
      12'h376: dout <= 8'b00011000; //  886 :  24 - 0x18
      12'h377: dout <= 8'b00000000; //  887 :   0 - 0x0
      12'h378: dout <= 8'b00000000; //  888 :   0 - 0x0 -- plane 1
      12'h379: dout <= 8'b00000000; //  889 :   0 - 0x0
      12'h37A: dout <= 8'b00000000; //  890 :   0 - 0x0
      12'h37B: dout <= 8'b00000000; //  891 :   0 - 0x0
      12'h37C: dout <= 8'b00000000; //  892 :   0 - 0x0
      12'h37D: dout <= 8'b00000000; //  893 :   0 - 0x0
      12'h37E: dout <= 8'b00000000; //  894 :   0 - 0x0
      12'h37F: dout <= 8'b00000000; //  895 :   0 - 0x0
      12'h380: dout <= 8'b00111100; //  896 :  60 - 0x3c -- Background 0x38
      12'h381: dout <= 8'b01100010; //  897 :  98 - 0x62
      12'h382: dout <= 8'b01110010; //  898 : 114 - 0x72
      12'h383: dout <= 8'b00111100; //  899 :  60 - 0x3c
      12'h384: dout <= 8'b01001111; //  900 :  79 - 0x4f
      12'h385: dout <= 8'b01000011; //  901 :  67 - 0x43
      12'h386: dout <= 8'b00111110; //  902 :  62 - 0x3e
      12'h387: dout <= 8'b00000000; //  903 :   0 - 0x0
      12'h388: dout <= 8'b00000000; //  904 :   0 - 0x0 -- plane 1
      12'h389: dout <= 8'b00000000; //  905 :   0 - 0x0
      12'h38A: dout <= 8'b00000000; //  906 :   0 - 0x0
      12'h38B: dout <= 8'b00000000; //  907 :   0 - 0x0
      12'h38C: dout <= 8'b00000000; //  908 :   0 - 0x0
      12'h38D: dout <= 8'b00000000; //  909 :   0 - 0x0
      12'h38E: dout <= 8'b00000000; //  910 :   0 - 0x0
      12'h38F: dout <= 8'b00000000; //  911 :   0 - 0x0
      12'h390: dout <= 8'b00111110; //  912 :  62 - 0x3e -- Background 0x39
      12'h391: dout <= 8'b01100011; //  913 :  99 - 0x63
      12'h392: dout <= 8'b01100011; //  914 :  99 - 0x63
      12'h393: dout <= 8'b00111111; //  915 :  63 - 0x3f
      12'h394: dout <= 8'b00000011; //  916 :   3 - 0x3
      12'h395: dout <= 8'b00000110; //  917 :   6 - 0x6
      12'h396: dout <= 8'b00111100; //  918 :  60 - 0x3c
      12'h397: dout <= 8'b00000000; //  919 :   0 - 0x0
      12'h398: dout <= 8'b00000000; //  920 :   0 - 0x0 -- plane 1
      12'h399: dout <= 8'b00000000; //  921 :   0 - 0x0
      12'h39A: dout <= 8'b00000000; //  922 :   0 - 0x0
      12'h39B: dout <= 8'b00000000; //  923 :   0 - 0x0
      12'h39C: dout <= 8'b00000000; //  924 :   0 - 0x0
      12'h39D: dout <= 8'b00000000; //  925 :   0 - 0x0
      12'h39E: dout <= 8'b00000000; //  926 :   0 - 0x0
      12'h39F: dout <= 8'b00000000; //  927 :   0 - 0x0
      12'h3A0: dout <= 8'b00000000; //  928 :   0 - 0x0 -- Background 0x3a
      12'h3A1: dout <= 8'b00000000; //  929 :   0 - 0x0
      12'h3A2: dout <= 8'b00000000; //  930 :   0 - 0x0
      12'h3A3: dout <= 8'b01111110; //  931 : 126 - 0x7e
      12'h3A4: dout <= 8'b00000000; //  932 :   0 - 0x0
      12'h3A5: dout <= 8'b00000000; //  933 :   0 - 0x0
      12'h3A6: dout <= 8'b00000000; //  934 :   0 - 0x0
      12'h3A7: dout <= 8'b00000000; //  935 :   0 - 0x0
      12'h3A8: dout <= 8'b00000000; //  936 :   0 - 0x0 -- plane 1
      12'h3A9: dout <= 8'b00000000; //  937 :   0 - 0x0
      12'h3AA: dout <= 8'b00000000; //  938 :   0 - 0x0
      12'h3AB: dout <= 8'b00000000; //  939 :   0 - 0x0
      12'h3AC: dout <= 8'b00000000; //  940 :   0 - 0x0
      12'h3AD: dout <= 8'b00000000; //  941 :   0 - 0x0
      12'h3AE: dout <= 8'b00000000; //  942 :   0 - 0x0
      12'h3AF: dout <= 8'b00000000; //  943 :   0 - 0x0
      12'h3B0: dout <= 8'b00000000; //  944 :   0 - 0x0 -- Background 0x3b
      12'h3B1: dout <= 8'b00000010; //  945 :   2 - 0x2
      12'h3B2: dout <= 8'b00000100; //  946 :   4 - 0x4
      12'h3B3: dout <= 8'b00001000; //  947 :   8 - 0x8
      12'h3B4: dout <= 8'b00010000; //  948 :  16 - 0x10
      12'h3B5: dout <= 8'b00100000; //  949 :  32 - 0x20
      12'h3B6: dout <= 8'b00000000; //  950 :   0 - 0x0
      12'h3B7: dout <= 8'b00000000; //  951 :   0 - 0x0
      12'h3B8: dout <= 8'b00000000; //  952 :   0 - 0x0 -- plane 1
      12'h3B9: dout <= 8'b00000000; //  953 :   0 - 0x0
      12'h3BA: dout <= 8'b00000000; //  954 :   0 - 0x0
      12'h3BB: dout <= 8'b00000000; //  955 :   0 - 0x0
      12'h3BC: dout <= 8'b00000000; //  956 :   0 - 0x0
      12'h3BD: dout <= 8'b00000000; //  957 :   0 - 0x0
      12'h3BE: dout <= 8'b00000000; //  958 :   0 - 0x0
      12'h3BF: dout <= 8'b00000000; //  959 :   0 - 0x0
      12'h3C0: dout <= 8'b00000000; //  960 :   0 - 0x0 -- Background 0x3c
      12'h3C1: dout <= 8'b00000111; //  961 :   7 - 0x7
      12'h3C2: dout <= 8'b00011111; //  962 :  31 - 0x1f
      12'h3C3: dout <= 8'b00111111; //  963 :  63 - 0x3f
      12'h3C4: dout <= 8'b00111111; //  964 :  63 - 0x3f
      12'h3C5: dout <= 8'b00001111; //  965 :  15 - 0xf
      12'h3C6: dout <= 8'b00000011; //  966 :   3 - 0x3
      12'h3C7: dout <= 8'b00000000; //  967 :   0 - 0x0
      12'h3C8: dout <= 8'b00000000; //  968 :   0 - 0x0 -- plane 1
      12'h3C9: dout <= 8'b00000111; //  969 :   7 - 0x7
      12'h3CA: dout <= 8'b00011111; //  970 :  31 - 0x1f
      12'h3CB: dout <= 8'b00111111; //  971 :  63 - 0x3f
      12'h3CC: dout <= 8'b00111111; //  972 :  63 - 0x3f
      12'h3CD: dout <= 8'b00001111; //  973 :  15 - 0xf
      12'h3CE: dout <= 8'b00000011; //  974 :   3 - 0x3
      12'h3CF: dout <= 8'b00000000; //  975 :   0 - 0x0
      12'h3D0: dout <= 8'b00000000; //  976 :   0 - 0x0 -- Background 0x3d
      12'h3D1: dout <= 8'b11000000; //  977 : 192 - 0xc0
      12'h3D2: dout <= 8'b11110000; //  978 : 240 - 0xf0
      12'h3D3: dout <= 8'b11111000; //  979 : 248 - 0xf8
      12'h3D4: dout <= 8'b11111000; //  980 : 248 - 0xf8
      12'h3D5: dout <= 8'b11111100; //  981 : 252 - 0xfc
      12'h3D6: dout <= 8'b11111100; //  982 : 252 - 0xfc
      12'h3D7: dout <= 8'b11111100; //  983 : 252 - 0xfc
      12'h3D8: dout <= 8'b00000000; //  984 :   0 - 0x0 -- plane 1
      12'h3D9: dout <= 8'b11000000; //  985 : 192 - 0xc0
      12'h3DA: dout <= 8'b11110000; //  986 : 240 - 0xf0
      12'h3DB: dout <= 8'b11111000; //  987 : 248 - 0xf8
      12'h3DC: dout <= 8'b11111000; //  988 : 248 - 0xf8
      12'h3DD: dout <= 8'b11111100; //  989 : 252 - 0xfc
      12'h3DE: dout <= 8'b11111100; //  990 : 252 - 0xfc
      12'h3DF: dout <= 8'b11111100; //  991 : 252 - 0xfc
      12'h3E0: dout <= 8'b00000000; //  992 :   0 - 0x0 -- Background 0x3e
      12'h3E1: dout <= 8'b00000011; //  993 :   3 - 0x3
      12'h3E2: dout <= 8'b00001111; //  994 :  15 - 0xf
      12'h3E3: dout <= 8'b00111111; //  995 :  63 - 0x3f
      12'h3E4: dout <= 8'b00111111; //  996 :  63 - 0x3f
      12'h3E5: dout <= 8'b00011111; //  997 :  31 - 0x1f
      12'h3E6: dout <= 8'b00000111; //  998 :   7 - 0x7
      12'h3E7: dout <= 8'b00000000; //  999 :   0 - 0x0
      12'h3E8: dout <= 8'b00000000; // 1000 :   0 - 0x0 -- plane 1
      12'h3E9: dout <= 8'b00000011; // 1001 :   3 - 0x3
      12'h3EA: dout <= 8'b00001111; // 1002 :  15 - 0xf
      12'h3EB: dout <= 8'b00111111; // 1003 :  63 - 0x3f
      12'h3EC: dout <= 8'b00111111; // 1004 :  63 - 0x3f
      12'h3ED: dout <= 8'b00011111; // 1005 :  31 - 0x1f
      12'h3EE: dout <= 8'b00000111; // 1006 :   7 - 0x7
      12'h3EF: dout <= 8'b00000000; // 1007 :   0 - 0x0
      12'h3F0: dout <= 8'b11111100; // 1008 : 252 - 0xfc -- Background 0x3f
      12'h3F1: dout <= 8'b11111100; // 1009 : 252 - 0xfc
      12'h3F2: dout <= 8'b11111100; // 1010 : 252 - 0xfc
      12'h3F3: dout <= 8'b11111000; // 1011 : 248 - 0xf8
      12'h3F4: dout <= 8'b11111000; // 1012 : 248 - 0xf8
      12'h3F5: dout <= 8'b11110000; // 1013 : 240 - 0xf0
      12'h3F6: dout <= 8'b11000000; // 1014 : 192 - 0xc0
      12'h3F7: dout <= 8'b00000000; // 1015 :   0 - 0x0
      12'h3F8: dout <= 8'b11111100; // 1016 : 252 - 0xfc -- plane 1
      12'h3F9: dout <= 8'b11111100; // 1017 : 252 - 0xfc
      12'h3FA: dout <= 8'b11111100; // 1018 : 252 - 0xfc
      12'h3FB: dout <= 8'b11111000; // 1019 : 248 - 0xf8
      12'h3FC: dout <= 8'b11111000; // 1020 : 248 - 0xf8
      12'h3FD: dout <= 8'b11110000; // 1021 : 240 - 0xf0
      12'h3FE: dout <= 8'b11000000; // 1022 : 192 - 0xc0
      12'h3FF: dout <= 8'b00000000; // 1023 :   0 - 0x0
      12'h400: dout <= 8'b00000000; // 1024 :   0 - 0x0 -- Background 0x40
      12'h401: dout <= 8'b00000000; // 1025 :   0 - 0x0
      12'h402: dout <= 8'b00000000; // 1026 :   0 - 0x0
      12'h403: dout <= 8'b00000000; // 1027 :   0 - 0x0
      12'h404: dout <= 8'b00000000; // 1028 :   0 - 0x0
      12'h405: dout <= 8'b00000000; // 1029 :   0 - 0x0
      12'h406: dout <= 8'b00000000; // 1030 :   0 - 0x0
      12'h407: dout <= 8'b00000000; // 1031 :   0 - 0x0
      12'h408: dout <= 8'b00000000; // 1032 :   0 - 0x0 -- plane 1
      12'h409: dout <= 8'b00000000; // 1033 :   0 - 0x0
      12'h40A: dout <= 8'b00000000; // 1034 :   0 - 0x0
      12'h40B: dout <= 8'b00000000; // 1035 :   0 - 0x0
      12'h40C: dout <= 8'b00000000; // 1036 :   0 - 0x0
      12'h40D: dout <= 8'b00000000; // 1037 :   0 - 0x0
      12'h40E: dout <= 8'b00000000; // 1038 :   0 - 0x0
      12'h40F: dout <= 8'b00000000; // 1039 :   0 - 0x0
      12'h410: dout <= 8'b00011100; // 1040 :  28 - 0x1c -- Background 0x41
      12'h411: dout <= 8'b00110110; // 1041 :  54 - 0x36
      12'h412: dout <= 8'b01100011; // 1042 :  99 - 0x63
      12'h413: dout <= 8'b01100011; // 1043 :  99 - 0x63
      12'h414: dout <= 8'b01111111; // 1044 : 127 - 0x7f
      12'h415: dout <= 8'b01100011; // 1045 :  99 - 0x63
      12'h416: dout <= 8'b01100011; // 1046 :  99 - 0x63
      12'h417: dout <= 8'b00000000; // 1047 :   0 - 0x0
      12'h418: dout <= 8'b00000000; // 1048 :   0 - 0x0 -- plane 1
      12'h419: dout <= 8'b00000000; // 1049 :   0 - 0x0
      12'h41A: dout <= 8'b00000000; // 1050 :   0 - 0x0
      12'h41B: dout <= 8'b00000000; // 1051 :   0 - 0x0
      12'h41C: dout <= 8'b00000000; // 1052 :   0 - 0x0
      12'h41D: dout <= 8'b00000000; // 1053 :   0 - 0x0
      12'h41E: dout <= 8'b00000000; // 1054 :   0 - 0x0
      12'h41F: dout <= 8'b00000000; // 1055 :   0 - 0x0
      12'h420: dout <= 8'b01111110; // 1056 : 126 - 0x7e -- Background 0x42
      12'h421: dout <= 8'b01100011; // 1057 :  99 - 0x63
      12'h422: dout <= 8'b01100011; // 1058 :  99 - 0x63
      12'h423: dout <= 8'b01111110; // 1059 : 126 - 0x7e
      12'h424: dout <= 8'b01100011; // 1060 :  99 - 0x63
      12'h425: dout <= 8'b01100011; // 1061 :  99 - 0x63
      12'h426: dout <= 8'b01111110; // 1062 : 126 - 0x7e
      12'h427: dout <= 8'b00000000; // 1063 :   0 - 0x0
      12'h428: dout <= 8'b00000000; // 1064 :   0 - 0x0 -- plane 1
      12'h429: dout <= 8'b00000000; // 1065 :   0 - 0x0
      12'h42A: dout <= 8'b00000000; // 1066 :   0 - 0x0
      12'h42B: dout <= 8'b00000000; // 1067 :   0 - 0x0
      12'h42C: dout <= 8'b00000000; // 1068 :   0 - 0x0
      12'h42D: dout <= 8'b00000000; // 1069 :   0 - 0x0
      12'h42E: dout <= 8'b00000000; // 1070 :   0 - 0x0
      12'h42F: dout <= 8'b00000000; // 1071 :   0 - 0x0
      12'h430: dout <= 8'b00011110; // 1072 :  30 - 0x1e -- Background 0x43
      12'h431: dout <= 8'b00110011; // 1073 :  51 - 0x33
      12'h432: dout <= 8'b01100000; // 1074 :  96 - 0x60
      12'h433: dout <= 8'b01100000; // 1075 :  96 - 0x60
      12'h434: dout <= 8'b01100000; // 1076 :  96 - 0x60
      12'h435: dout <= 8'b00110011; // 1077 :  51 - 0x33
      12'h436: dout <= 8'b00011110; // 1078 :  30 - 0x1e
      12'h437: dout <= 8'b00000000; // 1079 :   0 - 0x0
      12'h438: dout <= 8'b00000000; // 1080 :   0 - 0x0 -- plane 1
      12'h439: dout <= 8'b00000000; // 1081 :   0 - 0x0
      12'h43A: dout <= 8'b00000000; // 1082 :   0 - 0x0
      12'h43B: dout <= 8'b00000000; // 1083 :   0 - 0x0
      12'h43C: dout <= 8'b00000000; // 1084 :   0 - 0x0
      12'h43D: dout <= 8'b00000000; // 1085 :   0 - 0x0
      12'h43E: dout <= 8'b00000000; // 1086 :   0 - 0x0
      12'h43F: dout <= 8'b00000000; // 1087 :   0 - 0x0
      12'h440: dout <= 8'b01111100; // 1088 : 124 - 0x7c -- Background 0x44
      12'h441: dout <= 8'b01100110; // 1089 : 102 - 0x66
      12'h442: dout <= 8'b01100011; // 1090 :  99 - 0x63
      12'h443: dout <= 8'b01100011; // 1091 :  99 - 0x63
      12'h444: dout <= 8'b01100011; // 1092 :  99 - 0x63
      12'h445: dout <= 8'b01100110; // 1093 : 102 - 0x66
      12'h446: dout <= 8'b01111100; // 1094 : 124 - 0x7c
      12'h447: dout <= 8'b00000000; // 1095 :   0 - 0x0
      12'h448: dout <= 8'b00000000; // 1096 :   0 - 0x0 -- plane 1
      12'h449: dout <= 8'b00000000; // 1097 :   0 - 0x0
      12'h44A: dout <= 8'b00000000; // 1098 :   0 - 0x0
      12'h44B: dout <= 8'b00000000; // 1099 :   0 - 0x0
      12'h44C: dout <= 8'b00000000; // 1100 :   0 - 0x0
      12'h44D: dout <= 8'b00000000; // 1101 :   0 - 0x0
      12'h44E: dout <= 8'b00000000; // 1102 :   0 - 0x0
      12'h44F: dout <= 8'b00000000; // 1103 :   0 - 0x0
      12'h450: dout <= 8'b01111111; // 1104 : 127 - 0x7f -- Background 0x45
      12'h451: dout <= 8'b01100000; // 1105 :  96 - 0x60
      12'h452: dout <= 8'b01100000; // 1106 :  96 - 0x60
      12'h453: dout <= 8'b01111110; // 1107 : 126 - 0x7e
      12'h454: dout <= 8'b01100000; // 1108 :  96 - 0x60
      12'h455: dout <= 8'b01100000; // 1109 :  96 - 0x60
      12'h456: dout <= 8'b01111111; // 1110 : 127 - 0x7f
      12'h457: dout <= 8'b00000000; // 1111 :   0 - 0x0
      12'h458: dout <= 8'b00000000; // 1112 :   0 - 0x0 -- plane 1
      12'h459: dout <= 8'b00000000; // 1113 :   0 - 0x0
      12'h45A: dout <= 8'b00000000; // 1114 :   0 - 0x0
      12'h45B: dout <= 8'b00000000; // 1115 :   0 - 0x0
      12'h45C: dout <= 8'b00000000; // 1116 :   0 - 0x0
      12'h45D: dout <= 8'b00000000; // 1117 :   0 - 0x0
      12'h45E: dout <= 8'b00000000; // 1118 :   0 - 0x0
      12'h45F: dout <= 8'b00000000; // 1119 :   0 - 0x0
      12'h460: dout <= 8'b01111111; // 1120 : 127 - 0x7f -- Background 0x46
      12'h461: dout <= 8'b01100000; // 1121 :  96 - 0x60
      12'h462: dout <= 8'b01100000; // 1122 :  96 - 0x60
      12'h463: dout <= 8'b01111110; // 1123 : 126 - 0x7e
      12'h464: dout <= 8'b01100000; // 1124 :  96 - 0x60
      12'h465: dout <= 8'b01100000; // 1125 :  96 - 0x60
      12'h466: dout <= 8'b01100000; // 1126 :  96 - 0x60
      12'h467: dout <= 8'b00000000; // 1127 :   0 - 0x0
      12'h468: dout <= 8'b00000000; // 1128 :   0 - 0x0 -- plane 1
      12'h469: dout <= 8'b00000000; // 1129 :   0 - 0x0
      12'h46A: dout <= 8'b00000000; // 1130 :   0 - 0x0
      12'h46B: dout <= 8'b00000000; // 1131 :   0 - 0x0
      12'h46C: dout <= 8'b00000000; // 1132 :   0 - 0x0
      12'h46D: dout <= 8'b00000000; // 1133 :   0 - 0x0
      12'h46E: dout <= 8'b00000000; // 1134 :   0 - 0x0
      12'h46F: dout <= 8'b00000000; // 1135 :   0 - 0x0
      12'h470: dout <= 8'b00011111; // 1136 :  31 - 0x1f -- Background 0x47
      12'h471: dout <= 8'b00110000; // 1137 :  48 - 0x30
      12'h472: dout <= 8'b01100000; // 1138 :  96 - 0x60
      12'h473: dout <= 8'b01100111; // 1139 : 103 - 0x67
      12'h474: dout <= 8'b01100011; // 1140 :  99 - 0x63
      12'h475: dout <= 8'b00110011; // 1141 :  51 - 0x33
      12'h476: dout <= 8'b00011111; // 1142 :  31 - 0x1f
      12'h477: dout <= 8'b00000000; // 1143 :   0 - 0x0
      12'h478: dout <= 8'b00000000; // 1144 :   0 - 0x0 -- plane 1
      12'h479: dout <= 8'b00000000; // 1145 :   0 - 0x0
      12'h47A: dout <= 8'b00000000; // 1146 :   0 - 0x0
      12'h47B: dout <= 8'b00000000; // 1147 :   0 - 0x0
      12'h47C: dout <= 8'b00000000; // 1148 :   0 - 0x0
      12'h47D: dout <= 8'b00000000; // 1149 :   0 - 0x0
      12'h47E: dout <= 8'b00000000; // 1150 :   0 - 0x0
      12'h47F: dout <= 8'b00000000; // 1151 :   0 - 0x0
      12'h480: dout <= 8'b01100011; // 1152 :  99 - 0x63 -- Background 0x48
      12'h481: dout <= 8'b01100011; // 1153 :  99 - 0x63
      12'h482: dout <= 8'b01100011; // 1154 :  99 - 0x63
      12'h483: dout <= 8'b01111111; // 1155 : 127 - 0x7f
      12'h484: dout <= 8'b01100011; // 1156 :  99 - 0x63
      12'h485: dout <= 8'b01100011; // 1157 :  99 - 0x63
      12'h486: dout <= 8'b01100011; // 1158 :  99 - 0x63
      12'h487: dout <= 8'b00000000; // 1159 :   0 - 0x0
      12'h488: dout <= 8'b00000000; // 1160 :   0 - 0x0 -- plane 1
      12'h489: dout <= 8'b00000000; // 1161 :   0 - 0x0
      12'h48A: dout <= 8'b00000000; // 1162 :   0 - 0x0
      12'h48B: dout <= 8'b00000000; // 1163 :   0 - 0x0
      12'h48C: dout <= 8'b00000000; // 1164 :   0 - 0x0
      12'h48D: dout <= 8'b00000000; // 1165 :   0 - 0x0
      12'h48E: dout <= 8'b00000000; // 1166 :   0 - 0x0
      12'h48F: dout <= 8'b00000000; // 1167 :   0 - 0x0
      12'h490: dout <= 8'b00111111; // 1168 :  63 - 0x3f -- Background 0x49
      12'h491: dout <= 8'b00001100; // 1169 :  12 - 0xc
      12'h492: dout <= 8'b00001100; // 1170 :  12 - 0xc
      12'h493: dout <= 8'b00001100; // 1171 :  12 - 0xc
      12'h494: dout <= 8'b00001100; // 1172 :  12 - 0xc
      12'h495: dout <= 8'b00001100; // 1173 :  12 - 0xc
      12'h496: dout <= 8'b00111111; // 1174 :  63 - 0x3f
      12'h497: dout <= 8'b00000000; // 1175 :   0 - 0x0
      12'h498: dout <= 8'b00000000; // 1176 :   0 - 0x0 -- plane 1
      12'h499: dout <= 8'b00000000; // 1177 :   0 - 0x0
      12'h49A: dout <= 8'b00000000; // 1178 :   0 - 0x0
      12'h49B: dout <= 8'b00000000; // 1179 :   0 - 0x0
      12'h49C: dout <= 8'b00000000; // 1180 :   0 - 0x0
      12'h49D: dout <= 8'b00000000; // 1181 :   0 - 0x0
      12'h49E: dout <= 8'b00000000; // 1182 :   0 - 0x0
      12'h49F: dout <= 8'b00000000; // 1183 :   0 - 0x0
      12'h4A0: dout <= 8'b00000011; // 1184 :   3 - 0x3 -- Background 0x4a
      12'h4A1: dout <= 8'b00000011; // 1185 :   3 - 0x3
      12'h4A2: dout <= 8'b00000011; // 1186 :   3 - 0x3
      12'h4A3: dout <= 8'b00000011; // 1187 :   3 - 0x3
      12'h4A4: dout <= 8'b00000011; // 1188 :   3 - 0x3
      12'h4A5: dout <= 8'b01100011; // 1189 :  99 - 0x63
      12'h4A6: dout <= 8'b00111110; // 1190 :  62 - 0x3e
      12'h4A7: dout <= 8'b00000000; // 1191 :   0 - 0x0
      12'h4A8: dout <= 8'b00000000; // 1192 :   0 - 0x0 -- plane 1
      12'h4A9: dout <= 8'b00000000; // 1193 :   0 - 0x0
      12'h4AA: dout <= 8'b00000000; // 1194 :   0 - 0x0
      12'h4AB: dout <= 8'b00000000; // 1195 :   0 - 0x0
      12'h4AC: dout <= 8'b00000000; // 1196 :   0 - 0x0
      12'h4AD: dout <= 8'b00000000; // 1197 :   0 - 0x0
      12'h4AE: dout <= 8'b00000000; // 1198 :   0 - 0x0
      12'h4AF: dout <= 8'b00000000; // 1199 :   0 - 0x0
      12'h4B0: dout <= 8'b01100011; // 1200 :  99 - 0x63 -- Background 0x4b
      12'h4B1: dout <= 8'b01100110; // 1201 : 102 - 0x66
      12'h4B2: dout <= 8'b01101100; // 1202 : 108 - 0x6c
      12'h4B3: dout <= 8'b01111000; // 1203 : 120 - 0x78
      12'h4B4: dout <= 8'b01111100; // 1204 : 124 - 0x7c
      12'h4B5: dout <= 8'b01100110; // 1205 : 102 - 0x66
      12'h4B6: dout <= 8'b01100011; // 1206 :  99 - 0x63
      12'h4B7: dout <= 8'b00000000; // 1207 :   0 - 0x0
      12'h4B8: dout <= 8'b00000000; // 1208 :   0 - 0x0 -- plane 1
      12'h4B9: dout <= 8'b00000000; // 1209 :   0 - 0x0
      12'h4BA: dout <= 8'b00000000; // 1210 :   0 - 0x0
      12'h4BB: dout <= 8'b00000000; // 1211 :   0 - 0x0
      12'h4BC: dout <= 8'b00000000; // 1212 :   0 - 0x0
      12'h4BD: dout <= 8'b00000000; // 1213 :   0 - 0x0
      12'h4BE: dout <= 8'b00000000; // 1214 :   0 - 0x0
      12'h4BF: dout <= 8'b00000000; // 1215 :   0 - 0x0
      12'h4C0: dout <= 8'b01100000; // 1216 :  96 - 0x60 -- Background 0x4c
      12'h4C1: dout <= 8'b01100000; // 1217 :  96 - 0x60
      12'h4C2: dout <= 8'b01100000; // 1218 :  96 - 0x60
      12'h4C3: dout <= 8'b01100000; // 1219 :  96 - 0x60
      12'h4C4: dout <= 8'b01100000; // 1220 :  96 - 0x60
      12'h4C5: dout <= 8'b01100000; // 1221 :  96 - 0x60
      12'h4C6: dout <= 8'b01111111; // 1222 : 127 - 0x7f
      12'h4C7: dout <= 8'b00000000; // 1223 :   0 - 0x0
      12'h4C8: dout <= 8'b00000000; // 1224 :   0 - 0x0 -- plane 1
      12'h4C9: dout <= 8'b00000000; // 1225 :   0 - 0x0
      12'h4CA: dout <= 8'b00000000; // 1226 :   0 - 0x0
      12'h4CB: dout <= 8'b00000000; // 1227 :   0 - 0x0
      12'h4CC: dout <= 8'b00000000; // 1228 :   0 - 0x0
      12'h4CD: dout <= 8'b00000000; // 1229 :   0 - 0x0
      12'h4CE: dout <= 8'b00000000; // 1230 :   0 - 0x0
      12'h4CF: dout <= 8'b00000000; // 1231 :   0 - 0x0
      12'h4D0: dout <= 8'b01100011; // 1232 :  99 - 0x63 -- Background 0x4d
      12'h4D1: dout <= 8'b01110111; // 1233 : 119 - 0x77
      12'h4D2: dout <= 8'b01111111; // 1234 : 127 - 0x7f
      12'h4D3: dout <= 8'b01111111; // 1235 : 127 - 0x7f
      12'h4D4: dout <= 8'b01101011; // 1236 : 107 - 0x6b
      12'h4D5: dout <= 8'b01100011; // 1237 :  99 - 0x63
      12'h4D6: dout <= 8'b01100011; // 1238 :  99 - 0x63
      12'h4D7: dout <= 8'b00000000; // 1239 :   0 - 0x0
      12'h4D8: dout <= 8'b00000000; // 1240 :   0 - 0x0 -- plane 1
      12'h4D9: dout <= 8'b00000000; // 1241 :   0 - 0x0
      12'h4DA: dout <= 8'b00000000; // 1242 :   0 - 0x0
      12'h4DB: dout <= 8'b00000000; // 1243 :   0 - 0x0
      12'h4DC: dout <= 8'b00000000; // 1244 :   0 - 0x0
      12'h4DD: dout <= 8'b00000000; // 1245 :   0 - 0x0
      12'h4DE: dout <= 8'b00000000; // 1246 :   0 - 0x0
      12'h4DF: dout <= 8'b00000000; // 1247 :   0 - 0x0
      12'h4E0: dout <= 8'b01100011; // 1248 :  99 - 0x63 -- Background 0x4e
      12'h4E1: dout <= 8'b01110011; // 1249 : 115 - 0x73
      12'h4E2: dout <= 8'b01111011; // 1250 : 123 - 0x7b
      12'h4E3: dout <= 8'b01111111; // 1251 : 127 - 0x7f
      12'h4E4: dout <= 8'b01101111; // 1252 : 111 - 0x6f
      12'h4E5: dout <= 8'b01100111; // 1253 : 103 - 0x67
      12'h4E6: dout <= 8'b01100011; // 1254 :  99 - 0x63
      12'h4E7: dout <= 8'b00000000; // 1255 :   0 - 0x0
      12'h4E8: dout <= 8'b00000000; // 1256 :   0 - 0x0 -- plane 1
      12'h4E9: dout <= 8'b00000000; // 1257 :   0 - 0x0
      12'h4EA: dout <= 8'b00000000; // 1258 :   0 - 0x0
      12'h4EB: dout <= 8'b00000000; // 1259 :   0 - 0x0
      12'h4EC: dout <= 8'b00000000; // 1260 :   0 - 0x0
      12'h4ED: dout <= 8'b00000000; // 1261 :   0 - 0x0
      12'h4EE: dout <= 8'b00000000; // 1262 :   0 - 0x0
      12'h4EF: dout <= 8'b00000000; // 1263 :   0 - 0x0
      12'h4F0: dout <= 8'b00111110; // 1264 :  62 - 0x3e -- Background 0x4f
      12'h4F1: dout <= 8'b01100011; // 1265 :  99 - 0x63
      12'h4F2: dout <= 8'b01100011; // 1266 :  99 - 0x63
      12'h4F3: dout <= 8'b01100011; // 1267 :  99 - 0x63
      12'h4F4: dout <= 8'b01100011; // 1268 :  99 - 0x63
      12'h4F5: dout <= 8'b01100011; // 1269 :  99 - 0x63
      12'h4F6: dout <= 8'b00111110; // 1270 :  62 - 0x3e
      12'h4F7: dout <= 8'b00000000; // 1271 :   0 - 0x0
      12'h4F8: dout <= 8'b00000000; // 1272 :   0 - 0x0 -- plane 1
      12'h4F9: dout <= 8'b00000000; // 1273 :   0 - 0x0
      12'h4FA: dout <= 8'b00000000; // 1274 :   0 - 0x0
      12'h4FB: dout <= 8'b00000000; // 1275 :   0 - 0x0
      12'h4FC: dout <= 8'b00000000; // 1276 :   0 - 0x0
      12'h4FD: dout <= 8'b00000000; // 1277 :   0 - 0x0
      12'h4FE: dout <= 8'b00000000; // 1278 :   0 - 0x0
      12'h4FF: dout <= 8'b00000000; // 1279 :   0 - 0x0
      12'h500: dout <= 8'b01111110; // 1280 : 126 - 0x7e -- Background 0x50
      12'h501: dout <= 8'b01100011; // 1281 :  99 - 0x63
      12'h502: dout <= 8'b01100011; // 1282 :  99 - 0x63
      12'h503: dout <= 8'b01100011; // 1283 :  99 - 0x63
      12'h504: dout <= 8'b01111110; // 1284 : 126 - 0x7e
      12'h505: dout <= 8'b01100000; // 1285 :  96 - 0x60
      12'h506: dout <= 8'b01100000; // 1286 :  96 - 0x60
      12'h507: dout <= 8'b00000000; // 1287 :   0 - 0x0
      12'h508: dout <= 8'b00000000; // 1288 :   0 - 0x0 -- plane 1
      12'h509: dout <= 8'b00000000; // 1289 :   0 - 0x0
      12'h50A: dout <= 8'b00000000; // 1290 :   0 - 0x0
      12'h50B: dout <= 8'b00000000; // 1291 :   0 - 0x0
      12'h50C: dout <= 8'b00000000; // 1292 :   0 - 0x0
      12'h50D: dout <= 8'b00000000; // 1293 :   0 - 0x0
      12'h50E: dout <= 8'b00000000; // 1294 :   0 - 0x0
      12'h50F: dout <= 8'b00000000; // 1295 :   0 - 0x0
      12'h510: dout <= 8'b00111110; // 1296 :  62 - 0x3e -- Background 0x51
      12'h511: dout <= 8'b01100011; // 1297 :  99 - 0x63
      12'h512: dout <= 8'b01100011; // 1298 :  99 - 0x63
      12'h513: dout <= 8'b01100011; // 1299 :  99 - 0x63
      12'h514: dout <= 8'b01101111; // 1300 : 111 - 0x6f
      12'h515: dout <= 8'b01100110; // 1301 : 102 - 0x66
      12'h516: dout <= 8'b00111101; // 1302 :  61 - 0x3d
      12'h517: dout <= 8'b00000000; // 1303 :   0 - 0x0
      12'h518: dout <= 8'b00000000; // 1304 :   0 - 0x0 -- plane 1
      12'h519: dout <= 8'b00000000; // 1305 :   0 - 0x0
      12'h51A: dout <= 8'b00000000; // 1306 :   0 - 0x0
      12'h51B: dout <= 8'b00000000; // 1307 :   0 - 0x0
      12'h51C: dout <= 8'b00000000; // 1308 :   0 - 0x0
      12'h51D: dout <= 8'b00000000; // 1309 :   0 - 0x0
      12'h51E: dout <= 8'b00000000; // 1310 :   0 - 0x0
      12'h51F: dout <= 8'b00000000; // 1311 :   0 - 0x0
      12'h520: dout <= 8'b01111110; // 1312 : 126 - 0x7e -- Background 0x52
      12'h521: dout <= 8'b01100011; // 1313 :  99 - 0x63
      12'h522: dout <= 8'b01100011; // 1314 :  99 - 0x63
      12'h523: dout <= 8'b01100111; // 1315 : 103 - 0x67
      12'h524: dout <= 8'b01111100; // 1316 : 124 - 0x7c
      12'h525: dout <= 8'b01101110; // 1317 : 110 - 0x6e
      12'h526: dout <= 8'b01100111; // 1318 : 103 - 0x67
      12'h527: dout <= 8'b00000000; // 1319 :   0 - 0x0
      12'h528: dout <= 8'b00000000; // 1320 :   0 - 0x0 -- plane 1
      12'h529: dout <= 8'b00000000; // 1321 :   0 - 0x0
      12'h52A: dout <= 8'b00000000; // 1322 :   0 - 0x0
      12'h52B: dout <= 8'b00000000; // 1323 :   0 - 0x0
      12'h52C: dout <= 8'b00000000; // 1324 :   0 - 0x0
      12'h52D: dout <= 8'b00000000; // 1325 :   0 - 0x0
      12'h52E: dout <= 8'b00000000; // 1326 :   0 - 0x0
      12'h52F: dout <= 8'b00000000; // 1327 :   0 - 0x0
      12'h530: dout <= 8'b00111100; // 1328 :  60 - 0x3c -- Background 0x53
      12'h531: dout <= 8'b01100110; // 1329 : 102 - 0x66
      12'h532: dout <= 8'b01100000; // 1330 :  96 - 0x60
      12'h533: dout <= 8'b00111110; // 1331 :  62 - 0x3e
      12'h534: dout <= 8'b00000011; // 1332 :   3 - 0x3
      12'h535: dout <= 8'b01100011; // 1333 :  99 - 0x63
      12'h536: dout <= 8'b00111110; // 1334 :  62 - 0x3e
      12'h537: dout <= 8'b00000000; // 1335 :   0 - 0x0
      12'h538: dout <= 8'b00000000; // 1336 :   0 - 0x0 -- plane 1
      12'h539: dout <= 8'b00000000; // 1337 :   0 - 0x0
      12'h53A: dout <= 8'b00000000; // 1338 :   0 - 0x0
      12'h53B: dout <= 8'b00000000; // 1339 :   0 - 0x0
      12'h53C: dout <= 8'b00000000; // 1340 :   0 - 0x0
      12'h53D: dout <= 8'b00000000; // 1341 :   0 - 0x0
      12'h53E: dout <= 8'b00000000; // 1342 :   0 - 0x0
      12'h53F: dout <= 8'b00000000; // 1343 :   0 - 0x0
      12'h540: dout <= 8'b00111111; // 1344 :  63 - 0x3f -- Background 0x54
      12'h541: dout <= 8'b00001100; // 1345 :  12 - 0xc
      12'h542: dout <= 8'b00001100; // 1346 :  12 - 0xc
      12'h543: dout <= 8'b00001100; // 1347 :  12 - 0xc
      12'h544: dout <= 8'b00001100; // 1348 :  12 - 0xc
      12'h545: dout <= 8'b00001100; // 1349 :  12 - 0xc
      12'h546: dout <= 8'b00001100; // 1350 :  12 - 0xc
      12'h547: dout <= 8'b00000000; // 1351 :   0 - 0x0
      12'h548: dout <= 8'b00000000; // 1352 :   0 - 0x0 -- plane 1
      12'h549: dout <= 8'b00000000; // 1353 :   0 - 0x0
      12'h54A: dout <= 8'b00000000; // 1354 :   0 - 0x0
      12'h54B: dout <= 8'b00000000; // 1355 :   0 - 0x0
      12'h54C: dout <= 8'b00000000; // 1356 :   0 - 0x0
      12'h54D: dout <= 8'b00000000; // 1357 :   0 - 0x0
      12'h54E: dout <= 8'b00000000; // 1358 :   0 - 0x0
      12'h54F: dout <= 8'b00000000; // 1359 :   0 - 0x0
      12'h550: dout <= 8'b01100011; // 1360 :  99 - 0x63 -- Background 0x55
      12'h551: dout <= 8'b01100011; // 1361 :  99 - 0x63
      12'h552: dout <= 8'b01100011; // 1362 :  99 - 0x63
      12'h553: dout <= 8'b01100011; // 1363 :  99 - 0x63
      12'h554: dout <= 8'b01100011; // 1364 :  99 - 0x63
      12'h555: dout <= 8'b01100011; // 1365 :  99 - 0x63
      12'h556: dout <= 8'b00111110; // 1366 :  62 - 0x3e
      12'h557: dout <= 8'b00000000; // 1367 :   0 - 0x0
      12'h558: dout <= 8'b00000000; // 1368 :   0 - 0x0 -- plane 1
      12'h559: dout <= 8'b00000000; // 1369 :   0 - 0x0
      12'h55A: dout <= 8'b00000000; // 1370 :   0 - 0x0
      12'h55B: dout <= 8'b00000000; // 1371 :   0 - 0x0
      12'h55C: dout <= 8'b00000000; // 1372 :   0 - 0x0
      12'h55D: dout <= 8'b00000000; // 1373 :   0 - 0x0
      12'h55E: dout <= 8'b00000000; // 1374 :   0 - 0x0
      12'h55F: dout <= 8'b00000000; // 1375 :   0 - 0x0
      12'h560: dout <= 8'b01100011; // 1376 :  99 - 0x63 -- Background 0x56
      12'h561: dout <= 8'b01100011; // 1377 :  99 - 0x63
      12'h562: dout <= 8'b01100011; // 1378 :  99 - 0x63
      12'h563: dout <= 8'b01110111; // 1379 : 119 - 0x77
      12'h564: dout <= 8'b00111110; // 1380 :  62 - 0x3e
      12'h565: dout <= 8'b00011100; // 1381 :  28 - 0x1c
      12'h566: dout <= 8'b00001000; // 1382 :   8 - 0x8
      12'h567: dout <= 8'b00000000; // 1383 :   0 - 0x0
      12'h568: dout <= 8'b00000000; // 1384 :   0 - 0x0 -- plane 1
      12'h569: dout <= 8'b00000000; // 1385 :   0 - 0x0
      12'h56A: dout <= 8'b00000000; // 1386 :   0 - 0x0
      12'h56B: dout <= 8'b00000000; // 1387 :   0 - 0x0
      12'h56C: dout <= 8'b00000000; // 1388 :   0 - 0x0
      12'h56D: dout <= 8'b00000000; // 1389 :   0 - 0x0
      12'h56E: dout <= 8'b00000000; // 1390 :   0 - 0x0
      12'h56F: dout <= 8'b00000000; // 1391 :   0 - 0x0
      12'h570: dout <= 8'b01100011; // 1392 :  99 - 0x63 -- Background 0x57
      12'h571: dout <= 8'b01100011; // 1393 :  99 - 0x63
      12'h572: dout <= 8'b01101011; // 1394 : 107 - 0x6b
      12'h573: dout <= 8'b01111111; // 1395 : 127 - 0x7f
      12'h574: dout <= 8'b01111111; // 1396 : 127 - 0x7f
      12'h575: dout <= 8'b01110111; // 1397 : 119 - 0x77
      12'h576: dout <= 8'b01100011; // 1398 :  99 - 0x63
      12'h577: dout <= 8'b00000000; // 1399 :   0 - 0x0
      12'h578: dout <= 8'b00000000; // 1400 :   0 - 0x0 -- plane 1
      12'h579: dout <= 8'b00000000; // 1401 :   0 - 0x0
      12'h57A: dout <= 8'b00000000; // 1402 :   0 - 0x0
      12'h57B: dout <= 8'b00000000; // 1403 :   0 - 0x0
      12'h57C: dout <= 8'b00000000; // 1404 :   0 - 0x0
      12'h57D: dout <= 8'b00000000; // 1405 :   0 - 0x0
      12'h57E: dout <= 8'b00000000; // 1406 :   0 - 0x0
      12'h57F: dout <= 8'b00000000; // 1407 :   0 - 0x0
      12'h580: dout <= 8'b01100011; // 1408 :  99 - 0x63 -- Background 0x58
      12'h581: dout <= 8'b01110111; // 1409 : 119 - 0x77
      12'h582: dout <= 8'b00111110; // 1410 :  62 - 0x3e
      12'h583: dout <= 8'b00011100; // 1411 :  28 - 0x1c
      12'h584: dout <= 8'b00111110; // 1412 :  62 - 0x3e
      12'h585: dout <= 8'b01110111; // 1413 : 119 - 0x77
      12'h586: dout <= 8'b01100011; // 1414 :  99 - 0x63
      12'h587: dout <= 8'b00000000; // 1415 :   0 - 0x0
      12'h588: dout <= 8'b00000000; // 1416 :   0 - 0x0 -- plane 1
      12'h589: dout <= 8'b00000000; // 1417 :   0 - 0x0
      12'h58A: dout <= 8'b00000000; // 1418 :   0 - 0x0
      12'h58B: dout <= 8'b00000000; // 1419 :   0 - 0x0
      12'h58C: dout <= 8'b00000000; // 1420 :   0 - 0x0
      12'h58D: dout <= 8'b00000000; // 1421 :   0 - 0x0
      12'h58E: dout <= 8'b00000000; // 1422 :   0 - 0x0
      12'h58F: dout <= 8'b00000000; // 1423 :   0 - 0x0
      12'h590: dout <= 8'b00110011; // 1424 :  51 - 0x33 -- Background 0x59
      12'h591: dout <= 8'b00110011; // 1425 :  51 - 0x33
      12'h592: dout <= 8'b00110011; // 1426 :  51 - 0x33
      12'h593: dout <= 8'b00011110; // 1427 :  30 - 0x1e
      12'h594: dout <= 8'b00001100; // 1428 :  12 - 0xc
      12'h595: dout <= 8'b00001100; // 1429 :  12 - 0xc
      12'h596: dout <= 8'b00001100; // 1430 :  12 - 0xc
      12'h597: dout <= 8'b00000000; // 1431 :   0 - 0x0
      12'h598: dout <= 8'b00000000; // 1432 :   0 - 0x0 -- plane 1
      12'h599: dout <= 8'b00000000; // 1433 :   0 - 0x0
      12'h59A: dout <= 8'b00000000; // 1434 :   0 - 0x0
      12'h59B: dout <= 8'b00000000; // 1435 :   0 - 0x0
      12'h59C: dout <= 8'b00000000; // 1436 :   0 - 0x0
      12'h59D: dout <= 8'b00000000; // 1437 :   0 - 0x0
      12'h59E: dout <= 8'b00000000; // 1438 :   0 - 0x0
      12'h59F: dout <= 8'b00000000; // 1439 :   0 - 0x0
      12'h5A0: dout <= 8'b01111111; // 1440 : 127 - 0x7f -- Background 0x5a
      12'h5A1: dout <= 8'b00000111; // 1441 :   7 - 0x7
      12'h5A2: dout <= 8'b00001110; // 1442 :  14 - 0xe
      12'h5A3: dout <= 8'b00011100; // 1443 :  28 - 0x1c
      12'h5A4: dout <= 8'b00111000; // 1444 :  56 - 0x38
      12'h5A5: dout <= 8'b01110000; // 1445 : 112 - 0x70
      12'h5A6: dout <= 8'b01111111; // 1446 : 127 - 0x7f
      12'h5A7: dout <= 8'b00000000; // 1447 :   0 - 0x0
      12'h5A8: dout <= 8'b00000000; // 1448 :   0 - 0x0 -- plane 1
      12'h5A9: dout <= 8'b00000000; // 1449 :   0 - 0x0
      12'h5AA: dout <= 8'b00000000; // 1450 :   0 - 0x0
      12'h5AB: dout <= 8'b00000000; // 1451 :   0 - 0x0
      12'h5AC: dout <= 8'b00000000; // 1452 :   0 - 0x0
      12'h5AD: dout <= 8'b00000000; // 1453 :   0 - 0x0
      12'h5AE: dout <= 8'b00000000; // 1454 :   0 - 0x0
      12'h5AF: dout <= 8'b00000000; // 1455 :   0 - 0x0
      12'h5B0: dout <= 8'b00000000; // 1456 :   0 - 0x0 -- Background 0x5b
      12'h5B1: dout <= 8'b00000000; // 1457 :   0 - 0x0
      12'h5B2: dout <= 8'b00000000; // 1458 :   0 - 0x0
      12'h5B3: dout <= 8'b00000000; // 1459 :   0 - 0x0
      12'h5B4: dout <= 8'b00000000; // 1460 :   0 - 0x0
      12'h5B5: dout <= 8'b00110000; // 1461 :  48 - 0x30
      12'h5B6: dout <= 8'b00110000; // 1462 :  48 - 0x30
      12'h5B7: dout <= 8'b00000000; // 1463 :   0 - 0x0
      12'h5B8: dout <= 8'b00000000; // 1464 :   0 - 0x0 -- plane 1
      12'h5B9: dout <= 8'b00000000; // 1465 :   0 - 0x0
      12'h5BA: dout <= 8'b00000000; // 1466 :   0 - 0x0
      12'h5BB: dout <= 8'b00000000; // 1467 :   0 - 0x0
      12'h5BC: dout <= 8'b00000000; // 1468 :   0 - 0x0
      12'h5BD: dout <= 8'b00000000; // 1469 :   0 - 0x0
      12'h5BE: dout <= 8'b00000000; // 1470 :   0 - 0x0
      12'h5BF: dout <= 8'b00000000; // 1471 :   0 - 0x0
      12'h5C0: dout <= 8'b11000000; // 1472 : 192 - 0xc0 -- Background 0x5c
      12'h5C1: dout <= 8'b11110000; // 1473 : 240 - 0xf0
      12'h5C2: dout <= 8'b11111100; // 1474 : 252 - 0xfc
      12'h5C3: dout <= 8'b11111111; // 1475 : 255 - 0xff
      12'h5C4: dout <= 8'b11111100; // 1476 : 252 - 0xfc
      12'h5C5: dout <= 8'b11110000; // 1477 : 240 - 0xf0
      12'h5C6: dout <= 8'b11000000; // 1478 : 192 - 0xc0
      12'h5C7: dout <= 8'b00000000; // 1479 :   0 - 0x0
      12'h5C8: dout <= 8'b00000000; // 1480 :   0 - 0x0 -- plane 1
      12'h5C9: dout <= 8'b00000000; // 1481 :   0 - 0x0
      12'h5CA: dout <= 8'b00000000; // 1482 :   0 - 0x0
      12'h5CB: dout <= 8'b00000000; // 1483 :   0 - 0x0
      12'h5CC: dout <= 8'b00000000; // 1484 :   0 - 0x0
      12'h5CD: dout <= 8'b00000000; // 1485 :   0 - 0x0
      12'h5CE: dout <= 8'b00000000; // 1486 :   0 - 0x0
      12'h5CF: dout <= 8'b00000000; // 1487 :   0 - 0x0
      12'h5D0: dout <= 8'b00111100; // 1488 :  60 - 0x3c -- Background 0x5d
      12'h5D1: dout <= 8'b01000010; // 1489 :  66 - 0x42
      12'h5D2: dout <= 8'b10011001; // 1490 : 153 - 0x99
      12'h5D3: dout <= 8'b10100001; // 1491 : 161 - 0xa1
      12'h5D4: dout <= 8'b10100001; // 1492 : 161 - 0xa1
      12'h5D5: dout <= 8'b10011001; // 1493 : 153 - 0x99
      12'h5D6: dout <= 8'b01000010; // 1494 :  66 - 0x42
      12'h5D7: dout <= 8'b00111100; // 1495 :  60 - 0x3c
      12'h5D8: dout <= 8'b00000000; // 1496 :   0 - 0x0 -- plane 1
      12'h5D9: dout <= 8'b00000000; // 1497 :   0 - 0x0
      12'h5DA: dout <= 8'b00000000; // 1498 :   0 - 0x0
      12'h5DB: dout <= 8'b00000000; // 1499 :   0 - 0x0
      12'h5DC: dout <= 8'b00000000; // 1500 :   0 - 0x0
      12'h5DD: dout <= 8'b00000000; // 1501 :   0 - 0x0
      12'h5DE: dout <= 8'b00000000; // 1502 :   0 - 0x0
      12'h5DF: dout <= 8'b00000000; // 1503 :   0 - 0x0
      12'h5E0: dout <= 8'b00000000; // 1504 :   0 - 0x0 -- Background 0x5e
      12'h5E1: dout <= 8'b00000000; // 1505 :   0 - 0x0
      12'h5E2: dout <= 8'b00010000; // 1506 :  16 - 0x10
      12'h5E3: dout <= 8'b00010000; // 1507 :  16 - 0x10
      12'h5E4: dout <= 8'b00010000; // 1508 :  16 - 0x10
      12'h5E5: dout <= 8'b00010000; // 1509 :  16 - 0x10
      12'h5E6: dout <= 8'b00000000; // 1510 :   0 - 0x0
      12'h5E7: dout <= 8'b00000000; // 1511 :   0 - 0x0
      12'h5E8: dout <= 8'b00000000; // 1512 :   0 - 0x0 -- plane 1
      12'h5E9: dout <= 8'b00000000; // 1513 :   0 - 0x0
      12'h5EA: dout <= 8'b00010000; // 1514 :  16 - 0x10
      12'h5EB: dout <= 8'b00010000; // 1515 :  16 - 0x10
      12'h5EC: dout <= 8'b00010000; // 1516 :  16 - 0x10
      12'h5ED: dout <= 8'b00010000; // 1517 :  16 - 0x10
      12'h5EE: dout <= 8'b00000000; // 1518 :   0 - 0x0
      12'h5EF: dout <= 8'b00000000; // 1519 :   0 - 0x0
      12'h5F0: dout <= 8'b00110110; // 1520 :  54 - 0x36 -- Background 0x5f
      12'h5F1: dout <= 8'b00110110; // 1521 :  54 - 0x36
      12'h5F2: dout <= 8'b00010010; // 1522 :  18 - 0x12
      12'h5F3: dout <= 8'b00000000; // 1523 :   0 - 0x0
      12'h5F4: dout <= 8'b00000000; // 1524 :   0 - 0x0
      12'h5F5: dout <= 8'b00000000; // 1525 :   0 - 0x0
      12'h5F6: dout <= 8'b00000000; // 1526 :   0 - 0x0
      12'h5F7: dout <= 8'b00000000; // 1527 :   0 - 0x0
      12'h5F8: dout <= 8'b00000000; // 1528 :   0 - 0x0 -- plane 1
      12'h5F9: dout <= 8'b00000000; // 1529 :   0 - 0x0
      12'h5FA: dout <= 8'b00000000; // 1530 :   0 - 0x0
      12'h5FB: dout <= 8'b00000000; // 1531 :   0 - 0x0
      12'h5FC: dout <= 8'b00000000; // 1532 :   0 - 0x0
      12'h5FD: dout <= 8'b00000000; // 1533 :   0 - 0x0
      12'h5FE: dout <= 8'b00000000; // 1534 :   0 - 0x0
      12'h5FF: dout <= 8'b00000000; // 1535 :   0 - 0x0
      12'h600: dout <= 8'b00000000; // 1536 :   0 - 0x0 -- Background 0x60
      12'h601: dout <= 8'b00000000; // 1537 :   0 - 0x0
      12'h602: dout <= 8'b00000000; // 1538 :   0 - 0x0
      12'h603: dout <= 8'b00000000; // 1539 :   0 - 0x0
      12'h604: dout <= 8'b00000000; // 1540 :   0 - 0x0
      12'h605: dout <= 8'b00000001; // 1541 :   1 - 0x1
      12'h606: dout <= 8'b00011110; // 1542 :  30 - 0x1e
      12'h607: dout <= 8'b00111011; // 1543 :  59 - 0x3b
      12'h608: dout <= 8'b00000000; // 1544 :   0 - 0x0 -- plane 1
      12'h609: dout <= 8'b00000000; // 1545 :   0 - 0x0
      12'h60A: dout <= 8'b00000000; // 1546 :   0 - 0x0
      12'h60B: dout <= 8'b00000000; // 1547 :   0 - 0x0
      12'h60C: dout <= 8'b00000000; // 1548 :   0 - 0x0
      12'h60D: dout <= 8'b00000000; // 1549 :   0 - 0x0
      12'h60E: dout <= 8'b00000000; // 1550 :   0 - 0x0
      12'h60F: dout <= 8'b00000000; // 1551 :   0 - 0x0
      12'h610: dout <= 8'b00000000; // 1552 :   0 - 0x0 -- Background 0x61
      12'h611: dout <= 8'b00000000; // 1553 :   0 - 0x0
      12'h612: dout <= 8'b00001100; // 1554 :  12 - 0xc
      12'h613: dout <= 8'b00111100; // 1555 :  60 - 0x3c
      12'h614: dout <= 8'b11010000; // 1556 : 208 - 0xd0
      12'h615: dout <= 8'b00010000; // 1557 :  16 - 0x10
      12'h616: dout <= 8'b00100000; // 1558 :  32 - 0x20
      12'h617: dout <= 8'b01000000; // 1559 :  64 - 0x40
      12'h618: dout <= 8'b00000000; // 1560 :   0 - 0x0 -- plane 1
      12'h619: dout <= 8'b00000000; // 1561 :   0 - 0x0
      12'h61A: dout <= 8'b00000000; // 1562 :   0 - 0x0
      12'h61B: dout <= 8'b00000000; // 1563 :   0 - 0x0
      12'h61C: dout <= 8'b00000000; // 1564 :   0 - 0x0
      12'h61D: dout <= 8'b00000000; // 1565 :   0 - 0x0
      12'h61E: dout <= 8'b00000000; // 1566 :   0 - 0x0
      12'h61F: dout <= 8'b00000000; // 1567 :   0 - 0x0
      12'h620: dout <= 8'b00111110; // 1568 :  62 - 0x3e -- Background 0x62
      12'h621: dout <= 8'b00101101; // 1569 :  45 - 0x2d
      12'h622: dout <= 8'b00110101; // 1570 :  53 - 0x35
      12'h623: dout <= 8'b00011101; // 1571 :  29 - 0x1d
      12'h624: dout <= 8'b00000001; // 1572 :   1 - 0x1
      12'h625: dout <= 8'b00000000; // 1573 :   0 - 0x0
      12'h626: dout <= 8'b00000000; // 1574 :   0 - 0x0
      12'h627: dout <= 8'b00000000; // 1575 :   0 - 0x0
      12'h628: dout <= 8'b00000000; // 1576 :   0 - 0x0 -- plane 1
      12'h629: dout <= 8'b00000000; // 1577 :   0 - 0x0
      12'h62A: dout <= 8'b00000000; // 1578 :   0 - 0x0
      12'h62B: dout <= 8'b00000000; // 1579 :   0 - 0x0
      12'h62C: dout <= 8'b00000000; // 1580 :   0 - 0x0
      12'h62D: dout <= 8'b00000000; // 1581 :   0 - 0x0
      12'h62E: dout <= 8'b00000000; // 1582 :   0 - 0x0
      12'h62F: dout <= 8'b00000000; // 1583 :   0 - 0x0
      12'h630: dout <= 8'b10110000; // 1584 : 176 - 0xb0 -- Background 0x63
      12'h631: dout <= 8'b10111000; // 1585 : 184 - 0xb8
      12'h632: dout <= 8'b11111000; // 1586 : 248 - 0xf8
      12'h633: dout <= 8'b01111000; // 1587 : 120 - 0x78
      12'h634: dout <= 8'b10011000; // 1588 : 152 - 0x98
      12'h635: dout <= 8'b11110000; // 1589 : 240 - 0xf0
      12'h636: dout <= 8'b00000000; // 1590 :   0 - 0x0
      12'h637: dout <= 8'b00000000; // 1591 :   0 - 0x0
      12'h638: dout <= 8'b00000000; // 1592 :   0 - 0x0 -- plane 1
      12'h639: dout <= 8'b00000000; // 1593 :   0 - 0x0
      12'h63A: dout <= 8'b00000000; // 1594 :   0 - 0x0
      12'h63B: dout <= 8'b00000000; // 1595 :   0 - 0x0
      12'h63C: dout <= 8'b00000000; // 1596 :   0 - 0x0
      12'h63D: dout <= 8'b00000000; // 1597 :   0 - 0x0
      12'h63E: dout <= 8'b00000000; // 1598 :   0 - 0x0
      12'h63F: dout <= 8'b00000000; // 1599 :   0 - 0x0
      12'h640: dout <= 8'b00000000; // 1600 :   0 - 0x0 -- Background 0x64
      12'h641: dout <= 8'b00000000; // 1601 :   0 - 0x0
      12'h642: dout <= 8'b00000111; // 1602 :   7 - 0x7
      12'h643: dout <= 8'b00000011; // 1603 :   3 - 0x3
      12'h644: dout <= 8'b00001101; // 1604 :  13 - 0xd
      12'h645: dout <= 8'b00011110; // 1605 :  30 - 0x1e
      12'h646: dout <= 8'b00010111; // 1606 :  23 - 0x17
      12'h647: dout <= 8'b00011101; // 1607 :  29 - 0x1d
      12'h648: dout <= 8'b00000000; // 1608 :   0 - 0x0 -- plane 1
      12'h649: dout <= 8'b00000000; // 1609 :   0 - 0x0
      12'h64A: dout <= 8'b00000000; // 1610 :   0 - 0x0
      12'h64B: dout <= 8'b00000000; // 1611 :   0 - 0x0
      12'h64C: dout <= 8'b00000000; // 1612 :   0 - 0x0
      12'h64D: dout <= 8'b00000000; // 1613 :   0 - 0x0
      12'h64E: dout <= 8'b00000000; // 1614 :   0 - 0x0
      12'h64F: dout <= 8'b00000000; // 1615 :   0 - 0x0
      12'h650: dout <= 8'b00000000; // 1616 :   0 - 0x0 -- Background 0x65
      12'h651: dout <= 8'b10000000; // 1617 : 128 - 0x80
      12'h652: dout <= 8'b01110000; // 1618 : 112 - 0x70
      12'h653: dout <= 8'b11100000; // 1619 : 224 - 0xe0
      12'h654: dout <= 8'b11011000; // 1620 : 216 - 0xd8
      12'h655: dout <= 8'b10111100; // 1621 : 188 - 0xbc
      12'h656: dout <= 8'b01110100; // 1622 : 116 - 0x74
      12'h657: dout <= 8'b11011100; // 1623 : 220 - 0xdc
      12'h658: dout <= 8'b00000000; // 1624 :   0 - 0x0 -- plane 1
      12'h659: dout <= 8'b00000000; // 1625 :   0 - 0x0
      12'h65A: dout <= 8'b00000000; // 1626 :   0 - 0x0
      12'h65B: dout <= 8'b00000000; // 1627 :   0 - 0x0
      12'h65C: dout <= 8'b00000000; // 1628 :   0 - 0x0
      12'h65D: dout <= 8'b00000000; // 1629 :   0 - 0x0
      12'h65E: dout <= 8'b00000000; // 1630 :   0 - 0x0
      12'h65F: dout <= 8'b00000000; // 1631 :   0 - 0x0
      12'h660: dout <= 8'b00011111; // 1632 :  31 - 0x1f -- Background 0x66
      12'h661: dout <= 8'b00001011; // 1633 :  11 - 0xb
      12'h662: dout <= 8'b00001111; // 1634 :  15 - 0xf
      12'h663: dout <= 8'b00000101; // 1635 :   5 - 0x5
      12'h664: dout <= 8'b00000011; // 1636 :   3 - 0x3
      12'h665: dout <= 8'b00000001; // 1637 :   1 - 0x1
      12'h666: dout <= 8'b00000000; // 1638 :   0 - 0x0
      12'h667: dout <= 8'b00000000; // 1639 :   0 - 0x0
      12'h668: dout <= 8'b00000000; // 1640 :   0 - 0x0 -- plane 1
      12'h669: dout <= 8'b00000000; // 1641 :   0 - 0x0
      12'h66A: dout <= 8'b00000000; // 1642 :   0 - 0x0
      12'h66B: dout <= 8'b00000000; // 1643 :   0 - 0x0
      12'h66C: dout <= 8'b00000000; // 1644 :   0 - 0x0
      12'h66D: dout <= 8'b00000000; // 1645 :   0 - 0x0
      12'h66E: dout <= 8'b00000000; // 1646 :   0 - 0x0
      12'h66F: dout <= 8'b00000000; // 1647 :   0 - 0x0
      12'h670: dout <= 8'b11111100; // 1648 : 252 - 0xfc -- Background 0x67
      12'h671: dout <= 8'b01101000; // 1649 : 104 - 0x68
      12'h672: dout <= 8'b11111000; // 1650 : 248 - 0xf8
      12'h673: dout <= 8'b10110000; // 1651 : 176 - 0xb0
      12'h674: dout <= 8'b11100000; // 1652 : 224 - 0xe0
      12'h675: dout <= 8'b10000000; // 1653 : 128 - 0x80
      12'h676: dout <= 8'b00000000; // 1654 :   0 - 0x0
      12'h677: dout <= 8'b00000000; // 1655 :   0 - 0x0
      12'h678: dout <= 8'b00000000; // 1656 :   0 - 0x0 -- plane 1
      12'h679: dout <= 8'b00000000; // 1657 :   0 - 0x0
      12'h67A: dout <= 8'b00000000; // 1658 :   0 - 0x0
      12'h67B: dout <= 8'b00000000; // 1659 :   0 - 0x0
      12'h67C: dout <= 8'b00000000; // 1660 :   0 - 0x0
      12'h67D: dout <= 8'b00000000; // 1661 :   0 - 0x0
      12'h67E: dout <= 8'b00000000; // 1662 :   0 - 0x0
      12'h67F: dout <= 8'b00000000; // 1663 :   0 - 0x0
      12'h680: dout <= 8'b00000000; // 1664 :   0 - 0x0 -- Background 0x68
      12'h681: dout <= 8'b00000000; // 1665 :   0 - 0x0
      12'h682: dout <= 8'b00000000; // 1666 :   0 - 0x0
      12'h683: dout <= 8'b00000000; // 1667 :   0 - 0x0
      12'h684: dout <= 8'b00000000; // 1668 :   0 - 0x0
      12'h685: dout <= 8'b00000000; // 1669 :   0 - 0x0
      12'h686: dout <= 8'b00000000; // 1670 :   0 - 0x0
      12'h687: dout <= 8'b00000000; // 1671 :   0 - 0x0
      12'h688: dout <= 8'b00000000; // 1672 :   0 - 0x0 -- plane 1
      12'h689: dout <= 8'b00000000; // 1673 :   0 - 0x0
      12'h68A: dout <= 8'b00000000; // 1674 :   0 - 0x0
      12'h68B: dout <= 8'b00000001; // 1675 :   1 - 0x1
      12'h68C: dout <= 8'b00000001; // 1676 :   1 - 0x1
      12'h68D: dout <= 8'b00001011; // 1677 :  11 - 0xb
      12'h68E: dout <= 8'b00011100; // 1678 :  28 - 0x1c
      12'h68F: dout <= 8'b00111111; // 1679 :  63 - 0x3f
      12'h690: dout <= 8'b00000000; // 1680 :   0 - 0x0 -- Background 0x69
      12'h691: dout <= 8'b00000000; // 1681 :   0 - 0x0
      12'h692: dout <= 8'b00000000; // 1682 :   0 - 0x0
      12'h693: dout <= 8'b00000000; // 1683 :   0 - 0x0
      12'h694: dout <= 8'b00000000; // 1684 :   0 - 0x0
      12'h695: dout <= 8'b00000000; // 1685 :   0 - 0x0
      12'h696: dout <= 8'b00000000; // 1686 :   0 - 0x0
      12'h697: dout <= 8'b00000000; // 1687 :   0 - 0x0
      12'h698: dout <= 8'b00000000; // 1688 :   0 - 0x0 -- plane 1
      12'h699: dout <= 8'b00000000; // 1689 :   0 - 0x0
      12'h69A: dout <= 8'b00110000; // 1690 :  48 - 0x30
      12'h69B: dout <= 8'b01111000; // 1691 : 120 - 0x78
      12'h69C: dout <= 8'b10000000; // 1692 : 128 - 0x80
      12'h69D: dout <= 8'b11110000; // 1693 : 240 - 0xf0
      12'h69E: dout <= 8'b11111000; // 1694 : 248 - 0xf8
      12'h69F: dout <= 8'b11111100; // 1695 : 252 - 0xfc
      12'h6A0: dout <= 8'b00000000; // 1696 :   0 - 0x0 -- Background 0x6a
      12'h6A1: dout <= 8'b00000000; // 1697 :   0 - 0x0
      12'h6A2: dout <= 8'b00000000; // 1698 :   0 - 0x0
      12'h6A3: dout <= 8'b00000000; // 1699 :   0 - 0x0
      12'h6A4: dout <= 8'b00000000; // 1700 :   0 - 0x0
      12'h6A5: dout <= 8'b00000000; // 1701 :   0 - 0x0
      12'h6A6: dout <= 8'b00000000; // 1702 :   0 - 0x0
      12'h6A7: dout <= 8'b00000000; // 1703 :   0 - 0x0
      12'h6A8: dout <= 8'b00111111; // 1704 :  63 - 0x3f -- plane 1
      12'h6A9: dout <= 8'b00111111; // 1705 :  63 - 0x3f
      12'h6AA: dout <= 8'b00111111; // 1706 :  63 - 0x3f
      12'h6AB: dout <= 8'b00011111; // 1707 :  31 - 0x1f
      12'h6AC: dout <= 8'b00011111; // 1708 :  31 - 0x1f
      12'h6AD: dout <= 8'b00000111; // 1709 :   7 - 0x7
      12'h6AE: dout <= 8'b00000000; // 1710 :   0 - 0x0
      12'h6AF: dout <= 8'b00000000; // 1711 :   0 - 0x0
      12'h6B0: dout <= 8'b00000000; // 1712 :   0 - 0x0 -- Background 0x6b
      12'h6B1: dout <= 8'b00000000; // 1713 :   0 - 0x0
      12'h6B2: dout <= 8'b00000000; // 1714 :   0 - 0x0
      12'h6B3: dout <= 8'b00000000; // 1715 :   0 - 0x0
      12'h6B4: dout <= 8'b00000000; // 1716 :   0 - 0x0
      12'h6B5: dout <= 8'b00000000; // 1717 :   0 - 0x0
      12'h6B6: dout <= 8'b00000000; // 1718 :   0 - 0x0
      12'h6B7: dout <= 8'b00000000; // 1719 :   0 - 0x0
      12'h6B8: dout <= 8'b11111100; // 1720 : 252 - 0xfc -- plane 1
      12'h6B9: dout <= 8'b11101100; // 1721 : 236 - 0xec
      12'h6BA: dout <= 8'b11101100; // 1722 : 236 - 0xec
      12'h6BB: dout <= 8'b11011000; // 1723 : 216 - 0xd8
      12'h6BC: dout <= 8'b11111000; // 1724 : 248 - 0xf8
      12'h6BD: dout <= 8'b11100000; // 1725 : 224 - 0xe0
      12'h6BE: dout <= 8'b00000000; // 1726 :   0 - 0x0
      12'h6BF: dout <= 8'b00000000; // 1727 :   0 - 0x0
      12'h6C0: dout <= 8'b00000000; // 1728 :   0 - 0x0 -- Background 0x6c
      12'h6C1: dout <= 8'b00000000; // 1729 :   0 - 0x0
      12'h6C2: dout <= 8'b00000001; // 1730 :   1 - 0x1
      12'h6C3: dout <= 8'b00011101; // 1731 :  29 - 0x1d
      12'h6C4: dout <= 8'b00111110; // 1732 :  62 - 0x3e
      12'h6C5: dout <= 8'b00111111; // 1733 :  63 - 0x3f
      12'h6C6: dout <= 8'b00111111; // 1734 :  63 - 0x3f
      12'h6C7: dout <= 8'b00111111; // 1735 :  63 - 0x3f
      12'h6C8: dout <= 8'b00000000; // 1736 :   0 - 0x0 -- plane 1
      12'h6C9: dout <= 8'b00000000; // 1737 :   0 - 0x0
      12'h6CA: dout <= 8'b00000001; // 1738 :   1 - 0x1
      12'h6CB: dout <= 8'b00011101; // 1739 :  29 - 0x1d
      12'h6CC: dout <= 8'b00111110; // 1740 :  62 - 0x3e
      12'h6CD: dout <= 8'b00111111; // 1741 :  63 - 0x3f
      12'h6CE: dout <= 8'b00111111; // 1742 :  63 - 0x3f
      12'h6CF: dout <= 8'b00111111; // 1743 :  63 - 0x3f
      12'h6D0: dout <= 8'b00000000; // 1744 :   0 - 0x0 -- Background 0x6d
      12'h6D1: dout <= 8'b10000000; // 1745 : 128 - 0x80
      12'h6D2: dout <= 8'b00000000; // 1746 :   0 - 0x0
      12'h6D3: dout <= 8'b01110000; // 1747 : 112 - 0x70
      12'h6D4: dout <= 8'b11111000; // 1748 : 248 - 0xf8
      12'h6D5: dout <= 8'b11111100; // 1749 : 252 - 0xfc
      12'h6D6: dout <= 8'b11111100; // 1750 : 252 - 0xfc
      12'h6D7: dout <= 8'b11111100; // 1751 : 252 - 0xfc
      12'h6D8: dout <= 8'b00000000; // 1752 :   0 - 0x0 -- plane 1
      12'h6D9: dout <= 8'b10000000; // 1753 : 128 - 0x80
      12'h6DA: dout <= 8'b00000000; // 1754 :   0 - 0x0
      12'h6DB: dout <= 8'b01110000; // 1755 : 112 - 0x70
      12'h6DC: dout <= 8'b11111000; // 1756 : 248 - 0xf8
      12'h6DD: dout <= 8'b11111100; // 1757 : 252 - 0xfc
      12'h6DE: dout <= 8'b11111100; // 1758 : 252 - 0xfc
      12'h6DF: dout <= 8'b11111100; // 1759 : 252 - 0xfc
      12'h6E0: dout <= 8'b00111111; // 1760 :  63 - 0x3f -- Background 0x6e
      12'h6E1: dout <= 8'b00111111; // 1761 :  63 - 0x3f
      12'h6E2: dout <= 8'b00011111; // 1762 :  31 - 0x1f
      12'h6E3: dout <= 8'b00011111; // 1763 :  31 - 0x1f
      12'h6E4: dout <= 8'b00001111; // 1764 :  15 - 0xf
      12'h6E5: dout <= 8'b00000110; // 1765 :   6 - 0x6
      12'h6E6: dout <= 8'b00000000; // 1766 :   0 - 0x0
      12'h6E7: dout <= 8'b00000000; // 1767 :   0 - 0x0
      12'h6E8: dout <= 8'b00111111; // 1768 :  63 - 0x3f -- plane 1
      12'h6E9: dout <= 8'b00111111; // 1769 :  63 - 0x3f
      12'h6EA: dout <= 8'b00011111; // 1770 :  31 - 0x1f
      12'h6EB: dout <= 8'b00011111; // 1771 :  31 - 0x1f
      12'h6EC: dout <= 8'b00001111; // 1772 :  15 - 0xf
      12'h6ED: dout <= 8'b00000110; // 1773 :   6 - 0x6
      12'h6EE: dout <= 8'b00000000; // 1774 :   0 - 0x0
      12'h6EF: dout <= 8'b00000000; // 1775 :   0 - 0x0
      12'h6F0: dout <= 8'b11101100; // 1776 : 236 - 0xec -- Background 0x6f
      12'h6F1: dout <= 8'b11101100; // 1777 : 236 - 0xec
      12'h6F2: dout <= 8'b11011000; // 1778 : 216 - 0xd8
      12'h6F3: dout <= 8'b11111000; // 1779 : 248 - 0xf8
      12'h6F4: dout <= 8'b11110000; // 1780 : 240 - 0xf0
      12'h6F5: dout <= 8'b11100000; // 1781 : 224 - 0xe0
      12'h6F6: dout <= 8'b00000000; // 1782 :   0 - 0x0
      12'h6F7: dout <= 8'b00000000; // 1783 :   0 - 0x0
      12'h6F8: dout <= 8'b11101100; // 1784 : 236 - 0xec -- plane 1
      12'h6F9: dout <= 8'b11101100; // 1785 : 236 - 0xec
      12'h6FA: dout <= 8'b11011000; // 1786 : 216 - 0xd8
      12'h6FB: dout <= 8'b11111000; // 1787 : 248 - 0xf8
      12'h6FC: dout <= 8'b11110000; // 1788 : 240 - 0xf0
      12'h6FD: dout <= 8'b11100000; // 1789 : 224 - 0xe0
      12'h6FE: dout <= 8'b00000000; // 1790 :   0 - 0x0
      12'h6FF: dout <= 8'b00000000; // 1791 :   0 - 0x0
      12'h700: dout <= 8'b00000000; // 1792 :   0 - 0x0 -- Background 0x70
      12'h701: dout <= 8'b00000100; // 1793 :   4 - 0x4
      12'h702: dout <= 8'b00000011; // 1794 :   3 - 0x3
      12'h703: dout <= 8'b00000000; // 1795 :   0 - 0x0
      12'h704: dout <= 8'b00000001; // 1796 :   1 - 0x1
      12'h705: dout <= 8'b00000111; // 1797 :   7 - 0x7
      12'h706: dout <= 8'b00001111; // 1798 :  15 - 0xf
      12'h707: dout <= 8'b00001100; // 1799 :  12 - 0xc
      12'h708: dout <= 8'b00000000; // 1800 :   0 - 0x0 -- plane 1
      12'h709: dout <= 8'b00000000; // 1801 :   0 - 0x0
      12'h70A: dout <= 8'b00000000; // 1802 :   0 - 0x0
      12'h70B: dout <= 8'b00000000; // 1803 :   0 - 0x0
      12'h70C: dout <= 8'b00000000; // 1804 :   0 - 0x0
      12'h70D: dout <= 8'b00000000; // 1805 :   0 - 0x0
      12'h70E: dout <= 8'b00000000; // 1806 :   0 - 0x0
      12'h70F: dout <= 8'b00000000; // 1807 :   0 - 0x0
      12'h710: dout <= 8'b00000000; // 1808 :   0 - 0x0 -- Background 0x71
      12'h711: dout <= 8'b00000000; // 1809 :   0 - 0x0
      12'h712: dout <= 8'b11100000; // 1810 : 224 - 0xe0
      12'h713: dout <= 8'b10000000; // 1811 : 128 - 0x80
      12'h714: dout <= 8'b01000000; // 1812 :  64 - 0x40
      12'h715: dout <= 8'b11110000; // 1813 : 240 - 0xf0
      12'h716: dout <= 8'b10011000; // 1814 : 152 - 0x98
      12'h717: dout <= 8'b11111000; // 1815 : 248 - 0xf8
      12'h718: dout <= 8'b00000000; // 1816 :   0 - 0x0 -- plane 1
      12'h719: dout <= 8'b00000000; // 1817 :   0 - 0x0
      12'h71A: dout <= 8'b00000000; // 1818 :   0 - 0x0
      12'h71B: dout <= 8'b00000000; // 1819 :   0 - 0x0
      12'h71C: dout <= 8'b00000000; // 1820 :   0 - 0x0
      12'h71D: dout <= 8'b00000000; // 1821 :   0 - 0x0
      12'h71E: dout <= 8'b00000000; // 1822 :   0 - 0x0
      12'h71F: dout <= 8'b00000000; // 1823 :   0 - 0x0
      12'h720: dout <= 8'b00011111; // 1824 :  31 - 0x1f -- Background 0x72
      12'h721: dout <= 8'b00010011; // 1825 :  19 - 0x13
      12'h722: dout <= 8'b00011111; // 1826 :  31 - 0x1f
      12'h723: dout <= 8'b00001111; // 1827 :  15 - 0xf
      12'h724: dout <= 8'b00001001; // 1828 :   9 - 0x9
      12'h725: dout <= 8'b00000111; // 1829 :   7 - 0x7
      12'h726: dout <= 8'b00000001; // 1830 :   1 - 0x1
      12'h727: dout <= 8'b00000000; // 1831 :   0 - 0x0
      12'h728: dout <= 8'b00000000; // 1832 :   0 - 0x0 -- plane 1
      12'h729: dout <= 8'b00000000; // 1833 :   0 - 0x0
      12'h72A: dout <= 8'b00000000; // 1834 :   0 - 0x0
      12'h72B: dout <= 8'b00000000; // 1835 :   0 - 0x0
      12'h72C: dout <= 8'b00000000; // 1836 :   0 - 0x0
      12'h72D: dout <= 8'b00000000; // 1837 :   0 - 0x0
      12'h72E: dout <= 8'b00000000; // 1838 :   0 - 0x0
      12'h72F: dout <= 8'b00000000; // 1839 :   0 - 0x0
      12'h730: dout <= 8'b11100100; // 1840 : 228 - 0xe4 -- Background 0x73
      12'h731: dout <= 8'b00111100; // 1841 :  60 - 0x3c
      12'h732: dout <= 8'b11100100; // 1842 : 228 - 0xe4
      12'h733: dout <= 8'b00111000; // 1843 :  56 - 0x38
      12'h734: dout <= 8'b11111000; // 1844 : 248 - 0xf8
      12'h735: dout <= 8'b11110000; // 1845 : 240 - 0xf0
      12'h736: dout <= 8'b11000000; // 1846 : 192 - 0xc0
      12'h737: dout <= 8'b00000000; // 1847 :   0 - 0x0
      12'h738: dout <= 8'b00000000; // 1848 :   0 - 0x0 -- plane 1
      12'h739: dout <= 8'b00000000; // 1849 :   0 - 0x0
      12'h73A: dout <= 8'b00000000; // 1850 :   0 - 0x0
      12'h73B: dout <= 8'b00000000; // 1851 :   0 - 0x0
      12'h73C: dout <= 8'b00000000; // 1852 :   0 - 0x0
      12'h73D: dout <= 8'b00000000; // 1853 :   0 - 0x0
      12'h73E: dout <= 8'b00000000; // 1854 :   0 - 0x0
      12'h73F: dout <= 8'b00000000; // 1855 :   0 - 0x0
      12'h740: dout <= 8'b00000000; // 1856 :   0 - 0x0 -- Background 0x74
      12'h741: dout <= 8'b00000000; // 1857 :   0 - 0x0
      12'h742: dout <= 8'b00000000; // 1858 :   0 - 0x0
      12'h743: dout <= 8'b00000000; // 1859 :   0 - 0x0
      12'h744: dout <= 8'b00000000; // 1860 :   0 - 0x0
      12'h745: dout <= 8'b00000000; // 1861 :   0 - 0x0
      12'h746: dout <= 8'b00000000; // 1862 :   0 - 0x0
      12'h747: dout <= 8'b00000000; // 1863 :   0 - 0x0
      12'h748: dout <= 8'b00000000; // 1864 :   0 - 0x0 -- plane 1
      12'h749: dout <= 8'b00000000; // 1865 :   0 - 0x0
      12'h74A: dout <= 8'b00000000; // 1866 :   0 - 0x0
      12'h74B: dout <= 8'b00000000; // 1867 :   0 - 0x0
      12'h74C: dout <= 8'b00010001; // 1868 :  17 - 0x11
      12'h74D: dout <= 8'b00010011; // 1869 :  19 - 0x13
      12'h74E: dout <= 8'b00011111; // 1870 :  31 - 0x1f
      12'h74F: dout <= 8'b00011111; // 1871 :  31 - 0x1f
      12'h750: dout <= 8'b00000000; // 1872 :   0 - 0x0 -- Background 0x75
      12'h751: dout <= 8'b00000000; // 1873 :   0 - 0x0
      12'h752: dout <= 8'b00000000; // 1874 :   0 - 0x0
      12'h753: dout <= 8'b00000000; // 1875 :   0 - 0x0
      12'h754: dout <= 8'b00000000; // 1876 :   0 - 0x0
      12'h755: dout <= 8'b00000000; // 1877 :   0 - 0x0
      12'h756: dout <= 8'b00000000; // 1878 :   0 - 0x0
      12'h757: dout <= 8'b00000000; // 1879 :   0 - 0x0
      12'h758: dout <= 8'b00000000; // 1880 :   0 - 0x0 -- plane 1
      12'h759: dout <= 8'b00000000; // 1881 :   0 - 0x0
      12'h75A: dout <= 8'b00000000; // 1882 :   0 - 0x0
      12'h75B: dout <= 8'b10000000; // 1883 : 128 - 0x80
      12'h75C: dout <= 8'b11000100; // 1884 : 196 - 0xc4
      12'h75D: dout <= 8'b11100100; // 1885 : 228 - 0xe4
      12'h75E: dout <= 8'b11111100; // 1886 : 252 - 0xfc
      12'h75F: dout <= 8'b11111100; // 1887 : 252 - 0xfc
      12'h760: dout <= 8'b00000000; // 1888 :   0 - 0x0 -- Background 0x76
      12'h761: dout <= 8'b00000000; // 1889 :   0 - 0x0
      12'h762: dout <= 8'b00000000; // 1890 :   0 - 0x0
      12'h763: dout <= 8'b00000000; // 1891 :   0 - 0x0
      12'h764: dout <= 8'b00000000; // 1892 :   0 - 0x0
      12'h765: dout <= 8'b00000000; // 1893 :   0 - 0x0
      12'h766: dout <= 8'b00000000; // 1894 :   0 - 0x0
      12'h767: dout <= 8'b00000000; // 1895 :   0 - 0x0
      12'h768: dout <= 8'b00011111; // 1896 :  31 - 0x1f -- plane 1
      12'h769: dout <= 8'b00001110; // 1897 :  14 - 0xe
      12'h76A: dout <= 8'b00000110; // 1898 :   6 - 0x6
      12'h76B: dout <= 8'b00000010; // 1899 :   2 - 0x2
      12'h76C: dout <= 8'b00000000; // 1900 :   0 - 0x0
      12'h76D: dout <= 8'b00000000; // 1901 :   0 - 0x0
      12'h76E: dout <= 8'b00000000; // 1902 :   0 - 0x0
      12'h76F: dout <= 8'b00000000; // 1903 :   0 - 0x0
      12'h770: dout <= 8'b00000000; // 1904 :   0 - 0x0 -- Background 0x77
      12'h771: dout <= 8'b00000000; // 1905 :   0 - 0x0
      12'h772: dout <= 8'b00000000; // 1906 :   0 - 0x0
      12'h773: dout <= 8'b00000000; // 1907 :   0 - 0x0
      12'h774: dout <= 8'b00000000; // 1908 :   0 - 0x0
      12'h775: dout <= 8'b00000000; // 1909 :   0 - 0x0
      12'h776: dout <= 8'b00000000; // 1910 :   0 - 0x0
      12'h777: dout <= 8'b00000000; // 1911 :   0 - 0x0
      12'h778: dout <= 8'b11111100; // 1912 : 252 - 0xfc -- plane 1
      12'h779: dout <= 8'b10111000; // 1913 : 184 - 0xb8
      12'h77A: dout <= 8'b10110000; // 1914 : 176 - 0xb0
      12'h77B: dout <= 8'b10100000; // 1915 : 160 - 0xa0
      12'h77C: dout <= 8'b10000000; // 1916 : 128 - 0x80
      12'h77D: dout <= 8'b00000000; // 1917 :   0 - 0x0
      12'h77E: dout <= 8'b00000000; // 1918 :   0 - 0x0
      12'h77F: dout <= 8'b00000000; // 1919 :   0 - 0x0
      12'h780: dout <= 8'b00000000; // 1920 :   0 - 0x0 -- Background 0x78
      12'h781: dout <= 8'b00000000; // 1921 :   0 - 0x0
      12'h782: dout <= 8'b00000000; // 1922 :   0 - 0x0
      12'h783: dout <= 8'b00000000; // 1923 :   0 - 0x0
      12'h784: dout <= 8'b00000000; // 1924 :   0 - 0x0
      12'h785: dout <= 8'b00000000; // 1925 :   0 - 0x0
      12'h786: dout <= 8'b00000000; // 1926 :   0 - 0x0
      12'h787: dout <= 8'b00000000; // 1927 :   0 - 0x0
      12'h788: dout <= 8'b00000000; // 1928 :   0 - 0x0 -- plane 1
      12'h789: dout <= 8'b00000000; // 1929 :   0 - 0x0
      12'h78A: dout <= 8'b00000000; // 1930 :   0 - 0x0
      12'h78B: dout <= 8'b00000001; // 1931 :   1 - 0x1
      12'h78C: dout <= 8'b00000011; // 1932 :   3 - 0x3
      12'h78D: dout <= 8'b00000110; // 1933 :   6 - 0x6
      12'h78E: dout <= 8'b00000110; // 1934 :   6 - 0x6
      12'h78F: dout <= 8'b00001111; // 1935 :  15 - 0xf
      12'h790: dout <= 8'b00000000; // 1936 :   0 - 0x0 -- Background 0x79
      12'h791: dout <= 8'b00000000; // 1937 :   0 - 0x0
      12'h792: dout <= 8'b00000000; // 1938 :   0 - 0x0
      12'h793: dout <= 8'b00000000; // 1939 :   0 - 0x0
      12'h794: dout <= 8'b00000000; // 1940 :   0 - 0x0
      12'h795: dout <= 8'b00000000; // 1941 :   0 - 0x0
      12'h796: dout <= 8'b00000000; // 1942 :   0 - 0x0
      12'h797: dout <= 8'b00000000; // 1943 :   0 - 0x0
      12'h798: dout <= 8'b00000000; // 1944 :   0 - 0x0 -- plane 1
      12'h799: dout <= 8'b00011000; // 1945 :  24 - 0x18
      12'h79A: dout <= 8'b11110100; // 1946 : 244 - 0xf4
      12'h79B: dout <= 8'b11111000; // 1947 : 248 - 0xf8
      12'h79C: dout <= 8'b00111000; // 1948 :  56 - 0x38
      12'h79D: dout <= 8'b01111100; // 1949 : 124 - 0x7c
      12'h79E: dout <= 8'b11111100; // 1950 : 252 - 0xfc
      12'h79F: dout <= 8'b11111100; // 1951 : 252 - 0xfc
      12'h7A0: dout <= 8'b00000000; // 1952 :   0 - 0x0 -- Background 0x7a
      12'h7A1: dout <= 8'b00000000; // 1953 :   0 - 0x0
      12'h7A2: dout <= 8'b00000000; // 1954 :   0 - 0x0
      12'h7A3: dout <= 8'b00000000; // 1955 :   0 - 0x0
      12'h7A4: dout <= 8'b00000000; // 1956 :   0 - 0x0
      12'h7A5: dout <= 8'b00000000; // 1957 :   0 - 0x0
      12'h7A6: dout <= 8'b00000000; // 1958 :   0 - 0x0
      12'h7A7: dout <= 8'b00000000; // 1959 :   0 - 0x0
      12'h7A8: dout <= 8'b00001111; // 1960 :  15 - 0xf -- plane 1
      12'h7A9: dout <= 8'b00011111; // 1961 :  31 - 0x1f
      12'h7AA: dout <= 8'b00110000; // 1962 :  48 - 0x30
      12'h7AB: dout <= 8'b00111000; // 1963 :  56 - 0x38
      12'h7AC: dout <= 8'b00011101; // 1964 :  29 - 0x1d
      12'h7AD: dout <= 8'b00000011; // 1965 :   3 - 0x3
      12'h7AE: dout <= 8'b00000011; // 1966 :   3 - 0x3
      12'h7AF: dout <= 8'b00000000; // 1967 :   0 - 0x0
      12'h7B0: dout <= 8'b00000000; // 1968 :   0 - 0x0 -- Background 0x7b
      12'h7B1: dout <= 8'b00000000; // 1969 :   0 - 0x0
      12'h7B2: dout <= 8'b00000000; // 1970 :   0 - 0x0
      12'h7B3: dout <= 8'b00000000; // 1971 :   0 - 0x0
      12'h7B4: dout <= 8'b00000000; // 1972 :   0 - 0x0
      12'h7B5: dout <= 8'b00000000; // 1973 :   0 - 0x0
      12'h7B6: dout <= 8'b00000000; // 1974 :   0 - 0x0
      12'h7B7: dout <= 8'b00000000; // 1975 :   0 - 0x0
      12'h7B8: dout <= 8'b11111100; // 1976 : 252 - 0xfc -- plane 1
      12'h7B9: dout <= 8'b11111100; // 1977 : 252 - 0xfc
      12'h7BA: dout <= 8'b01111100; // 1978 : 124 - 0x7c
      12'h7BB: dout <= 8'b10001110; // 1979 : 142 - 0x8e
      12'h7BC: dout <= 8'b10000110; // 1980 : 134 - 0x86
      12'h7BD: dout <= 8'b10011100; // 1981 : 156 - 0x9c
      12'h7BE: dout <= 8'b01111000; // 1982 : 120 - 0x78
      12'h7BF: dout <= 8'b00000000; // 1983 :   0 - 0x0
      12'h7C0: dout <= 8'b00000000; // 1984 :   0 - 0x0 -- Background 0x7c
      12'h7C1: dout <= 8'b00000001; // 1985 :   1 - 0x1
      12'h7C2: dout <= 8'b00000110; // 1986 :   6 - 0x6
      12'h7C3: dout <= 8'b00000111; // 1987 :   7 - 0x7
      12'h7C4: dout <= 8'b00000111; // 1988 :   7 - 0x7
      12'h7C5: dout <= 8'b00000111; // 1989 :   7 - 0x7
      12'h7C6: dout <= 8'b00000001; // 1990 :   1 - 0x1
      12'h7C7: dout <= 8'b00000011; // 1991 :   3 - 0x3
      12'h7C8: dout <= 8'b00000000; // 1992 :   0 - 0x0 -- plane 1
      12'h7C9: dout <= 8'b00000001; // 1993 :   1 - 0x1
      12'h7CA: dout <= 8'b00000110; // 1994 :   6 - 0x6
      12'h7CB: dout <= 8'b00000111; // 1995 :   7 - 0x7
      12'h7CC: dout <= 8'b00000111; // 1996 :   7 - 0x7
      12'h7CD: dout <= 8'b00000111; // 1997 :   7 - 0x7
      12'h7CE: dout <= 8'b00000001; // 1998 :   1 - 0x1
      12'h7CF: dout <= 8'b00000011; // 1999 :   3 - 0x3
      12'h7D0: dout <= 8'b00000000; // 2000 :   0 - 0x0 -- Background 0x7d
      12'h7D1: dout <= 8'b11000000; // 2001 : 192 - 0xc0
      12'h7D2: dout <= 8'b00110000; // 2002 :  48 - 0x30
      12'h7D3: dout <= 8'b11110000; // 2003 : 240 - 0xf0
      12'h7D4: dout <= 8'b11110000; // 2004 : 240 - 0xf0
      12'h7D5: dout <= 8'b11110000; // 2005 : 240 - 0xf0
      12'h7D6: dout <= 8'b01000000; // 2006 :  64 - 0x40
      12'h7D7: dout <= 8'b01000000; // 2007 :  64 - 0x40
      12'h7D8: dout <= 8'b00000000; // 2008 :   0 - 0x0 -- plane 1
      12'h7D9: dout <= 8'b11000000; // 2009 : 192 - 0xc0
      12'h7DA: dout <= 8'b00110000; // 2010 :  48 - 0x30
      12'h7DB: dout <= 8'b11110000; // 2011 : 240 - 0xf0
      12'h7DC: dout <= 8'b11110000; // 2012 : 240 - 0xf0
      12'h7DD: dout <= 8'b11110000; // 2013 : 240 - 0xf0
      12'h7DE: dout <= 8'b01000000; // 2014 :  64 - 0x40
      12'h7DF: dout <= 8'b01000000; // 2015 :  64 - 0x40
      12'h7E0: dout <= 8'b00000001; // 2016 :   1 - 0x1 -- Background 0x7e
      12'h7E1: dout <= 8'b00000000; // 2017 :   0 - 0x0
      12'h7E2: dout <= 8'b00000001; // 2018 :   1 - 0x1
      12'h7E3: dout <= 8'b00000011; // 2019 :   3 - 0x3
      12'h7E4: dout <= 8'b00000001; // 2020 :   1 - 0x1
      12'h7E5: dout <= 8'b00000000; // 2021 :   0 - 0x0
      12'h7E6: dout <= 8'b00000000; // 2022 :   0 - 0x0
      12'h7E7: dout <= 8'b00000000; // 2023 :   0 - 0x0
      12'h7E8: dout <= 8'b00000001; // 2024 :   1 - 0x1 -- plane 1
      12'h7E9: dout <= 8'b00000000; // 2025 :   0 - 0x0
      12'h7EA: dout <= 8'b00000001; // 2026 :   1 - 0x1
      12'h7EB: dout <= 8'b00000011; // 2027 :   3 - 0x3
      12'h7EC: dout <= 8'b00000001; // 2028 :   1 - 0x1
      12'h7ED: dout <= 8'b00000000; // 2029 :   0 - 0x0
      12'h7EE: dout <= 8'b00000000; // 2030 :   0 - 0x0
      12'h7EF: dout <= 8'b00000000; // 2031 :   0 - 0x0
      12'h7F0: dout <= 8'b01000000; // 2032 :  64 - 0x40 -- Background 0x7f
      12'h7F1: dout <= 8'b01000000; // 2033 :  64 - 0x40
      12'h7F2: dout <= 8'b01000000; // 2034 :  64 - 0x40
      12'h7F3: dout <= 8'b01000000; // 2035 :  64 - 0x40
      12'h7F4: dout <= 8'b01000000; // 2036 :  64 - 0x40
      12'h7F5: dout <= 8'b10000000; // 2037 : 128 - 0x80
      12'h7F6: dout <= 8'b00000000; // 2038 :   0 - 0x0
      12'h7F7: dout <= 8'b00000000; // 2039 :   0 - 0x0
      12'h7F8: dout <= 8'b01000000; // 2040 :  64 - 0x40 -- plane 1
      12'h7F9: dout <= 8'b01000000; // 2041 :  64 - 0x40
      12'h7FA: dout <= 8'b01000000; // 2042 :  64 - 0x40
      12'h7FB: dout <= 8'b01000000; // 2043 :  64 - 0x40
      12'h7FC: dout <= 8'b01000000; // 2044 :  64 - 0x40
      12'h7FD: dout <= 8'b10000000; // 2045 : 128 - 0x80
      12'h7FE: dout <= 8'b00000000; // 2046 :   0 - 0x0
      12'h7FF: dout <= 8'b00000000; // 2047 :   0 - 0x0
      12'h800: dout <= 8'b11111111; // 2048 : 255 - 0xff -- Background 0x80
      12'h801: dout <= 8'b11111111; // 2049 : 255 - 0xff
      12'h802: dout <= 8'b11111111; // 2050 : 255 - 0xff
      12'h803: dout <= 8'b11111111; // 2051 : 255 - 0xff
      12'h804: dout <= 8'b11000000; // 2052 : 192 - 0xc0
      12'h805: dout <= 8'b11000000; // 2053 : 192 - 0xc0
      12'h806: dout <= 8'b11000000; // 2054 : 192 - 0xc0
      12'h807: dout <= 8'b11000111; // 2055 : 199 - 0xc7
      12'h808: dout <= 8'b00000000; // 2056 :   0 - 0x0 -- plane 1
      12'h809: dout <= 8'b00000000; // 2057 :   0 - 0x0
      12'h80A: dout <= 8'b00000000; // 2058 :   0 - 0x0
      12'h80B: dout <= 8'b00000000; // 2059 :   0 - 0x0
      12'h80C: dout <= 8'b00000000; // 2060 :   0 - 0x0
      12'h80D: dout <= 8'b00011111; // 2061 :  31 - 0x1f
      12'h80E: dout <= 8'b00010000; // 2062 :  16 - 0x10
      12'h80F: dout <= 8'b00010111; // 2063 :  23 - 0x17
      12'h810: dout <= 8'b11111111; // 2064 : 255 - 0xff -- Background 0x81
      12'h811: dout <= 8'b11111111; // 2065 : 255 - 0xff
      12'h812: dout <= 8'b11111111; // 2066 : 255 - 0xff
      12'h813: dout <= 8'b11111111; // 2067 : 255 - 0xff
      12'h814: dout <= 8'b00000000; // 2068 :   0 - 0x0
      12'h815: dout <= 8'b00000000; // 2069 :   0 - 0x0
      12'h816: dout <= 8'b00000000; // 2070 :   0 - 0x0
      12'h817: dout <= 8'b11111111; // 2071 : 255 - 0xff
      12'h818: dout <= 8'b00000000; // 2072 :   0 - 0x0 -- plane 1
      12'h819: dout <= 8'b00000000; // 2073 :   0 - 0x0
      12'h81A: dout <= 8'b00000000; // 2074 :   0 - 0x0
      12'h81B: dout <= 8'b00000000; // 2075 :   0 - 0x0
      12'h81C: dout <= 8'b00000000; // 2076 :   0 - 0x0
      12'h81D: dout <= 8'b11111111; // 2077 : 255 - 0xff
      12'h81E: dout <= 8'b00000000; // 2078 :   0 - 0x0
      12'h81F: dout <= 8'b11111111; // 2079 : 255 - 0xff
      12'h820: dout <= 8'b11111111; // 2080 : 255 - 0xff -- Background 0x82
      12'h821: dout <= 8'b11111111; // 2081 : 255 - 0xff
      12'h822: dout <= 8'b11111111; // 2082 : 255 - 0xff
      12'h823: dout <= 8'b11111111; // 2083 : 255 - 0xff
      12'h824: dout <= 8'b01111111; // 2084 : 127 - 0x7f
      12'h825: dout <= 8'b00111111; // 2085 :  63 - 0x3f
      12'h826: dout <= 8'b00011111; // 2086 :  31 - 0x1f
      12'h827: dout <= 8'b11001111; // 2087 : 207 - 0xcf
      12'h828: dout <= 8'b00000000; // 2088 :   0 - 0x0 -- plane 1
      12'h829: dout <= 8'b00000000; // 2089 :   0 - 0x0
      12'h82A: dout <= 8'b00000000; // 2090 :   0 - 0x0
      12'h82B: dout <= 8'b00000000; // 2091 :   0 - 0x0
      12'h82C: dout <= 8'b00000000; // 2092 :   0 - 0x0
      12'h82D: dout <= 8'b10000000; // 2093 : 128 - 0x80
      12'h82E: dout <= 8'b00000000; // 2094 :   0 - 0x0
      12'h82F: dout <= 8'b11000000; // 2095 : 192 - 0xc0
      12'h830: dout <= 8'b11111111; // 2096 : 255 - 0xff -- Background 0x83
      12'h831: dout <= 8'b11111111; // 2097 : 255 - 0xff
      12'h832: dout <= 8'b11111111; // 2098 : 255 - 0xff
      12'h833: dout <= 8'b11110111; // 2099 : 247 - 0xf7
      12'h834: dout <= 8'b11110111; // 2100 : 247 - 0xf7
      12'h835: dout <= 8'b11100010; // 2101 : 226 - 0xe2
      12'h836: dout <= 8'b11100000; // 2102 : 224 - 0xe0
      12'h837: dout <= 8'b11000110; // 2103 : 198 - 0xc6
      12'h838: dout <= 8'b00000000; // 2104 :   0 - 0x0 -- plane 1
      12'h839: dout <= 8'b00000000; // 2105 :   0 - 0x0
      12'h83A: dout <= 8'b00000000; // 2106 :   0 - 0x0
      12'h83B: dout <= 8'b00000000; // 2107 :   0 - 0x0
      12'h83C: dout <= 8'b00000000; // 2108 :   0 - 0x0
      12'h83D: dout <= 8'b00001000; // 2109 :   8 - 0x8
      12'h83E: dout <= 8'b00001000; // 2110 :   8 - 0x8
      12'h83F: dout <= 8'b00010110; // 2111 :  22 - 0x16
      12'h840: dout <= 8'b11111111; // 2112 : 255 - 0xff -- Background 0x84
      12'h841: dout <= 8'b11111111; // 2113 : 255 - 0xff
      12'h842: dout <= 8'b11111111; // 2114 : 255 - 0xff
      12'h843: dout <= 8'b11111111; // 2115 : 255 - 0xff
      12'h844: dout <= 8'b10111111; // 2116 : 191 - 0xbf
      12'h845: dout <= 8'b10111111; // 2117 : 191 - 0xbf
      12'h846: dout <= 8'b00011111; // 2118 :  31 - 0x1f
      12'h847: dout <= 8'b00011111; // 2119 :  31 - 0x1f
      12'h848: dout <= 8'b00000000; // 2120 :   0 - 0x0 -- plane 1
      12'h849: dout <= 8'b00000000; // 2121 :   0 - 0x0
      12'h84A: dout <= 8'b00000000; // 2122 :   0 - 0x0
      12'h84B: dout <= 8'b00000000; // 2123 :   0 - 0x0
      12'h84C: dout <= 8'b00000000; // 2124 :   0 - 0x0
      12'h84D: dout <= 8'b00000000; // 2125 :   0 - 0x0
      12'h84E: dout <= 8'b01000000; // 2126 :  64 - 0x40
      12'h84F: dout <= 8'b11000000; // 2127 : 192 - 0xc0
      12'h850: dout <= 8'b11111111; // 2128 : 255 - 0xff -- Background 0x85
      12'h851: dout <= 8'b11111111; // 2129 : 255 - 0xff
      12'h852: dout <= 8'b11111111; // 2130 : 255 - 0xff
      12'h853: dout <= 8'b11111111; // 2131 : 255 - 0xff
      12'h854: dout <= 8'b11111110; // 2132 : 254 - 0xfe
      12'h855: dout <= 8'b11111000; // 2133 : 248 - 0xf8
      12'h856: dout <= 8'b11100000; // 2134 : 224 - 0xe0
      12'h857: dout <= 8'b11000000; // 2135 : 192 - 0xc0
      12'h858: dout <= 8'b00000000; // 2136 :   0 - 0x0 -- plane 1
      12'h859: dout <= 8'b00000000; // 2137 :   0 - 0x0
      12'h85A: dout <= 8'b00000000; // 2138 :   0 - 0x0
      12'h85B: dout <= 8'b00000000; // 2139 :   0 - 0x0
      12'h85C: dout <= 8'b00000000; // 2140 :   0 - 0x0
      12'h85D: dout <= 8'b00000001; // 2141 :   1 - 0x1
      12'h85E: dout <= 8'b00000111; // 2142 :   7 - 0x7
      12'h85F: dout <= 8'b00001100; // 2143 :  12 - 0xc
      12'h860: dout <= 8'b11111111; // 2144 : 255 - 0xff -- Background 0x86
      12'h861: dout <= 8'b11111111; // 2145 : 255 - 0xff
      12'h862: dout <= 8'b11111111; // 2146 : 255 - 0xff
      12'h863: dout <= 8'b11111111; // 2147 : 255 - 0xff
      12'h864: dout <= 8'b00000111; // 2148 :   7 - 0x7
      12'h865: dout <= 8'b00000000; // 2149 :   0 - 0x0
      12'h866: dout <= 8'b00111111; // 2150 :  63 - 0x3f
      12'h867: dout <= 8'b11111111; // 2151 : 255 - 0xff
      12'h868: dout <= 8'b00000000; // 2152 :   0 - 0x0 -- plane 1
      12'h869: dout <= 8'b00000000; // 2153 :   0 - 0x0
      12'h86A: dout <= 8'b00000000; // 2154 :   0 - 0x0
      12'h86B: dout <= 8'b00000000; // 2155 :   0 - 0x0
      12'h86C: dout <= 8'b00000000; // 2156 :   0 - 0x0
      12'h86D: dout <= 8'b11000000; // 2157 : 192 - 0xc0
      12'h86E: dout <= 8'b00111111; // 2158 :  63 - 0x3f
      12'h86F: dout <= 8'b11111111; // 2159 : 255 - 0xff
      12'h870: dout <= 8'b11111111; // 2160 : 255 - 0xff -- Background 0x87
      12'h871: dout <= 8'b11111111; // 2161 : 255 - 0xff
      12'h872: dout <= 8'b11111111; // 2162 : 255 - 0xff
      12'h873: dout <= 8'b11111111; // 2163 : 255 - 0xff
      12'h874: dout <= 8'b11111111; // 2164 : 255 - 0xff
      12'h875: dout <= 8'b11111111; // 2165 : 255 - 0xff
      12'h876: dout <= 8'b00111111; // 2166 :  63 - 0x3f
      12'h877: dout <= 8'b11001111; // 2167 : 207 - 0xcf
      12'h878: dout <= 8'b00000000; // 2168 :   0 - 0x0 -- plane 1
      12'h879: dout <= 8'b00000000; // 2169 :   0 - 0x0
      12'h87A: dout <= 8'b00000000; // 2170 :   0 - 0x0
      12'h87B: dout <= 8'b00000000; // 2171 :   0 - 0x0
      12'h87C: dout <= 8'b00000000; // 2172 :   0 - 0x0
      12'h87D: dout <= 8'b00000000; // 2173 :   0 - 0x0
      12'h87E: dout <= 8'b00000000; // 2174 :   0 - 0x0
      12'h87F: dout <= 8'b11000000; // 2175 : 192 - 0xc0
      12'h880: dout <= 8'b11111111; // 2176 : 255 - 0xff -- Background 0x88
      12'h881: dout <= 8'b11111111; // 2177 : 255 - 0xff
      12'h882: dout <= 8'b11111111; // 2178 : 255 - 0xff
      12'h883: dout <= 8'b11111111; // 2179 : 255 - 0xff
      12'h884: dout <= 8'b11111111; // 2180 : 255 - 0xff
      12'h885: dout <= 8'b11111111; // 2181 : 255 - 0xff
      12'h886: dout <= 8'b11111111; // 2182 : 255 - 0xff
      12'h887: dout <= 8'b11111111; // 2183 : 255 - 0xff
      12'h888: dout <= 8'b00000000; // 2184 :   0 - 0x0 -- plane 1
      12'h889: dout <= 8'b00000000; // 2185 :   0 - 0x0
      12'h88A: dout <= 8'b00000000; // 2186 :   0 - 0x0
      12'h88B: dout <= 8'b00000000; // 2187 :   0 - 0x0
      12'h88C: dout <= 8'b00000000; // 2188 :   0 - 0x0
      12'h88D: dout <= 8'b00000000; // 2189 :   0 - 0x0
      12'h88E: dout <= 8'b00000000; // 2190 :   0 - 0x0
      12'h88F: dout <= 8'b00000000; // 2191 :   0 - 0x0
      12'h890: dout <= 8'b11111111; // 2192 : 255 - 0xff -- Background 0x89
      12'h891: dout <= 8'b11111111; // 2193 : 255 - 0xff
      12'h892: dout <= 8'b11111111; // 2194 : 255 - 0xff
      12'h893: dout <= 8'b01110111; // 2195 : 119 - 0x77
      12'h894: dout <= 8'b00010011; // 2196 :  19 - 0x13
      12'h895: dout <= 8'b00000001; // 2197 :   1 - 0x1
      12'h896: dout <= 8'b00010000; // 2198 :  16 - 0x10
      12'h897: dout <= 8'b00011000; // 2199 :  24 - 0x18
      12'h898: dout <= 8'b00000000; // 2200 :   0 - 0x0 -- plane 1
      12'h899: dout <= 8'b00000000; // 2201 :   0 - 0x0
      12'h89A: dout <= 8'b00000000; // 2202 :   0 - 0x0
      12'h89B: dout <= 8'b00000000; // 2203 :   0 - 0x0
      12'h89C: dout <= 8'b00000000; // 2204 :   0 - 0x0
      12'h89D: dout <= 8'b01000100; // 2205 :  68 - 0x44
      12'h89E: dout <= 8'b01010110; // 2206 :  86 - 0x56
      12'h89F: dout <= 8'b01011011; // 2207 :  91 - 0x5b
      12'h8A0: dout <= 8'b11111111; // 2208 : 255 - 0xff -- Background 0x8a
      12'h8A1: dout <= 8'b11111111; // 2209 : 255 - 0xff
      12'h8A2: dout <= 8'b11111111; // 2210 : 255 - 0xff
      12'h8A3: dout <= 8'b11111111; // 2211 : 255 - 0xff
      12'h8A4: dout <= 8'b11111111; // 2212 : 255 - 0xff
      12'h8A5: dout <= 8'b11111111; // 2213 : 255 - 0xff
      12'h8A6: dout <= 8'b11111111; // 2214 : 255 - 0xff
      12'h8A7: dout <= 8'b01111111; // 2215 : 127 - 0x7f
      12'h8A8: dout <= 8'b00000000; // 2216 :   0 - 0x0 -- plane 1
      12'h8A9: dout <= 8'b00000000; // 2217 :   0 - 0x0
      12'h8AA: dout <= 8'b00000000; // 2218 :   0 - 0x0
      12'h8AB: dout <= 8'b00000000; // 2219 :   0 - 0x0
      12'h8AC: dout <= 8'b00000000; // 2220 :   0 - 0x0
      12'h8AD: dout <= 8'b00000000; // 2221 :   0 - 0x0
      12'h8AE: dout <= 8'b00000000; // 2222 :   0 - 0x0
      12'h8AF: dout <= 8'b00000000; // 2223 :   0 - 0x0
      12'h8B0: dout <= 8'b11111111; // 2224 : 255 - 0xff -- Background 0x8b
      12'h8B1: dout <= 8'b11111111; // 2225 : 255 - 0xff
      12'h8B2: dout <= 8'b11111111; // 2226 : 255 - 0xff
      12'h8B3: dout <= 8'b11110111; // 2227 : 247 - 0xf7
      12'h8B4: dout <= 8'b11100101; // 2228 : 229 - 0xe5
      12'h8B5: dout <= 8'b11000001; // 2229 : 193 - 0xc1
      12'h8B6: dout <= 8'b10000100; // 2230 : 132 - 0x84
      12'h8B7: dout <= 8'b00001100; // 2231 :  12 - 0xc
      12'h8B8: dout <= 8'b00000000; // 2232 :   0 - 0x0 -- plane 1
      12'h8B9: dout <= 8'b00000000; // 2233 :   0 - 0x0
      12'h8BA: dout <= 8'b00000000; // 2234 :   0 - 0x0
      12'h8BB: dout <= 8'b00000000; // 2235 :   0 - 0x0
      12'h8BC: dout <= 8'b00000000; // 2236 :   0 - 0x0
      12'h8BD: dout <= 8'b00010000; // 2237 :  16 - 0x10
      12'h8BE: dout <= 8'b00110100; // 2238 :  52 - 0x34
      12'h8BF: dout <= 8'b01101101; // 2239 : 109 - 0x6d
      12'h8C0: dout <= 8'b11111111; // 2240 : 255 - 0xff -- Background 0x8c
      12'h8C1: dout <= 8'b11111111; // 2241 : 255 - 0xff
      12'h8C2: dout <= 8'b11111111; // 2242 : 255 - 0xff
      12'h8C3: dout <= 8'b11111111; // 2243 : 255 - 0xff
      12'h8C4: dout <= 8'b11111111; // 2244 : 255 - 0xff
      12'h8C5: dout <= 8'b01111111; // 2245 : 127 - 0x7f
      12'h8C6: dout <= 8'b01111110; // 2246 : 126 - 0x7e
      12'h8C7: dout <= 8'b01111110; // 2247 : 126 - 0x7e
      12'h8C8: dout <= 8'b00000000; // 2248 :   0 - 0x0 -- plane 1
      12'h8C9: dout <= 8'b00000000; // 2249 :   0 - 0x0
      12'h8CA: dout <= 8'b00000000; // 2250 :   0 - 0x0
      12'h8CB: dout <= 8'b00000000; // 2251 :   0 - 0x0
      12'h8CC: dout <= 8'b00000000; // 2252 :   0 - 0x0
      12'h8CD: dout <= 8'b00000000; // 2253 :   0 - 0x0
      12'h8CE: dout <= 8'b00000000; // 2254 :   0 - 0x0
      12'h8CF: dout <= 8'b00000000; // 2255 :   0 - 0x0
      12'h8D0: dout <= 8'b11111111; // 2256 : 255 - 0xff -- Background 0x8d
      12'h8D1: dout <= 8'b11111111; // 2257 : 255 - 0xff
      12'h8D2: dout <= 8'b10111111; // 2258 : 191 - 0xbf
      12'h8D3: dout <= 8'b10110111; // 2259 : 183 - 0xb7
      12'h8D4: dout <= 8'b00010111; // 2260 :  23 - 0x17
      12'h8D5: dout <= 8'b00000011; // 2261 :   3 - 0x3
      12'h8D6: dout <= 8'b00100011; // 2262 :  35 - 0x23
      12'h8D7: dout <= 8'b00100001; // 2263 :  33 - 0x21
      12'h8D8: dout <= 8'b00000000; // 2264 :   0 - 0x0 -- plane 1
      12'h8D9: dout <= 8'b00000000; // 2265 :   0 - 0x0
      12'h8DA: dout <= 8'b00000000; // 2266 :   0 - 0x0
      12'h8DB: dout <= 8'b00000000; // 2267 :   0 - 0x0
      12'h8DC: dout <= 8'b01000000; // 2268 :  64 - 0x40
      12'h8DD: dout <= 8'b01001000; // 2269 :  72 - 0x48
      12'h8DE: dout <= 8'b10101000; // 2270 : 168 - 0xa8
      12'h8DF: dout <= 8'b10101100; // 2271 : 172 - 0xac
      12'h8E0: dout <= 8'b11111111; // 2272 : 255 - 0xff -- Background 0x8e
      12'h8E1: dout <= 8'b11111111; // 2273 : 255 - 0xff
      12'h8E2: dout <= 8'b11111011; // 2274 : 251 - 0xfb
      12'h8E3: dout <= 8'b11111001; // 2275 : 249 - 0xf9
      12'h8E4: dout <= 8'b11111000; // 2276 : 248 - 0xf8
      12'h8E5: dout <= 8'b11111000; // 2277 : 248 - 0xf8
      12'h8E6: dout <= 8'b11111000; // 2278 : 248 - 0xf8
      12'h8E7: dout <= 8'b11111000; // 2279 : 248 - 0xf8
      12'h8E8: dout <= 8'b00000000; // 2280 :   0 - 0x0 -- plane 1
      12'h8E9: dout <= 8'b00000000; // 2281 :   0 - 0x0
      12'h8EA: dout <= 8'b00000000; // 2282 :   0 - 0x0
      12'h8EB: dout <= 8'b00000000; // 2283 :   0 - 0x0
      12'h8EC: dout <= 8'b00000010; // 2284 :   2 - 0x2
      12'h8ED: dout <= 8'b00000010; // 2285 :   2 - 0x2
      12'h8EE: dout <= 8'b00000010; // 2286 :   2 - 0x2
      12'h8EF: dout <= 8'b00000010; // 2287 :   2 - 0x2
      12'h8F0: dout <= 8'b11111111; // 2288 : 255 - 0xff -- Background 0x8f
      12'h8F1: dout <= 8'b11111111; // 2289 : 255 - 0xff
      12'h8F2: dout <= 8'b01111000; // 2290 : 120 - 0x78
      12'h8F3: dout <= 8'b00111000; // 2291 :  56 - 0x38
      12'h8F4: dout <= 8'b00011000; // 2292 :  24 - 0x18
      12'h8F5: dout <= 8'b00001000; // 2293 :   8 - 0x8
      12'h8F6: dout <= 8'b10000000; // 2294 : 128 - 0x80
      12'h8F7: dout <= 8'b11000000; // 2295 : 192 - 0xc0
      12'h8F8: dout <= 8'b00000000; // 2296 :   0 - 0x0 -- plane 1
      12'h8F9: dout <= 8'b00000000; // 2297 :   0 - 0x0
      12'h8FA: dout <= 8'b00000000; // 2298 :   0 - 0x0
      12'h8FB: dout <= 8'b00000011; // 2299 :   3 - 0x3
      12'h8FC: dout <= 8'b01000011; // 2300 :  67 - 0x43
      12'h8FD: dout <= 8'b01100010; // 2301 :  98 - 0x62
      12'h8FE: dout <= 8'b10110010; // 2302 : 178 - 0xb2
      12'h8FF: dout <= 8'b11011010; // 2303 : 218 - 0xda
      12'h900: dout <= 8'b11111111; // 2304 : 255 - 0xff -- Background 0x90
      12'h901: dout <= 8'b11111111; // 2305 : 255 - 0xff
      12'h902: dout <= 8'b00000001; // 2306 :   1 - 0x1
      12'h903: dout <= 8'b00000001; // 2307 :   1 - 0x1
      12'h904: dout <= 8'b00000001; // 2308 :   1 - 0x1
      12'h905: dout <= 8'b00000000; // 2309 :   0 - 0x0
      12'h906: dout <= 8'b11111111; // 2310 : 255 - 0xff
      12'h907: dout <= 8'b11111111; // 2311 : 255 - 0xff
      12'h908: dout <= 8'b00000000; // 2312 :   0 - 0x0 -- plane 1
      12'h909: dout <= 8'b00000000; // 2313 :   0 - 0x0
      12'h90A: dout <= 8'b00000000; // 2314 :   0 - 0x0
      12'h90B: dout <= 8'b11111100; // 2315 : 252 - 0xfc
      12'h90C: dout <= 8'b11111100; // 2316 : 252 - 0xfc
      12'h90D: dout <= 8'b00000000; // 2317 :   0 - 0x0
      12'h90E: dout <= 8'b11111111; // 2318 : 255 - 0xff
      12'h90F: dout <= 8'b11111111; // 2319 : 255 - 0xff
      12'h910: dout <= 8'b11111111; // 2320 : 255 - 0xff -- Background 0x91
      12'h911: dout <= 8'b11111111; // 2321 : 255 - 0xff
      12'h912: dout <= 8'b11111111; // 2322 : 255 - 0xff
      12'h913: dout <= 8'b11111111; // 2323 : 255 - 0xff
      12'h914: dout <= 8'b11111111; // 2324 : 255 - 0xff
      12'h915: dout <= 8'b11111111; // 2325 : 255 - 0xff
      12'h916: dout <= 8'b01111111; // 2326 : 127 - 0x7f
      12'h917: dout <= 8'b00111111; // 2327 :  63 - 0x3f
      12'h918: dout <= 8'b00000000; // 2328 :   0 - 0x0 -- plane 1
      12'h919: dout <= 8'b00000000; // 2329 :   0 - 0x0
      12'h91A: dout <= 8'b00000000; // 2330 :   0 - 0x0
      12'h91B: dout <= 8'b00000000; // 2331 :   0 - 0x0
      12'h91C: dout <= 8'b00000000; // 2332 :   0 - 0x0
      12'h91D: dout <= 8'b00000000; // 2333 :   0 - 0x0
      12'h91E: dout <= 8'b00000000; // 2334 :   0 - 0x0
      12'h91F: dout <= 8'b00000000; // 2335 :   0 - 0x0
      12'h920: dout <= 8'b11000111; // 2336 : 199 - 0xc7 -- Background 0x92
      12'h921: dout <= 8'b11000111; // 2337 : 199 - 0xc7
      12'h922: dout <= 8'b11000111; // 2338 : 199 - 0xc7
      12'h923: dout <= 8'b11000111; // 2339 : 199 - 0xc7
      12'h924: dout <= 8'b11000111; // 2340 : 199 - 0xc7
      12'h925: dout <= 8'b11000111; // 2341 : 199 - 0xc7
      12'h926: dout <= 8'b11000111; // 2342 : 199 - 0xc7
      12'h927: dout <= 8'b11000111; // 2343 : 199 - 0xc7
      12'h928: dout <= 8'b00010111; // 2344 :  23 - 0x17 -- plane 1
      12'h929: dout <= 8'b00010111; // 2345 :  23 - 0x17
      12'h92A: dout <= 8'b00010111; // 2346 :  23 - 0x17
      12'h92B: dout <= 8'b00010111; // 2347 :  23 - 0x17
      12'h92C: dout <= 8'b00010111; // 2348 :  23 - 0x17
      12'h92D: dout <= 8'b00010111; // 2349 :  23 - 0x17
      12'h92E: dout <= 8'b00010111; // 2350 :  23 - 0x17
      12'h92F: dout <= 8'b00010111; // 2351 :  23 - 0x17
      12'h930: dout <= 8'b11111111; // 2352 : 255 - 0xff -- Background 0x93
      12'h931: dout <= 8'b11111111; // 2353 : 255 - 0xff
      12'h932: dout <= 8'b11111111; // 2354 : 255 - 0xff
      12'h933: dout <= 8'b11111111; // 2355 : 255 - 0xff
      12'h934: dout <= 8'b11111001; // 2356 : 249 - 0xf9
      12'h935: dout <= 8'b11111001; // 2357 : 249 - 0xf9
      12'h936: dout <= 8'b11111111; // 2358 : 255 - 0xff
      12'h937: dout <= 8'b11111111; // 2359 : 255 - 0xff
      12'h938: dout <= 8'b11111111; // 2360 : 255 - 0xff -- plane 1
      12'h939: dout <= 8'b11111111; // 2361 : 255 - 0xff
      12'h93A: dout <= 8'b11111111; // 2362 : 255 - 0xff
      12'h93B: dout <= 8'b11111111; // 2363 : 255 - 0xff
      12'h93C: dout <= 8'b11111001; // 2364 : 249 - 0xf9
      12'h93D: dout <= 8'b11111001; // 2365 : 249 - 0xf9
      12'h93E: dout <= 8'b11111111; // 2366 : 255 - 0xff
      12'h93F: dout <= 8'b11111111; // 2367 : 255 - 0xff
      12'h940: dout <= 8'b11110111; // 2368 : 247 - 0xf7 -- Background 0x94
      12'h941: dout <= 8'b11111011; // 2369 : 251 - 0xfb
      12'h942: dout <= 8'b11111011; // 2370 : 251 - 0xfb
      12'h943: dout <= 8'b11111101; // 2371 : 253 - 0xfd
      12'h944: dout <= 8'b11111100; // 2372 : 252 - 0xfc
      12'h945: dout <= 8'b11111100; // 2373 : 252 - 0xfc
      12'h946: dout <= 8'b01111100; // 2374 : 124 - 0x7c
      12'h947: dout <= 8'b01111100; // 2375 : 124 - 0x7c
      12'h948: dout <= 8'b11110000; // 2376 : 240 - 0xf0 -- plane 1
      12'h949: dout <= 8'b11111000; // 2377 : 248 - 0xf8
      12'h94A: dout <= 8'b11111000; // 2378 : 248 - 0xf8
      12'h94B: dout <= 8'b11111100; // 2379 : 252 - 0xfc
      12'h94C: dout <= 8'b11111100; // 2380 : 252 - 0xfc
      12'h94D: dout <= 8'b11111100; // 2381 : 252 - 0xfc
      12'h94E: dout <= 8'b01111100; // 2382 : 124 - 0x7c
      12'h94F: dout <= 8'b01111100; // 2383 : 124 - 0x7c
      12'h950: dout <= 8'b11000111; // 2384 : 199 - 0xc7 -- Background 0x95
      12'h951: dout <= 8'b10001111; // 2385 : 143 - 0x8f
      12'h952: dout <= 8'b10001111; // 2386 : 143 - 0x8f
      12'h953: dout <= 8'b00011111; // 2387 :  31 - 0x1f
      12'h954: dout <= 8'b00011111; // 2388 :  31 - 0x1f
      12'h955: dout <= 8'b00111111; // 2389 :  63 - 0x3f
      12'h956: dout <= 8'b00111111; // 2390 :  63 - 0x3f
      12'h957: dout <= 8'b01111111; // 2391 : 127 - 0x7f
      12'h958: dout <= 8'b00010111; // 2392 :  23 - 0x17 -- plane 1
      12'h959: dout <= 8'b00101111; // 2393 :  47 - 0x2f
      12'h95A: dout <= 8'b00101111; // 2394 :  47 - 0x2f
      12'h95B: dout <= 8'b01011111; // 2395 :  95 - 0x5f
      12'h95C: dout <= 8'b01011111; // 2396 :  95 - 0x5f
      12'h95D: dout <= 8'b10111111; // 2397 : 191 - 0xbf
      12'h95E: dout <= 8'b10111111; // 2398 : 191 - 0xbf
      12'h95F: dout <= 8'b01111111; // 2399 : 127 - 0x7f
      12'h960: dout <= 8'b00001111; // 2400 :  15 - 0xf -- Background 0x96
      12'h961: dout <= 8'b00001111; // 2401 :  15 - 0xf
      12'h962: dout <= 8'b10000111; // 2402 : 135 - 0x87
      12'h963: dout <= 8'b10000111; // 2403 : 135 - 0x87
      12'h964: dout <= 8'b11000010; // 2404 : 194 - 0xc2
      12'h965: dout <= 8'b11000010; // 2405 : 194 - 0xc2
      12'h966: dout <= 8'b11100000; // 2406 : 224 - 0xe0
      12'h967: dout <= 8'b11100000; // 2407 : 224 - 0xe0
      12'h968: dout <= 8'b01100000; // 2408 :  96 - 0x60 -- plane 1
      12'h969: dout <= 8'b01100000; // 2409 :  96 - 0x60
      12'h96A: dout <= 8'b10110000; // 2410 : 176 - 0xb0
      12'h96B: dout <= 8'b10110000; // 2411 : 176 - 0xb0
      12'h96C: dout <= 8'b11011000; // 2412 : 216 - 0xd8
      12'h96D: dout <= 8'b11011000; // 2413 : 216 - 0xd8
      12'h96E: dout <= 8'b11101100; // 2414 : 236 - 0xec
      12'h96F: dout <= 8'b11101100; // 2415 : 236 - 0xec
      12'h970: dout <= 8'b10000011; // 2416 : 131 - 0x83 -- Background 0x97
      12'h971: dout <= 8'b10001111; // 2417 : 143 - 0x8f
      12'h972: dout <= 8'b00001111; // 2418 :  15 - 0xf
      12'h973: dout <= 8'b00011111; // 2419 :  31 - 0x1f
      12'h974: dout <= 8'b00011111; // 2420 :  31 - 0x1f
      12'h975: dout <= 8'b00111111; // 2421 :  63 - 0x3f
      12'h976: dout <= 8'b00111111; // 2422 :  63 - 0x3f
      12'h977: dout <= 8'b00111111; // 2423 :  63 - 0x3f
      12'h978: dout <= 8'b00110011; // 2424 :  51 - 0x33 -- plane 1
      12'h979: dout <= 8'b00101111; // 2425 :  47 - 0x2f
      12'h97A: dout <= 8'b01101111; // 2426 : 111 - 0x6f
      12'h97B: dout <= 8'b01011111; // 2427 :  95 - 0x5f
      12'h97C: dout <= 8'b11011111; // 2428 : 223 - 0xdf
      12'h97D: dout <= 8'b10111111; // 2429 : 191 - 0xbf
      12'h97E: dout <= 8'b10111111; // 2430 : 191 - 0xbf
      12'h97F: dout <= 8'b10111111; // 2431 : 191 - 0xbf
      12'h980: dout <= 8'b11111111; // 2432 : 255 - 0xff -- Background 0x98
      12'h981: dout <= 8'b11111111; // 2433 : 255 - 0xff
      12'h982: dout <= 8'b11111111; // 2434 : 255 - 0xff
      12'h983: dout <= 8'b11111110; // 2435 : 254 - 0xfe
      12'h984: dout <= 8'b11111001; // 2436 : 249 - 0xf9
      12'h985: dout <= 8'b11100111; // 2437 : 231 - 0xe7
      12'h986: dout <= 8'b11111100; // 2438 : 252 - 0xfc
      12'h987: dout <= 8'b11110000; // 2439 : 240 - 0xf0
      12'h988: dout <= 8'b11111111; // 2440 : 255 - 0xff -- plane 1
      12'h989: dout <= 8'b11111111; // 2441 : 255 - 0xff
      12'h98A: dout <= 8'b11111111; // 2442 : 255 - 0xff
      12'h98B: dout <= 8'b11111110; // 2443 : 254 - 0xfe
      12'h98C: dout <= 8'b11111001; // 2444 : 249 - 0xf9
      12'h98D: dout <= 8'b11100111; // 2445 : 231 - 0xe7
      12'h98E: dout <= 8'b11111100; // 2446 : 252 - 0xfc
      12'h98F: dout <= 8'b11110011; // 2447 : 243 - 0xf3
      12'h990: dout <= 8'b11110111; // 2448 : 247 - 0xf7 -- Background 0x99
      12'h991: dout <= 8'b11111011; // 2449 : 251 - 0xfb
      12'h992: dout <= 8'b11111011; // 2450 : 251 - 0xfb
      12'h993: dout <= 8'b01110011; // 2451 : 115 - 0x73
      12'h994: dout <= 8'b11000001; // 2452 : 193 - 0xc1
      12'h995: dout <= 8'b00000011; // 2453 :   3 - 0x3
      12'h996: dout <= 8'b00001111; // 2454 :  15 - 0xf
      12'h997: dout <= 8'b00111111; // 2455 :  63 - 0x3f
      12'h998: dout <= 8'b11110000; // 2456 : 240 - 0xf0 -- plane 1
      12'h999: dout <= 8'b11111000; // 2457 : 248 - 0xf8
      12'h99A: dout <= 8'b11111000; // 2458 : 248 - 0xf8
      12'h99B: dout <= 8'b01110000; // 2459 : 112 - 0x70
      12'h99C: dout <= 8'b11001100; // 2460 : 204 - 0xcc
      12'h99D: dout <= 8'b00110000; // 2461 :  48 - 0x30
      12'h99E: dout <= 8'b11000000; // 2462 : 192 - 0xc0
      12'h99F: dout <= 8'b00000000; // 2463 :   0 - 0x0
      12'h9A0: dout <= 8'b11111111; // 2464 : 255 - 0xff -- Background 0x9a
      12'h9A1: dout <= 8'b11111111; // 2465 : 255 - 0xff
      12'h9A2: dout <= 8'b11111111; // 2466 : 255 - 0xff
      12'h9A3: dout <= 8'b10000000; // 2467 : 128 - 0x80
      12'h9A4: dout <= 8'b10000000; // 2468 : 128 - 0x80
      12'h9A5: dout <= 8'b10000000; // 2469 : 128 - 0x80
      12'h9A6: dout <= 8'b10001111; // 2470 : 143 - 0x8f
      12'h9A7: dout <= 8'b10001111; // 2471 : 143 - 0x8f
      12'h9A8: dout <= 8'b00000000; // 2472 :   0 - 0x0 -- plane 1
      12'h9A9: dout <= 8'b00000000; // 2473 :   0 - 0x0
      12'h9AA: dout <= 8'b00000000; // 2474 :   0 - 0x0
      12'h9AB: dout <= 8'b00000000; // 2475 :   0 - 0x0
      12'h9AC: dout <= 8'b00111111; // 2476 :  63 - 0x3f
      12'h9AD: dout <= 8'b00100000; // 2477 :  32 - 0x20
      12'h9AE: dout <= 8'b00101111; // 2478 :  47 - 0x2f
      12'h9AF: dout <= 8'b00101111; // 2479 :  47 - 0x2f
      12'h9B0: dout <= 8'b11111111; // 2480 : 255 - 0xff -- Background 0x9b
      12'h9B1: dout <= 8'b11111111; // 2481 : 255 - 0xff
      12'h9B2: dout <= 8'b11111111; // 2482 : 255 - 0xff
      12'h9B3: dout <= 8'b00001111; // 2483 :  15 - 0xf
      12'h9B4: dout <= 8'b00001111; // 2484 :  15 - 0xf
      12'h9B5: dout <= 8'b00000111; // 2485 :   7 - 0x7
      12'h9B6: dout <= 8'b11110111; // 2486 : 247 - 0xf7
      12'h9B7: dout <= 8'b11110001; // 2487 : 241 - 0xf1
      12'h9B8: dout <= 8'b00000000; // 2488 :   0 - 0x0 -- plane 1
      12'h9B9: dout <= 8'b00000000; // 2489 :   0 - 0x0
      12'h9BA: dout <= 8'b00000000; // 2490 :   0 - 0x0
      12'h9BB: dout <= 8'b00000000; // 2491 :   0 - 0x0
      12'h9BC: dout <= 8'b11100000; // 2492 : 224 - 0xe0
      12'h9BD: dout <= 8'b00000000; // 2493 :   0 - 0x0
      12'h9BE: dout <= 8'b11110000; // 2494 : 240 - 0xf0
      12'h9BF: dout <= 8'b11110000; // 2495 : 240 - 0xf0
      12'h9C0: dout <= 8'b00011100; // 2496 :  28 - 0x1c -- Background 0x9c
      12'h9C1: dout <= 8'b00011110; // 2497 :  30 - 0x1e
      12'h9C2: dout <= 8'b00011111; // 2498 :  31 - 0x1f
      12'h9C3: dout <= 8'b00011111; // 2499 :  31 - 0x1f
      12'h9C4: dout <= 8'b00011111; // 2500 :  31 - 0x1f
      12'h9C5: dout <= 8'b00011111; // 2501 :  31 - 0x1f
      12'h9C6: dout <= 8'b00011111; // 2502 :  31 - 0x1f
      12'h9C7: dout <= 8'b00011111; // 2503 :  31 - 0x1f
      12'h9C8: dout <= 8'b01011101; // 2504 :  93 - 0x5d -- plane 1
      12'h9C9: dout <= 8'b01011110; // 2505 :  94 - 0x5e
      12'h9CA: dout <= 8'b01011111; // 2506 :  95 - 0x5f
      12'h9CB: dout <= 8'b01011111; // 2507 :  95 - 0x5f
      12'h9CC: dout <= 8'b01011111; // 2508 :  95 - 0x5f
      12'h9CD: dout <= 8'b01011111; // 2509 :  95 - 0x5f
      12'h9CE: dout <= 8'b01011111; // 2510 :  95 - 0x5f
      12'h9CF: dout <= 8'b01011111; // 2511 :  95 - 0x5f
      12'h9D0: dout <= 8'b00111110; // 2512 :  62 - 0x3e -- Background 0x9d
      12'h9D1: dout <= 8'b00011100; // 2513 :  28 - 0x1c
      12'h9D2: dout <= 8'b00001000; // 2514 :   8 - 0x8
      12'h9D3: dout <= 8'b10000000; // 2515 : 128 - 0x80
      12'h9D4: dout <= 8'b11000001; // 2516 : 193 - 0xc1
      12'h9D5: dout <= 8'b11100011; // 2517 : 227 - 0xe3
      12'h9D6: dout <= 8'b11110111; // 2518 : 247 - 0xf7
      12'h9D7: dout <= 8'b11111111; // 2519 : 255 - 0xff
      12'h9D8: dout <= 8'b10000000; // 2520 : 128 - 0x80 -- plane 1
      12'h9D9: dout <= 8'b11000001; // 2521 : 193 - 0xc1
      12'h9DA: dout <= 8'b01100011; // 2522 :  99 - 0x63
      12'h9DB: dout <= 8'b10110110; // 2523 : 182 - 0xb6
      12'h9DC: dout <= 8'b11011001; // 2524 : 217 - 0xd9
      12'h9DD: dout <= 8'b11101011; // 2525 : 235 - 0xeb
      12'h9DE: dout <= 8'b11110111; // 2526 : 247 - 0xf7
      12'h9DF: dout <= 8'b11111111; // 2527 : 255 - 0xff
      12'h9E0: dout <= 8'b00011100; // 2528 :  28 - 0x1c -- Background 0x9e
      12'h9E1: dout <= 8'b00111100; // 2529 :  60 - 0x3c
      12'h9E2: dout <= 8'b01111100; // 2530 : 124 - 0x7c
      12'h9E3: dout <= 8'b11111100; // 2531 : 252 - 0xfc
      12'h9E4: dout <= 8'b11111100; // 2532 : 252 - 0xfc
      12'h9E5: dout <= 8'b11111100; // 2533 : 252 - 0xfc
      12'h9E6: dout <= 8'b11111100; // 2534 : 252 - 0xfc
      12'h9E7: dout <= 8'b11111100; // 2535 : 252 - 0xfc
      12'h9E8: dout <= 8'b11011101; // 2536 : 221 - 0xdd -- plane 1
      12'h9E9: dout <= 8'b10111101; // 2537 : 189 - 0xbd
      12'h9EA: dout <= 8'b01111101; // 2538 : 125 - 0x7d
      12'h9EB: dout <= 8'b11111101; // 2539 : 253 - 0xfd
      12'h9EC: dout <= 8'b11111101; // 2540 : 253 - 0xfd
      12'h9ED: dout <= 8'b11111101; // 2541 : 253 - 0xfd
      12'h9EE: dout <= 8'b11111101; // 2542 : 253 - 0xfd
      12'h9EF: dout <= 8'b11111101; // 2543 : 253 - 0xfd
      12'h9F0: dout <= 8'b01111100; // 2544 : 124 - 0x7c -- Background 0x9f
      12'h9F1: dout <= 8'b01111100; // 2545 : 124 - 0x7c
      12'h9F2: dout <= 8'b01111000; // 2546 : 120 - 0x78
      12'h9F3: dout <= 8'b01111000; // 2547 : 120 - 0x78
      12'h9F4: dout <= 8'b01110001; // 2548 : 113 - 0x71
      12'h9F5: dout <= 8'b01110001; // 2549 : 113 - 0x71
      12'h9F6: dout <= 8'b01100011; // 2550 :  99 - 0x63
      12'h9F7: dout <= 8'b01100011; // 2551 :  99 - 0x63
      12'h9F8: dout <= 8'b00000001; // 2552 :   1 - 0x1 -- plane 1
      12'h9F9: dout <= 8'b00000001; // 2553 :   1 - 0x1
      12'h9FA: dout <= 8'b00000010; // 2554 :   2 - 0x2
      12'h9FB: dout <= 8'b00000010; // 2555 :   2 - 0x2
      12'h9FC: dout <= 8'b00000101; // 2556 :   5 - 0x5
      12'h9FD: dout <= 8'b00000101; // 2557 :   5 - 0x5
      12'h9FE: dout <= 8'b00001011; // 2558 :  11 - 0xb
      12'h9FF: dout <= 8'b00001011; // 2559 :  11 - 0xb
      12'hA00: dout <= 8'b01110001; // 2560 : 113 - 0x71 -- Background 0xa0
      12'hA01: dout <= 8'b01110000; // 2561 : 112 - 0x70
      12'hA02: dout <= 8'b11111000; // 2562 : 248 - 0xf8
      12'hA03: dout <= 8'b11111000; // 2563 : 248 - 0xf8
      12'hA04: dout <= 8'b11111100; // 2564 : 252 - 0xfc
      12'hA05: dout <= 8'b11111100; // 2565 : 252 - 0xfc
      12'hA06: dout <= 8'b11111110; // 2566 : 254 - 0xfe
      12'hA07: dout <= 8'b11111110; // 2567 : 254 - 0xfe
      12'hA08: dout <= 8'b01110100; // 2568 : 116 - 0x74 -- plane 1
      12'hA09: dout <= 8'b01110110; // 2569 : 118 - 0x76
      12'hA0A: dout <= 8'b11111010; // 2570 : 250 - 0xfa
      12'hA0B: dout <= 8'b11111011; // 2571 : 251 - 0xfb
      12'hA0C: dout <= 8'b11111101; // 2572 : 253 - 0xfd
      12'hA0D: dout <= 8'b11111101; // 2573 : 253 - 0xfd
      12'hA0E: dout <= 8'b11111110; // 2574 : 254 - 0xfe
      12'hA0F: dout <= 8'b11111110; // 2575 : 254 - 0xfe
      12'hA10: dout <= 8'b11111000; // 2576 : 248 - 0xf8 -- Background 0xa1
      12'hA11: dout <= 8'b11111000; // 2577 : 248 - 0xf8
      12'hA12: dout <= 8'b11111000; // 2578 : 248 - 0xf8
      12'hA13: dout <= 8'b01111000; // 2579 : 120 - 0x78
      12'hA14: dout <= 8'b01111000; // 2580 : 120 - 0x78
      12'hA15: dout <= 8'b00111000; // 2581 :  56 - 0x38
      12'hA16: dout <= 8'b00111000; // 2582 :  56 - 0x38
      12'hA17: dout <= 8'b00011000; // 2583 :  24 - 0x18
      12'hA18: dout <= 8'b00000010; // 2584 :   2 - 0x2 -- plane 1
      12'hA19: dout <= 8'b00000010; // 2585 :   2 - 0x2
      12'hA1A: dout <= 8'b00000010; // 2586 :   2 - 0x2
      12'hA1B: dout <= 8'b00000010; // 2587 :   2 - 0x2
      12'hA1C: dout <= 8'b00000010; // 2588 :   2 - 0x2
      12'hA1D: dout <= 8'b10000010; // 2589 : 130 - 0x82
      12'hA1E: dout <= 8'b10000010; // 2590 : 130 - 0x82
      12'hA1F: dout <= 8'b11000010; // 2591 : 194 - 0xc2
      12'hA20: dout <= 8'b11100000; // 2592 : 224 - 0xe0 -- Background 0xa2
      12'hA21: dout <= 8'b11110000; // 2593 : 240 - 0xf0
      12'hA22: dout <= 8'b11111000; // 2594 : 248 - 0xf8
      12'hA23: dout <= 8'b11111000; // 2595 : 248 - 0xf8
      12'hA24: dout <= 8'b11111100; // 2596 : 252 - 0xfc
      12'hA25: dout <= 8'b11111100; // 2597 : 252 - 0xfc
      12'hA26: dout <= 8'b11111110; // 2598 : 254 - 0xfe
      12'hA27: dout <= 8'b11111111; // 2599 : 255 - 0xff
      12'hA28: dout <= 8'b11101010; // 2600 : 234 - 0xea -- plane 1
      12'hA29: dout <= 8'b11110110; // 2601 : 246 - 0xf6
      12'hA2A: dout <= 8'b11111010; // 2602 : 250 - 0xfa
      12'hA2B: dout <= 8'b11111010; // 2603 : 250 - 0xfa
      12'hA2C: dout <= 8'b11111100; // 2604 : 252 - 0xfc
      12'hA2D: dout <= 8'b11111100; // 2605 : 252 - 0xfc
      12'hA2E: dout <= 8'b11111110; // 2606 : 254 - 0xfe
      12'hA2F: dout <= 8'b11111111; // 2607 : 255 - 0xff
      12'hA30: dout <= 8'b11111111; // 2608 : 255 - 0xff -- Background 0xa3
      12'hA31: dout <= 8'b11111111; // 2609 : 255 - 0xff
      12'hA32: dout <= 8'b11111111; // 2610 : 255 - 0xff
      12'hA33: dout <= 8'b11111111; // 2611 : 255 - 0xff
      12'hA34: dout <= 8'b11111111; // 2612 : 255 - 0xff
      12'hA35: dout <= 8'b11111111; // 2613 : 255 - 0xff
      12'hA36: dout <= 8'b11111111; // 2614 : 255 - 0xff
      12'hA37: dout <= 8'b11111111; // 2615 : 255 - 0xff
      12'hA38: dout <= 8'b11111111; // 2616 : 255 - 0xff -- plane 1
      12'hA39: dout <= 8'b11111111; // 2617 : 255 - 0xff
      12'hA3A: dout <= 8'b11111111; // 2618 : 255 - 0xff
      12'hA3B: dout <= 8'b11111111; // 2619 : 255 - 0xff
      12'hA3C: dout <= 8'b11111111; // 2620 : 255 - 0xff
      12'hA3D: dout <= 8'b11111111; // 2621 : 255 - 0xff
      12'hA3E: dout <= 8'b11111111; // 2622 : 255 - 0xff
      12'hA3F: dout <= 8'b11111111; // 2623 : 255 - 0xff
      12'hA40: dout <= 8'b00011111; // 2624 :  31 - 0x1f -- Background 0xa4
      12'hA41: dout <= 8'b00011111; // 2625 :  31 - 0x1f
      12'hA42: dout <= 8'b00011111; // 2626 :  31 - 0x1f
      12'hA43: dout <= 8'b00011111; // 2627 :  31 - 0x1f
      12'hA44: dout <= 8'b00011111; // 2628 :  31 - 0x1f
      12'hA45: dout <= 8'b00011111; // 2629 :  31 - 0x1f
      12'hA46: dout <= 8'b00011111; // 2630 :  31 - 0x1f
      12'hA47: dout <= 8'b00011111; // 2631 :  31 - 0x1f
      12'hA48: dout <= 8'b01000000; // 2632 :  64 - 0x40 -- plane 1
      12'hA49: dout <= 8'b01000000; // 2633 :  64 - 0x40
      12'hA4A: dout <= 8'b01000000; // 2634 :  64 - 0x40
      12'hA4B: dout <= 8'b01000000; // 2635 :  64 - 0x40
      12'hA4C: dout <= 8'b01000000; // 2636 :  64 - 0x40
      12'hA4D: dout <= 8'b01000000; // 2637 :  64 - 0x40
      12'hA4E: dout <= 8'b01000000; // 2638 :  64 - 0x40
      12'hA4F: dout <= 8'b01000000; // 2639 :  64 - 0x40
      12'hA50: dout <= 8'b11111000; // 2640 : 248 - 0xf8 -- Background 0xa5
      12'hA51: dout <= 8'b11111111; // 2641 : 255 - 0xff
      12'hA52: dout <= 8'b11111111; // 2642 : 255 - 0xff
      12'hA53: dout <= 8'b11111000; // 2643 : 248 - 0xf8
      12'hA54: dout <= 8'b11111000; // 2644 : 248 - 0xf8
      12'hA55: dout <= 8'b11111000; // 2645 : 248 - 0xf8
      12'hA56: dout <= 8'b11111000; // 2646 : 248 - 0xf8
      12'hA57: dout <= 8'b11111000; // 2647 : 248 - 0xf8
      12'hA58: dout <= 8'b11111000; // 2648 : 248 - 0xf8 -- plane 1
      12'hA59: dout <= 8'b11111111; // 2649 : 255 - 0xff
      12'hA5A: dout <= 8'b11111111; // 2650 : 255 - 0xff
      12'hA5B: dout <= 8'b11111000; // 2651 : 248 - 0xf8
      12'hA5C: dout <= 8'b11111011; // 2652 : 251 - 0xfb
      12'hA5D: dout <= 8'b11111010; // 2653 : 250 - 0xfa
      12'hA5E: dout <= 8'b11111010; // 2654 : 250 - 0xfa
      12'hA5F: dout <= 8'b11111010; // 2655 : 250 - 0xfa
      12'hA60: dout <= 8'b11111100; // 2656 : 252 - 0xfc -- Background 0xa6
      12'hA61: dout <= 8'b11111000; // 2657 : 248 - 0xf8
      12'hA62: dout <= 8'b11110000; // 2658 : 240 - 0xf0
      12'hA63: dout <= 8'b00000001; // 2659 :   1 - 0x1
      12'hA64: dout <= 8'b00000001; // 2660 :   1 - 0x1
      12'hA65: dout <= 8'b00000011; // 2661 :   3 - 0x3
      12'hA66: dout <= 8'b11000011; // 2662 : 195 - 0xc3
      12'hA67: dout <= 8'b10000111; // 2663 : 135 - 0x87
      12'hA68: dout <= 8'b11111100; // 2664 : 252 - 0xfc -- plane 1
      12'hA69: dout <= 8'b11111010; // 2665 : 250 - 0xfa
      12'hA6A: dout <= 8'b11110110; // 2666 : 246 - 0xf6
      12'hA6B: dout <= 8'b00001101; // 2667 :  13 - 0xd
      12'hA6C: dout <= 8'b11111001; // 2668 : 249 - 0xf9
      12'hA6D: dout <= 8'b00000011; // 2669 :   3 - 0x3
      12'hA6E: dout <= 8'b00010011; // 2670 :  19 - 0x13
      12'hA6F: dout <= 8'b00110111; // 2671 :  55 - 0x37
      12'hA70: dout <= 8'b01111111; // 2672 : 127 - 0x7f -- Background 0xa7
      12'hA71: dout <= 8'b11111001; // 2673 : 249 - 0xf9
      12'hA72: dout <= 8'b11111001; // 2674 : 249 - 0xf9
      12'hA73: dout <= 8'b11111111; // 2675 : 255 - 0xff
      12'hA74: dout <= 8'b11111110; // 2676 : 254 - 0xfe
      12'hA75: dout <= 8'b11111100; // 2677 : 252 - 0xfc
      12'hA76: dout <= 8'b11111111; // 2678 : 255 - 0xff
      12'hA77: dout <= 8'b11111111; // 2679 : 255 - 0xff
      12'hA78: dout <= 8'b01111111; // 2680 : 127 - 0x7f -- plane 1
      12'hA79: dout <= 8'b11111001; // 2681 : 249 - 0xf9
      12'hA7A: dout <= 8'b11111001; // 2682 : 249 - 0xf9
      12'hA7B: dout <= 8'b11111111; // 2683 : 255 - 0xff
      12'hA7C: dout <= 8'b11111110; // 2684 : 254 - 0xfe
      12'hA7D: dout <= 8'b11111100; // 2685 : 252 - 0xfc
      12'hA7E: dout <= 8'b11111111; // 2686 : 255 - 0xff
      12'hA7F: dout <= 8'b11111111; // 2687 : 255 - 0xff
      12'hA80: dout <= 8'b11110000; // 2688 : 240 - 0xf0 -- Background 0xa8
      12'hA81: dout <= 8'b11110000; // 2689 : 240 - 0xf0
      12'hA82: dout <= 8'b11111000; // 2690 : 248 - 0xf8
      12'hA83: dout <= 8'b01111000; // 2691 : 120 - 0x78
      12'hA84: dout <= 8'b11111100; // 2692 : 252 - 0xfc
      12'hA85: dout <= 8'b11110100; // 2693 : 244 - 0xf4
      12'hA86: dout <= 8'b11110110; // 2694 : 246 - 0xf6
      12'hA87: dout <= 8'b11111010; // 2695 : 250 - 0xfa
      12'hA88: dout <= 8'b11110110; // 2696 : 246 - 0xf6 -- plane 1
      12'hA89: dout <= 8'b11110110; // 2697 : 246 - 0xf6
      12'hA8A: dout <= 8'b11111011; // 2698 : 251 - 0xfb
      12'hA8B: dout <= 8'b01111011; // 2699 : 123 - 0x7b
      12'hA8C: dout <= 8'b11111101; // 2700 : 253 - 0xfd
      12'hA8D: dout <= 8'b11110101; // 2701 : 245 - 0xf5
      12'hA8E: dout <= 8'b11110110; // 2702 : 246 - 0xf6
      12'hA8F: dout <= 8'b11111010; // 2703 : 250 - 0xfa
      12'hA90: dout <= 8'b00111111; // 2704 :  63 - 0x3f -- Background 0xa9
      12'hA91: dout <= 8'b00111111; // 2705 :  63 - 0x3f
      12'hA92: dout <= 8'b00111111; // 2706 :  63 - 0x3f
      12'hA93: dout <= 8'b00111111; // 2707 :  63 - 0x3f
      12'hA94: dout <= 8'b00111111; // 2708 :  63 - 0x3f
      12'hA95: dout <= 8'b00011111; // 2709 :  31 - 0x1f
      12'hA96: dout <= 8'b00001111; // 2710 :  15 - 0xf
      12'hA97: dout <= 8'b00000111; // 2711 :   7 - 0x7
      12'hA98: dout <= 8'b10111111; // 2712 : 191 - 0xbf -- plane 1
      12'hA99: dout <= 8'b10111111; // 2713 : 191 - 0xbf
      12'hA9A: dout <= 8'b00111111; // 2714 :  63 - 0x3f
      12'hA9B: dout <= 8'b00111111; // 2715 :  63 - 0x3f
      12'hA9C: dout <= 8'b10111111; // 2716 : 191 - 0xbf
      12'hA9D: dout <= 8'b10011111; // 2717 : 159 - 0x9f
      12'hA9E: dout <= 8'b11001111; // 2718 : 207 - 0xcf
      12'hA9F: dout <= 8'b11010111; // 2719 : 215 - 0xd7
      12'hAA0: dout <= 8'b11100000; // 2720 : 224 - 0xe0 -- Background 0xaa
      12'hAA1: dout <= 8'b11111000; // 2721 : 248 - 0xf8
      12'hAA2: dout <= 8'b11111111; // 2722 : 255 - 0xff
      12'hAA3: dout <= 8'b11110011; // 2723 : 243 - 0xf3
      12'hAA4: dout <= 8'b11111100; // 2724 : 252 - 0xfc
      12'hAA5: dout <= 8'b11111111; // 2725 : 255 - 0xff
      12'hAA6: dout <= 8'b11111111; // 2726 : 255 - 0xff
      12'hAA7: dout <= 8'b11111111; // 2727 : 255 - 0xff
      12'hAA8: dout <= 8'b11100100; // 2728 : 228 - 0xe4 -- plane 1
      12'hAA9: dout <= 8'b11111000; // 2729 : 248 - 0xf8
      12'hAAA: dout <= 8'b11111111; // 2730 : 255 - 0xff
      12'hAAB: dout <= 8'b11110011; // 2731 : 243 - 0xf3
      12'hAAC: dout <= 8'b11111100; // 2732 : 252 - 0xfc
      12'hAAD: dout <= 8'b11111111; // 2733 : 255 - 0xff
      12'hAAE: dout <= 8'b11111111; // 2734 : 255 - 0xff
      12'hAAF: dout <= 8'b11111111; // 2735 : 255 - 0xff
      12'hAB0: dout <= 8'b11111111; // 2736 : 255 - 0xff -- Background 0xab
      12'hAB1: dout <= 8'b11111111; // 2737 : 255 - 0xff
      12'hAB2: dout <= 8'b00111111; // 2738 :  63 - 0x3f
      12'hAB3: dout <= 8'b11001111; // 2739 : 207 - 0xcf
      12'hAB4: dout <= 8'b11110011; // 2740 : 243 - 0xf3
      12'hAB5: dout <= 8'b00111101; // 2741 :  61 - 0x3d
      12'hAB6: dout <= 8'b11011000; // 2742 : 216 - 0xd8
      12'hAB7: dout <= 8'b10110000; // 2743 : 176 - 0xb0
      12'hAB8: dout <= 8'b00000000; // 2744 :   0 - 0x0 -- plane 1
      12'hAB9: dout <= 8'b00000000; // 2745 :   0 - 0x0
      12'hABA: dout <= 8'b00000000; // 2746 :   0 - 0x0
      12'hABB: dout <= 8'b11000000; // 2747 : 192 - 0xc0
      12'hABC: dout <= 8'b11110000; // 2748 : 240 - 0xf0
      12'hABD: dout <= 8'b00111100; // 2749 :  60 - 0x3c
      12'hABE: dout <= 8'b11011000; // 2750 : 216 - 0xd8
      12'hABF: dout <= 8'b10110110; // 2751 : 182 - 0xb6
      12'hAC0: dout <= 8'b10001111; // 2752 : 143 - 0x8f -- Background 0xac
      12'hAC1: dout <= 8'b11101111; // 2753 : 239 - 0xef
      12'hAC2: dout <= 8'b11100000; // 2754 : 224 - 0xe0
      12'hAC3: dout <= 8'b11111000; // 2755 : 248 - 0xf8
      12'hAC4: dout <= 8'b11111000; // 2756 : 248 - 0xf8
      12'hAC5: dout <= 8'b11111111; // 2757 : 255 - 0xff
      12'hAC6: dout <= 8'b11111111; // 2758 : 255 - 0xff
      12'hAC7: dout <= 8'b11111111; // 2759 : 255 - 0xff
      12'hAC8: dout <= 8'b00001111; // 2760 :  15 - 0xf -- plane 1
      12'hAC9: dout <= 8'b00001111; // 2761 :  15 - 0xf
      12'hACA: dout <= 8'b00000000; // 2762 :   0 - 0x0
      12'hACB: dout <= 8'b00000011; // 2763 :   3 - 0x3
      12'hACC: dout <= 8'b00000000; // 2764 :   0 - 0x0
      12'hACD: dout <= 8'b00000000; // 2765 :   0 - 0x0
      12'hACE: dout <= 8'b00000000; // 2766 :   0 - 0x0
      12'hACF: dout <= 8'b00000000; // 2767 :   0 - 0x0
      12'hAD0: dout <= 8'b11110001; // 2768 : 241 - 0xf1 -- Background 0xad
      12'hAD1: dout <= 8'b11110001; // 2769 : 241 - 0xf1
      12'hAD2: dout <= 8'b00000001; // 2770 :   1 - 0x1
      12'hAD3: dout <= 8'b00000001; // 2771 :   1 - 0x1
      12'hAD4: dout <= 8'b00000001; // 2772 :   1 - 0x1
      12'hAD5: dout <= 8'b11111111; // 2773 : 255 - 0xff
      12'hAD6: dout <= 8'b11111111; // 2774 : 255 - 0xff
      12'hAD7: dout <= 8'b11111111; // 2775 : 255 - 0xff
      12'hAD8: dout <= 8'b11110100; // 2776 : 244 - 0xf4 -- plane 1
      12'hAD9: dout <= 8'b11110100; // 2777 : 244 - 0xf4
      12'hADA: dout <= 8'b00000100; // 2778 :   4 - 0x4
      12'hADB: dout <= 8'b11111100; // 2779 : 252 - 0xfc
      12'hADC: dout <= 8'b00000000; // 2780 :   0 - 0x0
      12'hADD: dout <= 8'b00000000; // 2781 :   0 - 0x0
      12'hADE: dout <= 8'b00000000; // 2782 :   0 - 0x0
      12'hADF: dout <= 8'b00000000; // 2783 :   0 - 0x0
      12'hAE0: dout <= 8'b00011111; // 2784 :  31 - 0x1f -- Background 0xae
      12'hAE1: dout <= 8'b00011111; // 2785 :  31 - 0x1f
      12'hAE2: dout <= 8'b00011111; // 2786 :  31 - 0x1f
      12'hAE3: dout <= 8'b00011111; // 2787 :  31 - 0x1f
      12'hAE4: dout <= 8'b00011111; // 2788 :  31 - 0x1f
      12'hAE5: dout <= 8'b00011111; // 2789 :  31 - 0x1f
      12'hAE6: dout <= 8'b00011111; // 2790 :  31 - 0x1f
      12'hAE7: dout <= 8'b00011111; // 2791 :  31 - 0x1f
      12'hAE8: dout <= 8'b01011111; // 2792 :  95 - 0x5f -- plane 1
      12'hAE9: dout <= 8'b01011111; // 2793 :  95 - 0x5f
      12'hAEA: dout <= 8'b01011111; // 2794 :  95 - 0x5f
      12'hAEB: dout <= 8'b01011111; // 2795 :  95 - 0x5f
      12'hAEC: dout <= 8'b01011111; // 2796 :  95 - 0x5f
      12'hAED: dout <= 8'b01011111; // 2797 :  95 - 0x5f
      12'hAEE: dout <= 8'b01011111; // 2798 :  95 - 0x5f
      12'hAEF: dout <= 8'b01011111; // 2799 :  95 - 0x5f
      12'hAF0: dout <= 8'b11111100; // 2800 : 252 - 0xfc -- Background 0xaf
      12'hAF1: dout <= 8'b11111100; // 2801 : 252 - 0xfc
      12'hAF2: dout <= 8'b11111100; // 2802 : 252 - 0xfc
      12'hAF3: dout <= 8'b11111100; // 2803 : 252 - 0xfc
      12'hAF4: dout <= 8'b11110100; // 2804 : 244 - 0xf4
      12'hAF5: dout <= 8'b11110100; // 2805 : 244 - 0xf4
      12'hAF6: dout <= 8'b11110100; // 2806 : 244 - 0xf4
      12'hAF7: dout <= 8'b11110100; // 2807 : 244 - 0xf4
      12'hAF8: dout <= 8'b11111101; // 2808 : 253 - 0xfd -- plane 1
      12'hAF9: dout <= 8'b11111101; // 2809 : 253 - 0xfd
      12'hAFA: dout <= 8'b11111101; // 2810 : 253 - 0xfd
      12'hAFB: dout <= 8'b11111101; // 2811 : 253 - 0xfd
      12'hAFC: dout <= 8'b11110101; // 2812 : 245 - 0xf5
      12'hAFD: dout <= 8'b11110101; // 2813 : 245 - 0xf5
      12'hAFE: dout <= 8'b11110101; // 2814 : 245 - 0xf5
      12'hAFF: dout <= 8'b11110101; // 2815 : 245 - 0xf5
      12'hB00: dout <= 8'b00001100; // 2816 :  12 - 0xc -- Background 0xb0
      12'hB01: dout <= 8'b00011100; // 2817 :  28 - 0x1c
      12'hB02: dout <= 8'b00001100; // 2818 :  12 - 0xc
      12'hB03: dout <= 8'b00001100; // 2819 :  12 - 0xc
      12'hB04: dout <= 8'b00001100; // 2820 :  12 - 0xc
      12'hB05: dout <= 8'b00001100; // 2821 :  12 - 0xc
      12'hB06: dout <= 8'b00111111; // 2822 :  63 - 0x3f
      12'hB07: dout <= 8'b00000000; // 2823 :   0 - 0x0
      12'hB08: dout <= 8'b00001100; // 2824 :  12 - 0xc -- plane 1
      12'hB09: dout <= 8'b00011100; // 2825 :  28 - 0x1c
      12'hB0A: dout <= 8'b00001100; // 2826 :  12 - 0xc
      12'hB0B: dout <= 8'b00001100; // 2827 :  12 - 0xc
      12'hB0C: dout <= 8'b00001100; // 2828 :  12 - 0xc
      12'hB0D: dout <= 8'b00001100; // 2829 :  12 - 0xc
      12'hB0E: dout <= 8'b00111111; // 2830 :  63 - 0x3f
      12'hB0F: dout <= 8'b00000000; // 2831 :   0 - 0x0
      12'hB10: dout <= 8'b00111110; // 2832 :  62 - 0x3e -- Background 0xb1
      12'hB11: dout <= 8'b01100011; // 2833 :  99 - 0x63
      12'hB12: dout <= 8'b00000111; // 2834 :   7 - 0x7
      12'hB13: dout <= 8'b00011110; // 2835 :  30 - 0x1e
      12'hB14: dout <= 8'b00111100; // 2836 :  60 - 0x3c
      12'hB15: dout <= 8'b01110000; // 2837 : 112 - 0x70
      12'hB16: dout <= 8'b01111111; // 2838 : 127 - 0x7f
      12'hB17: dout <= 8'b00000000; // 2839 :   0 - 0x0
      12'hB18: dout <= 8'b00111110; // 2840 :  62 - 0x3e -- plane 1
      12'hB19: dout <= 8'b01100011; // 2841 :  99 - 0x63
      12'hB1A: dout <= 8'b00000111; // 2842 :   7 - 0x7
      12'hB1B: dout <= 8'b00011110; // 2843 :  30 - 0x1e
      12'hB1C: dout <= 8'b00111100; // 2844 :  60 - 0x3c
      12'hB1D: dout <= 8'b01110000; // 2845 : 112 - 0x70
      12'hB1E: dout <= 8'b01111111; // 2846 : 127 - 0x7f
      12'hB1F: dout <= 8'b00000000; // 2847 :   0 - 0x0
      12'hB20: dout <= 8'b01111110; // 2848 : 126 - 0x7e -- Background 0xb2
      12'hB21: dout <= 8'b01100011; // 2849 :  99 - 0x63
      12'hB22: dout <= 8'b01100011; // 2850 :  99 - 0x63
      12'hB23: dout <= 8'b01100011; // 2851 :  99 - 0x63
      12'hB24: dout <= 8'b01111110; // 2852 : 126 - 0x7e
      12'hB25: dout <= 8'b01100000; // 2853 :  96 - 0x60
      12'hB26: dout <= 8'b01100000; // 2854 :  96 - 0x60
      12'hB27: dout <= 8'b00000000; // 2855 :   0 - 0x0
      12'hB28: dout <= 8'b01111110; // 2856 : 126 - 0x7e -- plane 1
      12'hB29: dout <= 8'b01100011; // 2857 :  99 - 0x63
      12'hB2A: dout <= 8'b01100011; // 2858 :  99 - 0x63
      12'hB2B: dout <= 8'b01100011; // 2859 :  99 - 0x63
      12'hB2C: dout <= 8'b01111110; // 2860 : 126 - 0x7e
      12'hB2D: dout <= 8'b01100000; // 2861 :  96 - 0x60
      12'hB2E: dout <= 8'b01100000; // 2862 :  96 - 0x60
      12'hB2F: dout <= 8'b00000000; // 2863 :   0 - 0x0
      12'hB30: dout <= 8'b01100011; // 2864 :  99 - 0x63 -- Background 0xb3
      12'hB31: dout <= 8'b01100011; // 2865 :  99 - 0x63
      12'hB32: dout <= 8'b01100011; // 2866 :  99 - 0x63
      12'hB33: dout <= 8'b01100011; // 2867 :  99 - 0x63
      12'hB34: dout <= 8'b01100011; // 2868 :  99 - 0x63
      12'hB35: dout <= 8'b01100011; // 2869 :  99 - 0x63
      12'hB36: dout <= 8'b00111110; // 2870 :  62 - 0x3e
      12'hB37: dout <= 8'b00000000; // 2871 :   0 - 0x0
      12'hB38: dout <= 8'b01100011; // 2872 :  99 - 0x63 -- plane 1
      12'hB39: dout <= 8'b01100011; // 2873 :  99 - 0x63
      12'hB3A: dout <= 8'b01100011; // 2874 :  99 - 0x63
      12'hB3B: dout <= 8'b01100011; // 2875 :  99 - 0x63
      12'hB3C: dout <= 8'b01100011; // 2876 :  99 - 0x63
      12'hB3D: dout <= 8'b01100011; // 2877 :  99 - 0x63
      12'hB3E: dout <= 8'b00111110; // 2878 :  62 - 0x3e
      12'hB3F: dout <= 8'b00000000; // 2879 :   0 - 0x0
      12'hB40: dout <= 8'b01100011; // 2880 :  99 - 0x63 -- Background 0xb4
      12'hB41: dout <= 8'b01100011; // 2881 :  99 - 0x63
      12'hB42: dout <= 8'b01100011; // 2882 :  99 - 0x63
      12'hB43: dout <= 8'b01111111; // 2883 : 127 - 0x7f
      12'hB44: dout <= 8'b01100011; // 2884 :  99 - 0x63
      12'hB45: dout <= 8'b01100011; // 2885 :  99 - 0x63
      12'hB46: dout <= 8'b01100011; // 2886 :  99 - 0x63
      12'hB47: dout <= 8'b00000000; // 2887 :   0 - 0x0
      12'hB48: dout <= 8'b01100011; // 2888 :  99 - 0x63 -- plane 1
      12'hB49: dout <= 8'b01100011; // 2889 :  99 - 0x63
      12'hB4A: dout <= 8'b01100011; // 2890 :  99 - 0x63
      12'hB4B: dout <= 8'b01111111; // 2891 : 127 - 0x7f
      12'hB4C: dout <= 8'b01100011; // 2892 :  99 - 0x63
      12'hB4D: dout <= 8'b01100011; // 2893 :  99 - 0x63
      12'hB4E: dout <= 8'b01100011; // 2894 :  99 - 0x63
      12'hB4F: dout <= 8'b00000000; // 2895 :   0 - 0x0
      12'hB50: dout <= 8'b00111111; // 2896 :  63 - 0x3f -- Background 0xb5
      12'hB51: dout <= 8'b00001100; // 2897 :  12 - 0xc
      12'hB52: dout <= 8'b00001100; // 2898 :  12 - 0xc
      12'hB53: dout <= 8'b00001100; // 2899 :  12 - 0xc
      12'hB54: dout <= 8'b00001100; // 2900 :  12 - 0xc
      12'hB55: dout <= 8'b00001100; // 2901 :  12 - 0xc
      12'hB56: dout <= 8'b00111111; // 2902 :  63 - 0x3f
      12'hB57: dout <= 8'b00000000; // 2903 :   0 - 0x0
      12'hB58: dout <= 8'b00111111; // 2904 :  63 - 0x3f -- plane 1
      12'hB59: dout <= 8'b00001100; // 2905 :  12 - 0xc
      12'hB5A: dout <= 8'b00001100; // 2906 :  12 - 0xc
      12'hB5B: dout <= 8'b00001100; // 2907 :  12 - 0xc
      12'hB5C: dout <= 8'b00001100; // 2908 :  12 - 0xc
      12'hB5D: dout <= 8'b00001100; // 2909 :  12 - 0xc
      12'hB5E: dout <= 8'b00111111; // 2910 :  63 - 0x3f
      12'hB5F: dout <= 8'b00000000; // 2911 :   0 - 0x0
      12'hB60: dout <= 8'b00000000; // 2912 :   0 - 0x0 -- Background 0xb6
      12'hB61: dout <= 8'b00000000; // 2913 :   0 - 0x0
      12'hB62: dout <= 8'b00000000; // 2914 :   0 - 0x0
      12'hB63: dout <= 8'b01111110; // 2915 : 126 - 0x7e
      12'hB64: dout <= 8'b00000000; // 2916 :   0 - 0x0
      12'hB65: dout <= 8'b00000000; // 2917 :   0 - 0x0
      12'hB66: dout <= 8'b00000000; // 2918 :   0 - 0x0
      12'hB67: dout <= 8'b00000000; // 2919 :   0 - 0x0
      12'hB68: dout <= 8'b00000000; // 2920 :   0 - 0x0 -- plane 1
      12'hB69: dout <= 8'b00000000; // 2921 :   0 - 0x0
      12'hB6A: dout <= 8'b00000000; // 2922 :   0 - 0x0
      12'hB6B: dout <= 8'b01111110; // 2923 : 126 - 0x7e
      12'hB6C: dout <= 8'b00000000; // 2924 :   0 - 0x0
      12'hB6D: dout <= 8'b00000000; // 2925 :   0 - 0x0
      12'hB6E: dout <= 8'b00000000; // 2926 :   0 - 0x0
      12'hB6F: dout <= 8'b00000000; // 2927 :   0 - 0x0
      12'hB70: dout <= 8'b00111100; // 2928 :  60 - 0x3c -- Background 0xb7
      12'hB71: dout <= 8'b01100110; // 2929 : 102 - 0x66
      12'hB72: dout <= 8'b01100000; // 2930 :  96 - 0x60
      12'hB73: dout <= 8'b00111110; // 2931 :  62 - 0x3e
      12'hB74: dout <= 8'b00000011; // 2932 :   3 - 0x3
      12'hB75: dout <= 8'b01100011; // 2933 :  99 - 0x63
      12'hB76: dout <= 8'b00111110; // 2934 :  62 - 0x3e
      12'hB77: dout <= 8'b00000000; // 2935 :   0 - 0x0
      12'hB78: dout <= 8'b00111100; // 2936 :  60 - 0x3c -- plane 1
      12'hB79: dout <= 8'b01100110; // 2937 : 102 - 0x66
      12'hB7A: dout <= 8'b01100000; // 2938 :  96 - 0x60
      12'hB7B: dout <= 8'b00111110; // 2939 :  62 - 0x3e
      12'hB7C: dout <= 8'b00000011; // 2940 :   3 - 0x3
      12'hB7D: dout <= 8'b01100011; // 2941 :  99 - 0x63
      12'hB7E: dout <= 8'b00111110; // 2942 :  62 - 0x3e
      12'hB7F: dout <= 8'b00000000; // 2943 :   0 - 0x0
      12'hB80: dout <= 8'b00011110; // 2944 :  30 - 0x1e -- Background 0xb8
      12'hB81: dout <= 8'b00110011; // 2945 :  51 - 0x33
      12'hB82: dout <= 8'b01100000; // 2946 :  96 - 0x60
      12'hB83: dout <= 8'b01100000; // 2947 :  96 - 0x60
      12'hB84: dout <= 8'b01100000; // 2948 :  96 - 0x60
      12'hB85: dout <= 8'b00110011; // 2949 :  51 - 0x33
      12'hB86: dout <= 8'b00011110; // 2950 :  30 - 0x1e
      12'hB87: dout <= 8'b00000000; // 2951 :   0 - 0x0
      12'hB88: dout <= 8'b00011110; // 2952 :  30 - 0x1e -- plane 1
      12'hB89: dout <= 8'b00110011; // 2953 :  51 - 0x33
      12'hB8A: dout <= 8'b01100000; // 2954 :  96 - 0x60
      12'hB8B: dout <= 8'b01100000; // 2955 :  96 - 0x60
      12'hB8C: dout <= 8'b01100000; // 2956 :  96 - 0x60
      12'hB8D: dout <= 8'b00110011; // 2957 :  51 - 0x33
      12'hB8E: dout <= 8'b00011110; // 2958 :  30 - 0x1e
      12'hB8F: dout <= 8'b00000000; // 2959 :   0 - 0x0
      12'hB90: dout <= 8'b00111110; // 2960 :  62 - 0x3e -- Background 0xb9
      12'hB91: dout <= 8'b01100011; // 2961 :  99 - 0x63
      12'hB92: dout <= 8'b01100011; // 2962 :  99 - 0x63
      12'hB93: dout <= 8'b01100011; // 2963 :  99 - 0x63
      12'hB94: dout <= 8'b01100011; // 2964 :  99 - 0x63
      12'hB95: dout <= 8'b01100011; // 2965 :  99 - 0x63
      12'hB96: dout <= 8'b00111110; // 2966 :  62 - 0x3e
      12'hB97: dout <= 8'b00000000; // 2967 :   0 - 0x0
      12'hB98: dout <= 8'b00111110; // 2968 :  62 - 0x3e -- plane 1
      12'hB99: dout <= 8'b01100011; // 2969 :  99 - 0x63
      12'hB9A: dout <= 8'b01100011; // 2970 :  99 - 0x63
      12'hB9B: dout <= 8'b01100011; // 2971 :  99 - 0x63
      12'hB9C: dout <= 8'b01100011; // 2972 :  99 - 0x63
      12'hB9D: dout <= 8'b01100011; // 2973 :  99 - 0x63
      12'hB9E: dout <= 8'b00111110; // 2974 :  62 - 0x3e
      12'hB9F: dout <= 8'b00000000; // 2975 :   0 - 0x0
      12'hBA0: dout <= 8'b01111110; // 2976 : 126 - 0x7e -- Background 0xba
      12'hBA1: dout <= 8'b01100011; // 2977 :  99 - 0x63
      12'hBA2: dout <= 8'b01100011; // 2978 :  99 - 0x63
      12'hBA3: dout <= 8'b01100111; // 2979 : 103 - 0x67
      12'hBA4: dout <= 8'b01111100; // 2980 : 124 - 0x7c
      12'hBA5: dout <= 8'b01101110; // 2981 : 110 - 0x6e
      12'hBA6: dout <= 8'b01100111; // 2982 : 103 - 0x67
      12'hBA7: dout <= 8'b00000000; // 2983 :   0 - 0x0
      12'hBA8: dout <= 8'b01111110; // 2984 : 126 - 0x7e -- plane 1
      12'hBA9: dout <= 8'b01100011; // 2985 :  99 - 0x63
      12'hBAA: dout <= 8'b01100011; // 2986 :  99 - 0x63
      12'hBAB: dout <= 8'b01100111; // 2987 : 103 - 0x67
      12'hBAC: dout <= 8'b01111100; // 2988 : 124 - 0x7c
      12'hBAD: dout <= 8'b01101110; // 2989 : 110 - 0x6e
      12'hBAE: dout <= 8'b01100111; // 2990 : 103 - 0x67
      12'hBAF: dout <= 8'b00000000; // 2991 :   0 - 0x0
      12'hBB0: dout <= 8'b01111111; // 2992 : 127 - 0x7f -- Background 0xbb
      12'hBB1: dout <= 8'b01100000; // 2993 :  96 - 0x60
      12'hBB2: dout <= 8'b01100000; // 2994 :  96 - 0x60
      12'hBB3: dout <= 8'b01111110; // 2995 : 126 - 0x7e
      12'hBB4: dout <= 8'b01100000; // 2996 :  96 - 0x60
      12'hBB5: dout <= 8'b01100000; // 2997 :  96 - 0x60
      12'hBB6: dout <= 8'b01111111; // 2998 : 127 - 0x7f
      12'hBB7: dout <= 8'b00000000; // 2999 :   0 - 0x0
      12'hBB8: dout <= 8'b01111111; // 3000 : 127 - 0x7f -- plane 1
      12'hBB9: dout <= 8'b01100000; // 3001 :  96 - 0x60
      12'hBBA: dout <= 8'b01100000; // 3002 :  96 - 0x60
      12'hBBB: dout <= 8'b01111110; // 3003 : 126 - 0x7e
      12'hBBC: dout <= 8'b01100000; // 3004 :  96 - 0x60
      12'hBBD: dout <= 8'b01100000; // 3005 :  96 - 0x60
      12'hBBE: dout <= 8'b01111111; // 3006 : 127 - 0x7f
      12'hBBF: dout <= 8'b00000000; // 3007 :   0 - 0x0
      12'hBC0: dout <= 8'b00000000; // 3008 :   0 - 0x0 -- Background 0xbc
      12'hBC1: dout <= 8'b00100010; // 3009 :  34 - 0x22
      12'hBC2: dout <= 8'b01100101; // 3010 : 101 - 0x65
      12'hBC3: dout <= 8'b00100101; // 3011 :  37 - 0x25
      12'hBC4: dout <= 8'b00100101; // 3012 :  37 - 0x25
      12'hBC5: dout <= 8'b01110010; // 3013 : 114 - 0x72
      12'hBC6: dout <= 8'b00000000; // 3014 :   0 - 0x0
      12'hBC7: dout <= 8'b00000000; // 3015 :   0 - 0x0
      12'hBC8: dout <= 8'b00000000; // 3016 :   0 - 0x0 -- plane 1
      12'hBC9: dout <= 8'b00000000; // 3017 :   0 - 0x0
      12'hBCA: dout <= 8'b00000000; // 3018 :   0 - 0x0
      12'hBCB: dout <= 8'b00000000; // 3019 :   0 - 0x0
      12'hBCC: dout <= 8'b00000000; // 3020 :   0 - 0x0
      12'hBCD: dout <= 8'b00000000; // 3021 :   0 - 0x0
      12'hBCE: dout <= 8'b00000000; // 3022 :   0 - 0x0
      12'hBCF: dout <= 8'b00000000; // 3023 :   0 - 0x0
      12'hBD0: dout <= 8'b00000000; // 3024 :   0 - 0x0 -- Background 0xbd
      12'hBD1: dout <= 8'b01110010; // 3025 : 114 - 0x72
      12'hBD2: dout <= 8'b01000101; // 3026 :  69 - 0x45
      12'hBD3: dout <= 8'b01100101; // 3027 : 101 - 0x65
      12'hBD4: dout <= 8'b00010101; // 3028 :  21 - 0x15
      12'hBD5: dout <= 8'b01100010; // 3029 :  98 - 0x62
      12'hBD6: dout <= 8'b00000000; // 3030 :   0 - 0x0
      12'hBD7: dout <= 8'b00000000; // 3031 :   0 - 0x0
      12'hBD8: dout <= 8'b00000000; // 3032 :   0 - 0x0 -- plane 1
      12'hBD9: dout <= 8'b00000000; // 3033 :   0 - 0x0
      12'hBDA: dout <= 8'b00000000; // 3034 :   0 - 0x0
      12'hBDB: dout <= 8'b00000000; // 3035 :   0 - 0x0
      12'hBDC: dout <= 8'b00000000; // 3036 :   0 - 0x0
      12'hBDD: dout <= 8'b00000000; // 3037 :   0 - 0x0
      12'hBDE: dout <= 8'b00000000; // 3038 :   0 - 0x0
      12'hBDF: dout <= 8'b00000000; // 3039 :   0 - 0x0
      12'hBE0: dout <= 8'b00000000; // 3040 :   0 - 0x0 -- Background 0xbe
      12'hBE1: dout <= 8'b01100111; // 3041 : 103 - 0x67
      12'hBE2: dout <= 8'b01010010; // 3042 :  82 - 0x52
      12'hBE3: dout <= 8'b01100010; // 3043 :  98 - 0x62
      12'hBE4: dout <= 8'b01000010; // 3044 :  66 - 0x42
      12'hBE5: dout <= 8'b01000010; // 3045 :  66 - 0x42
      12'hBE6: dout <= 8'b00000000; // 3046 :   0 - 0x0
      12'hBE7: dout <= 8'b00000000; // 3047 :   0 - 0x0
      12'hBE8: dout <= 8'b00000000; // 3048 :   0 - 0x0 -- plane 1
      12'hBE9: dout <= 8'b00000000; // 3049 :   0 - 0x0
      12'hBEA: dout <= 8'b00000000; // 3050 :   0 - 0x0
      12'hBEB: dout <= 8'b00000000; // 3051 :   0 - 0x0
      12'hBEC: dout <= 8'b00000000; // 3052 :   0 - 0x0
      12'hBED: dout <= 8'b00000000; // 3053 :   0 - 0x0
      12'hBEE: dout <= 8'b00000000; // 3054 :   0 - 0x0
      12'hBEF: dout <= 8'b00000000; // 3055 :   0 - 0x0
      12'hBF0: dout <= 8'b00000000; // 3056 :   0 - 0x0 -- Background 0xbf
      12'hBF1: dout <= 8'b01100000; // 3057 :  96 - 0x60
      12'hBF2: dout <= 8'b10000000; // 3058 : 128 - 0x80
      12'hBF3: dout <= 8'b01000000; // 3059 :  64 - 0x40
      12'hBF4: dout <= 8'b00100000; // 3060 :  32 - 0x20
      12'hBF5: dout <= 8'b11000110; // 3061 : 198 - 0xc6
      12'hBF6: dout <= 8'b00000000; // 3062 :   0 - 0x0
      12'hBF7: dout <= 8'b00000000; // 3063 :   0 - 0x0
      12'hBF8: dout <= 8'b00000000; // 3064 :   0 - 0x0 -- plane 1
      12'hBF9: dout <= 8'b00000000; // 3065 :   0 - 0x0
      12'hBFA: dout <= 8'b00000000; // 3066 :   0 - 0x0
      12'hBFB: dout <= 8'b00000000; // 3067 :   0 - 0x0
      12'hBFC: dout <= 8'b00000000; // 3068 :   0 - 0x0
      12'hBFD: dout <= 8'b00000000; // 3069 :   0 - 0x0
      12'hBFE: dout <= 8'b00000000; // 3070 :   0 - 0x0
      12'hBFF: dout <= 8'b00000000; // 3071 :   0 - 0x0
      12'hC00: dout <= 8'b01100011; // 3072 :  99 - 0x63 -- Background 0xc0
      12'hC01: dout <= 8'b01100110; // 3073 : 102 - 0x66
      12'hC02: dout <= 8'b01101100; // 3074 : 108 - 0x6c
      12'hC03: dout <= 8'b01111000; // 3075 : 120 - 0x78
      12'hC04: dout <= 8'b01111100; // 3076 : 124 - 0x7c
      12'hC05: dout <= 8'b01100110; // 3077 : 102 - 0x66
      12'hC06: dout <= 8'b01100011; // 3078 :  99 - 0x63
      12'hC07: dout <= 8'b00000000; // 3079 :   0 - 0x0
      12'hC08: dout <= 8'b01100011; // 3080 :  99 - 0x63 -- plane 1
      12'hC09: dout <= 8'b01100110; // 3081 : 102 - 0x66
      12'hC0A: dout <= 8'b01101100; // 3082 : 108 - 0x6c
      12'hC0B: dout <= 8'b01111000; // 3083 : 120 - 0x78
      12'hC0C: dout <= 8'b01111100; // 3084 : 124 - 0x7c
      12'hC0D: dout <= 8'b01100110; // 3085 : 102 - 0x66
      12'hC0E: dout <= 8'b01100011; // 3086 :  99 - 0x63
      12'hC0F: dout <= 8'b00000000; // 3087 :   0 - 0x0
      12'hC10: dout <= 8'b00111111; // 3088 :  63 - 0x3f -- Background 0xc1
      12'hC11: dout <= 8'b00001100; // 3089 :  12 - 0xc
      12'hC12: dout <= 8'b00001100; // 3090 :  12 - 0xc
      12'hC13: dout <= 8'b00001100; // 3091 :  12 - 0xc
      12'hC14: dout <= 8'b00001100; // 3092 :  12 - 0xc
      12'hC15: dout <= 8'b00001100; // 3093 :  12 - 0xc
      12'hC16: dout <= 8'b00111111; // 3094 :  63 - 0x3f
      12'hC17: dout <= 8'b00000000; // 3095 :   0 - 0x0
      12'hC18: dout <= 8'b00111111; // 3096 :  63 - 0x3f -- plane 1
      12'hC19: dout <= 8'b00001100; // 3097 :  12 - 0xc
      12'hC1A: dout <= 8'b00001100; // 3098 :  12 - 0xc
      12'hC1B: dout <= 8'b00001100; // 3099 :  12 - 0xc
      12'hC1C: dout <= 8'b00001100; // 3100 :  12 - 0xc
      12'hC1D: dout <= 8'b00001100; // 3101 :  12 - 0xc
      12'hC1E: dout <= 8'b00111111; // 3102 :  63 - 0x3f
      12'hC1F: dout <= 8'b00000000; // 3103 :   0 - 0x0
      12'hC20: dout <= 8'b01100011; // 3104 :  99 - 0x63 -- Background 0xc2
      12'hC21: dout <= 8'b01110111; // 3105 : 119 - 0x77
      12'hC22: dout <= 8'b01111111; // 3106 : 127 - 0x7f
      12'hC23: dout <= 8'b01111111; // 3107 : 127 - 0x7f
      12'hC24: dout <= 8'b01101011; // 3108 : 107 - 0x6b
      12'hC25: dout <= 8'b01100011; // 3109 :  99 - 0x63
      12'hC26: dout <= 8'b01100011; // 3110 :  99 - 0x63
      12'hC27: dout <= 8'b00000000; // 3111 :   0 - 0x0
      12'hC28: dout <= 8'b01100011; // 3112 :  99 - 0x63 -- plane 1
      12'hC29: dout <= 8'b01110111; // 3113 : 119 - 0x77
      12'hC2A: dout <= 8'b01111111; // 3114 : 127 - 0x7f
      12'hC2B: dout <= 8'b01111111; // 3115 : 127 - 0x7f
      12'hC2C: dout <= 8'b01101011; // 3116 : 107 - 0x6b
      12'hC2D: dout <= 8'b01100011; // 3117 :  99 - 0x63
      12'hC2E: dout <= 8'b01100011; // 3118 :  99 - 0x63
      12'hC2F: dout <= 8'b00000000; // 3119 :   0 - 0x0
      12'hC30: dout <= 8'b00011100; // 3120 :  28 - 0x1c -- Background 0xc3
      12'hC31: dout <= 8'b00110110; // 3121 :  54 - 0x36
      12'hC32: dout <= 8'b01100011; // 3122 :  99 - 0x63
      12'hC33: dout <= 8'b01100011; // 3123 :  99 - 0x63
      12'hC34: dout <= 8'b01111111; // 3124 : 127 - 0x7f
      12'hC35: dout <= 8'b01100011; // 3125 :  99 - 0x63
      12'hC36: dout <= 8'b01100011; // 3126 :  99 - 0x63
      12'hC37: dout <= 8'b00000000; // 3127 :   0 - 0x0
      12'hC38: dout <= 8'b00011100; // 3128 :  28 - 0x1c -- plane 1
      12'hC39: dout <= 8'b00110110; // 3129 :  54 - 0x36
      12'hC3A: dout <= 8'b01100011; // 3130 :  99 - 0x63
      12'hC3B: dout <= 8'b01100011; // 3131 :  99 - 0x63
      12'hC3C: dout <= 8'b01111111; // 3132 : 127 - 0x7f
      12'hC3D: dout <= 8'b01100011; // 3133 :  99 - 0x63
      12'hC3E: dout <= 8'b01100011; // 3134 :  99 - 0x63
      12'hC3F: dout <= 8'b00000000; // 3135 :   0 - 0x0
      12'hC40: dout <= 8'b00011111; // 3136 :  31 - 0x1f -- Background 0xc4
      12'hC41: dout <= 8'b00110000; // 3137 :  48 - 0x30
      12'hC42: dout <= 8'b01100000; // 3138 :  96 - 0x60
      12'hC43: dout <= 8'b01100111; // 3139 : 103 - 0x67
      12'hC44: dout <= 8'b01100011; // 3140 :  99 - 0x63
      12'hC45: dout <= 8'b00110011; // 3141 :  51 - 0x33
      12'hC46: dout <= 8'b00011111; // 3142 :  31 - 0x1f
      12'hC47: dout <= 8'b00000000; // 3143 :   0 - 0x0
      12'hC48: dout <= 8'b00011111; // 3144 :  31 - 0x1f -- plane 1
      12'hC49: dout <= 8'b00110000; // 3145 :  48 - 0x30
      12'hC4A: dout <= 8'b01100000; // 3146 :  96 - 0x60
      12'hC4B: dout <= 8'b01100111; // 3147 : 103 - 0x67
      12'hC4C: dout <= 8'b01100011; // 3148 :  99 - 0x63
      12'hC4D: dout <= 8'b00110011; // 3149 :  51 - 0x33
      12'hC4E: dout <= 8'b00011111; // 3150 :  31 - 0x1f
      12'hC4F: dout <= 8'b00000000; // 3151 :   0 - 0x0
      12'hC50: dout <= 8'b01100011; // 3152 :  99 - 0x63 -- Background 0xc5
      12'hC51: dout <= 8'b01100011; // 3153 :  99 - 0x63
      12'hC52: dout <= 8'b01100011; // 3154 :  99 - 0x63
      12'hC53: dout <= 8'b01100011; // 3155 :  99 - 0x63
      12'hC54: dout <= 8'b01100011; // 3156 :  99 - 0x63
      12'hC55: dout <= 8'b01100011; // 3157 :  99 - 0x63
      12'hC56: dout <= 8'b00111110; // 3158 :  62 - 0x3e
      12'hC57: dout <= 8'b00000000; // 3159 :   0 - 0x0
      12'hC58: dout <= 8'b01100011; // 3160 :  99 - 0x63 -- plane 1
      12'hC59: dout <= 8'b01100011; // 3161 :  99 - 0x63
      12'hC5A: dout <= 8'b01100011; // 3162 :  99 - 0x63
      12'hC5B: dout <= 8'b01100011; // 3163 :  99 - 0x63
      12'hC5C: dout <= 8'b01100011; // 3164 :  99 - 0x63
      12'hC5D: dout <= 8'b01100011; // 3165 :  99 - 0x63
      12'hC5E: dout <= 8'b00111110; // 3166 :  62 - 0x3e
      12'hC5F: dout <= 8'b00000000; // 3167 :   0 - 0x0
      12'hC60: dout <= 8'b01111110; // 3168 : 126 - 0x7e -- Background 0xc6
      12'hC61: dout <= 8'b01100011; // 3169 :  99 - 0x63
      12'hC62: dout <= 8'b01100011; // 3170 :  99 - 0x63
      12'hC63: dout <= 8'b01100111; // 3171 : 103 - 0x67
      12'hC64: dout <= 8'b01111100; // 3172 : 124 - 0x7c
      12'hC65: dout <= 8'b01101110; // 3173 : 110 - 0x6e
      12'hC66: dout <= 8'b01100111; // 3174 : 103 - 0x67
      12'hC67: dout <= 8'b00000000; // 3175 :   0 - 0x0
      12'hC68: dout <= 8'b01111110; // 3176 : 126 - 0x7e -- plane 1
      12'hC69: dout <= 8'b01100011; // 3177 :  99 - 0x63
      12'hC6A: dout <= 8'b01100011; // 3178 :  99 - 0x63
      12'hC6B: dout <= 8'b01100111; // 3179 : 103 - 0x67
      12'hC6C: dout <= 8'b01111100; // 3180 : 124 - 0x7c
      12'hC6D: dout <= 8'b01101110; // 3181 : 110 - 0x6e
      12'hC6E: dout <= 8'b01100111; // 3182 : 103 - 0x67
      12'hC6F: dout <= 8'b00000000; // 3183 :   0 - 0x0
      12'hC70: dout <= 8'b01111111; // 3184 : 127 - 0x7f -- Background 0xc7
      12'hC71: dout <= 8'b01100000; // 3185 :  96 - 0x60
      12'hC72: dout <= 8'b01100000; // 3186 :  96 - 0x60
      12'hC73: dout <= 8'b01111110; // 3187 : 126 - 0x7e
      12'hC74: dout <= 8'b01100000; // 3188 :  96 - 0x60
      12'hC75: dout <= 8'b01100000; // 3189 :  96 - 0x60
      12'hC76: dout <= 8'b01111111; // 3190 : 127 - 0x7f
      12'hC77: dout <= 8'b00000000; // 3191 :   0 - 0x0
      12'hC78: dout <= 8'b01111111; // 3192 : 127 - 0x7f -- plane 1
      12'hC79: dout <= 8'b01100000; // 3193 :  96 - 0x60
      12'hC7A: dout <= 8'b01100000; // 3194 :  96 - 0x60
      12'hC7B: dout <= 8'b01111110; // 3195 : 126 - 0x7e
      12'hC7C: dout <= 8'b01100000; // 3196 :  96 - 0x60
      12'hC7D: dout <= 8'b01100000; // 3197 :  96 - 0x60
      12'hC7E: dout <= 8'b01111111; // 3198 : 127 - 0x7f
      12'hC7F: dout <= 8'b00000000; // 3199 :   0 - 0x0
      12'hC80: dout <= 8'b00110110; // 3200 :  54 - 0x36 -- Background 0xc8
      12'hC81: dout <= 8'b00110110; // 3201 :  54 - 0x36
      12'hC82: dout <= 8'b00010010; // 3202 :  18 - 0x12
      12'hC83: dout <= 8'b00000000; // 3203 :   0 - 0x0
      12'hC84: dout <= 8'b00000000; // 3204 :   0 - 0x0
      12'hC85: dout <= 8'b00000000; // 3205 :   0 - 0x0
      12'hC86: dout <= 8'b00000000; // 3206 :   0 - 0x0
      12'hC87: dout <= 8'b00000000; // 3207 :   0 - 0x0
      12'hC88: dout <= 8'b00110110; // 3208 :  54 - 0x36 -- plane 1
      12'hC89: dout <= 8'b00110110; // 3209 :  54 - 0x36
      12'hC8A: dout <= 8'b00010010; // 3210 :  18 - 0x12
      12'hC8B: dout <= 8'b00000000; // 3211 :   0 - 0x0
      12'hC8C: dout <= 8'b00000000; // 3212 :   0 - 0x0
      12'hC8D: dout <= 8'b00000000; // 3213 :   0 - 0x0
      12'hC8E: dout <= 8'b00000000; // 3214 :   0 - 0x0
      12'hC8F: dout <= 8'b00000000; // 3215 :   0 - 0x0
      12'hC90: dout <= 8'b00111110; // 3216 :  62 - 0x3e -- Background 0xc9
      12'hC91: dout <= 8'b01100011; // 3217 :  99 - 0x63
      12'hC92: dout <= 8'b01100011; // 3218 :  99 - 0x63
      12'hC93: dout <= 8'b01100011; // 3219 :  99 - 0x63
      12'hC94: dout <= 8'b01100011; // 3220 :  99 - 0x63
      12'hC95: dout <= 8'b01100011; // 3221 :  99 - 0x63
      12'hC96: dout <= 8'b00111110; // 3222 :  62 - 0x3e
      12'hC97: dout <= 8'b00000000; // 3223 :   0 - 0x0
      12'hC98: dout <= 8'b00111110; // 3224 :  62 - 0x3e -- plane 1
      12'hC99: dout <= 8'b01100011; // 3225 :  99 - 0x63
      12'hC9A: dout <= 8'b01100011; // 3226 :  99 - 0x63
      12'hC9B: dout <= 8'b01100011; // 3227 :  99 - 0x63
      12'hC9C: dout <= 8'b01100011; // 3228 :  99 - 0x63
      12'hC9D: dout <= 8'b01100011; // 3229 :  99 - 0x63
      12'hC9E: dout <= 8'b00111110; // 3230 :  62 - 0x3e
      12'hC9F: dout <= 8'b00000000; // 3231 :   0 - 0x0
      12'hCA0: dout <= 8'b00111100; // 3232 :  60 - 0x3c -- Background 0xca
      12'hCA1: dout <= 8'b01100110; // 3233 : 102 - 0x66
      12'hCA2: dout <= 8'b01100000; // 3234 :  96 - 0x60
      12'hCA3: dout <= 8'b00111110; // 3235 :  62 - 0x3e
      12'hCA4: dout <= 8'b00000011; // 3236 :   3 - 0x3
      12'hCA5: dout <= 8'b01100011; // 3237 :  99 - 0x63
      12'hCA6: dout <= 8'b00111110; // 3238 :  62 - 0x3e
      12'hCA7: dout <= 8'b00000000; // 3239 :   0 - 0x0
      12'hCA8: dout <= 8'b00111100; // 3240 :  60 - 0x3c -- plane 1
      12'hCA9: dout <= 8'b01100110; // 3241 : 102 - 0x66
      12'hCAA: dout <= 8'b01100000; // 3242 :  96 - 0x60
      12'hCAB: dout <= 8'b00111110; // 3243 :  62 - 0x3e
      12'hCAC: dout <= 8'b00000011; // 3244 :   3 - 0x3
      12'hCAD: dout <= 8'b01100011; // 3245 :  99 - 0x63
      12'hCAE: dout <= 8'b00111110; // 3246 :  62 - 0x3e
      12'hCAF: dout <= 8'b00000000; // 3247 :   0 - 0x0
      12'hCB0: dout <= 8'b00000000; // 3248 :   0 - 0x0 -- Background 0xcb
      12'hCB1: dout <= 8'b00000000; // 3249 :   0 - 0x0
      12'hCB2: dout <= 8'b00000000; // 3250 :   0 - 0x0
      12'hCB3: dout <= 8'b00000000; // 3251 :   0 - 0x0
      12'hCB4: dout <= 8'b00000000; // 3252 :   0 - 0x0
      12'hCB5: dout <= 8'b00000000; // 3253 :   0 - 0x0
      12'hCB6: dout <= 8'b00000000; // 3254 :   0 - 0x0
      12'hCB7: dout <= 8'b00000000; // 3255 :   0 - 0x0
      12'hCB8: dout <= 8'b00000000; // 3256 :   0 - 0x0 -- plane 1
      12'hCB9: dout <= 8'b00111000; // 3257 :  56 - 0x38
      12'hCBA: dout <= 8'b01111100; // 3258 : 124 - 0x7c
      12'hCBB: dout <= 8'b11111110; // 3259 : 254 - 0xfe
      12'hCBC: dout <= 8'b11111110; // 3260 : 254 - 0xfe
      12'hCBD: dout <= 8'b11111110; // 3261 : 254 - 0xfe
      12'hCBE: dout <= 8'b01111100; // 3262 : 124 - 0x7c
      12'hCBF: dout <= 8'b00111000; // 3263 :  56 - 0x38
      12'hCC0: dout <= 8'b00000000; // 3264 :   0 - 0x0 -- Background 0xcc
      12'hCC1: dout <= 8'b00000000; // 3265 :   0 - 0x0
      12'hCC2: dout <= 8'b00000000; // 3266 :   0 - 0x0
      12'hCC3: dout <= 8'b00000000; // 3267 :   0 - 0x0
      12'hCC4: dout <= 8'b00000000; // 3268 :   0 - 0x0
      12'hCC5: dout <= 8'b00000000; // 3269 :   0 - 0x0
      12'hCC6: dout <= 8'b00000000; // 3270 :   0 - 0x0
      12'hCC7: dout <= 8'b00000000; // 3271 :   0 - 0x0
      12'hCC8: dout <= 8'b00000000; // 3272 :   0 - 0x0 -- plane 1
      12'hCC9: dout <= 8'b00000000; // 3273 :   0 - 0x0
      12'hCCA: dout <= 8'b00000000; // 3274 :   0 - 0x0
      12'hCCB: dout <= 8'b00000000; // 3275 :   0 - 0x0
      12'hCCC: dout <= 8'b00000000; // 3276 :   0 - 0x0
      12'hCCD: dout <= 8'b00000000; // 3277 :   0 - 0x0
      12'hCCE: dout <= 8'b00000000; // 3278 :   0 - 0x0
      12'hCCF: dout <= 8'b00000000; // 3279 :   0 - 0x0
      12'hCD0: dout <= 8'b00000000; // 3280 :   0 - 0x0 -- Background 0xcd
      12'hCD1: dout <= 8'b00000000; // 3281 :   0 - 0x0
      12'hCD2: dout <= 8'b00000000; // 3282 :   0 - 0x0
      12'hCD3: dout <= 8'b00000000; // 3283 :   0 - 0x0
      12'hCD4: dout <= 8'b00000000; // 3284 :   0 - 0x0
      12'hCD5: dout <= 8'b00000000; // 3285 :   0 - 0x0
      12'hCD6: dout <= 8'b00000000; // 3286 :   0 - 0x0
      12'hCD7: dout <= 8'b00000000; // 3287 :   0 - 0x0
      12'hCD8: dout <= 8'b00000000; // 3288 :   0 - 0x0 -- plane 1
      12'hCD9: dout <= 8'b00000000; // 3289 :   0 - 0x0
      12'hCDA: dout <= 8'b00000000; // 3290 :   0 - 0x0
      12'hCDB: dout <= 8'b00000000; // 3291 :   0 - 0x0
      12'hCDC: dout <= 8'b00000000; // 3292 :   0 - 0x0
      12'hCDD: dout <= 8'b00000000; // 3293 :   0 - 0x0
      12'hCDE: dout <= 8'b00000000; // 3294 :   0 - 0x0
      12'hCDF: dout <= 8'b00000000; // 3295 :   0 - 0x0
      12'hCE0: dout <= 8'b00000000; // 3296 :   0 - 0x0 -- Background 0xce
      12'hCE1: dout <= 8'b00000000; // 3297 :   0 - 0x0
      12'hCE2: dout <= 8'b00000000; // 3298 :   0 - 0x0
      12'hCE3: dout <= 8'b00000000; // 3299 :   0 - 0x0
      12'hCE4: dout <= 8'b00000000; // 3300 :   0 - 0x0
      12'hCE5: dout <= 8'b00000000; // 3301 :   0 - 0x0
      12'hCE6: dout <= 8'b00000000; // 3302 :   0 - 0x0
      12'hCE7: dout <= 8'b00000000; // 3303 :   0 - 0x0
      12'hCE8: dout <= 8'b00000000; // 3304 :   0 - 0x0 -- plane 1
      12'hCE9: dout <= 8'b00000000; // 3305 :   0 - 0x0
      12'hCEA: dout <= 8'b00000000; // 3306 :   0 - 0x0
      12'hCEB: dout <= 8'b00000000; // 3307 :   0 - 0x0
      12'hCEC: dout <= 8'b00000000; // 3308 :   0 - 0x0
      12'hCED: dout <= 8'b00000000; // 3309 :   0 - 0x0
      12'hCEE: dout <= 8'b00000000; // 3310 :   0 - 0x0
      12'hCEF: dout <= 8'b00000000; // 3311 :   0 - 0x0
      12'hCF0: dout <= 8'b00000000; // 3312 :   0 - 0x0 -- Background 0xcf
      12'hCF1: dout <= 8'b00000000; // 3313 :   0 - 0x0
      12'hCF2: dout <= 8'b00000000; // 3314 :   0 - 0x0
      12'hCF3: dout <= 8'b00000000; // 3315 :   0 - 0x0
      12'hCF4: dout <= 8'b00000000; // 3316 :   0 - 0x0
      12'hCF5: dout <= 8'b00000000; // 3317 :   0 - 0x0
      12'hCF6: dout <= 8'b00000000; // 3318 :   0 - 0x0
      12'hCF7: dout <= 8'b00000000; // 3319 :   0 - 0x0
      12'hCF8: dout <= 8'b00000000; // 3320 :   0 - 0x0 -- plane 1
      12'hCF9: dout <= 8'b00000000; // 3321 :   0 - 0x0
      12'hCFA: dout <= 8'b00000000; // 3322 :   0 - 0x0
      12'hCFB: dout <= 8'b00000000; // 3323 :   0 - 0x0
      12'hCFC: dout <= 8'b00000000; // 3324 :   0 - 0x0
      12'hCFD: dout <= 8'b00000000; // 3325 :   0 - 0x0
      12'hCFE: dout <= 8'b00000000; // 3326 :   0 - 0x0
      12'hCFF: dout <= 8'b00000000; // 3327 :   0 - 0x0
      12'hD00: dout <= 8'b01000111; // 3328 :  71 - 0x47 -- Background 0xd0
      12'hD01: dout <= 8'b01000111; // 3329 :  71 - 0x47
      12'hD02: dout <= 8'b00001111; // 3330 :  15 - 0xf
      12'hD03: dout <= 8'b00001111; // 3331 :  15 - 0xf
      12'hD04: dout <= 8'b00011111; // 3332 :  31 - 0x1f
      12'hD05: dout <= 8'b00011111; // 3333 :  31 - 0x1f
      12'hD06: dout <= 8'b00111111; // 3334 :  63 - 0x3f
      12'hD07: dout <= 8'b00111111; // 3335 :  63 - 0x3f
      12'hD08: dout <= 8'b00010111; // 3336 :  23 - 0x17 -- plane 1
      12'hD09: dout <= 8'b00010111; // 3337 :  23 - 0x17
      12'hD0A: dout <= 8'b00101111; // 3338 :  47 - 0x2f
      12'hD0B: dout <= 8'b00101111; // 3339 :  47 - 0x2f
      12'hD0C: dout <= 8'b01011111; // 3340 :  95 - 0x5f
      12'hD0D: dout <= 8'b01011111; // 3341 :  95 - 0x5f
      12'hD0E: dout <= 8'b00111111; // 3342 :  63 - 0x3f
      12'hD0F: dout <= 8'b00111111; // 3343 :  63 - 0x3f
      12'hD10: dout <= 8'b11111111; // 3344 : 255 - 0xff -- Background 0xd1
      12'hD11: dout <= 8'b11001111; // 3345 : 207 - 0xcf
      12'hD12: dout <= 8'b11001111; // 3346 : 207 - 0xcf
      12'hD13: dout <= 8'b11111011; // 3347 : 251 - 0xfb
      12'hD14: dout <= 8'b11110111; // 3348 : 247 - 0xf7
      12'hD15: dout <= 8'b11100111; // 3349 : 231 - 0xe7
      12'hD16: dout <= 8'b11111111; // 3350 : 255 - 0xff
      12'hD17: dout <= 8'b11111111; // 3351 : 255 - 0xff
      12'hD18: dout <= 8'b11111111; // 3352 : 255 - 0xff -- plane 1
      12'hD19: dout <= 8'b11001111; // 3353 : 207 - 0xcf
      12'hD1A: dout <= 8'b11001111; // 3354 : 207 - 0xcf
      12'hD1B: dout <= 8'b11111011; // 3355 : 251 - 0xfb
      12'hD1C: dout <= 8'b11110111; // 3356 : 247 - 0xf7
      12'hD1D: dout <= 8'b11100111; // 3357 : 231 - 0xe7
      12'hD1E: dout <= 8'b11111111; // 3358 : 255 - 0xff
      12'hD1F: dout <= 8'b11111111; // 3359 : 255 - 0xff
      12'hD20: dout <= 8'b00011000; // 3360 :  24 - 0x18 -- Background 0xd2
      12'hD21: dout <= 8'b00001000; // 3361 :   8 - 0x8
      12'hD22: dout <= 8'b10001000; // 3362 : 136 - 0x88
      12'hD23: dout <= 8'b10000000; // 3363 : 128 - 0x80
      12'hD24: dout <= 8'b01000000; // 3364 :  64 - 0x40
      12'hD25: dout <= 8'b01000000; // 3365 :  64 - 0x40
      12'hD26: dout <= 8'b10100000; // 3366 : 160 - 0xa0
      12'hD27: dout <= 8'b10100000; // 3367 : 160 - 0xa0
      12'hD28: dout <= 8'b01000010; // 3368 :  66 - 0x42 -- plane 1
      12'hD29: dout <= 8'b01100010; // 3369 :  98 - 0x62
      12'hD2A: dout <= 8'b10100010; // 3370 : 162 - 0xa2
      12'hD2B: dout <= 8'b10110010; // 3371 : 178 - 0xb2
      12'hD2C: dout <= 8'b01010010; // 3372 :  82 - 0x52
      12'hD2D: dout <= 8'b01011010; // 3373 :  90 - 0x5a
      12'hD2E: dout <= 8'b10101010; // 3374 : 170 - 0xaa
      12'hD2F: dout <= 8'b10101100; // 3375 : 172 - 0xac
      12'hD30: dout <= 8'b11111111; // 3376 : 255 - 0xff -- Background 0xd3
      12'hD31: dout <= 8'b11111111; // 3377 : 255 - 0xff
      12'hD32: dout <= 8'b11111111; // 3378 : 255 - 0xff
      12'hD33: dout <= 8'b11111111; // 3379 : 255 - 0xff
      12'hD34: dout <= 8'b11111101; // 3380 : 253 - 0xfd
      12'hD35: dout <= 8'b11111101; // 3381 : 253 - 0xfd
      12'hD36: dout <= 8'b11111101; // 3382 : 253 - 0xfd
      12'hD37: dout <= 8'b11111101; // 3383 : 253 - 0xfd
      12'hD38: dout <= 8'b11111111; // 3384 : 255 - 0xff -- plane 1
      12'hD39: dout <= 8'b11111111; // 3385 : 255 - 0xff
      12'hD3A: dout <= 8'b11111111; // 3386 : 255 - 0xff
      12'hD3B: dout <= 8'b11111111; // 3387 : 255 - 0xff
      12'hD3C: dout <= 8'b11111101; // 3388 : 253 - 0xfd
      12'hD3D: dout <= 8'b11111101; // 3389 : 253 - 0xfd
      12'hD3E: dout <= 8'b11111101; // 3390 : 253 - 0xfd
      12'hD3F: dout <= 8'b11111101; // 3391 : 253 - 0xfd
      12'hD40: dout <= 8'b11000111; // 3392 : 199 - 0xc7 -- Background 0xd4
      12'hD41: dout <= 8'b11110111; // 3393 : 247 - 0xf7
      12'hD42: dout <= 8'b11110000; // 3394 : 240 - 0xf0
      12'hD43: dout <= 8'b11111000; // 3395 : 248 - 0xf8
      12'hD44: dout <= 8'b11111000; // 3396 : 248 - 0xf8
      12'hD45: dout <= 8'b11111111; // 3397 : 255 - 0xff
      12'hD46: dout <= 8'b11111111; // 3398 : 255 - 0xff
      12'hD47: dout <= 8'b11111111; // 3399 : 255 - 0xff
      12'hD48: dout <= 8'b00000111; // 3400 :   7 - 0x7 -- plane 1
      12'hD49: dout <= 8'b00000111; // 3401 :   7 - 0x7
      12'hD4A: dout <= 8'b00000000; // 3402 :   0 - 0x0
      12'hD4B: dout <= 8'b00000011; // 3403 :   3 - 0x3
      12'hD4C: dout <= 8'b00000000; // 3404 :   0 - 0x0
      12'hD4D: dout <= 8'b00000000; // 3405 :   0 - 0x0
      12'hD4E: dout <= 8'b00000000; // 3406 :   0 - 0x0
      12'hD4F: dout <= 8'b00000000; // 3407 :   0 - 0x0
      12'hD50: dout <= 8'b11111000; // 3408 : 248 - 0xf8 -- Background 0xd5
      12'hD51: dout <= 8'b11111000; // 3409 : 248 - 0xf8
      12'hD52: dout <= 8'b00000000; // 3410 :   0 - 0x0
      12'hD53: dout <= 8'b00000000; // 3411 :   0 - 0x0
      12'hD54: dout <= 8'b00000000; // 3412 :   0 - 0x0
      12'hD55: dout <= 8'b11111111; // 3413 : 255 - 0xff
      12'hD56: dout <= 8'b11111111; // 3414 : 255 - 0xff
      12'hD57: dout <= 8'b11111111; // 3415 : 255 - 0xff
      12'hD58: dout <= 8'b11111010; // 3416 : 250 - 0xfa -- plane 1
      12'hD59: dout <= 8'b11111010; // 3417 : 250 - 0xfa
      12'hD5A: dout <= 8'b00000010; // 3418 :   2 - 0x2
      12'hD5B: dout <= 8'b11111110; // 3419 : 254 - 0xfe
      12'hD5C: dout <= 8'b00000000; // 3420 :   0 - 0x0
      12'hD5D: dout <= 8'b00000000; // 3421 :   0 - 0x0
      12'hD5E: dout <= 8'b00000000; // 3422 :   0 - 0x0
      12'hD5F: dout <= 8'b00000000; // 3423 :   0 - 0x0
      12'hD60: dout <= 8'b10001111; // 3424 : 143 - 0x8f -- Background 0xd6
      12'hD61: dout <= 8'b11101111; // 3425 : 239 - 0xef
      12'hD62: dout <= 8'b11000000; // 3426 : 192 - 0xc0
      12'hD63: dout <= 8'b11110000; // 3427 : 240 - 0xf0
      12'hD64: dout <= 8'b11100000; // 3428 : 224 - 0xe0
      12'hD65: dout <= 8'b11111111; // 3429 : 255 - 0xff
      12'hD66: dout <= 8'b11111111; // 3430 : 255 - 0xff
      12'hD67: dout <= 8'b11111111; // 3431 : 255 - 0xff
      12'hD68: dout <= 8'b00001111; // 3432 :  15 - 0xf -- plane 1
      12'hD69: dout <= 8'b00001111; // 3433 :  15 - 0xf
      12'hD6A: dout <= 8'b00000000; // 3434 :   0 - 0x0
      12'hD6B: dout <= 8'b00000111; // 3435 :   7 - 0x7
      12'hD6C: dout <= 8'b00000000; // 3436 :   0 - 0x0
      12'hD6D: dout <= 8'b00000000; // 3437 :   0 - 0x0
      12'hD6E: dout <= 8'b00000000; // 3438 :   0 - 0x0
      12'hD6F: dout <= 8'b00000000; // 3439 :   0 - 0x0
      12'hD70: dout <= 8'b11111111; // 3440 : 255 - 0xff -- Background 0xd7
      12'hD71: dout <= 8'b11111111; // 3441 : 255 - 0xff
      12'hD72: dout <= 8'b00000000; // 3442 :   0 - 0x0
      12'hD73: dout <= 8'b00000000; // 3443 :   0 - 0x0
      12'hD74: dout <= 8'b00000000; // 3444 :   0 - 0x0
      12'hD75: dout <= 8'b11111111; // 3445 : 255 - 0xff
      12'hD76: dout <= 8'b11111111; // 3446 : 255 - 0xff
      12'hD77: dout <= 8'b11111111; // 3447 : 255 - 0xff
      12'hD78: dout <= 8'b11111111; // 3448 : 255 - 0xff -- plane 1
      12'hD79: dout <= 8'b11111111; // 3449 : 255 - 0xff
      12'hD7A: dout <= 8'b00000000; // 3450 :   0 - 0x0
      12'hD7B: dout <= 8'b11111111; // 3451 : 255 - 0xff
      12'hD7C: dout <= 8'b00000000; // 3452 :   0 - 0x0
      12'hD7D: dout <= 8'b00000000; // 3453 :   0 - 0x0
      12'hD7E: dout <= 8'b00000000; // 3454 :   0 - 0x0
      12'hD7F: dout <= 8'b00000000; // 3455 :   0 - 0x0
      12'hD80: dout <= 8'b11000011; // 3456 : 195 - 0xc3 -- Background 0xd8
      12'hD81: dout <= 8'b11111111; // 3457 : 255 - 0xff
      12'hD82: dout <= 8'b00000000; // 3458 :   0 - 0x0
      12'hD83: dout <= 8'b00000000; // 3459 :   0 - 0x0
      12'hD84: dout <= 8'b00000000; // 3460 :   0 - 0x0
      12'hD85: dout <= 8'b11111111; // 3461 : 255 - 0xff
      12'hD86: dout <= 8'b11111111; // 3462 : 255 - 0xff
      12'hD87: dout <= 8'b11111111; // 3463 : 255 - 0xff
      12'hD88: dout <= 8'b11000011; // 3464 : 195 - 0xc3 -- plane 1
      12'hD89: dout <= 8'b11111111; // 3465 : 255 - 0xff
      12'hD8A: dout <= 8'b00000000; // 3466 :   0 - 0x0
      12'hD8B: dout <= 8'b11111111; // 3467 : 255 - 0xff
      12'hD8C: dout <= 8'b00000000; // 3468 :   0 - 0x0
      12'hD8D: dout <= 8'b00000000; // 3469 :   0 - 0x0
      12'hD8E: dout <= 8'b00000000; // 3470 :   0 - 0x0
      12'hD8F: dout <= 8'b00000000; // 3471 :   0 - 0x0
      12'hD90: dout <= 8'b00000011; // 3472 :   3 - 0x3 -- Background 0xd9
      12'hD91: dout <= 8'b10000001; // 3473 : 129 - 0x81
      12'hD92: dout <= 8'b00000000; // 3474 :   0 - 0x0
      12'hD93: dout <= 8'b00000000; // 3475 :   0 - 0x0
      12'hD94: dout <= 8'b00000011; // 3476 :   3 - 0x3
      12'hD95: dout <= 8'b11111111; // 3477 : 255 - 0xff
      12'hD96: dout <= 8'b11111111; // 3478 : 255 - 0xff
      12'hD97: dout <= 8'b11111111; // 3479 : 255 - 0xff
      12'hD98: dout <= 8'b01101011; // 3480 : 107 - 0x6b -- plane 1
      12'hD99: dout <= 8'b10110101; // 3481 : 181 - 0xb5
      12'hD9A: dout <= 8'b00110110; // 3482 :  54 - 0x36
      12'hD9B: dout <= 8'b11111000; // 3483 : 248 - 0xf8
      12'hD9C: dout <= 8'b00000000; // 3484 :   0 - 0x0
      12'hD9D: dout <= 8'b00000000; // 3485 :   0 - 0x0
      12'hD9E: dout <= 8'b00000000; // 3486 :   0 - 0x0
      12'hD9F: dout <= 8'b00000000; // 3487 :   0 - 0x0
      12'hDA0: dout <= 8'b11111111; // 3488 : 255 - 0xff -- Background 0xda
      12'hDA1: dout <= 8'b11111111; // 3489 : 255 - 0xff
      12'hDA2: dout <= 8'b01111110; // 3490 : 126 - 0x7e
      12'hDA3: dout <= 8'b00000000; // 3491 :   0 - 0x0
      12'hDA4: dout <= 8'b00000000; // 3492 :   0 - 0x0
      12'hDA5: dout <= 8'b11100000; // 3493 : 224 - 0xe0
      12'hDA6: dout <= 8'b11111111; // 3494 : 255 - 0xff
      12'hDA7: dout <= 8'b11111111; // 3495 : 255 - 0xff
      12'hDA8: dout <= 8'b11111111; // 3496 : 255 - 0xff -- plane 1
      12'hDA9: dout <= 8'b11111111; // 3497 : 255 - 0xff
      12'hDAA: dout <= 8'b01111110; // 3498 : 126 - 0x7e
      12'hDAB: dout <= 8'b10000001; // 3499 : 129 - 0x81
      12'hDAC: dout <= 8'b00011111; // 3500 :  31 - 0x1f
      12'hDAD: dout <= 8'b00000000; // 3501 :   0 - 0x0
      12'hDAE: dout <= 8'b00000000; // 3502 :   0 - 0x0
      12'hDAF: dout <= 8'b00000000; // 3503 :   0 - 0x0
      12'hDB0: dout <= 8'b01100001; // 3504 :  97 - 0x61 -- Background 0xdb
      12'hDB1: dout <= 8'b11000011; // 3505 : 195 - 0xc3
      12'hDB2: dout <= 8'b00000111; // 3506 :   7 - 0x7
      12'hDB3: dout <= 8'b00001111; // 3507 :  15 - 0xf
      12'hDB4: dout <= 8'b00011111; // 3508 :  31 - 0x1f
      12'hDB5: dout <= 8'b01111111; // 3509 : 127 - 0x7f
      12'hDB6: dout <= 8'b11111111; // 3510 : 255 - 0xff
      12'hDB7: dout <= 8'b11111111; // 3511 : 255 - 0xff
      12'hDB8: dout <= 8'b01101100; // 3512 : 108 - 0x6c -- plane 1
      12'hDB9: dout <= 8'b11011000; // 3513 : 216 - 0xd8
      12'hDBA: dout <= 8'b00110000; // 3514 :  48 - 0x30
      12'hDBB: dout <= 8'b11100000; // 3515 : 224 - 0xe0
      12'hDBC: dout <= 8'b10000000; // 3516 : 128 - 0x80
      12'hDBD: dout <= 8'b00000000; // 3517 :   0 - 0x0
      12'hDBE: dout <= 8'b00000000; // 3518 :   0 - 0x0
      12'hDBF: dout <= 8'b00000000; // 3519 :   0 - 0x0
      12'hDC0: dout <= 8'b00011111; // 3520 :  31 - 0x1f -- Background 0xdc
      12'hDC1: dout <= 8'b11011111; // 3521 : 223 - 0xdf
      12'hDC2: dout <= 8'b11000000; // 3522 : 192 - 0xc0
      12'hDC3: dout <= 8'b11110000; // 3523 : 240 - 0xf0
      12'hDC4: dout <= 8'b11110000; // 3524 : 240 - 0xf0
      12'hDC5: dout <= 8'b11111111; // 3525 : 255 - 0xff
      12'hDC6: dout <= 8'b11111111; // 3526 : 255 - 0xff
      12'hDC7: dout <= 8'b11111111; // 3527 : 255 - 0xff
      12'hDC8: dout <= 8'b00011111; // 3528 :  31 - 0x1f -- plane 1
      12'hDC9: dout <= 8'b00011111; // 3529 :  31 - 0x1f
      12'hDCA: dout <= 8'b00000000; // 3530 :   0 - 0x0
      12'hDCB: dout <= 8'b00000111; // 3531 :   7 - 0x7
      12'hDCC: dout <= 8'b00000000; // 3532 :   0 - 0x0
      12'hDCD: dout <= 8'b00000000; // 3533 :   0 - 0x0
      12'hDCE: dout <= 8'b00000000; // 3534 :   0 - 0x0
      12'hDCF: dout <= 8'b00000000; // 3535 :   0 - 0x0
      12'hDD0: dout <= 8'b10000100; // 3536 : 132 - 0x84 -- Background 0xdd
      12'hDD1: dout <= 8'b11111100; // 3537 : 252 - 0xfc
      12'hDD2: dout <= 8'b00000000; // 3538 :   0 - 0x0
      12'hDD3: dout <= 8'b00000000; // 3539 :   0 - 0x0
      12'hDD4: dout <= 8'b00000000; // 3540 :   0 - 0x0
      12'hDD5: dout <= 8'b11111111; // 3541 : 255 - 0xff
      12'hDD6: dout <= 8'b11111111; // 3542 : 255 - 0xff
      12'hDD7: dout <= 8'b11111111; // 3543 : 255 - 0xff
      12'hDD8: dout <= 8'b10000101; // 3544 : 133 - 0x85 -- plane 1
      12'hDD9: dout <= 8'b11111101; // 3545 : 253 - 0xfd
      12'hDDA: dout <= 8'b00000001; // 3546 :   1 - 0x1
      12'hDDB: dout <= 8'b11111111; // 3547 : 255 - 0xff
      12'hDDC: dout <= 8'b00000000; // 3548 :   0 - 0x0
      12'hDDD: dout <= 8'b00000000; // 3549 :   0 - 0x0
      12'hDDE: dout <= 8'b00000000; // 3550 :   0 - 0x0
      12'hDDF: dout <= 8'b00000000; // 3551 :   0 - 0x0
      12'hDE0: dout <= 8'b01111111; // 3552 : 127 - 0x7f -- Background 0xde
      12'hDE1: dout <= 8'b01111111; // 3553 : 127 - 0x7f
      12'hDE2: dout <= 8'b00000000; // 3554 :   0 - 0x0
      12'hDE3: dout <= 8'b00000000; // 3555 :   0 - 0x0
      12'hDE4: dout <= 8'b00000000; // 3556 :   0 - 0x0
      12'hDE5: dout <= 8'b11111111; // 3557 : 255 - 0xff
      12'hDE6: dout <= 8'b11111111; // 3558 : 255 - 0xff
      12'hDE7: dout <= 8'b11111111; // 3559 : 255 - 0xff
      12'hDE8: dout <= 8'b01111111; // 3560 : 127 - 0x7f -- plane 1
      12'hDE9: dout <= 8'b01111111; // 3561 : 127 - 0x7f
      12'hDEA: dout <= 8'b00000000; // 3562 :   0 - 0x0
      12'hDEB: dout <= 8'b01011111; // 3563 :  95 - 0x5f
      12'hDEC: dout <= 8'b00000000; // 3564 :   0 - 0x0
      12'hDED: dout <= 8'b00000000; // 3565 :   0 - 0x0
      12'hDEE: dout <= 8'b00000000; // 3566 :   0 - 0x0
      12'hDEF: dout <= 8'b00000000; // 3567 :   0 - 0x0
      12'hDF0: dout <= 8'b11111100; // 3568 : 252 - 0xfc -- Background 0xdf
      12'hDF1: dout <= 8'b11111111; // 3569 : 255 - 0xff
      12'hDF2: dout <= 8'b00000000; // 3570 :   0 - 0x0
      12'hDF3: dout <= 8'b00000000; // 3571 :   0 - 0x0
      12'hDF4: dout <= 8'b00000000; // 3572 :   0 - 0x0
      12'hDF5: dout <= 8'b11111111; // 3573 : 255 - 0xff
      12'hDF6: dout <= 8'b11111111; // 3574 : 255 - 0xff
      12'hDF7: dout <= 8'b11111111; // 3575 : 255 - 0xff
      12'hDF8: dout <= 8'b11111100; // 3576 : 252 - 0xfc -- plane 1
      12'hDF9: dout <= 8'b11111111; // 3577 : 255 - 0xff
      12'hDFA: dout <= 8'b00000000; // 3578 :   0 - 0x0
      12'hDFB: dout <= 8'b11111111; // 3579 : 255 - 0xff
      12'hDFC: dout <= 8'b00000000; // 3580 :   0 - 0x0
      12'hDFD: dout <= 8'b00000000; // 3581 :   0 - 0x0
      12'hDFE: dout <= 8'b00000000; // 3582 :   0 - 0x0
      12'hDFF: dout <= 8'b00000000; // 3583 :   0 - 0x0
      12'hE00: dout <= 8'b00110000; // 3584 :  48 - 0x30 -- Background 0xe0
      12'hE01: dout <= 8'b11110000; // 3585 : 240 - 0xf0
      12'hE02: dout <= 8'b00000000; // 3586 :   0 - 0x0
      12'hE03: dout <= 8'b00000000; // 3587 :   0 - 0x0
      12'hE04: dout <= 8'b00000000; // 3588 :   0 - 0x0
      12'hE05: dout <= 8'b11111111; // 3589 : 255 - 0xff
      12'hE06: dout <= 8'b11111111; // 3590 : 255 - 0xff
      12'hE07: dout <= 8'b11111111; // 3591 : 255 - 0xff
      12'hE08: dout <= 8'b00110100; // 3592 :  52 - 0x34 -- plane 1
      12'hE09: dout <= 8'b11110110; // 3593 : 246 - 0xf6
      12'hE0A: dout <= 8'b00000010; // 3594 :   2 - 0x2
      12'hE0B: dout <= 8'b11111111; // 3595 : 255 - 0xff
      12'hE0C: dout <= 8'b00000000; // 3596 :   0 - 0x0
      12'hE0D: dout <= 8'b00000000; // 3597 :   0 - 0x0
      12'hE0E: dout <= 8'b00000000; // 3598 :   0 - 0x0
      12'hE0F: dout <= 8'b00000000; // 3599 :   0 - 0x0
      12'hE10: dout <= 8'b11111111; // 3600 : 255 - 0xff -- Background 0xe1
      12'hE11: dout <= 8'b11111111; // 3601 : 255 - 0xff
      12'hE12: dout <= 8'b00000000; // 3602 :   0 - 0x0
      12'hE13: dout <= 8'b00000000; // 3603 :   0 - 0x0
      12'hE14: dout <= 8'b00000000; // 3604 :   0 - 0x0
      12'hE15: dout <= 8'b11111111; // 3605 : 255 - 0xff
      12'hE16: dout <= 8'b11111111; // 3606 : 255 - 0xff
      12'hE17: dout <= 8'b11111111; // 3607 : 255 - 0xff
      12'hE18: dout <= 8'b11111111; // 3608 : 255 - 0xff -- plane 1
      12'hE19: dout <= 8'b11111111; // 3609 : 255 - 0xff
      12'hE1A: dout <= 8'b00000000; // 3610 :   0 - 0x0
      12'hE1B: dout <= 8'b01111111; // 3611 : 127 - 0x7f
      12'hE1C: dout <= 8'b00000000; // 3612 :   0 - 0x0
      12'hE1D: dout <= 8'b00000000; // 3613 :   0 - 0x0
      12'hE1E: dout <= 8'b00000000; // 3614 :   0 - 0x0
      12'hE1F: dout <= 8'b00000000; // 3615 :   0 - 0x0
      12'hE20: dout <= 8'b11100001; // 3616 : 225 - 0xe1 -- Background 0xe2
      12'hE21: dout <= 8'b11111111; // 3617 : 255 - 0xff
      12'hE22: dout <= 8'b00000000; // 3618 :   0 - 0x0
      12'hE23: dout <= 8'b00000000; // 3619 :   0 - 0x0
      12'hE24: dout <= 8'b00000000; // 3620 :   0 - 0x0
      12'hE25: dout <= 8'b11111111; // 3621 : 255 - 0xff
      12'hE26: dout <= 8'b11111111; // 3622 : 255 - 0xff
      12'hE27: dout <= 8'b11111111; // 3623 : 255 - 0xff
      12'hE28: dout <= 8'b11100001; // 3624 : 225 - 0xe1 -- plane 1
      12'hE29: dout <= 8'b11111111; // 3625 : 255 - 0xff
      12'hE2A: dout <= 8'b00000000; // 3626 :   0 - 0x0
      12'hE2B: dout <= 8'b11111111; // 3627 : 255 - 0xff
      12'hE2C: dout <= 8'b00000000; // 3628 :   0 - 0x0
      12'hE2D: dout <= 8'b00000000; // 3629 :   0 - 0x0
      12'hE2E: dout <= 8'b00000000; // 3630 :   0 - 0x0
      12'hE2F: dout <= 8'b00000000; // 3631 :   0 - 0x0
      12'hE30: dout <= 8'b00011111; // 3632 :  31 - 0x1f -- Background 0xe3
      12'hE31: dout <= 8'b00011111; // 3633 :  31 - 0x1f
      12'hE32: dout <= 8'b00011111; // 3634 :  31 - 0x1f
      12'hE33: dout <= 8'b00011111; // 3635 :  31 - 0x1f
      12'hE34: dout <= 8'b00011111; // 3636 :  31 - 0x1f
      12'hE35: dout <= 8'b11111111; // 3637 : 255 - 0xff
      12'hE36: dout <= 8'b11111111; // 3638 : 255 - 0xff
      12'hE37: dout <= 8'b11111111; // 3639 : 255 - 0xff
      12'hE38: dout <= 8'b01000000; // 3640 :  64 - 0x40 -- plane 1
      12'hE39: dout <= 8'b01000000; // 3641 :  64 - 0x40
      12'hE3A: dout <= 8'b01000000; // 3642 :  64 - 0x40
      12'hE3B: dout <= 8'b11000000; // 3643 : 192 - 0xc0
      12'hE3C: dout <= 8'b00000000; // 3644 :   0 - 0x0
      12'hE3D: dout <= 8'b00000000; // 3645 :   0 - 0x0
      12'hE3E: dout <= 8'b00000000; // 3646 :   0 - 0x0
      12'hE3F: dout <= 8'b00000000; // 3647 :   0 - 0x0
      12'hE40: dout <= 8'b00000000; // 3648 :   0 - 0x0 -- Background 0xe4
      12'hE41: dout <= 8'b00011111; // 3649 :  31 - 0x1f
      12'hE42: dout <= 8'b00111111; // 3650 :  63 - 0x3f
      12'hE43: dout <= 8'b01111000; // 3651 : 120 - 0x78
      12'hE44: dout <= 8'b01110111; // 3652 : 119 - 0x77
      12'hE45: dout <= 8'b01101111; // 3653 : 111 - 0x6f
      12'hE46: dout <= 8'b01101111; // 3654 : 111 - 0x6f
      12'hE47: dout <= 8'b01101111; // 3655 : 111 - 0x6f
      12'hE48: dout <= 8'b00000000; // 3656 :   0 - 0x0 -- plane 1
      12'hE49: dout <= 8'b00000000; // 3657 :   0 - 0x0
      12'hE4A: dout <= 8'b00000000; // 3658 :   0 - 0x0
      12'hE4B: dout <= 8'b00000000; // 3659 :   0 - 0x0
      12'hE4C: dout <= 8'b00000111; // 3660 :   7 - 0x7
      12'hE4D: dout <= 8'b00001111; // 3661 :  15 - 0xf
      12'hE4E: dout <= 8'b00001111; // 3662 :  15 - 0xf
      12'hE4F: dout <= 8'b00001111; // 3663 :  15 - 0xf
      12'hE50: dout <= 8'b00000000; // 3664 :   0 - 0x0 -- Background 0xe5
      12'hE51: dout <= 8'b11111000; // 3665 : 248 - 0xf8
      12'hE52: dout <= 8'b11111100; // 3666 : 252 - 0xfc
      12'hE53: dout <= 8'b00011110; // 3667 :  30 - 0x1e
      12'hE54: dout <= 8'b11101110; // 3668 : 238 - 0xee
      12'hE55: dout <= 8'b11110110; // 3669 : 246 - 0xf6
      12'hE56: dout <= 8'b11110110; // 3670 : 246 - 0xf6
      12'hE57: dout <= 8'b11110110; // 3671 : 246 - 0xf6
      12'hE58: dout <= 8'b00000000; // 3672 :   0 - 0x0 -- plane 1
      12'hE59: dout <= 8'b00000000; // 3673 :   0 - 0x0
      12'hE5A: dout <= 8'b00000000; // 3674 :   0 - 0x0
      12'hE5B: dout <= 8'b00000000; // 3675 :   0 - 0x0
      12'hE5C: dout <= 8'b11100000; // 3676 : 224 - 0xe0
      12'hE5D: dout <= 8'b11110000; // 3677 : 240 - 0xf0
      12'hE5E: dout <= 8'b11110000; // 3678 : 240 - 0xf0
      12'hE5F: dout <= 8'b11110000; // 3679 : 240 - 0xf0
      12'hE60: dout <= 8'b11110110; // 3680 : 246 - 0xf6 -- Background 0xe6
      12'hE61: dout <= 8'b11110110; // 3681 : 246 - 0xf6
      12'hE62: dout <= 8'b11110110; // 3682 : 246 - 0xf6
      12'hE63: dout <= 8'b11101110; // 3683 : 238 - 0xee
      12'hE64: dout <= 8'b00011110; // 3684 :  30 - 0x1e
      12'hE65: dout <= 8'b11111100; // 3685 : 252 - 0xfc
      12'hE66: dout <= 8'b11111000; // 3686 : 248 - 0xf8
      12'hE67: dout <= 8'b00000000; // 3687 :   0 - 0x0
      12'hE68: dout <= 8'b11110000; // 3688 : 240 - 0xf0 -- plane 1
      12'hE69: dout <= 8'b11110000; // 3689 : 240 - 0xf0
      12'hE6A: dout <= 8'b11110000; // 3690 : 240 - 0xf0
      12'hE6B: dout <= 8'b11100000; // 3691 : 224 - 0xe0
      12'hE6C: dout <= 8'b00000000; // 3692 :   0 - 0x0
      12'hE6D: dout <= 8'b00000000; // 3693 :   0 - 0x0
      12'hE6E: dout <= 8'b00000000; // 3694 :   0 - 0x0
      12'hE6F: dout <= 8'b00000000; // 3695 :   0 - 0x0
      12'hE70: dout <= 8'b01101111; // 3696 : 111 - 0x6f -- Background 0xe7
      12'hE71: dout <= 8'b01101111; // 3697 : 111 - 0x6f
      12'hE72: dout <= 8'b01101111; // 3698 : 111 - 0x6f
      12'hE73: dout <= 8'b01110111; // 3699 : 119 - 0x77
      12'hE74: dout <= 8'b01111000; // 3700 : 120 - 0x78
      12'hE75: dout <= 8'b00111111; // 3701 :  63 - 0x3f
      12'hE76: dout <= 8'b00011111; // 3702 :  31 - 0x1f
      12'hE77: dout <= 8'b00000000; // 3703 :   0 - 0x0
      12'hE78: dout <= 8'b00001111; // 3704 :  15 - 0xf -- plane 1
      12'hE79: dout <= 8'b00001111; // 3705 :  15 - 0xf
      12'hE7A: dout <= 8'b00001111; // 3706 :  15 - 0xf
      12'hE7B: dout <= 8'b00000111; // 3707 :   7 - 0x7
      12'hE7C: dout <= 8'b00000000; // 3708 :   0 - 0x0
      12'hE7D: dout <= 8'b00000000; // 3709 :   0 - 0x0
      12'hE7E: dout <= 8'b00000000; // 3710 :   0 - 0x0
      12'hE7F: dout <= 8'b00000000; // 3711 :   0 - 0x0
      12'hE80: dout <= 8'b00000000; // 3712 :   0 - 0x0 -- Background 0xe8
      12'hE81: dout <= 8'b11111111; // 3713 : 255 - 0xff
      12'hE82: dout <= 8'b11111111; // 3714 : 255 - 0xff
      12'hE83: dout <= 8'b00000000; // 3715 :   0 - 0x0
      12'hE84: dout <= 8'b11111111; // 3716 : 255 - 0xff
      12'hE85: dout <= 8'b11111111; // 3717 : 255 - 0xff
      12'hE86: dout <= 8'b11111111; // 3718 : 255 - 0xff
      12'hE87: dout <= 8'b11111111; // 3719 : 255 - 0xff
      12'hE88: dout <= 8'b00000000; // 3720 :   0 - 0x0 -- plane 1
      12'hE89: dout <= 8'b00000000; // 3721 :   0 - 0x0
      12'hE8A: dout <= 8'b00000000; // 3722 :   0 - 0x0
      12'hE8B: dout <= 8'b00000000; // 3723 :   0 - 0x0
      12'hE8C: dout <= 8'b11111111; // 3724 : 255 - 0xff
      12'hE8D: dout <= 8'b11111111; // 3725 : 255 - 0xff
      12'hE8E: dout <= 8'b11111111; // 3726 : 255 - 0xff
      12'hE8F: dout <= 8'b11111111; // 3727 : 255 - 0xff
      12'hE90: dout <= 8'b11110110; // 3728 : 246 - 0xf6 -- Background 0xe9
      12'hE91: dout <= 8'b11110110; // 3729 : 246 - 0xf6
      12'hE92: dout <= 8'b11110110; // 3730 : 246 - 0xf6
      12'hE93: dout <= 8'b11110110; // 3731 : 246 - 0xf6
      12'hE94: dout <= 8'b11110110; // 3732 : 246 - 0xf6
      12'hE95: dout <= 8'b11110110; // 3733 : 246 - 0xf6
      12'hE96: dout <= 8'b11110110; // 3734 : 246 - 0xf6
      12'hE97: dout <= 8'b11110110; // 3735 : 246 - 0xf6
      12'hE98: dout <= 8'b11110000; // 3736 : 240 - 0xf0 -- plane 1
      12'hE99: dout <= 8'b11110000; // 3737 : 240 - 0xf0
      12'hE9A: dout <= 8'b11110000; // 3738 : 240 - 0xf0
      12'hE9B: dout <= 8'b11110000; // 3739 : 240 - 0xf0
      12'hE9C: dout <= 8'b11110000; // 3740 : 240 - 0xf0
      12'hE9D: dout <= 8'b11110000; // 3741 : 240 - 0xf0
      12'hE9E: dout <= 8'b11110000; // 3742 : 240 - 0xf0
      12'hE9F: dout <= 8'b11110000; // 3743 : 240 - 0xf0
      12'hEA0: dout <= 8'b11111111; // 3744 : 255 - 0xff -- Background 0xea
      12'hEA1: dout <= 8'b11111111; // 3745 : 255 - 0xff
      12'hEA2: dout <= 8'b11111111; // 3746 : 255 - 0xff
      12'hEA3: dout <= 8'b11111111; // 3747 : 255 - 0xff
      12'hEA4: dout <= 8'b00000000; // 3748 :   0 - 0x0
      12'hEA5: dout <= 8'b11111111; // 3749 : 255 - 0xff
      12'hEA6: dout <= 8'b11111111; // 3750 : 255 - 0xff
      12'hEA7: dout <= 8'b00000000; // 3751 :   0 - 0x0
      12'hEA8: dout <= 8'b11111111; // 3752 : 255 - 0xff -- plane 1
      12'hEA9: dout <= 8'b11111111; // 3753 : 255 - 0xff
      12'hEAA: dout <= 8'b11111111; // 3754 : 255 - 0xff
      12'hEAB: dout <= 8'b11111111; // 3755 : 255 - 0xff
      12'hEAC: dout <= 8'b00000000; // 3756 :   0 - 0x0
      12'hEAD: dout <= 8'b00000000; // 3757 :   0 - 0x0
      12'hEAE: dout <= 8'b00000000; // 3758 :   0 - 0x0
      12'hEAF: dout <= 8'b00000000; // 3759 :   0 - 0x0
      12'hEB0: dout <= 8'b01101111; // 3760 : 111 - 0x6f -- Background 0xeb
      12'hEB1: dout <= 8'b01101111; // 3761 : 111 - 0x6f
      12'hEB2: dout <= 8'b01101111; // 3762 : 111 - 0x6f
      12'hEB3: dout <= 8'b01101111; // 3763 : 111 - 0x6f
      12'hEB4: dout <= 8'b01101111; // 3764 : 111 - 0x6f
      12'hEB5: dout <= 8'b01101111; // 3765 : 111 - 0x6f
      12'hEB6: dout <= 8'b01101111; // 3766 : 111 - 0x6f
      12'hEB7: dout <= 8'b01101111; // 3767 : 111 - 0x6f
      12'hEB8: dout <= 8'b00001111; // 3768 :  15 - 0xf -- plane 1
      12'hEB9: dout <= 8'b00001111; // 3769 :  15 - 0xf
      12'hEBA: dout <= 8'b00001111; // 3770 :  15 - 0xf
      12'hEBB: dout <= 8'b00001111; // 3771 :  15 - 0xf
      12'hEBC: dout <= 8'b00001111; // 3772 :  15 - 0xf
      12'hEBD: dout <= 8'b00001111; // 3773 :  15 - 0xf
      12'hEBE: dout <= 8'b00001111; // 3774 :  15 - 0xf
      12'hEBF: dout <= 8'b00001111; // 3775 :  15 - 0xf
      12'hEC0: dout <= 8'b00000000; // 3776 :   0 - 0x0 -- Background 0xec
      12'hEC1: dout <= 8'b00000000; // 3777 :   0 - 0x0
      12'hEC2: dout <= 8'b00000000; // 3778 :   0 - 0x0
      12'hEC3: dout <= 8'b00000000; // 3779 :   0 - 0x0
      12'hEC4: dout <= 8'b00000000; // 3780 :   0 - 0x0
      12'hEC5: dout <= 8'b00000000; // 3781 :   0 - 0x0
      12'hEC6: dout <= 8'b00000000; // 3782 :   0 - 0x0
      12'hEC7: dout <= 8'b00000000; // 3783 :   0 - 0x0
      12'hEC8: dout <= 8'b00000000; // 3784 :   0 - 0x0 -- plane 1
      12'hEC9: dout <= 8'b00000000; // 3785 :   0 - 0x0
      12'hECA: dout <= 8'b00000000; // 3786 :   0 - 0x0
      12'hECB: dout <= 8'b00000000; // 3787 :   0 - 0x0
      12'hECC: dout <= 8'b00000000; // 3788 :   0 - 0x0
      12'hECD: dout <= 8'b00000000; // 3789 :   0 - 0x0
      12'hECE: dout <= 8'b00000000; // 3790 :   0 - 0x0
      12'hECF: dout <= 8'b00000000; // 3791 :   0 - 0x0
      12'hED0: dout <= 8'b00000000; // 3792 :   0 - 0x0 -- Background 0xed
      12'hED1: dout <= 8'b00000000; // 3793 :   0 - 0x0
      12'hED2: dout <= 8'b00000000; // 3794 :   0 - 0x0
      12'hED3: dout <= 8'b00000000; // 3795 :   0 - 0x0
      12'hED4: dout <= 8'b00000000; // 3796 :   0 - 0x0
      12'hED5: dout <= 8'b00000000; // 3797 :   0 - 0x0
      12'hED6: dout <= 8'b00000000; // 3798 :   0 - 0x0
      12'hED7: dout <= 8'b00000000; // 3799 :   0 - 0x0
      12'hED8: dout <= 8'b00000000; // 3800 :   0 - 0x0 -- plane 1
      12'hED9: dout <= 8'b00000000; // 3801 :   0 - 0x0
      12'hEDA: dout <= 8'b00000000; // 3802 :   0 - 0x0
      12'hEDB: dout <= 8'b00000000; // 3803 :   0 - 0x0
      12'hEDC: dout <= 8'b00000000; // 3804 :   0 - 0x0
      12'hEDD: dout <= 8'b00000000; // 3805 :   0 - 0x0
      12'hEDE: dout <= 8'b00000000; // 3806 :   0 - 0x0
      12'hEDF: dout <= 8'b00000000; // 3807 :   0 - 0x0
      12'hEE0: dout <= 8'b00000000; // 3808 :   0 - 0x0 -- Background 0xee
      12'hEE1: dout <= 8'b00000000; // 3809 :   0 - 0x0
      12'hEE2: dout <= 8'b00000000; // 3810 :   0 - 0x0
      12'hEE3: dout <= 8'b00000000; // 3811 :   0 - 0x0
      12'hEE4: dout <= 8'b00000000; // 3812 :   0 - 0x0
      12'hEE5: dout <= 8'b00000000; // 3813 :   0 - 0x0
      12'hEE6: dout <= 8'b00000000; // 3814 :   0 - 0x0
      12'hEE7: dout <= 8'b00000000; // 3815 :   0 - 0x0
      12'hEE8: dout <= 8'b00000000; // 3816 :   0 - 0x0 -- plane 1
      12'hEE9: dout <= 8'b00000000; // 3817 :   0 - 0x0
      12'hEEA: dout <= 8'b00000000; // 3818 :   0 - 0x0
      12'hEEB: dout <= 8'b00000000; // 3819 :   0 - 0x0
      12'hEEC: dout <= 8'b00000000; // 3820 :   0 - 0x0
      12'hEED: dout <= 8'b00000000; // 3821 :   0 - 0x0
      12'hEEE: dout <= 8'b00000000; // 3822 :   0 - 0x0
      12'hEEF: dout <= 8'b00000000; // 3823 :   0 - 0x0
      12'hEF0: dout <= 8'b00000000; // 3824 :   0 - 0x0 -- Background 0xef
      12'hEF1: dout <= 8'b00000000; // 3825 :   0 - 0x0
      12'hEF2: dout <= 8'b00000000; // 3826 :   0 - 0x0
      12'hEF3: dout <= 8'b00000000; // 3827 :   0 - 0x0
      12'hEF4: dout <= 8'b00000000; // 3828 :   0 - 0x0
      12'hEF5: dout <= 8'b00000000; // 3829 :   0 - 0x0
      12'hEF6: dout <= 8'b00000000; // 3830 :   0 - 0x0
      12'hEF7: dout <= 8'b00000000; // 3831 :   0 - 0x0
      12'hEF8: dout <= 8'b00000000; // 3832 :   0 - 0x0 -- plane 1
      12'hEF9: dout <= 8'b00000000; // 3833 :   0 - 0x0
      12'hEFA: dout <= 8'b00000000; // 3834 :   0 - 0x0
      12'hEFB: dout <= 8'b00000000; // 3835 :   0 - 0x0
      12'hEFC: dout <= 8'b00000000; // 3836 :   0 - 0x0
      12'hEFD: dout <= 8'b00000000; // 3837 :   0 - 0x0
      12'hEFE: dout <= 8'b00000000; // 3838 :   0 - 0x0
      12'hEFF: dout <= 8'b00000000; // 3839 :   0 - 0x0
      12'hF00: dout <= 8'b11111111; // 3840 : 255 - 0xff -- Background 0xf0
      12'hF01: dout <= 8'b11111111; // 3841 : 255 - 0xff
      12'hF02: dout <= 8'b11111111; // 3842 : 255 - 0xff
      12'hF03: dout <= 8'b11111111; // 3843 : 255 - 0xff
      12'hF04: dout <= 8'b11111111; // 3844 : 255 - 0xff
      12'hF05: dout <= 8'b11111111; // 3845 : 255 - 0xff
      12'hF06: dout <= 8'b11111111; // 3846 : 255 - 0xff
      12'hF07: dout <= 8'b11111111; // 3847 : 255 - 0xff
      12'hF08: dout <= 8'b11111111; // 3848 : 255 - 0xff -- plane 1
      12'hF09: dout <= 8'b11111111; // 3849 : 255 - 0xff
      12'hF0A: dout <= 8'b11111111; // 3850 : 255 - 0xff
      12'hF0B: dout <= 8'b11111111; // 3851 : 255 - 0xff
      12'hF0C: dout <= 8'b11111111; // 3852 : 255 - 0xff
      12'hF0D: dout <= 8'b11111111; // 3853 : 255 - 0xff
      12'hF0E: dout <= 8'b11111111; // 3854 : 255 - 0xff
      12'hF0F: dout <= 8'b11111111; // 3855 : 255 - 0xff
      12'hF10: dout <= 8'b11111111; // 3856 : 255 - 0xff -- Background 0xf1
      12'hF11: dout <= 8'b11111111; // 3857 : 255 - 0xff
      12'hF12: dout <= 8'b11111111; // 3858 : 255 - 0xff
      12'hF13: dout <= 8'b11111111; // 3859 : 255 - 0xff
      12'hF14: dout <= 8'b11111111; // 3860 : 255 - 0xff
      12'hF15: dout <= 8'b11111111; // 3861 : 255 - 0xff
      12'hF16: dout <= 8'b11111111; // 3862 : 255 - 0xff
      12'hF17: dout <= 8'b11111111; // 3863 : 255 - 0xff
      12'hF18: dout <= 8'b11111111; // 3864 : 255 - 0xff -- plane 1
      12'hF19: dout <= 8'b11111111; // 3865 : 255 - 0xff
      12'hF1A: dout <= 8'b11111111; // 3866 : 255 - 0xff
      12'hF1B: dout <= 8'b11111111; // 3867 : 255 - 0xff
      12'hF1C: dout <= 8'b11111111; // 3868 : 255 - 0xff
      12'hF1D: dout <= 8'b11111111; // 3869 : 255 - 0xff
      12'hF1E: dout <= 8'b11111111; // 3870 : 255 - 0xff
      12'hF1F: dout <= 8'b11111111; // 3871 : 255 - 0xff
      12'hF20: dout <= 8'b11111111; // 3872 : 255 - 0xff -- Background 0xf2
      12'hF21: dout <= 8'b11111111; // 3873 : 255 - 0xff
      12'hF22: dout <= 8'b11111111; // 3874 : 255 - 0xff
      12'hF23: dout <= 8'b11111111; // 3875 : 255 - 0xff
      12'hF24: dout <= 8'b11111111; // 3876 : 255 - 0xff
      12'hF25: dout <= 8'b11111111; // 3877 : 255 - 0xff
      12'hF26: dout <= 8'b11111111; // 3878 : 255 - 0xff
      12'hF27: dout <= 8'b11111111; // 3879 : 255 - 0xff
      12'hF28: dout <= 8'b11111111; // 3880 : 255 - 0xff -- plane 1
      12'hF29: dout <= 8'b11111111; // 3881 : 255 - 0xff
      12'hF2A: dout <= 8'b11111111; // 3882 : 255 - 0xff
      12'hF2B: dout <= 8'b11111111; // 3883 : 255 - 0xff
      12'hF2C: dout <= 8'b11111111; // 3884 : 255 - 0xff
      12'hF2D: dout <= 8'b11111111; // 3885 : 255 - 0xff
      12'hF2E: dout <= 8'b11111111; // 3886 : 255 - 0xff
      12'hF2F: dout <= 8'b11111111; // 3887 : 255 - 0xff
      12'hF30: dout <= 8'b11111111; // 3888 : 255 - 0xff -- Background 0xf3
      12'hF31: dout <= 8'b11111111; // 3889 : 255 - 0xff
      12'hF32: dout <= 8'b11111111; // 3890 : 255 - 0xff
      12'hF33: dout <= 8'b11111111; // 3891 : 255 - 0xff
      12'hF34: dout <= 8'b11111111; // 3892 : 255 - 0xff
      12'hF35: dout <= 8'b11111111; // 3893 : 255 - 0xff
      12'hF36: dout <= 8'b11111111; // 3894 : 255 - 0xff
      12'hF37: dout <= 8'b11111111; // 3895 : 255 - 0xff
      12'hF38: dout <= 8'b11111111; // 3896 : 255 - 0xff -- plane 1
      12'hF39: dout <= 8'b11111111; // 3897 : 255 - 0xff
      12'hF3A: dout <= 8'b11111111; // 3898 : 255 - 0xff
      12'hF3B: dout <= 8'b11111111; // 3899 : 255 - 0xff
      12'hF3C: dout <= 8'b11111111; // 3900 : 255 - 0xff
      12'hF3D: dout <= 8'b11111111; // 3901 : 255 - 0xff
      12'hF3E: dout <= 8'b11111111; // 3902 : 255 - 0xff
      12'hF3F: dout <= 8'b11111111; // 3903 : 255 - 0xff
      12'hF40: dout <= 8'b11111111; // 3904 : 255 - 0xff -- Background 0xf4
      12'hF41: dout <= 8'b11111111; // 3905 : 255 - 0xff
      12'hF42: dout <= 8'b11111111; // 3906 : 255 - 0xff
      12'hF43: dout <= 8'b11111111; // 3907 : 255 - 0xff
      12'hF44: dout <= 8'b11111111; // 3908 : 255 - 0xff
      12'hF45: dout <= 8'b11111111; // 3909 : 255 - 0xff
      12'hF46: dout <= 8'b11111111; // 3910 : 255 - 0xff
      12'hF47: dout <= 8'b11111111; // 3911 : 255 - 0xff
      12'hF48: dout <= 8'b11111111; // 3912 : 255 - 0xff -- plane 1
      12'hF49: dout <= 8'b11111111; // 3913 : 255 - 0xff
      12'hF4A: dout <= 8'b11111111; // 3914 : 255 - 0xff
      12'hF4B: dout <= 8'b11111111; // 3915 : 255 - 0xff
      12'hF4C: dout <= 8'b11111111; // 3916 : 255 - 0xff
      12'hF4D: dout <= 8'b11111111; // 3917 : 255 - 0xff
      12'hF4E: dout <= 8'b11111111; // 3918 : 255 - 0xff
      12'hF4F: dout <= 8'b11111111; // 3919 : 255 - 0xff
      12'hF50: dout <= 8'b11111111; // 3920 : 255 - 0xff -- Background 0xf5
      12'hF51: dout <= 8'b11111111; // 3921 : 255 - 0xff
      12'hF52: dout <= 8'b11111111; // 3922 : 255 - 0xff
      12'hF53: dout <= 8'b11111111; // 3923 : 255 - 0xff
      12'hF54: dout <= 8'b11111111; // 3924 : 255 - 0xff
      12'hF55: dout <= 8'b11111111; // 3925 : 255 - 0xff
      12'hF56: dout <= 8'b11111111; // 3926 : 255 - 0xff
      12'hF57: dout <= 8'b11111111; // 3927 : 255 - 0xff
      12'hF58: dout <= 8'b11111111; // 3928 : 255 - 0xff -- plane 1
      12'hF59: dout <= 8'b11111111; // 3929 : 255 - 0xff
      12'hF5A: dout <= 8'b11111111; // 3930 : 255 - 0xff
      12'hF5B: dout <= 8'b11111111; // 3931 : 255 - 0xff
      12'hF5C: dout <= 8'b11111111; // 3932 : 255 - 0xff
      12'hF5D: dout <= 8'b11111111; // 3933 : 255 - 0xff
      12'hF5E: dout <= 8'b11111111; // 3934 : 255 - 0xff
      12'hF5F: dout <= 8'b11111111; // 3935 : 255 - 0xff
      12'hF60: dout <= 8'b11111111; // 3936 : 255 - 0xff -- Background 0xf6
      12'hF61: dout <= 8'b11111111; // 3937 : 255 - 0xff
      12'hF62: dout <= 8'b11111111; // 3938 : 255 - 0xff
      12'hF63: dout <= 8'b11111111; // 3939 : 255 - 0xff
      12'hF64: dout <= 8'b11111111; // 3940 : 255 - 0xff
      12'hF65: dout <= 8'b11111111; // 3941 : 255 - 0xff
      12'hF66: dout <= 8'b11111111; // 3942 : 255 - 0xff
      12'hF67: dout <= 8'b11111111; // 3943 : 255 - 0xff
      12'hF68: dout <= 8'b11111111; // 3944 : 255 - 0xff -- plane 1
      12'hF69: dout <= 8'b11111111; // 3945 : 255 - 0xff
      12'hF6A: dout <= 8'b11111111; // 3946 : 255 - 0xff
      12'hF6B: dout <= 8'b11111111; // 3947 : 255 - 0xff
      12'hF6C: dout <= 8'b11111111; // 3948 : 255 - 0xff
      12'hF6D: dout <= 8'b11111111; // 3949 : 255 - 0xff
      12'hF6E: dout <= 8'b11111111; // 3950 : 255 - 0xff
      12'hF6F: dout <= 8'b11111111; // 3951 : 255 - 0xff
      12'hF70: dout <= 8'b11111111; // 3952 : 255 - 0xff -- Background 0xf7
      12'hF71: dout <= 8'b11111111; // 3953 : 255 - 0xff
      12'hF72: dout <= 8'b11111111; // 3954 : 255 - 0xff
      12'hF73: dout <= 8'b11111111; // 3955 : 255 - 0xff
      12'hF74: dout <= 8'b11111111; // 3956 : 255 - 0xff
      12'hF75: dout <= 8'b11111111; // 3957 : 255 - 0xff
      12'hF76: dout <= 8'b11111111; // 3958 : 255 - 0xff
      12'hF77: dout <= 8'b11111111; // 3959 : 255 - 0xff
      12'hF78: dout <= 8'b11111111; // 3960 : 255 - 0xff -- plane 1
      12'hF79: dout <= 8'b11111111; // 3961 : 255 - 0xff
      12'hF7A: dout <= 8'b11111111; // 3962 : 255 - 0xff
      12'hF7B: dout <= 8'b11111111; // 3963 : 255 - 0xff
      12'hF7C: dout <= 8'b11111111; // 3964 : 255 - 0xff
      12'hF7D: dout <= 8'b11111111; // 3965 : 255 - 0xff
      12'hF7E: dout <= 8'b11111111; // 3966 : 255 - 0xff
      12'hF7F: dout <= 8'b11111111; // 3967 : 255 - 0xff
      12'hF80: dout <= 8'b11111111; // 3968 : 255 - 0xff -- Background 0xf8
      12'hF81: dout <= 8'b11111111; // 3969 : 255 - 0xff
      12'hF82: dout <= 8'b11111111; // 3970 : 255 - 0xff
      12'hF83: dout <= 8'b11111111; // 3971 : 255 - 0xff
      12'hF84: dout <= 8'b11111111; // 3972 : 255 - 0xff
      12'hF85: dout <= 8'b11111111; // 3973 : 255 - 0xff
      12'hF86: dout <= 8'b11111111; // 3974 : 255 - 0xff
      12'hF87: dout <= 8'b11111111; // 3975 : 255 - 0xff
      12'hF88: dout <= 8'b11111111; // 3976 : 255 - 0xff -- plane 1
      12'hF89: dout <= 8'b11111111; // 3977 : 255 - 0xff
      12'hF8A: dout <= 8'b11111111; // 3978 : 255 - 0xff
      12'hF8B: dout <= 8'b11111111; // 3979 : 255 - 0xff
      12'hF8C: dout <= 8'b11111111; // 3980 : 255 - 0xff
      12'hF8D: dout <= 8'b11111111; // 3981 : 255 - 0xff
      12'hF8E: dout <= 8'b11111111; // 3982 : 255 - 0xff
      12'hF8F: dout <= 8'b11111111; // 3983 : 255 - 0xff
      12'hF90: dout <= 8'b11111111; // 3984 : 255 - 0xff -- Background 0xf9
      12'hF91: dout <= 8'b11111111; // 3985 : 255 - 0xff
      12'hF92: dout <= 8'b11111111; // 3986 : 255 - 0xff
      12'hF93: dout <= 8'b11111111; // 3987 : 255 - 0xff
      12'hF94: dout <= 8'b11111111; // 3988 : 255 - 0xff
      12'hF95: dout <= 8'b11111111; // 3989 : 255 - 0xff
      12'hF96: dout <= 8'b11111111; // 3990 : 255 - 0xff
      12'hF97: dout <= 8'b11111111; // 3991 : 255 - 0xff
      12'hF98: dout <= 8'b11111111; // 3992 : 255 - 0xff -- plane 1
      12'hF99: dout <= 8'b11111111; // 3993 : 255 - 0xff
      12'hF9A: dout <= 8'b11111111; // 3994 : 255 - 0xff
      12'hF9B: dout <= 8'b11111111; // 3995 : 255 - 0xff
      12'hF9C: dout <= 8'b11111111; // 3996 : 255 - 0xff
      12'hF9D: dout <= 8'b11111111; // 3997 : 255 - 0xff
      12'hF9E: dout <= 8'b11111111; // 3998 : 255 - 0xff
      12'hF9F: dout <= 8'b11111111; // 3999 : 255 - 0xff
      12'hFA0: dout <= 8'b11111111; // 4000 : 255 - 0xff -- Background 0xfa
      12'hFA1: dout <= 8'b11111111; // 4001 : 255 - 0xff
      12'hFA2: dout <= 8'b11111111; // 4002 : 255 - 0xff
      12'hFA3: dout <= 8'b11111111; // 4003 : 255 - 0xff
      12'hFA4: dout <= 8'b11111111; // 4004 : 255 - 0xff
      12'hFA5: dout <= 8'b11111111; // 4005 : 255 - 0xff
      12'hFA6: dout <= 8'b11111111; // 4006 : 255 - 0xff
      12'hFA7: dout <= 8'b11111111; // 4007 : 255 - 0xff
      12'hFA8: dout <= 8'b11111111; // 4008 : 255 - 0xff -- plane 1
      12'hFA9: dout <= 8'b11111111; // 4009 : 255 - 0xff
      12'hFAA: dout <= 8'b11111111; // 4010 : 255 - 0xff
      12'hFAB: dout <= 8'b11111111; // 4011 : 255 - 0xff
      12'hFAC: dout <= 8'b11111111; // 4012 : 255 - 0xff
      12'hFAD: dout <= 8'b11111111; // 4013 : 255 - 0xff
      12'hFAE: dout <= 8'b11111111; // 4014 : 255 - 0xff
      12'hFAF: dout <= 8'b11111111; // 4015 : 255 - 0xff
      12'hFB0: dout <= 8'b11111111; // 4016 : 255 - 0xff -- Background 0xfb
      12'hFB1: dout <= 8'b11111111; // 4017 : 255 - 0xff
      12'hFB2: dout <= 8'b11111111; // 4018 : 255 - 0xff
      12'hFB3: dout <= 8'b11111111; // 4019 : 255 - 0xff
      12'hFB4: dout <= 8'b11111111; // 4020 : 255 - 0xff
      12'hFB5: dout <= 8'b11111111; // 4021 : 255 - 0xff
      12'hFB6: dout <= 8'b11111111; // 4022 : 255 - 0xff
      12'hFB7: dout <= 8'b11111111; // 4023 : 255 - 0xff
      12'hFB8: dout <= 8'b11111111; // 4024 : 255 - 0xff -- plane 1
      12'hFB9: dout <= 8'b11111111; // 4025 : 255 - 0xff
      12'hFBA: dout <= 8'b11111111; // 4026 : 255 - 0xff
      12'hFBB: dout <= 8'b11111111; // 4027 : 255 - 0xff
      12'hFBC: dout <= 8'b11111111; // 4028 : 255 - 0xff
      12'hFBD: dout <= 8'b11111111; // 4029 : 255 - 0xff
      12'hFBE: dout <= 8'b11111111; // 4030 : 255 - 0xff
      12'hFBF: dout <= 8'b11111111; // 4031 : 255 - 0xff
      12'hFC0: dout <= 8'b11111111; // 4032 : 255 - 0xff -- Background 0xfc
      12'hFC1: dout <= 8'b11111111; // 4033 : 255 - 0xff
      12'hFC2: dout <= 8'b11111111; // 4034 : 255 - 0xff
      12'hFC3: dout <= 8'b11111111; // 4035 : 255 - 0xff
      12'hFC4: dout <= 8'b11111111; // 4036 : 255 - 0xff
      12'hFC5: dout <= 8'b11111111; // 4037 : 255 - 0xff
      12'hFC6: dout <= 8'b11111111; // 4038 : 255 - 0xff
      12'hFC7: dout <= 8'b11111111; // 4039 : 255 - 0xff
      12'hFC8: dout <= 8'b11111111; // 4040 : 255 - 0xff -- plane 1
      12'hFC9: dout <= 8'b11111111; // 4041 : 255 - 0xff
      12'hFCA: dout <= 8'b11111111; // 4042 : 255 - 0xff
      12'hFCB: dout <= 8'b11111111; // 4043 : 255 - 0xff
      12'hFCC: dout <= 8'b11111111; // 4044 : 255 - 0xff
      12'hFCD: dout <= 8'b11111111; // 4045 : 255 - 0xff
      12'hFCE: dout <= 8'b11111111; // 4046 : 255 - 0xff
      12'hFCF: dout <= 8'b11111111; // 4047 : 255 - 0xff
      12'hFD0: dout <= 8'b11111111; // 4048 : 255 - 0xff -- Background 0xfd
      12'hFD1: dout <= 8'b11111111; // 4049 : 255 - 0xff
      12'hFD2: dout <= 8'b11111111; // 4050 : 255 - 0xff
      12'hFD3: dout <= 8'b11111111; // 4051 : 255 - 0xff
      12'hFD4: dout <= 8'b11111111; // 4052 : 255 - 0xff
      12'hFD5: dout <= 8'b11111111; // 4053 : 255 - 0xff
      12'hFD6: dout <= 8'b11111111; // 4054 : 255 - 0xff
      12'hFD7: dout <= 8'b11111111; // 4055 : 255 - 0xff
      12'hFD8: dout <= 8'b11111111; // 4056 : 255 - 0xff -- plane 1
      12'hFD9: dout <= 8'b11111111; // 4057 : 255 - 0xff
      12'hFDA: dout <= 8'b11111111; // 4058 : 255 - 0xff
      12'hFDB: dout <= 8'b11111111; // 4059 : 255 - 0xff
      12'hFDC: dout <= 8'b11111111; // 4060 : 255 - 0xff
      12'hFDD: dout <= 8'b11111111; // 4061 : 255 - 0xff
      12'hFDE: dout <= 8'b11111111; // 4062 : 255 - 0xff
      12'hFDF: dout <= 8'b11111111; // 4063 : 255 - 0xff
      12'hFE0: dout <= 8'b11111111; // 4064 : 255 - 0xff -- Background 0xfe
      12'hFE1: dout <= 8'b11111111; // 4065 : 255 - 0xff
      12'hFE2: dout <= 8'b11111111; // 4066 : 255 - 0xff
      12'hFE3: dout <= 8'b11111111; // 4067 : 255 - 0xff
      12'hFE4: dout <= 8'b11111111; // 4068 : 255 - 0xff
      12'hFE5: dout <= 8'b11111111; // 4069 : 255 - 0xff
      12'hFE6: dout <= 8'b11111111; // 4070 : 255 - 0xff
      12'hFE7: dout <= 8'b11111111; // 4071 : 255 - 0xff
      12'hFE8: dout <= 8'b11111111; // 4072 : 255 - 0xff -- plane 1
      12'hFE9: dout <= 8'b11111111; // 4073 : 255 - 0xff
      12'hFEA: dout <= 8'b11111111; // 4074 : 255 - 0xff
      12'hFEB: dout <= 8'b11111111; // 4075 : 255 - 0xff
      12'hFEC: dout <= 8'b11111111; // 4076 : 255 - 0xff
      12'hFED: dout <= 8'b11111111; // 4077 : 255 - 0xff
      12'hFEE: dout <= 8'b11111111; // 4078 : 255 - 0xff
      12'hFEF: dout <= 8'b11111111; // 4079 : 255 - 0xff
      12'hFF0: dout <= 8'b11111111; // 4080 : 255 - 0xff -- Background 0xff
      12'hFF1: dout <= 8'b11111111; // 4081 : 255 - 0xff
      12'hFF2: dout <= 8'b11111111; // 4082 : 255 - 0xff
      12'hFF3: dout <= 8'b11111111; // 4083 : 255 - 0xff
      12'hFF4: dout <= 8'b11111111; // 4084 : 255 - 0xff
      12'hFF5: dout <= 8'b11111111; // 4085 : 255 - 0xff
      12'hFF6: dout <= 8'b11111111; // 4086 : 255 - 0xff
      12'hFF7: dout <= 8'b11111111; // 4087 : 255 - 0xff
      12'hFF8: dout <= 8'b11111111; // 4088 : 255 - 0xff -- plane 1
      12'hFF9: dout <= 8'b11111111; // 4089 : 255 - 0xff
      12'hFFA: dout <= 8'b11111111; // 4090 : 255 - 0xff
      12'hFFB: dout <= 8'b11111111; // 4091 : 255 - 0xff
      12'hFFC: dout <= 8'b11111111; // 4092 : 255 - 0xff
      12'hFFD: dout <= 8'b11111111; // 4093 : 255 - 0xff
      12'hFFE: dout <= 8'b11111111; // 4094 : 255 - 0xff
      12'hFFF: dout <= 8'b11111111; // 4095 : 255 - 0xff
    endcase
  end

endmodule
