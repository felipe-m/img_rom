//-   Sprites Pattern table COLOR PLANE 0
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
//- Autcmatically generated verilog ROM from a NES memory file----


//-  Original memory dump file name: nova_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_PTABLE_NOVA_SPR_PLN0
  (
     input     clk,   // clock
     input      [11-1:0] addr,  //2048 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Sprite pattern Table COLOR PLANE 0
      11'h0: dout <= 8'b11111111; //    0 : 255 - 0xff -- Sprite 0x0
      11'h1: dout <= 8'b11111111; //    1 : 255 - 0xff
      11'h2: dout <= 8'b11000000; //    2 : 192 - 0xc0
      11'h3: dout <= 8'b11000000; //    3 : 192 - 0xc0
      11'h4: dout <= 8'b11000000; //    4 : 192 - 0xc0
      11'h5: dout <= 8'b11000000; //    5 : 192 - 0xc0
      11'h6: dout <= 8'b11010101; //    6 : 213 - 0xd5
      11'h7: dout <= 8'b11111111; //    7 : 255 - 0xff
      11'h8: dout <= 8'b11111111; //    8 : 255 - 0xff -- Sprite 0x1
      11'h9: dout <= 8'b11111111; //    9 : 255 - 0xff
      11'hA: dout <= 8'b11001110; //   10 : 206 - 0xce
      11'hB: dout <= 8'b11000110; //   11 : 198 - 0xc6
      11'hC: dout <= 8'b11001110; //   12 : 206 - 0xce
      11'hD: dout <= 8'b11000110; //   13 : 198 - 0xc6
      11'hE: dout <= 8'b11101110; //   14 : 238 - 0xee
      11'hF: dout <= 8'b11111111; //   15 : 255 - 0xff
      11'h10: dout <= 8'b11111111; //   16 : 255 - 0xff -- Sprite 0x2
      11'h11: dout <= 8'b11111111; //   17 : 255 - 0xff
      11'h12: dout <= 8'b01110001; //   18 : 113 - 0x71
      11'h13: dout <= 8'b00110011; //   19 :  51 - 0x33
      11'h14: dout <= 8'b01110001; //   20 : 113 - 0x71
      11'h15: dout <= 8'b00110011; //   21 :  51 - 0x33
      11'h16: dout <= 8'b01110101; //   22 : 117 - 0x75
      11'h17: dout <= 8'b11111111; //   23 : 255 - 0xff
      11'h18: dout <= 8'b11111111; //   24 : 255 - 0xff -- Sprite 0x3
      11'h19: dout <= 8'b11111111; //   25 : 255 - 0xff
      11'h1A: dout <= 8'b00000011; //   26 :   3 - 0x3
      11'h1B: dout <= 8'b00000001; //   27 :   1 - 0x1
      11'h1C: dout <= 8'b00000011; //   28 :   3 - 0x3
      11'h1D: dout <= 8'b00000001; //   29 :   1 - 0x1
      11'h1E: dout <= 8'b10101011; //   30 : 171 - 0xab
      11'h1F: dout <= 8'b11111111; //   31 : 255 - 0xff
      11'h20: dout <= 8'b11111111; //   32 : 255 - 0xff -- Sprite 0x4
      11'h21: dout <= 8'b11111111; //   33 : 255 - 0xff
      11'h22: dout <= 8'b11100000; //   34 : 224 - 0xe0
      11'h23: dout <= 8'b11000110; //   35 : 198 - 0xc6
      11'h24: dout <= 8'b11000110; //   36 : 198 - 0xc6
      11'h25: dout <= 8'b11110110; //   37 : 246 - 0xf6
      11'h26: dout <= 8'b11110000; //   38 : 240 - 0xf0
      11'h27: dout <= 8'b11110001; //   39 : 241 - 0xf1
      11'h28: dout <= 8'b11000111; //   40 : 199 - 0xc7 -- Sprite 0x5
      11'h29: dout <= 8'b11001111; //   41 : 207 - 0xcf
      11'h2A: dout <= 8'b11011111; //   42 : 223 - 0xdf
      11'h2B: dout <= 8'b11011111; //   43 : 223 - 0xdf
      11'h2C: dout <= 8'b11001110; //   44 : 206 - 0xce
      11'h2D: dout <= 8'b11100000; //   45 : 224 - 0xe0
      11'h2E: dout <= 8'b11111111; //   46 : 255 - 0xff
      11'h2F: dout <= 8'b11111111; //   47 : 255 - 0xff
      11'h30: dout <= 8'b11111111; //   48 : 255 - 0xff -- Sprite 0x6
      11'h31: dout <= 8'b11111111; //   49 : 255 - 0xff
      11'h32: dout <= 8'b00000111; //   50 :   7 - 0x7
      11'h33: dout <= 8'b01100011; //   51 :  99 - 0x63
      11'h34: dout <= 8'b01100011; //   52 :  99 - 0x63
      11'h35: dout <= 8'b01101111; //   53 : 111 - 0x6f
      11'h36: dout <= 8'b00001111; //   54 :  15 - 0xf
      11'h37: dout <= 8'b10001111; //   55 : 143 - 0x8f
      11'h38: dout <= 8'b11100011; //   56 : 227 - 0xe3 -- Sprite 0x7
      11'h39: dout <= 8'b11110011; //   57 : 243 - 0xf3
      11'h3A: dout <= 8'b11111011; //   58 : 251 - 0xfb
      11'h3B: dout <= 8'b11111011; //   59 : 251 - 0xfb
      11'h3C: dout <= 8'b01110011; //   60 : 115 - 0x73
      11'h3D: dout <= 8'b00000111; //   61 :   7 - 0x7
      11'h3E: dout <= 8'b11111111; //   62 : 255 - 0xff
      11'h3F: dout <= 8'b11111111; //   63 : 255 - 0xff
      11'h40: dout <= 8'b11111111; //   64 : 255 - 0xff -- Sprite 0x8
      11'h41: dout <= 8'b11010101; //   65 : 213 - 0xd5
      11'h42: dout <= 8'b10101010; //   66 : 170 - 0xaa
      11'h43: dout <= 8'b11010101; //   67 : 213 - 0xd5
      11'h44: dout <= 8'b10101010; //   68 : 170 - 0xaa
      11'h45: dout <= 8'b11010101; //   69 : 213 - 0xd5
      11'h46: dout <= 8'b10101010; //   70 : 170 - 0xaa
      11'h47: dout <= 8'b11010101; //   71 : 213 - 0xd5
      11'h48: dout <= 8'b10101010; //   72 : 170 - 0xaa -- Sprite 0x9
      11'h49: dout <= 8'b11010101; //   73 : 213 - 0xd5
      11'h4A: dout <= 8'b10101010; //   74 : 170 - 0xaa
      11'h4B: dout <= 8'b11010101; //   75 : 213 - 0xd5
      11'h4C: dout <= 8'b10101010; //   76 : 170 - 0xaa
      11'h4D: dout <= 8'b11110101; //   77 : 245 - 0xf5
      11'h4E: dout <= 8'b10101010; //   78 : 170 - 0xaa
      11'h4F: dout <= 8'b11111111; //   79 : 255 - 0xff
      11'h50: dout <= 8'b11111111; //   80 : 255 - 0xff -- Sprite 0xa
      11'h51: dout <= 8'b01010101; //   81 :  85 - 0x55
      11'h52: dout <= 8'b10101111; //   82 : 175 - 0xaf
      11'h53: dout <= 8'b01010101; //   83 :  85 - 0x55
      11'h54: dout <= 8'b10101011; //   84 : 171 - 0xab
      11'h55: dout <= 8'b01010101; //   85 :  85 - 0x55
      11'h56: dout <= 8'b10101011; //   86 : 171 - 0xab
      11'h57: dout <= 8'b01010101; //   87 :  85 - 0x55
      11'h58: dout <= 8'b10101011; //   88 : 171 - 0xab -- Sprite 0xb
      11'h59: dout <= 8'b01010101; //   89 :  85 - 0x55
      11'h5A: dout <= 8'b10101011; //   90 : 171 - 0xab
      11'h5B: dout <= 8'b01010101; //   91 :  85 - 0x55
      11'h5C: dout <= 8'b10101011; //   92 : 171 - 0xab
      11'h5D: dout <= 8'b01010101; //   93 :  85 - 0x55
      11'h5E: dout <= 8'b10101011; //   94 : 171 - 0xab
      11'h5F: dout <= 8'b11111111; //   95 : 255 - 0xff
      11'h60: dout <= 8'b11111111; //   96 : 255 - 0xff -- Sprite 0xc
      11'h61: dout <= 8'b11010101; //   97 : 213 - 0xd5
      11'h62: dout <= 8'b10100000; //   98 : 160 - 0xa0
      11'h63: dout <= 8'b11010000; //   99 : 208 - 0xd0
      11'h64: dout <= 8'b10001111; //  100 : 143 - 0x8f
      11'h65: dout <= 8'b11001000; //  101 : 200 - 0xc8
      11'h66: dout <= 8'b10001000; //  102 : 136 - 0x88
      11'h67: dout <= 8'b11001000; //  103 : 200 - 0xc8
      11'h68: dout <= 8'b10001000; //  104 : 136 - 0x88 -- Sprite 0xd
      11'h69: dout <= 8'b11001000; //  105 : 200 - 0xc8
      11'h6A: dout <= 8'b10001000; //  106 : 136 - 0x88
      11'h6B: dout <= 8'b11001111; //  107 : 207 - 0xcf
      11'h6C: dout <= 8'b10010000; //  108 : 144 - 0x90
      11'h6D: dout <= 8'b11100000; //  109 : 224 - 0xe0
      11'h6E: dout <= 8'b11101010; //  110 : 234 - 0xea
      11'h6F: dout <= 8'b11111111; //  111 : 255 - 0xff
      11'h70: dout <= 8'b11111111; //  112 : 255 - 0xff -- Sprite 0xe
      11'h71: dout <= 8'b01011011; //  113 :  91 - 0x5b
      11'h72: dout <= 8'b00000111; //  114 :   7 - 0x7
      11'h73: dout <= 8'b00001001; //  115 :   9 - 0x9
      11'h74: dout <= 8'b11110011; //  116 : 243 - 0xf3
      11'h75: dout <= 8'b00010001; //  117 :  17 - 0x11
      11'h76: dout <= 8'b00010011; //  118 :  19 - 0x13
      11'h77: dout <= 8'b00010001; //  119 :  17 - 0x11
      11'h78: dout <= 8'b00010011; //  120 :  19 - 0x13 -- Sprite 0xf
      11'h79: dout <= 8'b00010001; //  121 :  17 - 0x11
      11'h7A: dout <= 8'b00010011; //  122 :  19 - 0x13
      11'h7B: dout <= 8'b11110001; //  123 : 241 - 0xf1
      11'h7C: dout <= 8'b00001011; //  124 :  11 - 0xb
      11'h7D: dout <= 8'b00000101; //  125 :   5 - 0x5
      11'h7E: dout <= 8'b10101011; //  126 : 171 - 0xab
      11'h7F: dout <= 8'b11111111; //  127 : 255 - 0xff
      11'h80: dout <= 8'b11010000; //  128 : 208 - 0xd0 -- Sprite 0x10
      11'h81: dout <= 8'b10010000; //  129 : 144 - 0x90
      11'h82: dout <= 8'b11011111; //  130 : 223 - 0xdf
      11'h83: dout <= 8'b10011010; //  131 : 154 - 0x9a
      11'h84: dout <= 8'b11010101; //  132 : 213 - 0xd5
      11'h85: dout <= 8'b10011111; //  133 : 159 - 0x9f
      11'h86: dout <= 8'b11010000; //  134 : 208 - 0xd0
      11'h87: dout <= 8'b10010000; //  135 : 144 - 0x90
      11'h88: dout <= 8'b00001001; //  136 :   9 - 0x9 -- Sprite 0x11
      11'h89: dout <= 8'b00001011; //  137 :  11 - 0xb
      11'h8A: dout <= 8'b11111001; //  138 : 249 - 0xf9
      11'h8B: dout <= 8'b10101011; //  139 : 171 - 0xab
      11'h8C: dout <= 8'b01011001; //  140 :  89 - 0x59
      11'h8D: dout <= 8'b11111011; //  141 : 251 - 0xfb
      11'h8E: dout <= 8'b00001001; //  142 :   9 - 0x9
      11'h8F: dout <= 8'b00001011; //  143 :  11 - 0xb
      11'h90: dout <= 8'b00011000; //  144 :  24 - 0x18 -- Sprite 0x12
      11'h91: dout <= 8'b00010100; //  145 :  20 - 0x14
      11'h92: dout <= 8'b00010100; //  146 :  20 - 0x14
      11'h93: dout <= 8'b00111010; //  147 :  58 - 0x3a
      11'h94: dout <= 8'b00111010; //  148 :  58 - 0x3a
      11'h95: dout <= 8'b01111010; //  149 : 122 - 0x7a
      11'h96: dout <= 8'b01111010; //  150 : 122 - 0x7a
      11'h97: dout <= 8'b01111010; //  151 : 122 - 0x7a
      11'h98: dout <= 8'b11111011; //  152 : 251 - 0xfb -- Sprite 0x13
      11'h99: dout <= 8'b11111101; //  153 : 253 - 0xfd
      11'h9A: dout <= 8'b11111101; //  154 : 253 - 0xfd
      11'h9B: dout <= 8'b11111101; //  155 : 253 - 0xfd
      11'h9C: dout <= 8'b11111101; //  156 : 253 - 0xfd
      11'h9D: dout <= 8'b11111101; //  157 : 253 - 0xfd
      11'h9E: dout <= 8'b10000001; //  158 : 129 - 0x81
      11'h9F: dout <= 8'b11111111; //  159 : 255 - 0xff
      11'hA0: dout <= 8'b00000000; //  160 :   0 - 0x0 -- Sprite 0x14
      11'hA1: dout <= 8'b00000111; //  161 :   7 - 0x7
      11'hA2: dout <= 8'b00000010; //  162 :   2 - 0x2
      11'hA3: dout <= 8'b00000100; //  163 :   4 - 0x4
      11'hA4: dout <= 8'b00000011; //  164 :   3 - 0x3
      11'hA5: dout <= 8'b00000011; //  165 :   3 - 0x3
      11'hA6: dout <= 8'b00001101; //  166 :  13 - 0xd
      11'hA7: dout <= 8'b00010111; //  167 :  23 - 0x17
      11'hA8: dout <= 8'b00101111; //  168 :  47 - 0x2f -- Sprite 0x15
      11'hA9: dout <= 8'b01001111; //  169 :  79 - 0x4f
      11'hAA: dout <= 8'b01001111; //  170 :  79 - 0x4f
      11'hAB: dout <= 8'b01001111; //  171 :  79 - 0x4f
      11'hAC: dout <= 8'b01001111; //  172 :  79 - 0x4f
      11'hAD: dout <= 8'b00100111; //  173 :  39 - 0x27
      11'hAE: dout <= 8'b00010000; //  174 :  16 - 0x10
      11'hAF: dout <= 8'b00001111; //  175 :  15 - 0xf
      11'hB0: dout <= 8'b00000000; //  176 :   0 - 0x0 -- Sprite 0x16
      11'hB1: dout <= 8'b11100000; //  177 : 224 - 0xe0
      11'hB2: dout <= 8'b10100000; //  178 : 160 - 0xa0
      11'hB3: dout <= 8'b00100000; //  179 :  32 - 0x20
      11'hB4: dout <= 8'b11000000; //  180 : 192 - 0xc0
      11'hB5: dout <= 8'b01000000; //  181 :  64 - 0x40
      11'hB6: dout <= 8'b00110000; //  182 :  48 - 0x30
      11'hB7: dout <= 8'b11101000; //  183 : 232 - 0xe8
      11'hB8: dout <= 8'b11110100; //  184 : 244 - 0xf4 -- Sprite 0x17
      11'hB9: dout <= 8'b11110010; //  185 : 242 - 0xf2
      11'hBA: dout <= 8'b11110010; //  186 : 242 - 0xf2
      11'hBB: dout <= 8'b11110010; //  187 : 242 - 0xf2
      11'hBC: dout <= 8'b11110010; //  188 : 242 - 0xf2
      11'hBD: dout <= 8'b11100100; //  189 : 228 - 0xe4
      11'hBE: dout <= 8'b00001000; //  190 :   8 - 0x8
      11'hBF: dout <= 8'b11110000; //  191 : 240 - 0xf0
      11'hC0: dout <= 8'b00111111; //  192 :  63 - 0x3f -- Sprite 0x18
      11'hC1: dout <= 8'b01000000; //  193 :  64 - 0x40
      11'hC2: dout <= 8'b01000000; //  194 :  64 - 0x40
      11'hC3: dout <= 8'b10000000; //  195 : 128 - 0x80
      11'hC4: dout <= 8'b10000000; //  196 : 128 - 0x80
      11'hC5: dout <= 8'b01111111; //  197 : 127 - 0x7f
      11'hC6: dout <= 8'b00000001; //  198 :   1 - 0x1
      11'hC7: dout <= 8'b01111111; //  199 : 127 - 0x7f
      11'hC8: dout <= 8'b11111100; //  200 : 252 - 0xfc -- Sprite 0x19
      11'hC9: dout <= 8'b00000010; //  201 :   2 - 0x2
      11'hCA: dout <= 8'b00000010; //  202 :   2 - 0x2
      11'hCB: dout <= 8'b00000001; //  203 :   1 - 0x1
      11'hCC: dout <= 8'b00000001; //  204 :   1 - 0x1
      11'hCD: dout <= 8'b11111110; //  205 : 254 - 0xfe
      11'hCE: dout <= 8'b10000000; //  206 : 128 - 0x80
      11'hCF: dout <= 8'b11111110; //  207 : 254 - 0xfe
      11'hD0: dout <= 8'b00000000; //  208 :   0 - 0x0 -- Sprite 0x1a
      11'hD1: dout <= 8'b00000000; //  209 :   0 - 0x0
      11'hD2: dout <= 8'b00111111; //  210 :  63 - 0x3f
      11'hD3: dout <= 8'b01000000; //  211 :  64 - 0x40
      11'hD4: dout <= 8'b01000000; //  212 :  64 - 0x40
      11'hD5: dout <= 8'b10000000; //  213 : 128 - 0x80
      11'hD6: dout <= 8'b10000000; //  214 : 128 - 0x80
      11'hD7: dout <= 8'b01111111; //  215 : 127 - 0x7f
      11'hD8: dout <= 8'b00000000; //  216 :   0 - 0x0 -- Sprite 0x1b
      11'hD9: dout <= 8'b00000000; //  217 :   0 - 0x0
      11'hDA: dout <= 8'b11111100; //  218 : 252 - 0xfc
      11'hDB: dout <= 8'b00000010; //  219 :   2 - 0x2
      11'hDC: dout <= 8'b00000010; //  220 :   2 - 0x2
      11'hDD: dout <= 8'b00000001; //  221 :   1 - 0x1
      11'hDE: dout <= 8'b00000001; //  222 :   1 - 0x1
      11'hDF: dout <= 8'b11111110; //  223 : 254 - 0xfe
      11'hE0: dout <= 8'b01111111; //  224 : 127 - 0x7f -- Sprite 0x1c
      11'hE1: dout <= 8'b10000000; //  225 : 128 - 0x80
      11'hE2: dout <= 8'b10000000; //  226 : 128 - 0x80
      11'hE3: dout <= 8'b10000000; //  227 : 128 - 0x80
      11'hE4: dout <= 8'b10011011; //  228 : 155 - 0x9b
      11'hE5: dout <= 8'b10100100; //  229 : 164 - 0xa4
      11'hE6: dout <= 8'b10100110; //  230 : 166 - 0xa6
      11'hE7: dout <= 8'b10000000; //  231 : 128 - 0x80
      11'hE8: dout <= 8'b10000000; //  232 : 128 - 0x80 -- Sprite 0x1d
      11'hE9: dout <= 8'b01111111; //  233 : 127 - 0x7f
      11'hEA: dout <= 8'b00000010; //  234 :   2 - 0x2
      11'hEB: dout <= 8'b00000010; //  235 :   2 - 0x2
      11'hEC: dout <= 8'b00000010; //  236 :   2 - 0x2
      11'hED: dout <= 8'b00000010; //  237 :   2 - 0x2
      11'hEE: dout <= 8'b00000010; //  238 :   2 - 0x2
      11'hEF: dout <= 8'b00001111; //  239 :  15 - 0xf
      11'hF0: dout <= 8'b11111110; //  240 : 254 - 0xfe -- Sprite 0x1e
      11'hF1: dout <= 8'b00000001; //  241 :   1 - 0x1
      11'hF2: dout <= 8'b00000001; //  242 :   1 - 0x1
      11'hF3: dout <= 8'b00000001; //  243 :   1 - 0x1
      11'hF4: dout <= 8'b01000001; //  244 :  65 - 0x41
      11'hF5: dout <= 8'b11110101; //  245 : 245 - 0xf5
      11'hF6: dout <= 8'b00011101; //  246 :  29 - 0x1d
      11'hF7: dout <= 8'b00000001; //  247 :   1 - 0x1
      11'hF8: dout <= 8'b00000001; //  248 :   1 - 0x1 -- Sprite 0x1f
      11'hF9: dout <= 8'b11111110; //  249 : 254 - 0xfe
      11'hFA: dout <= 8'b01000000; //  250 :  64 - 0x40
      11'hFB: dout <= 8'b01000000; //  251 :  64 - 0x40
      11'hFC: dout <= 8'b01000000; //  252 :  64 - 0x40
      11'hFD: dout <= 8'b01000000; //  253 :  64 - 0x40
      11'hFE: dout <= 8'b01000000; //  254 :  64 - 0x40
      11'hFF: dout <= 8'b11110000; //  255 : 240 - 0xf0
      11'h100: dout <= 8'b00000111; //  256 :   7 - 0x7 -- Sprite 0x20
      11'h101: dout <= 8'b00011111; //  257 :  31 - 0x1f
      11'h102: dout <= 8'b00111111; //  258 :  63 - 0x3f
      11'h103: dout <= 8'b01111111; //  259 : 127 - 0x7f
      11'h104: dout <= 8'b01111111; //  260 : 127 - 0x7f
      11'h105: dout <= 8'b11111111; //  261 : 255 - 0xff
      11'h106: dout <= 8'b11111111; //  262 : 255 - 0xff
      11'h107: dout <= 8'b11111111; //  263 : 255 - 0xff
      11'h108: dout <= 8'b11100000; //  264 : 224 - 0xe0 -- Sprite 0x21
      11'h109: dout <= 8'b11111000; //  265 : 248 - 0xf8
      11'h10A: dout <= 8'b11111100; //  266 : 252 - 0xfc
      11'h10B: dout <= 8'b11111110; //  267 : 254 - 0xfe
      11'h10C: dout <= 8'b11111110; //  268 : 254 - 0xfe
      11'h10D: dout <= 8'b11111111; //  269 : 255 - 0xff
      11'h10E: dout <= 8'b11111111; //  270 : 255 - 0xff
      11'h10F: dout <= 8'b11111111; //  271 : 255 - 0xff
      11'h110: dout <= 8'b00000111; //  272 :   7 - 0x7 -- Sprite 0x22
      11'h111: dout <= 8'b00011111; //  273 :  31 - 0x1f
      11'h112: dout <= 8'b00111111; //  274 :  63 - 0x3f
      11'h113: dout <= 8'b01111111; //  275 : 127 - 0x7f
      11'h114: dout <= 8'b01111111; //  276 : 127 - 0x7f
      11'h115: dout <= 8'b11111111; //  277 : 255 - 0xff
      11'h116: dout <= 8'b11111111; //  278 : 255 - 0xff
      11'h117: dout <= 8'b11111111; //  279 : 255 - 0xff
      11'h118: dout <= 8'b11100000; //  280 : 224 - 0xe0 -- Sprite 0x23
      11'h119: dout <= 8'b11111000; //  281 : 248 - 0xf8
      11'h11A: dout <= 8'b11111100; //  282 : 252 - 0xfc
      11'h11B: dout <= 8'b11111110; //  283 : 254 - 0xfe
      11'h11C: dout <= 8'b11111110; //  284 : 254 - 0xfe
      11'h11D: dout <= 8'b11111111; //  285 : 255 - 0xff
      11'h11E: dout <= 8'b11111111; //  286 : 255 - 0xff
      11'h11F: dout <= 8'b11111111; //  287 : 255 - 0xff
      11'h120: dout <= 8'b00000000; //  288 :   0 - 0x0 -- Sprite 0x24
      11'h121: dout <= 8'b00000000; //  289 :   0 - 0x0
      11'h122: dout <= 8'b00000000; //  290 :   0 - 0x0
      11'h123: dout <= 8'b00000000; //  291 :   0 - 0x0
      11'h124: dout <= 8'b00000000; //  292 :   0 - 0x0
      11'h125: dout <= 8'b00000000; //  293 :   0 - 0x0
      11'h126: dout <= 8'b00000000; //  294 :   0 - 0x0
      11'h127: dout <= 8'b00000000; //  295 :   0 - 0x0
      11'h128: dout <= 8'b00101111; //  296 :  47 - 0x2f -- Sprite 0x25
      11'h129: dout <= 8'b01001111; //  297 :  79 - 0x4f
      11'h12A: dout <= 8'b01001111; //  298 :  79 - 0x4f
      11'h12B: dout <= 8'b01001111; //  299 :  79 - 0x4f
      11'h12C: dout <= 8'b01001111; //  300 :  79 - 0x4f
      11'h12D: dout <= 8'b00100111; //  301 :  39 - 0x27
      11'h12E: dout <= 8'b00010000; //  302 :  16 - 0x10
      11'h12F: dout <= 8'b00001111; //  303 :  15 - 0xf
      11'h130: dout <= 8'b00000000; //  304 :   0 - 0x0 -- Sprite 0x26
      11'h131: dout <= 8'b11100000; //  305 : 224 - 0xe0
      11'h132: dout <= 8'b10100000; //  306 : 160 - 0xa0
      11'h133: dout <= 8'b00100000; //  307 :  32 - 0x20
      11'h134: dout <= 8'b11000000; //  308 : 192 - 0xc0
      11'h135: dout <= 8'b01000000; //  309 :  64 - 0x40
      11'h136: dout <= 8'b00110000; //  310 :  48 - 0x30
      11'h137: dout <= 8'b11101000; //  311 : 232 - 0xe8
      11'h138: dout <= 8'b11110100; //  312 : 244 - 0xf4 -- Sprite 0x27
      11'h139: dout <= 8'b11110010; //  313 : 242 - 0xf2
      11'h13A: dout <= 8'b11110010; //  314 : 242 - 0xf2
      11'h13B: dout <= 8'b11110010; //  315 : 242 - 0xf2
      11'h13C: dout <= 8'b11110010; //  316 : 242 - 0xf2
      11'h13D: dout <= 8'b11100100; //  317 : 228 - 0xe4
      11'h13E: dout <= 8'b00001000; //  318 :   8 - 0x8
      11'h13F: dout <= 8'b11110000; //  319 : 240 - 0xf0
      11'h140: dout <= 8'b11111111; //  320 : 255 - 0xff -- Sprite 0x28
      11'h141: dout <= 8'b11010101; //  321 : 213 - 0xd5
      11'h142: dout <= 8'b10100011; //  322 : 163 - 0xa3
      11'h143: dout <= 8'b11010111; //  323 : 215 - 0xd7
      11'h144: dout <= 8'b10001111; //  324 : 143 - 0x8f
      11'h145: dout <= 8'b11001111; //  325 : 207 - 0xcf
      11'h146: dout <= 8'b10001011; //  326 : 139 - 0x8b
      11'h147: dout <= 8'b11001011; //  327 : 203 - 0xcb
      11'h148: dout <= 8'b10001111; //  328 : 143 - 0x8f -- Sprite 0x29
      11'h149: dout <= 8'b11001111; //  329 : 207 - 0xcf
      11'h14A: dout <= 8'b10001111; //  330 : 143 - 0x8f
      11'h14B: dout <= 8'b11001111; //  331 : 207 - 0xcf
      11'h14C: dout <= 8'b10010000; //  332 : 144 - 0x90
      11'h14D: dout <= 8'b11100000; //  333 : 224 - 0xe0
      11'h14E: dout <= 8'b11101010; //  334 : 234 - 0xea
      11'h14F: dout <= 8'b11111111; //  335 : 255 - 0xff
      11'h150: dout <= 8'b11111111; //  336 : 255 - 0xff -- Sprite 0x2a
      11'h151: dout <= 8'b11011011; //  337 : 219 - 0xdb
      11'h152: dout <= 8'b11000111; //  338 : 199 - 0xc7
      11'h153: dout <= 8'b11101001; //  339 : 233 - 0xe9
      11'h154: dout <= 8'b11110011; //  340 : 243 - 0xf3
      11'h155: dout <= 8'b11110001; //  341 : 241 - 0xf1
      11'h156: dout <= 8'b11010011; //  342 : 211 - 0xd3
      11'h157: dout <= 8'b11010001; //  343 : 209 - 0xd1
      11'h158: dout <= 8'b11110011; //  344 : 243 - 0xf3 -- Sprite 0x2b
      11'h159: dout <= 8'b11110001; //  345 : 241 - 0xf1
      11'h15A: dout <= 8'b11110011; //  346 : 243 - 0xf3
      11'h15B: dout <= 8'b11110001; //  347 : 241 - 0xf1
      11'h15C: dout <= 8'b00001011; //  348 :  11 - 0xb
      11'h15D: dout <= 8'b00000101; //  349 :   5 - 0x5
      11'h15E: dout <= 8'b10101011; //  350 : 171 - 0xab
      11'h15F: dout <= 8'b11111111; //  351 : 255 - 0xff
      11'h160: dout <= 8'b00000000; //  352 :   0 - 0x0 -- Sprite 0x2c
      11'h161: dout <= 8'b00000000; //  353 :   0 - 0x0
      11'h162: dout <= 8'b00000000; //  354 :   0 - 0x0
      11'h163: dout <= 8'b00000000; //  355 :   0 - 0x0
      11'h164: dout <= 8'b00000000; //  356 :   0 - 0x0
      11'h165: dout <= 8'b00000000; //  357 :   0 - 0x0
      11'h166: dout <= 8'b00000000; //  358 :   0 - 0x0
      11'h167: dout <= 8'b00000000; //  359 :   0 - 0x0
      11'h168: dout <= 8'b00101111; //  360 :  47 - 0x2f -- Sprite 0x2d
      11'h169: dout <= 8'b01001111; //  361 :  79 - 0x4f
      11'h16A: dout <= 8'b01001111; //  362 :  79 - 0x4f
      11'h16B: dout <= 8'b01001111; //  363 :  79 - 0x4f
      11'h16C: dout <= 8'b01001111; //  364 :  79 - 0x4f
      11'h16D: dout <= 8'b00100111; //  365 :  39 - 0x27
      11'h16E: dout <= 8'b00010000; //  366 :  16 - 0x10
      11'h16F: dout <= 8'b00001111; //  367 :  15 - 0xf
      11'h170: dout <= 8'b00000000; //  368 :   0 - 0x0 -- Sprite 0x2e
      11'h171: dout <= 8'b00000000; //  369 :   0 - 0x0
      11'h172: dout <= 8'b00000000; //  370 :   0 - 0x0
      11'h173: dout <= 8'b00000000; //  371 :   0 - 0x0
      11'h174: dout <= 8'b00000000; //  372 :   0 - 0x0
      11'h175: dout <= 8'b00000000; //  373 :   0 - 0x0
      11'h176: dout <= 8'b00000000; //  374 :   0 - 0x0
      11'h177: dout <= 8'b00000000; //  375 :   0 - 0x0
      11'h178: dout <= 8'b11110100; //  376 : 244 - 0xf4 -- Sprite 0x2f
      11'h179: dout <= 8'b11110010; //  377 : 242 - 0xf2
      11'h17A: dout <= 8'b11110010; //  378 : 242 - 0xf2
      11'h17B: dout <= 8'b11110010; //  379 : 242 - 0xf2
      11'h17C: dout <= 8'b11110010; //  380 : 242 - 0xf2
      11'h17D: dout <= 8'b11100100; //  381 : 228 - 0xe4
      11'h17E: dout <= 8'b00001000; //  382 :   8 - 0x8
      11'h17F: dout <= 8'b11110000; //  383 : 240 - 0xf0
      11'h180: dout <= 8'b00011000; //  384 :  24 - 0x18 -- Sprite 0x30
      11'h181: dout <= 8'b00100100; //  385 :  36 - 0x24
      11'h182: dout <= 8'b01000010; //  386 :  66 - 0x42
      11'h183: dout <= 8'b10100101; //  387 : 165 - 0xa5
      11'h184: dout <= 8'b11100111; //  388 : 231 - 0xe7
      11'h185: dout <= 8'b00100100; //  389 :  36 - 0x24
      11'h186: dout <= 8'b00100100; //  390 :  36 - 0x24
      11'h187: dout <= 8'b00111100; //  391 :  60 - 0x3c
      11'h188: dout <= 8'b00111100; //  392 :  60 - 0x3c -- Sprite 0x31
      11'h189: dout <= 8'b00100100; //  393 :  36 - 0x24
      11'h18A: dout <= 8'b00100100; //  394 :  36 - 0x24
      11'h18B: dout <= 8'b01100110; //  395 : 102 - 0x66
      11'h18C: dout <= 8'b10100101; //  396 : 165 - 0xa5
      11'h18D: dout <= 8'b01000010; //  397 :  66 - 0x42
      11'h18E: dout <= 8'b00100100; //  398 :  36 - 0x24
      11'h18F: dout <= 8'b00011000; //  399 :  24 - 0x18
      11'h190: dout <= 8'b00000010; //  400 :   2 - 0x2 -- Sprite 0x32
      11'h191: dout <= 8'b00000010; //  401 :   2 - 0x2
      11'h192: dout <= 8'b00000011; //  402 :   3 - 0x3
      11'h193: dout <= 8'b00000010; //  403 :   2 - 0x2
      11'h194: dout <= 8'b00000010; //  404 :   2 - 0x2
      11'h195: dout <= 8'b00000010; //  405 :   2 - 0x2
      11'h196: dout <= 8'b00000011; //  406 :   3 - 0x3
      11'h197: dout <= 8'b00000010; //  407 :   2 - 0x2
      11'h198: dout <= 8'b01000000; //  408 :  64 - 0x40 -- Sprite 0x33
      11'h199: dout <= 8'b11000000; //  409 : 192 - 0xc0
      11'h19A: dout <= 8'b01000000; //  410 :  64 - 0x40
      11'h19B: dout <= 8'b01000000; //  411 :  64 - 0x40
      11'h19C: dout <= 8'b01000000; //  412 :  64 - 0x40
      11'h19D: dout <= 8'b11000000; //  413 : 192 - 0xc0
      11'h19E: dout <= 8'b01000000; //  414 :  64 - 0x40
      11'h19F: dout <= 8'b01000000; //  415 :  64 - 0x40
      11'h1A0: dout <= 8'b00000000; //  416 :   0 - 0x0 -- Sprite 0x34
      11'h1A1: dout <= 8'b00011000; //  417 :  24 - 0x18
      11'h1A2: dout <= 8'b00111100; //  418 :  60 - 0x3c
      11'h1A3: dout <= 8'b01100010; //  419 :  98 - 0x62
      11'h1A4: dout <= 8'b01100001; //  420 :  97 - 0x61
      11'h1A5: dout <= 8'b11000000; //  421 : 192 - 0xc0
      11'h1A6: dout <= 8'b11000000; //  422 : 192 - 0xc0
      11'h1A7: dout <= 8'b11000000; //  423 : 192 - 0xc0
      11'h1A8: dout <= 8'b01100000; //  424 :  96 - 0x60 -- Sprite 0x35
      11'h1A9: dout <= 8'b01100000; //  425 :  96 - 0x60
      11'h1AA: dout <= 8'b00110000; //  426 :  48 - 0x30
      11'h1AB: dout <= 8'b00011000; //  427 :  24 - 0x18
      11'h1AC: dout <= 8'b00001100; //  428 :  12 - 0xc
      11'h1AD: dout <= 8'b00000110; //  429 :   6 - 0x6
      11'h1AE: dout <= 8'b00000010; //  430 :   2 - 0x2
      11'h1AF: dout <= 8'b00000001; //  431 :   1 - 0x1
      11'h1B0: dout <= 8'b00000000; //  432 :   0 - 0x0 -- Sprite 0x36
      11'h1B1: dout <= 8'b00011000; //  433 :  24 - 0x18
      11'h1B2: dout <= 8'b00100100; //  434 :  36 - 0x24
      11'h1B3: dout <= 8'b01000010; //  435 :  66 - 0x42
      11'h1B4: dout <= 8'b10000010; //  436 : 130 - 0x82
      11'h1B5: dout <= 8'b00000001; //  437 :   1 - 0x1
      11'h1B6: dout <= 8'b00000001; //  438 :   1 - 0x1
      11'h1B7: dout <= 8'b00000001; //  439 :   1 - 0x1
      11'h1B8: dout <= 8'b00000010; //  440 :   2 - 0x2 -- Sprite 0x37
      11'h1B9: dout <= 8'b00000010; //  441 :   2 - 0x2
      11'h1BA: dout <= 8'b00000100; //  442 :   4 - 0x4
      11'h1BB: dout <= 8'b00001000; //  443 :   8 - 0x8
      11'h1BC: dout <= 8'b00010000; //  444 :  16 - 0x10
      11'h1BD: dout <= 8'b00100000; //  445 :  32 - 0x20
      11'h1BE: dout <= 8'b01000000; //  446 :  64 - 0x40
      11'h1BF: dout <= 8'b10000000; //  447 : 128 - 0x80
      11'h1C0: dout <= 8'b00000000; //  448 :   0 - 0x0 -- Sprite 0x38
      11'h1C1: dout <= 8'b00000110; //  449 :   6 - 0x6
      11'h1C2: dout <= 8'b00001101; //  450 :  13 - 0xd
      11'h1C3: dout <= 8'b00001100; //  451 :  12 - 0xc
      11'h1C4: dout <= 8'b00001100; //  452 :  12 - 0xc
      11'h1C5: dout <= 8'b00000110; //  453 :   6 - 0x6
      11'h1C6: dout <= 8'b00000010; //  454 :   2 - 0x2
      11'h1C7: dout <= 8'b00000001; //  455 :   1 - 0x1
      11'h1C8: dout <= 8'b11111111; //  456 : 255 - 0xff -- Sprite 0x39
      11'h1C9: dout <= 8'b00000000; //  457 :   0 - 0x0
      11'h1CA: dout <= 8'b00000000; //  458 :   0 - 0x0
      11'h1CB: dout <= 8'b00000000; //  459 :   0 - 0x0
      11'h1CC: dout <= 8'b00000000; //  460 :   0 - 0x0
      11'h1CD: dout <= 8'b00000000; //  461 :   0 - 0x0
      11'h1CE: dout <= 8'b00000000; //  462 :   0 - 0x0
      11'h1CF: dout <= 8'b00000000; //  463 :   0 - 0x0
      11'h1D0: dout <= 8'b00000000; //  464 :   0 - 0x0 -- Sprite 0x3a
      11'h1D1: dout <= 8'b01100000; //  465 :  96 - 0x60
      11'h1D2: dout <= 8'b10010000; //  466 : 144 - 0x90
      11'h1D3: dout <= 8'b00010000; //  467 :  16 - 0x10
      11'h1D4: dout <= 8'b00010000; //  468 :  16 - 0x10
      11'h1D5: dout <= 8'b00100000; //  469 :  32 - 0x20
      11'h1D6: dout <= 8'b01000000; //  470 :  64 - 0x40
      11'h1D7: dout <= 8'b10000000; //  471 : 128 - 0x80
      11'h1D8: dout <= 8'b00000000; //  472 :   0 - 0x0 -- Sprite 0x3b
      11'h1D9: dout <= 8'b01010100; //  473 :  84 - 0x54
      11'h1DA: dout <= 8'b00000010; //  474 :   2 - 0x2
      11'h1DB: dout <= 8'b01000000; //  475 :  64 - 0x40
      11'h1DC: dout <= 8'b00000010; //  476 :   2 - 0x2
      11'h1DD: dout <= 8'b01000000; //  477 :  64 - 0x40
      11'h1DE: dout <= 8'b00101010; //  478 :  42 - 0x2a
      11'h1DF: dout <= 8'b00000000; //  479 :   0 - 0x0
      11'h1E0: dout <= 8'b11111111; //  480 : 255 - 0xff -- Sprite 0x3c
      11'h1E1: dout <= 8'b11111111; //  481 : 255 - 0xff
      11'h1E2: dout <= 8'b11111111; //  482 : 255 - 0xff
      11'h1E3: dout <= 8'b11111111; //  483 : 255 - 0xff
      11'h1E4: dout <= 8'b11111111; //  484 : 255 - 0xff
      11'h1E5: dout <= 8'b11111111; //  485 : 255 - 0xff
      11'h1E6: dout <= 8'b11111111; //  486 : 255 - 0xff
      11'h1E7: dout <= 8'b11111111; //  487 : 255 - 0xff
      11'h1E8: dout <= 8'b00000000; //  488 :   0 - 0x0 -- Sprite 0x3d
      11'h1E9: dout <= 8'b00000000; //  489 :   0 - 0x0
      11'h1EA: dout <= 8'b00000000; //  490 :   0 - 0x0
      11'h1EB: dout <= 8'b00000000; //  491 :   0 - 0x0
      11'h1EC: dout <= 8'b00000000; //  492 :   0 - 0x0
      11'h1ED: dout <= 8'b00000000; //  493 :   0 - 0x0
      11'h1EE: dout <= 8'b00000000; //  494 :   0 - 0x0
      11'h1EF: dout <= 8'b00000000; //  495 :   0 - 0x0
      11'h1F0: dout <= 8'b11111111; //  496 : 255 - 0xff -- Sprite 0x3e
      11'h1F1: dout <= 8'b11111111; //  497 : 255 - 0xff
      11'h1F2: dout <= 8'b11111111; //  498 : 255 - 0xff
      11'h1F3: dout <= 8'b11111111; //  499 : 255 - 0xff
      11'h1F4: dout <= 8'b11111111; //  500 : 255 - 0xff
      11'h1F5: dout <= 8'b11111111; //  501 : 255 - 0xff
      11'h1F6: dout <= 8'b11111111; //  502 : 255 - 0xff
      11'h1F7: dout <= 8'b11111111; //  503 : 255 - 0xff
      11'h1F8: dout <= 8'b00000000; //  504 :   0 - 0x0 -- Sprite 0x3f
      11'h1F9: dout <= 8'b00000000; //  505 :   0 - 0x0
      11'h1FA: dout <= 8'b00000000; //  506 :   0 - 0x0
      11'h1FB: dout <= 8'b00000000; //  507 :   0 - 0x0
      11'h1FC: dout <= 8'b00000000; //  508 :   0 - 0x0
      11'h1FD: dout <= 8'b00000000; //  509 :   0 - 0x0
      11'h1FE: dout <= 8'b00000000; //  510 :   0 - 0x0
      11'h1FF: dout <= 8'b00000000; //  511 :   0 - 0x0
      11'h200: dout <= 8'b00111100; //  512 :  60 - 0x3c -- Sprite 0x40
      11'h201: dout <= 8'b01000010; //  513 :  66 - 0x42
      11'h202: dout <= 8'b10011001; //  514 : 153 - 0x99
      11'h203: dout <= 8'b10100101; //  515 : 165 - 0xa5
      11'h204: dout <= 8'b10100101; //  516 : 165 - 0xa5
      11'h205: dout <= 8'b10011010; //  517 : 154 - 0x9a
      11'h206: dout <= 8'b01000000; //  518 :  64 - 0x40
      11'h207: dout <= 8'b00111100; //  519 :  60 - 0x3c
      11'h208: dout <= 8'b00001100; //  520 :  12 - 0xc -- Sprite 0x41
      11'h209: dout <= 8'b00010010; //  521 :  18 - 0x12
      11'h20A: dout <= 8'b00100010; //  522 :  34 - 0x22
      11'h20B: dout <= 8'b00100010; //  523 :  34 - 0x22
      11'h20C: dout <= 8'b01111110; //  524 : 126 - 0x7e
      11'h20D: dout <= 8'b00100010; //  525 :  34 - 0x22
      11'h20E: dout <= 8'b00100100; //  526 :  36 - 0x24
      11'h20F: dout <= 8'b00000000; //  527 :   0 - 0x0
      11'h210: dout <= 8'b00111100; //  528 :  60 - 0x3c -- Sprite 0x42
      11'h211: dout <= 8'b01000010; //  529 :  66 - 0x42
      11'h212: dout <= 8'b01010010; //  530 :  82 - 0x52
      11'h213: dout <= 8'b00011100; //  531 :  28 - 0x1c
      11'h214: dout <= 8'b00010010; //  532 :  18 - 0x12
      11'h215: dout <= 8'b00110010; //  533 :  50 - 0x32
      11'h216: dout <= 8'b00011100; //  534 :  28 - 0x1c
      11'h217: dout <= 8'b00000000; //  535 :   0 - 0x0
      11'h218: dout <= 8'b00011000; //  536 :  24 - 0x18 -- Sprite 0x43
      11'h219: dout <= 8'b00100100; //  537 :  36 - 0x24
      11'h21A: dout <= 8'b01010100; //  538 :  84 - 0x54
      11'h21B: dout <= 8'b01001000; //  539 :  72 - 0x48
      11'h21C: dout <= 8'b01000010; //  540 :  66 - 0x42
      11'h21D: dout <= 8'b00100100; //  541 :  36 - 0x24
      11'h21E: dout <= 8'b00011000; //  542 :  24 - 0x18
      11'h21F: dout <= 8'b00000000; //  543 :   0 - 0x0
      11'h220: dout <= 8'b01011000; //  544 :  88 - 0x58 -- Sprite 0x44
      11'h221: dout <= 8'b11100100; //  545 : 228 - 0xe4
      11'h222: dout <= 8'b01000010; //  546 :  66 - 0x42
      11'h223: dout <= 8'b01000010; //  547 :  66 - 0x42
      11'h224: dout <= 8'b00100010; //  548 :  34 - 0x22
      11'h225: dout <= 8'b01100100; //  549 : 100 - 0x64
      11'h226: dout <= 8'b00111000; //  550 :  56 - 0x38
      11'h227: dout <= 8'b00000000; //  551 :   0 - 0x0
      11'h228: dout <= 8'b00011100; //  552 :  28 - 0x1c -- Sprite 0x45
      11'h229: dout <= 8'b00100000; //  553 :  32 - 0x20
      11'h22A: dout <= 8'b00100000; //  554 :  32 - 0x20
      11'h22B: dout <= 8'b00101100; //  555 :  44 - 0x2c
      11'h22C: dout <= 8'b01110000; //  556 : 112 - 0x70
      11'h22D: dout <= 8'b00100010; //  557 :  34 - 0x22
      11'h22E: dout <= 8'b00011100; //  558 :  28 - 0x1c
      11'h22F: dout <= 8'b00000000; //  559 :   0 - 0x0
      11'h230: dout <= 8'b00011100; //  560 :  28 - 0x1c -- Sprite 0x46
      11'h231: dout <= 8'b00100000; //  561 :  32 - 0x20
      11'h232: dout <= 8'b00100000; //  562 :  32 - 0x20
      11'h233: dout <= 8'b00101100; //  563 :  44 - 0x2c
      11'h234: dout <= 8'b01110000; //  564 : 112 - 0x70
      11'h235: dout <= 8'b00010000; //  565 :  16 - 0x10
      11'h236: dout <= 8'b00010000; //  566 :  16 - 0x10
      11'h237: dout <= 8'b00000000; //  567 :   0 - 0x0
      11'h238: dout <= 8'b00011000; //  568 :  24 - 0x18 -- Sprite 0x47
      11'h239: dout <= 8'b00100100; //  569 :  36 - 0x24
      11'h23A: dout <= 8'b01000000; //  570 :  64 - 0x40
      11'h23B: dout <= 8'b01001110; //  571 :  78 - 0x4e
      11'h23C: dout <= 8'b01000010; //  572 :  66 - 0x42
      11'h23D: dout <= 8'b00100100; //  573 :  36 - 0x24
      11'h23E: dout <= 8'b00011000; //  574 :  24 - 0x18
      11'h23F: dout <= 8'b00000000; //  575 :   0 - 0x0
      11'h240: dout <= 8'b00100000; //  576 :  32 - 0x20 -- Sprite 0x48
      11'h241: dout <= 8'b01000100; //  577 :  68 - 0x44
      11'h242: dout <= 8'b01000100; //  578 :  68 - 0x44
      11'h243: dout <= 8'b01000100; //  579 :  68 - 0x44
      11'h244: dout <= 8'b11111100; //  580 : 252 - 0xfc
      11'h245: dout <= 8'b01000100; //  581 :  68 - 0x44
      11'h246: dout <= 8'b01001000; //  582 :  72 - 0x48
      11'h247: dout <= 8'b00000000; //  583 :   0 - 0x0
      11'h248: dout <= 8'b00010000; //  584 :  16 - 0x10 -- Sprite 0x49
      11'h249: dout <= 8'b00010000; //  585 :  16 - 0x10
      11'h24A: dout <= 8'b00010000; //  586 :  16 - 0x10
      11'h24B: dout <= 8'b00010000; //  587 :  16 - 0x10
      11'h24C: dout <= 8'b00010000; //  588 :  16 - 0x10
      11'h24D: dout <= 8'b00001000; //  589 :   8 - 0x8
      11'h24E: dout <= 8'b00001000; //  590 :   8 - 0x8
      11'h24F: dout <= 8'b00000000; //  591 :   0 - 0x0
      11'h250: dout <= 8'b00001000; //  592 :   8 - 0x8 -- Sprite 0x4a
      11'h251: dout <= 8'b00001000; //  593 :   8 - 0x8
      11'h252: dout <= 8'b00000100; //  594 :   4 - 0x4
      11'h253: dout <= 8'b00000100; //  595 :   4 - 0x4
      11'h254: dout <= 8'b01000100; //  596 :  68 - 0x44
      11'h255: dout <= 8'b01001000; //  597 :  72 - 0x48
      11'h256: dout <= 8'b00110000; //  598 :  48 - 0x30
      11'h257: dout <= 8'b00000000; //  599 :   0 - 0x0
      11'h258: dout <= 8'b01000100; //  600 :  68 - 0x44 -- Sprite 0x4b
      11'h259: dout <= 8'b01000100; //  601 :  68 - 0x44
      11'h25A: dout <= 8'b01001000; //  602 :  72 - 0x48
      11'h25B: dout <= 8'b01110000; //  603 : 112 - 0x70
      11'h25C: dout <= 8'b01001000; //  604 :  72 - 0x48
      11'h25D: dout <= 8'b00100100; //  605 :  36 - 0x24
      11'h25E: dout <= 8'b00100010; //  606 :  34 - 0x22
      11'h25F: dout <= 8'b00000000; //  607 :   0 - 0x0
      11'h260: dout <= 8'b00010000; //  608 :  16 - 0x10 -- Sprite 0x4c
      11'h261: dout <= 8'b00100000; //  609 :  32 - 0x20
      11'h262: dout <= 8'b00100000; //  610 :  32 - 0x20
      11'h263: dout <= 8'b00100000; //  611 :  32 - 0x20
      11'h264: dout <= 8'b01000000; //  612 :  64 - 0x40
      11'h265: dout <= 8'b01000000; //  613 :  64 - 0x40
      11'h266: dout <= 8'b01000110; //  614 :  70 - 0x46
      11'h267: dout <= 8'b00111000; //  615 :  56 - 0x38
      11'h268: dout <= 8'b00100100; //  616 :  36 - 0x24 -- Sprite 0x4d
      11'h269: dout <= 8'b01011010; //  617 :  90 - 0x5a
      11'h26A: dout <= 8'b01011010; //  618 :  90 - 0x5a
      11'h26B: dout <= 8'b01011010; //  619 :  90 - 0x5a
      11'h26C: dout <= 8'b01000010; //  620 :  66 - 0x42
      11'h26D: dout <= 8'b01000010; //  621 :  66 - 0x42
      11'h26E: dout <= 8'b00100010; //  622 :  34 - 0x22
      11'h26F: dout <= 8'b00000000; //  623 :   0 - 0x0
      11'h270: dout <= 8'b00100100; //  624 :  36 - 0x24 -- Sprite 0x4e
      11'h271: dout <= 8'b01010010; //  625 :  82 - 0x52
      11'h272: dout <= 8'b01010010; //  626 :  82 - 0x52
      11'h273: dout <= 8'b01010010; //  627 :  82 - 0x52
      11'h274: dout <= 8'b01010010; //  628 :  82 - 0x52
      11'h275: dout <= 8'b01010010; //  629 :  82 - 0x52
      11'h276: dout <= 8'b01001100; //  630 :  76 - 0x4c
      11'h277: dout <= 8'b00000000; //  631 :   0 - 0x0
      11'h278: dout <= 8'b00111000; //  632 :  56 - 0x38 -- Sprite 0x4f
      11'h279: dout <= 8'b01000100; //  633 :  68 - 0x44
      11'h27A: dout <= 8'b10000010; //  634 : 130 - 0x82
      11'h27B: dout <= 8'b10000010; //  635 : 130 - 0x82
      11'h27C: dout <= 8'b10000010; //  636 : 130 - 0x82
      11'h27D: dout <= 8'b01000100; //  637 :  68 - 0x44
      11'h27E: dout <= 8'b00111000; //  638 :  56 - 0x38
      11'h27F: dout <= 8'b00000000; //  639 :   0 - 0x0
      11'h280: dout <= 8'b01111111; //  640 : 127 - 0x7f -- Sprite 0x50
      11'h281: dout <= 8'b11000000; //  641 : 192 - 0xc0
      11'h282: dout <= 8'b10000000; //  642 : 128 - 0x80
      11'h283: dout <= 8'b10000000; //  643 : 128 - 0x80
      11'h284: dout <= 8'b10000000; //  644 : 128 - 0x80
      11'h285: dout <= 8'b11000011; //  645 : 195 - 0xc3
      11'h286: dout <= 8'b11111111; //  646 : 255 - 0xff
      11'h287: dout <= 8'b11111111; //  647 : 255 - 0xff
      11'h288: dout <= 8'b11111110; //  648 : 254 - 0xfe -- Sprite 0x51
      11'h289: dout <= 8'b00000011; //  649 :   3 - 0x3
      11'h28A: dout <= 8'b00000001; //  650 :   1 - 0x1
      11'h28B: dout <= 8'b00000001; //  651 :   1 - 0x1
      11'h28C: dout <= 8'b00000001; //  652 :   1 - 0x1
      11'h28D: dout <= 8'b11000011; //  653 : 195 - 0xc3
      11'h28E: dout <= 8'b11111111; //  654 : 255 - 0xff
      11'h28F: dout <= 8'b11111111; //  655 : 255 - 0xff
      11'h290: dout <= 8'b00000000; //  656 :   0 - 0x0 -- Sprite 0x52
      11'h291: dout <= 8'b00000111; //  657 :   7 - 0x7
      11'h292: dout <= 8'b00001100; //  658 :  12 - 0xc
      11'h293: dout <= 8'b00011000; //  659 :  24 - 0x18
      11'h294: dout <= 8'b00110000; //  660 :  48 - 0x30
      11'h295: dout <= 8'b01100000; //  661 :  96 - 0x60
      11'h296: dout <= 8'b01000000; //  662 :  64 - 0x40
      11'h297: dout <= 8'b01001111; //  663 :  79 - 0x4f
      11'h298: dout <= 8'b00000000; //  664 :   0 - 0x0 -- Sprite 0x53
      11'h299: dout <= 8'b11110000; //  665 : 240 - 0xf0
      11'h29A: dout <= 8'b01010000; //  666 :  80 - 0x50
      11'h29B: dout <= 8'b01001000; //  667 :  72 - 0x48
      11'h29C: dout <= 8'b01001100; //  668 :  76 - 0x4c
      11'h29D: dout <= 8'b01000100; //  669 :  68 - 0x44
      11'h29E: dout <= 8'b10000010; //  670 : 130 - 0x82
      11'h29F: dout <= 8'b10000011; //  671 : 131 - 0x83
      11'h2A0: dout <= 8'b01111111; //  672 : 127 - 0x7f -- Sprite 0x54
      11'h2A1: dout <= 8'b11011110; //  673 : 222 - 0xde
      11'h2A2: dout <= 8'b10001110; //  674 : 142 - 0x8e
      11'h2A3: dout <= 8'b11000101; //  675 : 197 - 0xc5
      11'h2A4: dout <= 8'b10010010; //  676 : 146 - 0x92
      11'h2A5: dout <= 8'b11000111; //  677 : 199 - 0xc7
      11'h2A6: dout <= 8'b11100010; //  678 : 226 - 0xe2
      11'h2A7: dout <= 8'b11010000; //  679 : 208 - 0xd0
      11'h2A8: dout <= 8'b11111111; //  680 : 255 - 0xff -- Sprite 0x55
      11'h2A9: dout <= 8'b11011110; //  681 : 222 - 0xde
      11'h2AA: dout <= 8'b10001110; //  682 : 142 - 0x8e
      11'h2AB: dout <= 8'b11000101; //  683 : 197 - 0xc5
      11'h2AC: dout <= 8'b10010010; //  684 : 146 - 0x92
      11'h2AD: dout <= 8'b01000111; //  685 :  71 - 0x47
      11'h2AE: dout <= 8'b11100010; //  686 : 226 - 0xe2
      11'h2AF: dout <= 8'b01010000; //  687 :  80 - 0x50
      11'h2B0: dout <= 8'b11111110; //  688 : 254 - 0xfe -- Sprite 0x56
      11'h2B1: dout <= 8'b11011111; //  689 : 223 - 0xdf
      11'h2B2: dout <= 8'b10001111; //  690 : 143 - 0x8f
      11'h2B3: dout <= 8'b11000101; //  691 : 197 - 0xc5
      11'h2B4: dout <= 8'b10010011; //  692 : 147 - 0x93
      11'h2B5: dout <= 8'b01000111; //  693 :  71 - 0x47
      11'h2B6: dout <= 8'b11100011; //  694 : 227 - 0xe3
      11'h2B7: dout <= 8'b01010001; //  695 :  81 - 0x51
      11'h2B8: dout <= 8'b01111111; //  696 : 127 - 0x7f -- Sprite 0x57
      11'h2B9: dout <= 8'b10000000; //  697 : 128 - 0x80
      11'h2BA: dout <= 8'b10110011; //  698 : 179 - 0xb3
      11'h2BB: dout <= 8'b01001100; //  699 :  76 - 0x4c
      11'h2BC: dout <= 8'b00111111; //  700 :  63 - 0x3f
      11'h2BD: dout <= 8'b00000011; //  701 :   3 - 0x3
      11'h2BE: dout <= 8'b00000000; //  702 :   0 - 0x0
      11'h2BF: dout <= 8'b00000000; //  703 :   0 - 0x0
      11'h2C0: dout <= 8'b11111111; //  704 : 255 - 0xff -- Sprite 0x58
      11'h2C1: dout <= 8'b00000000; //  705 :   0 - 0x0
      11'h2C2: dout <= 8'b00110011; //  706 :  51 - 0x33
      11'h2C3: dout <= 8'b11001100; //  707 : 204 - 0xcc
      11'h2C4: dout <= 8'b00110011; //  708 :  51 - 0x33
      11'h2C5: dout <= 8'b11111111; //  709 : 255 - 0xff
      11'h2C6: dout <= 8'b00000000; //  710 :   0 - 0x0
      11'h2C7: dout <= 8'b00000000; //  711 :   0 - 0x0
      11'h2C8: dout <= 8'b11111110; //  712 : 254 - 0xfe -- Sprite 0x59
      11'h2C9: dout <= 8'b00000001; //  713 :   1 - 0x1
      11'h2CA: dout <= 8'b00110011; //  714 :  51 - 0x33
      11'h2CB: dout <= 8'b11001110; //  715 : 206 - 0xce
      11'h2CC: dout <= 8'b00111100; //  716 :  60 - 0x3c
      11'h2CD: dout <= 8'b11000000; //  717 : 192 - 0xc0
      11'h2CE: dout <= 8'b00000000; //  718 :   0 - 0x0
      11'h2CF: dout <= 8'b00000000; //  719 :   0 - 0x0
      11'h2D0: dout <= 8'b00000000; //  720 :   0 - 0x0 -- Sprite 0x5a
      11'h2D1: dout <= 8'b00000000; //  721 :   0 - 0x0
      11'h2D2: dout <= 8'b00000000; //  722 :   0 - 0x0
      11'h2D3: dout <= 8'b00000000; //  723 :   0 - 0x0
      11'h2D4: dout <= 8'b00000000; //  724 :   0 - 0x0
      11'h2D5: dout <= 8'b00000000; //  725 :   0 - 0x0
      11'h2D6: dout <= 8'b00000000; //  726 :   0 - 0x0
      11'h2D7: dout <= 8'b00000000; //  727 :   0 - 0x0
      11'h2D8: dout <= 8'b00000000; //  728 :   0 - 0x0 -- Sprite 0x5b
      11'h2D9: dout <= 8'b00000000; //  729 :   0 - 0x0
      11'h2DA: dout <= 8'b00000000; //  730 :   0 - 0x0
      11'h2DB: dout <= 8'b00000001; //  731 :   1 - 0x1
      11'h2DC: dout <= 8'b00000011; //  732 :   3 - 0x3
      11'h2DD: dout <= 8'b00000011; //  733 :   3 - 0x3
      11'h2DE: dout <= 8'b00000111; //  734 :   7 - 0x7
      11'h2DF: dout <= 8'b00111111; //  735 :  63 - 0x3f
      11'h2E0: dout <= 8'b00000000; //  736 :   0 - 0x0 -- Sprite 0x5c
      11'h2E1: dout <= 8'b00000001; //  737 :   1 - 0x1
      11'h2E2: dout <= 8'b01111111; //  738 : 127 - 0x7f
      11'h2E3: dout <= 8'b11111111; //  739 : 255 - 0xff
      11'h2E4: dout <= 8'b11111111; //  740 : 255 - 0xff
      11'h2E5: dout <= 8'b11111111; //  741 : 255 - 0xff
      11'h2E6: dout <= 8'b11111111; //  742 : 255 - 0xff
      11'h2E7: dout <= 8'b11111111; //  743 : 255 - 0xff
      11'h2E8: dout <= 8'b11111111; //  744 : 255 - 0xff -- Sprite 0x5d
      11'h2E9: dout <= 8'b11111111; //  745 : 255 - 0xff
      11'h2EA: dout <= 8'b11111111; //  746 : 255 - 0xff
      11'h2EB: dout <= 8'b11111111; //  747 : 255 - 0xff
      11'h2EC: dout <= 8'b11111111; //  748 : 255 - 0xff
      11'h2ED: dout <= 8'b11111111; //  749 : 255 - 0xff
      11'h2EE: dout <= 8'b11111111; //  750 : 255 - 0xff
      11'h2EF: dout <= 8'b11111111; //  751 : 255 - 0xff
      11'h2F0: dout <= 8'b00000000; //  752 :   0 - 0x0 -- Sprite 0x5e
      11'h2F1: dout <= 8'b10000000; //  753 : 128 - 0x80
      11'h2F2: dout <= 8'b11111110; //  754 : 254 - 0xfe
      11'h2F3: dout <= 8'b11111111; //  755 : 255 - 0xff
      11'h2F4: dout <= 8'b11111111; //  756 : 255 - 0xff
      11'h2F5: dout <= 8'b11111111; //  757 : 255 - 0xff
      11'h2F6: dout <= 8'b11111111; //  758 : 255 - 0xff
      11'h2F7: dout <= 8'b11111111; //  759 : 255 - 0xff
      11'h2F8: dout <= 8'b00000000; //  760 :   0 - 0x0 -- Sprite 0x5f
      11'h2F9: dout <= 8'b00000000; //  761 :   0 - 0x0
      11'h2FA: dout <= 8'b00000000; //  762 :   0 - 0x0
      11'h2FB: dout <= 8'b10000000; //  763 : 128 - 0x80
      11'h2FC: dout <= 8'b11000000; //  764 : 192 - 0xc0
      11'h2FD: dout <= 8'b11000000; //  765 : 192 - 0xc0
      11'h2FE: dout <= 8'b11100000; //  766 : 224 - 0xe0
      11'h2FF: dout <= 8'b11111000; //  767 : 248 - 0xf8
      11'h300: dout <= 8'b11111111; //  768 : 255 - 0xff -- Sprite 0x60
      11'h301: dout <= 8'b11111111; //  769 : 255 - 0xff
      11'h302: dout <= 8'b11111111; //  770 : 255 - 0xff
      11'h303: dout <= 8'b11111111; //  771 : 255 - 0xff
      11'h304: dout <= 8'b11111111; //  772 : 255 - 0xff
      11'h305: dout <= 8'b11111111; //  773 : 255 - 0xff
      11'h306: dout <= 8'b11111111; //  774 : 255 - 0xff
      11'h307: dout <= 8'b11111111; //  775 : 255 - 0xff
      11'h308: dout <= 8'b11111111; //  776 : 255 - 0xff -- Sprite 0x61
      11'h309: dout <= 8'b11111111; //  777 : 255 - 0xff
      11'h30A: dout <= 8'b11111111; //  778 : 255 - 0xff
      11'h30B: dout <= 8'b11111111; //  779 : 255 - 0xff
      11'h30C: dout <= 8'b11111111; //  780 : 255 - 0xff
      11'h30D: dout <= 8'b11111111; //  781 : 255 - 0xff
      11'h30E: dout <= 8'b11111111; //  782 : 255 - 0xff
      11'h30F: dout <= 8'b11111111; //  783 : 255 - 0xff
      11'h310: dout <= 8'b01111000; //  784 : 120 - 0x78 -- Sprite 0x62
      11'h311: dout <= 8'b01100000; //  785 :  96 - 0x60
      11'h312: dout <= 8'b01000000; //  786 :  64 - 0x40
      11'h313: dout <= 8'b01000000; //  787 :  64 - 0x40
      11'h314: dout <= 8'b01000000; //  788 :  64 - 0x40
      11'h315: dout <= 8'b01100000; //  789 :  96 - 0x60
      11'h316: dout <= 8'b00110000; //  790 :  48 - 0x30
      11'h317: dout <= 8'b00011111; //  791 :  31 - 0x1f
      11'h318: dout <= 8'b10000001; //  792 : 129 - 0x81 -- Sprite 0x63
      11'h319: dout <= 8'b10000011; //  793 : 131 - 0x83
      11'h31A: dout <= 8'b11000001; //  794 : 193 - 0xc1
      11'h31B: dout <= 8'b01000011; //  795 :  67 - 0x43
      11'h31C: dout <= 8'b01000001; //  796 :  65 - 0x41
      11'h31D: dout <= 8'b01100011; //  797 :  99 - 0x63
      11'h31E: dout <= 8'b00100110; //  798 :  38 - 0x26
      11'h31F: dout <= 8'b11111000; //  799 : 248 - 0xf8
      11'h320: dout <= 8'b10111001; //  800 : 185 - 0xb9 -- Sprite 0x64
      11'h321: dout <= 8'b10010100; //  801 : 148 - 0x94
      11'h322: dout <= 8'b10001110; //  802 : 142 - 0x8e
      11'h323: dout <= 8'b11000101; //  803 : 197 - 0xc5
      11'h324: dout <= 8'b10010010; //  804 : 146 - 0x92
      11'h325: dout <= 8'b11000111; //  805 : 199 - 0xc7
      11'h326: dout <= 8'b11100010; //  806 : 226 - 0xe2
      11'h327: dout <= 8'b11010000; //  807 : 208 - 0xd0
      11'h328: dout <= 8'b10111001; //  808 : 185 - 0xb9 -- Sprite 0x65
      11'h329: dout <= 8'b00010100; //  809 :  20 - 0x14
      11'h32A: dout <= 8'b10001110; //  810 : 142 - 0x8e
      11'h32B: dout <= 8'b11000101; //  811 : 197 - 0xc5
      11'h32C: dout <= 8'b10010010; //  812 : 146 - 0x92
      11'h32D: dout <= 8'b01000111; //  813 :  71 - 0x47
      11'h32E: dout <= 8'b11100010; //  814 : 226 - 0xe2
      11'h32F: dout <= 8'b01010000; //  815 :  80 - 0x50
      11'h330: dout <= 8'b10111001; //  816 : 185 - 0xb9 -- Sprite 0x66
      11'h331: dout <= 8'b00010101; //  817 :  21 - 0x15
      11'h332: dout <= 8'b10001111; //  818 : 143 - 0x8f
      11'h333: dout <= 8'b11000101; //  819 : 197 - 0xc5
      11'h334: dout <= 8'b10010011; //  820 : 147 - 0x93
      11'h335: dout <= 8'b01000111; //  821 :  71 - 0x47
      11'h336: dout <= 8'b11100011; //  822 : 227 - 0xe3
      11'h337: dout <= 8'b01010001; //  823 :  81 - 0x51
      11'h338: dout <= 8'b01111111; //  824 : 127 - 0x7f -- Sprite 0x67
      11'h339: dout <= 8'b10000000; //  825 : 128 - 0x80
      11'h33A: dout <= 8'b11001100; //  826 : 204 - 0xcc
      11'h33B: dout <= 8'b01111111; //  827 : 127 - 0x7f
      11'h33C: dout <= 8'b00111111; //  828 :  63 - 0x3f
      11'h33D: dout <= 8'b00000011; //  829 :   3 - 0x3
      11'h33E: dout <= 8'b00000000; //  830 :   0 - 0x0
      11'h33F: dout <= 8'b00000000; //  831 :   0 - 0x0
      11'h340: dout <= 8'b11111111; //  832 : 255 - 0xff -- Sprite 0x68
      11'h341: dout <= 8'b00000000; //  833 :   0 - 0x0
      11'h342: dout <= 8'b11001100; //  834 : 204 - 0xcc
      11'h343: dout <= 8'b00110011; //  835 :  51 - 0x33
      11'h344: dout <= 8'b11111111; //  836 : 255 - 0xff
      11'h345: dout <= 8'b11111111; //  837 : 255 - 0xff
      11'h346: dout <= 8'b00000000; //  838 :   0 - 0x0
      11'h347: dout <= 8'b00000000; //  839 :   0 - 0x0
      11'h348: dout <= 8'b11111110; //  840 : 254 - 0xfe -- Sprite 0x69
      11'h349: dout <= 8'b00000001; //  841 :   1 - 0x1
      11'h34A: dout <= 8'b11001101; //  842 : 205 - 0xcd
      11'h34B: dout <= 8'b00111110; //  843 :  62 - 0x3e
      11'h34C: dout <= 8'b11111100; //  844 : 252 - 0xfc
      11'h34D: dout <= 8'b11000000; //  845 : 192 - 0xc0
      11'h34E: dout <= 8'b00000000; //  846 :   0 - 0x0
      11'h34F: dout <= 8'b00000000; //  847 :   0 - 0x0
      11'h350: dout <= 8'b00000000; //  848 :   0 - 0x0 -- Sprite 0x6a
      11'h351: dout <= 8'b00000000; //  849 :   0 - 0x0
      11'h352: dout <= 8'b00000000; //  850 :   0 - 0x0
      11'h353: dout <= 8'b00000000; //  851 :   0 - 0x0
      11'h354: dout <= 8'b00000000; //  852 :   0 - 0x0
      11'h355: dout <= 8'b00000000; //  853 :   0 - 0x0
      11'h356: dout <= 8'b00000000; //  854 :   0 - 0x0
      11'h357: dout <= 8'b00000000; //  855 :   0 - 0x0
      11'h358: dout <= 8'b01111111; //  856 : 127 - 0x7f -- Sprite 0x6b
      11'h359: dout <= 8'b11111111; //  857 : 255 - 0xff
      11'h35A: dout <= 8'b11111111; //  858 : 255 - 0xff
      11'h35B: dout <= 8'b11111111; //  859 : 255 - 0xff
      11'h35C: dout <= 8'b01111111; //  860 : 127 - 0x7f
      11'h35D: dout <= 8'b00110000; //  861 :  48 - 0x30
      11'h35E: dout <= 8'b00001111; //  862 :  15 - 0xf
      11'h35F: dout <= 8'b00000000; //  863 :   0 - 0x0
      11'h360: dout <= 8'b11111111; //  864 : 255 - 0xff -- Sprite 0x6c
      11'h361: dout <= 8'b11111111; //  865 : 255 - 0xff
      11'h362: dout <= 8'b11111111; //  866 : 255 - 0xff
      11'h363: dout <= 8'b11111111; //  867 : 255 - 0xff
      11'h364: dout <= 8'b11111111; //  868 : 255 - 0xff
      11'h365: dout <= 8'b11111110; //  869 : 254 - 0xfe
      11'h366: dout <= 8'b00000001; //  870 :   1 - 0x1
      11'h367: dout <= 8'b11111110; //  871 : 254 - 0xfe
      11'h368: dout <= 8'b00000000; //  872 :   0 - 0x0 -- Sprite 0x6d
      11'h369: dout <= 8'b00000000; //  873 :   0 - 0x0
      11'h36A: dout <= 8'b00000000; //  874 :   0 - 0x0
      11'h36B: dout <= 8'b00000000; //  875 :   0 - 0x0
      11'h36C: dout <= 8'b00000000; //  876 :   0 - 0x0
      11'h36D: dout <= 8'b00000000; //  877 :   0 - 0x0
      11'h36E: dout <= 8'b00000000; //  878 :   0 - 0x0
      11'h36F: dout <= 8'b00000000; //  879 :   0 - 0x0
      11'h370: dout <= 8'b00000000; //  880 :   0 - 0x0 -- Sprite 0x6e
      11'h371: dout <= 8'b00000000; //  881 :   0 - 0x0
      11'h372: dout <= 8'b00000000; //  882 :   0 - 0x0
      11'h373: dout <= 8'b00000000; //  883 :   0 - 0x0
      11'h374: dout <= 8'b00000000; //  884 :   0 - 0x0
      11'h375: dout <= 8'b00000000; //  885 :   0 - 0x0
      11'h376: dout <= 8'b00000000; //  886 :   0 - 0x0
      11'h377: dout <= 8'b00000000; //  887 :   0 - 0x0
      11'h378: dout <= 8'b11111100; //  888 : 252 - 0xfc -- Sprite 0x6f
      11'h379: dout <= 8'b11111110; //  889 : 254 - 0xfe
      11'h37A: dout <= 8'b11111111; //  890 : 255 - 0xff
      11'h37B: dout <= 8'b11111111; //  891 : 255 - 0xff
      11'h37C: dout <= 8'b11110010; //  892 : 242 - 0xf2
      11'h37D: dout <= 8'b00001100; //  893 :  12 - 0xc
      11'h37E: dout <= 8'b11110000; //  894 : 240 - 0xf0
      11'h37F: dout <= 8'b00000000; //  895 :   0 - 0x0
      11'h380: dout <= 8'b01111111; //  896 : 127 - 0x7f -- Sprite 0x70
      11'h381: dout <= 8'b11000000; //  897 : 192 - 0xc0
      11'h382: dout <= 8'b10000000; //  898 : 128 - 0x80
      11'h383: dout <= 8'b10000000; //  899 : 128 - 0x80
      11'h384: dout <= 8'b11100011; //  900 : 227 - 0xe3
      11'h385: dout <= 8'b11111111; //  901 : 255 - 0xff
      11'h386: dout <= 8'b11111111; //  902 : 255 - 0xff
      11'h387: dout <= 8'b11111111; //  903 : 255 - 0xff
      11'h388: dout <= 8'b11111111; //  904 : 255 - 0xff -- Sprite 0x71
      11'h389: dout <= 8'b00000000; //  905 :   0 - 0x0
      11'h38A: dout <= 8'b00000000; //  906 :   0 - 0x0
      11'h38B: dout <= 8'b00000000; //  907 :   0 - 0x0
      11'h38C: dout <= 8'b00000000; //  908 :   0 - 0x0
      11'h38D: dout <= 8'b11000011; //  909 : 195 - 0xc3
      11'h38E: dout <= 8'b11111111; //  910 : 255 - 0xff
      11'h38F: dout <= 8'b11111111; //  911 : 255 - 0xff
      11'h390: dout <= 8'b11111110; //  912 : 254 - 0xfe -- Sprite 0x72
      11'h391: dout <= 8'b00000011; //  913 :   3 - 0x3
      11'h392: dout <= 8'b00000001; //  914 :   1 - 0x1
      11'h393: dout <= 8'b00000001; //  915 :   1 - 0x1
      11'h394: dout <= 8'b11000111; //  916 : 199 - 0xc7
      11'h395: dout <= 8'b11111111; //  917 : 255 - 0xff
      11'h396: dout <= 8'b11111111; //  918 : 255 - 0xff
      11'h397: dout <= 8'b11111111; //  919 : 255 - 0xff
      11'h398: dout <= 8'b11111111; //  920 : 255 - 0xff -- Sprite 0x73
      11'h399: dout <= 8'b11111111; //  921 : 255 - 0xff
      11'h39A: dout <= 8'b11111111; //  922 : 255 - 0xff
      11'h39B: dout <= 8'b11111111; //  923 : 255 - 0xff
      11'h39C: dout <= 8'b11111111; //  924 : 255 - 0xff
      11'h39D: dout <= 8'b11111111; //  925 : 255 - 0xff
      11'h39E: dout <= 8'b11111111; //  926 : 255 - 0xff
      11'h39F: dout <= 8'b11111111; //  927 : 255 - 0xff
      11'h3A0: dout <= 8'b10111001; //  928 : 185 - 0xb9 -- Sprite 0x74
      11'h3A1: dout <= 8'b10010100; //  929 : 148 - 0x94
      11'h3A2: dout <= 8'b10001110; //  930 : 142 - 0x8e
      11'h3A3: dout <= 8'b11000101; //  931 : 197 - 0xc5
      11'h3A4: dout <= 8'b10010010; //  932 : 146 - 0x92
      11'h3A5: dout <= 8'b11000111; //  933 : 199 - 0xc7
      11'h3A6: dout <= 8'b11100010; //  934 : 226 - 0xe2
      11'h3A7: dout <= 8'b01111111; //  935 : 127 - 0x7f
      11'h3A8: dout <= 8'b10111001; //  936 : 185 - 0xb9 -- Sprite 0x75
      11'h3A9: dout <= 8'b00010100; //  937 :  20 - 0x14
      11'h3AA: dout <= 8'b10001110; //  938 : 142 - 0x8e
      11'h3AB: dout <= 8'b11000101; //  939 : 197 - 0xc5
      11'h3AC: dout <= 8'b10010010; //  940 : 146 - 0x92
      11'h3AD: dout <= 8'b01000111; //  941 :  71 - 0x47
      11'h3AE: dout <= 8'b11100010; //  942 : 226 - 0xe2
      11'h3AF: dout <= 8'b11111111; //  943 : 255 - 0xff
      11'h3B0: dout <= 8'b10111001; //  944 : 185 - 0xb9 -- Sprite 0x76
      11'h3B1: dout <= 8'b00010101; //  945 :  21 - 0x15
      11'h3B2: dout <= 8'b10001111; //  946 : 143 - 0x8f
      11'h3B3: dout <= 8'b11000101; //  947 : 197 - 0xc5
      11'h3B4: dout <= 8'b10010011; //  948 : 147 - 0x93
      11'h3B5: dout <= 8'b01000111; //  949 :  71 - 0x47
      11'h3B6: dout <= 8'b11100011; //  950 : 227 - 0xe3
      11'h3B7: dout <= 8'b11111110; //  951 : 254 - 0xfe
      11'h3B8: dout <= 8'b11111111; //  952 : 255 - 0xff -- Sprite 0x77
      11'h3B9: dout <= 8'b11111111; //  953 : 255 - 0xff
      11'h3BA: dout <= 8'b11111111; //  954 : 255 - 0xff
      11'h3BB: dout <= 8'b11111111; //  955 : 255 - 0xff
      11'h3BC: dout <= 8'b11111111; //  956 : 255 - 0xff
      11'h3BD: dout <= 8'b11111111; //  957 : 255 - 0xff
      11'h3BE: dout <= 8'b11111111; //  958 : 255 - 0xff
      11'h3BF: dout <= 8'b11111111; //  959 : 255 - 0xff
      11'h3C0: dout <= 8'b00000000; //  960 :   0 - 0x0 -- Sprite 0x78
      11'h3C1: dout <= 8'b00000000; //  961 :   0 - 0x0
      11'h3C2: dout <= 8'b00000000; //  962 :   0 - 0x0
      11'h3C3: dout <= 8'b00000000; //  963 :   0 - 0x0
      11'h3C4: dout <= 8'b00000000; //  964 :   0 - 0x0
      11'h3C5: dout <= 8'b00000000; //  965 :   0 - 0x0
      11'h3C6: dout <= 8'b00000000; //  966 :   0 - 0x0
      11'h3C7: dout <= 8'b00000000; //  967 :   0 - 0x0
      11'h3C8: dout <= 8'b00000000; //  968 :   0 - 0x0 -- Sprite 0x79
      11'h3C9: dout <= 8'b00000000; //  969 :   0 - 0x0
      11'h3CA: dout <= 8'b00000000; //  970 :   0 - 0x0
      11'h3CB: dout <= 8'b00000000; //  971 :   0 - 0x0
      11'h3CC: dout <= 8'b00000000; //  972 :   0 - 0x0
      11'h3CD: dout <= 8'b00000000; //  973 :   0 - 0x0
      11'h3CE: dout <= 8'b00000000; //  974 :   0 - 0x0
      11'h3CF: dout <= 8'b00000000; //  975 :   0 - 0x0
      11'h3D0: dout <= 8'b00000000; //  976 :   0 - 0x0 -- Sprite 0x7a
      11'h3D1: dout <= 8'b00000000; //  977 :   0 - 0x0
      11'h3D2: dout <= 8'b00000000; //  978 :   0 - 0x0
      11'h3D3: dout <= 8'b00000000; //  979 :   0 - 0x0
      11'h3D4: dout <= 8'b00000000; //  980 :   0 - 0x0
      11'h3D5: dout <= 8'b00000000; //  981 :   0 - 0x0
      11'h3D6: dout <= 8'b00000000; //  982 :   0 - 0x0
      11'h3D7: dout <= 8'b00000000; //  983 :   0 - 0x0
      11'h3D8: dout <= 8'b00000000; //  984 :   0 - 0x0 -- Sprite 0x7b
      11'h3D9: dout <= 8'b00000000; //  985 :   0 - 0x0
      11'h3DA: dout <= 8'b00000000; //  986 :   0 - 0x0
      11'h3DB: dout <= 8'b00000000; //  987 :   0 - 0x0
      11'h3DC: dout <= 8'b00000000; //  988 :   0 - 0x0
      11'h3DD: dout <= 8'b00000000; //  989 :   0 - 0x0
      11'h3DE: dout <= 8'b00000000; //  990 :   0 - 0x0
      11'h3DF: dout <= 8'b00000000; //  991 :   0 - 0x0
      11'h3E0: dout <= 8'b00100010; //  992 :  34 - 0x22 -- Sprite 0x7c
      11'h3E1: dout <= 8'b01010101; //  993 :  85 - 0x55
      11'h3E2: dout <= 8'b10101010; //  994 : 170 - 0xaa
      11'h3E3: dout <= 8'b00000101; //  995 :   5 - 0x5
      11'h3E4: dout <= 8'b00000100; //  996 :   4 - 0x4
      11'h3E5: dout <= 8'b00001010; //  997 :  10 - 0xa
      11'h3E6: dout <= 8'b01010000; //  998 :  80 - 0x50
      11'h3E7: dout <= 8'b00000010; //  999 :   2 - 0x2
      11'h3E8: dout <= 8'b01110011; // 1000 : 115 - 0x73 -- Sprite 0x7d
      11'h3E9: dout <= 8'b11111111; // 1001 : 255 - 0xff
      11'h3EA: dout <= 8'b11111111; // 1002 : 255 - 0xff
      11'h3EB: dout <= 8'b10111101; // 1003 : 189 - 0xbd
      11'h3EC: dout <= 8'b01101110; // 1004 : 110 - 0x6e
      11'h3ED: dout <= 8'b00001010; // 1005 :  10 - 0xa
      11'h3EE: dout <= 8'b01010000; // 1006 :  80 - 0x50
      11'h3EF: dout <= 8'b00000010; // 1007 :   2 - 0x2
      11'h3F0: dout <= 8'b00100000; // 1008 :  32 - 0x20 -- Sprite 0x7e
      11'h3F1: dout <= 8'b01010000; // 1009 :  80 - 0x50
      11'h3F2: dout <= 8'b10000100; // 1010 : 132 - 0x84
      11'h3F3: dout <= 8'b00000000; // 1011 :   0 - 0x0
      11'h3F4: dout <= 8'b00100100; // 1012 :  36 - 0x24
      11'h3F5: dout <= 8'b01011010; // 1013 :  90 - 0x5a
      11'h3F6: dout <= 8'b00010000; // 1014 :  16 - 0x10
      11'h3F7: dout <= 8'b00000000; // 1015 :   0 - 0x0
      11'h3F8: dout <= 8'b11111111; // 1016 : 255 - 0xff -- Sprite 0x7f
      11'h3F9: dout <= 8'b01010000; // 1017 :  80 - 0x50
      11'h3FA: dout <= 8'b10000100; // 1018 : 132 - 0x84
      11'h3FB: dout <= 8'b00000000; // 1019 :   0 - 0x0
      11'h3FC: dout <= 8'b00100100; // 1020 :  36 - 0x24
      11'h3FD: dout <= 8'b01011010; // 1021 :  90 - 0x5a
      11'h3FE: dout <= 8'b00010000; // 1022 :  16 - 0x10
      11'h3FF: dout <= 8'b00000000; // 1023 :   0 - 0x0
      11'h400: dout <= 8'b11111111; // 1024 : 255 - 0xff -- Sprite 0x80
      11'h401: dout <= 8'b10000000; // 1025 : 128 - 0x80
      11'h402: dout <= 8'b11001111; // 1026 : 207 - 0xcf
      11'h403: dout <= 8'b01001000; // 1027 :  72 - 0x48
      11'h404: dout <= 8'b11001111; // 1028 : 207 - 0xcf
      11'h405: dout <= 8'b10000000; // 1029 : 128 - 0x80
      11'h406: dout <= 8'b11001111; // 1030 : 207 - 0xcf
      11'h407: dout <= 8'b01001000; // 1031 :  72 - 0x48
      11'h408: dout <= 8'b11111111; // 1032 : 255 - 0xff -- Sprite 0x81
      11'h409: dout <= 8'b10000000; // 1033 : 128 - 0x80
      11'h40A: dout <= 8'b11111111; // 1034 : 255 - 0xff
      11'h40B: dout <= 8'b10000000; // 1035 : 128 - 0x80
      11'h40C: dout <= 8'b10000000; // 1036 : 128 - 0x80
      11'h40D: dout <= 8'b11011111; // 1037 : 223 - 0xdf
      11'h40E: dout <= 8'b10110000; // 1038 : 176 - 0xb0
      11'h40F: dout <= 8'b11000000; // 1039 : 192 - 0xc0
      11'h410: dout <= 8'b11111111; // 1040 : 255 - 0xff -- Sprite 0x82
      11'h411: dout <= 8'b00000001; // 1041 :   1 - 0x1
      11'h412: dout <= 8'b11110011; // 1042 : 243 - 0xf3
      11'h413: dout <= 8'b00010010; // 1043 :  18 - 0x12
      11'h414: dout <= 8'b11110011; // 1044 : 243 - 0xf3
      11'h415: dout <= 8'b00000001; // 1045 :   1 - 0x1
      11'h416: dout <= 8'b11110011; // 1046 : 243 - 0xf3
      11'h417: dout <= 8'b00010010; // 1047 :  18 - 0x12
      11'h418: dout <= 8'b11111111; // 1048 : 255 - 0xff -- Sprite 0x83
      11'h419: dout <= 8'b00000000; // 1049 :   0 - 0x0
      11'h41A: dout <= 8'b11111111; // 1050 : 255 - 0xff
      11'h41B: dout <= 8'b00000000; // 1051 :   0 - 0x0
      11'h41C: dout <= 8'b00000000; // 1052 :   0 - 0x0
      11'h41D: dout <= 8'b11111111; // 1053 : 255 - 0xff
      11'h41E: dout <= 8'b00000000; // 1054 :   0 - 0x0
      11'h41F: dout <= 8'b00000000; // 1055 :   0 - 0x0
      11'h420: dout <= 8'b11111111; // 1056 : 255 - 0xff -- Sprite 0x84
      11'h421: dout <= 8'b10000010; // 1057 : 130 - 0x82
      11'h422: dout <= 8'b00010000; // 1058 :  16 - 0x10
      11'h423: dout <= 8'b00000000; // 1059 :   0 - 0x0
      11'h424: dout <= 8'b00000000; // 1060 :   0 - 0x0
      11'h425: dout <= 8'b00010000; // 1061 :  16 - 0x10
      11'h426: dout <= 8'b01000100; // 1062 :  68 - 0x44
      11'h427: dout <= 8'b11111111; // 1063 : 255 - 0xff
      11'h428: dout <= 8'b11111111; // 1064 : 255 - 0xff -- Sprite 0x85
      11'h429: dout <= 8'b00000001; // 1065 :   1 - 0x1
      11'h42A: dout <= 8'b11111111; // 1066 : 255 - 0xff
      11'h42B: dout <= 8'b00000001; // 1067 :   1 - 0x1
      11'h42C: dout <= 8'b00000001; // 1068 :   1 - 0x1
      11'h42D: dout <= 8'b11110011; // 1069 : 243 - 0xf3
      11'h42E: dout <= 8'b00001101; // 1070 :  13 - 0xd
      11'h42F: dout <= 8'b00000011; // 1071 :   3 - 0x3
      11'h430: dout <= 8'b00000000; // 1072 :   0 - 0x0 -- Sprite 0x86
      11'h431: dout <= 8'b00000000; // 1073 :   0 - 0x0
      11'h432: dout <= 8'b00000000; // 1074 :   0 - 0x0
      11'h433: dout <= 8'b00000000; // 1075 :   0 - 0x0
      11'h434: dout <= 8'b00000000; // 1076 :   0 - 0x0
      11'h435: dout <= 8'b00000000; // 1077 :   0 - 0x0
      11'h436: dout <= 8'b00000000; // 1078 :   0 - 0x0
      11'h437: dout <= 8'b00000000; // 1079 :   0 - 0x0
      11'h438: dout <= 8'b00000000; // 1080 :   0 - 0x0 -- Sprite 0x87
      11'h439: dout <= 8'b00000000; // 1081 :   0 - 0x0
      11'h43A: dout <= 8'b00000000; // 1082 :   0 - 0x0
      11'h43B: dout <= 8'b00000000; // 1083 :   0 - 0x0
      11'h43C: dout <= 8'b00000000; // 1084 :   0 - 0x0
      11'h43D: dout <= 8'b00000000; // 1085 :   0 - 0x0
      11'h43E: dout <= 8'b00000000; // 1086 :   0 - 0x0
      11'h43F: dout <= 8'b00000000; // 1087 :   0 - 0x0
      11'h440: dout <= 8'b00000111; // 1088 :   7 - 0x7 -- Sprite 0x88
      11'h441: dout <= 8'b00011110; // 1089 :  30 - 0x1e
      11'h442: dout <= 8'b00101111; // 1090 :  47 - 0x2f
      11'h443: dout <= 8'b01010011; // 1091 :  83 - 0x53
      11'h444: dout <= 8'b01101110; // 1092 : 110 - 0x6e
      11'h445: dout <= 8'b11011011; // 1093 : 219 - 0xdb
      11'h446: dout <= 8'b11111010; // 1094 : 250 - 0xfa
      11'h447: dout <= 8'b11010101; // 1095 : 213 - 0xd5
      11'h448: dout <= 8'b10111011; // 1096 : 187 - 0xbb -- Sprite 0x89
      11'h449: dout <= 8'b11110010; // 1097 : 242 - 0xf2
      11'h44A: dout <= 8'b11011101; // 1098 : 221 - 0xdd
      11'h44B: dout <= 8'b01001111; // 1099 :  79 - 0x4f
      11'h44C: dout <= 8'b01111011; // 1100 : 123 - 0x7b
      11'h44D: dout <= 8'b00110010; // 1101 :  50 - 0x32
      11'h44E: dout <= 8'b00011111; // 1102 :  31 - 0x1f
      11'h44F: dout <= 8'b00000111; // 1103 :   7 - 0x7
      11'h450: dout <= 8'b11100000; // 1104 : 224 - 0xe0 -- Sprite 0x8a
      11'h451: dout <= 8'b11011000; // 1105 : 216 - 0xd8
      11'h452: dout <= 8'b01010100; // 1106 :  84 - 0x54
      11'h453: dout <= 8'b11101010; // 1107 : 234 - 0xea
      11'h454: dout <= 8'b10111010; // 1108 : 186 - 0xba
      11'h455: dout <= 8'b10010011; // 1109 : 147 - 0x93
      11'h456: dout <= 8'b11011111; // 1110 : 223 - 0xdf
      11'h457: dout <= 8'b10111101; // 1111 : 189 - 0xbd
      11'h458: dout <= 8'b01101011; // 1112 : 107 - 0x6b -- Sprite 0x8b
      11'h459: dout <= 8'b10011111; // 1113 : 159 - 0x9f
      11'h45A: dout <= 8'b01011101; // 1114 :  93 - 0x5d
      11'h45B: dout <= 8'b10110110; // 1115 : 182 - 0xb6
      11'h45C: dout <= 8'b11101010; // 1116 : 234 - 0xea
      11'h45D: dout <= 8'b11001100; // 1117 : 204 - 0xcc
      11'h45E: dout <= 8'b01111000; // 1118 : 120 - 0x78
      11'h45F: dout <= 8'b11100000; // 1119 : 224 - 0xe0
      11'h460: dout <= 8'b00000111; // 1120 :   7 - 0x7 -- Sprite 0x8c
      11'h461: dout <= 8'b00011000; // 1121 :  24 - 0x18
      11'h462: dout <= 8'b00100011; // 1122 :  35 - 0x23
      11'h463: dout <= 8'b01001100; // 1123 :  76 - 0x4c
      11'h464: dout <= 8'b01110000; // 1124 : 112 - 0x70
      11'h465: dout <= 8'b10100001; // 1125 : 161 - 0xa1
      11'h466: dout <= 8'b10100110; // 1126 : 166 - 0xa6
      11'h467: dout <= 8'b10101000; // 1127 : 168 - 0xa8
      11'h468: dout <= 8'b10100101; // 1128 : 165 - 0xa5 -- Sprite 0x8d
      11'h469: dout <= 8'b10100010; // 1129 : 162 - 0xa2
      11'h46A: dout <= 8'b10010000; // 1130 : 144 - 0x90
      11'h46B: dout <= 8'b01001000; // 1131 :  72 - 0x48
      11'h46C: dout <= 8'b01000111; // 1132 :  71 - 0x47
      11'h46D: dout <= 8'b00100000; // 1133 :  32 - 0x20
      11'h46E: dout <= 8'b00011001; // 1134 :  25 - 0x19
      11'h46F: dout <= 8'b00000111; // 1135 :   7 - 0x7
      11'h470: dout <= 8'b11100000; // 1136 : 224 - 0xe0 -- Sprite 0x8e
      11'h471: dout <= 8'b00011000; // 1137 :  24 - 0x18
      11'h472: dout <= 8'b00000100; // 1138 :   4 - 0x4
      11'h473: dout <= 8'b11000010; // 1139 : 194 - 0xc2
      11'h474: dout <= 8'b00110010; // 1140 :  50 - 0x32
      11'h475: dout <= 8'b00001001; // 1141 :   9 - 0x9
      11'h476: dout <= 8'b11000101; // 1142 : 197 - 0xc5
      11'h477: dout <= 8'b00100101; // 1143 :  37 - 0x25
      11'h478: dout <= 8'b10100101; // 1144 : 165 - 0xa5 -- Sprite 0x8f
      11'h479: dout <= 8'b01100101; // 1145 : 101 - 0x65
      11'h47A: dout <= 8'b01000101; // 1146 :  69 - 0x45
      11'h47B: dout <= 8'b10001010; // 1147 : 138 - 0x8a
      11'h47C: dout <= 8'b10010010; // 1148 : 146 - 0x92
      11'h47D: dout <= 8'b00100100; // 1149 :  36 - 0x24
      11'h47E: dout <= 8'b11011000; // 1150 : 216 - 0xd8
      11'h47F: dout <= 8'b11100000; // 1151 : 224 - 0xe0
      11'h480: dout <= 8'b00000000; // 1152 :   0 - 0x0 -- Sprite 0x90
      11'h481: dout <= 8'b00000000; // 1153 :   0 - 0x0
      11'h482: dout <= 8'b00100000; // 1154 :  32 - 0x20
      11'h483: dout <= 8'b00110000; // 1155 :  48 - 0x30
      11'h484: dout <= 8'b00101100; // 1156 :  44 - 0x2c
      11'h485: dout <= 8'b00100010; // 1157 :  34 - 0x22
      11'h486: dout <= 8'b00010001; // 1158 :  17 - 0x11
      11'h487: dout <= 8'b00001000; // 1159 :   8 - 0x8
      11'h488: dout <= 8'b00000100; // 1160 :   4 - 0x4 -- Sprite 0x91
      11'h489: dout <= 8'b11110010; // 1161 : 242 - 0xf2
      11'h48A: dout <= 8'b11001111; // 1162 : 207 - 0xcf
      11'h48B: dout <= 8'b00110000; // 1163 :  48 - 0x30
      11'h48C: dout <= 8'b00001100; // 1164 :  12 - 0xc
      11'h48D: dout <= 8'b11111111; // 1165 : 255 - 0xff
      11'h48E: dout <= 8'b10000000; // 1166 : 128 - 0x80
      11'h48F: dout <= 8'b11111111; // 1167 : 255 - 0xff
      11'h490: dout <= 8'b01000010; // 1168 :  66 - 0x42 -- Sprite 0x92
      11'h491: dout <= 8'b10100101; // 1169 : 165 - 0xa5
      11'h492: dout <= 8'b10100101; // 1170 : 165 - 0xa5
      11'h493: dout <= 8'b10011001; // 1171 : 153 - 0x99
      11'h494: dout <= 8'b10011001; // 1172 : 153 - 0x99
      11'h495: dout <= 8'b10011001; // 1173 : 153 - 0x99
      11'h496: dout <= 8'b00000001; // 1174 :   1 - 0x1
      11'h497: dout <= 8'b00000000; // 1175 :   0 - 0x0
      11'h498: dout <= 8'b11111111; // 1176 : 255 - 0xff -- Sprite 0x93
      11'h499: dout <= 8'b11111111; // 1177 : 255 - 0xff
      11'h49A: dout <= 8'b11111111; // 1178 : 255 - 0xff
      11'h49B: dout <= 8'b10000001; // 1179 : 129 - 0x81
      11'h49C: dout <= 8'b11111111; // 1180 : 255 - 0xff
      11'h49D: dout <= 8'b11111111; // 1181 : 255 - 0xff
      11'h49E: dout <= 8'b11111111; // 1182 : 255 - 0xff
      11'h49F: dout <= 8'b10000001; // 1183 : 129 - 0x81
      11'h4A0: dout <= 8'b00000000; // 1184 :   0 - 0x0 -- Sprite 0x94
      11'h4A1: dout <= 8'b00000000; // 1185 :   0 - 0x0
      11'h4A2: dout <= 8'b00000100; // 1186 :   4 - 0x4
      11'h4A3: dout <= 8'b00001100; // 1187 :  12 - 0xc
      11'h4A4: dout <= 8'b00110100; // 1188 :  52 - 0x34
      11'h4A5: dout <= 8'b01000100; // 1189 :  68 - 0x44
      11'h4A6: dout <= 8'b10001000; // 1190 : 136 - 0x88
      11'h4A7: dout <= 8'b00010000; // 1191 :  16 - 0x10
      11'h4A8: dout <= 8'b00100000; // 1192 :  32 - 0x20 -- Sprite 0x95
      11'h4A9: dout <= 8'b01001111; // 1193 :  79 - 0x4f
      11'h4AA: dout <= 8'b11110011; // 1194 : 243 - 0xf3
      11'h4AB: dout <= 8'b00001100; // 1195 :  12 - 0xc
      11'h4AC: dout <= 8'b00110000; // 1196 :  48 - 0x30
      11'h4AD: dout <= 8'b11111111; // 1197 : 255 - 0xff
      11'h4AE: dout <= 8'b00000001; // 1198 :   1 - 0x1
      11'h4AF: dout <= 8'b11111111; // 1199 : 255 - 0xff
      11'h4B0: dout <= 8'b01111111; // 1200 : 127 - 0x7f -- Sprite 0x96
      11'h4B1: dout <= 8'b11111111; // 1201 : 255 - 0xff
      11'h4B2: dout <= 8'b11111111; // 1202 : 255 - 0xff
      11'h4B3: dout <= 8'b11111111; // 1203 : 255 - 0xff
      11'h4B4: dout <= 8'b11111011; // 1204 : 251 - 0xfb
      11'h4B5: dout <= 8'b11111111; // 1205 : 255 - 0xff
      11'h4B6: dout <= 8'b11111111; // 1206 : 255 - 0xff
      11'h4B7: dout <= 8'b11111111; // 1207 : 255 - 0xff
      11'h4B8: dout <= 8'b11111111; // 1208 : 255 - 0xff -- Sprite 0x97
      11'h4B9: dout <= 8'b11111111; // 1209 : 255 - 0xff
      11'h4BA: dout <= 8'b11111111; // 1210 : 255 - 0xff
      11'h4BB: dout <= 8'b11111111; // 1211 : 255 - 0xff
      11'h4BC: dout <= 8'b11111111; // 1212 : 255 - 0xff
      11'h4BD: dout <= 8'b11111111; // 1213 : 255 - 0xff
      11'h4BE: dout <= 8'b11111110; // 1214 : 254 - 0xfe
      11'h4BF: dout <= 8'b11111111; // 1215 : 255 - 0xff
      11'h4C0: dout <= 8'b11111111; // 1216 : 255 - 0xff -- Sprite 0x98
      11'h4C1: dout <= 8'b10111111; // 1217 : 191 - 0xbf
      11'h4C2: dout <= 8'b11111111; // 1218 : 255 - 0xff
      11'h4C3: dout <= 8'b11111111; // 1219 : 255 - 0xff
      11'h4C4: dout <= 8'b11111011; // 1220 : 251 - 0xfb
      11'h4C5: dout <= 8'b11111111; // 1221 : 255 - 0xff
      11'h4C6: dout <= 8'b11111111; // 1222 : 255 - 0xff
      11'h4C7: dout <= 8'b11111111; // 1223 : 255 - 0xff
      11'h4C8: dout <= 8'b11111111; // 1224 : 255 - 0xff -- Sprite 0x99
      11'h4C9: dout <= 8'b11111111; // 1225 : 255 - 0xff
      11'h4CA: dout <= 8'b11111111; // 1226 : 255 - 0xff
      11'h4CB: dout <= 8'b11111111; // 1227 : 255 - 0xff
      11'h4CC: dout <= 8'b11111111; // 1228 : 255 - 0xff
      11'h4CD: dout <= 8'b11111111; // 1229 : 255 - 0xff
      11'h4CE: dout <= 8'b11111110; // 1230 : 254 - 0xfe
      11'h4CF: dout <= 8'b11111111; // 1231 : 255 - 0xff
      11'h4D0: dout <= 8'b11111110; // 1232 : 254 - 0xfe -- Sprite 0x9a
      11'h4D1: dout <= 8'b11111111; // 1233 : 255 - 0xff
      11'h4D2: dout <= 8'b11111111; // 1234 : 255 - 0xff
      11'h4D3: dout <= 8'b11111111; // 1235 : 255 - 0xff
      11'h4D4: dout <= 8'b11111011; // 1236 : 251 - 0xfb
      11'h4D5: dout <= 8'b11111111; // 1237 : 255 - 0xff
      11'h4D6: dout <= 8'b11111111; // 1238 : 255 - 0xff
      11'h4D7: dout <= 8'b11111111; // 1239 : 255 - 0xff
      11'h4D8: dout <= 8'b11111111; // 1240 : 255 - 0xff -- Sprite 0x9b
      11'h4D9: dout <= 8'b11111111; // 1241 : 255 - 0xff
      11'h4DA: dout <= 8'b11111111; // 1242 : 255 - 0xff
      11'h4DB: dout <= 8'b11111111; // 1243 : 255 - 0xff
      11'h4DC: dout <= 8'b11111111; // 1244 : 255 - 0xff
      11'h4DD: dout <= 8'b11111111; // 1245 : 255 - 0xff
      11'h4DE: dout <= 8'b11111111; // 1246 : 255 - 0xff
      11'h4DF: dout <= 8'b11111111; // 1247 : 255 - 0xff
      11'h4E0: dout <= 8'b11111111; // 1248 : 255 - 0xff -- Sprite 0x9c
      11'h4E1: dout <= 8'b11111111; // 1249 : 255 - 0xff
      11'h4E2: dout <= 8'b10100000; // 1250 : 160 - 0xa0
      11'h4E3: dout <= 8'b10010000; // 1251 : 144 - 0x90
      11'h4E4: dout <= 8'b10001000; // 1252 : 136 - 0x88
      11'h4E5: dout <= 8'b10000100; // 1253 : 132 - 0x84
      11'h4E6: dout <= 8'b01101010; // 1254 : 106 - 0x6a
      11'h4E7: dout <= 8'b00111111; // 1255 :  63 - 0x3f
      11'h4E8: dout <= 8'b11111111; // 1256 : 255 - 0xff -- Sprite 0x9d
      11'h4E9: dout <= 8'b11111111; // 1257 : 255 - 0xff
      11'h4EA: dout <= 8'b00100001; // 1258 :  33 - 0x21
      11'h4EB: dout <= 8'b00010001; // 1259 :  17 - 0x11
      11'h4EC: dout <= 8'b00001001; // 1260 :   9 - 0x9
      11'h4ED: dout <= 8'b00000101; // 1261 :   5 - 0x5
      11'h4EE: dout <= 8'b10101010; // 1262 : 170 - 0xaa
      11'h4EF: dout <= 8'b11111100; // 1263 : 252 - 0xfc
      11'h4F0: dout <= 8'b11111111; // 1264 : 255 - 0xff -- Sprite 0x9e
      11'h4F1: dout <= 8'b11111111; // 1265 : 255 - 0xff
      11'h4F2: dout <= 8'b00100000; // 1266 :  32 - 0x20
      11'h4F3: dout <= 8'b00010000; // 1267 :  16 - 0x10
      11'h4F4: dout <= 8'b00001000; // 1268 :   8 - 0x8
      11'h4F5: dout <= 8'b00000100; // 1269 :   4 - 0x4
      11'h4F6: dout <= 8'b10101010; // 1270 : 170 - 0xaa
      11'h4F7: dout <= 8'b11111111; // 1271 : 255 - 0xff
      11'h4F8: dout <= 8'b00000000; // 1272 :   0 - 0x0 -- Sprite 0x9f
      11'h4F9: dout <= 8'b00000000; // 1273 :   0 - 0x0
      11'h4FA: dout <= 8'b00000000; // 1274 :   0 - 0x0
      11'h4FB: dout <= 8'b00000000; // 1275 :   0 - 0x0
      11'h4FC: dout <= 8'b00000000; // 1276 :   0 - 0x0
      11'h4FD: dout <= 8'b00000000; // 1277 :   0 - 0x0
      11'h4FE: dout <= 8'b00000000; // 1278 :   0 - 0x0
      11'h4FF: dout <= 8'b00000000; // 1279 :   0 - 0x0
      11'h500: dout <= 8'b11111111; // 1280 : 255 - 0xff -- Sprite 0xa0
      11'h501: dout <= 8'b11010101; // 1281 : 213 - 0xd5
      11'h502: dout <= 8'b11111111; // 1282 : 255 - 0xff
      11'h503: dout <= 8'b00000010; // 1283 :   2 - 0x2
      11'h504: dout <= 8'b00000010; // 1284 :   2 - 0x2
      11'h505: dout <= 8'b00000010; // 1285 :   2 - 0x2
      11'h506: dout <= 8'b00000010; // 1286 :   2 - 0x2
      11'h507: dout <= 8'b00000010; // 1287 :   2 - 0x2
      11'h508: dout <= 8'b00000010; // 1288 :   2 - 0x2 -- Sprite 0xa1
      11'h509: dout <= 8'b00000010; // 1289 :   2 - 0x2
      11'h50A: dout <= 8'b00000010; // 1290 :   2 - 0x2
      11'h50B: dout <= 8'b00000010; // 1291 :   2 - 0x2
      11'h50C: dout <= 8'b00000010; // 1292 :   2 - 0x2
      11'h50D: dout <= 8'b00000010; // 1293 :   2 - 0x2
      11'h50E: dout <= 8'b00000010; // 1294 :   2 - 0x2
      11'h50F: dout <= 8'b00000010; // 1295 :   2 - 0x2
      11'h510: dout <= 8'b11111111; // 1296 : 255 - 0xff -- Sprite 0xa2
      11'h511: dout <= 8'b01010101; // 1297 :  85 - 0x55
      11'h512: dout <= 8'b11111111; // 1298 : 255 - 0xff
      11'h513: dout <= 8'b01000000; // 1299 :  64 - 0x40
      11'h514: dout <= 8'b01000000; // 1300 :  64 - 0x40
      11'h515: dout <= 8'b01000000; // 1301 :  64 - 0x40
      11'h516: dout <= 8'b01000000; // 1302 :  64 - 0x40
      11'h517: dout <= 8'b01000000; // 1303 :  64 - 0x40
      11'h518: dout <= 8'b01000000; // 1304 :  64 - 0x40 -- Sprite 0xa3
      11'h519: dout <= 8'b01000000; // 1305 :  64 - 0x40
      11'h51A: dout <= 8'b01000000; // 1306 :  64 - 0x40
      11'h51B: dout <= 8'b01000000; // 1307 :  64 - 0x40
      11'h51C: dout <= 8'b01000000; // 1308 :  64 - 0x40
      11'h51D: dout <= 8'b01000000; // 1309 :  64 - 0x40
      11'h51E: dout <= 8'b01000000; // 1310 :  64 - 0x40
      11'h51F: dout <= 8'b01000000; // 1311 :  64 - 0x40
      11'h520: dout <= 8'b00110001; // 1312 :  49 - 0x31 -- Sprite 0xa4
      11'h521: dout <= 8'b01001000; // 1313 :  72 - 0x48
      11'h522: dout <= 8'b01000101; // 1314 :  69 - 0x45
      11'h523: dout <= 8'b10000101; // 1315 : 133 - 0x85
      11'h524: dout <= 8'b10000011; // 1316 : 131 - 0x83
      11'h525: dout <= 8'b10000010; // 1317 : 130 - 0x82
      11'h526: dout <= 8'b01100010; // 1318 :  98 - 0x62
      11'h527: dout <= 8'b00010010; // 1319 :  18 - 0x12
      11'h528: dout <= 8'b00110010; // 1320 :  50 - 0x32 -- Sprite 0xa5
      11'h529: dout <= 8'b00100010; // 1321 :  34 - 0x22
      11'h52A: dout <= 8'b01000010; // 1322 :  66 - 0x42
      11'h52B: dout <= 8'b01000000; // 1323 :  64 - 0x40
      11'h52C: dout <= 8'b01000000; // 1324 :  64 - 0x40
      11'h52D: dout <= 8'b00100000; // 1325 :  32 - 0x20
      11'h52E: dout <= 8'b00011110; // 1326 :  30 - 0x1e
      11'h52F: dout <= 8'b00000111; // 1327 :   7 - 0x7
      11'h530: dout <= 8'b10000000; // 1328 : 128 - 0x80 -- Sprite 0xa6
      11'h531: dout <= 8'b11100000; // 1329 : 224 - 0xe0
      11'h532: dout <= 8'b00111000; // 1330 :  56 - 0x38
      11'h533: dout <= 8'b00100100; // 1331 :  36 - 0x24
      11'h534: dout <= 8'b00000100; // 1332 :   4 - 0x4
      11'h535: dout <= 8'b00001000; // 1333 :   8 - 0x8
      11'h536: dout <= 8'b00110000; // 1334 :  48 - 0x30
      11'h537: dout <= 8'b00100000; // 1335 :  32 - 0x20
      11'h538: dout <= 8'b00110000; // 1336 :  48 - 0x30 -- Sprite 0xa7
      11'h539: dout <= 8'b00001000; // 1337 :   8 - 0x8
      11'h53A: dout <= 8'b00001000; // 1338 :   8 - 0x8
      11'h53B: dout <= 8'b00110000; // 1339 :  48 - 0x30
      11'h53C: dout <= 8'b00100000; // 1340 :  32 - 0x20
      11'h53D: dout <= 8'b00100000; // 1341 :  32 - 0x20
      11'h53E: dout <= 8'b00110000; // 1342 :  48 - 0x30
      11'h53F: dout <= 8'b11110000; // 1343 : 240 - 0xf0
      11'h540: dout <= 8'b11111111; // 1344 : 255 - 0xff -- Sprite 0xa8
      11'h541: dout <= 8'b11010010; // 1345 : 210 - 0xd2
      11'h542: dout <= 8'b11110100; // 1346 : 244 - 0xf4
      11'h543: dout <= 8'b11011000; // 1347 : 216 - 0xd8
      11'h544: dout <= 8'b11111000; // 1348 : 248 - 0xf8
      11'h545: dout <= 8'b11010100; // 1349 : 212 - 0xd4
      11'h546: dout <= 8'b11110010; // 1350 : 242 - 0xf2
      11'h547: dout <= 8'b11010001; // 1351 : 209 - 0xd1
      11'h548: dout <= 8'b11110001; // 1352 : 241 - 0xf1 -- Sprite 0xa9
      11'h549: dout <= 8'b11010010; // 1353 : 210 - 0xd2
      11'h54A: dout <= 8'b11110100; // 1354 : 244 - 0xf4
      11'h54B: dout <= 8'b11011000; // 1355 : 216 - 0xd8
      11'h54C: dout <= 8'b11111000; // 1356 : 248 - 0xf8
      11'h54D: dout <= 8'b11010100; // 1357 : 212 - 0xd4
      11'h54E: dout <= 8'b11110010; // 1358 : 242 - 0xf2
      11'h54F: dout <= 8'b11111111; // 1359 : 255 - 0xff
      11'h550: dout <= 8'b11111111; // 1360 : 255 - 0xff -- Sprite 0xaa
      11'h551: dout <= 8'b01000010; // 1361 :  66 - 0x42
      11'h552: dout <= 8'b00100100; // 1362 :  36 - 0x24
      11'h553: dout <= 8'b00011000; // 1363 :  24 - 0x18
      11'h554: dout <= 8'b00011000; // 1364 :  24 - 0x18
      11'h555: dout <= 8'b00100100; // 1365 :  36 - 0x24
      11'h556: dout <= 8'b01000010; // 1366 :  66 - 0x42
      11'h557: dout <= 8'b10000001; // 1367 : 129 - 0x81
      11'h558: dout <= 8'b10000001; // 1368 : 129 - 0x81 -- Sprite 0xab
      11'h559: dout <= 8'b01000010; // 1369 :  66 - 0x42
      11'h55A: dout <= 8'b00100100; // 1370 :  36 - 0x24
      11'h55B: dout <= 8'b00011000; // 1371 :  24 - 0x18
      11'h55C: dout <= 8'b00011000; // 1372 :  24 - 0x18
      11'h55D: dout <= 8'b00100100; // 1373 :  36 - 0x24
      11'h55E: dout <= 8'b01000010; // 1374 :  66 - 0x42
      11'h55F: dout <= 8'b11111111; // 1375 : 255 - 0xff
      11'h560: dout <= 8'b11111111; // 1376 : 255 - 0xff -- Sprite 0xac
      11'h561: dout <= 8'b01001101; // 1377 :  77 - 0x4d
      11'h562: dout <= 8'b00101111; // 1378 :  47 - 0x2f
      11'h563: dout <= 8'b00011101; // 1379 :  29 - 0x1d
      11'h564: dout <= 8'b00011111; // 1380 :  31 - 0x1f
      11'h565: dout <= 8'b00101101; // 1381 :  45 - 0x2d
      11'h566: dout <= 8'b01001111; // 1382 :  79 - 0x4f
      11'h567: dout <= 8'b10001101; // 1383 : 141 - 0x8d
      11'h568: dout <= 8'b10001111; // 1384 : 143 - 0x8f -- Sprite 0xad
      11'h569: dout <= 8'b01001101; // 1385 :  77 - 0x4d
      11'h56A: dout <= 8'b00101111; // 1386 :  47 - 0x2f
      11'h56B: dout <= 8'b00011101; // 1387 :  29 - 0x1d
      11'h56C: dout <= 8'b00011111; // 1388 :  31 - 0x1f
      11'h56D: dout <= 8'b00101101; // 1389 :  45 - 0x2d
      11'h56E: dout <= 8'b01001111; // 1390 :  79 - 0x4f
      11'h56F: dout <= 8'b11111111; // 1391 : 255 - 0xff
      11'h570: dout <= 8'b00000001; // 1392 :   1 - 0x1 -- Sprite 0xae
      11'h571: dout <= 8'b00000011; // 1393 :   3 - 0x3
      11'h572: dout <= 8'b00000110; // 1394 :   6 - 0x6
      11'h573: dout <= 8'b00000111; // 1395 :   7 - 0x7
      11'h574: dout <= 8'b00000111; // 1396 :   7 - 0x7
      11'h575: dout <= 8'b00000111; // 1397 :   7 - 0x7
      11'h576: dout <= 8'b00000110; // 1398 :   6 - 0x6
      11'h577: dout <= 8'b00000111; // 1399 :   7 - 0x7
      11'h578: dout <= 8'b00000110; // 1400 :   6 - 0x6 -- Sprite 0xaf
      11'h579: dout <= 8'b00000110; // 1401 :   6 - 0x6
      11'h57A: dout <= 8'b00001110; // 1402 :  14 - 0xe
      11'h57B: dout <= 8'b00001111; // 1403 :  15 - 0xf
      11'h57C: dout <= 8'b00001110; // 1404 :  14 - 0xe
      11'h57D: dout <= 8'b00011010; // 1405 :  26 - 0x1a
      11'h57E: dout <= 8'b00011011; // 1406 :  27 - 0x1b
      11'h57F: dout <= 8'b00001111; // 1407 :  15 - 0xf
      11'h580: dout <= 8'b00000000; // 1408 :   0 - 0x0 -- Sprite 0xb0
      11'h581: dout <= 8'b11000000; // 1409 : 192 - 0xc0
      11'h582: dout <= 8'b11110000; // 1410 : 240 - 0xf0
      11'h583: dout <= 8'b10001000; // 1411 : 136 - 0x88
      11'h584: dout <= 8'b00010100; // 1412 :  20 - 0x14
      11'h585: dout <= 8'b01101000; // 1413 : 104 - 0x68
      11'h586: dout <= 8'b10101000; // 1414 : 168 - 0xa8
      11'h587: dout <= 8'b00101100; // 1415 :  44 - 0x2c
      11'h588: dout <= 8'b00000100; // 1416 :   4 - 0x4 -- Sprite 0xb1
      11'h589: dout <= 8'b00111000; // 1417 :  56 - 0x38
      11'h58A: dout <= 8'b00010000; // 1418 :  16 - 0x10
      11'h58B: dout <= 8'b10100000; // 1419 : 160 - 0xa0
      11'h58C: dout <= 8'b01100000; // 1420 :  96 - 0x60
      11'h58D: dout <= 8'b00100000; // 1421 :  32 - 0x20
      11'h58E: dout <= 8'b00010000; // 1422 :  16 - 0x10
      11'h58F: dout <= 8'b10001000; // 1423 : 136 - 0x88
      11'h590: dout <= 8'b00001111; // 1424 :  15 - 0xf -- Sprite 0xb2
      11'h591: dout <= 8'b00011011; // 1425 :  27 - 0x1b
      11'h592: dout <= 8'b00011011; // 1426 :  27 - 0x1b
      11'h593: dout <= 8'b00001110; // 1427 :  14 - 0xe
      11'h594: dout <= 8'b00000110; // 1428 :   6 - 0x6
      11'h595: dout <= 8'b00001100; // 1429 :  12 - 0xc
      11'h596: dout <= 8'b00001100; // 1430 :  12 - 0xc
      11'h597: dout <= 8'b00111111; // 1431 :  63 - 0x3f
      11'h598: dout <= 8'b01111111; // 1432 : 127 - 0x7f -- Sprite 0xb3
      11'h599: dout <= 8'b01100000; // 1433 :  96 - 0x60
      11'h59A: dout <= 8'b01100000; // 1434 :  96 - 0x60
      11'h59B: dout <= 8'b01100000; // 1435 :  96 - 0x60
      11'h59C: dout <= 8'b01100000; // 1436 :  96 - 0x60
      11'h59D: dout <= 8'b01100000; // 1437 :  96 - 0x60
      11'h59E: dout <= 8'b01101010; // 1438 : 106 - 0x6a
      11'h59F: dout <= 8'b01111111; // 1439 : 127 - 0x7f
      11'h5A0: dout <= 8'b01001000; // 1440 :  72 - 0x48 -- Sprite 0xb4
      11'h5A1: dout <= 8'b00110000; // 1441 :  48 - 0x30
      11'h5A2: dout <= 8'b00010000; // 1442 :  16 - 0x10
      11'h5A3: dout <= 8'b00010000; // 1443 :  16 - 0x10
      11'h5A4: dout <= 8'b00001000; // 1444 :   8 - 0x8
      11'h5A5: dout <= 8'b00001000; // 1445 :   8 - 0x8
      11'h5A6: dout <= 8'b00001000; // 1446 :   8 - 0x8
      11'h5A7: dout <= 8'b11111100; // 1447 : 252 - 0xfc
      11'h5A8: dout <= 8'b11111110; // 1448 : 254 - 0xfe -- Sprite 0xb5
      11'h5A9: dout <= 8'b00000110; // 1449 :   6 - 0x6
      11'h5AA: dout <= 8'b00000010; // 1450 :   2 - 0x2
      11'h5AB: dout <= 8'b00000110; // 1451 :   6 - 0x6
      11'h5AC: dout <= 8'b00000010; // 1452 :   2 - 0x2
      11'h5AD: dout <= 8'b00000110; // 1453 :   6 - 0x6
      11'h5AE: dout <= 8'b10101010; // 1454 : 170 - 0xaa
      11'h5AF: dout <= 8'b11111110; // 1455 : 254 - 0xfe
      11'h5B0: dout <= 8'b11111111; // 1456 : 255 - 0xff -- Sprite 0xb6
      11'h5B1: dout <= 8'b10000000; // 1457 : 128 - 0x80
      11'h5B2: dout <= 8'b10000000; // 1458 : 128 - 0x80
      11'h5B3: dout <= 8'b10000000; // 1459 : 128 - 0x80
      11'h5B4: dout <= 8'b10000000; // 1460 : 128 - 0x80
      11'h5B5: dout <= 8'b10000000; // 1461 : 128 - 0x80
      11'h5B6: dout <= 8'b10010101; // 1462 : 149 - 0x95
      11'h5B7: dout <= 8'b11111111; // 1463 : 255 - 0xff
      11'h5B8: dout <= 8'b11111111; // 1464 : 255 - 0xff -- Sprite 0xb7
      11'h5B9: dout <= 8'b10000100; // 1465 : 132 - 0x84
      11'h5BA: dout <= 8'b10001100; // 1466 : 140 - 0x8c
      11'h5BB: dout <= 8'b10000100; // 1467 : 132 - 0x84
      11'h5BC: dout <= 8'b10001100; // 1468 : 140 - 0x8c
      11'h5BD: dout <= 8'b10000100; // 1469 : 132 - 0x84
      11'h5BE: dout <= 8'b10101100; // 1470 : 172 - 0xac
      11'h5BF: dout <= 8'b11111111; // 1471 : 255 - 0xff
      11'h5C0: dout <= 8'b11111111; // 1472 : 255 - 0xff -- Sprite 0xb8
      11'h5C1: dout <= 8'b00100001; // 1473 :  33 - 0x21
      11'h5C2: dout <= 8'b01100001; // 1474 :  97 - 0x61
      11'h5C3: dout <= 8'b00100011; // 1475 :  35 - 0x23
      11'h5C4: dout <= 8'b01100001; // 1476 :  97 - 0x61
      11'h5C5: dout <= 8'b00100011; // 1477 :  35 - 0x23
      11'h5C6: dout <= 8'b01100101; // 1478 : 101 - 0x65
      11'h5C7: dout <= 8'b11111111; // 1479 : 255 - 0xff
      11'h5C8: dout <= 8'b11111111; // 1480 : 255 - 0xff -- Sprite 0xb9
      11'h5C9: dout <= 8'b00000001; // 1481 :   1 - 0x1
      11'h5CA: dout <= 8'b00000011; // 1482 :   3 - 0x3
      11'h5CB: dout <= 8'b00000001; // 1483 :   1 - 0x1
      11'h5CC: dout <= 8'b00000011; // 1484 :   3 - 0x3
      11'h5CD: dout <= 8'b00000001; // 1485 :   1 - 0x1
      11'h5CE: dout <= 8'b10101011; // 1486 : 171 - 0xab
      11'h5CF: dout <= 8'b11111111; // 1487 : 255 - 0xff
      11'h5D0: dout <= 8'b11111111; // 1488 : 255 - 0xff -- Sprite 0xba
      11'h5D1: dout <= 8'b11010101; // 1489 : 213 - 0xd5
      11'h5D2: dout <= 8'b10101010; // 1490 : 170 - 0xaa
      11'h5D3: dout <= 8'b11111111; // 1491 : 255 - 0xff
      11'h5D4: dout <= 8'b10000000; // 1492 : 128 - 0x80
      11'h5D5: dout <= 8'b10000000; // 1493 : 128 - 0x80
      11'h5D6: dout <= 8'b10010101; // 1494 : 149 - 0x95
      11'h5D7: dout <= 8'b11111111; // 1495 : 255 - 0xff
      11'h5D8: dout <= 8'b00000000; // 1496 :   0 - 0x0 -- Sprite 0xbb
      11'h5D9: dout <= 8'b00000000; // 1497 :   0 - 0x0
      11'h5DA: dout <= 8'b00000000; // 1498 :   0 - 0x0
      11'h5DB: dout <= 8'b00000000; // 1499 :   0 - 0x0
      11'h5DC: dout <= 8'b00000000; // 1500 :   0 - 0x0
      11'h5DD: dout <= 8'b00000000; // 1501 :   0 - 0x0
      11'h5DE: dout <= 8'b00000000; // 1502 :   0 - 0x0
      11'h5DF: dout <= 8'b00000000; // 1503 :   0 - 0x0
      11'h5E0: dout <= 8'b11111111; // 1504 : 255 - 0xff -- Sprite 0xbc
      11'h5E1: dout <= 8'b01010101; // 1505 :  85 - 0x55
      11'h5E2: dout <= 8'b10101011; // 1506 : 171 - 0xab
      11'h5E3: dout <= 8'b11111111; // 1507 : 255 - 0xff
      11'h5E4: dout <= 8'b01100001; // 1508 :  97 - 0x61
      11'h5E5: dout <= 8'b00100011; // 1509 :  35 - 0x23
      11'h5E6: dout <= 8'b01100101; // 1510 : 101 - 0x65
      11'h5E7: dout <= 8'b11111111; // 1511 : 255 - 0xff
      11'h5E8: dout <= 8'b00000000; // 1512 :   0 - 0x0 -- Sprite 0xbd
      11'h5E9: dout <= 8'b00000000; // 1513 :   0 - 0x0
      11'h5EA: dout <= 8'b00000000; // 1514 :   0 - 0x0
      11'h5EB: dout <= 8'b00000000; // 1515 :   0 - 0x0
      11'h5EC: dout <= 8'b00000000; // 1516 :   0 - 0x0
      11'h5ED: dout <= 8'b00000000; // 1517 :   0 - 0x0
      11'h5EE: dout <= 8'b00000000; // 1518 :   0 - 0x0
      11'h5EF: dout <= 8'b00000000; // 1519 :   0 - 0x0
      11'h5F0: dout <= 8'b00000000; // 1520 :   0 - 0x0 -- Sprite 0xbe
      11'h5F1: dout <= 8'b00000000; // 1521 :   0 - 0x0
      11'h5F2: dout <= 8'b00000000; // 1522 :   0 - 0x0
      11'h5F3: dout <= 8'b00000000; // 1523 :   0 - 0x0
      11'h5F4: dout <= 8'b00000000; // 1524 :   0 - 0x0
      11'h5F5: dout <= 8'b00000000; // 1525 :   0 - 0x0
      11'h5F6: dout <= 8'b00000000; // 1526 :   0 - 0x0
      11'h5F7: dout <= 8'b00000000; // 1527 :   0 - 0x0
      11'h5F8: dout <= 8'b00000000; // 1528 :   0 - 0x0 -- Sprite 0xbf
      11'h5F9: dout <= 8'b00000000; // 1529 :   0 - 0x0
      11'h5FA: dout <= 8'b00000000; // 1530 :   0 - 0x0
      11'h5FB: dout <= 8'b00000000; // 1531 :   0 - 0x0
      11'h5FC: dout <= 8'b00000000; // 1532 :   0 - 0x0
      11'h5FD: dout <= 8'b00000000; // 1533 :   0 - 0x0
      11'h5FE: dout <= 8'b00000000; // 1534 :   0 - 0x0
      11'h5FF: dout <= 8'b00000000; // 1535 :   0 - 0x0
      11'h600: dout <= 8'b00000000; // 1536 :   0 - 0x0 -- Sprite 0xc0
      11'h601: dout <= 8'b00000000; // 1537 :   0 - 0x0
      11'h602: dout <= 8'b00000000; // 1538 :   0 - 0x0
      11'h603: dout <= 8'b00000000; // 1539 :   0 - 0x0
      11'h604: dout <= 8'b00000000; // 1540 :   0 - 0x0
      11'h605: dout <= 8'b00000000; // 1541 :   0 - 0x0
      11'h606: dout <= 8'b00000000; // 1542 :   0 - 0x0
      11'h607: dout <= 8'b00000000; // 1543 :   0 - 0x0
      11'h608: dout <= 8'b00000000; // 1544 :   0 - 0x0 -- Sprite 0xc1
      11'h609: dout <= 8'b00000000; // 1545 :   0 - 0x0
      11'h60A: dout <= 8'b00000000; // 1546 :   0 - 0x0
      11'h60B: dout <= 8'b00000000; // 1547 :   0 - 0x0
      11'h60C: dout <= 8'b00000000; // 1548 :   0 - 0x0
      11'h60D: dout <= 8'b00000000; // 1549 :   0 - 0x0
      11'h60E: dout <= 8'b00000000; // 1550 :   0 - 0x0
      11'h60F: dout <= 8'b00000000; // 1551 :   0 - 0x0
      11'h610: dout <= 8'b00000000; // 1552 :   0 - 0x0 -- Sprite 0xc2
      11'h611: dout <= 8'b00000000; // 1553 :   0 - 0x0
      11'h612: dout <= 8'b00000000; // 1554 :   0 - 0x0
      11'h613: dout <= 8'b00000000; // 1555 :   0 - 0x0
      11'h614: dout <= 8'b00000000; // 1556 :   0 - 0x0
      11'h615: dout <= 8'b00000000; // 1557 :   0 - 0x0
      11'h616: dout <= 8'b00000000; // 1558 :   0 - 0x0
      11'h617: dout <= 8'b00000000; // 1559 :   0 - 0x0
      11'h618: dout <= 8'b00000000; // 1560 :   0 - 0x0 -- Sprite 0xc3
      11'h619: dout <= 8'b00000000; // 1561 :   0 - 0x0
      11'h61A: dout <= 8'b00000000; // 1562 :   0 - 0x0
      11'h61B: dout <= 8'b00000000; // 1563 :   0 - 0x0
      11'h61C: dout <= 8'b00000000; // 1564 :   0 - 0x0
      11'h61D: dout <= 8'b00000000; // 1565 :   0 - 0x0
      11'h61E: dout <= 8'b00000000; // 1566 :   0 - 0x0
      11'h61F: dout <= 8'b00000000; // 1567 :   0 - 0x0
      11'h620: dout <= 8'b00000000; // 1568 :   0 - 0x0 -- Sprite 0xc4
      11'h621: dout <= 8'b00000000; // 1569 :   0 - 0x0
      11'h622: dout <= 8'b00000000; // 1570 :   0 - 0x0
      11'h623: dout <= 8'b00000000; // 1571 :   0 - 0x0
      11'h624: dout <= 8'b00000000; // 1572 :   0 - 0x0
      11'h625: dout <= 8'b00000000; // 1573 :   0 - 0x0
      11'h626: dout <= 8'b00000000; // 1574 :   0 - 0x0
      11'h627: dout <= 8'b00000000; // 1575 :   0 - 0x0
      11'h628: dout <= 8'b00000000; // 1576 :   0 - 0x0 -- Sprite 0xc5
      11'h629: dout <= 8'b00000000; // 1577 :   0 - 0x0
      11'h62A: dout <= 8'b00000001; // 1578 :   1 - 0x1
      11'h62B: dout <= 8'b00000110; // 1579 :   6 - 0x6
      11'h62C: dout <= 8'b00001010; // 1580 :  10 - 0xa
      11'h62D: dout <= 8'b00010100; // 1581 :  20 - 0x14
      11'h62E: dout <= 8'b00010000; // 1582 :  16 - 0x10
      11'h62F: dout <= 8'b00101000; // 1583 :  40 - 0x28
      11'h630: dout <= 8'b00011111; // 1584 :  31 - 0x1f -- Sprite 0xc6
      11'h631: dout <= 8'b01100000; // 1585 :  96 - 0x60
      11'h632: dout <= 8'b10100000; // 1586 : 160 - 0xa0
      11'h633: dout <= 8'b01000000; // 1587 :  64 - 0x40
      11'h634: dout <= 8'b00000000; // 1588 :   0 - 0x0
      11'h635: dout <= 8'b00000000; // 1589 :   0 - 0x0
      11'h636: dout <= 8'b00000000; // 1590 :   0 - 0x0
      11'h637: dout <= 8'b00000000; // 1591 :   0 - 0x0
      11'h638: dout <= 8'b00110000; // 1592 :  48 - 0x30 -- Sprite 0xc7
      11'h639: dout <= 8'b01000000; // 1593 :  64 - 0x40
      11'h63A: dout <= 8'b01100000; // 1594 :  96 - 0x60
      11'h63B: dout <= 8'b11000000; // 1595 : 192 - 0xc0
      11'h63C: dout <= 8'b10000000; // 1596 : 128 - 0x80
      11'h63D: dout <= 8'b10100000; // 1597 : 160 - 0xa0
      11'h63E: dout <= 8'b11000000; // 1598 : 192 - 0xc0
      11'h63F: dout <= 8'b10000000; // 1599 : 128 - 0x80
      11'h640: dout <= 8'b11111111; // 1600 : 255 - 0xff -- Sprite 0xc8
      11'h641: dout <= 8'b00000000; // 1601 :   0 - 0x0
      11'h642: dout <= 8'b00000000; // 1602 :   0 - 0x0
      11'h643: dout <= 8'b00000000; // 1603 :   0 - 0x0
      11'h644: dout <= 8'b00000000; // 1604 :   0 - 0x0
      11'h645: dout <= 8'b00000000; // 1605 :   0 - 0x0
      11'h646: dout <= 8'b00000000; // 1606 :   0 - 0x0
      11'h647: dout <= 8'b00000000; // 1607 :   0 - 0x0
      11'h648: dout <= 8'b00010100; // 1608 :  20 - 0x14 -- Sprite 0xc9
      11'h649: dout <= 8'b00101010; // 1609 :  42 - 0x2a
      11'h64A: dout <= 8'b00010110; // 1610 :  22 - 0x16
      11'h64B: dout <= 8'b00101011; // 1611 :  43 - 0x2b
      11'h64C: dout <= 8'b00010101; // 1612 :  21 - 0x15
      11'h64D: dout <= 8'b00101011; // 1613 :  43 - 0x2b
      11'h64E: dout <= 8'b00010101; // 1614 :  21 - 0x15
      11'h64F: dout <= 8'b00101011; // 1615 :  43 - 0x2b
      11'h650: dout <= 8'b00000000; // 1616 :   0 - 0x0 -- Sprite 0xca
      11'h651: dout <= 8'b00000100; // 1617 :   4 - 0x4
      11'h652: dout <= 8'b00000100; // 1618 :   4 - 0x4
      11'h653: dout <= 8'b00000101; // 1619 :   5 - 0x5
      11'h654: dout <= 8'b00010101; // 1620 :  21 - 0x15
      11'h655: dout <= 8'b00010101; // 1621 :  21 - 0x15
      11'h656: dout <= 8'b01010101; // 1622 :  85 - 0x55
      11'h657: dout <= 8'b01010101; // 1623 :  85 - 0x55
      11'h658: dout <= 8'b00000000; // 1624 :   0 - 0x0 -- Sprite 0xcb
      11'h659: dout <= 8'b00000000; // 1625 :   0 - 0x0
      11'h65A: dout <= 8'b00010000; // 1626 :  16 - 0x10
      11'h65B: dout <= 8'b00010000; // 1627 :  16 - 0x10
      11'h65C: dout <= 8'b01010001; // 1628 :  81 - 0x51
      11'h65D: dout <= 8'b01010101; // 1629 :  85 - 0x55
      11'h65E: dout <= 8'b01010101; // 1630 :  85 - 0x55
      11'h65F: dout <= 8'b01010101; // 1631 :  85 - 0x55
      11'h660: dout <= 8'b00000000; // 1632 :   0 - 0x0 -- Sprite 0xcc
      11'h661: dout <= 8'b00000000; // 1633 :   0 - 0x0
      11'h662: dout <= 8'b00000000; // 1634 :   0 - 0x0
      11'h663: dout <= 8'b00000101; // 1635 :   5 - 0x5
      11'h664: dout <= 8'b00001111; // 1636 :  15 - 0xf
      11'h665: dout <= 8'b00000111; // 1637 :   7 - 0x7
      11'h666: dout <= 8'b00000011; // 1638 :   3 - 0x3
      11'h667: dout <= 8'b00000001; // 1639 :   1 - 0x1
      11'h668: dout <= 8'b00000000; // 1640 :   0 - 0x0 -- Sprite 0xcd
      11'h669: dout <= 8'b00000000; // 1641 :   0 - 0x0
      11'h66A: dout <= 8'b10000000; // 1642 : 128 - 0x80
      11'h66B: dout <= 8'b11010000; // 1643 : 208 - 0xd0
      11'h66C: dout <= 8'b11111000; // 1644 : 248 - 0xf8
      11'h66D: dout <= 8'b11110000; // 1645 : 240 - 0xf0
      11'h66E: dout <= 8'b11100000; // 1646 : 224 - 0xe0
      11'h66F: dout <= 8'b11000000; // 1647 : 192 - 0xc0
      11'h670: dout <= 8'b00000000; // 1648 :   0 - 0x0 -- Sprite 0xce
      11'h671: dout <= 8'b00000000; // 1649 :   0 - 0x0
      11'h672: dout <= 8'b00000000; // 1650 :   0 - 0x0
      11'h673: dout <= 8'b01111000; // 1651 : 120 - 0x78
      11'h674: dout <= 8'b11001111; // 1652 : 207 - 0xcf
      11'h675: dout <= 8'b10000000; // 1653 : 128 - 0x80
      11'h676: dout <= 8'b11001111; // 1654 : 207 - 0xcf
      11'h677: dout <= 8'b01001000; // 1655 :  72 - 0x48
      11'h678: dout <= 8'b00000000; // 1656 :   0 - 0x0 -- Sprite 0xcf
      11'h679: dout <= 8'b00000000; // 1657 :   0 - 0x0
      11'h67A: dout <= 8'b00000000; // 1658 :   0 - 0x0
      11'h67B: dout <= 8'b00011110; // 1659 :  30 - 0x1e
      11'h67C: dout <= 8'b11110011; // 1660 : 243 - 0xf3
      11'h67D: dout <= 8'b00000001; // 1661 :   1 - 0x1
      11'h67E: dout <= 8'b11110011; // 1662 : 243 - 0xf3
      11'h67F: dout <= 8'b00010010; // 1663 :  18 - 0x12
      11'h680: dout <= 8'b00000000; // 1664 :   0 - 0x0 -- Sprite 0xd0
      11'h681: dout <= 8'b00000000; // 1665 :   0 - 0x0
      11'h682: dout <= 8'b00000000; // 1666 :   0 - 0x0
      11'h683: dout <= 8'b00000000; // 1667 :   0 - 0x0
      11'h684: dout <= 8'b00000000; // 1668 :   0 - 0x0
      11'h685: dout <= 8'b00000000; // 1669 :   0 - 0x0
      11'h686: dout <= 8'b00000000; // 1670 :   0 - 0x0
      11'h687: dout <= 8'b00000000; // 1671 :   0 - 0x0
      11'h688: dout <= 8'b00000000; // 1672 :   0 - 0x0 -- Sprite 0xd1
      11'h689: dout <= 8'b00000000; // 1673 :   0 - 0x0
      11'h68A: dout <= 8'b00000000; // 1674 :   0 - 0x0
      11'h68B: dout <= 8'b00000000; // 1675 :   0 - 0x0
      11'h68C: dout <= 8'b00000000; // 1676 :   0 - 0x0
      11'h68D: dout <= 8'b00000000; // 1677 :   0 - 0x0
      11'h68E: dout <= 8'b00000000; // 1678 :   0 - 0x0
      11'h68F: dout <= 8'b00000000; // 1679 :   0 - 0x0
      11'h690: dout <= 8'b00001000; // 1680 :   8 - 0x8 -- Sprite 0xd2
      11'h691: dout <= 8'b00001100; // 1681 :  12 - 0xc
      11'h692: dout <= 8'b00001000; // 1682 :   8 - 0x8
      11'h693: dout <= 8'b00001000; // 1683 :   8 - 0x8
      11'h694: dout <= 8'b00001010; // 1684 :  10 - 0xa
      11'h695: dout <= 8'b00001000; // 1685 :   8 - 0x8
      11'h696: dout <= 8'b00001000; // 1686 :   8 - 0x8
      11'h697: dout <= 8'b00001100; // 1687 :  12 - 0xc
      11'h698: dout <= 8'b00010000; // 1688 :  16 - 0x10 -- Sprite 0xd3
      11'h699: dout <= 8'b00010000; // 1689 :  16 - 0x10
      11'h69A: dout <= 8'b00110000; // 1690 :  48 - 0x30
      11'h69B: dout <= 8'b00010000; // 1691 :  16 - 0x10
      11'h69C: dout <= 8'b01010000; // 1692 :  80 - 0x50
      11'h69D: dout <= 8'b00010000; // 1693 :  16 - 0x10
      11'h69E: dout <= 8'b00110000; // 1694 :  48 - 0x30
      11'h69F: dout <= 8'b00010000; // 1695 :  16 - 0x10
      11'h6A0: dout <= 8'b00000000; // 1696 :   0 - 0x0 -- Sprite 0xd4
      11'h6A1: dout <= 8'b00000000; // 1697 :   0 - 0x0
      11'h6A2: dout <= 8'b00000000; // 1698 :   0 - 0x0
      11'h6A3: dout <= 8'b00000000; // 1699 :   0 - 0x0
      11'h6A4: dout <= 8'b00000000; // 1700 :   0 - 0x0
      11'h6A5: dout <= 8'b00000000; // 1701 :   0 - 0x0
      11'h6A6: dout <= 8'b00000000; // 1702 :   0 - 0x0
      11'h6A7: dout <= 8'b00000000; // 1703 :   0 - 0x0
      11'h6A8: dout <= 8'b11111000; // 1704 : 248 - 0xf8 -- Sprite 0xd5
      11'h6A9: dout <= 8'b00000110; // 1705 :   6 - 0x6
      11'h6AA: dout <= 8'b00000001; // 1706 :   1 - 0x1
      11'h6AB: dout <= 8'b00000000; // 1707 :   0 - 0x0
      11'h6AC: dout <= 8'b00000000; // 1708 :   0 - 0x0
      11'h6AD: dout <= 8'b00000000; // 1709 :   0 - 0x0
      11'h6AE: dout <= 8'b00000000; // 1710 :   0 - 0x0
      11'h6AF: dout <= 8'b00000000; // 1711 :   0 - 0x0
      11'h6B0: dout <= 8'b00000000; // 1712 :   0 - 0x0 -- Sprite 0xd6
      11'h6B1: dout <= 8'b00000000; // 1713 :   0 - 0x0
      11'h6B2: dout <= 8'b10000000; // 1714 : 128 - 0x80
      11'h6B3: dout <= 8'b01100000; // 1715 :  96 - 0x60
      11'h6B4: dout <= 8'b01010000; // 1716 :  80 - 0x50
      11'h6B5: dout <= 8'b10101000; // 1717 : 168 - 0xa8
      11'h6B6: dout <= 8'b01011000; // 1718 :  88 - 0x58
      11'h6B7: dout <= 8'b00101100; // 1719 :  44 - 0x2c
      11'h6B8: dout <= 8'b10100000; // 1720 : 160 - 0xa0 -- Sprite 0xd7
      11'h6B9: dout <= 8'b11000000; // 1721 : 192 - 0xc0
      11'h6BA: dout <= 8'b10000000; // 1722 : 128 - 0x80
      11'h6BB: dout <= 8'b01010000; // 1723 :  80 - 0x50
      11'h6BC: dout <= 8'b01100000; // 1724 :  96 - 0x60
      11'h6BD: dout <= 8'b00111000; // 1725 :  56 - 0x38
      11'h6BE: dout <= 8'b00001000; // 1726 :   8 - 0x8
      11'h6BF: dout <= 8'b00000111; // 1727 :   7 - 0x7
      11'h6C0: dout <= 8'b00000000; // 1728 :   0 - 0x0 -- Sprite 0xd8
      11'h6C1: dout <= 8'b00000000; // 1729 :   0 - 0x0
      11'h6C2: dout <= 8'b00000000; // 1730 :   0 - 0x0
      11'h6C3: dout <= 8'b00000000; // 1731 :   0 - 0x0
      11'h6C4: dout <= 8'b00000000; // 1732 :   0 - 0x0
      11'h6C5: dout <= 8'b00000000; // 1733 :   0 - 0x0
      11'h6C6: dout <= 8'b00000000; // 1734 :   0 - 0x0
      11'h6C7: dout <= 8'b11111111; // 1735 : 255 - 0xff
      11'h6C8: dout <= 8'b00010101; // 1736 :  21 - 0x15 -- Sprite 0xd9
      11'h6C9: dout <= 8'b00101011; // 1737 :  43 - 0x2b
      11'h6CA: dout <= 8'b00010101; // 1738 :  21 - 0x15
      11'h6CB: dout <= 8'b00101010; // 1739 :  42 - 0x2a
      11'h6CC: dout <= 8'b01010110; // 1740 :  86 - 0x56
      11'h6CD: dout <= 8'b10101100; // 1741 : 172 - 0xac
      11'h6CE: dout <= 8'b01010000; // 1742 :  80 - 0x50
      11'h6CF: dout <= 8'b11100000; // 1743 : 224 - 0xe0
      11'h6D0: dout <= 8'b00000001; // 1744 :   1 - 0x1 -- Sprite 0xda
      11'h6D1: dout <= 8'b00001101; // 1745 :  13 - 0xd
      11'h6D2: dout <= 8'b00010011; // 1746 :  19 - 0x13
      11'h6D3: dout <= 8'b00001101; // 1747 :  13 - 0xd
      11'h6D4: dout <= 8'b00000001; // 1748 :   1 - 0x1
      11'h6D5: dout <= 8'b00000001; // 1749 :   1 - 0x1
      11'h6D6: dout <= 8'b00000001; // 1750 :   1 - 0x1
      11'h6D7: dout <= 8'b00000001; // 1751 :   1 - 0x1
      11'h6D8: dout <= 8'b11000000; // 1752 : 192 - 0xc0 -- Sprite 0xdb
      11'h6D9: dout <= 8'b01000000; // 1753 :  64 - 0x40
      11'h6DA: dout <= 8'b01000000; // 1754 :  64 - 0x40
      11'h6DB: dout <= 8'b01011000; // 1755 :  88 - 0x58
      11'h6DC: dout <= 8'b01100100; // 1756 : 100 - 0x64
      11'h6DD: dout <= 8'b01011000; // 1757 :  88 - 0x58
      11'h6DE: dout <= 8'b01000000; // 1758 :  64 - 0x40
      11'h6DF: dout <= 8'b01000000; // 1759 :  64 - 0x40
      11'h6E0: dout <= 8'b00000000; // 1760 :   0 - 0x0 -- Sprite 0xdc
      11'h6E1: dout <= 8'b00000000; // 1761 :   0 - 0x0
      11'h6E2: dout <= 8'b00000000; // 1762 :   0 - 0x0
      11'h6E3: dout <= 8'b00000110; // 1763 :   6 - 0x6
      11'h6E4: dout <= 8'b00000111; // 1764 :   7 - 0x7
      11'h6E5: dout <= 8'b00000111; // 1765 :   7 - 0x7
      11'h6E6: dout <= 8'b00000111; // 1766 :   7 - 0x7
      11'h6E7: dout <= 8'b00000011; // 1767 :   3 - 0x3
      11'h6E8: dout <= 8'b00000000; // 1768 :   0 - 0x0 -- Sprite 0xdd
      11'h6E9: dout <= 8'b00000000; // 1769 :   0 - 0x0
      11'h6EA: dout <= 8'b00000000; // 1770 :   0 - 0x0
      11'h6EB: dout <= 8'b10110000; // 1771 : 176 - 0xb0
      11'h6EC: dout <= 8'b11110000; // 1772 : 240 - 0xf0
      11'h6ED: dout <= 8'b11110000; // 1773 : 240 - 0xf0
      11'h6EE: dout <= 8'b11110000; // 1774 : 240 - 0xf0
      11'h6EF: dout <= 8'b11100000; // 1775 : 224 - 0xe0
      11'h6F0: dout <= 8'b11001111; // 1776 : 207 - 0xcf -- Sprite 0xde
      11'h6F1: dout <= 8'b10000000; // 1777 : 128 - 0x80
      11'h6F2: dout <= 8'b11001111; // 1778 : 207 - 0xcf
      11'h6F3: dout <= 8'b01001000; // 1779 :  72 - 0x48
      11'h6F4: dout <= 8'b01001000; // 1780 :  72 - 0x48
      11'h6F5: dout <= 8'b01001000; // 1781 :  72 - 0x48
      11'h6F6: dout <= 8'b01001000; // 1782 :  72 - 0x48
      11'h6F7: dout <= 8'b01001000; // 1783 :  72 - 0x48
      11'h6F8: dout <= 8'b11110011; // 1784 : 243 - 0xf3 -- Sprite 0xdf
      11'h6F9: dout <= 8'b00000001; // 1785 :   1 - 0x1
      11'h6FA: dout <= 8'b11110011; // 1786 : 243 - 0xf3
      11'h6FB: dout <= 8'b00010010; // 1787 :  18 - 0x12
      11'h6FC: dout <= 8'b00010010; // 1788 :  18 - 0x12
      11'h6FD: dout <= 8'b00010010; // 1789 :  18 - 0x12
      11'h6FE: dout <= 8'b00010010; // 1790 :  18 - 0x12
      11'h6FF: dout <= 8'b00010010; // 1791 :  18 - 0x12
      11'h700: dout <= 8'b00000000; // 1792 :   0 - 0x0 -- Sprite 0xe0
      11'h701: dout <= 8'b00000000; // 1793 :   0 - 0x0
      11'h702: dout <= 8'b00000000; // 1794 :   0 - 0x0
      11'h703: dout <= 8'b00000000; // 1795 :   0 - 0x0
      11'h704: dout <= 8'b00000000; // 1796 :   0 - 0x0
      11'h705: dout <= 8'b00000000; // 1797 :   0 - 0x0
      11'h706: dout <= 8'b00000000; // 1798 :   0 - 0x0
      11'h707: dout <= 8'b00000000; // 1799 :   0 - 0x0
      11'h708: dout <= 8'b00000000; // 1800 :   0 - 0x0 -- Sprite 0xe1
      11'h709: dout <= 8'b00000000; // 1801 :   0 - 0x0
      11'h70A: dout <= 8'b00000000; // 1802 :   0 - 0x0
      11'h70B: dout <= 8'b00000000; // 1803 :   0 - 0x0
      11'h70C: dout <= 8'b00000000; // 1804 :   0 - 0x0
      11'h70D: dout <= 8'b00000000; // 1805 :   0 - 0x0
      11'h70E: dout <= 8'b00000000; // 1806 :   0 - 0x0
      11'h70F: dout <= 8'b00000000; // 1807 :   0 - 0x0
      11'h710: dout <= 8'b00000000; // 1808 :   0 - 0x0 -- Sprite 0xe2
      11'h711: dout <= 8'b00000000; // 1809 :   0 - 0x0
      11'h712: dout <= 8'b00000000; // 1810 :   0 - 0x0
      11'h713: dout <= 8'b00000000; // 1811 :   0 - 0x0
      11'h714: dout <= 8'b00000000; // 1812 :   0 - 0x0
      11'h715: dout <= 8'b00000000; // 1813 :   0 - 0x0
      11'h716: dout <= 8'b00000000; // 1814 :   0 - 0x0
      11'h717: dout <= 8'b00000000; // 1815 :   0 - 0x0
      11'h718: dout <= 8'b00000000; // 1816 :   0 - 0x0 -- Sprite 0xe3
      11'h719: dout <= 8'b00000000; // 1817 :   0 - 0x0
      11'h71A: dout <= 8'b00000000; // 1818 :   0 - 0x0
      11'h71B: dout <= 8'b00000000; // 1819 :   0 - 0x0
      11'h71C: dout <= 8'b00000000; // 1820 :   0 - 0x0
      11'h71D: dout <= 8'b00000000; // 1821 :   0 - 0x0
      11'h71E: dout <= 8'b00000000; // 1822 :   0 - 0x0
      11'h71F: dout <= 8'b00000000; // 1823 :   0 - 0x0
      11'h720: dout <= 8'b00000000; // 1824 :   0 - 0x0 -- Sprite 0xe4
      11'h721: dout <= 8'b00000000; // 1825 :   0 - 0x0
      11'h722: dout <= 8'b00000000; // 1826 :   0 - 0x0
      11'h723: dout <= 8'b00000000; // 1827 :   0 - 0x0
      11'h724: dout <= 8'b00000000; // 1828 :   0 - 0x0
      11'h725: dout <= 8'b00000000; // 1829 :   0 - 0x0
      11'h726: dout <= 8'b00000000; // 1830 :   0 - 0x0
      11'h727: dout <= 8'b00000000; // 1831 :   0 - 0x0
      11'h728: dout <= 8'b00000000; // 1832 :   0 - 0x0 -- Sprite 0xe5
      11'h729: dout <= 8'b00000000; // 1833 :   0 - 0x0
      11'h72A: dout <= 8'b00000000; // 1834 :   0 - 0x0
      11'h72B: dout <= 8'b00000000; // 1835 :   0 - 0x0
      11'h72C: dout <= 8'b00000000; // 1836 :   0 - 0x0
      11'h72D: dout <= 8'b00000000; // 1837 :   0 - 0x0
      11'h72E: dout <= 8'b00000000; // 1838 :   0 - 0x0
      11'h72F: dout <= 8'b00000000; // 1839 :   0 - 0x0
      11'h730: dout <= 8'b00000000; // 1840 :   0 - 0x0 -- Sprite 0xe6
      11'h731: dout <= 8'b00000000; // 1841 :   0 - 0x0
      11'h732: dout <= 8'b00000000; // 1842 :   0 - 0x0
      11'h733: dout <= 8'b00000000; // 1843 :   0 - 0x0
      11'h734: dout <= 8'b00000000; // 1844 :   0 - 0x0
      11'h735: dout <= 8'b00000000; // 1845 :   0 - 0x0
      11'h736: dout <= 8'b00000000; // 1846 :   0 - 0x0
      11'h737: dout <= 8'b00000000; // 1847 :   0 - 0x0
      11'h738: dout <= 8'b00000000; // 1848 :   0 - 0x0 -- Sprite 0xe7
      11'h739: dout <= 8'b00000000; // 1849 :   0 - 0x0
      11'h73A: dout <= 8'b00000000; // 1850 :   0 - 0x0
      11'h73B: dout <= 8'b00000000; // 1851 :   0 - 0x0
      11'h73C: dout <= 8'b00000000; // 1852 :   0 - 0x0
      11'h73D: dout <= 8'b00000000; // 1853 :   0 - 0x0
      11'h73E: dout <= 8'b00000000; // 1854 :   0 - 0x0
      11'h73F: dout <= 8'b00000000; // 1855 :   0 - 0x0
      11'h740: dout <= 8'b00000000; // 1856 :   0 - 0x0 -- Sprite 0xe8
      11'h741: dout <= 8'b00000000; // 1857 :   0 - 0x0
      11'h742: dout <= 8'b00000000; // 1858 :   0 - 0x0
      11'h743: dout <= 8'b00000000; // 1859 :   0 - 0x0
      11'h744: dout <= 8'b00000000; // 1860 :   0 - 0x0
      11'h745: dout <= 8'b00000000; // 1861 :   0 - 0x0
      11'h746: dout <= 8'b00000000; // 1862 :   0 - 0x0
      11'h747: dout <= 8'b00000000; // 1863 :   0 - 0x0
      11'h748: dout <= 8'b00000000; // 1864 :   0 - 0x0 -- Sprite 0xe9
      11'h749: dout <= 8'b00000000; // 1865 :   0 - 0x0
      11'h74A: dout <= 8'b00000000; // 1866 :   0 - 0x0
      11'h74B: dout <= 8'b00000000; // 1867 :   0 - 0x0
      11'h74C: dout <= 8'b00000000; // 1868 :   0 - 0x0
      11'h74D: dout <= 8'b00000000; // 1869 :   0 - 0x0
      11'h74E: dout <= 8'b00000000; // 1870 :   0 - 0x0
      11'h74F: dout <= 8'b00000000; // 1871 :   0 - 0x0
      11'h750: dout <= 8'b00000000; // 1872 :   0 - 0x0 -- Sprite 0xea
      11'h751: dout <= 8'b00000000; // 1873 :   0 - 0x0
      11'h752: dout <= 8'b00000000; // 1874 :   0 - 0x0
      11'h753: dout <= 8'b00000000; // 1875 :   0 - 0x0
      11'h754: dout <= 8'b00000000; // 1876 :   0 - 0x0
      11'h755: dout <= 8'b00000000; // 1877 :   0 - 0x0
      11'h756: dout <= 8'b00000000; // 1878 :   0 - 0x0
      11'h757: dout <= 8'b00000000; // 1879 :   0 - 0x0
      11'h758: dout <= 8'b00000000; // 1880 :   0 - 0x0 -- Sprite 0xeb
      11'h759: dout <= 8'b00000000; // 1881 :   0 - 0x0
      11'h75A: dout <= 8'b00000000; // 1882 :   0 - 0x0
      11'h75B: dout <= 8'b00000000; // 1883 :   0 - 0x0
      11'h75C: dout <= 8'b00000000; // 1884 :   0 - 0x0
      11'h75D: dout <= 8'b00000000; // 1885 :   0 - 0x0
      11'h75E: dout <= 8'b00000000; // 1886 :   0 - 0x0
      11'h75F: dout <= 8'b00000000; // 1887 :   0 - 0x0
      11'h760: dout <= 8'b00000000; // 1888 :   0 - 0x0 -- Sprite 0xec
      11'h761: dout <= 8'b00000000; // 1889 :   0 - 0x0
      11'h762: dout <= 8'b00000000; // 1890 :   0 - 0x0
      11'h763: dout <= 8'b00000000; // 1891 :   0 - 0x0
      11'h764: dout <= 8'b00000000; // 1892 :   0 - 0x0
      11'h765: dout <= 8'b00000000; // 1893 :   0 - 0x0
      11'h766: dout <= 8'b00000000; // 1894 :   0 - 0x0
      11'h767: dout <= 8'b00000000; // 1895 :   0 - 0x0
      11'h768: dout <= 8'b00000000; // 1896 :   0 - 0x0 -- Sprite 0xed
      11'h769: dout <= 8'b00000000; // 1897 :   0 - 0x0
      11'h76A: dout <= 8'b00000000; // 1898 :   0 - 0x0
      11'h76B: dout <= 8'b00000000; // 1899 :   0 - 0x0
      11'h76C: dout <= 8'b00000000; // 1900 :   0 - 0x0
      11'h76D: dout <= 8'b00000000; // 1901 :   0 - 0x0
      11'h76E: dout <= 8'b00000000; // 1902 :   0 - 0x0
      11'h76F: dout <= 8'b00000000; // 1903 :   0 - 0x0
      11'h770: dout <= 8'b00000000; // 1904 :   0 - 0x0 -- Sprite 0xee
      11'h771: dout <= 8'b00000000; // 1905 :   0 - 0x0
      11'h772: dout <= 8'b00000000; // 1906 :   0 - 0x0
      11'h773: dout <= 8'b00000000; // 1907 :   0 - 0x0
      11'h774: dout <= 8'b00000000; // 1908 :   0 - 0x0
      11'h775: dout <= 8'b00000000; // 1909 :   0 - 0x0
      11'h776: dout <= 8'b00000000; // 1910 :   0 - 0x0
      11'h777: dout <= 8'b00000000; // 1911 :   0 - 0x0
      11'h778: dout <= 8'b00000000; // 1912 :   0 - 0x0 -- Sprite 0xef
      11'h779: dout <= 8'b00000000; // 1913 :   0 - 0x0
      11'h77A: dout <= 8'b00000000; // 1914 :   0 - 0x0
      11'h77B: dout <= 8'b00000000; // 1915 :   0 - 0x0
      11'h77C: dout <= 8'b00000000; // 1916 :   0 - 0x0
      11'h77D: dout <= 8'b00000000; // 1917 :   0 - 0x0
      11'h77E: dout <= 8'b00000000; // 1918 :   0 - 0x0
      11'h77F: dout <= 8'b00000000; // 1919 :   0 - 0x0
      11'h780: dout <= 8'b00000000; // 1920 :   0 - 0x0 -- Sprite 0xf0
      11'h781: dout <= 8'b00000000; // 1921 :   0 - 0x0
      11'h782: dout <= 8'b00000000; // 1922 :   0 - 0x0
      11'h783: dout <= 8'b00000000; // 1923 :   0 - 0x0
      11'h784: dout <= 8'b00000000; // 1924 :   0 - 0x0
      11'h785: dout <= 8'b00000000; // 1925 :   0 - 0x0
      11'h786: dout <= 8'b00000000; // 1926 :   0 - 0x0
      11'h787: dout <= 8'b00000000; // 1927 :   0 - 0x0
      11'h788: dout <= 8'b00000000; // 1928 :   0 - 0x0 -- Sprite 0xf1
      11'h789: dout <= 8'b00000000; // 1929 :   0 - 0x0
      11'h78A: dout <= 8'b00000000; // 1930 :   0 - 0x0
      11'h78B: dout <= 8'b00000000; // 1931 :   0 - 0x0
      11'h78C: dout <= 8'b00000000; // 1932 :   0 - 0x0
      11'h78D: dout <= 8'b00000000; // 1933 :   0 - 0x0
      11'h78E: dout <= 8'b00000000; // 1934 :   0 - 0x0
      11'h78F: dout <= 8'b00000000; // 1935 :   0 - 0x0
      11'h790: dout <= 8'b00000000; // 1936 :   0 - 0x0 -- Sprite 0xf2
      11'h791: dout <= 8'b00000000; // 1937 :   0 - 0x0
      11'h792: dout <= 8'b00000000; // 1938 :   0 - 0x0
      11'h793: dout <= 8'b00000000; // 1939 :   0 - 0x0
      11'h794: dout <= 8'b00000000; // 1940 :   0 - 0x0
      11'h795: dout <= 8'b00000000; // 1941 :   0 - 0x0
      11'h796: dout <= 8'b00000000; // 1942 :   0 - 0x0
      11'h797: dout <= 8'b00000000; // 1943 :   0 - 0x0
      11'h798: dout <= 8'b00000000; // 1944 :   0 - 0x0 -- Sprite 0xf3
      11'h799: dout <= 8'b00000000; // 1945 :   0 - 0x0
      11'h79A: dout <= 8'b00000000; // 1946 :   0 - 0x0
      11'h79B: dout <= 8'b00000000; // 1947 :   0 - 0x0
      11'h79C: dout <= 8'b00000000; // 1948 :   0 - 0x0
      11'h79D: dout <= 8'b00000000; // 1949 :   0 - 0x0
      11'h79E: dout <= 8'b00000000; // 1950 :   0 - 0x0
      11'h79F: dout <= 8'b00000000; // 1951 :   0 - 0x0
      11'h7A0: dout <= 8'b00000000; // 1952 :   0 - 0x0 -- Sprite 0xf4
      11'h7A1: dout <= 8'b00000000; // 1953 :   0 - 0x0
      11'h7A2: dout <= 8'b00000000; // 1954 :   0 - 0x0
      11'h7A3: dout <= 8'b00000000; // 1955 :   0 - 0x0
      11'h7A4: dout <= 8'b00000000; // 1956 :   0 - 0x0
      11'h7A5: dout <= 8'b00000000; // 1957 :   0 - 0x0
      11'h7A6: dout <= 8'b00000000; // 1958 :   0 - 0x0
      11'h7A7: dout <= 8'b00000000; // 1959 :   0 - 0x0
      11'h7A8: dout <= 8'b00000000; // 1960 :   0 - 0x0 -- Sprite 0xf5
      11'h7A9: dout <= 8'b00000000; // 1961 :   0 - 0x0
      11'h7AA: dout <= 8'b00000000; // 1962 :   0 - 0x0
      11'h7AB: dout <= 8'b00000000; // 1963 :   0 - 0x0
      11'h7AC: dout <= 8'b00000000; // 1964 :   0 - 0x0
      11'h7AD: dout <= 8'b00000000; // 1965 :   0 - 0x0
      11'h7AE: dout <= 8'b00000000; // 1966 :   0 - 0x0
      11'h7AF: dout <= 8'b00000000; // 1967 :   0 - 0x0
      11'h7B0: dout <= 8'b00000000; // 1968 :   0 - 0x0 -- Sprite 0xf6
      11'h7B1: dout <= 8'b00000000; // 1969 :   0 - 0x0
      11'h7B2: dout <= 8'b00000000; // 1970 :   0 - 0x0
      11'h7B3: dout <= 8'b00000000; // 1971 :   0 - 0x0
      11'h7B4: dout <= 8'b00000000; // 1972 :   0 - 0x0
      11'h7B5: dout <= 8'b00000000; // 1973 :   0 - 0x0
      11'h7B6: dout <= 8'b00000000; // 1974 :   0 - 0x0
      11'h7B7: dout <= 8'b00000000; // 1975 :   0 - 0x0
      11'h7B8: dout <= 8'b00000000; // 1976 :   0 - 0x0 -- Sprite 0xf7
      11'h7B9: dout <= 8'b00000000; // 1977 :   0 - 0x0
      11'h7BA: dout <= 8'b00000000; // 1978 :   0 - 0x0
      11'h7BB: dout <= 8'b00000000; // 1979 :   0 - 0x0
      11'h7BC: dout <= 8'b00000000; // 1980 :   0 - 0x0
      11'h7BD: dout <= 8'b00000000; // 1981 :   0 - 0x0
      11'h7BE: dout <= 8'b00000000; // 1982 :   0 - 0x0
      11'h7BF: dout <= 8'b00000000; // 1983 :   0 - 0x0
      11'h7C0: dout <= 8'b00000000; // 1984 :   0 - 0x0 -- Sprite 0xf8
      11'h7C1: dout <= 8'b00000000; // 1985 :   0 - 0x0
      11'h7C2: dout <= 8'b00000000; // 1986 :   0 - 0x0
      11'h7C3: dout <= 8'b00000000; // 1987 :   0 - 0x0
      11'h7C4: dout <= 8'b00000000; // 1988 :   0 - 0x0
      11'h7C5: dout <= 8'b00000000; // 1989 :   0 - 0x0
      11'h7C6: dout <= 8'b00000000; // 1990 :   0 - 0x0
      11'h7C7: dout <= 8'b00000000; // 1991 :   0 - 0x0
      11'h7C8: dout <= 8'b00000000; // 1992 :   0 - 0x0 -- Sprite 0xf9
      11'h7C9: dout <= 8'b00000000; // 1993 :   0 - 0x0
      11'h7CA: dout <= 8'b00000000; // 1994 :   0 - 0x0
      11'h7CB: dout <= 8'b00000000; // 1995 :   0 - 0x0
      11'h7CC: dout <= 8'b00000000; // 1996 :   0 - 0x0
      11'h7CD: dout <= 8'b00000000; // 1997 :   0 - 0x0
      11'h7CE: dout <= 8'b00000000; // 1998 :   0 - 0x0
      11'h7CF: dout <= 8'b00000000; // 1999 :   0 - 0x0
      11'h7D0: dout <= 8'b00000000; // 2000 :   0 - 0x0 -- Sprite 0xfa
      11'h7D1: dout <= 8'b00000000; // 2001 :   0 - 0x0
      11'h7D2: dout <= 8'b00000000; // 2002 :   0 - 0x0
      11'h7D3: dout <= 8'b00000000; // 2003 :   0 - 0x0
      11'h7D4: dout <= 8'b00000000; // 2004 :   0 - 0x0
      11'h7D5: dout <= 8'b00000000; // 2005 :   0 - 0x0
      11'h7D6: dout <= 8'b00000000; // 2006 :   0 - 0x0
      11'h7D7: dout <= 8'b00000000; // 2007 :   0 - 0x0
      11'h7D8: dout <= 8'b00000000; // 2008 :   0 - 0x0 -- Sprite 0xfb
      11'h7D9: dout <= 8'b00000000; // 2009 :   0 - 0x0
      11'h7DA: dout <= 8'b00000000; // 2010 :   0 - 0x0
      11'h7DB: dout <= 8'b00000000; // 2011 :   0 - 0x0
      11'h7DC: dout <= 8'b00000000; // 2012 :   0 - 0x0
      11'h7DD: dout <= 8'b00000000; // 2013 :   0 - 0x0
      11'h7DE: dout <= 8'b00000000; // 2014 :   0 - 0x0
      11'h7DF: dout <= 8'b00000000; // 2015 :   0 - 0x0
      11'h7E0: dout <= 8'b00000000; // 2016 :   0 - 0x0 -- Sprite 0xfc
      11'h7E1: dout <= 8'b00000000; // 2017 :   0 - 0x0
      11'h7E2: dout <= 8'b10001110; // 2018 : 142 - 0x8e
      11'h7E3: dout <= 8'b10001010; // 2019 : 138 - 0x8a
      11'h7E4: dout <= 8'b10001010; // 2020 : 138 - 0x8a
      11'h7E5: dout <= 8'b10001010; // 2021 : 138 - 0x8a
      11'h7E6: dout <= 8'b10001010; // 2022 : 138 - 0x8a
      11'h7E7: dout <= 8'b11101110; // 2023 : 238 - 0xee
      11'h7E8: dout <= 8'b00000000; // 2024 :   0 - 0x0 -- Sprite 0xfd
      11'h7E9: dout <= 8'b00000000; // 2025 :   0 - 0x0
      11'h7EA: dout <= 8'b01001100; // 2026 :  76 - 0x4c
      11'h7EB: dout <= 8'b10101010; // 2027 : 170 - 0xaa
      11'h7EC: dout <= 8'b10101010; // 2028 : 170 - 0xaa
      11'h7ED: dout <= 8'b11101010; // 2029 : 234 - 0xea
      11'h7EE: dout <= 8'b10101010; // 2030 : 170 - 0xaa
      11'h7EF: dout <= 8'b10101100; // 2031 : 172 - 0xac
      11'h7F0: dout <= 8'b00000000; // 2032 :   0 - 0x0 -- Sprite 0xfe
      11'h7F1: dout <= 8'b00000000; // 2033 :   0 - 0x0
      11'h7F2: dout <= 8'b11101100; // 2034 : 236 - 0xec
      11'h7F3: dout <= 8'b01001010; // 2035 :  74 - 0x4a
      11'h7F4: dout <= 8'b01001010; // 2036 :  74 - 0x4a
      11'h7F5: dout <= 8'b01001010; // 2037 :  74 - 0x4a
      11'h7F6: dout <= 8'b01001010; // 2038 :  74 - 0x4a
      11'h7F7: dout <= 8'b11101010; // 2039 : 234 - 0xea
      11'h7F8: dout <= 8'b00000000; // 2040 :   0 - 0x0 -- Sprite 0xff
      11'h7F9: dout <= 8'b00000000; // 2041 :   0 - 0x0
      11'h7FA: dout <= 8'b01100000; // 2042 :  96 - 0x60
      11'h7FB: dout <= 8'b10001000; // 2043 : 136 - 0x88
      11'h7FC: dout <= 8'b10100000; // 2044 : 160 - 0xa0
      11'h7FD: dout <= 8'b10100000; // 2045 : 160 - 0xa0
      11'h7FE: dout <= 8'b10101000; // 2046 : 168 - 0xa8
      11'h7FF: dout <= 8'b01000000; // 2047 :  64 - 0x40
    endcase
  end

endmodule
