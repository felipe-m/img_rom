//- Autcmatically generated verilog ROM from a NES memory file----
//-   PATTERN TABLE
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


//-  Original memory dump file name: smario_traspas_patron.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_PTABLE_SMARIO_TRASPAS
  (
     //input     clk,   // clock
     input      [13-1:0] addr,  //8192 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Pattern Table 0---------
      13'h0: dout  = 8'b00000011; //    0 :   3 - 0x3 -- Sprite 0x0
      13'h1: dout  = 8'b00001111; //    1 :  15 - 0xf
      13'h2: dout  = 8'b00011111; //    2 :  31 - 0x1f
      13'h3: dout  = 8'b00011111; //    3 :  31 - 0x1f
      13'h4: dout  = 8'b00011100; //    4 :  28 - 0x1c
      13'h5: dout  = 8'b00100100; //    5 :  36 - 0x24
      13'h6: dout  = 8'b00100110; //    6 :  38 - 0x26
      13'h7: dout  = 8'b01100110; //    7 : 102 - 0x66
      13'h8: dout  = 8'b00000000; //    8 :   0 - 0x0
      13'h9: dout  = 8'b00000000; //    9 :   0 - 0x0
      13'hA: dout  = 8'b00000000; //   10 :   0 - 0x0
      13'hB: dout  = 8'b00000000; //   11 :   0 - 0x0
      13'hC: dout  = 8'b00011111; //   12 :  31 - 0x1f
      13'hD: dout  = 8'b00111111; //   13 :  63 - 0x3f
      13'hE: dout  = 8'b00111111; //   14 :  63 - 0x3f
      13'hF: dout  = 8'b01111111; //   15 : 127 - 0x7f
      13'h10: dout  = 8'b11100000; //   16 : 224 - 0xe0 -- Sprite 0x1
      13'h11: dout  = 8'b11000000; //   17 : 192 - 0xc0
      13'h12: dout  = 8'b10000000; //   18 : 128 - 0x80
      13'h13: dout  = 8'b11111100; //   19 : 252 - 0xfc
      13'h14: dout  = 8'b10000000; //   20 : 128 - 0x80
      13'h15: dout  = 8'b11000000; //   21 : 192 - 0xc0
      13'h16: dout  = 8'b00000000; //   22 :   0 - 0x0
      13'h17: dout  = 8'b00100000; //   23 :  32 - 0x20
      13'h18: dout  = 8'b00000000; //   24 :   0 - 0x0
      13'h19: dout  = 8'b00100000; //   25 :  32 - 0x20
      13'h1A: dout  = 8'b01100000; //   26 :  96 - 0x60
      13'h1B: dout  = 8'b00000000; //   27 :   0 - 0x0
      13'h1C: dout  = 8'b11110000; //   28 : 240 - 0xf0
      13'h1D: dout  = 8'b11111100; //   29 : 252 - 0xfc
      13'h1E: dout  = 8'b11111110; //   30 : 254 - 0xfe
      13'h1F: dout  = 8'b11111110; //   31 : 254 - 0xfe
      13'h20: dout  = 8'b01100000; //   32 :  96 - 0x60 -- Sprite 0x2
      13'h21: dout  = 8'b01110000; //   33 : 112 - 0x70
      13'h22: dout  = 8'b00011000; //   34 :  24 - 0x18
      13'h23: dout  = 8'b00000111; //   35 :   7 - 0x7
      13'h24: dout  = 8'b00001111; //   36 :  15 - 0xf
      13'h25: dout  = 8'b00011111; //   37 :  31 - 0x1f
      13'h26: dout  = 8'b00111111; //   38 :  63 - 0x3f
      13'h27: dout  = 8'b01111111; //   39 : 127 - 0x7f
      13'h28: dout  = 8'b01111111; //   40 : 127 - 0x7f
      13'h29: dout  = 8'b01111111; //   41 : 127 - 0x7f
      13'h2A: dout  = 8'b00011111; //   42 :  31 - 0x1f
      13'h2B: dout  = 8'b00000111; //   43 :   7 - 0x7
      13'h2C: dout  = 8'b00000000; //   44 :   0 - 0x0
      13'h2D: dout  = 8'b00011110; //   45 :  30 - 0x1e
      13'h2E: dout  = 8'b00111111; //   46 :  63 - 0x3f
      13'h2F: dout  = 8'b01111111; //   47 : 127 - 0x7f
      13'h30: dout  = 8'b11111100; //   48 : 252 - 0xfc -- Sprite 0x3
      13'h31: dout  = 8'b01111100; //   49 : 124 - 0x7c
      13'h32: dout  = 8'b00000000; //   50 :   0 - 0x0
      13'h33: dout  = 8'b00000000; //   51 :   0 - 0x0
      13'h34: dout  = 8'b11100000; //   52 : 224 - 0xe0
      13'h35: dout  = 8'b11110000; //   53 : 240 - 0xf0
      13'h36: dout  = 8'b11111000; //   54 : 248 - 0xf8
      13'h37: dout  = 8'b11111000; //   55 : 248 - 0xf8
      13'h38: dout  = 8'b11111100; //   56 : 252 - 0xfc
      13'h39: dout  = 8'b11111100; //   57 : 252 - 0xfc
      13'h3A: dout  = 8'b11111000; //   58 : 248 - 0xf8
      13'h3B: dout  = 8'b11000000; //   59 : 192 - 0xc0
      13'h3C: dout  = 8'b11000010; //   60 : 194 - 0xc2
      13'h3D: dout  = 8'b01100111; //   61 : 103 - 0x67
      13'h3E: dout  = 8'b00101111; //   62 :  47 - 0x2f
      13'h3F: dout  = 8'b00110111; //   63 :  55 - 0x37
      13'h40: dout  = 8'b01111111; //   64 : 127 - 0x7f -- Sprite 0x4
      13'h41: dout  = 8'b01111111; //   65 : 127 - 0x7f
      13'h42: dout  = 8'b11111111; //   66 : 255 - 0xff
      13'h43: dout  = 8'b11111111; //   67 : 255 - 0xff
      13'h44: dout  = 8'b00000111; //   68 :   7 - 0x7
      13'h45: dout  = 8'b00000111; //   69 :   7 - 0x7
      13'h46: dout  = 8'b00001111; //   70 :  15 - 0xf
      13'h47: dout  = 8'b00001111; //   71 :  15 - 0xf
      13'h48: dout  = 8'b01111111; //   72 : 127 - 0x7f
      13'h49: dout  = 8'b01111110; //   73 : 126 - 0x7e
      13'h4A: dout  = 8'b11111100; //   74 : 252 - 0xfc
      13'h4B: dout  = 8'b11110000; //   75 : 240 - 0xf0
      13'h4C: dout  = 8'b11111000; //   76 : 248 - 0xf8
      13'h4D: dout  = 8'b11111000; //   77 : 248 - 0xf8
      13'h4E: dout  = 8'b11110000; //   78 : 240 - 0xf0
      13'h4F: dout  = 8'b01110000; //   79 : 112 - 0x70
      13'h50: dout  = 8'b11111101; //   80 : 253 - 0xfd -- Sprite 0x5
      13'h51: dout  = 8'b11111110; //   81 : 254 - 0xfe
      13'h52: dout  = 8'b10110100; //   82 : 180 - 0xb4
      13'h53: dout  = 8'b11111000; //   83 : 248 - 0xf8
      13'h54: dout  = 8'b11111000; //   84 : 248 - 0xf8
      13'h55: dout  = 8'b11111001; //   85 : 249 - 0xf9
      13'h56: dout  = 8'b11111011; //   86 : 251 - 0xfb
      13'h57: dout  = 8'b11111111; //   87 : 255 - 0xff
      13'h58: dout  = 8'b00110111; //   88 :  55 - 0x37
      13'h59: dout  = 8'b00110110; //   89 :  54 - 0x36
      13'h5A: dout  = 8'b01011100; //   90 :  92 - 0x5c
      13'h5B: dout  = 8'b00000000; //   91 :   0 - 0x0
      13'h5C: dout  = 8'b00000000; //   92 :   0 - 0x0
      13'h5D: dout  = 8'b00000001; //   93 :   1 - 0x1
      13'h5E: dout  = 8'b00000011; //   94 :   3 - 0x3
      13'h5F: dout  = 8'b00011111; //   95 :  31 - 0x1f
      13'h60: dout  = 8'b00011111; //   96 :  31 - 0x1f -- Sprite 0x6
      13'h61: dout  = 8'b00111111; //   97 :  63 - 0x3f
      13'h62: dout  = 8'b11111111; //   98 : 255 - 0xff
      13'h63: dout  = 8'b11111111; //   99 : 255 - 0xff
      13'h64: dout  = 8'b11111100; //  100 : 252 - 0xfc
      13'h65: dout  = 8'b01110000; //  101 : 112 - 0x70
      13'h66: dout  = 8'b01110000; //  102 : 112 - 0x70
      13'h67: dout  = 8'b00111000; //  103 :  56 - 0x38
      13'h68: dout  = 8'b00001000; //  104 :   8 - 0x8
      13'h69: dout  = 8'b00100100; //  105 :  36 - 0x24
      13'h6A: dout  = 8'b11100011; //  106 : 227 - 0xe3
      13'h6B: dout  = 8'b11110000; //  107 : 240 - 0xf0
      13'h6C: dout  = 8'b11111000; //  108 : 248 - 0xf8
      13'h6D: dout  = 8'b01110000; //  109 : 112 - 0x70
      13'h6E: dout  = 8'b01110000; //  110 : 112 - 0x70
      13'h6F: dout  = 8'b00111000; //  111 :  56 - 0x38
      13'h70: dout  = 8'b11111111; //  112 : 255 - 0xff -- Sprite 0x7
      13'h71: dout  = 8'b11111111; //  113 : 255 - 0xff
      13'h72: dout  = 8'b11111111; //  114 : 255 - 0xff
      13'h73: dout  = 8'b00011111; //  115 :  31 - 0x1f
      13'h74: dout  = 8'b00000000; //  116 :   0 - 0x0
      13'h75: dout  = 8'b00000000; //  117 :   0 - 0x0
      13'h76: dout  = 8'b00000000; //  118 :   0 - 0x0
      13'h77: dout  = 8'b00000000; //  119 :   0 - 0x0
      13'h78: dout  = 8'b00011111; //  120 :  31 - 0x1f
      13'h79: dout  = 8'b00011111; //  121 :  31 - 0x1f
      13'h7A: dout  = 8'b00011111; //  122 :  31 - 0x1f
      13'h7B: dout  = 8'b00011111; //  123 :  31 - 0x1f
      13'h7C: dout  = 8'b00000000; //  124 :   0 - 0x0
      13'h7D: dout  = 8'b00000000; //  125 :   0 - 0x0
      13'h7E: dout  = 8'b00000000; //  126 :   0 - 0x0
      13'h7F: dout  = 8'b00000000; //  127 :   0 - 0x0
      13'h80: dout  = 8'b00000000; //  128 :   0 - 0x0 -- Sprite 0x8
      13'h81: dout  = 8'b00000000; //  129 :   0 - 0x0
      13'h82: dout  = 8'b00000001; //  130 :   1 - 0x1
      13'h83: dout  = 8'b00000111; //  131 :   7 - 0x7
      13'h84: dout  = 8'b00001111; //  132 :  15 - 0xf
      13'h85: dout  = 8'b00001111; //  133 :  15 - 0xf
      13'h86: dout  = 8'b00001110; //  134 :  14 - 0xe
      13'h87: dout  = 8'b00010010; //  135 :  18 - 0x12
      13'h88: dout  = 8'b00000000; //  136 :   0 - 0x0
      13'h89: dout  = 8'b00000000; //  137 :   0 - 0x0
      13'h8A: dout  = 8'b00000000; //  138 :   0 - 0x0
      13'h8B: dout  = 8'b00000000; //  139 :   0 - 0x0
      13'h8C: dout  = 8'b00000000; //  140 :   0 - 0x0
      13'h8D: dout  = 8'b00000000; //  141 :   0 - 0x0
      13'h8E: dout  = 8'b00001111; //  142 :  15 - 0xf
      13'h8F: dout  = 8'b00011111; //  143 :  31 - 0x1f
      13'h90: dout  = 8'b00000000; //  144 :   0 - 0x0 -- Sprite 0x9
      13'h91: dout  = 8'b00000000; //  145 :   0 - 0x0
      13'h92: dout  = 8'b11110000; //  146 : 240 - 0xf0
      13'h93: dout  = 8'b11100000; //  147 : 224 - 0xe0
      13'h94: dout  = 8'b11000000; //  148 : 192 - 0xc0
      13'h95: dout  = 8'b11111110; //  149 : 254 - 0xfe
      13'h96: dout  = 8'b01000000; //  150 :  64 - 0x40
      13'h97: dout  = 8'b01100000; //  151 :  96 - 0x60
      13'h98: dout  = 8'b00000000; //  152 :   0 - 0x0
      13'h99: dout  = 8'b00000000; //  153 :   0 - 0x0
      13'h9A: dout  = 8'b00000000; //  154 :   0 - 0x0
      13'h9B: dout  = 8'b00010000; //  155 :  16 - 0x10
      13'h9C: dout  = 8'b00110000; //  156 :  48 - 0x30
      13'h9D: dout  = 8'b00000000; //  157 :   0 - 0x0
      13'h9E: dout  = 8'b11111000; //  158 : 248 - 0xf8
      13'h9F: dout  = 8'b11111110; //  159 : 254 - 0xfe
      13'hA0: dout  = 8'b00010011; //  160 :  19 - 0x13 -- Sprite 0xa
      13'hA1: dout  = 8'b00110011; //  161 :  51 - 0x33
      13'hA2: dout  = 8'b00110000; //  162 :  48 - 0x30
      13'hA3: dout  = 8'b00011000; //  163 :  24 - 0x18
      13'hA4: dout  = 8'b00000100; //  164 :   4 - 0x4
      13'hA5: dout  = 8'b00001111; //  165 :  15 - 0xf
      13'hA6: dout  = 8'b00011111; //  166 :  31 - 0x1f
      13'hA7: dout  = 8'b00011111; //  167 :  31 - 0x1f
      13'hA8: dout  = 8'b00011111; //  168 :  31 - 0x1f
      13'hA9: dout  = 8'b00111111; //  169 :  63 - 0x3f
      13'hAA: dout  = 8'b00111111; //  170 :  63 - 0x3f
      13'hAB: dout  = 8'b00011111; //  171 :  31 - 0x1f
      13'hAC: dout  = 8'b00000111; //  172 :   7 - 0x7
      13'hAD: dout  = 8'b00001000; //  173 :   8 - 0x8
      13'hAE: dout  = 8'b00010111; //  174 :  23 - 0x17
      13'hAF: dout  = 8'b00010111; //  175 :  23 - 0x17
      13'hB0: dout  = 8'b00000000; //  176 :   0 - 0x0 -- Sprite 0xb
      13'hB1: dout  = 8'b00010000; //  177 :  16 - 0x10
      13'hB2: dout  = 8'b01111110; //  178 : 126 - 0x7e
      13'hB3: dout  = 8'b00111110; //  179 :  62 - 0x3e
      13'hB4: dout  = 8'b00000000; //  180 :   0 - 0x0
      13'hB5: dout  = 8'b00000000; //  181 :   0 - 0x0
      13'hB6: dout  = 8'b11000000; //  182 : 192 - 0xc0
      13'hB7: dout  = 8'b11100000; //  183 : 224 - 0xe0
      13'hB8: dout  = 8'b11111111; //  184 : 255 - 0xff
      13'hB9: dout  = 8'b11111111; //  185 : 255 - 0xff
      13'hBA: dout  = 8'b11111110; //  186 : 254 - 0xfe
      13'hBB: dout  = 8'b11111110; //  187 : 254 - 0xfe
      13'hBC: dout  = 8'b11111100; //  188 : 252 - 0xfc
      13'hBD: dout  = 8'b11100000; //  189 : 224 - 0xe0
      13'hBE: dout  = 8'b01000000; //  190 :  64 - 0x40
      13'hBF: dout  = 8'b10100000; //  191 : 160 - 0xa0
      13'hC0: dout  = 8'b00111111; //  192 :  63 - 0x3f -- Sprite 0xc
      13'hC1: dout  = 8'b00111111; //  193 :  63 - 0x3f
      13'hC2: dout  = 8'b00111111; //  194 :  63 - 0x3f
      13'hC3: dout  = 8'b00011111; //  195 :  31 - 0x1f
      13'hC4: dout  = 8'b00011111; //  196 :  31 - 0x1f
      13'hC5: dout  = 8'b00011111; //  197 :  31 - 0x1f
      13'hC6: dout  = 8'b00011111; //  198 :  31 - 0x1f
      13'hC7: dout  = 8'b00011111; //  199 :  31 - 0x1f
      13'hC8: dout  = 8'b00110111; //  200 :  55 - 0x37
      13'hC9: dout  = 8'b00100111; //  201 :  39 - 0x27
      13'hCA: dout  = 8'b00100011; //  202 :  35 - 0x23
      13'hCB: dout  = 8'b00000011; //  203 :   3 - 0x3
      13'hCC: dout  = 8'b00000001; //  204 :   1 - 0x1
      13'hCD: dout  = 8'b00000000; //  205 :   0 - 0x0
      13'hCE: dout  = 8'b00000000; //  206 :   0 - 0x0
      13'hCF: dout  = 8'b00000000; //  207 :   0 - 0x0
      13'hD0: dout  = 8'b11110000; //  208 : 240 - 0xf0 -- Sprite 0xd
      13'hD1: dout  = 8'b11110000; //  209 : 240 - 0xf0
      13'hD2: dout  = 8'b11110000; //  210 : 240 - 0xf0
      13'hD3: dout  = 8'b11111000; //  211 : 248 - 0xf8
      13'hD4: dout  = 8'b11111000; //  212 : 248 - 0xf8
      13'hD5: dout  = 8'b11111000; //  213 : 248 - 0xf8
      13'hD6: dout  = 8'b11111000; //  214 : 248 - 0xf8
      13'hD7: dout  = 8'b11111000; //  215 : 248 - 0xf8
      13'hD8: dout  = 8'b11001100; //  216 : 204 - 0xcc
      13'hD9: dout  = 8'b11111111; //  217 : 255 - 0xff
      13'hDA: dout  = 8'b11111111; //  218 : 255 - 0xff
      13'hDB: dout  = 8'b11111111; //  219 : 255 - 0xff
      13'hDC: dout  = 8'b11111111; //  220 : 255 - 0xff
      13'hDD: dout  = 8'b01110000; //  221 : 112 - 0x70
      13'hDE: dout  = 8'b00000000; //  222 :   0 - 0x0
      13'hDF: dout  = 8'b00001000; //  223 :   8 - 0x8
      13'hE0: dout  = 8'b11111111; //  224 : 255 - 0xff -- Sprite 0xe
      13'hE1: dout  = 8'b11111111; //  225 : 255 - 0xff
      13'hE2: dout  = 8'b11111111; //  226 : 255 - 0xff
      13'hE3: dout  = 8'b11111110; //  227 : 254 - 0xfe
      13'hE4: dout  = 8'b11110000; //  228 : 240 - 0xf0
      13'hE5: dout  = 8'b11000000; //  229 : 192 - 0xc0
      13'hE6: dout  = 8'b10000000; //  230 : 128 - 0x80
      13'hE7: dout  = 8'b00000000; //  231 :   0 - 0x0
      13'hE8: dout  = 8'b11110000; //  232 : 240 - 0xf0
      13'hE9: dout  = 8'b11110000; //  233 : 240 - 0xf0
      13'hEA: dout  = 8'b11110000; //  234 : 240 - 0xf0
      13'hEB: dout  = 8'b11110000; //  235 : 240 - 0xf0
      13'hEC: dout  = 8'b11110000; //  236 : 240 - 0xf0
      13'hED: dout  = 8'b11000000; //  237 : 192 - 0xc0
      13'hEE: dout  = 8'b10000000; //  238 : 128 - 0x80
      13'hEF: dout  = 8'b00000000; //  239 :   0 - 0x0
      13'hF0: dout  = 8'b11111100; //  240 : 252 - 0xfc -- Sprite 0xf
      13'hF1: dout  = 8'b11111100; //  241 : 252 - 0xfc
      13'hF2: dout  = 8'b11111000; //  242 : 248 - 0xf8
      13'hF3: dout  = 8'b01111000; //  243 : 120 - 0x78
      13'hF4: dout  = 8'b01111000; //  244 : 120 - 0x78
      13'hF5: dout  = 8'b01111000; //  245 : 120 - 0x78
      13'hF6: dout  = 8'b01111110; //  246 : 126 - 0x7e
      13'hF7: dout  = 8'b01111110; //  247 : 126 - 0x7e
      13'hF8: dout  = 8'b00010000; //  248 :  16 - 0x10
      13'hF9: dout  = 8'b01100000; //  249 :  96 - 0x60
      13'hFA: dout  = 8'b10000000; //  250 : 128 - 0x80
      13'hFB: dout  = 8'b00000000; //  251 :   0 - 0x0
      13'hFC: dout  = 8'b01111000; //  252 : 120 - 0x78
      13'hFD: dout  = 8'b01111000; //  253 : 120 - 0x78
      13'hFE: dout  = 8'b01111110; //  254 : 126 - 0x7e
      13'hFF: dout  = 8'b01111110; //  255 : 126 - 0x7e
      13'h100: dout  = 8'b00000000; //  256 :   0 - 0x0 -- Sprite 0x10
      13'h101: dout  = 8'b00000011; //  257 :   3 - 0x3
      13'h102: dout  = 8'b00001111; //  258 :  15 - 0xf
      13'h103: dout  = 8'b00011111; //  259 :  31 - 0x1f
      13'h104: dout  = 8'b00011111; //  260 :  31 - 0x1f
      13'h105: dout  = 8'b00011100; //  261 :  28 - 0x1c
      13'h106: dout  = 8'b00100100; //  262 :  36 - 0x24
      13'h107: dout  = 8'b00100110; //  263 :  38 - 0x26
      13'h108: dout  = 8'b00000000; //  264 :   0 - 0x0
      13'h109: dout  = 8'b00000000; //  265 :   0 - 0x0
      13'h10A: dout  = 8'b00000000; //  266 :   0 - 0x0
      13'h10B: dout  = 8'b00000000; //  267 :   0 - 0x0
      13'h10C: dout  = 8'b00000000; //  268 :   0 - 0x0
      13'h10D: dout  = 8'b00011111; //  269 :  31 - 0x1f
      13'h10E: dout  = 8'b00111111; //  270 :  63 - 0x3f
      13'h10F: dout  = 8'b00111111; //  271 :  63 - 0x3f
      13'h110: dout  = 8'b00000000; //  272 :   0 - 0x0 -- Sprite 0x11
      13'h111: dout  = 8'b11100000; //  273 : 224 - 0xe0
      13'h112: dout  = 8'b11000000; //  274 : 192 - 0xc0
      13'h113: dout  = 8'b10000000; //  275 : 128 - 0x80
      13'h114: dout  = 8'b11111100; //  276 : 252 - 0xfc
      13'h115: dout  = 8'b10000000; //  277 : 128 - 0x80
      13'h116: dout  = 8'b11000000; //  278 : 192 - 0xc0
      13'h117: dout  = 8'b00000000; //  279 :   0 - 0x0
      13'h118: dout  = 8'b00000000; //  280 :   0 - 0x0
      13'h119: dout  = 8'b00000000; //  281 :   0 - 0x0
      13'h11A: dout  = 8'b00100000; //  282 :  32 - 0x20
      13'h11B: dout  = 8'b01100000; //  283 :  96 - 0x60
      13'h11C: dout  = 8'b00000000; //  284 :   0 - 0x0
      13'h11D: dout  = 8'b11110000; //  285 : 240 - 0xf0
      13'h11E: dout  = 8'b11111100; //  286 : 252 - 0xfc
      13'h11F: dout  = 8'b11111110; //  287 : 254 - 0xfe
      13'h120: dout  = 8'b01100110; //  288 : 102 - 0x66 -- Sprite 0x12
      13'h121: dout  = 8'b01100000; //  289 :  96 - 0x60
      13'h122: dout  = 8'b00110000; //  290 :  48 - 0x30
      13'h123: dout  = 8'b00011000; //  291 :  24 - 0x18
      13'h124: dout  = 8'b00001111; //  292 :  15 - 0xf
      13'h125: dout  = 8'b00011111; //  293 :  31 - 0x1f
      13'h126: dout  = 8'b00111111; //  294 :  63 - 0x3f
      13'h127: dout  = 8'b00111111; //  295 :  63 - 0x3f
      13'h128: dout  = 8'b01111111; //  296 : 127 - 0x7f
      13'h129: dout  = 8'b01111111; //  297 : 127 - 0x7f
      13'h12A: dout  = 8'b00111111; //  298 :  63 - 0x3f
      13'h12B: dout  = 8'b00011111; //  299 :  31 - 0x1f
      13'h12C: dout  = 8'b00000000; //  300 :   0 - 0x0
      13'h12D: dout  = 8'b00010110; //  301 :  22 - 0x16
      13'h12E: dout  = 8'b00101111; //  302 :  47 - 0x2f
      13'h12F: dout  = 8'b00101111; //  303 :  47 - 0x2f
      13'h130: dout  = 8'b00100000; //  304 :  32 - 0x20 -- Sprite 0x13
      13'h131: dout  = 8'b11111100; //  305 : 252 - 0xfc
      13'h132: dout  = 8'b01111100; //  306 : 124 - 0x7c
      13'h133: dout  = 8'b00000000; //  307 :   0 - 0x0
      13'h134: dout  = 8'b00000000; //  308 :   0 - 0x0
      13'h135: dout  = 8'b11100000; //  309 : 224 - 0xe0
      13'h136: dout  = 8'b11100000; //  310 : 224 - 0xe0
      13'h137: dout  = 8'b11110000; //  311 : 240 - 0xf0
      13'h138: dout  = 8'b11111110; //  312 : 254 - 0xfe
      13'h139: dout  = 8'b11111100; //  313 : 252 - 0xfc
      13'h13A: dout  = 8'b11111100; //  314 : 252 - 0xfc
      13'h13B: dout  = 8'b11111000; //  315 : 248 - 0xf8
      13'h13C: dout  = 8'b11000000; //  316 : 192 - 0xc0
      13'h13D: dout  = 8'b01100000; //  317 :  96 - 0x60
      13'h13E: dout  = 8'b00100000; //  318 :  32 - 0x20
      13'h13F: dout  = 8'b00110000; //  319 :  48 - 0x30
      13'h140: dout  = 8'b00111111; //  320 :  63 - 0x3f -- Sprite 0x14
      13'h141: dout  = 8'b00111111; //  321 :  63 - 0x3f
      13'h142: dout  = 8'b00111111; //  322 :  63 - 0x3f
      13'h143: dout  = 8'b00111111; //  323 :  63 - 0x3f
      13'h144: dout  = 8'b00111111; //  324 :  63 - 0x3f
      13'h145: dout  = 8'b00111111; //  325 :  63 - 0x3f
      13'h146: dout  = 8'b00111111; //  326 :  63 - 0x3f
      13'h147: dout  = 8'b00011111; //  327 :  31 - 0x1f
      13'h148: dout  = 8'b00101111; //  328 :  47 - 0x2f
      13'h149: dout  = 8'b00101111; //  329 :  47 - 0x2f
      13'h14A: dout  = 8'b00101111; //  330 :  47 - 0x2f
      13'h14B: dout  = 8'b00001111; //  331 :  15 - 0xf
      13'h14C: dout  = 8'b00000111; //  332 :   7 - 0x7
      13'h14D: dout  = 8'b00000011; //  333 :   3 - 0x3
      13'h14E: dout  = 8'b00000000; //  334 :   0 - 0x0
      13'h14F: dout  = 8'b00000000; //  335 :   0 - 0x0
      13'h150: dout  = 8'b11110000; //  336 : 240 - 0xf0 -- Sprite 0x15
      13'h151: dout  = 8'b10010000; //  337 : 144 - 0x90
      13'h152: dout  = 8'b00000000; //  338 :   0 - 0x0
      13'h153: dout  = 8'b00001000; //  339 :   8 - 0x8
      13'h154: dout  = 8'b00001100; //  340 :  12 - 0xc
      13'h155: dout  = 8'b00011100; //  341 :  28 - 0x1c
      13'h156: dout  = 8'b11111100; //  342 : 252 - 0xfc
      13'h157: dout  = 8'b11111000; //  343 : 248 - 0xf8
      13'h158: dout  = 8'b00010000; //  344 :  16 - 0x10
      13'h159: dout  = 8'b11110000; //  345 : 240 - 0xf0
      13'h15A: dout  = 8'b11110000; //  346 : 240 - 0xf0
      13'h15B: dout  = 8'b11110000; //  347 : 240 - 0xf0
      13'h15C: dout  = 8'b11110000; //  348 : 240 - 0xf0
      13'h15D: dout  = 8'b11100000; //  349 : 224 - 0xe0
      13'h15E: dout  = 8'b11000000; //  350 : 192 - 0xc0
      13'h15F: dout  = 8'b11100000; //  351 : 224 - 0xe0
      13'h160: dout  = 8'b00001111; //  352 :  15 - 0xf -- Sprite 0x16
      13'h161: dout  = 8'b00001111; //  353 :  15 - 0xf
      13'h162: dout  = 8'b00000111; //  354 :   7 - 0x7
      13'h163: dout  = 8'b00000111; //  355 :   7 - 0x7
      13'h164: dout  = 8'b00000111; //  356 :   7 - 0x7
      13'h165: dout  = 8'b00001111; //  357 :  15 - 0xf
      13'h166: dout  = 8'b00001111; //  358 :  15 - 0xf
      13'h167: dout  = 8'b00000011; //  359 :   3 - 0x3
      13'h168: dout  = 8'b00000001; //  360 :   1 - 0x1
      13'h169: dout  = 8'b00000011; //  361 :   3 - 0x3
      13'h16A: dout  = 8'b00000001; //  362 :   1 - 0x1
      13'h16B: dout  = 8'b00000100; //  363 :   4 - 0x4
      13'h16C: dout  = 8'b00000111; //  364 :   7 - 0x7
      13'h16D: dout  = 8'b00001111; //  365 :  15 - 0xf
      13'h16E: dout  = 8'b00001111; //  366 :  15 - 0xf
      13'h16F: dout  = 8'b00000011; //  367 :   3 - 0x3
      13'h170: dout  = 8'b11111000; //  368 : 248 - 0xf8 -- Sprite 0x17
      13'h171: dout  = 8'b11110000; //  369 : 240 - 0xf0
      13'h172: dout  = 8'b11100000; //  370 : 224 - 0xe0
      13'h173: dout  = 8'b11110000; //  371 : 240 - 0xf0
      13'h174: dout  = 8'b10110000; //  372 : 176 - 0xb0
      13'h175: dout  = 8'b10000000; //  373 : 128 - 0x80
      13'h176: dout  = 8'b11100000; //  374 : 224 - 0xe0
      13'h177: dout  = 8'b11100000; //  375 : 224 - 0xe0
      13'h178: dout  = 8'b11111000; //  376 : 248 - 0xf8
      13'h179: dout  = 8'b11110000; //  377 : 240 - 0xf0
      13'h17A: dout  = 8'b11100000; //  378 : 224 - 0xe0
      13'h17B: dout  = 8'b01110000; //  379 : 112 - 0x70
      13'h17C: dout  = 8'b10110000; //  380 : 176 - 0xb0
      13'h17D: dout  = 8'b10000000; //  381 : 128 - 0x80
      13'h17E: dout  = 8'b11100000; //  382 : 224 - 0xe0
      13'h17F: dout  = 8'b11100000; //  383 : 224 - 0xe0
      13'h180: dout  = 8'b00000011; //  384 :   3 - 0x3 -- Sprite 0x18
      13'h181: dout  = 8'b00111111; //  385 :  63 - 0x3f
      13'h182: dout  = 8'b01111111; //  386 : 127 - 0x7f
      13'h183: dout  = 8'b00011001; //  387 :  25 - 0x19
      13'h184: dout  = 8'b00001001; //  388 :   9 - 0x9
      13'h185: dout  = 8'b00001001; //  389 :   9 - 0x9
      13'h186: dout  = 8'b00101000; //  390 :  40 - 0x28
      13'h187: dout  = 8'b01011100; //  391 :  92 - 0x5c
      13'h188: dout  = 8'b00000000; //  392 :   0 - 0x0
      13'h189: dout  = 8'b00110000; //  393 :  48 - 0x30
      13'h18A: dout  = 8'b01110000; //  394 : 112 - 0x70
      13'h18B: dout  = 8'b01111111; //  395 : 127 - 0x7f
      13'h18C: dout  = 8'b11111111; //  396 : 255 - 0xff
      13'h18D: dout  = 8'b11111111; //  397 : 255 - 0xff
      13'h18E: dout  = 8'b11110111; //  398 : 247 - 0xf7
      13'h18F: dout  = 8'b11110011; //  399 : 243 - 0xf3
      13'h190: dout  = 8'b11111000; //  400 : 248 - 0xf8 -- Sprite 0x19
      13'h191: dout  = 8'b11100000; //  401 : 224 - 0xe0
      13'h192: dout  = 8'b11100000; //  402 : 224 - 0xe0
      13'h193: dout  = 8'b11111100; //  403 : 252 - 0xfc
      13'h194: dout  = 8'b00100110; //  404 :  38 - 0x26
      13'h195: dout  = 8'b00110000; //  405 :  48 - 0x30
      13'h196: dout  = 8'b10000000; //  406 : 128 - 0x80
      13'h197: dout  = 8'b00010000; //  407 :  16 - 0x10
      13'h198: dout  = 8'b00000000; //  408 :   0 - 0x0
      13'h199: dout  = 8'b00011000; //  409 :  24 - 0x18
      13'h19A: dout  = 8'b00010000; //  410 :  16 - 0x10
      13'h19B: dout  = 8'b00000000; //  411 :   0 - 0x0
      13'h19C: dout  = 8'b11111000; //  412 : 248 - 0xf8
      13'h19D: dout  = 8'b11111000; //  413 : 248 - 0xf8
      13'h19E: dout  = 8'b11111110; //  414 : 254 - 0xfe
      13'h19F: dout  = 8'b11111111; //  415 : 255 - 0xff
      13'h1A0: dout  = 8'b00111110; //  416 :  62 - 0x3e -- Sprite 0x1a
      13'h1A1: dout  = 8'b00011110; //  417 :  30 - 0x1e
      13'h1A2: dout  = 8'b00111111; //  418 :  63 - 0x3f
      13'h1A3: dout  = 8'b00111000; //  419 :  56 - 0x38
      13'h1A4: dout  = 8'b00110000; //  420 :  48 - 0x30
      13'h1A5: dout  = 8'b00110000; //  421 :  48 - 0x30
      13'h1A6: dout  = 8'b00000000; //  422 :   0 - 0x0
      13'h1A7: dout  = 8'b00111010; //  423 :  58 - 0x3a
      13'h1A8: dout  = 8'b11100111; //  424 : 231 - 0xe7
      13'h1A9: dout  = 8'b00001111; //  425 :  15 - 0xf
      13'h1AA: dout  = 8'b00001111; //  426 :  15 - 0xf
      13'h1AB: dout  = 8'b00011111; //  427 :  31 - 0x1f
      13'h1AC: dout  = 8'b00011111; //  428 :  31 - 0x1f
      13'h1AD: dout  = 8'b00011111; //  429 :  31 - 0x1f
      13'h1AE: dout  = 8'b00001111; //  430 :  15 - 0xf
      13'h1AF: dout  = 8'b00000111; //  431 :   7 - 0x7
      13'h1B0: dout  = 8'b01111000; //  432 : 120 - 0x78 -- Sprite 0x1b
      13'h1B1: dout  = 8'b00011110; //  433 :  30 - 0x1e
      13'h1B2: dout  = 8'b10000000; //  434 : 128 - 0x80
      13'h1B3: dout  = 8'b11111110; //  435 : 254 - 0xfe
      13'h1B4: dout  = 8'b01111110; //  436 : 126 - 0x7e
      13'h1B5: dout  = 8'b01111110; //  437 : 126 - 0x7e
      13'h1B6: dout  = 8'b01111111; //  438 : 127 - 0x7f
      13'h1B7: dout  = 8'b01111111; //  439 : 127 - 0x7f
      13'h1B8: dout  = 8'b11111111; //  440 : 255 - 0xff
      13'h1B9: dout  = 8'b11111110; //  441 : 254 - 0xfe
      13'h1BA: dout  = 8'b11111100; //  442 : 252 - 0xfc
      13'h1BB: dout  = 8'b11000110; //  443 : 198 - 0xc6
      13'h1BC: dout  = 8'b10001110; //  444 : 142 - 0x8e
      13'h1BD: dout  = 8'b11101110; //  445 : 238 - 0xee
      13'h1BE: dout  = 8'b11111111; //  446 : 255 - 0xff
      13'h1BF: dout  = 8'b11111111; //  447 : 255 - 0xff
      13'h1C0: dout  = 8'b00111100; //  448 :  60 - 0x3c -- Sprite 0x1c
      13'h1C1: dout  = 8'b00111111; //  449 :  63 - 0x3f
      13'h1C2: dout  = 8'b00011111; //  450 :  31 - 0x1f
      13'h1C3: dout  = 8'b00001111; //  451 :  15 - 0xf
      13'h1C4: dout  = 8'b00000111; //  452 :   7 - 0x7
      13'h1C5: dout  = 8'b00111111; //  453 :  63 - 0x3f
      13'h1C6: dout  = 8'b00100001; //  454 :  33 - 0x21
      13'h1C7: dout  = 8'b00100000; //  455 :  32 - 0x20
      13'h1C8: dout  = 8'b00000011; //  456 :   3 - 0x3
      13'h1C9: dout  = 8'b00000000; //  457 :   0 - 0x0
      13'h1CA: dout  = 8'b00000000; //  458 :   0 - 0x0
      13'h1CB: dout  = 8'b00001110; //  459 :  14 - 0xe
      13'h1CC: dout  = 8'b00000111; //  460 :   7 - 0x7
      13'h1CD: dout  = 8'b00111111; //  461 :  63 - 0x3f
      13'h1CE: dout  = 8'b00111111; //  462 :  63 - 0x3f
      13'h1CF: dout  = 8'b00111111; //  463 :  63 - 0x3f
      13'h1D0: dout  = 8'b11111111; //  464 : 255 - 0xff -- Sprite 0x1d
      13'h1D1: dout  = 8'b11111111; //  465 : 255 - 0xff
      13'h1D2: dout  = 8'b11111111; //  466 : 255 - 0xff
      13'h1D3: dout  = 8'b11111110; //  467 : 254 - 0xfe
      13'h1D4: dout  = 8'b11111110; //  468 : 254 - 0xfe
      13'h1D5: dout  = 8'b11111110; //  469 : 254 - 0xfe
      13'h1D6: dout  = 8'b11111100; //  470 : 252 - 0xfc
      13'h1D7: dout  = 8'b01110000; //  471 : 112 - 0x70
      13'h1D8: dout  = 8'b11111111; //  472 : 255 - 0xff
      13'h1D9: dout  = 8'b01111111; //  473 : 127 - 0x7f
      13'h1DA: dout  = 8'b00111111; //  474 :  63 - 0x3f
      13'h1DB: dout  = 8'b00001110; //  475 :  14 - 0xe
      13'h1DC: dout  = 8'b11000000; //  476 : 192 - 0xc0
      13'h1DD: dout  = 8'b11000000; //  477 : 192 - 0xc0
      13'h1DE: dout  = 8'b11100000; //  478 : 224 - 0xe0
      13'h1DF: dout  = 8'b11100000; //  479 : 224 - 0xe0
      13'h1E0: dout  = 8'b00001111; //  480 :  15 - 0xf -- Sprite 0x1e
      13'h1E1: dout  = 8'b10011111; //  481 : 159 - 0x9f
      13'h1E2: dout  = 8'b11001111; //  482 : 207 - 0xcf
      13'h1E3: dout  = 8'b11111111; //  483 : 255 - 0xff
      13'h1E4: dout  = 8'b01111111; //  484 : 127 - 0x7f
      13'h1E5: dout  = 8'b00111111; //  485 :  63 - 0x3f
      13'h1E6: dout  = 8'b00011110; //  486 :  30 - 0x1e
      13'h1E7: dout  = 8'b00001110; //  487 :  14 - 0xe
      13'h1E8: dout  = 8'b00000000; //  488 :   0 - 0x0
      13'h1E9: dout  = 8'b10000000; //  489 : 128 - 0x80
      13'h1EA: dout  = 8'b11001000; //  490 : 200 - 0xc8
      13'h1EB: dout  = 8'b11111110; //  491 : 254 - 0xfe
      13'h1EC: dout  = 8'b01111111; //  492 : 127 - 0x7f
      13'h1ED: dout  = 8'b00111111; //  493 :  63 - 0x3f
      13'h1EE: dout  = 8'b00011110; //  494 :  30 - 0x1e
      13'h1EF: dout  = 8'b00001110; //  495 :  14 - 0xe
      13'h1F0: dout  = 8'b00100000; //  496 :  32 - 0x20 -- Sprite 0x1f
      13'h1F1: dout  = 8'b11000000; //  497 : 192 - 0xc0
      13'h1F2: dout  = 8'b10000000; //  498 : 128 - 0x80
      13'h1F3: dout  = 8'b10000000; //  499 : 128 - 0x80
      13'h1F4: dout  = 8'b00000000; //  500 :   0 - 0x0
      13'h1F5: dout  = 8'b00000000; //  501 :   0 - 0x0
      13'h1F6: dout  = 8'b00000000; //  502 :   0 - 0x0
      13'h1F7: dout  = 8'b00000000; //  503 :   0 - 0x0
      13'h1F8: dout  = 8'b11100000; //  504 : 224 - 0xe0
      13'h1F9: dout  = 8'b00000000; //  505 :   0 - 0x0
      13'h1FA: dout  = 8'b00000000; //  506 :   0 - 0x0
      13'h1FB: dout  = 8'b00000000; //  507 :   0 - 0x0
      13'h1FC: dout  = 8'b00000000; //  508 :   0 - 0x0
      13'h1FD: dout  = 8'b00000000; //  509 :   0 - 0x0
      13'h1FE: dout  = 8'b00000000; //  510 :   0 - 0x0
      13'h1FF: dout  = 8'b00000000; //  511 :   0 - 0x0
      13'h200: dout  = 8'b00000000; //  512 :   0 - 0x0 -- Sprite 0x20
      13'h201: dout  = 8'b00000000; //  513 :   0 - 0x0
      13'h202: dout  = 8'b00000011; //  514 :   3 - 0x3
      13'h203: dout  = 8'b00001111; //  515 :  15 - 0xf
      13'h204: dout  = 8'b00011111; //  516 :  31 - 0x1f
      13'h205: dout  = 8'b00011111; //  517 :  31 - 0x1f
      13'h206: dout  = 8'b00011100; //  518 :  28 - 0x1c
      13'h207: dout  = 8'b00100100; //  519 :  36 - 0x24
      13'h208: dout  = 8'b00000000; //  520 :   0 - 0x0
      13'h209: dout  = 8'b00000000; //  521 :   0 - 0x0
      13'h20A: dout  = 8'b00000000; //  522 :   0 - 0x0
      13'h20B: dout  = 8'b00000000; //  523 :   0 - 0x0
      13'h20C: dout  = 8'b00000000; //  524 :   0 - 0x0
      13'h20D: dout  = 8'b00000000; //  525 :   0 - 0x0
      13'h20E: dout  = 8'b00011111; //  526 :  31 - 0x1f
      13'h20F: dout  = 8'b00111111; //  527 :  63 - 0x3f
      13'h210: dout  = 8'b00000000; //  528 :   0 - 0x0 -- Sprite 0x21
      13'h211: dout  = 8'b00000100; //  529 :   4 - 0x4
      13'h212: dout  = 8'b11100110; //  530 : 230 - 0xe6
      13'h213: dout  = 8'b11100000; //  531 : 224 - 0xe0
      13'h214: dout  = 8'b11111111; //  532 : 255 - 0xff
      13'h215: dout  = 8'b11111111; //  533 : 255 - 0xff
      13'h216: dout  = 8'b10001111; //  534 : 143 - 0x8f
      13'h217: dout  = 8'b10000011; //  535 : 131 - 0x83
      13'h218: dout  = 8'b00001110; //  536 :  14 - 0xe
      13'h219: dout  = 8'b00011111; //  537 :  31 - 0x1f
      13'h21A: dout  = 8'b00011111; //  538 :  31 - 0x1f
      13'h21B: dout  = 8'b00011111; //  539 :  31 - 0x1f
      13'h21C: dout  = 8'b00011111; //  540 :  31 - 0x1f
      13'h21D: dout  = 8'b00000011; //  541 :   3 - 0x3
      13'h21E: dout  = 8'b11111111; //  542 : 255 - 0xff
      13'h21F: dout  = 8'b11111111; //  543 : 255 - 0xff
      13'h220: dout  = 8'b00100110; //  544 :  38 - 0x26 -- Sprite 0x22
      13'h221: dout  = 8'b00100110; //  545 :  38 - 0x26
      13'h222: dout  = 8'b01100000; //  546 :  96 - 0x60
      13'h223: dout  = 8'b01111000; //  547 : 120 - 0x78
      13'h224: dout  = 8'b00011000; //  548 :  24 - 0x18
      13'h225: dout  = 8'b00001111; //  549 :  15 - 0xf
      13'h226: dout  = 8'b01111111; //  550 : 127 - 0x7f
      13'h227: dout  = 8'b11111111; //  551 : 255 - 0xff
      13'h228: dout  = 8'b00111111; //  552 :  63 - 0x3f
      13'h229: dout  = 8'b00111111; //  553 :  63 - 0x3f
      13'h22A: dout  = 8'b01111111; //  554 : 127 - 0x7f
      13'h22B: dout  = 8'b01111111; //  555 : 127 - 0x7f
      13'h22C: dout  = 8'b00011111; //  556 :  31 - 0x1f
      13'h22D: dout  = 8'b00000000; //  557 :   0 - 0x0
      13'h22E: dout  = 8'b01111110; //  558 : 126 - 0x7e
      13'h22F: dout  = 8'b11111111; //  559 : 255 - 0xff
      13'h230: dout  = 8'b00000001; //  560 :   1 - 0x1 -- Sprite 0x23
      13'h231: dout  = 8'b00100001; //  561 :  33 - 0x21
      13'h232: dout  = 8'b11111110; //  562 : 254 - 0xfe
      13'h233: dout  = 8'b01111010; //  563 : 122 - 0x7a
      13'h234: dout  = 8'b00000110; //  564 :   6 - 0x6
      13'h235: dout  = 8'b11111110; //  565 : 254 - 0xfe
      13'h236: dout  = 8'b11111100; //  566 : 252 - 0xfc
      13'h237: dout  = 8'b11111100; //  567 : 252 - 0xfc
      13'h238: dout  = 8'b11111111; //  568 : 255 - 0xff
      13'h239: dout  = 8'b11111111; //  569 : 255 - 0xff
      13'h23A: dout  = 8'b11111110; //  570 : 254 - 0xfe
      13'h23B: dout  = 8'b11111110; //  571 : 254 - 0xfe
      13'h23C: dout  = 8'b11111110; //  572 : 254 - 0xfe
      13'h23D: dout  = 8'b11011110; //  573 : 222 - 0xde
      13'h23E: dout  = 8'b01011100; //  574 :  92 - 0x5c
      13'h23F: dout  = 8'b01101100; //  575 : 108 - 0x6c
      13'h240: dout  = 8'b11111111; //  576 : 255 - 0xff -- Sprite 0x24
      13'h241: dout  = 8'b11001111; //  577 : 207 - 0xcf
      13'h242: dout  = 8'b10000111; //  578 : 135 - 0x87
      13'h243: dout  = 8'b00000111; //  579 :   7 - 0x7
      13'h244: dout  = 8'b00000111; //  580 :   7 - 0x7
      13'h245: dout  = 8'b00001111; //  581 :  15 - 0xf
      13'h246: dout  = 8'b00011111; //  582 :  31 - 0x1f
      13'h247: dout  = 8'b00011111; //  583 :  31 - 0x1f
      13'h248: dout  = 8'b11111111; //  584 : 255 - 0xff
      13'h249: dout  = 8'b11111111; //  585 : 255 - 0xff
      13'h24A: dout  = 8'b11111110; //  586 : 254 - 0xfe
      13'h24B: dout  = 8'b11111100; //  587 : 252 - 0xfc
      13'h24C: dout  = 8'b11111000; //  588 : 248 - 0xf8
      13'h24D: dout  = 8'b10110000; //  589 : 176 - 0xb0
      13'h24E: dout  = 8'b01100000; //  590 :  96 - 0x60
      13'h24F: dout  = 8'b00000000; //  591 :   0 - 0x0
      13'h250: dout  = 8'b11111000; //  592 : 248 - 0xf8 -- Sprite 0x25
      13'h251: dout  = 8'b11111000; //  593 : 248 - 0xf8
      13'h252: dout  = 8'b11110000; //  594 : 240 - 0xf0
      13'h253: dout  = 8'b10111000; //  595 : 184 - 0xb8
      13'h254: dout  = 8'b11111000; //  596 : 248 - 0xf8
      13'h255: dout  = 8'b11111001; //  597 : 249 - 0xf9
      13'h256: dout  = 8'b11111011; //  598 : 251 - 0xfb
      13'h257: dout  = 8'b11111111; //  599 : 255 - 0xff
      13'h258: dout  = 8'b00101000; //  600 :  40 - 0x28
      13'h259: dout  = 8'b00110000; //  601 :  48 - 0x30
      13'h25A: dout  = 8'b00011000; //  602 :  24 - 0x18
      13'h25B: dout  = 8'b01000000; //  603 :  64 - 0x40
      13'h25C: dout  = 8'b00000000; //  604 :   0 - 0x0
      13'h25D: dout  = 8'b00000001; //  605 :   1 - 0x1
      13'h25E: dout  = 8'b00000011; //  606 :   3 - 0x3
      13'h25F: dout  = 8'b00001111; //  607 :  15 - 0xf
      13'h260: dout  = 8'b00011111; //  608 :  31 - 0x1f -- Sprite 0x26
      13'h261: dout  = 8'b11111111; //  609 : 255 - 0xff
      13'h262: dout  = 8'b11111111; //  610 : 255 - 0xff
      13'h263: dout  = 8'b11111111; //  611 : 255 - 0xff
      13'h264: dout  = 8'b11111111; //  612 : 255 - 0xff
      13'h265: dout  = 8'b11111110; //  613 : 254 - 0xfe
      13'h266: dout  = 8'b11000000; //  614 : 192 - 0xc0
      13'h267: dout  = 8'b10000000; //  615 : 128 - 0x80
      13'h268: dout  = 8'b00010000; //  616 :  16 - 0x10
      13'h269: dout  = 8'b11101100; //  617 : 236 - 0xec
      13'h26A: dout  = 8'b11100011; //  618 : 227 - 0xe3
      13'h26B: dout  = 8'b11100000; //  619 : 224 - 0xe0
      13'h26C: dout  = 8'b11100000; //  620 : 224 - 0xe0
      13'h26D: dout  = 8'b11100000; //  621 : 224 - 0xe0
      13'h26E: dout  = 8'b11000000; //  622 : 192 - 0xc0
      13'h26F: dout  = 8'b10000000; //  623 : 128 - 0x80
      13'h270: dout  = 8'b11111111; //  624 : 255 - 0xff -- Sprite 0x27
      13'h271: dout  = 8'b11111111; //  625 : 255 - 0xff
      13'h272: dout  = 8'b11111111; //  626 : 255 - 0xff
      13'h273: dout  = 8'b00111111; //  627 :  63 - 0x3f
      13'h274: dout  = 8'b00000000; //  628 :   0 - 0x0
      13'h275: dout  = 8'b00000000; //  629 :   0 - 0x0
      13'h276: dout  = 8'b00000000; //  630 :   0 - 0x0
      13'h277: dout  = 8'b00000000; //  631 :   0 - 0x0
      13'h278: dout  = 8'b00001111; //  632 :  15 - 0xf
      13'h279: dout  = 8'b00001111; //  633 :  15 - 0xf
      13'h27A: dout  = 8'b00001111; //  634 :  15 - 0xf
      13'h27B: dout  = 8'b00001111; //  635 :  15 - 0xf
      13'h27C: dout  = 8'b00000000; //  636 :   0 - 0x0
      13'h27D: dout  = 8'b00000000; //  637 :   0 - 0x0
      13'h27E: dout  = 8'b00000000; //  638 :   0 - 0x0
      13'h27F: dout  = 8'b00000000; //  639 :   0 - 0x0
      13'h280: dout  = 8'b00010011; //  640 :  19 - 0x13 -- Sprite 0x28
      13'h281: dout  = 8'b00110011; //  641 :  51 - 0x33
      13'h282: dout  = 8'b00110000; //  642 :  48 - 0x30
      13'h283: dout  = 8'b00011000; //  643 :  24 - 0x18
      13'h284: dout  = 8'b00000100; //  644 :   4 - 0x4
      13'h285: dout  = 8'b00001111; //  645 :  15 - 0xf
      13'h286: dout  = 8'b00011111; //  646 :  31 - 0x1f
      13'h287: dout  = 8'b00011111; //  647 :  31 - 0x1f
      13'h288: dout  = 8'b00011111; //  648 :  31 - 0x1f
      13'h289: dout  = 8'b00111111; //  649 :  63 - 0x3f
      13'h28A: dout  = 8'b00111111; //  650 :  63 - 0x3f
      13'h28B: dout  = 8'b00011111; //  651 :  31 - 0x1f
      13'h28C: dout  = 8'b00000111; //  652 :   7 - 0x7
      13'h28D: dout  = 8'b00001001; //  653 :   9 - 0x9
      13'h28E: dout  = 8'b00010011; //  654 :  19 - 0x13
      13'h28F: dout  = 8'b00010111; //  655 :  23 - 0x17
      13'h290: dout  = 8'b00000000; //  656 :   0 - 0x0 -- Sprite 0x29
      13'h291: dout  = 8'b00010000; //  657 :  16 - 0x10
      13'h292: dout  = 8'b01111110; //  658 : 126 - 0x7e
      13'h293: dout  = 8'b00110000; //  659 :  48 - 0x30
      13'h294: dout  = 8'b11100000; //  660 : 224 - 0xe0
      13'h295: dout  = 8'b11110000; //  661 : 240 - 0xf0
      13'h296: dout  = 8'b11110000; //  662 : 240 - 0xf0
      13'h297: dout  = 8'b11100000; //  663 : 224 - 0xe0
      13'h298: dout  = 8'b11111111; //  664 : 255 - 0xff
      13'h299: dout  = 8'b11111111; //  665 : 255 - 0xff
      13'h29A: dout  = 8'b11111110; //  666 : 254 - 0xfe
      13'h29B: dout  = 8'b11111111; //  667 : 255 - 0xff
      13'h29C: dout  = 8'b11111110; //  668 : 254 - 0xfe
      13'h29D: dout  = 8'b11111100; //  669 : 252 - 0xfc
      13'h29E: dout  = 8'b11111000; //  670 : 248 - 0xf8
      13'h29F: dout  = 8'b11100000; //  671 : 224 - 0xe0
      13'h2A0: dout  = 8'b00011111; //  672 :  31 - 0x1f -- Sprite 0x2a
      13'h2A1: dout  = 8'b00011111; //  673 :  31 - 0x1f
      13'h2A2: dout  = 8'b00001111; //  674 :  15 - 0xf
      13'h2A3: dout  = 8'b00001111; //  675 :  15 - 0xf
      13'h2A4: dout  = 8'b00001111; //  676 :  15 - 0xf
      13'h2A5: dout  = 8'b00011111; //  677 :  31 - 0x1f
      13'h2A6: dout  = 8'b00011111; //  678 :  31 - 0x1f
      13'h2A7: dout  = 8'b00011111; //  679 :  31 - 0x1f
      13'h2A8: dout  = 8'b00010111; //  680 :  23 - 0x17
      13'h2A9: dout  = 8'b00010111; //  681 :  23 - 0x17
      13'h2AA: dout  = 8'b00000011; //  682 :   3 - 0x3
      13'h2AB: dout  = 8'b00000000; //  683 :   0 - 0x0
      13'h2AC: dout  = 8'b00000000; //  684 :   0 - 0x0
      13'h2AD: dout  = 8'b00000000; //  685 :   0 - 0x0
      13'h2AE: dout  = 8'b00000000; //  686 :   0 - 0x0
      13'h2AF: dout  = 8'b00000000; //  687 :   0 - 0x0
      13'h2B0: dout  = 8'b11110000; //  688 : 240 - 0xf0 -- Sprite 0x2b
      13'h2B1: dout  = 8'b11110000; //  689 : 240 - 0xf0
      13'h2B2: dout  = 8'b11111000; //  690 : 248 - 0xf8
      13'h2B3: dout  = 8'b11111000; //  691 : 248 - 0xf8
      13'h2B4: dout  = 8'b10111000; //  692 : 184 - 0xb8
      13'h2B5: dout  = 8'b11111000; //  693 : 248 - 0xf8
      13'h2B6: dout  = 8'b11111000; //  694 : 248 - 0xf8
      13'h2B7: dout  = 8'b11111000; //  695 : 248 - 0xf8
      13'h2B8: dout  = 8'b11010000; //  696 : 208 - 0xd0
      13'h2B9: dout  = 8'b10010000; //  697 : 144 - 0x90
      13'h2BA: dout  = 8'b00011000; //  698 :  24 - 0x18
      13'h2BB: dout  = 8'b00001000; //  699 :   8 - 0x8
      13'h2BC: dout  = 8'b01000000; //  700 :  64 - 0x40
      13'h2BD: dout  = 8'b00000000; //  701 :   0 - 0x0
      13'h2BE: dout  = 8'b00000000; //  702 :   0 - 0x0
      13'h2BF: dout  = 8'b00000000; //  703 :   0 - 0x0
      13'h2C0: dout  = 8'b00111111; //  704 :  63 - 0x3f -- Sprite 0x2c
      13'h2C1: dout  = 8'b11111111; //  705 : 255 - 0xff
      13'h2C2: dout  = 8'b11111111; //  706 : 255 - 0xff
      13'h2C3: dout  = 8'b11111111; //  707 : 255 - 0xff
      13'h2C4: dout  = 8'b11110110; //  708 : 246 - 0xf6
      13'h2C5: dout  = 8'b11000110; //  709 : 198 - 0xc6
      13'h2C6: dout  = 8'b10000100; //  710 : 132 - 0x84
      13'h2C7: dout  = 8'b00000000; //  711 :   0 - 0x0
      13'h2C8: dout  = 8'b00110000; //  712 :  48 - 0x30
      13'h2C9: dout  = 8'b11110000; //  713 : 240 - 0xf0
      13'h2CA: dout  = 8'b11110000; //  714 : 240 - 0xf0
      13'h2CB: dout  = 8'b11110001; //  715 : 241 - 0xf1
      13'h2CC: dout  = 8'b11110110; //  716 : 246 - 0xf6
      13'h2CD: dout  = 8'b11000110; //  717 : 198 - 0xc6
      13'h2CE: dout  = 8'b10000100; //  718 : 132 - 0x84
      13'h2CF: dout  = 8'b00000000; //  719 :   0 - 0x0
      13'h2D0: dout  = 8'b11110000; //  720 : 240 - 0xf0 -- Sprite 0x2d
      13'h2D1: dout  = 8'b11100000; //  721 : 224 - 0xe0
      13'h2D2: dout  = 8'b10000000; //  722 : 128 - 0x80
      13'h2D3: dout  = 8'b00000000; //  723 :   0 - 0x0
      13'h2D4: dout  = 8'b00000000; //  724 :   0 - 0x0
      13'h2D5: dout  = 8'b00000000; //  725 :   0 - 0x0
      13'h2D6: dout  = 8'b00000000; //  726 :   0 - 0x0
      13'h2D7: dout  = 8'b00000000; //  727 :   0 - 0x0
      13'h2D8: dout  = 8'b00000000; //  728 :   0 - 0x0
      13'h2D9: dout  = 8'b00000000; //  729 :   0 - 0x0
      13'h2DA: dout  = 8'b00000000; //  730 :   0 - 0x0
      13'h2DB: dout  = 8'b00000000; //  731 :   0 - 0x0
      13'h2DC: dout  = 8'b00000000; //  732 :   0 - 0x0
      13'h2DD: dout  = 8'b00000000; //  733 :   0 - 0x0
      13'h2DE: dout  = 8'b00000000; //  734 :   0 - 0x0
      13'h2DF: dout  = 8'b00000000; //  735 :   0 - 0x0
      13'h2E0: dout  = 8'b00011111; //  736 :  31 - 0x1f -- Sprite 0x2e
      13'h2E1: dout  = 8'b00011111; //  737 :  31 - 0x1f
      13'h2E2: dout  = 8'b00111111; //  738 :  63 - 0x3f
      13'h2E3: dout  = 8'b00111111; //  739 :  63 - 0x3f
      13'h2E4: dout  = 8'b00011111; //  740 :  31 - 0x1f
      13'h2E5: dout  = 8'b00001111; //  741 :  15 - 0xf
      13'h2E6: dout  = 8'b00001111; //  742 :  15 - 0xf
      13'h2E7: dout  = 8'b00011111; //  743 :  31 - 0x1f
      13'h2E8: dout  = 8'b00011111; //  744 :  31 - 0x1f
      13'h2E9: dout  = 8'b00011111; //  745 :  31 - 0x1f
      13'h2EA: dout  = 8'b00111111; //  746 :  63 - 0x3f
      13'h2EB: dout  = 8'b00111110; //  747 :  62 - 0x3e
      13'h2EC: dout  = 8'b01111100; //  748 : 124 - 0x7c
      13'h2ED: dout  = 8'b01111000; //  749 : 120 - 0x78
      13'h2EE: dout  = 8'b11110000; //  750 : 240 - 0xf0
      13'h2EF: dout  = 8'b11100000; //  751 : 224 - 0xe0
      13'h2F0: dout  = 8'b11110000; //  752 : 240 - 0xf0 -- Sprite 0x2f
      13'h2F1: dout  = 8'b11110000; //  753 : 240 - 0xf0
      13'h2F2: dout  = 8'b11111000; //  754 : 248 - 0xf8
      13'h2F3: dout  = 8'b11111000; //  755 : 248 - 0xf8
      13'h2F4: dout  = 8'b10111000; //  756 : 184 - 0xb8
      13'h2F5: dout  = 8'b11111000; //  757 : 248 - 0xf8
      13'h2F6: dout  = 8'b11111000; //  758 : 248 - 0xf8
      13'h2F7: dout  = 8'b11110000; //  759 : 240 - 0xf0
      13'h2F8: dout  = 8'b10110000; //  760 : 176 - 0xb0
      13'h2F9: dout  = 8'b10010000; //  761 : 144 - 0x90
      13'h2FA: dout  = 8'b00011000; //  762 :  24 - 0x18
      13'h2FB: dout  = 8'b00001000; //  763 :   8 - 0x8
      13'h2FC: dout  = 8'b01000000; //  764 :  64 - 0x40
      13'h2FD: dout  = 8'b00000000; //  765 :   0 - 0x0
      13'h2FE: dout  = 8'b00000000; //  766 :   0 - 0x0
      13'h2FF: dout  = 8'b00000000; //  767 :   0 - 0x0
      13'h300: dout  = 8'b11100000; //  768 : 224 - 0xe0 -- Sprite 0x30
      13'h301: dout  = 8'b11110000; //  769 : 240 - 0xf0
      13'h302: dout  = 8'b11110000; //  770 : 240 - 0xf0
      13'h303: dout  = 8'b11110000; //  771 : 240 - 0xf0
      13'h304: dout  = 8'b11110000; //  772 : 240 - 0xf0
      13'h305: dout  = 8'b11110000; //  773 : 240 - 0xf0
      13'h306: dout  = 8'b11111000; //  774 : 248 - 0xf8
      13'h307: dout  = 8'b11110000; //  775 : 240 - 0xf0
      13'h308: dout  = 8'b11000000; //  776 : 192 - 0xc0
      13'h309: dout  = 8'b11100000; //  777 : 224 - 0xe0
      13'h30A: dout  = 8'b11111100; //  778 : 252 - 0xfc
      13'h30B: dout  = 8'b11111110; //  779 : 254 - 0xfe
      13'h30C: dout  = 8'b11111111; //  780 : 255 - 0xff
      13'h30D: dout  = 8'b01111111; //  781 : 127 - 0x7f
      13'h30E: dout  = 8'b00000011; //  782 :   3 - 0x3
      13'h30F: dout  = 8'b00000000; //  783 :   0 - 0x0
      13'h310: dout  = 8'b00011111; //  784 :  31 - 0x1f -- Sprite 0x31
      13'h311: dout  = 8'b00011111; //  785 :  31 - 0x1f
      13'h312: dout  = 8'b00011111; //  786 :  31 - 0x1f
      13'h313: dout  = 8'b00111111; //  787 :  63 - 0x3f
      13'h314: dout  = 8'b00111110; //  788 :  62 - 0x3e
      13'h315: dout  = 8'b00111100; //  789 :  60 - 0x3c
      13'h316: dout  = 8'b00111000; //  790 :  56 - 0x38
      13'h317: dout  = 8'b00011000; //  791 :  24 - 0x18
      13'h318: dout  = 8'b00000000; //  792 :   0 - 0x0
      13'h319: dout  = 8'b00000000; //  793 :   0 - 0x0
      13'h31A: dout  = 8'b00010000; //  794 :  16 - 0x10
      13'h31B: dout  = 8'b00111000; //  795 :  56 - 0x38
      13'h31C: dout  = 8'b00111110; //  796 :  62 - 0x3e
      13'h31D: dout  = 8'b00111100; //  797 :  60 - 0x3c
      13'h31E: dout  = 8'b00111000; //  798 :  56 - 0x38
      13'h31F: dout  = 8'b00011000; //  799 :  24 - 0x18
      13'h320: dout  = 8'b00000000; //  800 :   0 - 0x0 -- Sprite 0x32
      13'h321: dout  = 8'b00000011; //  801 :   3 - 0x3
      13'h322: dout  = 8'b00000111; //  802 :   7 - 0x7
      13'h323: dout  = 8'b00000111; //  803 :   7 - 0x7
      13'h324: dout  = 8'b00001010; //  804 :  10 - 0xa
      13'h325: dout  = 8'b00001011; //  805 :  11 - 0xb
      13'h326: dout  = 8'b00001100; //  806 :  12 - 0xc
      13'h327: dout  = 8'b00000000; //  807 :   0 - 0x0
      13'h328: dout  = 8'b00000000; //  808 :   0 - 0x0
      13'h329: dout  = 8'b00000000; //  809 :   0 - 0x0
      13'h32A: dout  = 8'b00000000; //  810 :   0 - 0x0
      13'h32B: dout  = 8'b00000111; //  811 :   7 - 0x7
      13'h32C: dout  = 8'b00001111; //  812 :  15 - 0xf
      13'h32D: dout  = 8'b00001111; //  813 :  15 - 0xf
      13'h32E: dout  = 8'b00001111; //  814 :  15 - 0xf
      13'h32F: dout  = 8'b00000011; //  815 :   3 - 0x3
      13'h330: dout  = 8'b00000000; //  816 :   0 - 0x0 -- Sprite 0x33
      13'h331: dout  = 8'b11100000; //  817 : 224 - 0xe0
      13'h332: dout  = 8'b11111100; //  818 : 252 - 0xfc
      13'h333: dout  = 8'b00100000; //  819 :  32 - 0x20
      13'h334: dout  = 8'b00100000; //  820 :  32 - 0x20
      13'h335: dout  = 8'b00010000; //  821 :  16 - 0x10
      13'h336: dout  = 8'b00111100; //  822 :  60 - 0x3c
      13'h337: dout  = 8'b00000000; //  823 :   0 - 0x0
      13'h338: dout  = 8'b00000000; //  824 :   0 - 0x0
      13'h339: dout  = 8'b00000000; //  825 :   0 - 0x0
      13'h33A: dout  = 8'b00000000; //  826 :   0 - 0x0
      13'h33B: dout  = 8'b11110000; //  827 : 240 - 0xf0
      13'h33C: dout  = 8'b11111100; //  828 : 252 - 0xfc
      13'h33D: dout  = 8'b11111110; //  829 : 254 - 0xfe
      13'h33E: dout  = 8'b11111100; //  830 : 252 - 0xfc
      13'h33F: dout  = 8'b11111000; //  831 : 248 - 0xf8
      13'h340: dout  = 8'b00000111; //  832 :   7 - 0x7 -- Sprite 0x34
      13'h341: dout  = 8'b00000111; //  833 :   7 - 0x7
      13'h342: dout  = 8'b00000111; //  834 :   7 - 0x7
      13'h343: dout  = 8'b00011111; //  835 :  31 - 0x1f
      13'h344: dout  = 8'b00011111; //  836 :  31 - 0x1f
      13'h345: dout  = 8'b00111110; //  837 :  62 - 0x3e
      13'h346: dout  = 8'b00100001; //  838 :  33 - 0x21
      13'h347: dout  = 8'b00000001; //  839 :   1 - 0x1
      13'h348: dout  = 8'b00000111; //  840 :   7 - 0x7
      13'h349: dout  = 8'b00001111; //  841 :  15 - 0xf
      13'h34A: dout  = 8'b00011011; //  842 :  27 - 0x1b
      13'h34B: dout  = 8'b00011000; //  843 :  24 - 0x18
      13'h34C: dout  = 8'b00010000; //  844 :  16 - 0x10
      13'h34D: dout  = 8'b00110000; //  845 :  48 - 0x30
      13'h34E: dout  = 8'b00100001; //  846 :  33 - 0x21
      13'h34F: dout  = 8'b00000001; //  847 :   1 - 0x1
      13'h350: dout  = 8'b11100000; //  848 : 224 - 0xe0 -- Sprite 0x35
      13'h351: dout  = 8'b11100000; //  849 : 224 - 0xe0
      13'h352: dout  = 8'b11100000; //  850 : 224 - 0xe0
      13'h353: dout  = 8'b11110000; //  851 : 240 - 0xf0
      13'h354: dout  = 8'b11110000; //  852 : 240 - 0xf0
      13'h355: dout  = 8'b11100000; //  853 : 224 - 0xe0
      13'h356: dout  = 8'b11000000; //  854 : 192 - 0xc0
      13'h357: dout  = 8'b11100000; //  855 : 224 - 0xe0
      13'h358: dout  = 8'b10101000; //  856 : 168 - 0xa8
      13'h359: dout  = 8'b11111100; //  857 : 252 - 0xfc
      13'h35A: dout  = 8'b11111000; //  858 : 248 - 0xf8
      13'h35B: dout  = 8'b00000000; //  859 :   0 - 0x0
      13'h35C: dout  = 8'b00000000; //  860 :   0 - 0x0
      13'h35D: dout  = 8'b00000000; //  861 :   0 - 0x0
      13'h35E: dout  = 8'b11000000; //  862 : 192 - 0xc0
      13'h35F: dout  = 8'b11100000; //  863 : 224 - 0xe0
      13'h360: dout  = 8'b00000111; //  864 :   7 - 0x7 -- Sprite 0x36
      13'h361: dout  = 8'b00001111; //  865 :  15 - 0xf
      13'h362: dout  = 8'b00001110; //  866 :  14 - 0xe
      13'h363: dout  = 8'b00010100; //  867 :  20 - 0x14
      13'h364: dout  = 8'b00010110; //  868 :  22 - 0x16
      13'h365: dout  = 8'b00011000; //  869 :  24 - 0x18
      13'h366: dout  = 8'b00000000; //  870 :   0 - 0x0
      13'h367: dout  = 8'b00111111; //  871 :  63 - 0x3f
      13'h368: dout  = 8'b00000000; //  872 :   0 - 0x0
      13'h369: dout  = 8'b00000000; //  873 :   0 - 0x0
      13'h36A: dout  = 8'b00001111; //  874 :  15 - 0xf
      13'h36B: dout  = 8'b00011111; //  875 :  31 - 0x1f
      13'h36C: dout  = 8'b00011111; //  876 :  31 - 0x1f
      13'h36D: dout  = 8'b00011111; //  877 :  31 - 0x1f
      13'h36E: dout  = 8'b00000111; //  878 :   7 - 0x7
      13'h36F: dout  = 8'b00111100; //  879 :  60 - 0x3c
      13'h370: dout  = 8'b11000000; //  880 : 192 - 0xc0 -- Sprite 0x37
      13'h371: dout  = 8'b11111000; //  881 : 248 - 0xf8
      13'h372: dout  = 8'b01000000; //  882 :  64 - 0x40
      13'h373: dout  = 8'b01000000; //  883 :  64 - 0x40
      13'h374: dout  = 8'b00100000; //  884 :  32 - 0x20
      13'h375: dout  = 8'b01111000; //  885 : 120 - 0x78
      13'h376: dout  = 8'b00000000; //  886 :   0 - 0x0
      13'h377: dout  = 8'b11000000; //  887 : 192 - 0xc0
      13'h378: dout  = 8'b00000000; //  888 :   0 - 0x0
      13'h379: dout  = 8'b00000000; //  889 :   0 - 0x0
      13'h37A: dout  = 8'b11100000; //  890 : 224 - 0xe0
      13'h37B: dout  = 8'b11111000; //  891 : 248 - 0xf8
      13'h37C: dout  = 8'b11111100; //  892 : 252 - 0xfc
      13'h37D: dout  = 8'b11111000; //  893 : 248 - 0xf8
      13'h37E: dout  = 8'b11110000; //  894 : 240 - 0xf0
      13'h37F: dout  = 8'b11000000; //  895 : 192 - 0xc0
      13'h380: dout  = 8'b00111111; //  896 :  63 - 0x3f -- Sprite 0x38
      13'h381: dout  = 8'b00001110; //  897 :  14 - 0xe
      13'h382: dout  = 8'b00001111; //  898 :  15 - 0xf
      13'h383: dout  = 8'b00011111; //  899 :  31 - 0x1f
      13'h384: dout  = 8'b00111111; //  900 :  63 - 0x3f
      13'h385: dout  = 8'b01111100; //  901 : 124 - 0x7c
      13'h386: dout  = 8'b01110000; //  902 : 112 - 0x70
      13'h387: dout  = 8'b00111000; //  903 :  56 - 0x38
      13'h388: dout  = 8'b11111100; //  904 : 252 - 0xfc
      13'h389: dout  = 8'b11101101; //  905 : 237 - 0xed
      13'h38A: dout  = 8'b11000000; //  906 : 192 - 0xc0
      13'h38B: dout  = 8'b00000000; //  907 :   0 - 0x0
      13'h38C: dout  = 8'b00000000; //  908 :   0 - 0x0
      13'h38D: dout  = 8'b01100000; //  909 :  96 - 0x60
      13'h38E: dout  = 8'b01110000; //  910 : 112 - 0x70
      13'h38F: dout  = 8'b00111000; //  911 :  56 - 0x38
      13'h390: dout  = 8'b11110000; //  912 : 240 - 0xf0 -- Sprite 0x39
      13'h391: dout  = 8'b11111000; //  913 : 248 - 0xf8
      13'h392: dout  = 8'b11100100; //  914 : 228 - 0xe4
      13'h393: dout  = 8'b11111100; //  915 : 252 - 0xfc
      13'h394: dout  = 8'b11111100; //  916 : 252 - 0xfc
      13'h395: dout  = 8'b01111100; //  917 : 124 - 0x7c
      13'h396: dout  = 8'b00000000; //  918 :   0 - 0x0
      13'h397: dout  = 8'b00000000; //  919 :   0 - 0x0
      13'h398: dout  = 8'b01111110; //  920 : 126 - 0x7e
      13'h399: dout  = 8'b00011110; //  921 :  30 - 0x1e
      13'h39A: dout  = 8'b00000100; //  922 :   4 - 0x4
      13'h39B: dout  = 8'b00001100; //  923 :  12 - 0xc
      13'h39C: dout  = 8'b00001100; //  924 :  12 - 0xc
      13'h39D: dout  = 8'b00001100; //  925 :  12 - 0xc
      13'h39E: dout  = 8'b00000000; //  926 :   0 - 0x0
      13'h39F: dout  = 8'b00000000; //  927 :   0 - 0x0
      13'h3A0: dout  = 8'b00000111; //  928 :   7 - 0x7 -- Sprite 0x3a
      13'h3A1: dout  = 8'b00001111; //  929 :  15 - 0xf
      13'h3A2: dout  = 8'b00001110; //  930 :  14 - 0xe
      13'h3A3: dout  = 8'b00010100; //  931 :  20 - 0x14
      13'h3A4: dout  = 8'b00010110; //  932 :  22 - 0x16
      13'h3A5: dout  = 8'b00011000; //  933 :  24 - 0x18
      13'h3A6: dout  = 8'b00000000; //  934 :   0 - 0x0
      13'h3A7: dout  = 8'b00001111; //  935 :  15 - 0xf
      13'h3A8: dout  = 8'b00000000; //  936 :   0 - 0x0
      13'h3A9: dout  = 8'b00000000; //  937 :   0 - 0x0
      13'h3AA: dout  = 8'b00001111; //  938 :  15 - 0xf
      13'h3AB: dout  = 8'b00011111; //  939 :  31 - 0x1f
      13'h3AC: dout  = 8'b00011111; //  940 :  31 - 0x1f
      13'h3AD: dout  = 8'b00011111; //  941 :  31 - 0x1f
      13'h3AE: dout  = 8'b00000111; //  942 :   7 - 0x7
      13'h3AF: dout  = 8'b00001101; //  943 :  13 - 0xd
      13'h3B0: dout  = 8'b00011111; //  944 :  31 - 0x1f -- Sprite 0x3b
      13'h3B1: dout  = 8'b00011111; //  945 :  31 - 0x1f
      13'h3B2: dout  = 8'b00011111; //  946 :  31 - 0x1f
      13'h3B3: dout  = 8'b00011100; //  947 :  28 - 0x1c
      13'h3B4: dout  = 8'b00001100; //  948 :  12 - 0xc
      13'h3B5: dout  = 8'b00000111; //  949 :   7 - 0x7
      13'h3B6: dout  = 8'b00000111; //  950 :   7 - 0x7
      13'h3B7: dout  = 8'b00000111; //  951 :   7 - 0x7
      13'h3B8: dout  = 8'b00011110; //  952 :  30 - 0x1e
      13'h3B9: dout  = 8'b00011100; //  953 :  28 - 0x1c
      13'h3BA: dout  = 8'b00011110; //  954 :  30 - 0x1e
      13'h3BB: dout  = 8'b00001111; //  955 :  15 - 0xf
      13'h3BC: dout  = 8'b00000111; //  956 :   7 - 0x7
      13'h3BD: dout  = 8'b00000000; //  957 :   0 - 0x0
      13'h3BE: dout  = 8'b00000111; //  958 :   7 - 0x7
      13'h3BF: dout  = 8'b00000111; //  959 :   7 - 0x7
      13'h3C0: dout  = 8'b11100000; //  960 : 224 - 0xe0 -- Sprite 0x3c
      13'h3C1: dout  = 8'b01100000; //  961 :  96 - 0x60
      13'h3C2: dout  = 8'b11110000; //  962 : 240 - 0xf0
      13'h3C3: dout  = 8'b01110000; //  963 : 112 - 0x70
      13'h3C4: dout  = 8'b11100000; //  964 : 224 - 0xe0
      13'h3C5: dout  = 8'b11100000; //  965 : 224 - 0xe0
      13'h3C6: dout  = 8'b11110000; //  966 : 240 - 0xf0
      13'h3C7: dout  = 8'b10000000; //  967 : 128 - 0x80
      13'h3C8: dout  = 8'b01100000; //  968 :  96 - 0x60
      13'h3C9: dout  = 8'b10010000; //  969 : 144 - 0x90
      13'h3CA: dout  = 8'b00000000; //  970 :   0 - 0x0
      13'h3CB: dout  = 8'b10000000; //  971 : 128 - 0x80
      13'h3CC: dout  = 8'b00000000; //  972 :   0 - 0x0
      13'h3CD: dout  = 8'b11100000; //  973 : 224 - 0xe0
      13'h3CE: dout  = 8'b11110000; //  974 : 240 - 0xf0
      13'h3CF: dout  = 8'b10000000; //  975 : 128 - 0x80
      13'h3D0: dout  = 8'b00000111; //  976 :   7 - 0x7 -- Sprite 0x3d
      13'h3D1: dout  = 8'b00011111; //  977 :  31 - 0x1f
      13'h3D2: dout  = 8'b00111111; //  978 :  63 - 0x3f
      13'h3D3: dout  = 8'b00010010; //  979 :  18 - 0x12
      13'h3D4: dout  = 8'b00010011; //  980 :  19 - 0x13
      13'h3D5: dout  = 8'b00001000; //  981 :   8 - 0x8
      13'h3D6: dout  = 8'b00011111; //  982 :  31 - 0x1f
      13'h3D7: dout  = 8'b00110001; //  983 :  49 - 0x31
      13'h3D8: dout  = 8'b00000000; //  984 :   0 - 0x0
      13'h3D9: dout  = 8'b00010000; //  985 :  16 - 0x10
      13'h3DA: dout  = 8'b00111111; //  986 :  63 - 0x3f
      13'h3DB: dout  = 8'b01111111; //  987 : 127 - 0x7f
      13'h3DC: dout  = 8'b01111111; //  988 : 127 - 0x7f
      13'h3DD: dout  = 8'b00111111; //  989 :  63 - 0x3f
      13'h3DE: dout  = 8'b00000011; //  990 :   3 - 0x3
      13'h3DF: dout  = 8'b00001111; //  991 :  15 - 0xf
      13'h3E0: dout  = 8'b11000000; //  992 : 192 - 0xc0 -- Sprite 0x3e
      13'h3E1: dout  = 8'b11110000; //  993 : 240 - 0xf0
      13'h3E2: dout  = 8'b01000000; //  994 :  64 - 0x40
      13'h3E3: dout  = 8'b00000000; //  995 :   0 - 0x0
      13'h3E4: dout  = 8'b00110000; //  996 :  48 - 0x30
      13'h3E5: dout  = 8'b00011000; //  997 :  24 - 0x18
      13'h3E6: dout  = 8'b11000000; //  998 : 192 - 0xc0
      13'h3E7: dout  = 8'b11111000; //  999 : 248 - 0xf8
      13'h3E8: dout  = 8'b00000000; // 1000 :   0 - 0x0
      13'h3E9: dout  = 8'b00000000; // 1001 :   0 - 0x0
      13'h3EA: dout  = 8'b11100000; // 1002 : 224 - 0xe0
      13'h3EB: dout  = 8'b11111000; // 1003 : 248 - 0xf8
      13'h3EC: dout  = 8'b11111100; // 1004 : 252 - 0xfc
      13'h3ED: dout  = 8'b11111000; // 1005 : 248 - 0xf8
      13'h3EE: dout  = 8'b10110000; // 1006 : 176 - 0xb0
      13'h3EF: dout  = 8'b00111000; // 1007 :  56 - 0x38
      13'h3F0: dout  = 8'b00110001; // 1008 :  49 - 0x31 -- Sprite 0x3f
      13'h3F1: dout  = 8'b00111001; // 1009 :  57 - 0x39
      13'h3F2: dout  = 8'b00011111; // 1010 :  31 - 0x1f
      13'h3F3: dout  = 8'b00011111; // 1011 :  31 - 0x1f
      13'h3F4: dout  = 8'b00001111; // 1012 :  15 - 0xf
      13'h3F5: dout  = 8'b01011111; // 1013 :  95 - 0x5f
      13'h3F6: dout  = 8'b01111110; // 1014 : 126 - 0x7e
      13'h3F7: dout  = 8'b00111100; // 1015 :  60 - 0x3c
      13'h3F8: dout  = 8'b00011111; // 1016 :  31 - 0x1f
      13'h3F9: dout  = 8'b00000111; // 1017 :   7 - 0x7
      13'h3FA: dout  = 8'b00000000; // 1018 :   0 - 0x0
      13'h3FB: dout  = 8'b00001110; // 1019 :  14 - 0xe
      13'h3FC: dout  = 8'b00001111; // 1020 :  15 - 0xf
      13'h3FD: dout  = 8'b01010011; // 1021 :  83 - 0x53
      13'h3FE: dout  = 8'b01111100; // 1022 : 124 - 0x7c
      13'h3FF: dout  = 8'b00111100; // 1023 :  60 - 0x3c
      13'h400: dout  = 8'b11111000; // 1024 : 248 - 0xf8 -- Sprite 0x40
      13'h401: dout  = 8'b11111000; // 1025 : 248 - 0xf8
      13'h402: dout  = 8'b11110000; // 1026 : 240 - 0xf0
      13'h403: dout  = 8'b11100000; // 1027 : 224 - 0xe0
      13'h404: dout  = 8'b11100000; // 1028 : 224 - 0xe0
      13'h405: dout  = 8'b11000000; // 1029 : 192 - 0xc0
      13'h406: dout  = 8'b00000000; // 1030 :   0 - 0x0
      13'h407: dout  = 8'b00000000; // 1031 :   0 - 0x0
      13'h408: dout  = 8'b11111000; // 1032 : 248 - 0xf8
      13'h409: dout  = 8'b11111000; // 1033 : 248 - 0xf8
      13'h40A: dout  = 8'b11110000; // 1034 : 240 - 0xf0
      13'h40B: dout  = 8'b00000000; // 1035 :   0 - 0x0
      13'h40C: dout  = 8'b00000000; // 1036 :   0 - 0x0
      13'h40D: dout  = 8'b10000000; // 1037 : 128 - 0x80
      13'h40E: dout  = 8'b00000000; // 1038 :   0 - 0x0
      13'h40F: dout  = 8'b00000000; // 1039 :   0 - 0x0
      13'h410: dout  = 8'b00000000; // 1040 :   0 - 0x0 -- Sprite 0x41
      13'h411: dout  = 8'b11100000; // 1041 : 224 - 0xe0
      13'h412: dout  = 8'b11111100; // 1042 : 252 - 0xfc
      13'h413: dout  = 8'b00100111; // 1043 :  39 - 0x27
      13'h414: dout  = 8'b00100111; // 1044 :  39 - 0x27
      13'h415: dout  = 8'b00010001; // 1045 :  17 - 0x11
      13'h416: dout  = 8'b00111110; // 1046 :  62 - 0x3e
      13'h417: dout  = 8'b00000100; // 1047 :   4 - 0x4
      13'h418: dout  = 8'b00000111; // 1048 :   7 - 0x7
      13'h419: dout  = 8'b00000111; // 1049 :   7 - 0x7
      13'h41A: dout  = 8'b00000011; // 1050 :   3 - 0x3
      13'h41B: dout  = 8'b11110111; // 1051 : 247 - 0xf7
      13'h41C: dout  = 8'b11111111; // 1052 : 255 - 0xff
      13'h41D: dout  = 8'b11111111; // 1053 : 255 - 0xff
      13'h41E: dout  = 8'b11111110; // 1054 : 254 - 0xfe
      13'h41F: dout  = 8'b11111100; // 1055 : 252 - 0xfc
      13'h420: dout  = 8'b00111111; // 1056 :  63 - 0x3f -- Sprite 0x42
      13'h421: dout  = 8'b01111111; // 1057 : 127 - 0x7f
      13'h422: dout  = 8'b00111111; // 1058 :  63 - 0x3f
      13'h423: dout  = 8'b00001111; // 1059 :  15 - 0xf
      13'h424: dout  = 8'b00011111; // 1060 :  31 - 0x1f
      13'h425: dout  = 8'b00111111; // 1061 :  63 - 0x3f
      13'h426: dout  = 8'b01111111; // 1062 : 127 - 0x7f
      13'h427: dout  = 8'b01001111; // 1063 :  79 - 0x4f
      13'h428: dout  = 8'b00111110; // 1064 :  62 - 0x3e
      13'h429: dout  = 8'b01111111; // 1065 : 127 - 0x7f
      13'h42A: dout  = 8'b11111111; // 1066 : 255 - 0xff
      13'h42B: dout  = 8'b11100010; // 1067 : 226 - 0xe2
      13'h42C: dout  = 8'b01010000; // 1068 :  80 - 0x50
      13'h42D: dout  = 8'b00111000; // 1069 :  56 - 0x38
      13'h42E: dout  = 8'b01110000; // 1070 : 112 - 0x70
      13'h42F: dout  = 8'b01000000; // 1071 :  64 - 0x40
      13'h430: dout  = 8'b11111000; // 1072 : 248 - 0xf8 -- Sprite 0x43
      13'h431: dout  = 8'b11111001; // 1073 : 249 - 0xf9
      13'h432: dout  = 8'b11111001; // 1074 : 249 - 0xf9
      13'h433: dout  = 8'b10110111; // 1075 : 183 - 0xb7
      13'h434: dout  = 8'b11111111; // 1076 : 255 - 0xff
      13'h435: dout  = 8'b11111111; // 1077 : 255 - 0xff
      13'h436: dout  = 8'b11100000; // 1078 : 224 - 0xe0
      13'h437: dout  = 8'b00000000; // 1079 :   0 - 0x0
      13'h438: dout  = 8'b11101000; // 1080 : 232 - 0xe8
      13'h439: dout  = 8'b01110001; // 1081 : 113 - 0x71
      13'h43A: dout  = 8'b00000001; // 1082 :   1 - 0x1
      13'h43B: dout  = 8'b01001011; // 1083 :  75 - 0x4b
      13'h43C: dout  = 8'b00000011; // 1084 :   3 - 0x3
      13'h43D: dout  = 8'b00000011; // 1085 :   3 - 0x3
      13'h43E: dout  = 8'b00000000; // 1086 :   0 - 0x0
      13'h43F: dout  = 8'b00000000; // 1087 :   0 - 0x0
      13'h440: dout  = 8'b00000111; // 1088 :   7 - 0x7 -- Sprite 0x44
      13'h441: dout  = 8'b00000111; // 1089 :   7 - 0x7
      13'h442: dout  = 8'b00001111; // 1090 :  15 - 0xf
      13'h443: dout  = 8'b00111111; // 1091 :  63 - 0x3f
      13'h444: dout  = 8'b00111111; // 1092 :  63 - 0x3f
      13'h445: dout  = 8'b00111111; // 1093 :  63 - 0x3f
      13'h446: dout  = 8'b00100110; // 1094 :  38 - 0x26
      13'h447: dout  = 8'b00000100; // 1095 :   4 - 0x4
      13'h448: dout  = 8'b00000101; // 1096 :   5 - 0x5
      13'h449: dout  = 8'b00000011; // 1097 :   3 - 0x3
      13'h44A: dout  = 8'b00000001; // 1098 :   1 - 0x1
      13'h44B: dout  = 8'b00110000; // 1099 :  48 - 0x30
      13'h44C: dout  = 8'b00110000; // 1100 :  48 - 0x30
      13'h44D: dout  = 8'b00110000; // 1101 :  48 - 0x30
      13'h44E: dout  = 8'b00100110; // 1102 :  38 - 0x26
      13'h44F: dout  = 8'b00000100; // 1103 :   4 - 0x4
      13'h450: dout  = 8'b11110000; // 1104 : 240 - 0xf0 -- Sprite 0x45
      13'h451: dout  = 8'b11110000; // 1105 : 240 - 0xf0
      13'h452: dout  = 8'b11110000; // 1106 : 240 - 0xf0
      13'h453: dout  = 8'b11100000; // 1107 : 224 - 0xe0
      13'h454: dout  = 8'b11000000; // 1108 : 192 - 0xc0
      13'h455: dout  = 8'b00000000; // 1109 :   0 - 0x0
      13'h456: dout  = 8'b00000000; // 1110 :   0 - 0x0
      13'h457: dout  = 8'b00000000; // 1111 :   0 - 0x0
      13'h458: dout  = 8'b11111110; // 1112 : 254 - 0xfe
      13'h459: dout  = 8'b11111100; // 1113 : 252 - 0xfc
      13'h45A: dout  = 8'b11100000; // 1114 : 224 - 0xe0
      13'h45B: dout  = 8'b00000000; // 1115 :   0 - 0x0
      13'h45C: dout  = 8'b00000000; // 1116 :   0 - 0x0
      13'h45D: dout  = 8'b00000000; // 1117 :   0 - 0x0
      13'h45E: dout  = 8'b00000000; // 1118 :   0 - 0x0
      13'h45F: dout  = 8'b00000000; // 1119 :   0 - 0x0
      13'h460: dout  = 8'b00000111; // 1120 :   7 - 0x7 -- Sprite 0x46
      13'h461: dout  = 8'b00000111; // 1121 :   7 - 0x7
      13'h462: dout  = 8'b00001111; // 1122 :  15 - 0xf
      13'h463: dout  = 8'b00011111; // 1123 :  31 - 0x1f
      13'h464: dout  = 8'b00111111; // 1124 :  63 - 0x3f
      13'h465: dout  = 8'b00001111; // 1125 :  15 - 0xf
      13'h466: dout  = 8'b00011100; // 1126 :  28 - 0x1c
      13'h467: dout  = 8'b00011000; // 1127 :  24 - 0x18
      13'h468: dout  = 8'b00000101; // 1128 :   5 - 0x5
      13'h469: dout  = 8'b00000011; // 1129 :   3 - 0x3
      13'h46A: dout  = 8'b00000001; // 1130 :   1 - 0x1
      13'h46B: dout  = 8'b00010000; // 1131 :  16 - 0x10
      13'h46C: dout  = 8'b00110000; // 1132 :  48 - 0x30
      13'h46D: dout  = 8'b00001100; // 1133 :  12 - 0xc
      13'h46E: dout  = 8'b00011100; // 1134 :  28 - 0x1c
      13'h46F: dout  = 8'b00011000; // 1135 :  24 - 0x18
      13'h470: dout  = 8'b11100000; // 1136 : 224 - 0xe0 -- Sprite 0x47
      13'h471: dout  = 8'b11100000; // 1137 : 224 - 0xe0
      13'h472: dout  = 8'b11100000; // 1138 : 224 - 0xe0
      13'h473: dout  = 8'b11100000; // 1139 : 224 - 0xe0
      13'h474: dout  = 8'b11000000; // 1140 : 192 - 0xc0
      13'h475: dout  = 8'b10000000; // 1141 : 128 - 0x80
      13'h476: dout  = 8'b00000000; // 1142 :   0 - 0x0
      13'h477: dout  = 8'b00000000; // 1143 :   0 - 0x0
      13'h478: dout  = 8'b11000000; // 1144 : 192 - 0xc0
      13'h479: dout  = 8'b11100000; // 1145 : 224 - 0xe0
      13'h47A: dout  = 8'b11110000; // 1146 : 240 - 0xf0
      13'h47B: dout  = 8'b01111000; // 1147 : 120 - 0x78
      13'h47C: dout  = 8'b00011000; // 1148 :  24 - 0x18
      13'h47D: dout  = 8'b00001000; // 1149 :   8 - 0x8
      13'h47E: dout  = 8'b00000000; // 1150 :   0 - 0x0
      13'h47F: dout  = 8'b00000000; // 1151 :   0 - 0x0
      13'h480: dout  = 8'b00000111; // 1152 :   7 - 0x7 -- Sprite 0x48
      13'h481: dout  = 8'b00001111; // 1153 :  15 - 0xf
      13'h482: dout  = 8'b00011111; // 1154 :  31 - 0x1f
      13'h483: dout  = 8'b00001111; // 1155 :  15 - 0xf
      13'h484: dout  = 8'b00111111; // 1156 :  63 - 0x3f
      13'h485: dout  = 8'b00001111; // 1157 :  15 - 0xf
      13'h486: dout  = 8'b00011100; // 1158 :  28 - 0x1c
      13'h487: dout  = 8'b00011000; // 1159 :  24 - 0x18
      13'h488: dout  = 8'b00000111; // 1160 :   7 - 0x7
      13'h489: dout  = 8'b00001111; // 1161 :  15 - 0xf
      13'h48A: dout  = 8'b00111110; // 1162 :  62 - 0x3e
      13'h48B: dout  = 8'b01111100; // 1163 : 124 - 0x7c
      13'h48C: dout  = 8'b00110000; // 1164 :  48 - 0x30
      13'h48D: dout  = 8'b00001100; // 1165 :  12 - 0xc
      13'h48E: dout  = 8'b00011100; // 1166 :  28 - 0x1c
      13'h48F: dout  = 8'b00011000; // 1167 :  24 - 0x18
      13'h490: dout  = 8'b11100000; // 1168 : 224 - 0xe0 -- Sprite 0x49
      13'h491: dout  = 8'b11100000; // 1169 : 224 - 0xe0
      13'h492: dout  = 8'b11100000; // 1170 : 224 - 0xe0
      13'h493: dout  = 8'b01000000; // 1171 :  64 - 0x40
      13'h494: dout  = 8'b11000000; // 1172 : 192 - 0xc0
      13'h495: dout  = 8'b10000000; // 1173 : 128 - 0x80
      13'h496: dout  = 8'b00000000; // 1174 :   0 - 0x0
      13'h497: dout  = 8'b00000000; // 1175 :   0 - 0x0
      13'h498: dout  = 8'b01100000; // 1176 :  96 - 0x60
      13'h499: dout  = 8'b01100000; // 1177 :  96 - 0x60
      13'h49A: dout  = 8'b01100000; // 1178 :  96 - 0x60
      13'h49B: dout  = 8'b10000000; // 1179 : 128 - 0x80
      13'h49C: dout  = 8'b00000000; // 1180 :   0 - 0x0
      13'h49D: dout  = 8'b00000000; // 1181 :   0 - 0x0
      13'h49E: dout  = 8'b00000000; // 1182 :   0 - 0x0
      13'h49F: dout  = 8'b00000000; // 1183 :   0 - 0x0
      13'h4A0: dout  = 8'b01111111; // 1184 : 127 - 0x7f -- Sprite 0x4a
      13'h4A1: dout  = 8'b11111111; // 1185 : 255 - 0xff
      13'h4A2: dout  = 8'b11111111; // 1186 : 255 - 0xff
      13'h4A3: dout  = 8'b11111011; // 1187 : 251 - 0xfb
      13'h4A4: dout  = 8'b00001111; // 1188 :  15 - 0xf
      13'h4A5: dout  = 8'b00001111; // 1189 :  15 - 0xf
      13'h4A6: dout  = 8'b00001111; // 1190 :  15 - 0xf
      13'h4A7: dout  = 8'b00011111; // 1191 :  31 - 0x1f
      13'h4A8: dout  = 8'b01110011; // 1192 : 115 - 0x73
      13'h4A9: dout  = 8'b11110011; // 1193 : 243 - 0xf3
      13'h4AA: dout  = 8'b11110000; // 1194 : 240 - 0xf0
      13'h4AB: dout  = 8'b11110100; // 1195 : 244 - 0xf4
      13'h4AC: dout  = 8'b11110000; // 1196 : 240 - 0xf0
      13'h4AD: dout  = 8'b11110000; // 1197 : 240 - 0xf0
      13'h4AE: dout  = 8'b01110000; // 1198 : 112 - 0x70
      13'h4AF: dout  = 8'b01100000; // 1199 :  96 - 0x60
      13'h4B0: dout  = 8'b00111111; // 1200 :  63 - 0x3f -- Sprite 0x4b
      13'h4B1: dout  = 8'b01111110; // 1201 : 126 - 0x7e
      13'h4B2: dout  = 8'b01111100; // 1202 : 124 - 0x7c
      13'h4B3: dout  = 8'b01111100; // 1203 : 124 - 0x7c
      13'h4B4: dout  = 8'b00111100; // 1204 :  60 - 0x3c
      13'h4B5: dout  = 8'b00111100; // 1205 :  60 - 0x3c
      13'h4B6: dout  = 8'b11111100; // 1206 : 252 - 0xfc
      13'h4B7: dout  = 8'b11111100; // 1207 : 252 - 0xfc
      13'h4B8: dout  = 8'b00000000; // 1208 :   0 - 0x0
      13'h4B9: dout  = 8'b00000000; // 1209 :   0 - 0x0
      13'h4BA: dout  = 8'b00000000; // 1210 :   0 - 0x0
      13'h4BB: dout  = 8'b00000000; // 1211 :   0 - 0x0
      13'h4BC: dout  = 8'b00111100; // 1212 :  60 - 0x3c
      13'h4BD: dout  = 8'b00111100; // 1213 :  60 - 0x3c
      13'h4BE: dout  = 8'b11111100; // 1214 : 252 - 0xfc
      13'h4BF: dout  = 8'b11111100; // 1215 : 252 - 0xfc
      13'h4C0: dout  = 8'b01100000; // 1216 :  96 - 0x60 -- Sprite 0x4c
      13'h4C1: dout  = 8'b01110000; // 1217 : 112 - 0x70
      13'h4C2: dout  = 8'b00011000; // 1218 :  24 - 0x18
      13'h4C3: dout  = 8'b00001000; // 1219 :   8 - 0x8
      13'h4C4: dout  = 8'b00001111; // 1220 :  15 - 0xf
      13'h4C5: dout  = 8'b00011111; // 1221 :  31 - 0x1f
      13'h4C6: dout  = 8'b00111111; // 1222 :  63 - 0x3f
      13'h4C7: dout  = 8'b01111111; // 1223 : 127 - 0x7f
      13'h4C8: dout  = 8'b01111111; // 1224 : 127 - 0x7f
      13'h4C9: dout  = 8'b01111111; // 1225 : 127 - 0x7f
      13'h4CA: dout  = 8'b00011111; // 1226 :  31 - 0x1f
      13'h4CB: dout  = 8'b00000111; // 1227 :   7 - 0x7
      13'h4CC: dout  = 8'b00001011; // 1228 :  11 - 0xb
      13'h4CD: dout  = 8'b00011011; // 1229 :  27 - 0x1b
      13'h4CE: dout  = 8'b00111011; // 1230 :  59 - 0x3b
      13'h4CF: dout  = 8'b01111011; // 1231 : 123 - 0x7b
      13'h4D0: dout  = 8'b11111100; // 1232 : 252 - 0xfc -- Sprite 0x4d
      13'h4D1: dout  = 8'b01111100; // 1233 : 124 - 0x7c
      13'h4D2: dout  = 8'b00000000; // 1234 :   0 - 0x0
      13'h4D3: dout  = 8'b00100000; // 1235 :  32 - 0x20
      13'h4D4: dout  = 8'b11110000; // 1236 : 240 - 0xf0
      13'h4D5: dout  = 8'b11111000; // 1237 : 248 - 0xf8
      13'h4D6: dout  = 8'b11111100; // 1238 : 252 - 0xfc
      13'h4D7: dout  = 8'b11111110; // 1239 : 254 - 0xfe
      13'h4D8: dout  = 8'b11111100; // 1240 : 252 - 0xfc
      13'h4D9: dout  = 8'b11111100; // 1241 : 252 - 0xfc
      13'h4DA: dout  = 8'b11111000; // 1242 : 248 - 0xf8
      13'h4DB: dout  = 8'b11100000; // 1243 : 224 - 0xe0
      13'h4DC: dout  = 8'b11010000; // 1244 : 208 - 0xd0
      13'h4DD: dout  = 8'b11011000; // 1245 : 216 - 0xd8
      13'h4DE: dout  = 8'b11011100; // 1246 : 220 - 0xdc
      13'h4DF: dout  = 8'b11011110; // 1247 : 222 - 0xde
      13'h4E0: dout  = 8'b00001011; // 1248 :  11 - 0xb -- Sprite 0x4e
      13'h4E1: dout  = 8'b00001111; // 1249 :  15 - 0xf
      13'h4E2: dout  = 8'b00011111; // 1250 :  31 - 0x1f
      13'h4E3: dout  = 8'b00011110; // 1251 :  30 - 0x1e
      13'h4E4: dout  = 8'b00111100; // 1252 :  60 - 0x3c
      13'h4E5: dout  = 8'b00111100; // 1253 :  60 - 0x3c
      13'h4E6: dout  = 8'b00111100; // 1254 :  60 - 0x3c
      13'h4E7: dout  = 8'b01111100; // 1255 : 124 - 0x7c
      13'h4E8: dout  = 8'b11000100; // 1256 : 196 - 0xc4
      13'h4E9: dout  = 8'b11100000; // 1257 : 224 - 0xe0
      13'h4EA: dout  = 8'b11100000; // 1258 : 224 - 0xe0
      13'h4EB: dout  = 8'b01000000; // 1259 :  64 - 0x40
      13'h4EC: dout  = 8'b00000000; // 1260 :   0 - 0x0
      13'h4ED: dout  = 8'b00111100; // 1261 :  60 - 0x3c
      13'h4EE: dout  = 8'b00111100; // 1262 :  60 - 0x3c
      13'h4EF: dout  = 8'b01111100; // 1263 : 124 - 0x7c
      13'h4F0: dout  = 8'b00011111; // 1264 :  31 - 0x1f -- Sprite 0x4f
      13'h4F1: dout  = 8'b00111111; // 1265 :  63 - 0x3f
      13'h4F2: dout  = 8'b00001101; // 1266 :  13 - 0xd
      13'h4F3: dout  = 8'b00000111; // 1267 :   7 - 0x7
      13'h4F4: dout  = 8'b00001111; // 1268 :  15 - 0xf
      13'h4F5: dout  = 8'b00001110; // 1269 :  14 - 0xe
      13'h4F6: dout  = 8'b00011100; // 1270 :  28 - 0x1c
      13'h4F7: dout  = 8'b00111100; // 1271 :  60 - 0x3c
      13'h4F8: dout  = 8'b00011101; // 1272 :  29 - 0x1d
      13'h4F9: dout  = 8'b00111100; // 1273 :  60 - 0x3c
      13'h4FA: dout  = 8'b00111010; // 1274 :  58 - 0x3a
      13'h4FB: dout  = 8'b00111000; // 1275 :  56 - 0x38
      13'h4FC: dout  = 8'b00110000; // 1276 :  48 - 0x30
      13'h4FD: dout  = 8'b00000000; // 1277 :   0 - 0x0
      13'h4FE: dout  = 8'b00011100; // 1278 :  28 - 0x1c
      13'h4FF: dout  = 8'b00111100; // 1279 :  60 - 0x3c
      13'h500: dout  = 8'b00000000; // 1280 :   0 - 0x0 -- Sprite 0x50
      13'h501: dout  = 8'b00000000; // 1281 :   0 - 0x0
      13'h502: dout  = 8'b00000000; // 1282 :   0 - 0x0
      13'h503: dout  = 8'b00000000; // 1283 :   0 - 0x0
      13'h504: dout  = 8'b00000000; // 1284 :   0 - 0x0
      13'h505: dout  = 8'b00000000; // 1285 :   0 - 0x0
      13'h506: dout  = 8'b00000000; // 1286 :   0 - 0x0
      13'h507: dout  = 8'b00000000; // 1287 :   0 - 0x0
      13'h508: dout  = 8'b00100010; // 1288 :  34 - 0x22
      13'h509: dout  = 8'b01010101; // 1289 :  85 - 0x55
      13'h50A: dout  = 8'b01010101; // 1290 :  85 - 0x55
      13'h50B: dout  = 8'b01010101; // 1291 :  85 - 0x55
      13'h50C: dout  = 8'b01010101; // 1292 :  85 - 0x55
      13'h50D: dout  = 8'b01010101; // 1293 :  85 - 0x55
      13'h50E: dout  = 8'b01110111; // 1294 : 119 - 0x77
      13'h50F: dout  = 8'b00100010; // 1295 :  34 - 0x22
      13'h510: dout  = 8'b00000000; // 1296 :   0 - 0x0 -- Sprite 0x51
      13'h511: dout  = 8'b00000111; // 1297 :   7 - 0x7
      13'h512: dout  = 8'b00011111; // 1298 :  31 - 0x1f
      13'h513: dout  = 8'b11111111; // 1299 : 255 - 0xff
      13'h514: dout  = 8'b00000111; // 1300 :   7 - 0x7
      13'h515: dout  = 8'b00011111; // 1301 :  31 - 0x1f
      13'h516: dout  = 8'b00001111; // 1302 :  15 - 0xf
      13'h517: dout  = 8'b00000110; // 1303 :   6 - 0x6
      13'h518: dout  = 8'b00000000; // 1304 :   0 - 0x0
      13'h519: dout  = 8'b00000000; // 1305 :   0 - 0x0
      13'h51A: dout  = 8'b00000000; // 1306 :   0 - 0x0
      13'h51B: dout  = 8'b00000000; // 1307 :   0 - 0x0
      13'h51C: dout  = 8'b00000000; // 1308 :   0 - 0x0
      13'h51D: dout  = 8'b00000000; // 1309 :   0 - 0x0
      13'h51E: dout  = 8'b00000000; // 1310 :   0 - 0x0
      13'h51F: dout  = 8'b00000000; // 1311 :   0 - 0x0
      13'h520: dout  = 8'b00111111; // 1312 :  63 - 0x3f -- Sprite 0x52
      13'h521: dout  = 8'b11111111; // 1313 : 255 - 0xff
      13'h522: dout  = 8'b11111111; // 1314 : 255 - 0xff
      13'h523: dout  = 8'b11111111; // 1315 : 255 - 0xff
      13'h524: dout  = 8'b11111111; // 1316 : 255 - 0xff
      13'h525: dout  = 8'b11111111; // 1317 : 255 - 0xff
      13'h526: dout  = 8'b11111011; // 1318 : 251 - 0xfb
      13'h527: dout  = 8'b01110110; // 1319 : 118 - 0x76
      13'h528: dout  = 8'b00000000; // 1320 :   0 - 0x0
      13'h529: dout  = 8'b00000000; // 1321 :   0 - 0x0
      13'h52A: dout  = 8'b11001111; // 1322 : 207 - 0xcf
      13'h52B: dout  = 8'b00000111; // 1323 :   7 - 0x7
      13'h52C: dout  = 8'b01111111; // 1324 : 127 - 0x7f
      13'h52D: dout  = 8'b00000000; // 1325 :   0 - 0x0
      13'h52E: dout  = 8'b00000000; // 1326 :   0 - 0x0
      13'h52F: dout  = 8'b00000000; // 1327 :   0 - 0x0
      13'h530: dout  = 8'b00100000; // 1328 :  32 - 0x20 -- Sprite 0x53
      13'h531: dout  = 8'b11111000; // 1329 : 248 - 0xf8
      13'h532: dout  = 8'b11111111; // 1330 : 255 - 0xff
      13'h533: dout  = 8'b11000011; // 1331 : 195 - 0xc3
      13'h534: dout  = 8'b11111101; // 1332 : 253 - 0xfd
      13'h535: dout  = 8'b11111110; // 1333 : 254 - 0xfe
      13'h536: dout  = 8'b11110000; // 1334 : 240 - 0xf0
      13'h537: dout  = 8'b01000000; // 1335 :  64 - 0x40
      13'h538: dout  = 8'b00000000; // 1336 :   0 - 0x0
      13'h539: dout  = 8'b00000000; // 1337 :   0 - 0x0
      13'h53A: dout  = 8'b00111100; // 1338 :  60 - 0x3c
      13'h53B: dout  = 8'b11111100; // 1339 : 252 - 0xfc
      13'h53C: dout  = 8'b11111110; // 1340 : 254 - 0xfe
      13'h53D: dout  = 8'b11100000; // 1341 : 224 - 0xe0
      13'h53E: dout  = 8'b00000000; // 1342 :   0 - 0x0
      13'h53F: dout  = 8'b00000000; // 1343 :   0 - 0x0
      13'h540: dout  = 8'b01000000; // 1344 :  64 - 0x40 -- Sprite 0x54
      13'h541: dout  = 8'b11100000; // 1345 : 224 - 0xe0
      13'h542: dout  = 8'b01000000; // 1346 :  64 - 0x40
      13'h543: dout  = 8'b01000000; // 1347 :  64 - 0x40
      13'h544: dout  = 8'b01000001; // 1348 :  65 - 0x41
      13'h545: dout  = 8'b01000001; // 1349 :  65 - 0x41
      13'h546: dout  = 8'b01001111; // 1350 :  79 - 0x4f
      13'h547: dout  = 8'b01000111; // 1351 :  71 - 0x47
      13'h548: dout  = 8'b01000000; // 1352 :  64 - 0x40
      13'h549: dout  = 8'b11100000; // 1353 : 224 - 0xe0
      13'h54A: dout  = 8'b01000000; // 1354 :  64 - 0x40
      13'h54B: dout  = 8'b00111111; // 1355 :  63 - 0x3f
      13'h54C: dout  = 8'b00111110; // 1356 :  62 - 0x3e
      13'h54D: dout  = 8'b00111110; // 1357 :  62 - 0x3e
      13'h54E: dout  = 8'b00110000; // 1358 :  48 - 0x30
      13'h54F: dout  = 8'b00111000; // 1359 :  56 - 0x38
      13'h550: dout  = 8'b00000000; // 1360 :   0 - 0x0 -- Sprite 0x55
      13'h551: dout  = 8'b00000000; // 1361 :   0 - 0x0
      13'h552: dout  = 8'b00000000; // 1362 :   0 - 0x0
      13'h553: dout  = 8'b00000000; // 1363 :   0 - 0x0
      13'h554: dout  = 8'b00000000; // 1364 :   0 - 0x0
      13'h555: dout  = 8'b00000000; // 1365 :   0 - 0x0
      13'h556: dout  = 8'b11100000; // 1366 : 224 - 0xe0
      13'h557: dout  = 8'b11000000; // 1367 : 192 - 0xc0
      13'h558: dout  = 8'b00000000; // 1368 :   0 - 0x0
      13'h559: dout  = 8'b00000000; // 1369 :   0 - 0x0
      13'h55A: dout  = 8'b00000000; // 1370 :   0 - 0x0
      13'h55B: dout  = 8'b11111000; // 1371 : 248 - 0xf8
      13'h55C: dout  = 8'b11111000; // 1372 : 248 - 0xf8
      13'h55D: dout  = 8'b11111000; // 1373 : 248 - 0xf8
      13'h55E: dout  = 8'b00011000; // 1374 :  24 - 0x18
      13'h55F: dout  = 8'b00111000; // 1375 :  56 - 0x38
      13'h560: dout  = 8'b01000011; // 1376 :  67 - 0x43 -- Sprite 0x56
      13'h561: dout  = 8'b01000110; // 1377 :  70 - 0x46
      13'h562: dout  = 8'b01000100; // 1378 :  68 - 0x44
      13'h563: dout  = 8'b01000000; // 1379 :  64 - 0x40
      13'h564: dout  = 8'b01000000; // 1380 :  64 - 0x40
      13'h565: dout  = 8'b01000000; // 1381 :  64 - 0x40
      13'h566: dout  = 8'b01000000; // 1382 :  64 - 0x40
      13'h567: dout  = 8'b01000000; // 1383 :  64 - 0x40
      13'h568: dout  = 8'b00111100; // 1384 :  60 - 0x3c
      13'h569: dout  = 8'b00111001; // 1385 :  57 - 0x39
      13'h56A: dout  = 8'b00111011; // 1386 :  59 - 0x3b
      13'h56B: dout  = 8'b00111111; // 1387 :  63 - 0x3f
      13'h56C: dout  = 8'b00000000; // 1388 :   0 - 0x0
      13'h56D: dout  = 8'b00000000; // 1389 :   0 - 0x0
      13'h56E: dout  = 8'b00000000; // 1390 :   0 - 0x0
      13'h56F: dout  = 8'b00000000; // 1391 :   0 - 0x0
      13'h570: dout  = 8'b10000000; // 1392 : 128 - 0x80 -- Sprite 0x57
      13'h571: dout  = 8'b11000000; // 1393 : 192 - 0xc0
      13'h572: dout  = 8'b01000000; // 1394 :  64 - 0x40
      13'h573: dout  = 8'b00000000; // 1395 :   0 - 0x0
      13'h574: dout  = 8'b00000000; // 1396 :   0 - 0x0
      13'h575: dout  = 8'b00000000; // 1397 :   0 - 0x0
      13'h576: dout  = 8'b00000000; // 1398 :   0 - 0x0
      13'h577: dout  = 8'b00000000; // 1399 :   0 - 0x0
      13'h578: dout  = 8'b01111000; // 1400 : 120 - 0x78
      13'h579: dout  = 8'b00111000; // 1401 :  56 - 0x38
      13'h57A: dout  = 8'b10111000; // 1402 : 184 - 0xb8
      13'h57B: dout  = 8'b11111000; // 1403 : 248 - 0xf8
      13'h57C: dout  = 8'b00000000; // 1404 :   0 - 0x0
      13'h57D: dout  = 8'b00000000; // 1405 :   0 - 0x0
      13'h57E: dout  = 8'b00000000; // 1406 :   0 - 0x0
      13'h57F: dout  = 8'b00000000; // 1407 :   0 - 0x0
      13'h580: dout  = 8'b00110001; // 1408 :  49 - 0x31 -- Sprite 0x58
      13'h581: dout  = 8'b00110000; // 1409 :  48 - 0x30
      13'h582: dout  = 8'b00111000; // 1410 :  56 - 0x38
      13'h583: dout  = 8'b01111100; // 1411 : 124 - 0x7c
      13'h584: dout  = 8'b01111111; // 1412 : 127 - 0x7f
      13'h585: dout  = 8'b11111111; // 1413 : 255 - 0xff
      13'h586: dout  = 8'b11111111; // 1414 : 255 - 0xff
      13'h587: dout  = 8'b11111011; // 1415 : 251 - 0xfb
      13'h588: dout  = 8'b00111111; // 1416 :  63 - 0x3f
      13'h589: dout  = 8'b00111111; // 1417 :  63 - 0x3f
      13'h58A: dout  = 8'b00001111; // 1418 :  15 - 0xf
      13'h58B: dout  = 8'b01110111; // 1419 : 119 - 0x77
      13'h58C: dout  = 8'b01110111; // 1420 : 119 - 0x77
      13'h58D: dout  = 8'b11110111; // 1421 : 247 - 0xf7
      13'h58E: dout  = 8'b11110111; // 1422 : 247 - 0xf7
      13'h58F: dout  = 8'b11110111; // 1423 : 247 - 0xf7
      13'h590: dout  = 8'b00010000; // 1424 :  16 - 0x10 -- Sprite 0x59
      13'h591: dout  = 8'b01111110; // 1425 : 126 - 0x7e
      13'h592: dout  = 8'b00111110; // 1426 :  62 - 0x3e
      13'h593: dout  = 8'b00000000; // 1427 :   0 - 0x0
      13'h594: dout  = 8'b00011110; // 1428 :  30 - 0x1e
      13'h595: dout  = 8'b11111110; // 1429 : 254 - 0xfe
      13'h596: dout  = 8'b11111111; // 1430 : 255 - 0xff
      13'h597: dout  = 8'b11111111; // 1431 : 255 - 0xff
      13'h598: dout  = 8'b11111111; // 1432 : 255 - 0xff
      13'h599: dout  = 8'b11111110; // 1433 : 254 - 0xfe
      13'h59A: dout  = 8'b11111110; // 1434 : 254 - 0xfe
      13'h59B: dout  = 8'b11111110; // 1435 : 254 - 0xfe
      13'h59C: dout  = 8'b11111010; // 1436 : 250 - 0xfa
      13'h59D: dout  = 8'b11111010; // 1437 : 250 - 0xfa
      13'h59E: dout  = 8'b11110011; // 1438 : 243 - 0xf3
      13'h59F: dout  = 8'b11100111; // 1439 : 231 - 0xe7
      13'h5A0: dout  = 8'b11111111; // 1440 : 255 - 0xff -- Sprite 0x5a
      13'h5A1: dout  = 8'b11111111; // 1441 : 255 - 0xff
      13'h5A2: dout  = 8'b11100011; // 1442 : 227 - 0xe3
      13'h5A3: dout  = 8'b11000011; // 1443 : 195 - 0xc3
      13'h5A4: dout  = 8'b10000111; // 1444 : 135 - 0x87
      13'h5A5: dout  = 8'b01001000; // 1445 :  72 - 0x48
      13'h5A6: dout  = 8'b00111100; // 1446 :  60 - 0x3c
      13'h5A7: dout  = 8'b11111100; // 1447 : 252 - 0xfc
      13'h5A8: dout  = 8'b11110000; // 1448 : 240 - 0xf0
      13'h5A9: dout  = 8'b11111000; // 1449 : 248 - 0xf8
      13'h5AA: dout  = 8'b11111100; // 1450 : 252 - 0xfc
      13'h5AB: dout  = 8'b01111100; // 1451 : 124 - 0x7c
      13'h5AC: dout  = 8'b01111000; // 1452 : 120 - 0x78
      13'h5AD: dout  = 8'b00111000; // 1453 :  56 - 0x38
      13'h5AE: dout  = 8'b00111100; // 1454 :  60 - 0x3c
      13'h5AF: dout  = 8'b11111100; // 1455 : 252 - 0xfc
      13'h5B0: dout  = 8'b00000000; // 1456 :   0 - 0x0 -- Sprite 0x5b
      13'h5B1: dout  = 8'b11111111; // 1457 : 255 - 0xff
      13'h5B2: dout  = 8'b11000011; // 1458 : 195 - 0xc3
      13'h5B3: dout  = 8'b10000011; // 1459 : 131 - 0x83
      13'h5B4: dout  = 8'b10000011; // 1460 : 131 - 0x83
      13'h5B5: dout  = 8'b11111111; // 1461 : 255 - 0xff
      13'h5B6: dout  = 8'b11111111; // 1462 : 255 - 0xff
      13'h5B7: dout  = 8'b11111111; // 1463 : 255 - 0xff
      13'h5B8: dout  = 8'b11111111; // 1464 : 255 - 0xff
      13'h5B9: dout  = 8'b00000000; // 1465 :   0 - 0x0
      13'h5BA: dout  = 8'b11000011; // 1466 : 195 - 0xc3
      13'h5BB: dout  = 8'b10000001; // 1467 : 129 - 0x81
      13'h5BC: dout  = 8'b10000001; // 1468 : 129 - 0x81
      13'h5BD: dout  = 8'b11000011; // 1469 : 195 - 0xc3
      13'h5BE: dout  = 8'b11111111; // 1470 : 255 - 0xff
      13'h5BF: dout  = 8'b00000000; // 1471 :   0 - 0x0
      13'h5C0: dout  = 8'b00011111; // 1472 :  31 - 0x1f -- Sprite 0x5c
      13'h5C1: dout  = 8'b00011111; // 1473 :  31 - 0x1f
      13'h5C2: dout  = 8'b00001111; // 1474 :  15 - 0xf
      13'h5C3: dout  = 8'b00000111; // 1475 :   7 - 0x7
      13'h5C4: dout  = 8'b00000001; // 1476 :   1 - 0x1
      13'h5C5: dout  = 8'b00000000; // 1477 :   0 - 0x0
      13'h5C6: dout  = 8'b00000000; // 1478 :   0 - 0x0
      13'h5C7: dout  = 8'b00000000; // 1479 :   0 - 0x0
      13'h5C8: dout  = 8'b00000000; // 1480 :   0 - 0x0
      13'h5C9: dout  = 8'b00000000; // 1481 :   0 - 0x0
      13'h5CA: dout  = 8'b00000000; // 1482 :   0 - 0x0
      13'h5CB: dout  = 8'b00000000; // 1483 :   0 - 0x0
      13'h5CC: dout  = 8'b00000000; // 1484 :   0 - 0x0
      13'h5CD: dout  = 8'b00000000; // 1485 :   0 - 0x0
      13'h5CE: dout  = 8'b00000000; // 1486 :   0 - 0x0
      13'h5CF: dout  = 8'b00000000; // 1487 :   0 - 0x0
      13'h5D0: dout  = 8'b11110000; // 1488 : 240 - 0xf0 -- Sprite 0x5d
      13'h5D1: dout  = 8'b11111011; // 1489 : 251 - 0xfb
      13'h5D2: dout  = 8'b11111111; // 1490 : 255 - 0xff
      13'h5D3: dout  = 8'b11111111; // 1491 : 255 - 0xff
      13'h5D4: dout  = 8'b11111110; // 1492 : 254 - 0xfe
      13'h5D5: dout  = 8'b00111110; // 1493 :  62 - 0x3e
      13'h5D6: dout  = 8'b00001100; // 1494 :  12 - 0xc
      13'h5D7: dout  = 8'b00000100; // 1495 :   4 - 0x4
      13'h5D8: dout  = 8'b00000000; // 1496 :   0 - 0x0
      13'h5D9: dout  = 8'b00001011; // 1497 :  11 - 0xb
      13'h5DA: dout  = 8'b00011111; // 1498 :  31 - 0x1f
      13'h5DB: dout  = 8'b00011111; // 1499 :  31 - 0x1f
      13'h5DC: dout  = 8'b00011110; // 1500 :  30 - 0x1e
      13'h5DD: dout  = 8'b00111110; // 1501 :  62 - 0x3e
      13'h5DE: dout  = 8'b00001100; // 1502 :  12 - 0xc
      13'h5DF: dout  = 8'b00000100; // 1503 :   4 - 0x4
      13'h5E0: dout  = 8'b00011111; // 1504 :  31 - 0x1f -- Sprite 0x5e
      13'h5E1: dout  = 8'b00011111; // 1505 :  31 - 0x1f
      13'h5E2: dout  = 8'b00001111; // 1506 :  15 - 0xf
      13'h5E3: dout  = 8'b00001111; // 1507 :  15 - 0xf
      13'h5E4: dout  = 8'b00000111; // 1508 :   7 - 0x7
      13'h5E5: dout  = 8'b00000000; // 1509 :   0 - 0x0
      13'h5E6: dout  = 8'b00000000; // 1510 :   0 - 0x0
      13'h5E7: dout  = 8'b00000000; // 1511 :   0 - 0x0
      13'h5E8: dout  = 8'b00000000; // 1512 :   0 - 0x0
      13'h5E9: dout  = 8'b00000000; // 1513 :   0 - 0x0
      13'h5EA: dout  = 8'b00000000; // 1514 :   0 - 0x0
      13'h5EB: dout  = 8'b00000000; // 1515 :   0 - 0x0
      13'h5EC: dout  = 8'b00000000; // 1516 :   0 - 0x0
      13'h5ED: dout  = 8'b00000000; // 1517 :   0 - 0x0
      13'h5EE: dout  = 8'b00000000; // 1518 :   0 - 0x0
      13'h5EF: dout  = 8'b00000000; // 1519 :   0 - 0x0
      13'h5F0: dout  = 8'b11111011; // 1520 : 251 - 0xfb -- Sprite 0x5f
      13'h5F1: dout  = 8'b11111111; // 1521 : 255 - 0xff
      13'h5F2: dout  = 8'b11111111; // 1522 : 255 - 0xff
      13'h5F3: dout  = 8'b11111111; // 1523 : 255 - 0xff
      13'h5F4: dout  = 8'b11111111; // 1524 : 255 - 0xff
      13'h5F5: dout  = 8'b00000000; // 1525 :   0 - 0x0
      13'h5F6: dout  = 8'b00000000; // 1526 :   0 - 0x0
      13'h5F7: dout  = 8'b00000000; // 1527 :   0 - 0x0
      13'h5F8: dout  = 8'b00000011; // 1528 :   3 - 0x3
      13'h5F9: dout  = 8'b00001111; // 1529 :  15 - 0xf
      13'h5FA: dout  = 8'b00001111; // 1530 :  15 - 0xf
      13'h5FB: dout  = 8'b00001111; // 1531 :  15 - 0xf
      13'h5FC: dout  = 8'b00001111; // 1532 :  15 - 0xf
      13'h5FD: dout  = 8'b00000000; // 1533 :   0 - 0x0
      13'h5FE: dout  = 8'b00000000; // 1534 :   0 - 0x0
      13'h5FF: dout  = 8'b00000000; // 1535 :   0 - 0x0
      13'h600: dout  = 8'b00000000; // 1536 :   0 - 0x0 -- Sprite 0x60
      13'h601: dout  = 8'b00011000; // 1537 :  24 - 0x18
      13'h602: dout  = 8'b00111100; // 1538 :  60 - 0x3c
      13'h603: dout  = 8'b01111110; // 1539 : 126 - 0x7e
      13'h604: dout  = 8'b01101110; // 1540 : 110 - 0x6e
      13'h605: dout  = 8'b11011111; // 1541 : 223 - 0xdf
      13'h606: dout  = 8'b11011111; // 1542 : 223 - 0xdf
      13'h607: dout  = 8'b11011111; // 1543 : 223 - 0xdf
      13'h608: dout  = 8'b00000000; // 1544 :   0 - 0x0
      13'h609: dout  = 8'b00011000; // 1545 :  24 - 0x18
      13'h60A: dout  = 8'b00111100; // 1546 :  60 - 0x3c
      13'h60B: dout  = 8'b01111110; // 1547 : 126 - 0x7e
      13'h60C: dout  = 8'b01110110; // 1548 : 118 - 0x76
      13'h60D: dout  = 8'b11111011; // 1549 : 251 - 0xfb
      13'h60E: dout  = 8'b11111011; // 1550 : 251 - 0xfb
      13'h60F: dout  = 8'b11111011; // 1551 : 251 - 0xfb
      13'h610: dout  = 8'b00000000; // 1552 :   0 - 0x0 -- Sprite 0x61
      13'h611: dout  = 8'b00011000; // 1553 :  24 - 0x18
      13'h612: dout  = 8'b00011000; // 1554 :  24 - 0x18
      13'h613: dout  = 8'b00111100; // 1555 :  60 - 0x3c
      13'h614: dout  = 8'b00111100; // 1556 :  60 - 0x3c
      13'h615: dout  = 8'b00111100; // 1557 :  60 - 0x3c
      13'h616: dout  = 8'b00111100; // 1558 :  60 - 0x3c
      13'h617: dout  = 8'b00011100; // 1559 :  28 - 0x1c
      13'h618: dout  = 8'b00000000; // 1560 :   0 - 0x0
      13'h619: dout  = 8'b00010000; // 1561 :  16 - 0x10
      13'h61A: dout  = 8'b00010000; // 1562 :  16 - 0x10
      13'h61B: dout  = 8'b00100000; // 1563 :  32 - 0x20
      13'h61C: dout  = 8'b00100000; // 1564 :  32 - 0x20
      13'h61D: dout  = 8'b00100000; // 1565 :  32 - 0x20
      13'h61E: dout  = 8'b00100000; // 1566 :  32 - 0x20
      13'h61F: dout  = 8'b00100000; // 1567 :  32 - 0x20
      13'h620: dout  = 8'b00000000; // 1568 :   0 - 0x0 -- Sprite 0x62
      13'h621: dout  = 8'b00001000; // 1569 :   8 - 0x8
      13'h622: dout  = 8'b00001000; // 1570 :   8 - 0x8
      13'h623: dout  = 8'b00001000; // 1571 :   8 - 0x8
      13'h624: dout  = 8'b00001000; // 1572 :   8 - 0x8
      13'h625: dout  = 8'b00001000; // 1573 :   8 - 0x8
      13'h626: dout  = 8'b00001000; // 1574 :   8 - 0x8
      13'h627: dout  = 8'b00000000; // 1575 :   0 - 0x0
      13'h628: dout  = 8'b00000000; // 1576 :   0 - 0x0
      13'h629: dout  = 8'b00001000; // 1577 :   8 - 0x8
      13'h62A: dout  = 8'b00001000; // 1578 :   8 - 0x8
      13'h62B: dout  = 8'b00001000; // 1579 :   8 - 0x8
      13'h62C: dout  = 8'b00001000; // 1580 :   8 - 0x8
      13'h62D: dout  = 8'b00001000; // 1581 :   8 - 0x8
      13'h62E: dout  = 8'b00001000; // 1582 :   8 - 0x8
      13'h62F: dout  = 8'b00001000; // 1583 :   8 - 0x8
      13'h630: dout  = 8'b00000000; // 1584 :   0 - 0x0 -- Sprite 0x63
      13'h631: dout  = 8'b00001000; // 1585 :   8 - 0x8
      13'h632: dout  = 8'b00001000; // 1586 :   8 - 0x8
      13'h633: dout  = 8'b00000100; // 1587 :   4 - 0x4
      13'h634: dout  = 8'b00000100; // 1588 :   4 - 0x4
      13'h635: dout  = 8'b00000100; // 1589 :   4 - 0x4
      13'h636: dout  = 8'b00000100; // 1590 :   4 - 0x4
      13'h637: dout  = 8'b00000100; // 1591 :   4 - 0x4
      13'h638: dout  = 8'b00000000; // 1592 :   0 - 0x0
      13'h639: dout  = 8'b00010000; // 1593 :  16 - 0x10
      13'h63A: dout  = 8'b00010000; // 1594 :  16 - 0x10
      13'h63B: dout  = 8'b00111000; // 1595 :  56 - 0x38
      13'h63C: dout  = 8'b00111000; // 1596 :  56 - 0x38
      13'h63D: dout  = 8'b00111000; // 1597 :  56 - 0x38
      13'h63E: dout  = 8'b00111000; // 1598 :  56 - 0x38
      13'h63F: dout  = 8'b00111000; // 1599 :  56 - 0x38
      13'h640: dout  = 8'b00111100; // 1600 :  60 - 0x3c -- Sprite 0x64
      13'h641: dout  = 8'b01111110; // 1601 : 126 - 0x7e
      13'h642: dout  = 8'b01110111; // 1602 : 119 - 0x77
      13'h643: dout  = 8'b11111011; // 1603 : 251 - 0xfb
      13'h644: dout  = 8'b10011111; // 1604 : 159 - 0x9f
      13'h645: dout  = 8'b01011111; // 1605 :  95 - 0x5f
      13'h646: dout  = 8'b10001110; // 1606 : 142 - 0x8e
      13'h647: dout  = 8'b00100000; // 1607 :  32 - 0x20
      13'h648: dout  = 8'b00000000; // 1608 :   0 - 0x0
      13'h649: dout  = 8'b00011000; // 1609 :  24 - 0x18
      13'h64A: dout  = 8'b00111100; // 1610 :  60 - 0x3c
      13'h64B: dout  = 8'b00001110; // 1611 :  14 - 0xe
      13'h64C: dout  = 8'b00001110; // 1612 :  14 - 0xe
      13'h64D: dout  = 8'b00000100; // 1613 :   4 - 0x4
      13'h64E: dout  = 8'b00000000; // 1614 :   0 - 0x0
      13'h64F: dout  = 8'b00000000; // 1615 :   0 - 0x0
      13'h650: dout  = 8'b01011100; // 1616 :  92 - 0x5c -- Sprite 0x65
      13'h651: dout  = 8'b00101110; // 1617 :  46 - 0x2e
      13'h652: dout  = 8'b10001111; // 1618 : 143 - 0x8f
      13'h653: dout  = 8'b00111111; // 1619 :  63 - 0x3f
      13'h654: dout  = 8'b01111011; // 1620 : 123 - 0x7b
      13'h655: dout  = 8'b01110111; // 1621 : 119 - 0x77
      13'h656: dout  = 8'b01111110; // 1622 : 126 - 0x7e
      13'h657: dout  = 8'b00111100; // 1623 :  60 - 0x3c
      13'h658: dout  = 8'b00000000; // 1624 :   0 - 0x0
      13'h659: dout  = 8'b00000000; // 1625 :   0 - 0x0
      13'h65A: dout  = 8'b00000100; // 1626 :   4 - 0x4
      13'h65B: dout  = 8'b00000110; // 1627 :   6 - 0x6
      13'h65C: dout  = 8'b00011110; // 1628 :  30 - 0x1e
      13'h65D: dout  = 8'b00111100; // 1629 :  60 - 0x3c
      13'h65E: dout  = 8'b00011000; // 1630 :  24 - 0x18
      13'h65F: dout  = 8'b00000000; // 1631 :   0 - 0x0
      13'h660: dout  = 8'b00010011; // 1632 :  19 - 0x13 -- Sprite 0x66
      13'h661: dout  = 8'b01001111; // 1633 :  79 - 0x4f
      13'h662: dout  = 8'b00111111; // 1634 :  63 - 0x3f
      13'h663: dout  = 8'b10111111; // 1635 : 191 - 0xbf
      13'h664: dout  = 8'b00111111; // 1636 :  63 - 0x3f
      13'h665: dout  = 8'b01111010; // 1637 : 122 - 0x7a
      13'h666: dout  = 8'b11111000; // 1638 : 248 - 0xf8
      13'h667: dout  = 8'b11111000; // 1639 : 248 - 0xf8
      13'h668: dout  = 8'b00000000; // 1640 :   0 - 0x0
      13'h669: dout  = 8'b00000000; // 1641 :   0 - 0x0
      13'h66A: dout  = 8'b00000001; // 1642 :   1 - 0x1
      13'h66B: dout  = 8'b00001010; // 1643 :  10 - 0xa
      13'h66C: dout  = 8'b00010111; // 1644 :  23 - 0x17
      13'h66D: dout  = 8'b00001111; // 1645 :  15 - 0xf
      13'h66E: dout  = 8'b00101111; // 1646 :  47 - 0x2f
      13'h66F: dout  = 8'b00011111; // 1647 :  31 - 0x1f
      13'h670: dout  = 8'b00000000; // 1648 :   0 - 0x0 -- Sprite 0x67
      13'h671: dout  = 8'b00001000; // 1649 :   8 - 0x8
      13'h672: dout  = 8'b00000101; // 1650 :   5 - 0x5
      13'h673: dout  = 8'b00001111; // 1651 :  15 - 0xf
      13'h674: dout  = 8'b00101111; // 1652 :  47 - 0x2f
      13'h675: dout  = 8'b00011101; // 1653 :  29 - 0x1d
      13'h676: dout  = 8'b00011100; // 1654 :  28 - 0x1c
      13'h677: dout  = 8'b00111100; // 1655 :  60 - 0x3c
      13'h678: dout  = 8'b00000000; // 1656 :   0 - 0x0
      13'h679: dout  = 8'b00000000; // 1657 :   0 - 0x0
      13'h67A: dout  = 8'b00000000; // 1658 :   0 - 0x0
      13'h67B: dout  = 8'b00000000; // 1659 :   0 - 0x0
      13'h67C: dout  = 8'b00000101; // 1660 :   5 - 0x5
      13'h67D: dout  = 8'b00000111; // 1661 :   7 - 0x7
      13'h67E: dout  = 8'b00001111; // 1662 :  15 - 0xf
      13'h67F: dout  = 8'b00000111; // 1663 :   7 - 0x7
      13'h680: dout  = 8'b00000000; // 1664 :   0 - 0x0 -- Sprite 0x68
      13'h681: dout  = 8'b00000000; // 1665 :   0 - 0x0
      13'h682: dout  = 8'b00000000; // 1666 :   0 - 0x0
      13'h683: dout  = 8'b00000000; // 1667 :   0 - 0x0
      13'h684: dout  = 8'b00000010; // 1668 :   2 - 0x2
      13'h685: dout  = 8'b00001011; // 1669 :  11 - 0xb
      13'h686: dout  = 8'b00000111; // 1670 :   7 - 0x7
      13'h687: dout  = 8'b00001111; // 1671 :  15 - 0xf
      13'h688: dout  = 8'b00000000; // 1672 :   0 - 0x0
      13'h689: dout  = 8'b00000000; // 1673 :   0 - 0x0
      13'h68A: dout  = 8'b00000000; // 1674 :   0 - 0x0
      13'h68B: dout  = 8'b00000000; // 1675 :   0 - 0x0
      13'h68C: dout  = 8'b00000000; // 1676 :   0 - 0x0
      13'h68D: dout  = 8'b00000000; // 1677 :   0 - 0x0
      13'h68E: dout  = 8'b00000001; // 1678 :   1 - 0x1
      13'h68F: dout  = 8'b00000011; // 1679 :   3 - 0x3
      13'h690: dout  = 8'b00000000; // 1680 :   0 - 0x0 -- Sprite 0x69
      13'h691: dout  = 8'b00000000; // 1681 :   0 - 0x0
      13'h692: dout  = 8'b00000000; // 1682 :   0 - 0x0
      13'h693: dout  = 8'b00000000; // 1683 :   0 - 0x0
      13'h694: dout  = 8'b00000000; // 1684 :   0 - 0x0
      13'h695: dout  = 8'b00001000; // 1685 :   8 - 0x8
      13'h696: dout  = 8'b00000100; // 1686 :   4 - 0x4
      13'h697: dout  = 8'b00000100; // 1687 :   4 - 0x4
      13'h698: dout  = 8'b00000000; // 1688 :   0 - 0x0
      13'h699: dout  = 8'b01100000; // 1689 :  96 - 0x60
      13'h69A: dout  = 8'b11110000; // 1690 : 240 - 0xf0
      13'h69B: dout  = 8'b11111000; // 1691 : 248 - 0xf8
      13'h69C: dout  = 8'b01111100; // 1692 : 124 - 0x7c
      13'h69D: dout  = 8'b00111110; // 1693 :  62 - 0x3e
      13'h69E: dout  = 8'b01111110; // 1694 : 126 - 0x7e
      13'h69F: dout  = 8'b01111111; // 1695 : 127 - 0x7f
      13'h6A0: dout  = 8'b00000010; // 1696 :   2 - 0x2 -- Sprite 0x6a
      13'h6A1: dout  = 8'b00000010; // 1697 :   2 - 0x2
      13'h6A2: dout  = 8'b00000010; // 1698 :   2 - 0x2
      13'h6A3: dout  = 8'b00000101; // 1699 :   5 - 0x5
      13'h6A4: dout  = 8'b01110001; // 1700 : 113 - 0x71
      13'h6A5: dout  = 8'b01111111; // 1701 : 127 - 0x7f
      13'h6A6: dout  = 8'b01111111; // 1702 : 127 - 0x7f
      13'h6A7: dout  = 8'b01111111; // 1703 : 127 - 0x7f
      13'h6A8: dout  = 8'b00111111; // 1704 :  63 - 0x3f
      13'h6A9: dout  = 8'b01011111; // 1705 :  95 - 0x5f
      13'h6AA: dout  = 8'b01111111; // 1706 : 127 - 0x7f
      13'h6AB: dout  = 8'b00111110; // 1707 :  62 - 0x3e
      13'h6AC: dout  = 8'b00001110; // 1708 :  14 - 0xe
      13'h6AD: dout  = 8'b00001010; // 1709 :  10 - 0xa
      13'h6AE: dout  = 8'b01010001; // 1710 :  81 - 0x51
      13'h6AF: dout  = 8'b00100000; // 1711 :  32 - 0x20
      13'h6B0: dout  = 8'b00000000; // 1712 :   0 - 0x0 -- Sprite 0x6b
      13'h6B1: dout  = 8'b00000000; // 1713 :   0 - 0x0
      13'h6B2: dout  = 8'b00000000; // 1714 :   0 - 0x0
      13'h6B3: dout  = 8'b00000000; // 1715 :   0 - 0x0
      13'h6B4: dout  = 8'b00000000; // 1716 :   0 - 0x0
      13'h6B5: dout  = 8'b00000000; // 1717 :   0 - 0x0
      13'h6B6: dout  = 8'b00000000; // 1718 :   0 - 0x0
      13'h6B7: dout  = 8'b00000100; // 1719 :   4 - 0x4
      13'h6B8: dout  = 8'b00000000; // 1720 :   0 - 0x0
      13'h6B9: dout  = 8'b00000000; // 1721 :   0 - 0x0
      13'h6BA: dout  = 8'b00000000; // 1722 :   0 - 0x0
      13'h6BB: dout  = 8'b00000000; // 1723 :   0 - 0x0
      13'h6BC: dout  = 8'b00000000; // 1724 :   0 - 0x0
      13'h6BD: dout  = 8'b00000000; // 1725 :   0 - 0x0
      13'h6BE: dout  = 8'b00001110; // 1726 :  14 - 0xe
      13'h6BF: dout  = 8'b00011111; // 1727 :  31 - 0x1f
      13'h6C0: dout  = 8'b00000010; // 1728 :   2 - 0x2 -- Sprite 0x6c
      13'h6C1: dout  = 8'b00000010; // 1729 :   2 - 0x2
      13'h6C2: dout  = 8'b00000000; // 1730 :   0 - 0x0
      13'h6C3: dout  = 8'b00000001; // 1731 :   1 - 0x1
      13'h6C4: dout  = 8'b00010011; // 1732 :  19 - 0x13
      13'h6C5: dout  = 8'b00111111; // 1733 :  63 - 0x3f
      13'h6C6: dout  = 8'b01111111; // 1734 : 127 - 0x7f
      13'h6C7: dout  = 8'b01111111; // 1735 : 127 - 0x7f
      13'h6C8: dout  = 8'b00111111; // 1736 :  63 - 0x3f
      13'h6C9: dout  = 8'b01111111; // 1737 : 127 - 0x7f
      13'h6CA: dout  = 8'b01111111; // 1738 : 127 - 0x7f
      13'h6CB: dout  = 8'b11111110; // 1739 : 254 - 0xfe
      13'h6CC: dout  = 8'b11101100; // 1740 : 236 - 0xec
      13'h6CD: dout  = 8'b11001010; // 1741 : 202 - 0xca
      13'h6CE: dout  = 8'b01010001; // 1742 :  81 - 0x51
      13'h6CF: dout  = 8'b00100000; // 1743 :  32 - 0x20
      13'h6D0: dout  = 8'b00000000; // 1744 :   0 - 0x0 -- Sprite 0x6d
      13'h6D1: dout  = 8'b01000000; // 1745 :  64 - 0x40
      13'h6D2: dout  = 8'b01100000; // 1746 :  96 - 0x60
      13'h6D3: dout  = 8'b01110000; // 1747 : 112 - 0x70
      13'h6D4: dout  = 8'b01110011; // 1748 : 115 - 0x73
      13'h6D5: dout  = 8'b00100111; // 1749 :  39 - 0x27
      13'h6D6: dout  = 8'b00001111; // 1750 :  15 - 0xf
      13'h6D7: dout  = 8'b00011111; // 1751 :  31 - 0x1f
      13'h6D8: dout  = 8'b00000000; // 1752 :   0 - 0x0
      13'h6D9: dout  = 8'b01000000; // 1753 :  64 - 0x40
      13'h6DA: dout  = 8'b01100011; // 1754 :  99 - 0x63
      13'h6DB: dout  = 8'b01110111; // 1755 : 119 - 0x77
      13'h6DC: dout  = 8'b01111100; // 1756 : 124 - 0x7c
      13'h6DD: dout  = 8'b00111000; // 1757 :  56 - 0x38
      13'h6DE: dout  = 8'b11111000; // 1758 : 248 - 0xf8
      13'h6DF: dout  = 8'b11100100; // 1759 : 228 - 0xe4
      13'h6E0: dout  = 8'b00000000; // 1760 :   0 - 0x0 -- Sprite 0x6e
      13'h6E1: dout  = 8'b00000000; // 1761 :   0 - 0x0
      13'h6E2: dout  = 8'b00000000; // 1762 :   0 - 0x0
      13'h6E3: dout  = 8'b00000000; // 1763 :   0 - 0x0
      13'h6E4: dout  = 8'b00000011; // 1764 :   3 - 0x3
      13'h6E5: dout  = 8'b00000111; // 1765 :   7 - 0x7
      13'h6E6: dout  = 8'b00001111; // 1766 :  15 - 0xf
      13'h6E7: dout  = 8'b00011111; // 1767 :  31 - 0x1f
      13'h6E8: dout  = 8'b00000000; // 1768 :   0 - 0x0
      13'h6E9: dout  = 8'b00000000; // 1769 :   0 - 0x0
      13'h6EA: dout  = 8'b00000011; // 1770 :   3 - 0x3
      13'h6EB: dout  = 8'b00000111; // 1771 :   7 - 0x7
      13'h6EC: dout  = 8'b00001100; // 1772 :  12 - 0xc
      13'h6ED: dout  = 8'b00011000; // 1773 :  24 - 0x18
      13'h6EE: dout  = 8'b11111000; // 1774 : 248 - 0xf8
      13'h6EF: dout  = 8'b11100100; // 1775 : 228 - 0xe4
      13'h6F0: dout  = 8'b01111111; // 1776 : 127 - 0x7f -- Sprite 0x6f
      13'h6F1: dout  = 8'b01111111; // 1777 : 127 - 0x7f
      13'h6F2: dout  = 8'b00111111; // 1778 :  63 - 0x3f
      13'h6F3: dout  = 8'b00111111; // 1779 :  63 - 0x3f
      13'h6F4: dout  = 8'b00011111; // 1780 :  31 - 0x1f
      13'h6F5: dout  = 8'b00011111; // 1781 :  31 - 0x1f
      13'h6F6: dout  = 8'b00001111; // 1782 :  15 - 0xf
      13'h6F7: dout  = 8'b00000111; // 1783 :   7 - 0x7
      13'h6F8: dout  = 8'b00000011; // 1784 :   3 - 0x3
      13'h6F9: dout  = 8'b01000100; // 1785 :  68 - 0x44
      13'h6FA: dout  = 8'b00101000; // 1786 :  40 - 0x28
      13'h6FB: dout  = 8'b00010000; // 1787 :  16 - 0x10
      13'h6FC: dout  = 8'b00001000; // 1788 :   8 - 0x8
      13'h6FD: dout  = 8'b00000100; // 1789 :   4 - 0x4
      13'h6FE: dout  = 8'b00000011; // 1790 :   3 - 0x3
      13'h6FF: dout  = 8'b00000100; // 1791 :   4 - 0x4
      13'h700: dout  = 8'b00000011; // 1792 :   3 - 0x3 -- Sprite 0x70
      13'h701: dout  = 8'b00000111; // 1793 :   7 - 0x7
      13'h702: dout  = 8'b00001111; // 1794 :  15 - 0xf
      13'h703: dout  = 8'b00011111; // 1795 :  31 - 0x1f
      13'h704: dout  = 8'b00111111; // 1796 :  63 - 0x3f
      13'h705: dout  = 8'b01110111; // 1797 : 119 - 0x77
      13'h706: dout  = 8'b01110111; // 1798 : 119 - 0x77
      13'h707: dout  = 8'b11110101; // 1799 : 245 - 0xf5
      13'h708: dout  = 8'b00000011; // 1800 :   3 - 0x3
      13'h709: dout  = 8'b00000111; // 1801 :   7 - 0x7
      13'h70A: dout  = 8'b00001111; // 1802 :  15 - 0xf
      13'h70B: dout  = 8'b00011111; // 1803 :  31 - 0x1f
      13'h70C: dout  = 8'b00100111; // 1804 :  39 - 0x27
      13'h70D: dout  = 8'b01111011; // 1805 : 123 - 0x7b
      13'h70E: dout  = 8'b01111000; // 1806 : 120 - 0x78
      13'h70F: dout  = 8'b11111011; // 1807 : 251 - 0xfb
      13'h710: dout  = 8'b11000000; // 1808 : 192 - 0xc0 -- Sprite 0x71
      13'h711: dout  = 8'b11100000; // 1809 : 224 - 0xe0
      13'h712: dout  = 8'b11110000; // 1810 : 240 - 0xf0
      13'h713: dout  = 8'b11111000; // 1811 : 248 - 0xf8
      13'h714: dout  = 8'b11111100; // 1812 : 252 - 0xfc
      13'h715: dout  = 8'b11101110; // 1813 : 238 - 0xee
      13'h716: dout  = 8'b11101110; // 1814 : 238 - 0xee
      13'h717: dout  = 8'b10101111; // 1815 : 175 - 0xaf
      13'h718: dout  = 8'b11000000; // 1816 : 192 - 0xc0
      13'h719: dout  = 8'b11100000; // 1817 : 224 - 0xe0
      13'h71A: dout  = 8'b11110000; // 1818 : 240 - 0xf0
      13'h71B: dout  = 8'b11111000; // 1819 : 248 - 0xf8
      13'h71C: dout  = 8'b11100100; // 1820 : 228 - 0xe4
      13'h71D: dout  = 8'b11011110; // 1821 : 222 - 0xde
      13'h71E: dout  = 8'b00011110; // 1822 :  30 - 0x1e
      13'h71F: dout  = 8'b11011111; // 1823 : 223 - 0xdf
      13'h720: dout  = 8'b11110001; // 1824 : 241 - 0xf1 -- Sprite 0x72
      13'h721: dout  = 8'b11111111; // 1825 : 255 - 0xff
      13'h722: dout  = 8'b01111000; // 1826 : 120 - 0x78
      13'h723: dout  = 8'b00000000; // 1827 :   0 - 0x0
      13'h724: dout  = 8'b00000000; // 1828 :   0 - 0x0
      13'h725: dout  = 8'b00011000; // 1829 :  24 - 0x18
      13'h726: dout  = 8'b00011100; // 1830 :  28 - 0x1c
      13'h727: dout  = 8'b00001110; // 1831 :  14 - 0xe
      13'h728: dout  = 8'b11111111; // 1832 : 255 - 0xff
      13'h729: dout  = 8'b11111111; // 1833 : 255 - 0xff
      13'h72A: dout  = 8'b01111111; // 1834 : 127 - 0x7f
      13'h72B: dout  = 8'b00001111; // 1835 :  15 - 0xf
      13'h72C: dout  = 8'b00001111; // 1836 :  15 - 0xf
      13'h72D: dout  = 8'b00000111; // 1837 :   7 - 0x7
      13'h72E: dout  = 8'b00000011; // 1838 :   3 - 0x3
      13'h72F: dout  = 8'b00000000; // 1839 :   0 - 0x0
      13'h730: dout  = 8'b10001111; // 1840 : 143 - 0x8f -- Sprite 0x73
      13'h731: dout  = 8'b11111111; // 1841 : 255 - 0xff
      13'h732: dout  = 8'b00011110; // 1842 :  30 - 0x1e
      13'h733: dout  = 8'b00000000; // 1843 :   0 - 0x0
      13'h734: dout  = 8'b00001100; // 1844 :  12 - 0xc
      13'h735: dout  = 8'b00111110; // 1845 :  62 - 0x3e
      13'h736: dout  = 8'b01111110; // 1846 : 126 - 0x7e
      13'h737: dout  = 8'b01111100; // 1847 : 124 - 0x7c
      13'h738: dout  = 8'b11111111; // 1848 : 255 - 0xff
      13'h739: dout  = 8'b11111111; // 1849 : 255 - 0xff
      13'h73A: dout  = 8'b11111110; // 1850 : 254 - 0xfe
      13'h73B: dout  = 8'b11110000; // 1851 : 240 - 0xf0
      13'h73C: dout  = 8'b11110000; // 1852 : 240 - 0xf0
      13'h73D: dout  = 8'b11000000; // 1853 : 192 - 0xc0
      13'h73E: dout  = 8'b10000000; // 1854 : 128 - 0x80
      13'h73F: dout  = 8'b00000000; // 1855 :   0 - 0x0
      13'h740: dout  = 8'b00000000; // 1856 :   0 - 0x0 -- Sprite 0x74
      13'h741: dout  = 8'b00000000; // 1857 :   0 - 0x0
      13'h742: dout  = 8'b00000000; // 1858 :   0 - 0x0
      13'h743: dout  = 8'b00000000; // 1859 :   0 - 0x0
      13'h744: dout  = 8'b00000000; // 1860 :   0 - 0x0
      13'h745: dout  = 8'b00000000; // 1861 :   0 - 0x0
      13'h746: dout  = 8'b00000000; // 1862 :   0 - 0x0
      13'h747: dout  = 8'b00000000; // 1863 :   0 - 0x0
      13'h748: dout  = 8'b00000000; // 1864 :   0 - 0x0
      13'h749: dout  = 8'b00000000; // 1865 :   0 - 0x0
      13'h74A: dout  = 8'b00011000; // 1866 :  24 - 0x18
      13'h74B: dout  = 8'b00100100; // 1867 :  36 - 0x24
      13'h74C: dout  = 8'b00100100; // 1868 :  36 - 0x24
      13'h74D: dout  = 8'b00011000; // 1869 :  24 - 0x18
      13'h74E: dout  = 8'b00000000; // 1870 :   0 - 0x0
      13'h74F: dout  = 8'b00000000; // 1871 :   0 - 0x0
      13'h750: dout  = 8'b00000000; // 1872 :   0 - 0x0 -- Sprite 0x75
      13'h751: dout  = 8'b00000010; // 1873 :   2 - 0x2
      13'h752: dout  = 8'b01000001; // 1874 :  65 - 0x41
      13'h753: dout  = 8'b01000001; // 1875 :  65 - 0x41
      13'h754: dout  = 8'b01100001; // 1876 :  97 - 0x61
      13'h755: dout  = 8'b00110011; // 1877 :  51 - 0x33
      13'h756: dout  = 8'b00000110; // 1878 :   6 - 0x6
      13'h757: dout  = 8'b00111100; // 1879 :  60 - 0x3c
      13'h758: dout  = 8'b00111100; // 1880 :  60 - 0x3c
      13'h759: dout  = 8'b01111110; // 1881 : 126 - 0x7e
      13'h75A: dout  = 8'b11111111; // 1882 : 255 - 0xff
      13'h75B: dout  = 8'b11111111; // 1883 : 255 - 0xff
      13'h75C: dout  = 8'b11111111; // 1884 : 255 - 0xff
      13'h75D: dout  = 8'b11111111; // 1885 : 255 - 0xff
      13'h75E: dout  = 8'b01111110; // 1886 : 126 - 0x7e
      13'h75F: dout  = 8'b00111100; // 1887 :  60 - 0x3c
      13'h760: dout  = 8'b00000011; // 1888 :   3 - 0x3 -- Sprite 0x76
      13'h761: dout  = 8'b00000111; // 1889 :   7 - 0x7
      13'h762: dout  = 8'b00001111; // 1890 :  15 - 0xf
      13'h763: dout  = 8'b00011111; // 1891 :  31 - 0x1f
      13'h764: dout  = 8'b00111111; // 1892 :  63 - 0x3f
      13'h765: dout  = 8'b01111111; // 1893 : 127 - 0x7f
      13'h766: dout  = 8'b01111111; // 1894 : 127 - 0x7f
      13'h767: dout  = 8'b11111111; // 1895 : 255 - 0xff
      13'h768: dout  = 8'b00000011; // 1896 :   3 - 0x3
      13'h769: dout  = 8'b00000111; // 1897 :   7 - 0x7
      13'h76A: dout  = 8'b00001111; // 1898 :  15 - 0xf
      13'h76B: dout  = 8'b00011111; // 1899 :  31 - 0x1f
      13'h76C: dout  = 8'b00111111; // 1900 :  63 - 0x3f
      13'h76D: dout  = 8'b01100011; // 1901 :  99 - 0x63
      13'h76E: dout  = 8'b01000001; // 1902 :  65 - 0x41
      13'h76F: dout  = 8'b11000001; // 1903 : 193 - 0xc1
      13'h770: dout  = 8'b11000000; // 1904 : 192 - 0xc0 -- Sprite 0x77
      13'h771: dout  = 8'b11100000; // 1905 : 224 - 0xe0
      13'h772: dout  = 8'b11110000; // 1906 : 240 - 0xf0
      13'h773: dout  = 8'b11111000; // 1907 : 248 - 0xf8
      13'h774: dout  = 8'b11111100; // 1908 : 252 - 0xfc
      13'h775: dout  = 8'b11111110; // 1909 : 254 - 0xfe
      13'h776: dout  = 8'b11111110; // 1910 : 254 - 0xfe
      13'h777: dout  = 8'b11111111; // 1911 : 255 - 0xff
      13'h778: dout  = 8'b11000000; // 1912 : 192 - 0xc0
      13'h779: dout  = 8'b10000000; // 1913 : 128 - 0x80
      13'h77A: dout  = 8'b00000000; // 1914 :   0 - 0x0
      13'h77B: dout  = 8'b00000000; // 1915 :   0 - 0x0
      13'h77C: dout  = 8'b10001100; // 1916 : 140 - 0x8c
      13'h77D: dout  = 8'b11111110; // 1917 : 254 - 0xfe
      13'h77E: dout  = 8'b11111110; // 1918 : 254 - 0xfe
      13'h77F: dout  = 8'b11110011; // 1919 : 243 - 0xf3
      13'h780: dout  = 8'b11111111; // 1920 : 255 - 0xff -- Sprite 0x78
      13'h781: dout  = 8'b11111111; // 1921 : 255 - 0xff
      13'h782: dout  = 8'b11111111; // 1922 : 255 - 0xff
      13'h783: dout  = 8'b01111000; // 1923 : 120 - 0x78
      13'h784: dout  = 8'b00000000; // 1924 :   0 - 0x0
      13'h785: dout  = 8'b00000000; // 1925 :   0 - 0x0
      13'h786: dout  = 8'b00000000; // 1926 :   0 - 0x0
      13'h787: dout  = 8'b00000000; // 1927 :   0 - 0x0
      13'h788: dout  = 8'b11000001; // 1928 : 193 - 0xc1
      13'h789: dout  = 8'b11100011; // 1929 : 227 - 0xe3
      13'h78A: dout  = 8'b11111111; // 1930 : 255 - 0xff
      13'h78B: dout  = 8'b01000111; // 1931 :  71 - 0x47
      13'h78C: dout  = 8'b00001111; // 1932 :  15 - 0xf
      13'h78D: dout  = 8'b00001111; // 1933 :  15 - 0xf
      13'h78E: dout  = 8'b00001111; // 1934 :  15 - 0xf
      13'h78F: dout  = 8'b00000111; // 1935 :   7 - 0x7
      13'h790: dout  = 8'b11111111; // 1936 : 255 - 0xff -- Sprite 0x79
      13'h791: dout  = 8'b11111111; // 1937 : 255 - 0xff
      13'h792: dout  = 8'b11111111; // 1938 : 255 - 0xff
      13'h793: dout  = 8'b00011110; // 1939 :  30 - 0x1e
      13'h794: dout  = 8'b00000000; // 1940 :   0 - 0x0
      13'h795: dout  = 8'b00100000; // 1941 :  32 - 0x20
      13'h796: dout  = 8'b00100000; // 1942 :  32 - 0x20
      13'h797: dout  = 8'b01000000; // 1943 :  64 - 0x40
      13'h798: dout  = 8'b11110001; // 1944 : 241 - 0xf1
      13'h799: dout  = 8'b11111001; // 1945 : 249 - 0xf9
      13'h79A: dout  = 8'b11111111; // 1946 : 255 - 0xff
      13'h79B: dout  = 8'b11100010; // 1947 : 226 - 0xe2
      13'h79C: dout  = 8'b11110000; // 1948 : 240 - 0xf0
      13'h79D: dout  = 8'b11110000; // 1949 : 240 - 0xf0
      13'h79E: dout  = 8'b11110000; // 1950 : 240 - 0xf0
      13'h79F: dout  = 8'b11100000; // 1951 : 224 - 0xe0
      13'h7A0: dout  = 8'b00010110; // 1952 :  22 - 0x16 -- Sprite 0x7a
      13'h7A1: dout  = 8'b00011111; // 1953 :  31 - 0x1f
      13'h7A2: dout  = 8'b00111111; // 1954 :  63 - 0x3f
      13'h7A3: dout  = 8'b01111111; // 1955 : 127 - 0x7f
      13'h7A4: dout  = 8'b00111101; // 1956 :  61 - 0x3d
      13'h7A5: dout  = 8'b00011101; // 1957 :  29 - 0x1d
      13'h7A6: dout  = 8'b00111111; // 1958 :  63 - 0x3f
      13'h7A7: dout  = 8'b00011111; // 1959 :  31 - 0x1f
      13'h7A8: dout  = 8'b00010110; // 1960 :  22 - 0x16
      13'h7A9: dout  = 8'b00011111; // 1961 :  31 - 0x1f
      13'h7AA: dout  = 8'b00000000; // 1962 :   0 - 0x0
      13'h7AB: dout  = 8'b00000000; // 1963 :   0 - 0x0
      13'h7AC: dout  = 8'b00000101; // 1964 :   5 - 0x5
      13'h7AD: dout  = 8'b00001101; // 1965 :  13 - 0xd
      13'h7AE: dout  = 8'b00111111; // 1966 :  63 - 0x3f
      13'h7AF: dout  = 8'b00011111; // 1967 :  31 - 0x1f
      13'h7B0: dout  = 8'b10000000; // 1968 : 128 - 0x80 -- Sprite 0x7b
      13'h7B1: dout  = 8'b10000000; // 1969 : 128 - 0x80
      13'h7B2: dout  = 8'b11000000; // 1970 : 192 - 0xc0
      13'h7B3: dout  = 8'b11100000; // 1971 : 224 - 0xe0
      13'h7B4: dout  = 8'b11110000; // 1972 : 240 - 0xf0
      13'h7B5: dout  = 8'b11110000; // 1973 : 240 - 0xf0
      13'h7B6: dout  = 8'b11110000; // 1974 : 240 - 0xf0
      13'h7B7: dout  = 8'b11111000; // 1975 : 248 - 0xf8
      13'h7B8: dout  = 8'b10000000; // 1976 : 128 - 0x80
      13'h7B9: dout  = 8'b10000000; // 1977 : 128 - 0x80
      13'h7BA: dout  = 8'b00000000; // 1978 :   0 - 0x0
      13'h7BB: dout  = 8'b00000000; // 1979 :   0 - 0x0
      13'h7BC: dout  = 8'b00000000; // 1980 :   0 - 0x0
      13'h7BD: dout  = 8'b10100000; // 1981 : 160 - 0xa0
      13'h7BE: dout  = 8'b10100000; // 1982 : 160 - 0xa0
      13'h7BF: dout  = 8'b11100000; // 1983 : 224 - 0xe0
      13'h7C0: dout  = 8'b00111100; // 1984 :  60 - 0x3c -- Sprite 0x7c
      13'h7C1: dout  = 8'b11111010; // 1985 : 250 - 0xfa
      13'h7C2: dout  = 8'b10110001; // 1986 : 177 - 0xb1
      13'h7C3: dout  = 8'b01110010; // 1987 : 114 - 0x72
      13'h7C4: dout  = 8'b11110010; // 1988 : 242 - 0xf2
      13'h7C5: dout  = 8'b11011011; // 1989 : 219 - 0xdb
      13'h7C6: dout  = 8'b11011111; // 1990 : 223 - 0xdf
      13'h7C7: dout  = 8'b01011111; // 1991 :  95 - 0x5f
      13'h7C8: dout  = 8'b00000000; // 1992 :   0 - 0x0
      13'h7C9: dout  = 8'b00000100; // 1993 :   4 - 0x4
      13'h7CA: dout  = 8'b01001110; // 1994 :  78 - 0x4e
      13'h7CB: dout  = 8'b10001100; // 1995 : 140 - 0x8c
      13'h7CC: dout  = 8'b00001100; // 1996 :  12 - 0xc
      13'h7CD: dout  = 8'b01111111; // 1997 : 127 - 0x7f
      13'h7CE: dout  = 8'b11111111; // 1998 : 255 - 0xff
      13'h7CF: dout  = 8'b11111111; // 1999 : 255 - 0xff
      13'h7D0: dout  = 8'b00000000; // 2000 :   0 - 0x0 -- Sprite 0x7d
      13'h7D1: dout  = 8'b00000000; // 2001 :   0 - 0x0
      13'h7D2: dout  = 8'b00000000; // 2002 :   0 - 0x0
      13'h7D3: dout  = 8'b00000001; // 2003 :   1 - 0x1
      13'h7D4: dout  = 8'b00000001; // 2004 :   1 - 0x1
      13'h7D5: dout  = 8'b00000001; // 2005 :   1 - 0x1
      13'h7D6: dout  = 8'b00000110; // 2006 :   6 - 0x6
      13'h7D7: dout  = 8'b00011110; // 2007 :  30 - 0x1e
      13'h7D8: dout  = 8'b00000000; // 2008 :   0 - 0x0
      13'h7D9: dout  = 8'b00000000; // 2009 :   0 - 0x0
      13'h7DA: dout  = 8'b00000000; // 2010 :   0 - 0x0
      13'h7DB: dout  = 8'b00000000; // 2011 :   0 - 0x0
      13'h7DC: dout  = 8'b00000000; // 2012 :   0 - 0x0
      13'h7DD: dout  = 8'b00000000; // 2013 :   0 - 0x0
      13'h7DE: dout  = 8'b00000001; // 2014 :   1 - 0x1
      13'h7DF: dout  = 8'b00000001; // 2015 :   1 - 0x1
      13'h7E0: dout  = 8'b00000000; // 2016 :   0 - 0x0 -- Sprite 0x7e
      13'h7E1: dout  = 8'b00000000; // 2017 :   0 - 0x0
      13'h7E2: dout  = 8'b00000000; // 2018 :   0 - 0x0
      13'h7E3: dout  = 8'b00000000; // 2019 :   0 - 0x0
      13'h7E4: dout  = 8'b00000000; // 2020 :   0 - 0x0
      13'h7E5: dout  = 8'b00000000; // 2021 :   0 - 0x0
      13'h7E6: dout  = 8'b00000000; // 2022 :   0 - 0x0
      13'h7E7: dout  = 8'b00000000; // 2023 :   0 - 0x0
      13'h7E8: dout  = 8'b11111111; // 2024 : 255 - 0xff
      13'h7E9: dout  = 8'b01111111; // 2025 : 127 - 0x7f
      13'h7EA: dout  = 8'b00111111; // 2026 :  63 - 0x3f
      13'h7EB: dout  = 8'b00011111; // 2027 :  31 - 0x1f
      13'h7EC: dout  = 8'b00001111; // 2028 :  15 - 0xf
      13'h7ED: dout  = 8'b00000111; // 2029 :   7 - 0x7
      13'h7EE: dout  = 8'b00000011; // 2030 :   3 - 0x3
      13'h7EF: dout  = 8'b00000001; // 2031 :   1 - 0x1
      13'h7F0: dout  = 8'b00000000; // 2032 :   0 - 0x0 -- Sprite 0x7f
      13'h7F1: dout  = 8'b01111100; // 2033 : 124 - 0x7c
      13'h7F2: dout  = 8'b11010110; // 2034 : 214 - 0xd6
      13'h7F3: dout  = 8'b10010010; // 2035 : 146 - 0x92
      13'h7F4: dout  = 8'b10111010; // 2036 : 186 - 0xba
      13'h7F5: dout  = 8'b11101110; // 2037 : 238 - 0xee
      13'h7F6: dout  = 8'b11111110; // 2038 : 254 - 0xfe
      13'h7F7: dout  = 8'b00111000; // 2039 :  56 - 0x38
      13'h7F8: dout  = 8'b11111111; // 2040 : 255 - 0xff
      13'h7F9: dout  = 8'b10000011; // 2041 : 131 - 0x83
      13'h7FA: dout  = 8'b00101001; // 2042 :  41 - 0x29
      13'h7FB: dout  = 8'b01101101; // 2043 : 109 - 0x6d
      13'h7FC: dout  = 8'b01000101; // 2044 :  69 - 0x45
      13'h7FD: dout  = 8'b00010001; // 2045 :  17 - 0x11
      13'h7FE: dout  = 8'b00000001; // 2046 :   1 - 0x1
      13'h7FF: dout  = 8'b11000111; // 2047 : 199 - 0xc7
      13'h800: dout  = 8'b00000000; // 2048 :   0 - 0x0 -- Sprite 0x80
      13'h801: dout  = 8'b00010101; // 2049 :  21 - 0x15
      13'h802: dout  = 8'b00111111; // 2050 :  63 - 0x3f
      13'h803: dout  = 8'b01100010; // 2051 :  98 - 0x62
      13'h804: dout  = 8'b01011111; // 2052 :  95 - 0x5f
      13'h805: dout  = 8'b11111111; // 2053 : 255 - 0xff
      13'h806: dout  = 8'b10011111; // 2054 : 159 - 0x9f
      13'h807: dout  = 8'b01111101; // 2055 : 125 - 0x7d
      13'h808: dout  = 8'b00001000; // 2056 :   8 - 0x8
      13'h809: dout  = 8'b00001000; // 2057 :   8 - 0x8
      13'h80A: dout  = 8'b00000010; // 2058 :   2 - 0x2
      13'h80B: dout  = 8'b00011111; // 2059 :  31 - 0x1f
      13'h80C: dout  = 8'b00100010; // 2060 :  34 - 0x22
      13'h80D: dout  = 8'b00000010; // 2061 :   2 - 0x2
      13'h80E: dout  = 8'b00000010; // 2062 :   2 - 0x2
      13'h80F: dout  = 8'b00000000; // 2063 :   0 - 0x0
      13'h810: dout  = 8'b00000000; // 2064 :   0 - 0x0 -- Sprite 0x81
      13'h811: dout  = 8'b00000000; // 2065 :   0 - 0x0
      13'h812: dout  = 8'b00000000; // 2066 :   0 - 0x0
      13'h813: dout  = 8'b00000000; // 2067 :   0 - 0x0
      13'h814: dout  = 8'b00000000; // 2068 :   0 - 0x0
      13'h815: dout  = 8'b00000000; // 2069 :   0 - 0x0
      13'h816: dout  = 8'b00000000; // 2070 :   0 - 0x0
      13'h817: dout  = 8'b00000000; // 2071 :   0 - 0x0
      13'h818: dout  = 8'b00001000; // 2072 :   8 - 0x8
      13'h819: dout  = 8'b00001000; // 2073 :   8 - 0x8
      13'h81A: dout  = 8'b00001000; // 2074 :   8 - 0x8
      13'h81B: dout  = 8'b00001000; // 2075 :   8 - 0x8
      13'h81C: dout  = 8'b00001000; // 2076 :   8 - 0x8
      13'h81D: dout  = 8'b00001000; // 2077 :   8 - 0x8
      13'h81E: dout  = 8'b00001000; // 2078 :   8 - 0x8
      13'h81F: dout  = 8'b00001000; // 2079 :   8 - 0x8
      13'h820: dout  = 8'b00101111; // 2080 :  47 - 0x2f -- Sprite 0x82
      13'h821: dout  = 8'b00011110; // 2081 :  30 - 0x1e
      13'h822: dout  = 8'b00101111; // 2082 :  47 - 0x2f
      13'h823: dout  = 8'b00101111; // 2083 :  47 - 0x2f
      13'h824: dout  = 8'b00101111; // 2084 :  47 - 0x2f
      13'h825: dout  = 8'b00010101; // 2085 :  21 - 0x15
      13'h826: dout  = 8'b00001101; // 2086 :  13 - 0xd
      13'h827: dout  = 8'b00001110; // 2087 :  14 - 0xe
      13'h828: dout  = 8'b00010000; // 2088 :  16 - 0x10
      13'h829: dout  = 8'b00011110; // 2089 :  30 - 0x1e
      13'h82A: dout  = 8'b00010000; // 2090 :  16 - 0x10
      13'h82B: dout  = 8'b01010000; // 2091 :  80 - 0x50
      13'h82C: dout  = 8'b00010000; // 2092 :  16 - 0x10
      13'h82D: dout  = 8'b00001000; // 2093 :   8 - 0x8
      13'h82E: dout  = 8'b00000000; // 2094 :   0 - 0x0
      13'h82F: dout  = 8'b00000000; // 2095 :   0 - 0x0
      13'h830: dout  = 8'b00000000; // 2096 :   0 - 0x0 -- Sprite 0x83
      13'h831: dout  = 8'b00000000; // 2097 :   0 - 0x0
      13'h832: dout  = 8'b00000000; // 2098 :   0 - 0x0
      13'h833: dout  = 8'b00000000; // 2099 :   0 - 0x0
      13'h834: dout  = 8'b00000000; // 2100 :   0 - 0x0
      13'h835: dout  = 8'b00000000; // 2101 :   0 - 0x0
      13'h836: dout  = 8'b00000000; // 2102 :   0 - 0x0
      13'h837: dout  = 8'b00000000; // 2103 :   0 - 0x0
      13'h838: dout  = 8'b00000000; // 2104 :   0 - 0x0
      13'h839: dout  = 8'b00000000; // 2105 :   0 - 0x0
      13'h83A: dout  = 8'b00000000; // 2106 :   0 - 0x0
      13'h83B: dout  = 8'b11111110; // 2107 : 254 - 0xfe
      13'h83C: dout  = 8'b00000000; // 2108 :   0 - 0x0
      13'h83D: dout  = 8'b00000000; // 2109 :   0 - 0x0
      13'h83E: dout  = 8'b00000000; // 2110 :   0 - 0x0
      13'h83F: dout  = 8'b00000000; // 2111 :   0 - 0x0
      13'h840: dout  = 8'b00011100; // 2112 :  28 - 0x1c -- Sprite 0x84
      13'h841: dout  = 8'b00111110; // 2113 :  62 - 0x3e
      13'h842: dout  = 8'b01111111; // 2114 : 127 - 0x7f
      13'h843: dout  = 8'b11111111; // 2115 : 255 - 0xff
      13'h844: dout  = 8'b11111111; // 2116 : 255 - 0xff
      13'h845: dout  = 8'b11111110; // 2117 : 254 - 0xfe
      13'h846: dout  = 8'b01111100; // 2118 : 124 - 0x7c
      13'h847: dout  = 8'b00111000; // 2119 :  56 - 0x38
      13'h848: dout  = 8'b00011100; // 2120 :  28 - 0x1c
      13'h849: dout  = 8'b00101010; // 2121 :  42 - 0x2a
      13'h84A: dout  = 8'b01110111; // 2122 : 119 - 0x77
      13'h84B: dout  = 8'b11101110; // 2123 : 238 - 0xee
      13'h84C: dout  = 8'b11011101; // 2124 : 221 - 0xdd
      13'h84D: dout  = 8'b10101010; // 2125 : 170 - 0xaa
      13'h84E: dout  = 8'b01110100; // 2126 : 116 - 0x74
      13'h84F: dout  = 8'b00101000; // 2127 :  40 - 0x28
      13'h850: dout  = 8'b00000000; // 2128 :   0 - 0x0 -- Sprite 0x85
      13'h851: dout  = 8'b11111111; // 2129 : 255 - 0xff
      13'h852: dout  = 8'b11111111; // 2130 : 255 - 0xff
      13'h853: dout  = 8'b11111111; // 2131 : 255 - 0xff
      13'h854: dout  = 8'b11111111; // 2132 : 255 - 0xff
      13'h855: dout  = 8'b11111111; // 2133 : 255 - 0xff
      13'h856: dout  = 8'b11111111; // 2134 : 255 - 0xff
      13'h857: dout  = 8'b11111111; // 2135 : 255 - 0xff
      13'h858: dout  = 8'b11111111; // 2136 : 255 - 0xff
      13'h859: dout  = 8'b11111110; // 2137 : 254 - 0xfe
      13'h85A: dout  = 8'b11111110; // 2138 : 254 - 0xfe
      13'h85B: dout  = 8'b00000000; // 2139 :   0 - 0x0
      13'h85C: dout  = 8'b11101111; // 2140 : 239 - 0xef
      13'h85D: dout  = 8'b11101111; // 2141 : 239 - 0xef
      13'h85E: dout  = 8'b11101111; // 2142 : 239 - 0xef
      13'h85F: dout  = 8'b00000000; // 2143 :   0 - 0x0
      13'h860: dout  = 8'b11111111; // 2144 : 255 - 0xff -- Sprite 0x86
      13'h861: dout  = 8'b11111111; // 2145 : 255 - 0xff
      13'h862: dout  = 8'b11111111; // 2146 : 255 - 0xff
      13'h863: dout  = 8'b11111111; // 2147 : 255 - 0xff
      13'h864: dout  = 8'b11111111; // 2148 : 255 - 0xff
      13'h865: dout  = 8'b11111111; // 2149 : 255 - 0xff
      13'h866: dout  = 8'b11111111; // 2150 : 255 - 0xff
      13'h867: dout  = 8'b11111111; // 2151 : 255 - 0xff
      13'h868: dout  = 8'b11111110; // 2152 : 254 - 0xfe
      13'h869: dout  = 8'b11111110; // 2153 : 254 - 0xfe
      13'h86A: dout  = 8'b11111110; // 2154 : 254 - 0xfe
      13'h86B: dout  = 8'b00000000; // 2155 :   0 - 0x0
      13'h86C: dout  = 8'b11101111; // 2156 : 239 - 0xef
      13'h86D: dout  = 8'b11101111; // 2157 : 239 - 0xef
      13'h86E: dout  = 8'b11101111; // 2158 : 239 - 0xef
      13'h86F: dout  = 8'b00000000; // 2159 :   0 - 0x0
      13'h870: dout  = 8'b01111111; // 2160 : 127 - 0x7f -- Sprite 0x87
      13'h871: dout  = 8'b11111111; // 2161 : 255 - 0xff
      13'h872: dout  = 8'b11111111; // 2162 : 255 - 0xff
      13'h873: dout  = 8'b11111111; // 2163 : 255 - 0xff
      13'h874: dout  = 8'b11111111; // 2164 : 255 - 0xff
      13'h875: dout  = 8'b11111111; // 2165 : 255 - 0xff
      13'h876: dout  = 8'b11111111; // 2166 : 255 - 0xff
      13'h877: dout  = 8'b11111111; // 2167 : 255 - 0xff
      13'h878: dout  = 8'b00000000; // 2168 :   0 - 0x0
      13'h879: dout  = 8'b01111111; // 2169 : 127 - 0x7f
      13'h87A: dout  = 8'b01011111; // 2170 :  95 - 0x5f
      13'h87B: dout  = 8'b01111111; // 2171 : 127 - 0x7f
      13'h87C: dout  = 8'b01111111; // 2172 : 127 - 0x7f
      13'h87D: dout  = 8'b01111111; // 2173 : 127 - 0x7f
      13'h87E: dout  = 8'b01111111; // 2174 : 127 - 0x7f
      13'h87F: dout  = 8'b01111111; // 2175 : 127 - 0x7f
      13'h880: dout  = 8'b01101000; // 2176 : 104 - 0x68 -- Sprite 0x88
      13'h881: dout  = 8'b01001110; // 2177 :  78 - 0x4e
      13'h882: dout  = 8'b11100000; // 2178 : 224 - 0xe0
      13'h883: dout  = 8'b11100000; // 2179 : 224 - 0xe0
      13'h884: dout  = 8'b11100000; // 2180 : 224 - 0xe0
      13'h885: dout  = 8'b11110000; // 2181 : 240 - 0xf0
      13'h886: dout  = 8'b11111000; // 2182 : 248 - 0xf8
      13'h887: dout  = 8'b11111100; // 2183 : 252 - 0xfc
      13'h888: dout  = 8'b10111000; // 2184 : 184 - 0xb8
      13'h889: dout  = 8'b10011110; // 2185 : 158 - 0x9e
      13'h88A: dout  = 8'b10000000; // 2186 : 128 - 0x80
      13'h88B: dout  = 8'b11000000; // 2187 : 192 - 0xc0
      13'h88C: dout  = 8'b11100000; // 2188 : 224 - 0xe0
      13'h88D: dout  = 8'b11110000; // 2189 : 240 - 0xf0
      13'h88E: dout  = 8'b11111000; // 2190 : 248 - 0xf8
      13'h88F: dout  = 8'b01111100; // 2191 : 124 - 0x7c
      13'h890: dout  = 8'b00111111; // 2192 :  63 - 0x3f -- Sprite 0x89
      13'h891: dout  = 8'b01011100; // 2193 :  92 - 0x5c
      13'h892: dout  = 8'b00111001; // 2194 :  57 - 0x39
      13'h893: dout  = 8'b00111011; // 2195 :  59 - 0x3b
      13'h894: dout  = 8'b10111011; // 2196 : 187 - 0xbb
      13'h895: dout  = 8'b11111001; // 2197 : 249 - 0xf9
      13'h896: dout  = 8'b11111100; // 2198 : 252 - 0xfc
      13'h897: dout  = 8'b11111110; // 2199 : 254 - 0xfe
      13'h898: dout  = 8'b00000000; // 2200 :   0 - 0x0
      13'h899: dout  = 8'b00100011; // 2201 :  35 - 0x23
      13'h89A: dout  = 8'b01010111; // 2202 :  87 - 0x57
      13'h89B: dout  = 8'b01001111; // 2203 :  79 - 0x4f
      13'h89C: dout  = 8'b01010111; // 2204 :  87 - 0x57
      13'h89D: dout  = 8'b00100111; // 2205 :  39 - 0x27
      13'h89E: dout  = 8'b11000011; // 2206 : 195 - 0xc3
      13'h89F: dout  = 8'b00100001; // 2207 :  33 - 0x21
      13'h8A0: dout  = 8'b11000000; // 2208 : 192 - 0xc0 -- Sprite 0x8a
      13'h8A1: dout  = 8'b11110000; // 2209 : 240 - 0xf0
      13'h8A2: dout  = 8'b11110000; // 2210 : 240 - 0xf0
      13'h8A3: dout  = 8'b11110000; // 2211 : 240 - 0xf0
      13'h8A4: dout  = 8'b11110000; // 2212 : 240 - 0xf0
      13'h8A5: dout  = 8'b11100000; // 2213 : 224 - 0xe0
      13'h8A6: dout  = 8'b11000000; // 2214 : 192 - 0xc0
      13'h8A7: dout  = 8'b00000000; // 2215 :   0 - 0x0
      13'h8A8: dout  = 8'b00000000; // 2216 :   0 - 0x0
      13'h8A9: dout  = 8'b00110000; // 2217 :  48 - 0x30
      13'h8AA: dout  = 8'b01110000; // 2218 : 112 - 0x70
      13'h8AB: dout  = 8'b01110000; // 2219 : 112 - 0x70
      13'h8AC: dout  = 8'b11110000; // 2220 : 240 - 0xf0
      13'h8AD: dout  = 8'b11100000; // 2221 : 224 - 0xe0
      13'h8AE: dout  = 8'b11000000; // 2222 : 192 - 0xc0
      13'h8AF: dout  = 8'b00000000; // 2223 :   0 - 0x0
      13'h8B0: dout  = 8'b11111110; // 2224 : 254 - 0xfe -- Sprite 0x8b
      13'h8B1: dout  = 8'b11111100; // 2225 : 252 - 0xfc
      13'h8B2: dout  = 8'b01100001; // 2226 :  97 - 0x61
      13'h8B3: dout  = 8'b00001111; // 2227 :  15 - 0xf
      13'h8B4: dout  = 8'b11111111; // 2228 : 255 - 0xff
      13'h8B5: dout  = 8'b11111110; // 2229 : 254 - 0xfe
      13'h8B6: dout  = 8'b11110000; // 2230 : 240 - 0xf0
      13'h8B7: dout  = 8'b11100000; // 2231 : 224 - 0xe0
      13'h8B8: dout  = 8'b00010011; // 2232 :  19 - 0x13
      13'h8B9: dout  = 8'b00001111; // 2233 :  15 - 0xf
      13'h8BA: dout  = 8'b00011110; // 2234 :  30 - 0x1e
      13'h8BB: dout  = 8'b11110000; // 2235 : 240 - 0xf0
      13'h8BC: dout  = 8'b11111100; // 2236 : 252 - 0xfc
      13'h8BD: dout  = 8'b11111000; // 2237 : 248 - 0xf8
      13'h8BE: dout  = 8'b11110000; // 2238 : 240 - 0xf0
      13'h8BF: dout  = 8'b11100000; // 2239 : 224 - 0xe0
      13'h8C0: dout  = 8'b01101110; // 2240 : 110 - 0x6e -- Sprite 0x8c
      13'h8C1: dout  = 8'b01000000; // 2241 :  64 - 0x40
      13'h8C2: dout  = 8'b11100000; // 2242 : 224 - 0xe0
      13'h8C3: dout  = 8'b11100000; // 2243 : 224 - 0xe0
      13'h8C4: dout  = 8'b11100000; // 2244 : 224 - 0xe0
      13'h8C5: dout  = 8'b11100000; // 2245 : 224 - 0xe0
      13'h8C6: dout  = 8'b11100000; // 2246 : 224 - 0xe0
      13'h8C7: dout  = 8'b11000000; // 2247 : 192 - 0xc0
      13'h8C8: dout  = 8'b10111110; // 2248 : 190 - 0xbe
      13'h8C9: dout  = 8'b10010000; // 2249 : 144 - 0x90
      13'h8CA: dout  = 8'b10000000; // 2250 : 128 - 0x80
      13'h8CB: dout  = 8'b11000000; // 2251 : 192 - 0xc0
      13'h8CC: dout  = 8'b11000000; // 2252 : 192 - 0xc0
      13'h8CD: dout  = 8'b10000000; // 2253 : 128 - 0x80
      13'h8CE: dout  = 8'b00000000; // 2254 :   0 - 0x0
      13'h8CF: dout  = 8'b00000000; // 2255 :   0 - 0x0
      13'h8D0: dout  = 8'b00000001; // 2256 :   1 - 0x1 -- Sprite 0x8d
      13'h8D1: dout  = 8'b00000001; // 2257 :   1 - 0x1
      13'h8D2: dout  = 8'b00000011; // 2258 :   3 - 0x3
      13'h8D3: dout  = 8'b00000011; // 2259 :   3 - 0x3
      13'h8D4: dout  = 8'b00000111; // 2260 :   7 - 0x7
      13'h8D5: dout  = 8'b01111111; // 2261 : 127 - 0x7f
      13'h8D6: dout  = 8'b01111111; // 2262 : 127 - 0x7f
      13'h8D7: dout  = 8'b00111111; // 2263 :  63 - 0x3f
      13'h8D8: dout  = 8'b00000001; // 2264 :   1 - 0x1
      13'h8D9: dout  = 8'b00000001; // 2265 :   1 - 0x1
      13'h8DA: dout  = 8'b00000011; // 2266 :   3 - 0x3
      13'h8DB: dout  = 8'b00000011; // 2267 :   3 - 0x3
      13'h8DC: dout  = 8'b00000111; // 2268 :   7 - 0x7
      13'h8DD: dout  = 8'b01111111; // 2269 : 127 - 0x7f
      13'h8DE: dout  = 8'b01111101; // 2270 : 125 - 0x7d
      13'h8DF: dout  = 8'b00111101; // 2271 :  61 - 0x3d
      13'h8E0: dout  = 8'b00000110; // 2272 :   6 - 0x6 -- Sprite 0x8e
      13'h8E1: dout  = 8'b00000111; // 2273 :   7 - 0x7
      13'h8E2: dout  = 8'b00111111; // 2274 :  63 - 0x3f
      13'h8E3: dout  = 8'b00111100; // 2275 :  60 - 0x3c
      13'h8E4: dout  = 8'b00011001; // 2276 :  25 - 0x19
      13'h8E5: dout  = 8'b01111011; // 2277 : 123 - 0x7b
      13'h8E6: dout  = 8'b01111111; // 2278 : 127 - 0x7f
      13'h8E7: dout  = 8'b00111111; // 2279 :  63 - 0x3f
      13'h8E8: dout  = 8'b00000110; // 2280 :   6 - 0x6
      13'h8E9: dout  = 8'b00000100; // 2281 :   4 - 0x4
      13'h8EA: dout  = 8'b00110000; // 2282 :  48 - 0x30
      13'h8EB: dout  = 8'b00100011; // 2283 :  35 - 0x23
      13'h8EC: dout  = 8'b00000110; // 2284 :   6 - 0x6
      13'h8ED: dout  = 8'b01100100; // 2285 : 100 - 0x64
      13'h8EE: dout  = 8'b01100000; // 2286 :  96 - 0x60
      13'h8EF: dout  = 8'b00000000; // 2287 :   0 - 0x0
      13'h8F0: dout  = 8'b00111111; // 2288 :  63 - 0x3f -- Sprite 0x8f
      13'h8F1: dout  = 8'b01111111; // 2289 : 127 - 0x7f
      13'h8F2: dout  = 8'b01111111; // 2290 : 127 - 0x7f
      13'h8F3: dout  = 8'b00011111; // 2291 :  31 - 0x1f
      13'h8F4: dout  = 8'b00111111; // 2292 :  63 - 0x3f
      13'h8F5: dout  = 8'b00111111; // 2293 :  63 - 0x3f
      13'h8F6: dout  = 8'b00000111; // 2294 :   7 - 0x7
      13'h8F7: dout  = 8'b00000110; // 2295 :   6 - 0x6
      13'h8F8: dout  = 8'b00000000; // 2296 :   0 - 0x0
      13'h8F9: dout  = 8'b01100000; // 2297 :  96 - 0x60
      13'h8FA: dout  = 8'b01100000; // 2298 :  96 - 0x60
      13'h8FB: dout  = 8'b00000000; // 2299 :   0 - 0x0
      13'h8FC: dout  = 8'b00100000; // 2300 :  32 - 0x20
      13'h8FD: dout  = 8'b00110000; // 2301 :  48 - 0x30
      13'h8FE: dout  = 8'b00000100; // 2302 :   4 - 0x4
      13'h8FF: dout  = 8'b00000110; // 2303 :   6 - 0x6
      13'h900: dout  = 8'b00000011; // 2304 :   3 - 0x3 -- Sprite 0x90
      13'h901: dout  = 8'b00000111; // 2305 :   7 - 0x7
      13'h902: dout  = 8'b00001111; // 2306 :  15 - 0xf
      13'h903: dout  = 8'b00001111; // 2307 :  15 - 0xf
      13'h904: dout  = 8'b00001111; // 2308 :  15 - 0xf
      13'h905: dout  = 8'b00001111; // 2309 :  15 - 0xf
      13'h906: dout  = 8'b00000111; // 2310 :   7 - 0x7
      13'h907: dout  = 8'b00000011; // 2311 :   3 - 0x3
      13'h908: dout  = 8'b00000000; // 2312 :   0 - 0x0
      13'h909: dout  = 8'b00000001; // 2313 :   1 - 0x1
      13'h90A: dout  = 8'b00000001; // 2314 :   1 - 0x1
      13'h90B: dout  = 8'b00000000; // 2315 :   0 - 0x0
      13'h90C: dout  = 8'b00000000; // 2316 :   0 - 0x0
      13'h90D: dout  = 8'b00000000; // 2317 :   0 - 0x0
      13'h90E: dout  = 8'b00000000; // 2318 :   0 - 0x0
      13'h90F: dout  = 8'b00000000; // 2319 :   0 - 0x0
      13'h910: dout  = 8'b11111000; // 2320 : 248 - 0xf8 -- Sprite 0x91
      13'h911: dout  = 8'b11111000; // 2321 : 248 - 0xf8
      13'h912: dout  = 8'b11111000; // 2322 : 248 - 0xf8
      13'h913: dout  = 8'b10100000; // 2323 : 160 - 0xa0
      13'h914: dout  = 8'b11100001; // 2324 : 225 - 0xe1
      13'h915: dout  = 8'b11111111; // 2325 : 255 - 0xff
      13'h916: dout  = 8'b11111111; // 2326 : 255 - 0xff
      13'h917: dout  = 8'b11111111; // 2327 : 255 - 0xff
      13'h918: dout  = 8'b11111110; // 2328 : 254 - 0xfe
      13'h919: dout  = 8'b11111111; // 2329 : 255 - 0xff
      13'h91A: dout  = 8'b11111111; // 2330 : 255 - 0xff
      13'h91B: dout  = 8'b01000000; // 2331 :  64 - 0x40
      13'h91C: dout  = 8'b00000001; // 2332 :   1 - 0x1
      13'h91D: dout  = 8'b00000011; // 2333 :   3 - 0x3
      13'h91E: dout  = 8'b00000011; // 2334 :   3 - 0x3
      13'h91F: dout  = 8'b00000011; // 2335 :   3 - 0x3
      13'h920: dout  = 8'b00001111; // 2336 :  15 - 0xf -- Sprite 0x92
      13'h921: dout  = 8'b00001111; // 2337 :  15 - 0xf
      13'h922: dout  = 8'b00001111; // 2338 :  15 - 0xf
      13'h923: dout  = 8'b00011111; // 2339 :  31 - 0x1f
      13'h924: dout  = 8'b00011111; // 2340 :  31 - 0x1f
      13'h925: dout  = 8'b00011111; // 2341 :  31 - 0x1f
      13'h926: dout  = 8'b00001111; // 2342 :  15 - 0xf
      13'h927: dout  = 8'b00000111; // 2343 :   7 - 0x7
      13'h928: dout  = 8'b00000001; // 2344 :   1 - 0x1
      13'h929: dout  = 8'b00000001; // 2345 :   1 - 0x1
      13'h92A: dout  = 8'b00000000; // 2346 :   0 - 0x0
      13'h92B: dout  = 8'b00000000; // 2347 :   0 - 0x0
      13'h92C: dout  = 8'b00000000; // 2348 :   0 - 0x0
      13'h92D: dout  = 8'b00000000; // 2349 :   0 - 0x0
      13'h92E: dout  = 8'b00000000; // 2350 :   0 - 0x0
      13'h92F: dout  = 8'b00000000; // 2351 :   0 - 0x0
      13'h930: dout  = 8'b11100000; // 2352 : 224 - 0xe0 -- Sprite 0x93
      13'h931: dout  = 8'b11111000; // 2353 : 248 - 0xf8
      13'h932: dout  = 8'b11111000; // 2354 : 248 - 0xf8
      13'h933: dout  = 8'b11111000; // 2355 : 248 - 0xf8
      13'h934: dout  = 8'b11111111; // 2356 : 255 - 0xff
      13'h935: dout  = 8'b11111110; // 2357 : 254 - 0xfe
      13'h936: dout  = 8'b11110000; // 2358 : 240 - 0xf0
      13'h937: dout  = 8'b11000000; // 2359 : 192 - 0xc0
      13'h938: dout  = 8'b11100000; // 2360 : 224 - 0xe0
      13'h939: dout  = 8'b11111110; // 2361 : 254 - 0xfe
      13'h93A: dout  = 8'b11111111; // 2362 : 255 - 0xff
      13'h93B: dout  = 8'b01111111; // 2363 : 127 - 0x7f
      13'h93C: dout  = 8'b00000011; // 2364 :   3 - 0x3
      13'h93D: dout  = 8'b00000010; // 2365 :   2 - 0x2
      13'h93E: dout  = 8'b00000000; // 2366 :   0 - 0x0
      13'h93F: dout  = 8'b00000000; // 2367 :   0 - 0x0
      13'h940: dout  = 8'b00000001; // 2368 :   1 - 0x1 -- Sprite 0x94
      13'h941: dout  = 8'b00001111; // 2369 :  15 - 0xf
      13'h942: dout  = 8'b00001111; // 2370 :  15 - 0xf
      13'h943: dout  = 8'b00011111; // 2371 :  31 - 0x1f
      13'h944: dout  = 8'b00111001; // 2372 :  57 - 0x39
      13'h945: dout  = 8'b00110011; // 2373 :  51 - 0x33
      13'h946: dout  = 8'b00110111; // 2374 :  55 - 0x37
      13'h947: dout  = 8'b01111111; // 2375 : 127 - 0x7f
      13'h948: dout  = 8'b00000001; // 2376 :   1 - 0x1
      13'h949: dout  = 8'b00001101; // 2377 :  13 - 0xd
      13'h94A: dout  = 8'b00001000; // 2378 :   8 - 0x8
      13'h94B: dout  = 8'b00000000; // 2379 :   0 - 0x0
      13'h94C: dout  = 8'b00110110; // 2380 :  54 - 0x36
      13'h94D: dout  = 8'b00101100; // 2381 :  44 - 0x2c
      13'h94E: dout  = 8'b00001000; // 2382 :   8 - 0x8
      13'h94F: dout  = 8'b01100000; // 2383 :  96 - 0x60
      13'h950: dout  = 8'b01111111; // 2384 : 127 - 0x7f -- Sprite 0x95
      13'h951: dout  = 8'b00111111; // 2385 :  63 - 0x3f
      13'h952: dout  = 8'b00111111; // 2386 :  63 - 0x3f
      13'h953: dout  = 8'b00111111; // 2387 :  63 - 0x3f
      13'h954: dout  = 8'b00011111; // 2388 :  31 - 0x1f
      13'h955: dout  = 8'b00001111; // 2389 :  15 - 0xf
      13'h956: dout  = 8'b00001111; // 2390 :  15 - 0xf
      13'h957: dout  = 8'b00000001; // 2391 :   1 - 0x1
      13'h958: dout  = 8'b01100000; // 2392 :  96 - 0x60
      13'h959: dout  = 8'b00000000; // 2393 :   0 - 0x0
      13'h95A: dout  = 8'b00100000; // 2394 :  32 - 0x20
      13'h95B: dout  = 8'b00110000; // 2395 :  48 - 0x30
      13'h95C: dout  = 8'b00000000; // 2396 :   0 - 0x0
      13'h95D: dout  = 8'b00001000; // 2397 :   8 - 0x8
      13'h95E: dout  = 8'b00001101; // 2398 :  13 - 0xd
      13'h95F: dout  = 8'b00000001; // 2399 :   1 - 0x1
      13'h960: dout  = 8'b00000000; // 2400 :   0 - 0x0 -- Sprite 0x96
      13'h961: dout  = 8'b00000000; // 2401 :   0 - 0x0
      13'h962: dout  = 8'b00000011; // 2402 :   3 - 0x3
      13'h963: dout  = 8'b00000011; // 2403 :   3 - 0x3
      13'h964: dout  = 8'b01000111; // 2404 :  71 - 0x47
      13'h965: dout  = 8'b01100111; // 2405 : 103 - 0x67
      13'h966: dout  = 8'b01110111; // 2406 : 119 - 0x77
      13'h967: dout  = 8'b01110111; // 2407 : 119 - 0x77
      13'h968: dout  = 8'b00000001; // 2408 :   1 - 0x1
      13'h969: dout  = 8'b00000001; // 2409 :   1 - 0x1
      13'h96A: dout  = 8'b00000011; // 2410 :   3 - 0x3
      13'h96B: dout  = 8'b01000011; // 2411 :  67 - 0x43
      13'h96C: dout  = 8'b01100111; // 2412 : 103 - 0x67
      13'h96D: dout  = 8'b01110111; // 2413 : 119 - 0x77
      13'h96E: dout  = 8'b01111011; // 2414 : 123 - 0x7b
      13'h96F: dout  = 8'b01111000; // 2415 : 120 - 0x78
      13'h970: dout  = 8'b00000000; // 2416 :   0 - 0x0 -- Sprite 0x97
      13'h971: dout  = 8'b00000000; // 2417 :   0 - 0x0
      13'h972: dout  = 8'b00000000; // 2418 :   0 - 0x0
      13'h973: dout  = 8'b00000000; // 2419 :   0 - 0x0
      13'h974: dout  = 8'b10001000; // 2420 : 136 - 0x88
      13'h975: dout  = 8'b10011000; // 2421 : 152 - 0x98
      13'h976: dout  = 8'b11111000; // 2422 : 248 - 0xf8
      13'h977: dout  = 8'b11110000; // 2423 : 240 - 0xf0
      13'h978: dout  = 8'b00000000; // 2424 :   0 - 0x0
      13'h979: dout  = 8'b00000000; // 2425 :   0 - 0x0
      13'h97A: dout  = 8'b10000000; // 2426 : 128 - 0x80
      13'h97B: dout  = 8'b10000100; // 2427 : 132 - 0x84
      13'h97C: dout  = 8'b11001100; // 2428 : 204 - 0xcc
      13'h97D: dout  = 8'b11011100; // 2429 : 220 - 0xdc
      13'h97E: dout  = 8'b10111100; // 2430 : 188 - 0xbc
      13'h97F: dout  = 8'b00111100; // 2431 :  60 - 0x3c
      13'h980: dout  = 8'b01111110; // 2432 : 126 - 0x7e -- Sprite 0x98
      13'h981: dout  = 8'b01111111; // 2433 : 127 - 0x7f
      13'h982: dout  = 8'b11111111; // 2434 : 255 - 0xff
      13'h983: dout  = 8'b00011111; // 2435 :  31 - 0x1f
      13'h984: dout  = 8'b00000111; // 2436 :   7 - 0x7
      13'h985: dout  = 8'b00110000; // 2437 :  48 - 0x30
      13'h986: dout  = 8'b00011100; // 2438 :  28 - 0x1c
      13'h987: dout  = 8'b00001100; // 2439 :  12 - 0xc
      13'h988: dout  = 8'b00110011; // 2440 :  51 - 0x33
      13'h989: dout  = 8'b00000111; // 2441 :   7 - 0x7
      13'h98A: dout  = 8'b00000111; // 2442 :   7 - 0x7
      13'h98B: dout  = 8'b11100011; // 2443 : 227 - 0xe3
      13'h98C: dout  = 8'b00111000; // 2444 :  56 - 0x38
      13'h98D: dout  = 8'b00111111; // 2445 :  63 - 0x3f
      13'h98E: dout  = 8'b00011100; // 2446 :  28 - 0x1c
      13'h98F: dout  = 8'b00001100; // 2447 :  12 - 0xc
      13'h990: dout  = 8'b01111110; // 2448 : 126 - 0x7e -- Sprite 0x99
      13'h991: dout  = 8'b00111000; // 2449 :  56 - 0x38
      13'h992: dout  = 8'b11110110; // 2450 : 246 - 0xf6
      13'h993: dout  = 8'b11101101; // 2451 : 237 - 0xed
      13'h994: dout  = 8'b11011111; // 2452 : 223 - 0xdf
      13'h995: dout  = 8'b00111000; // 2453 :  56 - 0x38
      13'h996: dout  = 8'b01110000; // 2454 : 112 - 0x70
      13'h997: dout  = 8'b01100000; // 2455 :  96 - 0x60
      13'h998: dout  = 8'b10011000; // 2456 : 152 - 0x98
      13'h999: dout  = 8'b11000111; // 2457 : 199 - 0xc7
      13'h99A: dout  = 8'b11001000; // 2458 : 200 - 0xc8
      13'h99B: dout  = 8'b10010010; // 2459 : 146 - 0x92
      13'h99C: dout  = 8'b00110000; // 2460 :  48 - 0x30
      13'h99D: dout  = 8'b11111000; // 2461 : 248 - 0xf8
      13'h99E: dout  = 8'b01110000; // 2462 : 112 - 0x70
      13'h99F: dout  = 8'b01100000; // 2463 :  96 - 0x60
      13'h9A0: dout  = 8'b00000000; // 2464 :   0 - 0x0 -- Sprite 0x9a
      13'h9A1: dout  = 8'b00000000; // 2465 :   0 - 0x0
      13'h9A2: dout  = 8'b00000000; // 2466 :   0 - 0x0
      13'h9A3: dout  = 8'b00000011; // 2467 :   3 - 0x3
      13'h9A4: dout  = 8'b00000011; // 2468 :   3 - 0x3
      13'h9A5: dout  = 8'b01000111; // 2469 :  71 - 0x47
      13'h9A6: dout  = 8'b01100111; // 2470 : 103 - 0x67
      13'h9A7: dout  = 8'b01110111; // 2471 : 119 - 0x77
      13'h9A8: dout  = 8'b00000000; // 2472 :   0 - 0x0
      13'h9A9: dout  = 8'b00000001; // 2473 :   1 - 0x1
      13'h9AA: dout  = 8'b00000001; // 2474 :   1 - 0x1
      13'h9AB: dout  = 8'b00000011; // 2475 :   3 - 0x3
      13'h9AC: dout  = 8'b01000011; // 2476 :  67 - 0x43
      13'h9AD: dout  = 8'b01100111; // 2477 : 103 - 0x67
      13'h9AE: dout  = 8'b01110111; // 2478 : 119 - 0x77
      13'h9AF: dout  = 8'b01111011; // 2479 : 123 - 0x7b
      13'h9B0: dout  = 8'b00000000; // 2480 :   0 - 0x0 -- Sprite 0x9b
      13'h9B1: dout  = 8'b00000000; // 2481 :   0 - 0x0
      13'h9B2: dout  = 8'b00000000; // 2482 :   0 - 0x0
      13'h9B3: dout  = 8'b00000000; // 2483 :   0 - 0x0
      13'h9B4: dout  = 8'b00000000; // 2484 :   0 - 0x0
      13'h9B5: dout  = 8'b10001000; // 2485 : 136 - 0x88
      13'h9B6: dout  = 8'b10011000; // 2486 : 152 - 0x98
      13'h9B7: dout  = 8'b11111000; // 2487 : 248 - 0xf8
      13'h9B8: dout  = 8'b00000000; // 2488 :   0 - 0x0
      13'h9B9: dout  = 8'b00000000; // 2489 :   0 - 0x0
      13'h9BA: dout  = 8'b00000000; // 2490 :   0 - 0x0
      13'h9BB: dout  = 8'b10000000; // 2491 : 128 - 0x80
      13'h9BC: dout  = 8'b10000100; // 2492 : 132 - 0x84
      13'h9BD: dout  = 8'b11001100; // 2493 : 204 - 0xcc
      13'h9BE: dout  = 8'b11011100; // 2494 : 220 - 0xdc
      13'h9BF: dout  = 8'b10111100; // 2495 : 188 - 0xbc
      13'h9C0: dout  = 8'b01110111; // 2496 : 119 - 0x77 -- Sprite 0x9c
      13'h9C1: dout  = 8'b01111110; // 2497 : 126 - 0x7e
      13'h9C2: dout  = 8'b01111111; // 2498 : 127 - 0x7f
      13'h9C3: dout  = 8'b11111111; // 2499 : 255 - 0xff
      13'h9C4: dout  = 8'b00011111; // 2500 :  31 - 0x1f
      13'h9C5: dout  = 8'b00000111; // 2501 :   7 - 0x7
      13'h9C6: dout  = 8'b01110000; // 2502 : 112 - 0x70
      13'h9C7: dout  = 8'b11110000; // 2503 : 240 - 0xf0
      13'h9C8: dout  = 8'b01111000; // 2504 : 120 - 0x78
      13'h9C9: dout  = 8'b00110011; // 2505 :  51 - 0x33
      13'h9CA: dout  = 8'b00000111; // 2506 :   7 - 0x7
      13'h9CB: dout  = 8'b00000111; // 2507 :   7 - 0x7
      13'h9CC: dout  = 8'b11100011; // 2508 : 227 - 0xe3
      13'h9CD: dout  = 8'b00111000; // 2509 :  56 - 0x38
      13'h9CE: dout  = 8'b01111111; // 2510 : 127 - 0x7f
      13'h9CF: dout  = 8'b11110000; // 2511 : 240 - 0xf0
      13'h9D0: dout  = 8'b11110000; // 2512 : 240 - 0xf0 -- Sprite 0x9d
      13'h9D1: dout  = 8'b01111110; // 2513 : 126 - 0x7e
      13'h9D2: dout  = 8'b00111000; // 2514 :  56 - 0x38
      13'h9D3: dout  = 8'b11110110; // 2515 : 246 - 0xf6
      13'h9D4: dout  = 8'b11101101; // 2516 : 237 - 0xed
      13'h9D5: dout  = 8'b11011111; // 2517 : 223 - 0xdf
      13'h9D6: dout  = 8'b00111000; // 2518 :  56 - 0x38
      13'h9D7: dout  = 8'b00111100; // 2519 :  60 - 0x3c
      13'h9D8: dout  = 8'b00111100; // 2520 :  60 - 0x3c
      13'h9D9: dout  = 8'b10011000; // 2521 : 152 - 0x98
      13'h9DA: dout  = 8'b11000111; // 2522 : 199 - 0xc7
      13'h9DB: dout  = 8'b11001000; // 2523 : 200 - 0xc8
      13'h9DC: dout  = 8'b10010010; // 2524 : 146 - 0x92
      13'h9DD: dout  = 8'b00110000; // 2525 :  48 - 0x30
      13'h9DE: dout  = 8'b11111000; // 2526 : 248 - 0xf8
      13'h9DF: dout  = 8'b00111100; // 2527 :  60 - 0x3c
      13'h9E0: dout  = 8'b00000011; // 2528 :   3 - 0x3 -- Sprite 0x9e
      13'h9E1: dout  = 8'b00000111; // 2529 :   7 - 0x7
      13'h9E2: dout  = 8'b00001010; // 2530 :  10 - 0xa
      13'h9E3: dout  = 8'b00011010; // 2531 :  26 - 0x1a
      13'h9E4: dout  = 8'b00011100; // 2532 :  28 - 0x1c
      13'h9E5: dout  = 8'b00011110; // 2533 :  30 - 0x1e
      13'h9E6: dout  = 8'b00001011; // 2534 :  11 - 0xb
      13'h9E7: dout  = 8'b00001000; // 2535 :   8 - 0x8
      13'h9E8: dout  = 8'b00000000; // 2536 :   0 - 0x0
      13'h9E9: dout  = 8'b00010000; // 2537 :  16 - 0x10
      13'h9EA: dout  = 8'b01111111; // 2538 : 127 - 0x7f
      13'h9EB: dout  = 8'b01111111; // 2539 : 127 - 0x7f
      13'h9EC: dout  = 8'b01111111; // 2540 : 127 - 0x7f
      13'h9ED: dout  = 8'b00011111; // 2541 :  31 - 0x1f
      13'h9EE: dout  = 8'b00001111; // 2542 :  15 - 0xf
      13'h9EF: dout  = 8'b00001111; // 2543 :  15 - 0xf
      13'h9F0: dout  = 8'b00011100; // 2544 :  28 - 0x1c -- Sprite 0x9f
      13'h9F1: dout  = 8'b00111111; // 2545 :  63 - 0x3f
      13'h9F2: dout  = 8'b00111111; // 2546 :  63 - 0x3f
      13'h9F3: dout  = 8'b00111101; // 2547 :  61 - 0x3d
      13'h9F4: dout  = 8'b00111111; // 2548 :  63 - 0x3f
      13'h9F5: dout  = 8'b00011111; // 2549 :  31 - 0x1f
      13'h9F6: dout  = 8'b00000000; // 2550 :   0 - 0x0
      13'h9F7: dout  = 8'b00000000; // 2551 :   0 - 0x0
      13'h9F8: dout  = 8'b00000011; // 2552 :   3 - 0x3
      13'h9F9: dout  = 8'b00110011; // 2553 :  51 - 0x33
      13'h9FA: dout  = 8'b00111001; // 2554 :  57 - 0x39
      13'h9FB: dout  = 8'b00111010; // 2555 :  58 - 0x3a
      13'h9FC: dout  = 8'b00111000; // 2556 :  56 - 0x38
      13'h9FD: dout  = 8'b00011000; // 2557 :  24 - 0x18
      13'h9FE: dout  = 8'b00000000; // 2558 :   0 - 0x0
      13'h9FF: dout  = 8'b00000000; // 2559 :   0 - 0x0
      13'hA00: dout  = 8'b00000000; // 2560 :   0 - 0x0 -- Sprite 0xa0
      13'hA01: dout  = 8'b00000000; // 2561 :   0 - 0x0
      13'hA02: dout  = 8'b00000100; // 2562 :   4 - 0x4
      13'hA03: dout  = 8'b01001100; // 2563 :  76 - 0x4c
      13'hA04: dout  = 8'b01001110; // 2564 :  78 - 0x4e
      13'hA05: dout  = 8'b01001110; // 2565 :  78 - 0x4e
      13'hA06: dout  = 8'b01000110; // 2566 :  70 - 0x46
      13'hA07: dout  = 8'b01101111; // 2567 : 111 - 0x6f
      13'hA08: dout  = 8'b00010000; // 2568 :  16 - 0x10
      13'hA09: dout  = 8'b00111000; // 2569 :  56 - 0x38
      13'hA0A: dout  = 8'b00111100; // 2570 :  60 - 0x3c
      13'hA0B: dout  = 8'b01110100; // 2571 : 116 - 0x74
      13'hA0C: dout  = 8'b01110110; // 2572 : 118 - 0x76
      13'hA0D: dout  = 8'b01110110; // 2573 : 118 - 0x76
      13'hA0E: dout  = 8'b01111110; // 2574 : 126 - 0x7e
      13'hA0F: dout  = 8'b01111101; // 2575 : 125 - 0x7d
      13'hA10: dout  = 8'b00000000; // 2576 :   0 - 0x0 -- Sprite 0xa1
      13'hA11: dout  = 8'b00011111; // 2577 :  31 - 0x1f
      13'hA12: dout  = 8'b00111111; // 2578 :  63 - 0x3f
      13'hA13: dout  = 8'b00111111; // 2579 :  63 - 0x3f
      13'hA14: dout  = 8'b01001111; // 2580 :  79 - 0x4f
      13'hA15: dout  = 8'b01011111; // 2581 :  95 - 0x5f
      13'hA16: dout  = 8'b01111111; // 2582 : 127 - 0x7f
      13'hA17: dout  = 8'b01111111; // 2583 : 127 - 0x7f
      13'hA18: dout  = 8'b00000000; // 2584 :   0 - 0x0
      13'hA19: dout  = 8'b00000000; // 2585 :   0 - 0x0
      13'hA1A: dout  = 8'b00010001; // 2586 :  17 - 0x11
      13'hA1B: dout  = 8'b00001010; // 2587 :  10 - 0xa
      13'hA1C: dout  = 8'b00110100; // 2588 :  52 - 0x34
      13'hA1D: dout  = 8'b00101010; // 2589 :  42 - 0x2a
      13'hA1E: dout  = 8'b01010001; // 2590 :  81 - 0x51
      13'hA1F: dout  = 8'b00100000; // 2591 :  32 - 0x20
      13'hA20: dout  = 8'b01111111; // 2592 : 127 - 0x7f -- Sprite 0xa2
      13'hA21: dout  = 8'b01100111; // 2593 : 103 - 0x67
      13'hA22: dout  = 8'b10100011; // 2594 : 163 - 0xa3
      13'hA23: dout  = 8'b10110000; // 2595 : 176 - 0xb0
      13'hA24: dout  = 8'b11011000; // 2596 : 216 - 0xd8
      13'hA25: dout  = 8'b11011110; // 2597 : 222 - 0xde
      13'hA26: dout  = 8'b11011100; // 2598 : 220 - 0xdc
      13'hA27: dout  = 8'b11001000; // 2599 : 200 - 0xc8
      13'hA28: dout  = 8'b01111111; // 2600 : 127 - 0x7f
      13'hA29: dout  = 8'b01100111; // 2601 : 103 - 0x67
      13'hA2A: dout  = 8'b01100011; // 2602 :  99 - 0x63
      13'hA2B: dout  = 8'b01110000; // 2603 : 112 - 0x70
      13'hA2C: dout  = 8'b00111000; // 2604 :  56 - 0x38
      13'hA2D: dout  = 8'b00111110; // 2605 :  62 - 0x3e
      13'hA2E: dout  = 8'b01111100; // 2606 : 124 - 0x7c
      13'hA2F: dout  = 8'b10111000; // 2607 : 184 - 0xb8
      13'hA30: dout  = 8'b01111111; // 2608 : 127 - 0x7f -- Sprite 0xa3
      13'hA31: dout  = 8'b01111111; // 2609 : 127 - 0x7f
      13'hA32: dout  = 8'b01111111; // 2610 : 127 - 0x7f
      13'hA33: dout  = 8'b00011111; // 2611 :  31 - 0x1f
      13'hA34: dout  = 8'b01000111; // 2612 :  71 - 0x47
      13'hA35: dout  = 8'b01110000; // 2613 : 112 - 0x70
      13'hA36: dout  = 8'b01110000; // 2614 : 112 - 0x70
      13'hA37: dout  = 8'b00111001; // 2615 :  57 - 0x39
      13'hA38: dout  = 8'b01010001; // 2616 :  81 - 0x51
      13'hA39: dout  = 8'b00001010; // 2617 :  10 - 0xa
      13'hA3A: dout  = 8'b00000100; // 2618 :   4 - 0x4
      13'hA3B: dout  = 8'b11101010; // 2619 : 234 - 0xea
      13'hA3C: dout  = 8'b01111001; // 2620 : 121 - 0x79
      13'hA3D: dout  = 8'b01111111; // 2621 : 127 - 0x7f
      13'hA3E: dout  = 8'b01110000; // 2622 : 112 - 0x70
      13'hA3F: dout  = 8'b00111001; // 2623 :  57 - 0x39
      13'hA40: dout  = 8'b11101000; // 2624 : 232 - 0xe8 -- Sprite 0xa4
      13'hA41: dout  = 8'b11101000; // 2625 : 232 - 0xe8
      13'hA42: dout  = 8'b11100000; // 2626 : 224 - 0xe0
      13'hA43: dout  = 8'b11000000; // 2627 : 192 - 0xc0
      13'hA44: dout  = 8'b00010000; // 2628 :  16 - 0x10
      13'hA45: dout  = 8'b01110000; // 2629 : 112 - 0x70
      13'hA46: dout  = 8'b11100000; // 2630 : 224 - 0xe0
      13'hA47: dout  = 8'b11000000; // 2631 : 192 - 0xc0
      13'hA48: dout  = 8'b01011000; // 2632 :  88 - 0x58
      13'hA49: dout  = 8'b00111000; // 2633 :  56 - 0x38
      13'hA4A: dout  = 8'b00010000; // 2634 :  16 - 0x10
      13'hA4B: dout  = 8'b00110000; // 2635 :  48 - 0x30
      13'hA4C: dout  = 8'b11110000; // 2636 : 240 - 0xf0
      13'hA4D: dout  = 8'b11110000; // 2637 : 240 - 0xf0
      13'hA4E: dout  = 8'b11100000; // 2638 : 224 - 0xe0
      13'hA4F: dout  = 8'b11000000; // 2639 : 192 - 0xc0
      13'hA50: dout  = 8'b00000000; // 2640 :   0 - 0x0 -- Sprite 0xa5
      13'hA51: dout  = 8'b00000000; // 2641 :   0 - 0x0
      13'hA52: dout  = 8'b00000000; // 2642 :   0 - 0x0
      13'hA53: dout  = 8'b00100000; // 2643 :  32 - 0x20
      13'hA54: dout  = 8'b01100110; // 2644 : 102 - 0x66
      13'hA55: dout  = 8'b01100110; // 2645 : 102 - 0x66
      13'hA56: dout  = 8'b01100110; // 2646 : 102 - 0x66
      13'hA57: dout  = 8'b01100010; // 2647 :  98 - 0x62
      13'hA58: dout  = 8'b00000000; // 2648 :   0 - 0x0
      13'hA59: dout  = 8'b00001000; // 2649 :   8 - 0x8
      13'hA5A: dout  = 8'b00011100; // 2650 :  28 - 0x1c
      13'hA5B: dout  = 8'b00111100; // 2651 :  60 - 0x3c
      13'hA5C: dout  = 8'b01111010; // 2652 : 122 - 0x7a
      13'hA5D: dout  = 8'b01111010; // 2653 : 122 - 0x7a
      13'hA5E: dout  = 8'b01111010; // 2654 : 122 - 0x7a
      13'hA5F: dout  = 8'b01111110; // 2655 : 126 - 0x7e
      13'hA60: dout  = 8'b00000000; // 2656 :   0 - 0x0 -- Sprite 0xa6
      13'hA61: dout  = 8'b00000000; // 2657 :   0 - 0x0
      13'hA62: dout  = 8'b00011111; // 2658 :  31 - 0x1f
      13'hA63: dout  = 8'b00111111; // 2659 :  63 - 0x3f
      13'hA64: dout  = 8'b01111111; // 2660 : 127 - 0x7f
      13'hA65: dout  = 8'b01001111; // 2661 :  79 - 0x4f
      13'hA66: dout  = 8'b01011111; // 2662 :  95 - 0x5f
      13'hA67: dout  = 8'b01111111; // 2663 : 127 - 0x7f
      13'hA68: dout  = 8'b00000000; // 2664 :   0 - 0x0
      13'hA69: dout  = 8'b00000000; // 2665 :   0 - 0x0
      13'hA6A: dout  = 8'b00000000; // 2666 :   0 - 0x0
      13'hA6B: dout  = 8'b00010001; // 2667 :  17 - 0x11
      13'hA6C: dout  = 8'b00001010; // 2668 :  10 - 0xa
      13'hA6D: dout  = 8'b00110100; // 2669 :  52 - 0x34
      13'hA6E: dout  = 8'b00101010; // 2670 :  42 - 0x2a
      13'hA6F: dout  = 8'b01010001; // 2671 :  81 - 0x51
      13'hA70: dout  = 8'b01110111; // 2672 : 119 - 0x77 -- Sprite 0xa7
      13'hA71: dout  = 8'b01111111; // 2673 : 127 - 0x7f
      13'hA72: dout  = 8'b00111111; // 2674 :  63 - 0x3f
      13'hA73: dout  = 8'b10110111; // 2675 : 183 - 0xb7
      13'hA74: dout  = 8'b10110011; // 2676 : 179 - 0xb3
      13'hA75: dout  = 8'b11011011; // 2677 : 219 - 0xdb
      13'hA76: dout  = 8'b11011010; // 2678 : 218 - 0xda
      13'hA77: dout  = 8'b11011000; // 2679 : 216 - 0xd8
      13'hA78: dout  = 8'b01111111; // 2680 : 127 - 0x7f
      13'hA79: dout  = 8'b01111101; // 2681 : 125 - 0x7d
      13'hA7A: dout  = 8'b00111111; // 2682 :  63 - 0x3f
      13'hA7B: dout  = 8'b00110111; // 2683 :  55 - 0x37
      13'hA7C: dout  = 8'b00110011; // 2684 :  51 - 0x33
      13'hA7D: dout  = 8'b00111011; // 2685 :  59 - 0x3b
      13'hA7E: dout  = 8'b00111010; // 2686 :  58 - 0x3a
      13'hA7F: dout  = 8'b01111000; // 2687 : 120 - 0x78
      13'hA80: dout  = 8'b01111111; // 2688 : 127 - 0x7f -- Sprite 0xa8
      13'hA81: dout  = 8'b01111111; // 2689 : 127 - 0x7f
      13'hA82: dout  = 8'b01111111; // 2690 : 127 - 0x7f
      13'hA83: dout  = 8'b01111111; // 2691 : 127 - 0x7f
      13'hA84: dout  = 8'b00011111; // 2692 :  31 - 0x1f
      13'hA85: dout  = 8'b00000111; // 2693 :   7 - 0x7
      13'hA86: dout  = 8'b01110000; // 2694 : 112 - 0x70
      13'hA87: dout  = 8'b11110000; // 2695 : 240 - 0xf0
      13'hA88: dout  = 8'b00100000; // 2696 :  32 - 0x20
      13'hA89: dout  = 8'b01010001; // 2697 :  81 - 0x51
      13'hA8A: dout  = 8'b00001010; // 2698 :  10 - 0xa
      13'hA8B: dout  = 8'b00000100; // 2699 :   4 - 0x4
      13'hA8C: dout  = 8'b11101010; // 2700 : 234 - 0xea
      13'hA8D: dout  = 8'b00111001; // 2701 :  57 - 0x39
      13'hA8E: dout  = 8'b01111111; // 2702 : 127 - 0x7f
      13'hA8F: dout  = 8'b11110000; // 2703 : 240 - 0xf0
      13'hA90: dout  = 8'b11001100; // 2704 : 204 - 0xcc -- Sprite 0xa9
      13'hA91: dout  = 8'b11101000; // 2705 : 232 - 0xe8
      13'hA92: dout  = 8'b11101000; // 2706 : 232 - 0xe8
      13'hA93: dout  = 8'b11100000; // 2707 : 224 - 0xe0
      13'hA94: dout  = 8'b11000000; // 2708 : 192 - 0xc0
      13'hA95: dout  = 8'b00011000; // 2709 :  24 - 0x18
      13'hA96: dout  = 8'b01111100; // 2710 : 124 - 0x7c
      13'hA97: dout  = 8'b00111110; // 2711 :  62 - 0x3e
      13'hA98: dout  = 8'b10111100; // 2712 : 188 - 0xbc
      13'hA99: dout  = 8'b01011000; // 2713 :  88 - 0x58
      13'hA9A: dout  = 8'b00111000; // 2714 :  56 - 0x38
      13'hA9B: dout  = 8'b00010000; // 2715 :  16 - 0x10
      13'hA9C: dout  = 8'b00110000; // 2716 :  48 - 0x30
      13'hA9D: dout  = 8'b11111000; // 2717 : 248 - 0xf8
      13'hA9E: dout  = 8'b11111100; // 2718 : 252 - 0xfc
      13'hA9F: dout  = 8'b00111110; // 2719 :  62 - 0x3e
      13'hAA0: dout  = 8'b00000011; // 2720 :   3 - 0x3 -- Sprite 0xaa
      13'hAA1: dout  = 8'b00001111; // 2721 :  15 - 0xf
      13'hAA2: dout  = 8'b00011111; // 2722 :  31 - 0x1f
      13'hAA3: dout  = 8'b00111111; // 2723 :  63 - 0x3f
      13'hAA4: dout  = 8'b00111011; // 2724 :  59 - 0x3b
      13'hAA5: dout  = 8'b00111111; // 2725 :  63 - 0x3f
      13'hAA6: dout  = 8'b01111111; // 2726 : 127 - 0x7f
      13'hAA7: dout  = 8'b01111111; // 2727 : 127 - 0x7f
      13'hAA8: dout  = 8'b00000000; // 2728 :   0 - 0x0
      13'hAA9: dout  = 8'b00000000; // 2729 :   0 - 0x0
      13'hAAA: dout  = 8'b00000000; // 2730 :   0 - 0x0
      13'hAAB: dout  = 8'b00000110; // 2731 :   6 - 0x6
      13'hAAC: dout  = 8'b00001110; // 2732 :  14 - 0xe
      13'hAAD: dout  = 8'b00001100; // 2733 :  12 - 0xc
      13'hAAE: dout  = 8'b00000000; // 2734 :   0 - 0x0
      13'hAAF: dout  = 8'b00000000; // 2735 :   0 - 0x0
      13'hAB0: dout  = 8'b10000000; // 2736 : 128 - 0x80 -- Sprite 0xab
      13'hAB1: dout  = 8'b11110000; // 2737 : 240 - 0xf0
      13'hAB2: dout  = 8'b11111000; // 2738 : 248 - 0xf8
      13'hAB3: dout  = 8'b11111100; // 2739 : 252 - 0xfc
      13'hAB4: dout  = 8'b11111110; // 2740 : 254 - 0xfe
      13'hAB5: dout  = 8'b11111110; // 2741 : 254 - 0xfe
      13'hAB6: dout  = 8'b11111111; // 2742 : 255 - 0xff
      13'hAB7: dout  = 8'b11111110; // 2743 : 254 - 0xfe
      13'hAB8: dout  = 8'b00000000; // 2744 :   0 - 0x0
      13'hAB9: dout  = 8'b00000000; // 2745 :   0 - 0x0
      13'hABA: dout  = 8'b00000000; // 2746 :   0 - 0x0
      13'hABB: dout  = 8'b00000000; // 2747 :   0 - 0x0
      13'hABC: dout  = 8'b00000000; // 2748 :   0 - 0x0
      13'hABD: dout  = 8'b00000000; // 2749 :   0 - 0x0
      13'hABE: dout  = 8'b00001111; // 2750 :  15 - 0xf
      13'hABF: dout  = 8'b00011000; // 2751 :  24 - 0x18
      13'hAC0: dout  = 8'b01111111; // 2752 : 127 - 0x7f -- Sprite 0xac
      13'hAC1: dout  = 8'b01111111; // 2753 : 127 - 0x7f
      13'hAC2: dout  = 8'b01111111; // 2754 : 127 - 0x7f
      13'hAC3: dout  = 8'b01111111; // 2755 : 127 - 0x7f
      13'hAC4: dout  = 8'b11111111; // 2756 : 255 - 0xff
      13'hAC5: dout  = 8'b00001111; // 2757 :  15 - 0xf
      13'hAC6: dout  = 8'b00000011; // 2758 :   3 - 0x3
      13'hAC7: dout  = 8'b00000000; // 2759 :   0 - 0x0
      13'hAC8: dout  = 8'b00000000; // 2760 :   0 - 0x0
      13'hAC9: dout  = 8'b00000000; // 2761 :   0 - 0x0
      13'hACA: dout  = 8'b00000000; // 2762 :   0 - 0x0
      13'hACB: dout  = 8'b00000000; // 2763 :   0 - 0x0
      13'hACC: dout  = 8'b11111000; // 2764 : 248 - 0xf8
      13'hACD: dout  = 8'b00111110; // 2765 :  62 - 0x3e
      13'hACE: dout  = 8'b00111011; // 2766 :  59 - 0x3b
      13'hACF: dout  = 8'b00011000; // 2767 :  24 - 0x18
      13'hAD0: dout  = 8'b11111110; // 2768 : 254 - 0xfe -- Sprite 0xad
      13'hAD1: dout  = 8'b11111011; // 2769 : 251 - 0xfb
      13'hAD2: dout  = 8'b11111111; // 2770 : 255 - 0xff
      13'hAD3: dout  = 8'b11111111; // 2771 : 255 - 0xff
      13'hAD4: dout  = 8'b11110110; // 2772 : 246 - 0xf6
      13'hAD5: dout  = 8'b11100000; // 2773 : 224 - 0xe0
      13'hAD6: dout  = 8'b11000000; // 2774 : 192 - 0xc0
      13'hAD7: dout  = 8'b00000000; // 2775 :   0 - 0x0
      13'hAD8: dout  = 8'b00010000; // 2776 :  16 - 0x10
      13'hAD9: dout  = 8'b00010100; // 2777 :  20 - 0x14
      13'hADA: dout  = 8'b00010000; // 2778 :  16 - 0x10
      13'hADB: dout  = 8'b00010000; // 2779 :  16 - 0x10
      13'hADC: dout  = 8'b00111000; // 2780 :  56 - 0x38
      13'hADD: dout  = 8'b01111000; // 2781 : 120 - 0x78
      13'hADE: dout  = 8'b11111000; // 2782 : 248 - 0xf8
      13'hADF: dout  = 8'b00110000; // 2783 :  48 - 0x30
      13'hAE0: dout  = 8'b00000000; // 2784 :   0 - 0x0 -- Sprite 0xae
      13'hAE1: dout  = 8'b00000011; // 2785 :   3 - 0x3
      13'hAE2: dout  = 8'b00001111; // 2786 :  15 - 0xf
      13'hAE3: dout  = 8'b00011111; // 2787 :  31 - 0x1f
      13'hAE4: dout  = 8'b00111111; // 2788 :  63 - 0x3f
      13'hAE5: dout  = 8'b00111011; // 2789 :  59 - 0x3b
      13'hAE6: dout  = 8'b00111111; // 2790 :  63 - 0x3f
      13'hAE7: dout  = 8'b01111111; // 2791 : 127 - 0x7f
      13'hAE8: dout  = 8'b00000000; // 2792 :   0 - 0x0
      13'hAE9: dout  = 8'b00000000; // 2793 :   0 - 0x0
      13'hAEA: dout  = 8'b00000000; // 2794 :   0 - 0x0
      13'hAEB: dout  = 8'b00000000; // 2795 :   0 - 0x0
      13'hAEC: dout  = 8'b00000110; // 2796 :   6 - 0x6
      13'hAED: dout  = 8'b00001110; // 2797 :  14 - 0xe
      13'hAEE: dout  = 8'b00001100; // 2798 :  12 - 0xc
      13'hAEF: dout  = 8'b00000000; // 2799 :   0 - 0x0
      13'hAF0: dout  = 8'b00000000; // 2800 :   0 - 0x0 -- Sprite 0xaf
      13'hAF1: dout  = 8'b11000000; // 2801 : 192 - 0xc0
      13'hAF2: dout  = 8'b11110000; // 2802 : 240 - 0xf0
      13'hAF3: dout  = 8'b11111000; // 2803 : 248 - 0xf8
      13'hAF4: dout  = 8'b11111100; // 2804 : 252 - 0xfc
      13'hAF5: dout  = 8'b11111110; // 2805 : 254 - 0xfe
      13'hAF6: dout  = 8'b11111110; // 2806 : 254 - 0xfe
      13'hAF7: dout  = 8'b11111111; // 2807 : 255 - 0xff
      13'hAF8: dout  = 8'b00000000; // 2808 :   0 - 0x0
      13'hAF9: dout  = 8'b00000000; // 2809 :   0 - 0x0
      13'hAFA: dout  = 8'b00000000; // 2810 :   0 - 0x0
      13'hAFB: dout  = 8'b00000000; // 2811 :   0 - 0x0
      13'hAFC: dout  = 8'b00000000; // 2812 :   0 - 0x0
      13'hAFD: dout  = 8'b00000000; // 2813 :   0 - 0x0
      13'hAFE: dout  = 8'b00000000; // 2814 :   0 - 0x0
      13'hAFF: dout  = 8'b00001111; // 2815 :  15 - 0xf
      13'hB00: dout  = 8'b01111111; // 2816 : 127 - 0x7f -- Sprite 0xb0
      13'hB01: dout  = 8'b01111111; // 2817 : 127 - 0x7f
      13'hB02: dout  = 8'b01111111; // 2818 : 127 - 0x7f
      13'hB03: dout  = 8'b01111111; // 2819 : 127 - 0x7f
      13'hB04: dout  = 8'b01111111; // 2820 : 127 - 0x7f
      13'hB05: dout  = 8'b11111111; // 2821 : 255 - 0xff
      13'hB06: dout  = 8'b00001111; // 2822 :  15 - 0xf
      13'hB07: dout  = 8'b00000011; // 2823 :   3 - 0x3
      13'hB08: dout  = 8'b00000000; // 2824 :   0 - 0x0
      13'hB09: dout  = 8'b00000000; // 2825 :   0 - 0x0
      13'hB0A: dout  = 8'b00000000; // 2826 :   0 - 0x0
      13'hB0B: dout  = 8'b00000000; // 2827 :   0 - 0x0
      13'hB0C: dout  = 8'b00000000; // 2828 :   0 - 0x0
      13'hB0D: dout  = 8'b11111000; // 2829 : 248 - 0xf8
      13'hB0E: dout  = 8'b01111110; // 2830 : 126 - 0x7e
      13'hB0F: dout  = 8'b11110011; // 2831 : 243 - 0xf3
      13'hB10: dout  = 8'b11111110; // 2832 : 254 - 0xfe -- Sprite 0xb1
      13'hB11: dout  = 8'b11111110; // 2833 : 254 - 0xfe
      13'hB12: dout  = 8'b11111011; // 2834 : 251 - 0xfb
      13'hB13: dout  = 8'b11111111; // 2835 : 255 - 0xff
      13'hB14: dout  = 8'b11111111; // 2836 : 255 - 0xff
      13'hB15: dout  = 8'b11110110; // 2837 : 246 - 0xf6
      13'hB16: dout  = 8'b11100000; // 2838 : 224 - 0xe0
      13'hB17: dout  = 8'b11000000; // 2839 : 192 - 0xc0
      13'hB18: dout  = 8'b00011000; // 2840 :  24 - 0x18
      13'hB19: dout  = 8'b00010000; // 2841 :  16 - 0x10
      13'hB1A: dout  = 8'b00010100; // 2842 :  20 - 0x14
      13'hB1B: dout  = 8'b00010000; // 2843 :  16 - 0x10
      13'hB1C: dout  = 8'b00010000; // 2844 :  16 - 0x10
      13'hB1D: dout  = 8'b00111000; // 2845 :  56 - 0x38
      13'hB1E: dout  = 8'b01111100; // 2846 : 124 - 0x7c
      13'hB1F: dout  = 8'b11011110; // 2847 : 222 - 0xde
      13'hB20: dout  = 8'b00000000; // 2848 :   0 - 0x0 -- Sprite 0xb2
      13'hB21: dout  = 8'b00000001; // 2849 :   1 - 0x1
      13'hB22: dout  = 8'b00000001; // 2850 :   1 - 0x1
      13'hB23: dout  = 8'b00000001; // 2851 :   1 - 0x1
      13'hB24: dout  = 8'b00000001; // 2852 :   1 - 0x1
      13'hB25: dout  = 8'b00000000; // 2853 :   0 - 0x0
      13'hB26: dout  = 8'b00000000; // 2854 :   0 - 0x0
      13'hB27: dout  = 8'b00001000; // 2855 :   8 - 0x8
      13'hB28: dout  = 8'b00000000; // 2856 :   0 - 0x0
      13'hB29: dout  = 8'b00001101; // 2857 :  13 - 0xd
      13'hB2A: dout  = 8'b00011110; // 2858 :  30 - 0x1e
      13'hB2B: dout  = 8'b00011110; // 2859 :  30 - 0x1e
      13'hB2C: dout  = 8'b00011110; // 2860 :  30 - 0x1e
      13'hB2D: dout  = 8'b00011111; // 2861 :  31 - 0x1f
      13'hB2E: dout  = 8'b00001111; // 2862 :  15 - 0xf
      13'hB2F: dout  = 8'b00000111; // 2863 :   7 - 0x7
      13'hB30: dout  = 8'b01111000; // 2864 : 120 - 0x78 -- Sprite 0xb3
      13'hB31: dout  = 8'b11110000; // 2865 : 240 - 0xf0
      13'hB32: dout  = 8'b11111000; // 2866 : 248 - 0xf8
      13'hB33: dout  = 8'b11100100; // 2867 : 228 - 0xe4
      13'hB34: dout  = 8'b11000000; // 2868 : 192 - 0xc0
      13'hB35: dout  = 8'b11001010; // 2869 : 202 - 0xca
      13'hB36: dout  = 8'b11001010; // 2870 : 202 - 0xca
      13'hB37: dout  = 8'b11000000; // 2871 : 192 - 0xc0
      13'hB38: dout  = 8'b01111000; // 2872 : 120 - 0x78
      13'hB39: dout  = 8'b11110000; // 2873 : 240 - 0xf0
      13'hB3A: dout  = 8'b00000000; // 2874 :   0 - 0x0
      13'hB3B: dout  = 8'b00011010; // 2875 :  26 - 0x1a
      13'hB3C: dout  = 8'b00111111; // 2876 :  63 - 0x3f
      13'hB3D: dout  = 8'b00110101; // 2877 :  53 - 0x35
      13'hB3E: dout  = 8'b00110101; // 2878 :  53 - 0x35
      13'hB3F: dout  = 8'b00111111; // 2879 :  63 - 0x3f
      13'hB40: dout  = 8'b00001111; // 2880 :  15 - 0xf -- Sprite 0xb4
      13'hB41: dout  = 8'b00011111; // 2881 :  31 - 0x1f
      13'hB42: dout  = 8'b10011111; // 2882 : 159 - 0x9f
      13'hB43: dout  = 8'b11111111; // 2883 : 255 - 0xff
      13'hB44: dout  = 8'b11111111; // 2884 : 255 - 0xff
      13'hB45: dout  = 8'b01111111; // 2885 : 127 - 0x7f
      13'hB46: dout  = 8'b01110100; // 2886 : 116 - 0x74
      13'hB47: dout  = 8'b00100000; // 2887 :  32 - 0x20
      13'hB48: dout  = 8'b00000000; // 2888 :   0 - 0x0
      13'hB49: dout  = 8'b00000000; // 2889 :   0 - 0x0
      13'hB4A: dout  = 8'b10000000; // 2890 : 128 - 0x80
      13'hB4B: dout  = 8'b11100000; // 2891 : 224 - 0xe0
      13'hB4C: dout  = 8'b11100000; // 2892 : 224 - 0xe0
      13'hB4D: dout  = 8'b01110000; // 2893 : 112 - 0x70
      13'hB4E: dout  = 8'b01110011; // 2894 : 115 - 0x73
      13'hB4F: dout  = 8'b00100001; // 2895 :  33 - 0x21
      13'hB50: dout  = 8'b11100100; // 2896 : 228 - 0xe4 -- Sprite 0xb5
      13'hB51: dout  = 8'b11111111; // 2897 : 255 - 0xff
      13'hB52: dout  = 8'b11111110; // 2898 : 254 - 0xfe
      13'hB53: dout  = 8'b11111100; // 2899 : 252 - 0xfc
      13'hB54: dout  = 8'b10011100; // 2900 : 156 - 0x9c
      13'hB55: dout  = 8'b00011110; // 2901 :  30 - 0x1e
      13'hB56: dout  = 8'b00000000; // 2902 :   0 - 0x0
      13'hB57: dout  = 8'b00000000; // 2903 :   0 - 0x0
      13'hB58: dout  = 8'b00011010; // 2904 :  26 - 0x1a
      13'hB59: dout  = 8'b00000111; // 2905 :   7 - 0x7
      13'hB5A: dout  = 8'b00001100; // 2906 :  12 - 0xc
      13'hB5B: dout  = 8'b00011000; // 2907 :  24 - 0x18
      13'hB5C: dout  = 8'b01111000; // 2908 : 120 - 0x78
      13'hB5D: dout  = 8'b11111110; // 2909 : 254 - 0xfe
      13'hB5E: dout  = 8'b11111100; // 2910 : 252 - 0xfc
      13'hB5F: dout  = 8'b11110000; // 2911 : 240 - 0xf0
      13'hB60: dout  = 8'b00000000; // 2912 :   0 - 0x0 -- Sprite 0xb6
      13'hB61: dout  = 8'b00000001; // 2913 :   1 - 0x1
      13'hB62: dout  = 8'b00000011; // 2914 :   3 - 0x3
      13'hB63: dout  = 8'b00000011; // 2915 :   3 - 0x3
      13'hB64: dout  = 8'b00000111; // 2916 :   7 - 0x7
      13'hB65: dout  = 8'b00000011; // 2917 :   3 - 0x3
      13'hB66: dout  = 8'b00000001; // 2918 :   1 - 0x1
      13'hB67: dout  = 8'b00000000; // 2919 :   0 - 0x0
      13'hB68: dout  = 8'b00000000; // 2920 :   0 - 0x0
      13'hB69: dout  = 8'b00000001; // 2921 :   1 - 0x1
      13'hB6A: dout  = 8'b00000010; // 2922 :   2 - 0x2
      13'hB6B: dout  = 8'b00000000; // 2923 :   0 - 0x0
      13'hB6C: dout  = 8'b00111000; // 2924 :  56 - 0x38
      13'hB6D: dout  = 8'b01111100; // 2925 : 124 - 0x7c
      13'hB6E: dout  = 8'b01111110; // 2926 : 126 - 0x7e
      13'hB6F: dout  = 8'b00111111; // 2927 :  63 - 0x3f
      13'hB70: dout  = 8'b00000000; // 2928 :   0 - 0x0 -- Sprite 0xb7
      13'hB71: dout  = 8'b01011111; // 2929 :  95 - 0x5f
      13'hB72: dout  = 8'b01111111; // 2930 : 127 - 0x7f
      13'hB73: dout  = 8'b01111111; // 2931 : 127 - 0x7f
      13'hB74: dout  = 8'b00111111; // 2932 :  63 - 0x3f
      13'hB75: dout  = 8'b00111111; // 2933 :  63 - 0x3f
      13'hB76: dout  = 8'b00010100; // 2934 :  20 - 0x14
      13'hB77: dout  = 8'b00000000; // 2935 :   0 - 0x0
      13'hB78: dout  = 8'b00111111; // 2936 :  63 - 0x3f
      13'hB79: dout  = 8'b01000000; // 2937 :  64 - 0x40
      13'hB7A: dout  = 8'b01100000; // 2938 :  96 - 0x60
      13'hB7B: dout  = 8'b01100000; // 2939 :  96 - 0x60
      13'hB7C: dout  = 8'b00100000; // 2940 :  32 - 0x20
      13'hB7D: dout  = 8'b00110000; // 2941 :  48 - 0x30
      13'hB7E: dout  = 8'b00010011; // 2942 :  19 - 0x13
      13'hB7F: dout  = 8'b00000001; // 2943 :   1 - 0x1
      13'hB80: dout  = 8'b11000000; // 2944 : 192 - 0xc0 -- Sprite 0xb8
      13'hB81: dout  = 8'b11100000; // 2945 : 224 - 0xe0
      13'hB82: dout  = 8'b11110000; // 2946 : 240 - 0xf0
      13'hB83: dout  = 8'b00110000; // 2947 :  48 - 0x30
      13'hB84: dout  = 8'b00111000; // 2948 :  56 - 0x38
      13'hB85: dout  = 8'b00111100; // 2949 :  60 - 0x3c
      13'hB86: dout  = 8'b00111100; // 2950 :  60 - 0x3c
      13'hB87: dout  = 8'b11111100; // 2951 : 252 - 0xfc
      13'hB88: dout  = 8'b11000000; // 2952 : 192 - 0xc0
      13'hB89: dout  = 8'b11100000; // 2953 : 224 - 0xe0
      13'hB8A: dout  = 8'b00110000; // 2954 :  48 - 0x30
      13'hB8B: dout  = 8'b11010000; // 2955 : 208 - 0xd0
      13'hB8C: dout  = 8'b11010000; // 2956 : 208 - 0xd0
      13'hB8D: dout  = 8'b11010000; // 2957 : 208 - 0xd0
      13'hB8E: dout  = 8'b11010000; // 2958 : 208 - 0xd0
      13'hB8F: dout  = 8'b00000000; // 2959 :   0 - 0x0
      13'hB90: dout  = 8'b00000111; // 2960 :   7 - 0x7 -- Sprite 0xb9
      13'hB91: dout  = 8'b00001111; // 2961 :  15 - 0xf
      13'hB92: dout  = 8'b00011111; // 2962 :  31 - 0x1f
      13'hB93: dout  = 8'b00100010; // 2963 :  34 - 0x22
      13'hB94: dout  = 8'b00100000; // 2964 :  32 - 0x20
      13'hB95: dout  = 8'b00100101; // 2965 :  37 - 0x25
      13'hB96: dout  = 8'b00100101; // 2966 :  37 - 0x25
      13'hB97: dout  = 8'b00011111; // 2967 :  31 - 0x1f
      13'hB98: dout  = 8'b00000111; // 2968 :   7 - 0x7
      13'hB99: dout  = 8'b00001111; // 2969 :  15 - 0xf
      13'hB9A: dout  = 8'b00000010; // 2970 :   2 - 0x2
      13'hB9B: dout  = 8'b00011101; // 2971 :  29 - 0x1d
      13'hB9C: dout  = 8'b00011111; // 2972 :  31 - 0x1f
      13'hB9D: dout  = 8'b00011010; // 2973 :  26 - 0x1a
      13'hB9E: dout  = 8'b00011010; // 2974 :  26 - 0x1a
      13'hB9F: dout  = 8'b00000010; // 2975 :   2 - 0x2
      13'hBA0: dout  = 8'b11111110; // 2976 : 254 - 0xfe -- Sprite 0xba
      13'hBA1: dout  = 8'b11111110; // 2977 : 254 - 0xfe
      13'hBA2: dout  = 8'b01111110; // 2978 : 126 - 0x7e
      13'hBA3: dout  = 8'b00111010; // 2979 :  58 - 0x3a
      13'hBA4: dout  = 8'b00000010; // 2980 :   2 - 0x2
      13'hBA5: dout  = 8'b00000001; // 2981 :   1 - 0x1
      13'hBA6: dout  = 8'b01000001; // 2982 :  65 - 0x41
      13'hBA7: dout  = 8'b01000001; // 2983 :  65 - 0x41
      13'hBA8: dout  = 8'b00111000; // 2984 :  56 - 0x38
      13'hBA9: dout  = 8'b01111100; // 2985 : 124 - 0x7c
      13'hBAA: dout  = 8'b11111100; // 2986 : 252 - 0xfc
      13'hBAB: dout  = 8'b11111100; // 2987 : 252 - 0xfc
      13'hBAC: dout  = 8'b11111100; // 2988 : 252 - 0xfc
      13'hBAD: dout  = 8'b11111110; // 2989 : 254 - 0xfe
      13'hBAE: dout  = 8'b10111110; // 2990 : 190 - 0xbe
      13'hBAF: dout  = 8'b10111110; // 2991 : 190 - 0xbe
      13'hBB0: dout  = 8'b00011111; // 2992 :  31 - 0x1f -- Sprite 0xbb
      13'hBB1: dout  = 8'b00111111; // 2993 :  63 - 0x3f
      13'hBB2: dout  = 8'b01111110; // 2994 : 126 - 0x7e
      13'hBB3: dout  = 8'b01011100; // 2995 :  92 - 0x5c
      13'hBB4: dout  = 8'b01000000; // 2996 :  64 - 0x40
      13'hBB5: dout  = 8'b10000000; // 2997 : 128 - 0x80
      13'hBB6: dout  = 8'b10000010; // 2998 : 130 - 0x82
      13'hBB7: dout  = 8'b10000010; // 2999 : 130 - 0x82
      13'hBB8: dout  = 8'b00011100; // 3000 :  28 - 0x1c
      13'hBB9: dout  = 8'b00111110; // 3001 :  62 - 0x3e
      13'hBBA: dout  = 8'b00111111; // 3002 :  63 - 0x3f
      13'hBBB: dout  = 8'b00111111; // 3003 :  63 - 0x3f
      13'hBBC: dout  = 8'b00111111; // 3004 :  63 - 0x3f
      13'hBBD: dout  = 8'b01111111; // 3005 : 127 - 0x7f
      13'hBBE: dout  = 8'b01111101; // 3006 : 125 - 0x7d
      13'hBBF: dout  = 8'b01111101; // 3007 : 125 - 0x7d
      13'hBC0: dout  = 8'b10000010; // 3008 : 130 - 0x82 -- Sprite 0xbc
      13'hBC1: dout  = 8'b10000000; // 3009 : 128 - 0x80
      13'hBC2: dout  = 8'b10100000; // 3010 : 160 - 0xa0
      13'hBC3: dout  = 8'b01000100; // 3011 :  68 - 0x44
      13'hBC4: dout  = 8'b01000011; // 3012 :  67 - 0x43
      13'hBC5: dout  = 8'b01000000; // 3013 :  64 - 0x40
      13'hBC6: dout  = 8'b00100001; // 3014 :  33 - 0x21
      13'hBC7: dout  = 8'b00011110; // 3015 :  30 - 0x1e
      13'hBC8: dout  = 8'b01111101; // 3016 : 125 - 0x7d
      13'hBC9: dout  = 8'b01111111; // 3017 : 127 - 0x7f
      13'hBCA: dout  = 8'b01011111; // 3018 :  95 - 0x5f
      13'hBCB: dout  = 8'b00111011; // 3019 :  59 - 0x3b
      13'hBCC: dout  = 8'b00111100; // 3020 :  60 - 0x3c
      13'hBCD: dout  = 8'b00111111; // 3021 :  63 - 0x3f
      13'hBCE: dout  = 8'b00011110; // 3022 :  30 - 0x1e
      13'hBCF: dout  = 8'b00000000; // 3023 :   0 - 0x0
      13'hBD0: dout  = 8'b00011100; // 3024 :  28 - 0x1c -- Sprite 0xbd
      13'hBD1: dout  = 8'b00111111; // 3025 :  63 - 0x3f
      13'hBD2: dout  = 8'b00111110; // 3026 :  62 - 0x3e
      13'hBD3: dout  = 8'b00111100; // 3027 :  60 - 0x3c
      13'hBD4: dout  = 8'b01000000; // 3028 :  64 - 0x40
      13'hBD5: dout  = 8'b10000000; // 3029 : 128 - 0x80
      13'hBD6: dout  = 8'b10000010; // 3030 : 130 - 0x82
      13'hBD7: dout  = 8'b10000010; // 3031 : 130 - 0x82
      13'hBD8: dout  = 8'b00011100; // 3032 :  28 - 0x1c
      13'hBD9: dout  = 8'b00111110; // 3033 :  62 - 0x3e
      13'hBDA: dout  = 8'b00111111; // 3034 :  63 - 0x3f
      13'hBDB: dout  = 8'b00011111; // 3035 :  31 - 0x1f
      13'hBDC: dout  = 8'b00111111; // 3036 :  63 - 0x3f
      13'hBDD: dout  = 8'b01111111; // 3037 : 127 - 0x7f
      13'hBDE: dout  = 8'b01111101; // 3038 : 125 - 0x7d
      13'hBDF: dout  = 8'b01111101; // 3039 : 125 - 0x7d
      13'hBE0: dout  = 8'b00000000; // 3040 :   0 - 0x0 -- Sprite 0xbe
      13'hBE1: dout  = 8'b00000000; // 3041 :   0 - 0x0
      13'hBE2: dout  = 8'b10000000; // 3042 : 128 - 0x80
      13'hBE3: dout  = 8'b10000000; // 3043 : 128 - 0x80
      13'hBE4: dout  = 8'b10010010; // 3044 : 146 - 0x92
      13'hBE5: dout  = 8'b10011101; // 3045 : 157 - 0x9d
      13'hBE6: dout  = 8'b11000111; // 3046 : 199 - 0xc7
      13'hBE7: dout  = 8'b11101111; // 3047 : 239 - 0xef
      13'hBE8: dout  = 8'b00000000; // 3048 :   0 - 0x0
      13'hBE9: dout  = 8'b00000000; // 3049 :   0 - 0x0
      13'hBEA: dout  = 8'b00000000; // 3050 :   0 - 0x0
      13'hBEB: dout  = 8'b01100000; // 3051 :  96 - 0x60
      13'hBEC: dout  = 8'b01100010; // 3052 :  98 - 0x62
      13'hBED: dout  = 8'b01100101; // 3053 : 101 - 0x65
      13'hBEE: dout  = 8'b00111111; // 3054 :  63 - 0x3f
      13'hBEF: dout  = 8'b00011111; // 3055 :  31 - 0x1f
      13'hBF0: dout  = 8'b00000000; // 3056 :   0 - 0x0 -- Sprite 0xbf
      13'hBF1: dout  = 8'b00100011; // 3057 :  35 - 0x23
      13'hBF2: dout  = 8'b00110011; // 3058 :  51 - 0x33
      13'hBF3: dout  = 8'b00111111; // 3059 :  63 - 0x3f
      13'hBF4: dout  = 8'b00111111; // 3060 :  63 - 0x3f
      13'hBF5: dout  = 8'b01111111; // 3061 : 127 - 0x7f
      13'hBF6: dout  = 8'b01111111; // 3062 : 127 - 0x7f
      13'hBF7: dout  = 8'b01111111; // 3063 : 127 - 0x7f
      13'hBF8: dout  = 8'b01110000; // 3064 : 112 - 0x70
      13'hBF9: dout  = 8'b00111100; // 3065 :  60 - 0x3c
      13'hBFA: dout  = 8'b00111100; // 3066 :  60 - 0x3c
      13'hBFB: dout  = 8'b00011000; // 3067 :  24 - 0x18
      13'hBFC: dout  = 8'b00000000; // 3068 :   0 - 0x0
      13'hBFD: dout  = 8'b00000000; // 3069 :   0 - 0x0
      13'hBFE: dout  = 8'b00000010; // 3070 :   2 - 0x2
      13'hBFF: dout  = 8'b00000111; // 3071 :   7 - 0x7
      13'hC00: dout  = 8'b11111110; // 3072 : 254 - 0xfe -- Sprite 0xc0
      13'hC01: dout  = 8'b11111000; // 3073 : 248 - 0xf8
      13'hC02: dout  = 8'b10100000; // 3074 : 160 - 0xa0
      13'hC03: dout  = 8'b00000000; // 3075 :   0 - 0x0
      13'hC04: dout  = 8'b00000000; // 3076 :   0 - 0x0
      13'hC05: dout  = 8'b00000000; // 3077 :   0 - 0x0
      13'hC06: dout  = 8'b10000000; // 3078 : 128 - 0x80
      13'hC07: dout  = 8'b10000000; // 3079 : 128 - 0x80
      13'hC08: dout  = 8'b11001111; // 3080 : 207 - 0xcf
      13'hC09: dout  = 8'b01111010; // 3081 : 122 - 0x7a
      13'hC0A: dout  = 8'b01011010; // 3082 :  90 - 0x5a
      13'hC0B: dout  = 8'b00010000; // 3083 :  16 - 0x10
      13'hC0C: dout  = 8'b00000000; // 3084 :   0 - 0x0
      13'hC0D: dout  = 8'b00000000; // 3085 :   0 - 0x0
      13'hC0E: dout  = 8'b11000000; // 3086 : 192 - 0xc0
      13'hC0F: dout  = 8'b10000000; // 3087 : 128 - 0x80
      13'hC10: dout  = 8'b01111110; // 3088 : 126 - 0x7e -- Sprite 0xc1
      13'hC11: dout  = 8'b01111111; // 3089 : 127 - 0x7f
      13'hC12: dout  = 8'b01111101; // 3090 : 125 - 0x7d
      13'hC13: dout  = 8'b00111111; // 3091 :  63 - 0x3f
      13'hC14: dout  = 8'b00011110; // 3092 :  30 - 0x1e
      13'hC15: dout  = 8'b10001111; // 3093 : 143 - 0x8f
      13'hC16: dout  = 8'b10001111; // 3094 : 143 - 0x8f
      13'hC17: dout  = 8'b00011001; // 3095 :  25 - 0x19
      13'hC18: dout  = 8'b10000101; // 3096 : 133 - 0x85
      13'hC19: dout  = 8'b10000100; // 3097 : 132 - 0x84
      13'hC1A: dout  = 8'b10000110; // 3098 : 134 - 0x86
      13'hC1B: dout  = 8'b11000110; // 3099 : 198 - 0xc6
      13'hC1C: dout  = 8'b11100111; // 3100 : 231 - 0xe7
      13'hC1D: dout  = 8'b01110011; // 3101 : 115 - 0x73
      13'hC1E: dout  = 8'b01110011; // 3102 : 115 - 0x73
      13'hC1F: dout  = 8'b11100001; // 3103 : 225 - 0xe1
      13'hC20: dout  = 8'b11100000; // 3104 : 224 - 0xe0 -- Sprite 0xc2
      13'hC21: dout  = 8'b00001110; // 3105 :  14 - 0xe
      13'hC22: dout  = 8'b01110011; // 3106 : 115 - 0x73
      13'hC23: dout  = 8'b11110011; // 3107 : 243 - 0xf3
      13'hC24: dout  = 8'b11111001; // 3108 : 249 - 0xf9
      13'hC25: dout  = 8'b11111001; // 3109 : 249 - 0xf9
      13'hC26: dout  = 8'b11111000; // 3110 : 248 - 0xf8
      13'hC27: dout  = 8'b01110000; // 3111 : 112 - 0x70
      13'hC28: dout  = 8'b10000000; // 3112 : 128 - 0x80
      13'hC29: dout  = 8'b01001110; // 3113 :  78 - 0x4e
      13'hC2A: dout  = 8'b01110111; // 3114 : 119 - 0x77
      13'hC2B: dout  = 8'b11110011; // 3115 : 243 - 0xf3
      13'hC2C: dout  = 8'b11111011; // 3116 : 251 - 0xfb
      13'hC2D: dout  = 8'b11111001; // 3117 : 249 - 0xf9
      13'hC2E: dout  = 8'b11111010; // 3118 : 250 - 0xfa
      13'hC2F: dout  = 8'b01111000; // 3119 : 120 - 0x78
      13'hC30: dout  = 8'b00001110; // 3120 :  14 - 0xe -- Sprite 0xc3
      13'hC31: dout  = 8'b01100110; // 3121 : 102 - 0x66
      13'hC32: dout  = 8'b11100010; // 3122 : 226 - 0xe2
      13'hC33: dout  = 8'b11110110; // 3123 : 246 - 0xf6
      13'hC34: dout  = 8'b11111111; // 3124 : 255 - 0xff
      13'hC35: dout  = 8'b11111111; // 3125 : 255 - 0xff
      13'hC36: dout  = 8'b00011111; // 3126 :  31 - 0x1f
      13'hC37: dout  = 8'b10011000; // 3127 : 152 - 0x98
      13'hC38: dout  = 8'b00010001; // 3128 :  17 - 0x11
      13'hC39: dout  = 8'b00111001; // 3129 :  57 - 0x39
      13'hC3A: dout  = 8'b01111101; // 3130 : 125 - 0x7d
      13'hC3B: dout  = 8'b00111001; // 3131 :  57 - 0x39
      13'hC3C: dout  = 8'b00000000; // 3132 :   0 - 0x0
      13'hC3D: dout  = 8'b00000000; // 3133 :   0 - 0x0
      13'hC3E: dout  = 8'b11100000; // 3134 : 224 - 0xe0
      13'hC3F: dout  = 8'b11100111; // 3135 : 231 - 0xe7
      13'hC40: dout  = 8'b00000000; // 3136 :   0 - 0x0 -- Sprite 0xc4
      13'hC41: dout  = 8'b00000000; // 3137 :   0 - 0x0
      13'hC42: dout  = 8'b00000000; // 3138 :   0 - 0x0
      13'hC43: dout  = 8'b00000100; // 3139 :   4 - 0x4
      13'hC44: dout  = 8'b00001111; // 3140 :  15 - 0xf
      13'hC45: dout  = 8'b00001111; // 3141 :  15 - 0xf
      13'hC46: dout  = 8'b00011111; // 3142 :  31 - 0x1f
      13'hC47: dout  = 8'b00000111; // 3143 :   7 - 0x7
      13'hC48: dout  = 8'b00000000; // 3144 :   0 - 0x0
      13'hC49: dout  = 8'b00000000; // 3145 :   0 - 0x0
      13'hC4A: dout  = 8'b00000111; // 3146 :   7 - 0x7
      13'hC4B: dout  = 8'b00000111; // 3147 :   7 - 0x7
      13'hC4C: dout  = 8'b00010110; // 3148 :  22 - 0x16
      13'hC4D: dout  = 8'b00010000; // 3149 :  16 - 0x10
      13'hC4E: dout  = 8'b00000000; // 3150 :   0 - 0x0
      13'hC4F: dout  = 8'b00111000; // 3151 :  56 - 0x38
      13'hC50: dout  = 8'b11110011; // 3152 : 243 - 0xf3 -- Sprite 0xc5
      13'hC51: dout  = 8'b11100111; // 3153 : 231 - 0xe7
      13'hC52: dout  = 8'b11101110; // 3154 : 238 - 0xee
      13'hC53: dout  = 8'b11101100; // 3155 : 236 - 0xec
      13'hC54: dout  = 8'b11001101; // 3156 : 205 - 0xcd
      13'hC55: dout  = 8'b11001111; // 3157 : 207 - 0xcf
      13'hC56: dout  = 8'b11001111; // 3158 : 207 - 0xcf
      13'hC57: dout  = 8'b11011111; // 3159 : 223 - 0xdf
      13'hC58: dout  = 8'b11001111; // 3160 : 207 - 0xcf
      13'hC59: dout  = 8'b00011111; // 3161 :  31 - 0x1f
      13'hC5A: dout  = 8'b00010111; // 3162 :  23 - 0x17
      13'hC5B: dout  = 8'b00010000; // 3163 :  16 - 0x10
      13'hC5C: dout  = 8'b00110011; // 3164 :  51 - 0x33
      13'hC5D: dout  = 8'b00110000; // 3165 :  48 - 0x30
      13'hC5E: dout  = 8'b00110000; // 3166 :  48 - 0x30
      13'hC5F: dout  = 8'b00100000; // 3167 :  32 - 0x20
      13'hC60: dout  = 8'b00100111; // 3168 :  39 - 0x27 -- Sprite 0xc6
      13'hC61: dout  = 8'b00111111; // 3169 :  63 - 0x3f
      13'hC62: dout  = 8'b00111111; // 3170 :  63 - 0x3f
      13'hC63: dout  = 8'b01111000; // 3171 : 120 - 0x78
      13'hC64: dout  = 8'b00111100; // 3172 :  60 - 0x3c
      13'hC65: dout  = 8'b00011111; // 3173 :  31 - 0x1f
      13'hC66: dout  = 8'b00011111; // 3174 :  31 - 0x1f
      13'hC67: dout  = 8'b01110011; // 3175 : 115 - 0x73
      13'hC68: dout  = 8'b00111000; // 3176 :  56 - 0x38
      13'hC69: dout  = 8'b00110000; // 3177 :  48 - 0x30
      13'hC6A: dout  = 8'b01000000; // 3178 :  64 - 0x40
      13'hC6B: dout  = 8'b11000111; // 3179 : 199 - 0xc7
      13'hC6C: dout  = 8'b00000111; // 3180 :   7 - 0x7
      13'hC6D: dout  = 8'b01100110; // 3181 : 102 - 0x66
      13'hC6E: dout  = 8'b11100000; // 3182 : 224 - 0xe0
      13'hC6F: dout  = 8'b01101100; // 3183 : 108 - 0x6c
      13'hC70: dout  = 8'b10011111; // 3184 : 159 - 0x9f -- Sprite 0xc7
      13'hC71: dout  = 8'b00111110; // 3185 :  62 - 0x3e
      13'hC72: dout  = 8'b01111100; // 3186 : 124 - 0x7c
      13'hC73: dout  = 8'b11111100; // 3187 : 252 - 0xfc
      13'hC74: dout  = 8'b11111000; // 3188 : 248 - 0xf8
      13'hC75: dout  = 8'b11111000; // 3189 : 248 - 0xf8
      13'hC76: dout  = 8'b11000000; // 3190 : 192 - 0xc0
      13'hC77: dout  = 8'b01000000; // 3191 :  64 - 0x40
      13'hC78: dout  = 8'b01100000; // 3192 :  96 - 0x60
      13'hC79: dout  = 8'b11000000; // 3193 : 192 - 0xc0
      13'hC7A: dout  = 8'b10000000; // 3194 : 128 - 0x80
      13'hC7B: dout  = 8'b00000100; // 3195 :   4 - 0x4
      13'hC7C: dout  = 8'b10011110; // 3196 : 158 - 0x9e
      13'hC7D: dout  = 8'b11111111; // 3197 : 255 - 0xff
      13'hC7E: dout  = 8'b11110000; // 3198 : 240 - 0xf0
      13'hC7F: dout  = 8'b11111000; // 3199 : 248 - 0xf8
      13'hC80: dout  = 8'b01111111; // 3200 : 127 - 0x7f -- Sprite 0xc8
      13'hC81: dout  = 8'b01111110; // 3201 : 126 - 0x7e
      13'hC82: dout  = 8'b01111000; // 3202 : 120 - 0x78
      13'hC83: dout  = 8'b00000001; // 3203 :   1 - 0x1
      13'hC84: dout  = 8'b00000111; // 3204 :   7 - 0x7
      13'hC85: dout  = 8'b00011111; // 3205 :  31 - 0x1f
      13'hC86: dout  = 8'b00111100; // 3206 :  60 - 0x3c
      13'hC87: dout  = 8'b01111100; // 3207 : 124 - 0x7c
      13'hC88: dout  = 8'b00100100; // 3208 :  36 - 0x24
      13'hC89: dout  = 8'b00000001; // 3209 :   1 - 0x1
      13'hC8A: dout  = 8'b00000111; // 3210 :   7 - 0x7
      13'hC8B: dout  = 8'b11111110; // 3211 : 254 - 0xfe
      13'hC8C: dout  = 8'b11111111; // 3212 : 255 - 0xff
      13'hC8D: dout  = 8'b01111111; // 3213 : 127 - 0x7f
      13'hC8E: dout  = 8'b00111111; // 3214 :  63 - 0x3f
      13'hC8F: dout  = 8'b01111111; // 3215 : 127 - 0x7f
      13'hC90: dout  = 8'b11111100; // 3216 : 252 - 0xfc -- Sprite 0xc9
      13'hC91: dout  = 8'b11111000; // 3217 : 248 - 0xf8
      13'hC92: dout  = 8'b10100000; // 3218 : 160 - 0xa0
      13'hC93: dout  = 8'b11111110; // 3219 : 254 - 0xfe
      13'hC94: dout  = 8'b11111100; // 3220 : 252 - 0xfc
      13'hC95: dout  = 8'b11110000; // 3221 : 240 - 0xf0
      13'hC96: dout  = 8'b10000000; // 3222 : 128 - 0x80
      13'hC97: dout  = 8'b00000000; // 3223 :   0 - 0x0
      13'hC98: dout  = 8'b11001111; // 3224 : 207 - 0xcf
      13'hC99: dout  = 8'b01111010; // 3225 : 122 - 0x7a
      13'hC9A: dout  = 8'b00001010; // 3226 :  10 - 0xa
      13'hC9B: dout  = 8'b11111110; // 3227 : 254 - 0xfe
      13'hC9C: dout  = 8'b11111100; // 3228 : 252 - 0xfc
      13'hC9D: dout  = 8'b00000000; // 3229 :   0 - 0x0
      13'hC9E: dout  = 8'b00000000; // 3230 :   0 - 0x0
      13'hC9F: dout  = 8'b00000000; // 3231 :   0 - 0x0
      13'hCA0: dout  = 8'b01111110; // 3232 : 126 - 0x7e -- Sprite 0xca
      13'hCA1: dout  = 8'b01111111; // 3233 : 127 - 0x7f
      13'hCA2: dout  = 8'b01111111; // 3234 : 127 - 0x7f
      13'hCA3: dout  = 8'b00111111; // 3235 :  63 - 0x3f
      13'hCA4: dout  = 8'b00011111; // 3236 :  31 - 0x1f
      13'hCA5: dout  = 8'b10001111; // 3237 : 143 - 0x8f
      13'hCA6: dout  = 8'b10001111; // 3238 : 143 - 0x8f
      13'hCA7: dout  = 8'b00011000; // 3239 :  24 - 0x18
      13'hCA8: dout  = 8'b10000101; // 3240 : 133 - 0x85
      13'hCA9: dout  = 8'b10000110; // 3241 : 134 - 0x86
      13'hCAA: dout  = 8'b10000011; // 3242 : 131 - 0x83
      13'hCAB: dout  = 8'b11000011; // 3243 : 195 - 0xc3
      13'hCAC: dout  = 8'b11100001; // 3244 : 225 - 0xe1
      13'hCAD: dout  = 8'b01110000; // 3245 : 112 - 0x70
      13'hCAE: dout  = 8'b01110000; // 3246 : 112 - 0x70
      13'hCAF: dout  = 8'b11100000; // 3247 : 224 - 0xe0
      13'hCB0: dout  = 8'b10011111; // 3248 : 159 - 0x9f -- Sprite 0xcb
      13'hCB1: dout  = 8'b00111110; // 3249 :  62 - 0x3e
      13'hCB2: dout  = 8'b01111100; // 3250 : 124 - 0x7c
      13'hCB3: dout  = 8'b11111000; // 3251 : 248 - 0xf8
      13'hCB4: dout  = 8'b11111000; // 3252 : 248 - 0xf8
      13'hCB5: dout  = 8'b00111100; // 3253 :  60 - 0x3c
      13'hCB6: dout  = 8'b00011000; // 3254 :  24 - 0x18
      13'hCB7: dout  = 8'b11111000; // 3255 : 248 - 0xf8
      13'hCB8: dout  = 8'b01100000; // 3256 :  96 - 0x60
      13'hCB9: dout  = 8'b11000000; // 3257 : 192 - 0xc0
      13'hCBA: dout  = 8'b10000000; // 3258 : 128 - 0x80
      13'hCBB: dout  = 8'b00000000; // 3259 :   0 - 0x0
      13'hCBC: dout  = 8'b10011000; // 3260 : 152 - 0x98
      13'hCBD: dout  = 8'b11111100; // 3261 : 252 - 0xfc
      13'hCBE: dout  = 8'b11111110; // 3262 : 254 - 0xfe
      13'hCBF: dout  = 8'b11111111; // 3263 : 255 - 0xff
      13'hCC0: dout  = 8'b01111111; // 3264 : 127 - 0x7f -- Sprite 0xcc
      13'hCC1: dout  = 8'b01111111; // 3265 : 127 - 0x7f
      13'hCC2: dout  = 8'b01111000; // 3266 : 120 - 0x78
      13'hCC3: dout  = 8'b00000001; // 3267 :   1 - 0x1
      13'hCC4: dout  = 8'b00000111; // 3268 :   7 - 0x7
      13'hCC5: dout  = 8'b00010011; // 3269 :  19 - 0x13
      13'hCC6: dout  = 8'b11110001; // 3270 : 241 - 0xf1
      13'hCC7: dout  = 8'b00000011; // 3271 :   3 - 0x3
      13'hCC8: dout  = 8'b00100100; // 3272 :  36 - 0x24
      13'hCC9: dout  = 8'b00000000; // 3273 :   0 - 0x0
      13'hCCA: dout  = 8'b00000111; // 3274 :   7 - 0x7
      13'hCCB: dout  = 8'b11111110; // 3275 : 254 - 0xfe
      13'hCCC: dout  = 8'b11111111; // 3276 : 255 - 0xff
      13'hCCD: dout  = 8'b01111111; // 3277 : 127 - 0x7f
      13'hCCE: dout  = 8'b11111111; // 3278 : 255 - 0xff
      13'hCCF: dout  = 8'b00000011; // 3279 :   3 - 0x3
      13'hCD0: dout  = 8'b00000000; // 3280 :   0 - 0x0 -- Sprite 0xcd
      13'hCD1: dout  = 8'b00000000; // 3281 :   0 - 0x0
      13'hCD2: dout  = 8'b00011100; // 3282 :  28 - 0x1c
      13'hCD3: dout  = 8'b00011101; // 3283 :  29 - 0x1d
      13'hCD4: dout  = 8'b00011011; // 3284 :  27 - 0x1b
      13'hCD5: dout  = 8'b11000011; // 3285 : 195 - 0xc3
      13'hCD6: dout  = 8'b11100011; // 3286 : 227 - 0xe3
      13'hCD7: dout  = 8'b11100001; // 3287 : 225 - 0xe1
      13'hCD8: dout  = 8'b00000011; // 3288 :   3 - 0x3
      13'hCD9: dout  = 8'b00001111; // 3289 :  15 - 0xf
      13'hCDA: dout  = 8'b00100011; // 3290 :  35 - 0x23
      13'hCDB: dout  = 8'b01100010; // 3291 :  98 - 0x62
      13'hCDC: dout  = 8'b01100100; // 3292 : 100 - 0x64
      13'hCDD: dout  = 8'b00111100; // 3293 :  60 - 0x3c
      13'hCDE: dout  = 8'b00011100; // 3294 :  28 - 0x1c
      13'hCDF: dout  = 8'b00011110; // 3295 :  30 - 0x1e
      13'hCE0: dout  = 8'b11100000; // 3296 : 224 - 0xe0 -- Sprite 0xce
      13'hCE1: dout  = 8'b11001101; // 3297 : 205 - 0xcd
      13'hCE2: dout  = 8'b00011101; // 3298 :  29 - 0x1d
      13'hCE3: dout  = 8'b01001111; // 3299 :  79 - 0x4f
      13'hCE4: dout  = 8'b11101110; // 3300 : 238 - 0xee
      13'hCE5: dout  = 8'b11111111; // 3301 : 255 - 0xff
      13'hCE6: dout  = 8'b00111111; // 3302 :  63 - 0x3f
      13'hCE7: dout  = 8'b00111111; // 3303 :  63 - 0x3f
      13'hCE8: dout  = 8'b00011111; // 3304 :  31 - 0x1f
      13'hCE9: dout  = 8'b00111101; // 3305 :  61 - 0x3d
      13'hCEA: dout  = 8'b01101101; // 3306 : 109 - 0x6d
      13'hCEB: dout  = 8'b01001111; // 3307 :  79 - 0x4f
      13'hCEC: dout  = 8'b11101110; // 3308 : 238 - 0xee
      13'hCED: dout  = 8'b11110011; // 3309 : 243 - 0xf3
      13'hCEE: dout  = 8'b00100000; // 3310 :  32 - 0x20
      13'hCEF: dout  = 8'b00000011; // 3311 :   3 - 0x3
      13'hCF0: dout  = 8'b00111111; // 3312 :  63 - 0x3f -- Sprite 0xcf
      13'hCF1: dout  = 8'b00111111; // 3313 :  63 - 0x3f
      13'hCF2: dout  = 8'b00000000; // 3314 :   0 - 0x0
      13'hCF3: dout  = 8'b00000000; // 3315 :   0 - 0x0
      13'hCF4: dout  = 8'b01110000; // 3316 : 112 - 0x70
      13'hCF5: dout  = 8'b10111000; // 3317 : 184 - 0xb8
      13'hCF6: dout  = 8'b11111100; // 3318 : 252 - 0xfc
      13'hCF7: dout  = 8'b11111100; // 3319 : 252 - 0xfc
      13'hCF8: dout  = 8'b00000111; // 3320 :   7 - 0x7
      13'hCF9: dout  = 8'b00000111; // 3321 :   7 - 0x7
      13'hCFA: dout  = 8'b00011111; // 3322 :  31 - 0x1f
      13'hCFB: dout  = 8'b00111111; // 3323 :  63 - 0x3f
      13'hCFC: dout  = 8'b00001111; // 3324 :  15 - 0xf
      13'hCFD: dout  = 8'b01000111; // 3325 :  71 - 0x47
      13'hCFE: dout  = 8'b00000011; // 3326 :   3 - 0x3
      13'hCFF: dout  = 8'b00000000; // 3327 :   0 - 0x0
      13'hD00: dout  = 8'b00000111; // 3328 :   7 - 0x7 -- Sprite 0xd0
      13'hD01: dout  = 8'b00001111; // 3329 :  15 - 0xf
      13'hD02: dout  = 8'b00011111; // 3330 :  31 - 0x1f
      13'hD03: dout  = 8'b00111111; // 3331 :  63 - 0x3f
      13'hD04: dout  = 8'b00111110; // 3332 :  62 - 0x3e
      13'hD05: dout  = 8'b01111100; // 3333 : 124 - 0x7c
      13'hD06: dout  = 8'b01111000; // 3334 : 120 - 0x78
      13'hD07: dout  = 8'b01111000; // 3335 : 120 - 0x78
      13'hD08: dout  = 8'b00000000; // 3336 :   0 - 0x0
      13'hD09: dout  = 8'b00000000; // 3337 :   0 - 0x0
      13'hD0A: dout  = 8'b00000011; // 3338 :   3 - 0x3
      13'hD0B: dout  = 8'b00000111; // 3339 :   7 - 0x7
      13'hD0C: dout  = 8'b00001111; // 3340 :  15 - 0xf
      13'hD0D: dout  = 8'b00001111; // 3341 :  15 - 0xf
      13'hD0E: dout  = 8'b00011111; // 3342 :  31 - 0x1f
      13'hD0F: dout  = 8'b00011111; // 3343 :  31 - 0x1f
      13'hD10: dout  = 8'b00111111; // 3344 :  63 - 0x3f -- Sprite 0xd1
      13'hD11: dout  = 8'b01011100; // 3345 :  92 - 0x5c
      13'hD12: dout  = 8'b00111001; // 3346 :  57 - 0x39
      13'hD13: dout  = 8'b00111011; // 3347 :  59 - 0x3b
      13'hD14: dout  = 8'b10111111; // 3348 : 191 - 0xbf
      13'hD15: dout  = 8'b11111111; // 3349 : 255 - 0xff
      13'hD16: dout  = 8'b11111110; // 3350 : 254 - 0xfe
      13'hD17: dout  = 8'b11111110; // 3351 : 254 - 0xfe
      13'hD18: dout  = 8'b00000000; // 3352 :   0 - 0x0
      13'hD19: dout  = 8'b00100011; // 3353 :  35 - 0x23
      13'hD1A: dout  = 8'b01010111; // 3354 :  87 - 0x57
      13'hD1B: dout  = 8'b01001111; // 3355 :  79 - 0x4f
      13'hD1C: dout  = 8'b01010111; // 3356 :  87 - 0x57
      13'hD1D: dout  = 8'b00101111; // 3357 :  47 - 0x2f
      13'hD1E: dout  = 8'b11011111; // 3358 : 223 - 0xdf
      13'hD1F: dout  = 8'b00100001; // 3359 :  33 - 0x21
      13'hD20: dout  = 8'b11000000; // 3360 : 192 - 0xc0 -- Sprite 0xd2
      13'hD21: dout  = 8'b11000000; // 3361 : 192 - 0xc0
      13'hD22: dout  = 8'b10000000; // 3362 : 128 - 0x80
      13'hD23: dout  = 8'b10000000; // 3363 : 128 - 0x80
      13'hD24: dout  = 8'b10000000; // 3364 : 128 - 0x80
      13'hD25: dout  = 8'b10000000; // 3365 : 128 - 0x80
      13'hD26: dout  = 8'b00000000; // 3366 :   0 - 0x0
      13'hD27: dout  = 8'b00000000; // 3367 :   0 - 0x0
      13'hD28: dout  = 8'b00000000; // 3368 :   0 - 0x0
      13'hD29: dout  = 8'b00000000; // 3369 :   0 - 0x0
      13'hD2A: dout  = 8'b00000000; // 3370 :   0 - 0x0
      13'hD2B: dout  = 8'b00000000; // 3371 :   0 - 0x0
      13'hD2C: dout  = 8'b10000000; // 3372 : 128 - 0x80
      13'hD2D: dout  = 8'b10000000; // 3373 : 128 - 0x80
      13'hD2E: dout  = 8'b00000000; // 3374 :   0 - 0x0
      13'hD2F: dout  = 8'b00000000; // 3375 :   0 - 0x0
      13'hD30: dout  = 8'b11111110; // 3376 : 254 - 0xfe -- Sprite 0xd3
      13'hD31: dout  = 8'b11111100; // 3377 : 252 - 0xfc
      13'hD32: dout  = 8'b01100001; // 3378 :  97 - 0x61
      13'hD33: dout  = 8'b00001111; // 3379 :  15 - 0xf
      13'hD34: dout  = 8'b01111111; // 3380 : 127 - 0x7f
      13'hD35: dout  = 8'b00111111; // 3381 :  63 - 0x3f
      13'hD36: dout  = 8'b00011111; // 3382 :  31 - 0x1f
      13'hD37: dout  = 8'b00011110; // 3383 :  30 - 0x1e
      13'hD38: dout  = 8'b00100011; // 3384 :  35 - 0x23
      13'hD39: dout  = 8'b00001111; // 3385 :  15 - 0xf
      13'hD3A: dout  = 8'b00011110; // 3386 :  30 - 0x1e
      13'hD3B: dout  = 8'b11110000; // 3387 : 240 - 0xf0
      13'hD3C: dout  = 8'b00011100; // 3388 :  28 - 0x1c
      13'hD3D: dout  = 8'b00111111; // 3389 :  63 - 0x3f
      13'hD3E: dout  = 8'b00011111; // 3390 :  31 - 0x1f
      13'hD3F: dout  = 8'b00011110; // 3391 :  30 - 0x1e
      13'hD40: dout  = 8'b11110000; // 3392 : 240 - 0xf0 -- Sprite 0xd4
      13'hD41: dout  = 8'b01111000; // 3393 : 120 - 0x78
      13'hD42: dout  = 8'b11100100; // 3394 : 228 - 0xe4
      13'hD43: dout  = 8'b11001000; // 3395 : 200 - 0xc8
      13'hD44: dout  = 8'b11001100; // 3396 : 204 - 0xcc
      13'hD45: dout  = 8'b10111110; // 3397 : 190 - 0xbe
      13'hD46: dout  = 8'b10111110; // 3398 : 190 - 0xbe
      13'hD47: dout  = 8'b00111110; // 3399 :  62 - 0x3e
      13'hD48: dout  = 8'b00000000; // 3400 :   0 - 0x0
      13'hD49: dout  = 8'b10000000; // 3401 : 128 - 0x80
      13'hD4A: dout  = 8'b00011000; // 3402 :  24 - 0x18
      13'hD4B: dout  = 8'b00110000; // 3403 :  48 - 0x30
      13'hD4C: dout  = 8'b00110100; // 3404 :  52 - 0x34
      13'hD4D: dout  = 8'b11111110; // 3405 : 254 - 0xfe
      13'hD4E: dout  = 8'b11111110; // 3406 : 254 - 0xfe
      13'hD4F: dout  = 8'b11111110; // 3407 : 254 - 0xfe
      13'hD50: dout  = 8'b00000000; // 3408 :   0 - 0x0 -- Sprite 0xd5
      13'hD51: dout  = 8'b00000001; // 3409 :   1 - 0x1
      13'hD52: dout  = 8'b00000000; // 3410 :   0 - 0x0
      13'hD53: dout  = 8'b00000111; // 3411 :   7 - 0x7
      13'hD54: dout  = 8'b00000111; // 3412 :   7 - 0x7
      13'hD55: dout  = 8'b00000111; // 3413 :   7 - 0x7
      13'hD56: dout  = 8'b00000111; // 3414 :   7 - 0x7
      13'hD57: dout  = 8'b00011111; // 3415 :  31 - 0x1f
      13'hD58: dout  = 8'b00000000; // 3416 :   0 - 0x0
      13'hD59: dout  = 8'b00000000; // 3417 :   0 - 0x0
      13'hD5A: dout  = 8'b00000001; // 3418 :   1 - 0x1
      13'hD5B: dout  = 8'b00000100; // 3419 :   4 - 0x4
      13'hD5C: dout  = 8'b00000110; // 3420 :   6 - 0x6
      13'hD5D: dout  = 8'b00000110; // 3421 :   6 - 0x6
      13'hD5E: dout  = 8'b00000111; // 3422 :   7 - 0x7
      13'hD5F: dout  = 8'b00000111; // 3423 :   7 - 0x7
      13'hD60: dout  = 8'b00000000; // 3424 :   0 - 0x0 -- Sprite 0xd6
      13'hD61: dout  = 8'b00000000; // 3425 :   0 - 0x0
      13'hD62: dout  = 8'b00001111; // 3426 :  15 - 0xf
      13'hD63: dout  = 8'b00111111; // 3427 :  63 - 0x3f
      13'hD64: dout  = 8'b00111111; // 3428 :  63 - 0x3f
      13'hD65: dout  = 8'b00001111; // 3429 :  15 - 0xf
      13'hD66: dout  = 8'b00000000; // 3430 :   0 - 0x0
      13'hD67: dout  = 8'b00000000; // 3431 :   0 - 0x0
      13'hD68: dout  = 8'b00001111; // 3432 :  15 - 0xf
      13'hD69: dout  = 8'b00111111; // 3433 :  63 - 0x3f
      13'hD6A: dout  = 8'b01111111; // 3434 : 127 - 0x7f
      13'hD6B: dout  = 8'b11111000; // 3435 : 248 - 0xf8
      13'hD6C: dout  = 8'b11111000; // 3436 : 248 - 0xf8
      13'hD6D: dout  = 8'b01111111; // 3437 : 127 - 0x7f
      13'hD6E: dout  = 8'b00111111; // 3438 :  63 - 0x3f
      13'hD6F: dout  = 8'b00001111; // 3439 :  15 - 0xf
      13'hD70: dout  = 8'b01111000; // 3440 : 120 - 0x78 -- Sprite 0xd7
      13'hD71: dout  = 8'b01111100; // 3441 : 124 - 0x7c
      13'hD72: dout  = 8'b01111110; // 3442 : 126 - 0x7e
      13'hD73: dout  = 8'b01111111; // 3443 : 127 - 0x7f
      13'hD74: dout  = 8'b00111111; // 3444 :  63 - 0x3f
      13'hD75: dout  = 8'b00111111; // 3445 :  63 - 0x3f
      13'hD76: dout  = 8'b00011011; // 3446 :  27 - 0x1b
      13'hD77: dout  = 8'b00001001; // 3447 :   9 - 0x9
      13'hD78: dout  = 8'b00011111; // 3448 :  31 - 0x1f
      13'hD79: dout  = 8'b00011111; // 3449 :  31 - 0x1f
      13'hD7A: dout  = 8'b00011111; // 3450 :  31 - 0x1f
      13'hD7B: dout  = 8'b00001011; // 3451 :  11 - 0xb
      13'hD7C: dout  = 8'b00000001; // 3452 :   1 - 0x1
      13'hD7D: dout  = 8'b00000001; // 3453 :   1 - 0x1
      13'hD7E: dout  = 8'b00000000; // 3454 :   0 - 0x0
      13'hD7F: dout  = 8'b00000000; // 3455 :   0 - 0x0
      13'hD80: dout  = 8'b00001100; // 3456 :  12 - 0xc -- Sprite 0xd8
      13'hD81: dout  = 8'b00000000; // 3457 :   0 - 0x0
      13'hD82: dout  = 8'b00000000; // 3458 :   0 - 0x0
      13'hD83: dout  = 8'b00000000; // 3459 :   0 - 0x0
      13'hD84: dout  = 8'b00000111; // 3460 :   7 - 0x7
      13'hD85: dout  = 8'b01111111; // 3461 : 127 - 0x7f
      13'hD86: dout  = 8'b01111100; // 3462 : 124 - 0x7c
      13'hD87: dout  = 8'b00000000; // 3463 :   0 - 0x0
      13'hD88: dout  = 8'b00000011; // 3464 :   3 - 0x3
      13'hD89: dout  = 8'b00011111; // 3465 :  31 - 0x1f
      13'hD8A: dout  = 8'b00111111; // 3466 :  63 - 0x3f
      13'hD8B: dout  = 8'b00111111; // 3467 :  63 - 0x3f
      13'hD8C: dout  = 8'b01111000; // 3468 : 120 - 0x78
      13'hD8D: dout  = 8'b00000000; // 3469 :   0 - 0x0
      13'hD8E: dout  = 8'b00000011; // 3470 :   3 - 0x3
      13'hD8F: dout  = 8'b11111111; // 3471 : 255 - 0xff
      13'hD90: dout  = 8'b00000001; // 3472 :   1 - 0x1 -- Sprite 0xd9
      13'hD91: dout  = 8'b11100001; // 3473 : 225 - 0xe1
      13'hD92: dout  = 8'b01110001; // 3474 : 113 - 0x71
      13'hD93: dout  = 8'b01111001; // 3475 : 121 - 0x79
      13'hD94: dout  = 8'b00111101; // 3476 :  61 - 0x3d
      13'hD95: dout  = 8'b00111101; // 3477 :  61 - 0x3d
      13'hD96: dout  = 8'b00011111; // 3478 :  31 - 0x1f
      13'hD97: dout  = 8'b00000011; // 3479 :   3 - 0x3
      13'hD98: dout  = 8'b00000000; // 3480 :   0 - 0x0
      13'hD99: dout  = 8'b00000000; // 3481 :   0 - 0x0
      13'hD9A: dout  = 8'b00000000; // 3482 :   0 - 0x0
      13'hD9B: dout  = 8'b00000000; // 3483 :   0 - 0x0
      13'hD9C: dout  = 8'b00000000; // 3484 :   0 - 0x0
      13'hD9D: dout  = 8'b00000000; // 3485 :   0 - 0x0
      13'hD9E: dout  = 8'b00000000; // 3486 :   0 - 0x0
      13'hD9F: dout  = 8'b00000000; // 3487 :   0 - 0x0
      13'hDA0: dout  = 8'b00111111; // 3488 :  63 - 0x3f -- Sprite 0xda
      13'hDA1: dout  = 8'b00111111; // 3489 :  63 - 0x3f
      13'hDA2: dout  = 8'b00011111; // 3490 :  31 - 0x1f
      13'hDA3: dout  = 8'b00011011; // 3491 :  27 - 0x1b
      13'hDA4: dout  = 8'b00110110; // 3492 :  54 - 0x36
      13'hDA5: dout  = 8'b00110000; // 3493 :  48 - 0x30
      13'hDA6: dout  = 8'b01111111; // 3494 : 127 - 0x7f
      13'hDA7: dout  = 8'b00111111; // 3495 :  63 - 0x3f
      13'hDA8: dout  = 8'b00100011; // 3496 :  35 - 0x23
      13'hDA9: dout  = 8'b00100111; // 3497 :  39 - 0x27
      13'hDAA: dout  = 8'b00011111; // 3498 :  31 - 0x1f
      13'hDAB: dout  = 8'b00000111; // 3499 :   7 - 0x7
      13'hDAC: dout  = 8'b00001111; // 3500 :  15 - 0xf
      13'hDAD: dout  = 8'b00011111; // 3501 :  31 - 0x1f
      13'hDAE: dout  = 8'b01111111; // 3502 : 127 - 0x7f
      13'hDAF: dout  = 8'b00111111; // 3503 :  63 - 0x3f
      13'hDB0: dout  = 8'b11111000; // 3504 : 248 - 0xf8 -- Sprite 0xdb
      13'hDB1: dout  = 8'b11111000; // 3505 : 248 - 0xf8
      13'hDB2: dout  = 8'b11111000; // 3506 : 248 - 0xf8
      13'hDB3: dout  = 8'b10111000; // 3507 : 184 - 0xb8
      13'hDB4: dout  = 8'b00011000; // 3508 :  24 - 0x18
      13'hDB5: dout  = 8'b11011000; // 3509 : 216 - 0xd8
      13'hDB6: dout  = 8'b11011000; // 3510 : 216 - 0xd8
      13'hDB7: dout  = 8'b10111000; // 3511 : 184 - 0xb8
      13'hDB8: dout  = 8'b11100000; // 3512 : 224 - 0xe0
      13'hDB9: dout  = 8'b10000000; // 3513 : 128 - 0x80
      13'hDBA: dout  = 8'b10000000; // 3514 : 128 - 0x80
      13'hDBB: dout  = 8'b01000000; // 3515 :  64 - 0x40
      13'hDBC: dout  = 8'b11100000; // 3516 : 224 - 0xe0
      13'hDBD: dout  = 8'b11100000; // 3517 : 224 - 0xe0
      13'hDBE: dout  = 8'b11100000; // 3518 : 224 - 0xe0
      13'hDBF: dout  = 8'b11000000; // 3519 : 192 - 0xc0
      13'hDC0: dout  = 8'b00000001; // 3520 :   1 - 0x1 -- Sprite 0xdc
      13'hDC1: dout  = 8'b00000010; // 3521 :   2 - 0x2
      13'hDC2: dout  = 8'b00000100; // 3522 :   4 - 0x4
      13'hDC3: dout  = 8'b00000100; // 3523 :   4 - 0x4
      13'hDC4: dout  = 8'b00001000; // 3524 :   8 - 0x8
      13'hDC5: dout  = 8'b00001000; // 3525 :   8 - 0x8
      13'hDC6: dout  = 8'b00010000; // 3526 :  16 - 0x10
      13'hDC7: dout  = 8'b00010000; // 3527 :  16 - 0x10
      13'hDC8: dout  = 8'b00000011; // 3528 :   3 - 0x3
      13'hDC9: dout  = 8'b00000111; // 3529 :   7 - 0x7
      13'hDCA: dout  = 8'b00001111; // 3530 :  15 - 0xf
      13'hDCB: dout  = 8'b00011111; // 3531 :  31 - 0x1f
      13'hDCC: dout  = 8'b00111111; // 3532 :  63 - 0x3f
      13'hDCD: dout  = 8'b01111111; // 3533 : 127 - 0x7f
      13'hDCE: dout  = 8'b11111111; // 3534 : 255 - 0xff
      13'hDCF: dout  = 8'b00011111; // 3535 :  31 - 0x1f
      13'hDD0: dout  = 8'b00000000; // 3536 :   0 - 0x0 -- Sprite 0xdd
      13'hDD1: dout  = 8'b00001111; // 3537 :  15 - 0xf
      13'hDD2: dout  = 8'b00010011; // 3538 :  19 - 0x13
      13'hDD3: dout  = 8'b00001101; // 3539 :  13 - 0xd
      13'hDD4: dout  = 8'b00001101; // 3540 :  13 - 0xd
      13'hDD5: dout  = 8'b00010011; // 3541 :  19 - 0x13
      13'hDD6: dout  = 8'b00001100; // 3542 :  12 - 0xc
      13'hDD7: dout  = 8'b00100000; // 3543 :  32 - 0x20
      13'hDD8: dout  = 8'b00011111; // 3544 :  31 - 0x1f
      13'hDD9: dout  = 8'b00010000; // 3545 :  16 - 0x10
      13'hDDA: dout  = 8'b00001100; // 3546 :  12 - 0xc
      13'hDDB: dout  = 8'b00010010; // 3547 :  18 - 0x12
      13'hDDC: dout  = 8'b00010010; // 3548 :  18 - 0x12
      13'hDDD: dout  = 8'b00101100; // 3549 :  44 - 0x2c
      13'hDDE: dout  = 8'b00111111; // 3550 :  63 - 0x3f
      13'hDDF: dout  = 8'b00111111; // 3551 :  63 - 0x3f
      13'hDE0: dout  = 8'b00000000; // 3552 :   0 - 0x0 -- Sprite 0xde
      13'hDE1: dout  = 8'b00100100; // 3553 :  36 - 0x24
      13'hDE2: dout  = 8'b00000000; // 3554 :   0 - 0x0
      13'hDE3: dout  = 8'b00100100; // 3555 :  36 - 0x24
      13'hDE4: dout  = 8'b00000000; // 3556 :   0 - 0x0
      13'hDE5: dout  = 8'b00000100; // 3557 :   4 - 0x4
      13'hDE6: dout  = 8'b00000000; // 3558 :   0 - 0x0
      13'hDE7: dout  = 8'b00000000; // 3559 :   0 - 0x0
      13'hDE8: dout  = 8'b00110111; // 3560 :  55 - 0x37
      13'hDE9: dout  = 8'b00110110; // 3561 :  54 - 0x36
      13'hDEA: dout  = 8'b00110110; // 3562 :  54 - 0x36
      13'hDEB: dout  = 8'b00110110; // 3563 :  54 - 0x36
      13'hDEC: dout  = 8'b00010110; // 3564 :  22 - 0x16
      13'hDED: dout  = 8'b00010110; // 3565 :  22 - 0x16
      13'hDEE: dout  = 8'b00010010; // 3566 :  18 - 0x12
      13'hDEF: dout  = 8'b00000010; // 3567 :   2 - 0x2
      13'hDF0: dout  = 8'b00001111; // 3568 :  15 - 0xf -- Sprite 0xdf
      13'hDF1: dout  = 8'b01000001; // 3569 :  65 - 0x41
      13'hDF2: dout  = 8'b00000000; // 3570 :   0 - 0x0
      13'hDF3: dout  = 8'b10001000; // 3571 : 136 - 0x88
      13'hDF4: dout  = 8'b00000000; // 3572 :   0 - 0x0
      13'hDF5: dout  = 8'b01000100; // 3573 :  68 - 0x44
      13'hDF6: dout  = 8'b00000000; // 3574 :   0 - 0x0
      13'hDF7: dout  = 8'b00000000; // 3575 :   0 - 0x0
      13'hDF8: dout  = 8'b00010000; // 3576 :  16 - 0x10
      13'hDF9: dout  = 8'b01111110; // 3577 : 126 - 0x7e
      13'hDFA: dout  = 8'b11111111; // 3578 : 255 - 0xff
      13'hDFB: dout  = 8'b11111111; // 3579 : 255 - 0xff
      13'hDFC: dout  = 8'b11110110; // 3580 : 246 - 0xf6
      13'hDFD: dout  = 8'b01110110; // 3581 : 118 - 0x76
      13'hDFE: dout  = 8'b00111010; // 3582 :  58 - 0x3a
      13'hDFF: dout  = 8'b00011010; // 3583 :  26 - 0x1a
      13'hE00: dout  = 8'b00111000; // 3584 :  56 - 0x38 -- Sprite 0xe0
      13'hE01: dout  = 8'b01111100; // 3585 : 124 - 0x7c
      13'hE02: dout  = 8'b11111110; // 3586 : 254 - 0xfe
      13'hE03: dout  = 8'b11111110; // 3587 : 254 - 0xfe
      13'hE04: dout  = 8'b00111011; // 3588 :  59 - 0x3b
      13'hE05: dout  = 8'b00000011; // 3589 :   3 - 0x3
      13'hE06: dout  = 8'b00000011; // 3590 :   3 - 0x3
      13'hE07: dout  = 8'b00000011; // 3591 :   3 - 0x3
      13'hE08: dout  = 8'b00000000; // 3592 :   0 - 0x0
      13'hE09: dout  = 8'b00000000; // 3593 :   0 - 0x0
      13'hE0A: dout  = 8'b00111000; // 3594 :  56 - 0x38
      13'hE0B: dout  = 8'b00000100; // 3595 :   4 - 0x4
      13'hE0C: dout  = 8'b00000000; // 3596 :   0 - 0x0
      13'hE0D: dout  = 8'b00000000; // 3597 :   0 - 0x0
      13'hE0E: dout  = 8'b00000000; // 3598 :   0 - 0x0
      13'hE0F: dout  = 8'b00000000; // 3599 :   0 - 0x0
      13'hE10: dout  = 8'b00000011; // 3600 :   3 - 0x3 -- Sprite 0xe1
      13'hE11: dout  = 8'b00110011; // 3601 :  51 - 0x33
      13'hE12: dout  = 8'b01111011; // 3602 : 123 - 0x7b
      13'hE13: dout  = 8'b01111111; // 3603 : 127 - 0x7f
      13'hE14: dout  = 8'b11111111; // 3604 : 255 - 0xff
      13'hE15: dout  = 8'b11111011; // 3605 : 251 - 0xfb
      13'hE16: dout  = 8'b00000011; // 3606 :   3 - 0x3
      13'hE17: dout  = 8'b00000011; // 3607 :   3 - 0x3
      13'hE18: dout  = 8'b00000000; // 3608 :   0 - 0x0
      13'hE19: dout  = 8'b00000000; // 3609 :   0 - 0x0
      13'hE1A: dout  = 8'b00000000; // 3610 :   0 - 0x0
      13'hE1B: dout  = 8'b00111000; // 3611 :  56 - 0x38
      13'hE1C: dout  = 8'b01000000; // 3612 :  64 - 0x40
      13'hE1D: dout  = 8'b00000000; // 3613 :   0 - 0x0
      13'hE1E: dout  = 8'b00000000; // 3614 :   0 - 0x0
      13'hE1F: dout  = 8'b00000000; // 3615 :   0 - 0x0
      13'hE20: dout  = 8'b11011100; // 3616 : 220 - 0xdc -- Sprite 0xe2
      13'hE21: dout  = 8'b11000000; // 3617 : 192 - 0xc0
      13'hE22: dout  = 8'b11100000; // 3618 : 224 - 0xe0
      13'hE23: dout  = 8'b11100000; // 3619 : 224 - 0xe0
      13'hE24: dout  = 8'b11100000; // 3620 : 224 - 0xe0
      13'hE25: dout  = 8'b11100000; // 3621 : 224 - 0xe0
      13'hE26: dout  = 8'b11100000; // 3622 : 224 - 0xe0
      13'hE27: dout  = 8'b11000000; // 3623 : 192 - 0xc0
      13'hE28: dout  = 8'b11111100; // 3624 : 252 - 0xfc
      13'hE29: dout  = 8'b10100000; // 3625 : 160 - 0xa0
      13'hE2A: dout  = 8'b10000000; // 3626 : 128 - 0x80
      13'hE2B: dout  = 8'b10000000; // 3627 : 128 - 0x80
      13'hE2C: dout  = 8'b00000000; // 3628 :   0 - 0x0
      13'hE2D: dout  = 8'b00000000; // 3629 :   0 - 0x0
      13'hE2E: dout  = 8'b00000000; // 3630 :   0 - 0x0
      13'hE2F: dout  = 8'b00000000; // 3631 :   0 - 0x0
      13'hE30: dout  = 8'b00111111; // 3632 :  63 - 0x3f -- Sprite 0xe3
      13'hE31: dout  = 8'b01011111; // 3633 :  95 - 0x5f
      13'hE32: dout  = 8'b00111111; // 3634 :  63 - 0x3f
      13'hE33: dout  = 8'b00111111; // 3635 :  63 - 0x3f
      13'hE34: dout  = 8'b10111011; // 3636 : 187 - 0xbb
      13'hE35: dout  = 8'b11111000; // 3637 : 248 - 0xf8
      13'hE36: dout  = 8'b11111110; // 3638 : 254 - 0xfe
      13'hE37: dout  = 8'b11111110; // 3639 : 254 - 0xfe
      13'hE38: dout  = 8'b00000111; // 3640 :   7 - 0x7
      13'hE39: dout  = 8'b00100111; // 3641 :  39 - 0x27
      13'hE3A: dout  = 8'b01010111; // 3642 :  87 - 0x57
      13'hE3B: dout  = 8'b01001111; // 3643 :  79 - 0x4f
      13'hE3C: dout  = 8'b01010111; // 3644 :  87 - 0x57
      13'hE3D: dout  = 8'b00100111; // 3645 :  39 - 0x27
      13'hE3E: dout  = 8'b11000001; // 3646 : 193 - 0xc1
      13'hE3F: dout  = 8'b00100001; // 3647 :  33 - 0x21
      13'hE40: dout  = 8'b00011111; // 3648 :  31 - 0x1f -- Sprite 0xe4
      13'hE41: dout  = 8'b00001111; // 3649 :  15 - 0xf
      13'hE42: dout  = 8'b00001111; // 3650 :  15 - 0xf
      13'hE43: dout  = 8'b00011111; // 3651 :  31 - 0x1f
      13'hE44: dout  = 8'b00011111; // 3652 :  31 - 0x1f
      13'hE45: dout  = 8'b00011110; // 3653 :  30 - 0x1e
      13'hE46: dout  = 8'b00111000; // 3654 :  56 - 0x38
      13'hE47: dout  = 8'b00110000; // 3655 :  48 - 0x30
      13'hE48: dout  = 8'b00011101; // 3656 :  29 - 0x1d
      13'hE49: dout  = 8'b00001111; // 3657 :  15 - 0xf
      13'hE4A: dout  = 8'b00001111; // 3658 :  15 - 0xf
      13'hE4B: dout  = 8'b00011111; // 3659 :  31 - 0x1f
      13'hE4C: dout  = 8'b00011111; // 3660 :  31 - 0x1f
      13'hE4D: dout  = 8'b00011110; // 3661 :  30 - 0x1e
      13'hE4E: dout  = 8'b00111000; // 3662 :  56 - 0x38
      13'hE4F: dout  = 8'b00110000; // 3663 :  48 - 0x30
      13'hE50: dout  = 8'b00000000; // 3664 :   0 - 0x0 -- Sprite 0xe5
      13'hE51: dout  = 8'b00100000; // 3665 :  32 - 0x20
      13'hE52: dout  = 8'b01100000; // 3666 :  96 - 0x60
      13'hE53: dout  = 8'b01100000; // 3667 :  96 - 0x60
      13'hE54: dout  = 8'b01110000; // 3668 : 112 - 0x70
      13'hE55: dout  = 8'b11110000; // 3669 : 240 - 0xf0
      13'hE56: dout  = 8'b11111000; // 3670 : 248 - 0xf8
      13'hE57: dout  = 8'b11111000; // 3671 : 248 - 0xf8
      13'hE58: dout  = 8'b00000000; // 3672 :   0 - 0x0
      13'hE59: dout  = 8'b00000000; // 3673 :   0 - 0x0
      13'hE5A: dout  = 8'b00111000; // 3674 :  56 - 0x38
      13'hE5B: dout  = 8'b00010000; // 3675 :  16 - 0x10
      13'hE5C: dout  = 8'b01001100; // 3676 :  76 - 0x4c
      13'hE5D: dout  = 8'b00011000; // 3677 :  24 - 0x18
      13'hE5E: dout  = 8'b10000110; // 3678 : 134 - 0x86
      13'hE5F: dout  = 8'b00100100; // 3679 :  36 - 0x24
      13'hE60: dout  = 8'b11111000; // 3680 : 248 - 0xf8 -- Sprite 0xe6
      13'hE61: dout  = 8'b11111100; // 3681 : 252 - 0xfc
      13'hE62: dout  = 8'b11111100; // 3682 : 252 - 0xfc
      13'hE63: dout  = 8'b01111110; // 3683 : 126 - 0x7e
      13'hE64: dout  = 8'b01111110; // 3684 : 126 - 0x7e
      13'hE65: dout  = 8'b00111110; // 3685 :  62 - 0x3e
      13'hE66: dout  = 8'b00011111; // 3686 :  31 - 0x1f
      13'hE67: dout  = 8'b00000111; // 3687 :   7 - 0x7
      13'hE68: dout  = 8'b00000000; // 3688 :   0 - 0x0
      13'hE69: dout  = 8'b01000010; // 3689 :  66 - 0x42
      13'hE6A: dout  = 8'b00001010; // 3690 :  10 - 0xa
      13'hE6B: dout  = 8'b01000000; // 3691 :  64 - 0x40
      13'hE6C: dout  = 8'b00010000; // 3692 :  16 - 0x10
      13'hE6D: dout  = 8'b00000010; // 3693 :   2 - 0x2
      13'hE6E: dout  = 8'b00001000; // 3694 :   8 - 0x8
      13'hE6F: dout  = 8'b00000010; // 3695 :   2 - 0x2
      13'hE70: dout  = 8'b00000000; // 3696 :   0 - 0x0 -- Sprite 0xe7
      13'hE71: dout  = 8'b11000000; // 3697 : 192 - 0xc0
      13'hE72: dout  = 8'b01110000; // 3698 : 112 - 0x70
      13'hE73: dout  = 8'b10111000; // 3699 : 184 - 0xb8
      13'hE74: dout  = 8'b11110100; // 3700 : 244 - 0xf4
      13'hE75: dout  = 8'b11110010; // 3701 : 242 - 0xf2
      13'hE76: dout  = 8'b11110101; // 3702 : 245 - 0xf5
      13'hE77: dout  = 8'b01111011; // 3703 : 123 - 0x7b
      13'hE78: dout  = 8'b00000000; // 3704 :   0 - 0x0
      13'hE79: dout  = 8'b00000000; // 3705 :   0 - 0x0
      13'hE7A: dout  = 8'b10000000; // 3706 : 128 - 0x80
      13'hE7B: dout  = 8'b01000000; // 3707 :  64 - 0x40
      13'hE7C: dout  = 8'b00001000; // 3708 :   8 - 0x8
      13'hE7D: dout  = 8'b00001100; // 3709 :  12 - 0xc
      13'hE7E: dout  = 8'b00001010; // 3710 :  10 - 0xa
      13'hE7F: dout  = 8'b10000100; // 3711 : 132 - 0x84
      13'hE80: dout  = 8'b00000000; // 3712 :   0 - 0x0 -- Sprite 0xe8
      13'hE81: dout  = 8'b11011111; // 3713 : 223 - 0xdf
      13'hE82: dout  = 8'b00010000; // 3714 :  16 - 0x10
      13'hE83: dout  = 8'b11111111; // 3715 : 255 - 0xff
      13'hE84: dout  = 8'b11011111; // 3716 : 223 - 0xdf
      13'hE85: dout  = 8'b11111111; // 3717 : 255 - 0xff
      13'hE86: dout  = 8'b11111111; // 3718 : 255 - 0xff
      13'hE87: dout  = 8'b11111001; // 3719 : 249 - 0xf9
      13'hE88: dout  = 8'b00000000; // 3720 :   0 - 0x0
      13'hE89: dout  = 8'b00000000; // 3721 :   0 - 0x0
      13'hE8A: dout  = 8'b11001111; // 3722 : 207 - 0xcf
      13'hE8B: dout  = 8'b00100000; // 3723 :  32 - 0x20
      13'hE8C: dout  = 8'b00100000; // 3724 :  32 - 0x20
      13'hE8D: dout  = 8'b00100000; // 3725 :  32 - 0x20
      13'hE8E: dout  = 8'b00100110; // 3726 :  38 - 0x26
      13'hE8F: dout  = 8'b00101110; // 3727 :  46 - 0x2e
      13'hE90: dout  = 8'b00011111; // 3728 :  31 - 0x1f -- Sprite 0xe9
      13'hE91: dout  = 8'b00011111; // 3729 :  31 - 0x1f
      13'hE92: dout  = 8'b00111110; // 3730 :  62 - 0x3e
      13'hE93: dout  = 8'b11111100; // 3731 : 252 - 0xfc
      13'hE94: dout  = 8'b11111000; // 3732 : 248 - 0xf8
      13'hE95: dout  = 8'b11110000; // 3733 : 240 - 0xf0
      13'hE96: dout  = 8'b11000000; // 3734 : 192 - 0xc0
      13'hE97: dout  = 8'b00000000; // 3735 :   0 - 0x0
      13'hE98: dout  = 8'b11100000; // 3736 : 224 - 0xe0
      13'hE99: dout  = 8'b11100000; // 3737 : 224 - 0xe0
      13'hE9A: dout  = 8'b11000000; // 3738 : 192 - 0xc0
      13'hE9B: dout  = 8'b00000000; // 3739 :   0 - 0x0
      13'hE9C: dout  = 8'b00000000; // 3740 :   0 - 0x0
      13'hE9D: dout  = 8'b00000000; // 3741 :   0 - 0x0
      13'hE9E: dout  = 8'b00000000; // 3742 :   0 - 0x0
      13'hE9F: dout  = 8'b00000000; // 3743 :   0 - 0x0
      13'hEA0: dout  = 8'b11111000; // 3744 : 248 - 0xf8 -- Sprite 0xea
      13'hEA1: dout  = 8'b11111100; // 3745 : 252 - 0xfc
      13'hEA2: dout  = 8'b11111110; // 3746 : 254 - 0xfe
      13'hEA3: dout  = 8'b11111111; // 3747 : 255 - 0xff
      13'hEA4: dout  = 8'b11111111; // 3748 : 255 - 0xff
      13'hEA5: dout  = 8'b11011111; // 3749 : 223 - 0xdf
      13'hEA6: dout  = 8'b11011111; // 3750 : 223 - 0xdf
      13'hEA7: dout  = 8'b00000000; // 3751 :   0 - 0x0
      13'hEA8: dout  = 8'b00101111; // 3752 :  47 - 0x2f
      13'hEA9: dout  = 8'b00100011; // 3753 :  35 - 0x23
      13'hEAA: dout  = 8'b00100001; // 3754 :  33 - 0x21
      13'hEAB: dout  = 8'b00100000; // 3755 :  32 - 0x20
      13'hEAC: dout  = 8'b00100000; // 3756 :  32 - 0x20
      13'hEAD: dout  = 8'b00000000; // 3757 :   0 - 0x0
      13'hEAE: dout  = 8'b00000000; // 3758 :   0 - 0x0
      13'hEAF: dout  = 8'b00000000; // 3759 :   0 - 0x0
      13'hEB0: dout  = 8'b11000001; // 3760 : 193 - 0xc1 -- Sprite 0xeb
      13'hEB1: dout  = 8'b11110001; // 3761 : 241 - 0xf1
      13'hEB2: dout  = 8'b01111001; // 3762 : 121 - 0x79
      13'hEB3: dout  = 8'b01111101; // 3763 : 125 - 0x7d
      13'hEB4: dout  = 8'b00111101; // 3764 :  61 - 0x3d
      13'hEB5: dout  = 8'b00111111; // 3765 :  63 - 0x3f
      13'hEB6: dout  = 8'b00011111; // 3766 :  31 - 0x1f
      13'hEB7: dout  = 8'b00000011; // 3767 :   3 - 0x3
      13'hEB8: dout  = 8'b11000001; // 3768 : 193 - 0xc1
      13'hEB9: dout  = 8'b10110001; // 3769 : 177 - 0xb1
      13'hEBA: dout  = 8'b01011001; // 3770 :  89 - 0x59
      13'hEBB: dout  = 8'b01101101; // 3771 : 109 - 0x6d
      13'hEBC: dout  = 8'b00110101; // 3772 :  53 - 0x35
      13'hEBD: dout  = 8'b00111011; // 3773 :  59 - 0x3b
      13'hEBE: dout  = 8'b00011111; // 3774 :  31 - 0x1f
      13'hEBF: dout  = 8'b00000011; // 3775 :   3 - 0x3
      13'hEC0: dout  = 8'b00000010; // 3776 :   2 - 0x2 -- Sprite 0xec
      13'hEC1: dout  = 8'b00000110; // 3777 :   6 - 0x6
      13'hEC2: dout  = 8'b00001110; // 3778 :  14 - 0xe
      13'hEC3: dout  = 8'b00001110; // 3779 :  14 - 0xe
      13'hEC4: dout  = 8'b00011110; // 3780 :  30 - 0x1e
      13'hEC5: dout  = 8'b00011110; // 3781 :  30 - 0x1e
      13'hEC6: dout  = 8'b00111110; // 3782 :  62 - 0x3e
      13'hEC7: dout  = 8'b00111110; // 3783 :  62 - 0x3e
      13'hEC8: dout  = 8'b00000000; // 3784 :   0 - 0x0
      13'hEC9: dout  = 8'b00000010; // 3785 :   2 - 0x2
      13'hECA: dout  = 8'b00000000; // 3786 :   0 - 0x0
      13'hECB: dout  = 8'b00001000; // 3787 :   8 - 0x8
      13'hECC: dout  = 8'b00000010; // 3788 :   2 - 0x2
      13'hECD: dout  = 8'b00000000; // 3789 :   0 - 0x0
      13'hECE: dout  = 8'b00101000; // 3790 :  40 - 0x28
      13'hECF: dout  = 8'b00000000; // 3791 :   0 - 0x0
      13'hED0: dout  = 8'b00111110; // 3792 :  62 - 0x3e -- Sprite 0xed
      13'hED1: dout  = 8'b00111110; // 3793 :  62 - 0x3e
      13'hED2: dout  = 8'b00111110; // 3794 :  62 - 0x3e
      13'hED3: dout  = 8'b00111110; // 3795 :  62 - 0x3e
      13'hED4: dout  = 8'b00011110; // 3796 :  30 - 0x1e
      13'hED5: dout  = 8'b00011110; // 3797 :  30 - 0x1e
      13'hED6: dout  = 8'b00001110; // 3798 :  14 - 0xe
      13'hED7: dout  = 8'b00000010; // 3799 :   2 - 0x2
      13'hED8: dout  = 8'b00000100; // 3800 :   4 - 0x4
      13'hED9: dout  = 8'b00010000; // 3801 :  16 - 0x10
      13'hEDA: dout  = 8'b00000010; // 3802 :   2 - 0x2
      13'hEDB: dout  = 8'b00010000; // 3803 :  16 - 0x10
      13'hEDC: dout  = 8'b00000100; // 3804 :   4 - 0x4
      13'hEDD: dout  = 8'b00000000; // 3805 :   0 - 0x0
      13'hEDE: dout  = 8'b00001010; // 3806 :  10 - 0xa
      13'hEDF: dout  = 8'b00000000; // 3807 :   0 - 0x0
      13'hEE0: dout  = 8'b11000001; // 3808 : 193 - 0xc1 -- Sprite 0xee
      13'hEE1: dout  = 8'b11110001; // 3809 : 241 - 0xf1
      13'hEE2: dout  = 8'b01111001; // 3810 : 121 - 0x79
      13'hEE3: dout  = 8'b01111101; // 3811 : 125 - 0x7d
      13'hEE4: dout  = 8'b00111101; // 3812 :  61 - 0x3d
      13'hEE5: dout  = 8'b00111111; // 3813 :  63 - 0x3f
      13'hEE6: dout  = 8'b00011111; // 3814 :  31 - 0x1f
      13'hEE7: dout  = 8'b00000011; // 3815 :   3 - 0x3
      13'hEE8: dout  = 8'b11000001; // 3816 : 193 - 0xc1
      13'hEE9: dout  = 8'b10110001; // 3817 : 177 - 0xb1
      13'hEEA: dout  = 8'b01011001; // 3818 :  89 - 0x59
      13'hEEB: dout  = 8'b01101101; // 3819 : 109 - 0x6d
      13'hEEC: dout  = 8'b00110101; // 3820 :  53 - 0x35
      13'hEED: dout  = 8'b00111011; // 3821 :  59 - 0x3b
      13'hEEE: dout  = 8'b00011111; // 3822 :  31 - 0x1f
      13'hEEF: dout  = 8'b00000011; // 3823 :   3 - 0x3
      13'hEF0: dout  = 8'b01111100; // 3824 : 124 - 0x7c -- Sprite 0xef
      13'hEF1: dout  = 8'b00000000; // 3825 :   0 - 0x0
      13'hEF2: dout  = 8'b00000000; // 3826 :   0 - 0x0
      13'hEF3: dout  = 8'b11111111; // 3827 : 255 - 0xff
      13'hEF4: dout  = 8'b11000011; // 3828 : 195 - 0xc3
      13'hEF5: dout  = 8'b01111111; // 3829 : 127 - 0x7f
      13'hEF6: dout  = 8'b00011111; // 3830 :  31 - 0x1f
      13'hEF7: dout  = 8'b00000011; // 3831 :   3 - 0x3
      13'hEF8: dout  = 8'b00000000; // 3832 :   0 - 0x0
      13'hEF9: dout  = 8'b00001111; // 3833 :  15 - 0xf
      13'hEFA: dout  = 8'b00011111; // 3834 :  31 - 0x1f
      13'hEFB: dout  = 8'b11111111; // 3835 : 255 - 0xff
      13'hEFC: dout  = 8'b11111100; // 3836 : 252 - 0xfc
      13'hEFD: dout  = 8'b01100011; // 3837 :  99 - 0x63
      13'hEFE: dout  = 8'b00011111; // 3838 :  31 - 0x1f
      13'hEFF: dout  = 8'b00000011; // 3839 :   3 - 0x3
      13'hF00: dout  = 8'b11111111; // 3840 : 255 - 0xff -- Sprite 0xf0
      13'hF01: dout  = 8'b11111111; // 3841 : 255 - 0xff
      13'hF02: dout  = 8'b01111100; // 3842 : 124 - 0x7c
      13'hF03: dout  = 8'b00000000; // 3843 :   0 - 0x0
      13'hF04: dout  = 8'b00000000; // 3844 :   0 - 0x0
      13'hF05: dout  = 8'b01111100; // 3845 : 124 - 0x7c
      13'hF06: dout  = 8'b11111111; // 3846 : 255 - 0xff
      13'hF07: dout  = 8'b11111111; // 3847 : 255 - 0xff
      13'hF08: dout  = 8'b00000000; // 3848 :   0 - 0x0
      13'hF09: dout  = 8'b00000000; // 3849 :   0 - 0x0
      13'hF0A: dout  = 8'b11111110; // 3850 : 254 - 0xfe
      13'hF0B: dout  = 8'b11000110; // 3851 : 198 - 0xc6
      13'hF0C: dout  = 8'b11000110; // 3852 : 198 - 0xc6
      13'hF0D: dout  = 8'b11111110; // 3853 : 254 - 0xfe
      13'hF0E: dout  = 8'b00000000; // 3854 :   0 - 0x0
      13'hF0F: dout  = 8'b00000000; // 3855 :   0 - 0x0
      13'hF10: dout  = 8'b11111111; // 3856 : 255 - 0xff -- Sprite 0xf1
      13'hF11: dout  = 8'b11111111; // 3857 : 255 - 0xff
      13'hF12: dout  = 8'b00000000; // 3858 :   0 - 0x0
      13'hF13: dout  = 8'b00000100; // 3859 :   4 - 0x4
      13'hF14: dout  = 8'b00001100; // 3860 :  12 - 0xc
      13'hF15: dout  = 8'b00011000; // 3861 :  24 - 0x18
      13'hF16: dout  = 8'b00110000; // 3862 :  48 - 0x30
      13'hF17: dout  = 8'b00000000; // 3863 :   0 - 0x0
      13'hF18: dout  = 8'b00000000; // 3864 :   0 - 0x0
      13'hF19: dout  = 8'b00000000; // 3865 :   0 - 0x0
      13'hF1A: dout  = 8'b00000110; // 3866 :   6 - 0x6
      13'hF1B: dout  = 8'b00000110; // 3867 :   6 - 0x6
      13'hF1C: dout  = 8'b00001100; // 3868 :  12 - 0xc
      13'hF1D: dout  = 8'b00011000; // 3869 :  24 - 0x18
      13'hF1E: dout  = 8'b01110000; // 3870 : 112 - 0x70
      13'hF1F: dout  = 8'b01100000; // 3871 :  96 - 0x60
      13'hF20: dout  = 8'b11111111; // 3872 : 255 - 0xff -- Sprite 0xf2
      13'hF21: dout  = 8'b11111111; // 3873 : 255 - 0xff
      13'hF22: dout  = 8'b00000000; // 3874 :   0 - 0x0
      13'hF23: dout  = 8'b00000100; // 3875 :   4 - 0x4
      13'hF24: dout  = 8'b00000100; // 3876 :   4 - 0x4
      13'hF25: dout  = 8'b00000100; // 3877 :   4 - 0x4
      13'hF26: dout  = 8'b00001000; // 3878 :   8 - 0x8
      13'hF27: dout  = 8'b00001000; // 3879 :   8 - 0x8
      13'hF28: dout  = 8'b00000000; // 3880 :   0 - 0x0
      13'hF29: dout  = 8'b00000000; // 3881 :   0 - 0x0
      13'hF2A: dout  = 8'b00000110; // 3882 :   6 - 0x6
      13'hF2B: dout  = 8'b00000110; // 3883 :   6 - 0x6
      13'hF2C: dout  = 8'b00000100; // 3884 :   4 - 0x4
      13'hF2D: dout  = 8'b00000100; // 3885 :   4 - 0x4
      13'hF2E: dout  = 8'b00001000; // 3886 :   8 - 0x8
      13'hF2F: dout  = 8'b00001000; // 3887 :   8 - 0x8
      13'hF30: dout  = 8'b00001000; // 3888 :   8 - 0x8 -- Sprite 0xf3
      13'hF31: dout  = 8'b00010000; // 3889 :  16 - 0x10
      13'hF32: dout  = 8'b00010000; // 3890 :  16 - 0x10
      13'hF33: dout  = 8'b00000000; // 3891 :   0 - 0x0
      13'hF34: dout  = 8'b00000000; // 3892 :   0 - 0x0
      13'hF35: dout  = 8'b00010000; // 3893 :  16 - 0x10
      13'hF36: dout  = 8'b00010000; // 3894 :  16 - 0x10
      13'hF37: dout  = 8'b00001000; // 3895 :   8 - 0x8
      13'hF38: dout  = 8'b00001000; // 3896 :   8 - 0x8
      13'hF39: dout  = 8'b00010000; // 3897 :  16 - 0x10
      13'hF3A: dout  = 8'b00110000; // 3898 :  48 - 0x30
      13'hF3B: dout  = 8'b00110000; // 3899 :  48 - 0x30
      13'hF3C: dout  = 8'b00110000; // 3900 :  48 - 0x30
      13'hF3D: dout  = 8'b00110000; // 3901 :  48 - 0x30
      13'hF3E: dout  = 8'b00010000; // 3902 :  16 - 0x10
      13'hF3F: dout  = 8'b00001000; // 3903 :   8 - 0x8
      13'hF40: dout  = 8'b01111111; // 3904 : 127 - 0x7f -- Sprite 0xf4
      13'hF41: dout  = 8'b00111111; // 3905 :  63 - 0x3f
      13'hF42: dout  = 8'b00111111; // 3906 :  63 - 0x3f
      13'hF43: dout  = 8'b00111110; // 3907 :  62 - 0x3e
      13'hF44: dout  = 8'b00011111; // 3908 :  31 - 0x1f
      13'hF45: dout  = 8'b00001111; // 3909 :  15 - 0xf
      13'hF46: dout  = 8'b00000011; // 3910 :   3 - 0x3
      13'hF47: dout  = 8'b00000000; // 3911 :   0 - 0x0
      13'hF48: dout  = 8'b00000000; // 3912 :   0 - 0x0
      13'hF49: dout  = 8'b00000000; // 3913 :   0 - 0x0
      13'hF4A: dout  = 8'b00000001; // 3914 :   1 - 0x1
      13'hF4B: dout  = 8'b00000011; // 3915 :   3 - 0x3
      13'hF4C: dout  = 8'b00000001; // 3916 :   1 - 0x1
      13'hF4D: dout  = 8'b00000000; // 3917 :   0 - 0x0
      13'hF4E: dout  = 8'b00000000; // 3918 :   0 - 0x0
      13'hF4F: dout  = 8'b00000000; // 3919 :   0 - 0x0
      13'hF50: dout  = 8'b00000011; // 3920 :   3 - 0x3 -- Sprite 0xf5
      13'hF51: dout  = 8'b00001111; // 3921 :  15 - 0xf
      13'hF52: dout  = 8'b11111111; // 3922 : 255 - 0xff
      13'hF53: dout  = 8'b01111111; // 3923 : 127 - 0x7f
      13'hF54: dout  = 8'b01111111; // 3924 : 127 - 0x7f
      13'hF55: dout  = 8'b01111111; // 3925 : 127 - 0x7f
      13'hF56: dout  = 8'b01111111; // 3926 : 127 - 0x7f
      13'hF57: dout  = 8'b01111111; // 3927 : 127 - 0x7f
      13'hF58: dout  = 8'b00000011; // 3928 :   3 - 0x3
      13'hF59: dout  = 8'b00001110; // 3929 :  14 - 0xe
      13'hF5A: dout  = 8'b11111000; // 3930 : 248 - 0xf8
      13'hF5B: dout  = 8'b00000000; // 3931 :   0 - 0x0
      13'hF5C: dout  = 8'b00000000; // 3932 :   0 - 0x0
      13'hF5D: dout  = 8'b00000000; // 3933 :   0 - 0x0
      13'hF5E: dout  = 8'b00000000; // 3934 :   0 - 0x0
      13'hF5F: dout  = 8'b00000000; // 3935 :   0 - 0x0
      13'hF60: dout  = 8'b00000000; // 3936 :   0 - 0x0 -- Sprite 0xf6
      13'hF61: dout  = 8'b00000000; // 3937 :   0 - 0x0
      13'hF62: dout  = 8'b00000000; // 3938 :   0 - 0x0
      13'hF63: dout  = 8'b00000000; // 3939 :   0 - 0x0
      13'hF64: dout  = 8'b00000000; // 3940 :   0 - 0x0
      13'hF65: dout  = 8'b00000000; // 3941 :   0 - 0x0
      13'hF66: dout  = 8'b00000000; // 3942 :   0 - 0x0
      13'hF67: dout  = 8'b00000000; // 3943 :   0 - 0x0
      13'hF68: dout  = 8'b00100010; // 3944 :  34 - 0x22
      13'hF69: dout  = 8'b01100101; // 3945 : 101 - 0x65
      13'hF6A: dout  = 8'b00100101; // 3946 :  37 - 0x25
      13'hF6B: dout  = 8'b00100101; // 3947 :  37 - 0x25
      13'hF6C: dout  = 8'b00100101; // 3948 :  37 - 0x25
      13'hF6D: dout  = 8'b00100101; // 3949 :  37 - 0x25
      13'hF6E: dout  = 8'b01110111; // 3950 : 119 - 0x77
      13'hF6F: dout  = 8'b01110010; // 3951 : 114 - 0x72
      13'hF70: dout  = 8'b00000000; // 3952 :   0 - 0x0 -- Sprite 0xf7
      13'hF71: dout  = 8'b00000000; // 3953 :   0 - 0x0
      13'hF72: dout  = 8'b00000000; // 3954 :   0 - 0x0
      13'hF73: dout  = 8'b00000000; // 3955 :   0 - 0x0
      13'hF74: dout  = 8'b00000000; // 3956 :   0 - 0x0
      13'hF75: dout  = 8'b00000000; // 3957 :   0 - 0x0
      13'hF76: dout  = 8'b00000000; // 3958 :   0 - 0x0
      13'hF77: dout  = 8'b00000000; // 3959 :   0 - 0x0
      13'hF78: dout  = 8'b01100010; // 3960 :  98 - 0x62
      13'hF79: dout  = 8'b10010101; // 3961 : 149 - 0x95
      13'hF7A: dout  = 8'b00010101; // 3962 :  21 - 0x15
      13'hF7B: dout  = 8'b00100101; // 3963 :  37 - 0x25
      13'hF7C: dout  = 8'b01000101; // 3964 :  69 - 0x45
      13'hF7D: dout  = 8'b10000101; // 3965 : 133 - 0x85
      13'hF7E: dout  = 8'b11110111; // 3966 : 247 - 0xf7
      13'hF7F: dout  = 8'b11110010; // 3967 : 242 - 0xf2
      13'hF80: dout  = 8'b00000000; // 3968 :   0 - 0x0 -- Sprite 0xf8
      13'hF81: dout  = 8'b00000000; // 3969 :   0 - 0x0
      13'hF82: dout  = 8'b00000000; // 3970 :   0 - 0x0
      13'hF83: dout  = 8'b00000000; // 3971 :   0 - 0x0
      13'hF84: dout  = 8'b00000000; // 3972 :   0 - 0x0
      13'hF85: dout  = 8'b00000000; // 3973 :   0 - 0x0
      13'hF86: dout  = 8'b00000000; // 3974 :   0 - 0x0
      13'hF87: dout  = 8'b00000000; // 3975 :   0 - 0x0
      13'hF88: dout  = 8'b10100010; // 3976 : 162 - 0xa2
      13'hF89: dout  = 8'b10100101; // 3977 : 165 - 0xa5
      13'hF8A: dout  = 8'b10100101; // 3978 : 165 - 0xa5
      13'hF8B: dout  = 8'b10100101; // 3979 : 165 - 0xa5
      13'hF8C: dout  = 8'b11110101; // 3980 : 245 - 0xf5
      13'hF8D: dout  = 8'b11110101; // 3981 : 245 - 0xf5
      13'hF8E: dout  = 8'b00100111; // 3982 :  39 - 0x27
      13'hF8F: dout  = 8'b00100010; // 3983 :  34 - 0x22
      13'hF90: dout  = 8'b00000000; // 3984 :   0 - 0x0 -- Sprite 0xf9
      13'hF91: dout  = 8'b00000000; // 3985 :   0 - 0x0
      13'hF92: dout  = 8'b00000000; // 3986 :   0 - 0x0
      13'hF93: dout  = 8'b00000000; // 3987 :   0 - 0x0
      13'hF94: dout  = 8'b00000000; // 3988 :   0 - 0x0
      13'hF95: dout  = 8'b00000000; // 3989 :   0 - 0x0
      13'hF96: dout  = 8'b00000000; // 3990 :   0 - 0x0
      13'hF97: dout  = 8'b00000000; // 3991 :   0 - 0x0
      13'hF98: dout  = 8'b11110010; // 3992 : 242 - 0xf2
      13'hF99: dout  = 8'b10000101; // 3993 : 133 - 0x85
      13'hF9A: dout  = 8'b10000101; // 3994 : 133 - 0x85
      13'hF9B: dout  = 8'b11100101; // 3995 : 229 - 0xe5
      13'hF9C: dout  = 8'b00010101; // 3996 :  21 - 0x15
      13'hF9D: dout  = 8'b00010101; // 3997 :  21 - 0x15
      13'hF9E: dout  = 8'b11110111; // 3998 : 247 - 0xf7
      13'hF9F: dout  = 8'b11100010; // 3999 : 226 - 0xe2
      13'hFA0: dout  = 8'b00000000; // 4000 :   0 - 0x0 -- Sprite 0xfa
      13'hFA1: dout  = 8'b00000000; // 4001 :   0 - 0x0
      13'hFA2: dout  = 8'b00000000; // 4002 :   0 - 0x0
      13'hFA3: dout  = 8'b00000000; // 4003 :   0 - 0x0
      13'hFA4: dout  = 8'b00000000; // 4004 :   0 - 0x0
      13'hFA5: dout  = 8'b00000000; // 4005 :   0 - 0x0
      13'hFA6: dout  = 8'b00000000; // 4006 :   0 - 0x0
      13'hFA7: dout  = 8'b00000000; // 4007 :   0 - 0x0
      13'hFA8: dout  = 8'b01100010; // 4008 :  98 - 0x62
      13'hFA9: dout  = 8'b10010101; // 4009 : 149 - 0x95
      13'hFAA: dout  = 8'b01010101; // 4010 :  85 - 0x55
      13'hFAB: dout  = 8'b01100101; // 4011 : 101 - 0x65
      13'hFAC: dout  = 8'b10110101; // 4012 : 181 - 0xb5
      13'hFAD: dout  = 8'b10010101; // 4013 : 149 - 0x95
      13'hFAE: dout  = 8'b10010111; // 4014 : 151 - 0x97
      13'hFAF: dout  = 8'b01100010; // 4015 :  98 - 0x62
      13'hFB0: dout  = 8'b00000000; // 4016 :   0 - 0x0 -- Sprite 0xfb
      13'hFB1: dout  = 8'b00000000; // 4017 :   0 - 0x0
      13'hFB2: dout  = 8'b00000000; // 4018 :   0 - 0x0
      13'hFB3: dout  = 8'b00000000; // 4019 :   0 - 0x0
      13'hFB4: dout  = 8'b00000000; // 4020 :   0 - 0x0
      13'hFB5: dout  = 8'b00000000; // 4021 :   0 - 0x0
      13'hFB6: dout  = 8'b00000000; // 4022 :   0 - 0x0
      13'hFB7: dout  = 8'b00000000; // 4023 :   0 - 0x0
      13'hFB8: dout  = 8'b00100000; // 4024 :  32 - 0x20
      13'hFB9: dout  = 8'b01010000; // 4025 :  80 - 0x50
      13'hFBA: dout  = 8'b01010000; // 4026 :  80 - 0x50
      13'hFBB: dout  = 8'b01010000; // 4027 :  80 - 0x50
      13'hFBC: dout  = 8'b01010000; // 4028 :  80 - 0x50
      13'hFBD: dout  = 8'b01010000; // 4029 :  80 - 0x50
      13'hFBE: dout  = 8'b01110000; // 4030 : 112 - 0x70
      13'hFBF: dout  = 8'b00100000; // 4031 :  32 - 0x20
      13'hFC0: dout  = 8'b00000000; // 4032 :   0 - 0x0 -- Sprite 0xfc
      13'hFC1: dout  = 8'b00000000; // 4033 :   0 - 0x0
      13'hFC2: dout  = 8'b00000000; // 4034 :   0 - 0x0
      13'hFC3: dout  = 8'b00000000; // 4035 :   0 - 0x0
      13'hFC4: dout  = 8'b00000000; // 4036 :   0 - 0x0
      13'hFC5: dout  = 8'b00000000; // 4037 :   0 - 0x0
      13'hFC6: dout  = 8'b00000000; // 4038 :   0 - 0x0
      13'hFC7: dout  = 8'b00000000; // 4039 :   0 - 0x0
      13'hFC8: dout  = 8'b00000000; // 4040 :   0 - 0x0
      13'hFC9: dout  = 8'b00000000; // 4041 :   0 - 0x0
      13'hFCA: dout  = 8'b00000000; // 4042 :   0 - 0x0
      13'hFCB: dout  = 8'b00000000; // 4043 :   0 - 0x0
      13'hFCC: dout  = 8'b00000000; // 4044 :   0 - 0x0
      13'hFCD: dout  = 8'b00000000; // 4045 :   0 - 0x0
      13'hFCE: dout  = 8'b00000000; // 4046 :   0 - 0x0
      13'hFCF: dout  = 8'b00000000; // 4047 :   0 - 0x0
      13'hFD0: dout  = 8'b00000000; // 4048 :   0 - 0x0 -- Sprite 0xfd
      13'hFD1: dout  = 8'b00000000; // 4049 :   0 - 0x0
      13'hFD2: dout  = 8'b00000000; // 4050 :   0 - 0x0
      13'hFD3: dout  = 8'b00000000; // 4051 :   0 - 0x0
      13'hFD4: dout  = 8'b00000000; // 4052 :   0 - 0x0
      13'hFD5: dout  = 8'b00000000; // 4053 :   0 - 0x0
      13'hFD6: dout  = 8'b00000000; // 4054 :   0 - 0x0
      13'hFD7: dout  = 8'b00000000; // 4055 :   0 - 0x0
      13'hFD8: dout  = 8'b01100110; // 4056 : 102 - 0x66
      13'hFD9: dout  = 8'b11100110; // 4057 : 230 - 0xe6
      13'hFDA: dout  = 8'b01100110; // 4058 : 102 - 0x66
      13'hFDB: dout  = 8'b01100110; // 4059 : 102 - 0x66
      13'hFDC: dout  = 8'b01100110; // 4060 : 102 - 0x66
      13'hFDD: dout  = 8'b01100111; // 4061 : 103 - 0x67
      13'hFDE: dout  = 8'b11110011; // 4062 : 243 - 0xf3
      13'hFDF: dout  = 8'b00000000; // 4063 :   0 - 0x0
      13'hFE0: dout  = 8'b00000000; // 4064 :   0 - 0x0 -- Sprite 0xfe
      13'hFE1: dout  = 8'b00000000; // 4065 :   0 - 0x0
      13'hFE2: dout  = 8'b00000000; // 4066 :   0 - 0x0
      13'hFE3: dout  = 8'b00000000; // 4067 :   0 - 0x0
      13'hFE4: dout  = 8'b00000000; // 4068 :   0 - 0x0
      13'hFE5: dout  = 8'b00000000; // 4069 :   0 - 0x0
      13'hFE6: dout  = 8'b00000000; // 4070 :   0 - 0x0
      13'hFE7: dout  = 8'b00000000; // 4071 :   0 - 0x0
      13'hFE8: dout  = 8'b01011110; // 4072 :  94 - 0x5e
      13'hFE9: dout  = 8'b01011001; // 4073 :  89 - 0x59
      13'hFEA: dout  = 8'b01011001; // 4074 :  89 - 0x59
      13'hFEB: dout  = 8'b01011001; // 4075 :  89 - 0x59
      13'hFEC: dout  = 8'b01011110; // 4076 :  94 - 0x5e
      13'hFED: dout  = 8'b11011000; // 4077 : 216 - 0xd8
      13'hFEE: dout  = 8'b10011000; // 4078 : 152 - 0x98
      13'hFEF: dout  = 8'b00000000; // 4079 :   0 - 0x0
      13'hFF0: dout  = 8'b00000000; // 4080 :   0 - 0x0 -- Sprite 0xff
      13'hFF1: dout  = 8'b00000000; // 4081 :   0 - 0x0
      13'hFF2: dout  = 8'b00000000; // 4082 :   0 - 0x0
      13'hFF3: dout  = 8'b00000000; // 4083 :   0 - 0x0
      13'hFF4: dout  = 8'b00000000; // 4084 :   0 - 0x0
      13'hFF5: dout  = 8'b01111100; // 4085 : 124 - 0x7c
      13'hFF6: dout  = 8'b00111000; // 4086 :  56 - 0x38
      13'hFF7: dout  = 8'b00000000; // 4087 :   0 - 0x0
      13'hFF8: dout  = 8'b00000000; // 4088 :   0 - 0x0
      13'hFF9: dout  = 8'b00000000; // 4089 :   0 - 0x0
      13'hFFA: dout  = 8'b00000000; // 4090 :   0 - 0x0
      13'hFFB: dout  = 8'b00000000; // 4091 :   0 - 0x0
      13'hFFC: dout  = 8'b00000000; // 4092 :   0 - 0x0
      13'hFFD: dout  = 8'b00000100; // 4093 :   4 - 0x4
      13'hFFE: dout  = 8'b00001000; // 4094 :   8 - 0x8
      13'hFFF: dout  = 8'b00000000; // 4095 :   0 - 0x0
          // Pattern Table 1---------
      13'h1000: dout  = 8'b00111000; // 4096 :  56 - 0x38 -- Background 0x0
      13'h1001: dout  = 8'b01001100; // 4097 :  76 - 0x4c
      13'h1002: dout  = 8'b11000110; // 4098 : 198 - 0xc6
      13'h1003: dout  = 8'b11000110; // 4099 : 198 - 0xc6
      13'h1004: dout  = 8'b11000110; // 4100 : 198 - 0xc6
      13'h1005: dout  = 8'b01100100; // 4101 : 100 - 0x64
      13'h1006: dout  = 8'b00111000; // 4102 :  56 - 0x38
      13'h1007: dout  = 8'b00000000; // 4103 :   0 - 0x0
      13'h1008: dout  = 8'b00000000; // 4104 :   0 - 0x0
      13'h1009: dout  = 8'b00000000; // 4105 :   0 - 0x0
      13'h100A: dout  = 8'b00000000; // 4106 :   0 - 0x0
      13'h100B: dout  = 8'b00000000; // 4107 :   0 - 0x0
      13'h100C: dout  = 8'b00000000; // 4108 :   0 - 0x0
      13'h100D: dout  = 8'b00000000; // 4109 :   0 - 0x0
      13'h100E: dout  = 8'b00000000; // 4110 :   0 - 0x0
      13'h100F: dout  = 8'b00000000; // 4111 :   0 - 0x0
      13'h1010: dout  = 8'b00011000; // 4112 :  24 - 0x18 -- Background 0x1
      13'h1011: dout  = 8'b00111000; // 4113 :  56 - 0x38
      13'h1012: dout  = 8'b00011000; // 4114 :  24 - 0x18
      13'h1013: dout  = 8'b00011000; // 4115 :  24 - 0x18
      13'h1014: dout  = 8'b00011000; // 4116 :  24 - 0x18
      13'h1015: dout  = 8'b00011000; // 4117 :  24 - 0x18
      13'h1016: dout  = 8'b01111110; // 4118 : 126 - 0x7e
      13'h1017: dout  = 8'b00000000; // 4119 :   0 - 0x0
      13'h1018: dout  = 8'b00000000; // 4120 :   0 - 0x0
      13'h1019: dout  = 8'b00000000; // 4121 :   0 - 0x0
      13'h101A: dout  = 8'b00000000; // 4122 :   0 - 0x0
      13'h101B: dout  = 8'b00000000; // 4123 :   0 - 0x0
      13'h101C: dout  = 8'b00000000; // 4124 :   0 - 0x0
      13'h101D: dout  = 8'b00000000; // 4125 :   0 - 0x0
      13'h101E: dout  = 8'b00000000; // 4126 :   0 - 0x0
      13'h101F: dout  = 8'b00000000; // 4127 :   0 - 0x0
      13'h1020: dout  = 8'b01111100; // 4128 : 124 - 0x7c -- Background 0x2
      13'h1021: dout  = 8'b11000110; // 4129 : 198 - 0xc6
      13'h1022: dout  = 8'b00001110; // 4130 :  14 - 0xe
      13'h1023: dout  = 8'b00111100; // 4131 :  60 - 0x3c
      13'h1024: dout  = 8'b01111000; // 4132 : 120 - 0x78
      13'h1025: dout  = 8'b11100000; // 4133 : 224 - 0xe0
      13'h1026: dout  = 8'b11111110; // 4134 : 254 - 0xfe
      13'h1027: dout  = 8'b00000000; // 4135 :   0 - 0x0
      13'h1028: dout  = 8'b00000000; // 4136 :   0 - 0x0
      13'h1029: dout  = 8'b00000000; // 4137 :   0 - 0x0
      13'h102A: dout  = 8'b00000000; // 4138 :   0 - 0x0
      13'h102B: dout  = 8'b00000000; // 4139 :   0 - 0x0
      13'h102C: dout  = 8'b00000000; // 4140 :   0 - 0x0
      13'h102D: dout  = 8'b00000000; // 4141 :   0 - 0x0
      13'h102E: dout  = 8'b00000000; // 4142 :   0 - 0x0
      13'h102F: dout  = 8'b00000000; // 4143 :   0 - 0x0
      13'h1030: dout  = 8'b01111110; // 4144 : 126 - 0x7e -- Background 0x3
      13'h1031: dout  = 8'b00001100; // 4145 :  12 - 0xc
      13'h1032: dout  = 8'b00011000; // 4146 :  24 - 0x18
      13'h1033: dout  = 8'b00111100; // 4147 :  60 - 0x3c
      13'h1034: dout  = 8'b00000110; // 4148 :   6 - 0x6
      13'h1035: dout  = 8'b11000110; // 4149 : 198 - 0xc6
      13'h1036: dout  = 8'b01111100; // 4150 : 124 - 0x7c
      13'h1037: dout  = 8'b00000000; // 4151 :   0 - 0x0
      13'h1038: dout  = 8'b00000000; // 4152 :   0 - 0x0
      13'h1039: dout  = 8'b00000000; // 4153 :   0 - 0x0
      13'h103A: dout  = 8'b00000000; // 4154 :   0 - 0x0
      13'h103B: dout  = 8'b00000000; // 4155 :   0 - 0x0
      13'h103C: dout  = 8'b00000000; // 4156 :   0 - 0x0
      13'h103D: dout  = 8'b00000000; // 4157 :   0 - 0x0
      13'h103E: dout  = 8'b00000000; // 4158 :   0 - 0x0
      13'h103F: dout  = 8'b00000000; // 4159 :   0 - 0x0
      13'h1040: dout  = 8'b00011100; // 4160 :  28 - 0x1c -- Background 0x4
      13'h1041: dout  = 8'b00111100; // 4161 :  60 - 0x3c
      13'h1042: dout  = 8'b01101100; // 4162 : 108 - 0x6c
      13'h1043: dout  = 8'b11001100; // 4163 : 204 - 0xcc
      13'h1044: dout  = 8'b11111110; // 4164 : 254 - 0xfe
      13'h1045: dout  = 8'b00001100; // 4165 :  12 - 0xc
      13'h1046: dout  = 8'b00001100; // 4166 :  12 - 0xc
      13'h1047: dout  = 8'b00000000; // 4167 :   0 - 0x0
      13'h1048: dout  = 8'b00000000; // 4168 :   0 - 0x0
      13'h1049: dout  = 8'b00000000; // 4169 :   0 - 0x0
      13'h104A: dout  = 8'b00000000; // 4170 :   0 - 0x0
      13'h104B: dout  = 8'b00000000; // 4171 :   0 - 0x0
      13'h104C: dout  = 8'b00000000; // 4172 :   0 - 0x0
      13'h104D: dout  = 8'b00000000; // 4173 :   0 - 0x0
      13'h104E: dout  = 8'b00000000; // 4174 :   0 - 0x0
      13'h104F: dout  = 8'b00000000; // 4175 :   0 - 0x0
      13'h1050: dout  = 8'b11111100; // 4176 : 252 - 0xfc -- Background 0x5
      13'h1051: dout  = 8'b11000000; // 4177 : 192 - 0xc0
      13'h1052: dout  = 8'b11111100; // 4178 : 252 - 0xfc
      13'h1053: dout  = 8'b00000110; // 4179 :   6 - 0x6
      13'h1054: dout  = 8'b00000110; // 4180 :   6 - 0x6
      13'h1055: dout  = 8'b11000110; // 4181 : 198 - 0xc6
      13'h1056: dout  = 8'b01111100; // 4182 : 124 - 0x7c
      13'h1057: dout  = 8'b00000000; // 4183 :   0 - 0x0
      13'h1058: dout  = 8'b00000000; // 4184 :   0 - 0x0
      13'h1059: dout  = 8'b00000000; // 4185 :   0 - 0x0
      13'h105A: dout  = 8'b00000000; // 4186 :   0 - 0x0
      13'h105B: dout  = 8'b00000000; // 4187 :   0 - 0x0
      13'h105C: dout  = 8'b00000000; // 4188 :   0 - 0x0
      13'h105D: dout  = 8'b00000000; // 4189 :   0 - 0x0
      13'h105E: dout  = 8'b00000000; // 4190 :   0 - 0x0
      13'h105F: dout  = 8'b00000000; // 4191 :   0 - 0x0
      13'h1060: dout  = 8'b00111100; // 4192 :  60 - 0x3c -- Background 0x6
      13'h1061: dout  = 8'b01100000; // 4193 :  96 - 0x60
      13'h1062: dout  = 8'b11000000; // 4194 : 192 - 0xc0
      13'h1063: dout  = 8'b11111100; // 4195 : 252 - 0xfc
      13'h1064: dout  = 8'b11000110; // 4196 : 198 - 0xc6
      13'h1065: dout  = 8'b11000110; // 4197 : 198 - 0xc6
      13'h1066: dout  = 8'b01111100; // 4198 : 124 - 0x7c
      13'h1067: dout  = 8'b00000000; // 4199 :   0 - 0x0
      13'h1068: dout  = 8'b00000000; // 4200 :   0 - 0x0
      13'h1069: dout  = 8'b00000000; // 4201 :   0 - 0x0
      13'h106A: dout  = 8'b00000000; // 4202 :   0 - 0x0
      13'h106B: dout  = 8'b00000000; // 4203 :   0 - 0x0
      13'h106C: dout  = 8'b00000000; // 4204 :   0 - 0x0
      13'h106D: dout  = 8'b00000000; // 4205 :   0 - 0x0
      13'h106E: dout  = 8'b00000000; // 4206 :   0 - 0x0
      13'h106F: dout  = 8'b00000000; // 4207 :   0 - 0x0
      13'h1070: dout  = 8'b11111110; // 4208 : 254 - 0xfe -- Background 0x7
      13'h1071: dout  = 8'b11000110; // 4209 : 198 - 0xc6
      13'h1072: dout  = 8'b00001100; // 4210 :  12 - 0xc
      13'h1073: dout  = 8'b00011000; // 4211 :  24 - 0x18
      13'h1074: dout  = 8'b00110000; // 4212 :  48 - 0x30
      13'h1075: dout  = 8'b00110000; // 4213 :  48 - 0x30
      13'h1076: dout  = 8'b00110000; // 4214 :  48 - 0x30
      13'h1077: dout  = 8'b00000000; // 4215 :   0 - 0x0
      13'h1078: dout  = 8'b00000000; // 4216 :   0 - 0x0
      13'h1079: dout  = 8'b00000000; // 4217 :   0 - 0x0
      13'h107A: dout  = 8'b00000000; // 4218 :   0 - 0x0
      13'h107B: dout  = 8'b00000000; // 4219 :   0 - 0x0
      13'h107C: dout  = 8'b00000000; // 4220 :   0 - 0x0
      13'h107D: dout  = 8'b00000000; // 4221 :   0 - 0x0
      13'h107E: dout  = 8'b00000000; // 4222 :   0 - 0x0
      13'h107F: dout  = 8'b00000000; // 4223 :   0 - 0x0
      13'h1080: dout  = 8'b01111100; // 4224 : 124 - 0x7c -- Background 0x8
      13'h1081: dout  = 8'b11000110; // 4225 : 198 - 0xc6
      13'h1082: dout  = 8'b11000110; // 4226 : 198 - 0xc6
      13'h1083: dout  = 8'b01111100; // 4227 : 124 - 0x7c
      13'h1084: dout  = 8'b11000110; // 4228 : 198 - 0xc6
      13'h1085: dout  = 8'b11000110; // 4229 : 198 - 0xc6
      13'h1086: dout  = 8'b01111100; // 4230 : 124 - 0x7c
      13'h1087: dout  = 8'b00000000; // 4231 :   0 - 0x0
      13'h1088: dout  = 8'b00000000; // 4232 :   0 - 0x0
      13'h1089: dout  = 8'b00000000; // 4233 :   0 - 0x0
      13'h108A: dout  = 8'b00000000; // 4234 :   0 - 0x0
      13'h108B: dout  = 8'b00000000; // 4235 :   0 - 0x0
      13'h108C: dout  = 8'b00000000; // 4236 :   0 - 0x0
      13'h108D: dout  = 8'b00000000; // 4237 :   0 - 0x0
      13'h108E: dout  = 8'b00000000; // 4238 :   0 - 0x0
      13'h108F: dout  = 8'b00000000; // 4239 :   0 - 0x0
      13'h1090: dout  = 8'b01111100; // 4240 : 124 - 0x7c -- Background 0x9
      13'h1091: dout  = 8'b11000110; // 4241 : 198 - 0xc6
      13'h1092: dout  = 8'b11000110; // 4242 : 198 - 0xc6
      13'h1093: dout  = 8'b01111110; // 4243 : 126 - 0x7e
      13'h1094: dout  = 8'b00000110; // 4244 :   6 - 0x6
      13'h1095: dout  = 8'b00001100; // 4245 :  12 - 0xc
      13'h1096: dout  = 8'b01111000; // 4246 : 120 - 0x78
      13'h1097: dout  = 8'b00000000; // 4247 :   0 - 0x0
      13'h1098: dout  = 8'b00000000; // 4248 :   0 - 0x0
      13'h1099: dout  = 8'b00000000; // 4249 :   0 - 0x0
      13'h109A: dout  = 8'b00000000; // 4250 :   0 - 0x0
      13'h109B: dout  = 8'b00000000; // 4251 :   0 - 0x0
      13'h109C: dout  = 8'b00000000; // 4252 :   0 - 0x0
      13'h109D: dout  = 8'b00000000; // 4253 :   0 - 0x0
      13'h109E: dout  = 8'b00000000; // 4254 :   0 - 0x0
      13'h109F: dout  = 8'b00000000; // 4255 :   0 - 0x0
      13'h10A0: dout  = 8'b00111000; // 4256 :  56 - 0x38 -- Background 0xa
      13'h10A1: dout  = 8'b01101100; // 4257 : 108 - 0x6c
      13'h10A2: dout  = 8'b11000110; // 4258 : 198 - 0xc6
      13'h10A3: dout  = 8'b11000110; // 4259 : 198 - 0xc6
      13'h10A4: dout  = 8'b11111110; // 4260 : 254 - 0xfe
      13'h10A5: dout  = 8'b11000110; // 4261 : 198 - 0xc6
      13'h10A6: dout  = 8'b11000110; // 4262 : 198 - 0xc6
      13'h10A7: dout  = 8'b00000000; // 4263 :   0 - 0x0
      13'h10A8: dout  = 8'b00000000; // 4264 :   0 - 0x0
      13'h10A9: dout  = 8'b00000000; // 4265 :   0 - 0x0
      13'h10AA: dout  = 8'b00000000; // 4266 :   0 - 0x0
      13'h10AB: dout  = 8'b00000000; // 4267 :   0 - 0x0
      13'h10AC: dout  = 8'b00000000; // 4268 :   0 - 0x0
      13'h10AD: dout  = 8'b00000000; // 4269 :   0 - 0x0
      13'h10AE: dout  = 8'b00000000; // 4270 :   0 - 0x0
      13'h10AF: dout  = 8'b00000000; // 4271 :   0 - 0x0
      13'h10B0: dout  = 8'b11111100; // 4272 : 252 - 0xfc -- Background 0xb
      13'h10B1: dout  = 8'b11000110; // 4273 : 198 - 0xc6
      13'h10B2: dout  = 8'b11000110; // 4274 : 198 - 0xc6
      13'h10B3: dout  = 8'b11111100; // 4275 : 252 - 0xfc
      13'h10B4: dout  = 8'b11000110; // 4276 : 198 - 0xc6
      13'h10B5: dout  = 8'b11000110; // 4277 : 198 - 0xc6
      13'h10B6: dout  = 8'b11111100; // 4278 : 252 - 0xfc
      13'h10B7: dout  = 8'b00000000; // 4279 :   0 - 0x0
      13'h10B8: dout  = 8'b00000000; // 4280 :   0 - 0x0
      13'h10B9: dout  = 8'b00000000; // 4281 :   0 - 0x0
      13'h10BA: dout  = 8'b00000000; // 4282 :   0 - 0x0
      13'h10BB: dout  = 8'b00000000; // 4283 :   0 - 0x0
      13'h10BC: dout  = 8'b00000000; // 4284 :   0 - 0x0
      13'h10BD: dout  = 8'b00000000; // 4285 :   0 - 0x0
      13'h10BE: dout  = 8'b00000000; // 4286 :   0 - 0x0
      13'h10BF: dout  = 8'b00000000; // 4287 :   0 - 0x0
      13'h10C0: dout  = 8'b00111100; // 4288 :  60 - 0x3c -- Background 0xc
      13'h10C1: dout  = 8'b01100110; // 4289 : 102 - 0x66
      13'h10C2: dout  = 8'b11000000; // 4290 : 192 - 0xc0
      13'h10C3: dout  = 8'b11000000; // 4291 : 192 - 0xc0
      13'h10C4: dout  = 8'b11000000; // 4292 : 192 - 0xc0
      13'h10C5: dout  = 8'b01100110; // 4293 : 102 - 0x66
      13'h10C6: dout  = 8'b00111100; // 4294 :  60 - 0x3c
      13'h10C7: dout  = 8'b00000000; // 4295 :   0 - 0x0
      13'h10C8: dout  = 8'b00000000; // 4296 :   0 - 0x0
      13'h10C9: dout  = 8'b00000000; // 4297 :   0 - 0x0
      13'h10CA: dout  = 8'b00000000; // 4298 :   0 - 0x0
      13'h10CB: dout  = 8'b00000000; // 4299 :   0 - 0x0
      13'h10CC: dout  = 8'b00000000; // 4300 :   0 - 0x0
      13'h10CD: dout  = 8'b00000000; // 4301 :   0 - 0x0
      13'h10CE: dout  = 8'b00000000; // 4302 :   0 - 0x0
      13'h10CF: dout  = 8'b00000000; // 4303 :   0 - 0x0
      13'h10D0: dout  = 8'b11111000; // 4304 : 248 - 0xf8 -- Background 0xd
      13'h10D1: dout  = 8'b11001100; // 4305 : 204 - 0xcc
      13'h10D2: dout  = 8'b11000110; // 4306 : 198 - 0xc6
      13'h10D3: dout  = 8'b11000110; // 4307 : 198 - 0xc6
      13'h10D4: dout  = 8'b11000110; // 4308 : 198 - 0xc6
      13'h10D5: dout  = 8'b11001100; // 4309 : 204 - 0xcc
      13'h10D6: dout  = 8'b11111000; // 4310 : 248 - 0xf8
      13'h10D7: dout  = 8'b00000000; // 4311 :   0 - 0x0
      13'h10D8: dout  = 8'b00000000; // 4312 :   0 - 0x0
      13'h10D9: dout  = 8'b00000000; // 4313 :   0 - 0x0
      13'h10DA: dout  = 8'b00000000; // 4314 :   0 - 0x0
      13'h10DB: dout  = 8'b00000000; // 4315 :   0 - 0x0
      13'h10DC: dout  = 8'b00000000; // 4316 :   0 - 0x0
      13'h10DD: dout  = 8'b00000000; // 4317 :   0 - 0x0
      13'h10DE: dout  = 8'b00000000; // 4318 :   0 - 0x0
      13'h10DF: dout  = 8'b00000000; // 4319 :   0 - 0x0
      13'h10E0: dout  = 8'b11111110; // 4320 : 254 - 0xfe -- Background 0xe
      13'h10E1: dout  = 8'b11000000; // 4321 : 192 - 0xc0
      13'h10E2: dout  = 8'b11000000; // 4322 : 192 - 0xc0
      13'h10E3: dout  = 8'b11111100; // 4323 : 252 - 0xfc
      13'h10E4: dout  = 8'b11000000; // 4324 : 192 - 0xc0
      13'h10E5: dout  = 8'b11000000; // 4325 : 192 - 0xc0
      13'h10E6: dout  = 8'b11111110; // 4326 : 254 - 0xfe
      13'h10E7: dout  = 8'b00000000; // 4327 :   0 - 0x0
      13'h10E8: dout  = 8'b00000000; // 4328 :   0 - 0x0
      13'h10E9: dout  = 8'b00000000; // 4329 :   0 - 0x0
      13'h10EA: dout  = 8'b00000000; // 4330 :   0 - 0x0
      13'h10EB: dout  = 8'b00000000; // 4331 :   0 - 0x0
      13'h10EC: dout  = 8'b00000000; // 4332 :   0 - 0x0
      13'h10ED: dout  = 8'b00000000; // 4333 :   0 - 0x0
      13'h10EE: dout  = 8'b00000000; // 4334 :   0 - 0x0
      13'h10EF: dout  = 8'b00000000; // 4335 :   0 - 0x0
      13'h10F0: dout  = 8'b11111110; // 4336 : 254 - 0xfe -- Background 0xf
      13'h10F1: dout  = 8'b11000000; // 4337 : 192 - 0xc0
      13'h10F2: dout  = 8'b11000000; // 4338 : 192 - 0xc0
      13'h10F3: dout  = 8'b11111100; // 4339 : 252 - 0xfc
      13'h10F4: dout  = 8'b11000000; // 4340 : 192 - 0xc0
      13'h10F5: dout  = 8'b11000000; // 4341 : 192 - 0xc0
      13'h10F6: dout  = 8'b11000000; // 4342 : 192 - 0xc0
      13'h10F7: dout  = 8'b00000000; // 4343 :   0 - 0x0
      13'h10F8: dout  = 8'b00000000; // 4344 :   0 - 0x0
      13'h10F9: dout  = 8'b00000000; // 4345 :   0 - 0x0
      13'h10FA: dout  = 8'b00000000; // 4346 :   0 - 0x0
      13'h10FB: dout  = 8'b00000000; // 4347 :   0 - 0x0
      13'h10FC: dout  = 8'b00000000; // 4348 :   0 - 0x0
      13'h10FD: dout  = 8'b00000000; // 4349 :   0 - 0x0
      13'h10FE: dout  = 8'b00000000; // 4350 :   0 - 0x0
      13'h10FF: dout  = 8'b00000000; // 4351 :   0 - 0x0
      13'h1100: dout  = 8'b00111110; // 4352 :  62 - 0x3e -- Background 0x10
      13'h1101: dout  = 8'b01100000; // 4353 :  96 - 0x60
      13'h1102: dout  = 8'b11000000; // 4354 : 192 - 0xc0
      13'h1103: dout  = 8'b11001110; // 4355 : 206 - 0xce
      13'h1104: dout  = 8'b11000110; // 4356 : 198 - 0xc6
      13'h1105: dout  = 8'b01100110; // 4357 : 102 - 0x66
      13'h1106: dout  = 8'b00111110; // 4358 :  62 - 0x3e
      13'h1107: dout  = 8'b00000000; // 4359 :   0 - 0x0
      13'h1108: dout  = 8'b00000000; // 4360 :   0 - 0x0
      13'h1109: dout  = 8'b00000000; // 4361 :   0 - 0x0
      13'h110A: dout  = 8'b00000000; // 4362 :   0 - 0x0
      13'h110B: dout  = 8'b00000000; // 4363 :   0 - 0x0
      13'h110C: dout  = 8'b00000000; // 4364 :   0 - 0x0
      13'h110D: dout  = 8'b00000000; // 4365 :   0 - 0x0
      13'h110E: dout  = 8'b00000000; // 4366 :   0 - 0x0
      13'h110F: dout  = 8'b00000000; // 4367 :   0 - 0x0
      13'h1110: dout  = 8'b11000110; // 4368 : 198 - 0xc6 -- Background 0x11
      13'h1111: dout  = 8'b11000110; // 4369 : 198 - 0xc6
      13'h1112: dout  = 8'b11000110; // 4370 : 198 - 0xc6
      13'h1113: dout  = 8'b11111110; // 4371 : 254 - 0xfe
      13'h1114: dout  = 8'b11000110; // 4372 : 198 - 0xc6
      13'h1115: dout  = 8'b11000110; // 4373 : 198 - 0xc6
      13'h1116: dout  = 8'b11000110; // 4374 : 198 - 0xc6
      13'h1117: dout  = 8'b00000000; // 4375 :   0 - 0x0
      13'h1118: dout  = 8'b00000000; // 4376 :   0 - 0x0
      13'h1119: dout  = 8'b00000000; // 4377 :   0 - 0x0
      13'h111A: dout  = 8'b00000000; // 4378 :   0 - 0x0
      13'h111B: dout  = 8'b00000000; // 4379 :   0 - 0x0
      13'h111C: dout  = 8'b00000000; // 4380 :   0 - 0x0
      13'h111D: dout  = 8'b00000000; // 4381 :   0 - 0x0
      13'h111E: dout  = 8'b00000000; // 4382 :   0 - 0x0
      13'h111F: dout  = 8'b00000000; // 4383 :   0 - 0x0
      13'h1120: dout  = 8'b01111110; // 4384 : 126 - 0x7e -- Background 0x12
      13'h1121: dout  = 8'b00011000; // 4385 :  24 - 0x18
      13'h1122: dout  = 8'b00011000; // 4386 :  24 - 0x18
      13'h1123: dout  = 8'b00011000; // 4387 :  24 - 0x18
      13'h1124: dout  = 8'b00011000; // 4388 :  24 - 0x18
      13'h1125: dout  = 8'b00011000; // 4389 :  24 - 0x18
      13'h1126: dout  = 8'b01111110; // 4390 : 126 - 0x7e
      13'h1127: dout  = 8'b00000000; // 4391 :   0 - 0x0
      13'h1128: dout  = 8'b00000000; // 4392 :   0 - 0x0
      13'h1129: dout  = 8'b00000000; // 4393 :   0 - 0x0
      13'h112A: dout  = 8'b00000000; // 4394 :   0 - 0x0
      13'h112B: dout  = 8'b00000000; // 4395 :   0 - 0x0
      13'h112C: dout  = 8'b00000000; // 4396 :   0 - 0x0
      13'h112D: dout  = 8'b00000000; // 4397 :   0 - 0x0
      13'h112E: dout  = 8'b00000000; // 4398 :   0 - 0x0
      13'h112F: dout  = 8'b00000000; // 4399 :   0 - 0x0
      13'h1130: dout  = 8'b00011110; // 4400 :  30 - 0x1e -- Background 0x13
      13'h1131: dout  = 8'b00000110; // 4401 :   6 - 0x6
      13'h1132: dout  = 8'b00000110; // 4402 :   6 - 0x6
      13'h1133: dout  = 8'b00000110; // 4403 :   6 - 0x6
      13'h1134: dout  = 8'b11000110; // 4404 : 198 - 0xc6
      13'h1135: dout  = 8'b11000110; // 4405 : 198 - 0xc6
      13'h1136: dout  = 8'b01111100; // 4406 : 124 - 0x7c
      13'h1137: dout  = 8'b00000000; // 4407 :   0 - 0x0
      13'h1138: dout  = 8'b00000000; // 4408 :   0 - 0x0
      13'h1139: dout  = 8'b00000000; // 4409 :   0 - 0x0
      13'h113A: dout  = 8'b00000000; // 4410 :   0 - 0x0
      13'h113B: dout  = 8'b00000000; // 4411 :   0 - 0x0
      13'h113C: dout  = 8'b00000000; // 4412 :   0 - 0x0
      13'h113D: dout  = 8'b00000000; // 4413 :   0 - 0x0
      13'h113E: dout  = 8'b00000000; // 4414 :   0 - 0x0
      13'h113F: dout  = 8'b00000000; // 4415 :   0 - 0x0
      13'h1140: dout  = 8'b11000110; // 4416 : 198 - 0xc6 -- Background 0x14
      13'h1141: dout  = 8'b11001100; // 4417 : 204 - 0xcc
      13'h1142: dout  = 8'b11011000; // 4418 : 216 - 0xd8
      13'h1143: dout  = 8'b11110000; // 4419 : 240 - 0xf0
      13'h1144: dout  = 8'b11111000; // 4420 : 248 - 0xf8
      13'h1145: dout  = 8'b11011100; // 4421 : 220 - 0xdc
      13'h1146: dout  = 8'b11001110; // 4422 : 206 - 0xce
      13'h1147: dout  = 8'b00000000; // 4423 :   0 - 0x0
      13'h1148: dout  = 8'b00000000; // 4424 :   0 - 0x0
      13'h1149: dout  = 8'b00000000; // 4425 :   0 - 0x0
      13'h114A: dout  = 8'b00000000; // 4426 :   0 - 0x0
      13'h114B: dout  = 8'b00000000; // 4427 :   0 - 0x0
      13'h114C: dout  = 8'b00000000; // 4428 :   0 - 0x0
      13'h114D: dout  = 8'b00000000; // 4429 :   0 - 0x0
      13'h114E: dout  = 8'b00000000; // 4430 :   0 - 0x0
      13'h114F: dout  = 8'b00000000; // 4431 :   0 - 0x0
      13'h1150: dout  = 8'b01100000; // 4432 :  96 - 0x60 -- Background 0x15
      13'h1151: dout  = 8'b01100000; // 4433 :  96 - 0x60
      13'h1152: dout  = 8'b01100000; // 4434 :  96 - 0x60
      13'h1153: dout  = 8'b01100000; // 4435 :  96 - 0x60
      13'h1154: dout  = 8'b01100000; // 4436 :  96 - 0x60
      13'h1155: dout  = 8'b01100000; // 4437 :  96 - 0x60
      13'h1156: dout  = 8'b01111110; // 4438 : 126 - 0x7e
      13'h1157: dout  = 8'b00000000; // 4439 :   0 - 0x0
      13'h1158: dout  = 8'b00000000; // 4440 :   0 - 0x0
      13'h1159: dout  = 8'b00000000; // 4441 :   0 - 0x0
      13'h115A: dout  = 8'b00000000; // 4442 :   0 - 0x0
      13'h115B: dout  = 8'b00000000; // 4443 :   0 - 0x0
      13'h115C: dout  = 8'b00000000; // 4444 :   0 - 0x0
      13'h115D: dout  = 8'b00000000; // 4445 :   0 - 0x0
      13'h115E: dout  = 8'b00000000; // 4446 :   0 - 0x0
      13'h115F: dout  = 8'b00000000; // 4447 :   0 - 0x0
      13'h1160: dout  = 8'b11000110; // 4448 : 198 - 0xc6 -- Background 0x16
      13'h1161: dout  = 8'b11101110; // 4449 : 238 - 0xee
      13'h1162: dout  = 8'b11111110; // 4450 : 254 - 0xfe
      13'h1163: dout  = 8'b11111110; // 4451 : 254 - 0xfe
      13'h1164: dout  = 8'b11010110; // 4452 : 214 - 0xd6
      13'h1165: dout  = 8'b11000110; // 4453 : 198 - 0xc6
      13'h1166: dout  = 8'b11000110; // 4454 : 198 - 0xc6
      13'h1167: dout  = 8'b00000000; // 4455 :   0 - 0x0
      13'h1168: dout  = 8'b00000000; // 4456 :   0 - 0x0
      13'h1169: dout  = 8'b00000000; // 4457 :   0 - 0x0
      13'h116A: dout  = 8'b00000000; // 4458 :   0 - 0x0
      13'h116B: dout  = 8'b00000000; // 4459 :   0 - 0x0
      13'h116C: dout  = 8'b00000000; // 4460 :   0 - 0x0
      13'h116D: dout  = 8'b00000000; // 4461 :   0 - 0x0
      13'h116E: dout  = 8'b00000000; // 4462 :   0 - 0x0
      13'h116F: dout  = 8'b00000000; // 4463 :   0 - 0x0
      13'h1170: dout  = 8'b11000110; // 4464 : 198 - 0xc6 -- Background 0x17
      13'h1171: dout  = 8'b11100110; // 4465 : 230 - 0xe6
      13'h1172: dout  = 8'b11110110; // 4466 : 246 - 0xf6
      13'h1173: dout  = 8'b11111110; // 4467 : 254 - 0xfe
      13'h1174: dout  = 8'b11011110; // 4468 : 222 - 0xde
      13'h1175: dout  = 8'b11001110; // 4469 : 206 - 0xce
      13'h1176: dout  = 8'b11000110; // 4470 : 198 - 0xc6
      13'h1177: dout  = 8'b00000000; // 4471 :   0 - 0x0
      13'h1178: dout  = 8'b00000000; // 4472 :   0 - 0x0
      13'h1179: dout  = 8'b00000000; // 4473 :   0 - 0x0
      13'h117A: dout  = 8'b00000000; // 4474 :   0 - 0x0
      13'h117B: dout  = 8'b00000000; // 4475 :   0 - 0x0
      13'h117C: dout  = 8'b00000000; // 4476 :   0 - 0x0
      13'h117D: dout  = 8'b00000000; // 4477 :   0 - 0x0
      13'h117E: dout  = 8'b00000000; // 4478 :   0 - 0x0
      13'h117F: dout  = 8'b00000000; // 4479 :   0 - 0x0
      13'h1180: dout  = 8'b01111100; // 4480 : 124 - 0x7c -- Background 0x18
      13'h1181: dout  = 8'b11000110; // 4481 : 198 - 0xc6
      13'h1182: dout  = 8'b11000110; // 4482 : 198 - 0xc6
      13'h1183: dout  = 8'b11000110; // 4483 : 198 - 0xc6
      13'h1184: dout  = 8'b11000110; // 4484 : 198 - 0xc6
      13'h1185: dout  = 8'b11000110; // 4485 : 198 - 0xc6
      13'h1186: dout  = 8'b01111100; // 4486 : 124 - 0x7c
      13'h1187: dout  = 8'b00000000; // 4487 :   0 - 0x0
      13'h1188: dout  = 8'b00000000; // 4488 :   0 - 0x0
      13'h1189: dout  = 8'b00000000; // 4489 :   0 - 0x0
      13'h118A: dout  = 8'b00000000; // 4490 :   0 - 0x0
      13'h118B: dout  = 8'b00000000; // 4491 :   0 - 0x0
      13'h118C: dout  = 8'b00000000; // 4492 :   0 - 0x0
      13'h118D: dout  = 8'b00000000; // 4493 :   0 - 0x0
      13'h118E: dout  = 8'b00000000; // 4494 :   0 - 0x0
      13'h118F: dout  = 8'b00000000; // 4495 :   0 - 0x0
      13'h1190: dout  = 8'b11111100; // 4496 : 252 - 0xfc -- Background 0x19
      13'h1191: dout  = 8'b11000110; // 4497 : 198 - 0xc6
      13'h1192: dout  = 8'b11000110; // 4498 : 198 - 0xc6
      13'h1193: dout  = 8'b11000110; // 4499 : 198 - 0xc6
      13'h1194: dout  = 8'b11111100; // 4500 : 252 - 0xfc
      13'h1195: dout  = 8'b11000000; // 4501 : 192 - 0xc0
      13'h1196: dout  = 8'b11000000; // 4502 : 192 - 0xc0
      13'h1197: dout  = 8'b00000000; // 4503 :   0 - 0x0
      13'h1198: dout  = 8'b00000000; // 4504 :   0 - 0x0
      13'h1199: dout  = 8'b00000000; // 4505 :   0 - 0x0
      13'h119A: dout  = 8'b00000000; // 4506 :   0 - 0x0
      13'h119B: dout  = 8'b00000000; // 4507 :   0 - 0x0
      13'h119C: dout  = 8'b00000000; // 4508 :   0 - 0x0
      13'h119D: dout  = 8'b00000000; // 4509 :   0 - 0x0
      13'h119E: dout  = 8'b00000000; // 4510 :   0 - 0x0
      13'h119F: dout  = 8'b00000000; // 4511 :   0 - 0x0
      13'h11A0: dout  = 8'b01111100; // 4512 : 124 - 0x7c -- Background 0x1a
      13'h11A1: dout  = 8'b11000110; // 4513 : 198 - 0xc6
      13'h11A2: dout  = 8'b11000110; // 4514 : 198 - 0xc6
      13'h11A3: dout  = 8'b11000110; // 4515 : 198 - 0xc6
      13'h11A4: dout  = 8'b11011110; // 4516 : 222 - 0xde
      13'h11A5: dout  = 8'b11001100; // 4517 : 204 - 0xcc
      13'h11A6: dout  = 8'b01111010; // 4518 : 122 - 0x7a
      13'h11A7: dout  = 8'b00000000; // 4519 :   0 - 0x0
      13'h11A8: dout  = 8'b00000000; // 4520 :   0 - 0x0
      13'h11A9: dout  = 8'b00000000; // 4521 :   0 - 0x0
      13'h11AA: dout  = 8'b00000000; // 4522 :   0 - 0x0
      13'h11AB: dout  = 8'b00000000; // 4523 :   0 - 0x0
      13'h11AC: dout  = 8'b00000000; // 4524 :   0 - 0x0
      13'h11AD: dout  = 8'b00000000; // 4525 :   0 - 0x0
      13'h11AE: dout  = 8'b00000000; // 4526 :   0 - 0x0
      13'h11AF: dout  = 8'b00000000; // 4527 :   0 - 0x0
      13'h11B0: dout  = 8'b11111100; // 4528 : 252 - 0xfc -- Background 0x1b
      13'h11B1: dout  = 8'b11000110; // 4529 : 198 - 0xc6
      13'h11B2: dout  = 8'b11000110; // 4530 : 198 - 0xc6
      13'h11B3: dout  = 8'b11001110; // 4531 : 206 - 0xce
      13'h11B4: dout  = 8'b11111000; // 4532 : 248 - 0xf8
      13'h11B5: dout  = 8'b11011100; // 4533 : 220 - 0xdc
      13'h11B6: dout  = 8'b11001110; // 4534 : 206 - 0xce
      13'h11B7: dout  = 8'b00000000; // 4535 :   0 - 0x0
      13'h11B8: dout  = 8'b00000000; // 4536 :   0 - 0x0
      13'h11B9: dout  = 8'b00000000; // 4537 :   0 - 0x0
      13'h11BA: dout  = 8'b00000000; // 4538 :   0 - 0x0
      13'h11BB: dout  = 8'b00000000; // 4539 :   0 - 0x0
      13'h11BC: dout  = 8'b00000000; // 4540 :   0 - 0x0
      13'h11BD: dout  = 8'b00000000; // 4541 :   0 - 0x0
      13'h11BE: dout  = 8'b00000000; // 4542 :   0 - 0x0
      13'h11BF: dout  = 8'b00000000; // 4543 :   0 - 0x0
      13'h11C0: dout  = 8'b01111000; // 4544 : 120 - 0x78 -- Background 0x1c
      13'h11C1: dout  = 8'b11001100; // 4545 : 204 - 0xcc
      13'h11C2: dout  = 8'b11000000; // 4546 : 192 - 0xc0
      13'h11C3: dout  = 8'b01111100; // 4547 : 124 - 0x7c
      13'h11C4: dout  = 8'b00000110; // 4548 :   6 - 0x6
      13'h11C5: dout  = 8'b11000110; // 4549 : 198 - 0xc6
      13'h11C6: dout  = 8'b01111100; // 4550 : 124 - 0x7c
      13'h11C7: dout  = 8'b00000000; // 4551 :   0 - 0x0
      13'h11C8: dout  = 8'b00000000; // 4552 :   0 - 0x0
      13'h11C9: dout  = 8'b00000000; // 4553 :   0 - 0x0
      13'h11CA: dout  = 8'b00000000; // 4554 :   0 - 0x0
      13'h11CB: dout  = 8'b00000000; // 4555 :   0 - 0x0
      13'h11CC: dout  = 8'b00000000; // 4556 :   0 - 0x0
      13'h11CD: dout  = 8'b00000000; // 4557 :   0 - 0x0
      13'h11CE: dout  = 8'b00000000; // 4558 :   0 - 0x0
      13'h11CF: dout  = 8'b00000000; // 4559 :   0 - 0x0
      13'h11D0: dout  = 8'b01111110; // 4560 : 126 - 0x7e -- Background 0x1d
      13'h11D1: dout  = 8'b00011000; // 4561 :  24 - 0x18
      13'h11D2: dout  = 8'b00011000; // 4562 :  24 - 0x18
      13'h11D3: dout  = 8'b00011000; // 4563 :  24 - 0x18
      13'h11D4: dout  = 8'b00011000; // 4564 :  24 - 0x18
      13'h11D5: dout  = 8'b00011000; // 4565 :  24 - 0x18
      13'h11D6: dout  = 8'b00011000; // 4566 :  24 - 0x18
      13'h11D7: dout  = 8'b00000000; // 4567 :   0 - 0x0
      13'h11D8: dout  = 8'b00000000; // 4568 :   0 - 0x0
      13'h11D9: dout  = 8'b00000000; // 4569 :   0 - 0x0
      13'h11DA: dout  = 8'b00000000; // 4570 :   0 - 0x0
      13'h11DB: dout  = 8'b00000000; // 4571 :   0 - 0x0
      13'h11DC: dout  = 8'b00000000; // 4572 :   0 - 0x0
      13'h11DD: dout  = 8'b00000000; // 4573 :   0 - 0x0
      13'h11DE: dout  = 8'b00000000; // 4574 :   0 - 0x0
      13'h11DF: dout  = 8'b00000000; // 4575 :   0 - 0x0
      13'h11E0: dout  = 8'b11000110; // 4576 : 198 - 0xc6 -- Background 0x1e
      13'h11E1: dout  = 8'b11000110; // 4577 : 198 - 0xc6
      13'h11E2: dout  = 8'b11000110; // 4578 : 198 - 0xc6
      13'h11E3: dout  = 8'b11000110; // 4579 : 198 - 0xc6
      13'h11E4: dout  = 8'b11000110; // 4580 : 198 - 0xc6
      13'h11E5: dout  = 8'b11000110; // 4581 : 198 - 0xc6
      13'h11E6: dout  = 8'b01111100; // 4582 : 124 - 0x7c
      13'h11E7: dout  = 8'b00000000; // 4583 :   0 - 0x0
      13'h11E8: dout  = 8'b00000000; // 4584 :   0 - 0x0
      13'h11E9: dout  = 8'b00000000; // 4585 :   0 - 0x0
      13'h11EA: dout  = 8'b00000000; // 4586 :   0 - 0x0
      13'h11EB: dout  = 8'b00000000; // 4587 :   0 - 0x0
      13'h11EC: dout  = 8'b00000000; // 4588 :   0 - 0x0
      13'h11ED: dout  = 8'b00000000; // 4589 :   0 - 0x0
      13'h11EE: dout  = 8'b00000000; // 4590 :   0 - 0x0
      13'h11EF: dout  = 8'b00000000; // 4591 :   0 - 0x0
      13'h11F0: dout  = 8'b11000110; // 4592 : 198 - 0xc6 -- Background 0x1f
      13'h11F1: dout  = 8'b11000110; // 4593 : 198 - 0xc6
      13'h11F2: dout  = 8'b11000110; // 4594 : 198 - 0xc6
      13'h11F3: dout  = 8'b11101110; // 4595 : 238 - 0xee
      13'h11F4: dout  = 8'b01111100; // 4596 : 124 - 0x7c
      13'h11F5: dout  = 8'b00111000; // 4597 :  56 - 0x38
      13'h11F6: dout  = 8'b00010000; // 4598 :  16 - 0x10
      13'h11F7: dout  = 8'b00000000; // 4599 :   0 - 0x0
      13'h11F8: dout  = 8'b00000000; // 4600 :   0 - 0x0
      13'h11F9: dout  = 8'b00000000; // 4601 :   0 - 0x0
      13'h11FA: dout  = 8'b00000000; // 4602 :   0 - 0x0
      13'h11FB: dout  = 8'b00000000; // 4603 :   0 - 0x0
      13'h11FC: dout  = 8'b00000000; // 4604 :   0 - 0x0
      13'h11FD: dout  = 8'b00000000; // 4605 :   0 - 0x0
      13'h11FE: dout  = 8'b00000000; // 4606 :   0 - 0x0
      13'h11FF: dout  = 8'b00000000; // 4607 :   0 - 0x0
      13'h1200: dout  = 8'b11000110; // 4608 : 198 - 0xc6 -- Background 0x20
      13'h1201: dout  = 8'b11000110; // 4609 : 198 - 0xc6
      13'h1202: dout  = 8'b11010110; // 4610 : 214 - 0xd6
      13'h1203: dout  = 8'b11111110; // 4611 : 254 - 0xfe
      13'h1204: dout  = 8'b11111110; // 4612 : 254 - 0xfe
      13'h1205: dout  = 8'b11101110; // 4613 : 238 - 0xee
      13'h1206: dout  = 8'b11000110; // 4614 : 198 - 0xc6
      13'h1207: dout  = 8'b00000000; // 4615 :   0 - 0x0
      13'h1208: dout  = 8'b00000000; // 4616 :   0 - 0x0
      13'h1209: dout  = 8'b00000000; // 4617 :   0 - 0x0
      13'h120A: dout  = 8'b00000000; // 4618 :   0 - 0x0
      13'h120B: dout  = 8'b00000000; // 4619 :   0 - 0x0
      13'h120C: dout  = 8'b00000000; // 4620 :   0 - 0x0
      13'h120D: dout  = 8'b00000000; // 4621 :   0 - 0x0
      13'h120E: dout  = 8'b00000000; // 4622 :   0 - 0x0
      13'h120F: dout  = 8'b00000000; // 4623 :   0 - 0x0
      13'h1210: dout  = 8'b11000110; // 4624 : 198 - 0xc6 -- Background 0x21
      13'h1211: dout  = 8'b11101110; // 4625 : 238 - 0xee
      13'h1212: dout  = 8'b01111100; // 4626 : 124 - 0x7c
      13'h1213: dout  = 8'b00111000; // 4627 :  56 - 0x38
      13'h1214: dout  = 8'b01111100; // 4628 : 124 - 0x7c
      13'h1215: dout  = 8'b11101110; // 4629 : 238 - 0xee
      13'h1216: dout  = 8'b11000110; // 4630 : 198 - 0xc6
      13'h1217: dout  = 8'b00000000; // 4631 :   0 - 0x0
      13'h1218: dout  = 8'b00000000; // 4632 :   0 - 0x0
      13'h1219: dout  = 8'b00000000; // 4633 :   0 - 0x0
      13'h121A: dout  = 8'b00000000; // 4634 :   0 - 0x0
      13'h121B: dout  = 8'b00000000; // 4635 :   0 - 0x0
      13'h121C: dout  = 8'b00000000; // 4636 :   0 - 0x0
      13'h121D: dout  = 8'b00000000; // 4637 :   0 - 0x0
      13'h121E: dout  = 8'b00000000; // 4638 :   0 - 0x0
      13'h121F: dout  = 8'b00000000; // 4639 :   0 - 0x0
      13'h1220: dout  = 8'b01100110; // 4640 : 102 - 0x66 -- Background 0x22
      13'h1221: dout  = 8'b01100110; // 4641 : 102 - 0x66
      13'h1222: dout  = 8'b01100110; // 4642 : 102 - 0x66
      13'h1223: dout  = 8'b00111100; // 4643 :  60 - 0x3c
      13'h1224: dout  = 8'b00011000; // 4644 :  24 - 0x18
      13'h1225: dout  = 8'b00011000; // 4645 :  24 - 0x18
      13'h1226: dout  = 8'b00011000; // 4646 :  24 - 0x18
      13'h1227: dout  = 8'b00000000; // 4647 :   0 - 0x0
      13'h1228: dout  = 8'b00000000; // 4648 :   0 - 0x0
      13'h1229: dout  = 8'b00000000; // 4649 :   0 - 0x0
      13'h122A: dout  = 8'b00000000; // 4650 :   0 - 0x0
      13'h122B: dout  = 8'b00000000; // 4651 :   0 - 0x0
      13'h122C: dout  = 8'b00000000; // 4652 :   0 - 0x0
      13'h122D: dout  = 8'b00000000; // 4653 :   0 - 0x0
      13'h122E: dout  = 8'b00000000; // 4654 :   0 - 0x0
      13'h122F: dout  = 8'b00000000; // 4655 :   0 - 0x0
      13'h1230: dout  = 8'b11111110; // 4656 : 254 - 0xfe -- Background 0x23
      13'h1231: dout  = 8'b00001110; // 4657 :  14 - 0xe
      13'h1232: dout  = 8'b00011100; // 4658 :  28 - 0x1c
      13'h1233: dout  = 8'b00111000; // 4659 :  56 - 0x38
      13'h1234: dout  = 8'b01110000; // 4660 : 112 - 0x70
      13'h1235: dout  = 8'b11100000; // 4661 : 224 - 0xe0
      13'h1236: dout  = 8'b11111110; // 4662 : 254 - 0xfe
      13'h1237: dout  = 8'b00000000; // 4663 :   0 - 0x0
      13'h1238: dout  = 8'b00000000; // 4664 :   0 - 0x0
      13'h1239: dout  = 8'b00000000; // 4665 :   0 - 0x0
      13'h123A: dout  = 8'b00000000; // 4666 :   0 - 0x0
      13'h123B: dout  = 8'b00000000; // 4667 :   0 - 0x0
      13'h123C: dout  = 8'b00000000; // 4668 :   0 - 0x0
      13'h123D: dout  = 8'b00000000; // 4669 :   0 - 0x0
      13'h123E: dout  = 8'b00000000; // 4670 :   0 - 0x0
      13'h123F: dout  = 8'b00000000; // 4671 :   0 - 0x0
      13'h1240: dout  = 8'b00000000; // 4672 :   0 - 0x0 -- Background 0x24
      13'h1241: dout  = 8'b00000000; // 4673 :   0 - 0x0
      13'h1242: dout  = 8'b00000000; // 4674 :   0 - 0x0
      13'h1243: dout  = 8'b00000000; // 4675 :   0 - 0x0
      13'h1244: dout  = 8'b00000000; // 4676 :   0 - 0x0
      13'h1245: dout  = 8'b00000000; // 4677 :   0 - 0x0
      13'h1246: dout  = 8'b00000000; // 4678 :   0 - 0x0
      13'h1247: dout  = 8'b00000000; // 4679 :   0 - 0x0
      13'h1248: dout  = 8'b00000000; // 4680 :   0 - 0x0
      13'h1249: dout  = 8'b00000000; // 4681 :   0 - 0x0
      13'h124A: dout  = 8'b00000000; // 4682 :   0 - 0x0
      13'h124B: dout  = 8'b00000000; // 4683 :   0 - 0x0
      13'h124C: dout  = 8'b00000000; // 4684 :   0 - 0x0
      13'h124D: dout  = 8'b00000000; // 4685 :   0 - 0x0
      13'h124E: dout  = 8'b00000000; // 4686 :   0 - 0x0
      13'h124F: dout  = 8'b00000000; // 4687 :   0 - 0x0
      13'h1250: dout  = 8'b11111111; // 4688 : 255 - 0xff -- Background 0x25
      13'h1251: dout  = 8'b11111111; // 4689 : 255 - 0xff
      13'h1252: dout  = 8'b11111111; // 4690 : 255 - 0xff
      13'h1253: dout  = 8'b11111111; // 4691 : 255 - 0xff
      13'h1254: dout  = 8'b11111111; // 4692 : 255 - 0xff
      13'h1255: dout  = 8'b11111111; // 4693 : 255 - 0xff
      13'h1256: dout  = 8'b11111111; // 4694 : 255 - 0xff
      13'h1257: dout  = 8'b11111111; // 4695 : 255 - 0xff
      13'h1258: dout  = 8'b00000000; // 4696 :   0 - 0x0
      13'h1259: dout  = 8'b00000000; // 4697 :   0 - 0x0
      13'h125A: dout  = 8'b00000000; // 4698 :   0 - 0x0
      13'h125B: dout  = 8'b00000000; // 4699 :   0 - 0x0
      13'h125C: dout  = 8'b00000000; // 4700 :   0 - 0x0
      13'h125D: dout  = 8'b00000000; // 4701 :   0 - 0x0
      13'h125E: dout  = 8'b00000000; // 4702 :   0 - 0x0
      13'h125F: dout  = 8'b00000000; // 4703 :   0 - 0x0
      13'h1260: dout  = 8'b00000000; // 4704 :   0 - 0x0 -- Background 0x26
      13'h1261: dout  = 8'b00000000; // 4705 :   0 - 0x0
      13'h1262: dout  = 8'b00000000; // 4706 :   0 - 0x0
      13'h1263: dout  = 8'b00000000; // 4707 :   0 - 0x0
      13'h1264: dout  = 8'b00000000; // 4708 :   0 - 0x0
      13'h1265: dout  = 8'b00000000; // 4709 :   0 - 0x0
      13'h1266: dout  = 8'b00000000; // 4710 :   0 - 0x0
      13'h1267: dout  = 8'b00000000; // 4711 :   0 - 0x0
      13'h1268: dout  = 8'b11111111; // 4712 : 255 - 0xff
      13'h1269: dout  = 8'b11111111; // 4713 : 255 - 0xff
      13'h126A: dout  = 8'b11111111; // 4714 : 255 - 0xff
      13'h126B: dout  = 8'b11111111; // 4715 : 255 - 0xff
      13'h126C: dout  = 8'b11111111; // 4716 : 255 - 0xff
      13'h126D: dout  = 8'b11111111; // 4717 : 255 - 0xff
      13'h126E: dout  = 8'b11111111; // 4718 : 255 - 0xff
      13'h126F: dout  = 8'b11111111; // 4719 : 255 - 0xff
      13'h1270: dout  = 8'b11111111; // 4720 : 255 - 0xff -- Background 0x27
      13'h1271: dout  = 8'b11111111; // 4721 : 255 - 0xff
      13'h1272: dout  = 8'b11111111; // 4722 : 255 - 0xff
      13'h1273: dout  = 8'b11111111; // 4723 : 255 - 0xff
      13'h1274: dout  = 8'b11111111; // 4724 : 255 - 0xff
      13'h1275: dout  = 8'b11111111; // 4725 : 255 - 0xff
      13'h1276: dout  = 8'b11111111; // 4726 : 255 - 0xff
      13'h1277: dout  = 8'b11111111; // 4727 : 255 - 0xff
      13'h1278: dout  = 8'b11111111; // 4728 : 255 - 0xff
      13'h1279: dout  = 8'b11111111; // 4729 : 255 - 0xff
      13'h127A: dout  = 8'b11111111; // 4730 : 255 - 0xff
      13'h127B: dout  = 8'b11111111; // 4731 : 255 - 0xff
      13'h127C: dout  = 8'b11111111; // 4732 : 255 - 0xff
      13'h127D: dout  = 8'b11111111; // 4733 : 255 - 0xff
      13'h127E: dout  = 8'b11111111; // 4734 : 255 - 0xff
      13'h127F: dout  = 8'b11111111; // 4735 : 255 - 0xff
      13'h1280: dout  = 8'b00000000; // 4736 :   0 - 0x0 -- Background 0x28
      13'h1281: dout  = 8'b00000000; // 4737 :   0 - 0x0
      13'h1282: dout  = 8'b00000000; // 4738 :   0 - 0x0
      13'h1283: dout  = 8'b01111110; // 4739 : 126 - 0x7e
      13'h1284: dout  = 8'b01111110; // 4740 : 126 - 0x7e
      13'h1285: dout  = 8'b00000000; // 4741 :   0 - 0x0
      13'h1286: dout  = 8'b00000000; // 4742 :   0 - 0x0
      13'h1287: dout  = 8'b00000000; // 4743 :   0 - 0x0
      13'h1288: dout  = 8'b00000000; // 4744 :   0 - 0x0
      13'h1289: dout  = 8'b00000000; // 4745 :   0 - 0x0
      13'h128A: dout  = 8'b00000000; // 4746 :   0 - 0x0
      13'h128B: dout  = 8'b00000000; // 4747 :   0 - 0x0
      13'h128C: dout  = 8'b00000000; // 4748 :   0 - 0x0
      13'h128D: dout  = 8'b00000000; // 4749 :   0 - 0x0
      13'h128E: dout  = 8'b00000000; // 4750 :   0 - 0x0
      13'h128F: dout  = 8'b00000000; // 4751 :   0 - 0x0
      13'h1290: dout  = 8'b00000000; // 4752 :   0 - 0x0 -- Background 0x29
      13'h1291: dout  = 8'b00000000; // 4753 :   0 - 0x0
      13'h1292: dout  = 8'b01000100; // 4754 :  68 - 0x44
      13'h1293: dout  = 8'b00101000; // 4755 :  40 - 0x28
      13'h1294: dout  = 8'b00010000; // 4756 :  16 - 0x10
      13'h1295: dout  = 8'b00101000; // 4757 :  40 - 0x28
      13'h1296: dout  = 8'b01000100; // 4758 :  68 - 0x44
      13'h1297: dout  = 8'b00000000; // 4759 :   0 - 0x0
      13'h1298: dout  = 8'b00000000; // 4760 :   0 - 0x0
      13'h1299: dout  = 8'b00000000; // 4761 :   0 - 0x0
      13'h129A: dout  = 8'b00000000; // 4762 :   0 - 0x0
      13'h129B: dout  = 8'b00000000; // 4763 :   0 - 0x0
      13'h129C: dout  = 8'b00000000; // 4764 :   0 - 0x0
      13'h129D: dout  = 8'b00000000; // 4765 :   0 - 0x0
      13'h129E: dout  = 8'b00000000; // 4766 :   0 - 0x0
      13'h129F: dout  = 8'b00000000; // 4767 :   0 - 0x0
      13'h12A0: dout  = 8'b11111111; // 4768 : 255 - 0xff -- Background 0x2a
      13'h12A1: dout  = 8'b11111111; // 4769 : 255 - 0xff
      13'h12A2: dout  = 8'b11111111; // 4770 : 255 - 0xff
      13'h12A3: dout  = 8'b11111111; // 4771 : 255 - 0xff
      13'h12A4: dout  = 8'b11111111; // 4772 : 255 - 0xff
      13'h12A5: dout  = 8'b11111111; // 4773 : 255 - 0xff
      13'h12A6: dout  = 8'b11111111; // 4774 : 255 - 0xff
      13'h12A7: dout  = 8'b11111111; // 4775 : 255 - 0xff
      13'h12A8: dout  = 8'b01111111; // 4776 : 127 - 0x7f
      13'h12A9: dout  = 8'b01111111; // 4777 : 127 - 0x7f
      13'h12AA: dout  = 8'b01111111; // 4778 : 127 - 0x7f
      13'h12AB: dout  = 8'b01111111; // 4779 : 127 - 0x7f
      13'h12AC: dout  = 8'b01111111; // 4780 : 127 - 0x7f
      13'h12AD: dout  = 8'b01111111; // 4781 : 127 - 0x7f
      13'h12AE: dout  = 8'b01111111; // 4782 : 127 - 0x7f
      13'h12AF: dout  = 8'b01111111; // 4783 : 127 - 0x7f
      13'h12B0: dout  = 8'b00011000; // 4784 :  24 - 0x18 -- Background 0x2b
      13'h12B1: dout  = 8'b00111100; // 4785 :  60 - 0x3c
      13'h12B2: dout  = 8'b00111100; // 4786 :  60 - 0x3c
      13'h12B3: dout  = 8'b00111100; // 4787 :  60 - 0x3c
      13'h12B4: dout  = 8'b00011000; // 4788 :  24 - 0x18
      13'h12B5: dout  = 8'b00011000; // 4789 :  24 - 0x18
      13'h12B6: dout  = 8'b00000000; // 4790 :   0 - 0x0
      13'h12B7: dout  = 8'b00011000; // 4791 :  24 - 0x18
      13'h12B8: dout  = 8'b00000000; // 4792 :   0 - 0x0
      13'h12B9: dout  = 8'b00000000; // 4793 :   0 - 0x0
      13'h12BA: dout  = 8'b00000000; // 4794 :   0 - 0x0
      13'h12BB: dout  = 8'b00000000; // 4795 :   0 - 0x0
      13'h12BC: dout  = 8'b00000000; // 4796 :   0 - 0x0
      13'h12BD: dout  = 8'b00000000; // 4797 :   0 - 0x0
      13'h12BE: dout  = 8'b00000000; // 4798 :   0 - 0x0
      13'h12BF: dout  = 8'b00000000; // 4799 :   0 - 0x0
      13'h12C0: dout  = 8'b11111111; // 4800 : 255 - 0xff -- Background 0x2c
      13'h12C1: dout  = 8'b01111111; // 4801 : 127 - 0x7f
      13'h12C2: dout  = 8'b01111111; // 4802 : 127 - 0x7f
      13'h12C3: dout  = 8'b01111111; // 4803 : 127 - 0x7f
      13'h12C4: dout  = 8'b01111111; // 4804 : 127 - 0x7f
      13'h12C5: dout  = 8'b11111111; // 4805 : 255 - 0xff
      13'h12C6: dout  = 8'b11100011; // 4806 : 227 - 0xe3
      13'h12C7: dout  = 8'b11000001; // 4807 : 193 - 0xc1
      13'h12C8: dout  = 8'b11111111; // 4808 : 255 - 0xff
      13'h12C9: dout  = 8'b10000000; // 4809 : 128 - 0x80
      13'h12CA: dout  = 8'b10000000; // 4810 : 128 - 0x80
      13'h12CB: dout  = 8'b10000000; // 4811 : 128 - 0x80
      13'h12CC: dout  = 8'b10000000; // 4812 : 128 - 0x80
      13'h12CD: dout  = 8'b00000000; // 4813 :   0 - 0x0
      13'h12CE: dout  = 8'b00011100; // 4814 :  28 - 0x1c
      13'h12CF: dout  = 8'b00111110; // 4815 :  62 - 0x3e
      13'h12D0: dout  = 8'b10000000; // 4816 : 128 - 0x80 -- Background 0x2d
      13'h12D1: dout  = 8'b10000000; // 4817 : 128 - 0x80
      13'h12D2: dout  = 8'b10000000; // 4818 : 128 - 0x80
      13'h12D3: dout  = 8'b11000001; // 4819 : 193 - 0xc1
      13'h12D4: dout  = 8'b11100011; // 4820 : 227 - 0xe3
      13'h12D5: dout  = 8'b11111111; // 4821 : 255 - 0xff
      13'h12D6: dout  = 8'b11111111; // 4822 : 255 - 0xff
      13'h12D7: dout  = 8'b11111111; // 4823 : 255 - 0xff
      13'h12D8: dout  = 8'b01111111; // 4824 : 127 - 0x7f
      13'h12D9: dout  = 8'b01111111; // 4825 : 127 - 0x7f
      13'h12DA: dout  = 8'b01111111; // 4826 : 127 - 0x7f
      13'h12DB: dout  = 8'b00111110; // 4827 :  62 - 0x3e
      13'h12DC: dout  = 8'b00011100; // 4828 :  28 - 0x1c
      13'h12DD: dout  = 8'b00000000; // 4829 :   0 - 0x0
      13'h12DE: dout  = 8'b00000000; // 4830 :   0 - 0x0
      13'h12DF: dout  = 8'b11111111; // 4831 : 255 - 0xff
      13'h12E0: dout  = 8'b00111000; // 4832 :  56 - 0x38 -- Background 0x2e
      13'h12E1: dout  = 8'b01111100; // 4833 : 124 - 0x7c
      13'h12E2: dout  = 8'b01111100; // 4834 : 124 - 0x7c
      13'h12E3: dout  = 8'b01111100; // 4835 : 124 - 0x7c
      13'h12E4: dout  = 8'b01111100; // 4836 : 124 - 0x7c
      13'h12E5: dout  = 8'b01111100; // 4837 : 124 - 0x7c
      13'h12E6: dout  = 8'b00111000; // 4838 :  56 - 0x38
      13'h12E7: dout  = 8'b00000000; // 4839 :   0 - 0x0
      13'h12E8: dout  = 8'b00001000; // 4840 :   8 - 0x8
      13'h12E9: dout  = 8'b00000100; // 4841 :   4 - 0x4
      13'h12EA: dout  = 8'b00000100; // 4842 :   4 - 0x4
      13'h12EB: dout  = 8'b00000100; // 4843 :   4 - 0x4
      13'h12EC: dout  = 8'b00000100; // 4844 :   4 - 0x4
      13'h12ED: dout  = 8'b00000100; // 4845 :   4 - 0x4
      13'h12EE: dout  = 8'b00001000; // 4846 :   8 - 0x8
      13'h12EF: dout  = 8'b00000000; // 4847 :   0 - 0x0
      13'h12F0: dout  = 8'b00000011; // 4848 :   3 - 0x3 -- Background 0x2f
      13'h12F1: dout  = 8'b00000110; // 4849 :   6 - 0x6
      13'h12F2: dout  = 8'b00001100; // 4850 :  12 - 0xc
      13'h12F3: dout  = 8'b00001100; // 4851 :  12 - 0xc
      13'h12F4: dout  = 8'b00001000; // 4852 :   8 - 0x8
      13'h12F5: dout  = 8'b00001000; // 4853 :   8 - 0x8
      13'h12F6: dout  = 8'b00000100; // 4854 :   4 - 0x4
      13'h12F7: dout  = 8'b00000011; // 4855 :   3 - 0x3
      13'h12F8: dout  = 8'b00000011; // 4856 :   3 - 0x3
      13'h12F9: dout  = 8'b00000101; // 4857 :   5 - 0x5
      13'h12FA: dout  = 8'b00001011; // 4858 :  11 - 0xb
      13'h12FB: dout  = 8'b00001011; // 4859 :  11 - 0xb
      13'h12FC: dout  = 8'b00001111; // 4860 :  15 - 0xf
      13'h12FD: dout  = 8'b00001111; // 4861 :  15 - 0xf
      13'h12FE: dout  = 8'b00000111; // 4862 :   7 - 0x7
      13'h12FF: dout  = 8'b00000011; // 4863 :   3 - 0x3
      13'h1300: dout  = 8'b00000001; // 4864 :   1 - 0x1 -- Background 0x30
      13'h1301: dout  = 8'b00000010; // 4865 :   2 - 0x2
      13'h1302: dout  = 8'b00000100; // 4866 :   4 - 0x4
      13'h1303: dout  = 8'b00001000; // 4867 :   8 - 0x8
      13'h1304: dout  = 8'b00010000; // 4868 :  16 - 0x10
      13'h1305: dout  = 8'b00100000; // 4869 :  32 - 0x20
      13'h1306: dout  = 8'b01000000; // 4870 :  64 - 0x40
      13'h1307: dout  = 8'b10000000; // 4871 : 128 - 0x80
      13'h1308: dout  = 8'b00000001; // 4872 :   1 - 0x1
      13'h1309: dout  = 8'b00000011; // 4873 :   3 - 0x3
      13'h130A: dout  = 8'b00000111; // 4874 :   7 - 0x7
      13'h130B: dout  = 8'b00001111; // 4875 :  15 - 0xf
      13'h130C: dout  = 8'b00011111; // 4876 :  31 - 0x1f
      13'h130D: dout  = 8'b00111111; // 4877 :  63 - 0x3f
      13'h130E: dout  = 8'b01111111; // 4878 : 127 - 0x7f
      13'h130F: dout  = 8'b11111111; // 4879 : 255 - 0xff
      13'h1310: dout  = 8'b00000000; // 4880 :   0 - 0x0 -- Background 0x31
      13'h1311: dout  = 8'b00000000; // 4881 :   0 - 0x0
      13'h1312: dout  = 8'b00000000; // 4882 :   0 - 0x0
      13'h1313: dout  = 8'b00000000; // 4883 :   0 - 0x0
      13'h1314: dout  = 8'b00000000; // 4884 :   0 - 0x0
      13'h1315: dout  = 8'b00000111; // 4885 :   7 - 0x7
      13'h1316: dout  = 8'b00111000; // 4886 :  56 - 0x38
      13'h1317: dout  = 8'b11000000; // 4887 : 192 - 0xc0
      13'h1318: dout  = 8'b00000000; // 4888 :   0 - 0x0
      13'h1319: dout  = 8'b00000000; // 4889 :   0 - 0x0
      13'h131A: dout  = 8'b00000000; // 4890 :   0 - 0x0
      13'h131B: dout  = 8'b00000000; // 4891 :   0 - 0x0
      13'h131C: dout  = 8'b00000000; // 4892 :   0 - 0x0
      13'h131D: dout  = 8'b00000111; // 4893 :   7 - 0x7
      13'h131E: dout  = 8'b00111111; // 4894 :  63 - 0x3f
      13'h131F: dout  = 8'b11111111; // 4895 : 255 - 0xff
      13'h1320: dout  = 8'b00000000; // 4896 :   0 - 0x0 -- Background 0x32
      13'h1321: dout  = 8'b00000000; // 4897 :   0 - 0x0
      13'h1322: dout  = 8'b00000000; // 4898 :   0 - 0x0
      13'h1323: dout  = 8'b00000000; // 4899 :   0 - 0x0
      13'h1324: dout  = 8'b00000000; // 4900 :   0 - 0x0
      13'h1325: dout  = 8'b11100000; // 4901 : 224 - 0xe0
      13'h1326: dout  = 8'b00011100; // 4902 :  28 - 0x1c
      13'h1327: dout  = 8'b00000011; // 4903 :   3 - 0x3
      13'h1328: dout  = 8'b00000000; // 4904 :   0 - 0x0
      13'h1329: dout  = 8'b00000000; // 4905 :   0 - 0x0
      13'h132A: dout  = 8'b00000000; // 4906 :   0 - 0x0
      13'h132B: dout  = 8'b00000000; // 4907 :   0 - 0x0
      13'h132C: dout  = 8'b00000000; // 4908 :   0 - 0x0
      13'h132D: dout  = 8'b11100000; // 4909 : 224 - 0xe0
      13'h132E: dout  = 8'b11111100; // 4910 : 252 - 0xfc
      13'h132F: dout  = 8'b11111111; // 4911 : 255 - 0xff
      13'h1330: dout  = 8'b10000000; // 4912 : 128 - 0x80 -- Background 0x33
      13'h1331: dout  = 8'b01000000; // 4913 :  64 - 0x40
      13'h1332: dout  = 8'b00100000; // 4914 :  32 - 0x20
      13'h1333: dout  = 8'b00010000; // 4915 :  16 - 0x10
      13'h1334: dout  = 8'b00001000; // 4916 :   8 - 0x8
      13'h1335: dout  = 8'b00000100; // 4917 :   4 - 0x4
      13'h1336: dout  = 8'b00000010; // 4918 :   2 - 0x2
      13'h1337: dout  = 8'b00000001; // 4919 :   1 - 0x1
      13'h1338: dout  = 8'b10000000; // 4920 : 128 - 0x80
      13'h1339: dout  = 8'b11000000; // 4921 : 192 - 0xc0
      13'h133A: dout  = 8'b11100000; // 4922 : 224 - 0xe0
      13'h133B: dout  = 8'b11110000; // 4923 : 240 - 0xf0
      13'h133C: dout  = 8'b11111000; // 4924 : 248 - 0xf8
      13'h133D: dout  = 8'b11111100; // 4925 : 252 - 0xfc
      13'h133E: dout  = 8'b11111110; // 4926 : 254 - 0xfe
      13'h133F: dout  = 8'b11111111; // 4927 : 255 - 0xff
      13'h1340: dout  = 8'b00000100; // 4928 :   4 - 0x4 -- Background 0x34
      13'h1341: dout  = 8'b00001110; // 4929 :  14 - 0xe
      13'h1342: dout  = 8'b00001110; // 4930 :  14 - 0xe
      13'h1343: dout  = 8'b00001110; // 4931 :  14 - 0xe
      13'h1344: dout  = 8'b01101110; // 4932 : 110 - 0x6e
      13'h1345: dout  = 8'b01100100; // 4933 : 100 - 0x64
      13'h1346: dout  = 8'b01100000; // 4934 :  96 - 0x60
      13'h1347: dout  = 8'b01100000; // 4935 :  96 - 0x60
      13'h1348: dout  = 8'b11111111; // 4936 : 255 - 0xff
      13'h1349: dout  = 8'b11111111; // 4937 : 255 - 0xff
      13'h134A: dout  = 8'b11111111; // 4938 : 255 - 0xff
      13'h134B: dout  = 8'b11111111; // 4939 : 255 - 0xff
      13'h134C: dout  = 8'b11111111; // 4940 : 255 - 0xff
      13'h134D: dout  = 8'b11111111; // 4941 : 255 - 0xff
      13'h134E: dout  = 8'b11111111; // 4942 : 255 - 0xff
      13'h134F: dout  = 8'b11111111; // 4943 : 255 - 0xff
      13'h1350: dout  = 8'b00000111; // 4944 :   7 - 0x7 -- Background 0x35
      13'h1351: dout  = 8'b00001111; // 4945 :  15 - 0xf
      13'h1352: dout  = 8'b00011111; // 4946 :  31 - 0x1f
      13'h1353: dout  = 8'b00011111; // 4947 :  31 - 0x1f
      13'h1354: dout  = 8'b01111111; // 4948 : 127 - 0x7f
      13'h1355: dout  = 8'b11111111; // 4949 : 255 - 0xff
      13'h1356: dout  = 8'b11111111; // 4950 : 255 - 0xff
      13'h1357: dout  = 8'b01111111; // 4951 : 127 - 0x7f
      13'h1358: dout  = 8'b00000111; // 4952 :   7 - 0x7
      13'h1359: dout  = 8'b00001000; // 4953 :   8 - 0x8
      13'h135A: dout  = 8'b00010000; // 4954 :  16 - 0x10
      13'h135B: dout  = 8'b00000000; // 4955 :   0 - 0x0
      13'h135C: dout  = 8'b01100000; // 4956 :  96 - 0x60
      13'h135D: dout  = 8'b10000000; // 4957 : 128 - 0x80
      13'h135E: dout  = 8'b10000000; // 4958 : 128 - 0x80
      13'h135F: dout  = 8'b01000000; // 4959 :  64 - 0x40
      13'h1360: dout  = 8'b00000011; // 4960 :   3 - 0x3 -- Background 0x36
      13'h1361: dout  = 8'b00000111; // 4961 :   7 - 0x7
      13'h1362: dout  = 8'b00011111; // 4962 :  31 - 0x1f
      13'h1363: dout  = 8'b00111111; // 4963 :  63 - 0x3f
      13'h1364: dout  = 8'b00111111; // 4964 :  63 - 0x3f
      13'h1365: dout  = 8'b00111111; // 4965 :  63 - 0x3f
      13'h1366: dout  = 8'b01111001; // 4966 : 121 - 0x79
      13'h1367: dout  = 8'b11110111; // 4967 : 247 - 0xf7
      13'h1368: dout  = 8'b00000011; // 4968 :   3 - 0x3
      13'h1369: dout  = 8'b00000100; // 4969 :   4 - 0x4
      13'h136A: dout  = 8'b00011000; // 4970 :  24 - 0x18
      13'h136B: dout  = 8'b00100000; // 4971 :  32 - 0x20
      13'h136C: dout  = 8'b00100000; // 4972 :  32 - 0x20
      13'h136D: dout  = 8'b00100000; // 4973 :  32 - 0x20
      13'h136E: dout  = 8'b01000110; // 4974 :  70 - 0x46
      13'h136F: dout  = 8'b10001000; // 4975 : 136 - 0x88
      13'h1370: dout  = 8'b11000000; // 4976 : 192 - 0xc0 -- Background 0x37
      13'h1371: dout  = 8'b11100000; // 4977 : 224 - 0xe0
      13'h1372: dout  = 8'b11110000; // 4978 : 240 - 0xf0
      13'h1373: dout  = 8'b11110100; // 4979 : 244 - 0xf4
      13'h1374: dout  = 8'b11111110; // 4980 : 254 - 0xfe
      13'h1375: dout  = 8'b10111111; // 4981 : 191 - 0xbf
      13'h1376: dout  = 8'b11011111; // 4982 : 223 - 0xdf
      13'h1377: dout  = 8'b11111111; // 4983 : 255 - 0xff
      13'h1378: dout  = 8'b11000000; // 4984 : 192 - 0xc0
      13'h1379: dout  = 8'b00100000; // 4985 :  32 - 0x20
      13'h137A: dout  = 8'b00010000; // 4986 :  16 - 0x10
      13'h137B: dout  = 8'b00010100; // 4987 :  20 - 0x14
      13'h137C: dout  = 8'b00001010; // 4988 :  10 - 0xa
      13'h137D: dout  = 8'b01000001; // 4989 :  65 - 0x41
      13'h137E: dout  = 8'b00100001; // 4990 :  33 - 0x21
      13'h137F: dout  = 8'b00000001; // 4991 :   1 - 0x1
      13'h1380: dout  = 8'b10010000; // 4992 : 144 - 0x90 -- Background 0x38
      13'h1381: dout  = 8'b10111000; // 4993 : 184 - 0xb8
      13'h1382: dout  = 8'b11111000; // 4994 : 248 - 0xf8
      13'h1383: dout  = 8'b11111010; // 4995 : 250 - 0xfa
      13'h1384: dout  = 8'b11111111; // 4996 : 255 - 0xff
      13'h1385: dout  = 8'b11111111; // 4997 : 255 - 0xff
      13'h1386: dout  = 8'b11111111; // 4998 : 255 - 0xff
      13'h1387: dout  = 8'b11111110; // 4999 : 254 - 0xfe
      13'h1388: dout  = 8'b10010000; // 5000 : 144 - 0x90
      13'h1389: dout  = 8'b10101000; // 5001 : 168 - 0xa8
      13'h138A: dout  = 8'b01001000; // 5002 :  72 - 0x48
      13'h138B: dout  = 8'b00001010; // 5003 :  10 - 0xa
      13'h138C: dout  = 8'b00000101; // 5004 :   5 - 0x5
      13'h138D: dout  = 8'b00000001; // 5005 :   1 - 0x1
      13'h138E: dout  = 8'b00000001; // 5006 :   1 - 0x1
      13'h138F: dout  = 8'b00000010; // 5007 :   2 - 0x2
      13'h1390: dout  = 8'b00111011; // 5008 :  59 - 0x3b -- Background 0x39
      13'h1391: dout  = 8'b00011101; // 5009 :  29 - 0x1d
      13'h1392: dout  = 8'b00001110; // 5010 :  14 - 0xe
      13'h1393: dout  = 8'b00001111; // 5011 :  15 - 0xf
      13'h1394: dout  = 8'b00000111; // 5012 :   7 - 0x7
      13'h1395: dout  = 8'b00000000; // 5013 :   0 - 0x0
      13'h1396: dout  = 8'b00000000; // 5014 :   0 - 0x0
      13'h1397: dout  = 8'b00000000; // 5015 :   0 - 0x0
      13'h1398: dout  = 8'b00100100; // 5016 :  36 - 0x24
      13'h1399: dout  = 8'b00010010; // 5017 :  18 - 0x12
      13'h139A: dout  = 8'b00001001; // 5018 :   9 - 0x9
      13'h139B: dout  = 8'b00001000; // 5019 :   8 - 0x8
      13'h139C: dout  = 8'b00000111; // 5020 :   7 - 0x7
      13'h139D: dout  = 8'b00000000; // 5021 :   0 - 0x0
      13'h139E: dout  = 8'b00000000; // 5022 :   0 - 0x0
      13'h139F: dout  = 8'b00000000; // 5023 :   0 - 0x0
      13'h13A0: dout  = 8'b11111111; // 5024 : 255 - 0xff -- Background 0x3a
      13'h13A1: dout  = 8'b10111111; // 5025 : 191 - 0xbf
      13'h13A2: dout  = 8'b00011100; // 5026 :  28 - 0x1c
      13'h13A3: dout  = 8'b11000000; // 5027 : 192 - 0xc0
      13'h13A4: dout  = 8'b11110011; // 5028 : 243 - 0xf3
      13'h13A5: dout  = 8'b11111111; // 5029 : 255 - 0xff
      13'h13A6: dout  = 8'b01111110; // 5030 : 126 - 0x7e
      13'h13A7: dout  = 8'b00011100; // 5031 :  28 - 0x1c
      13'h13A8: dout  = 8'b00000000; // 5032 :   0 - 0x0
      13'h13A9: dout  = 8'b01000000; // 5033 :  64 - 0x40
      13'h13AA: dout  = 8'b11100011; // 5034 : 227 - 0xe3
      13'h13AB: dout  = 8'b00111111; // 5035 :  63 - 0x3f
      13'h13AC: dout  = 8'b00001100; // 5036 :  12 - 0xc
      13'h13AD: dout  = 8'b10000001; // 5037 : 129 - 0x81
      13'h13AE: dout  = 8'b01100010; // 5038 :  98 - 0x62
      13'h13AF: dout  = 8'b00011100; // 5039 :  28 - 0x1c
      13'h13B0: dout  = 8'b10111111; // 5040 : 191 - 0xbf -- Background 0x3b
      13'h13B1: dout  = 8'b01111111; // 5041 : 127 - 0x7f
      13'h13B2: dout  = 8'b00111101; // 5042 :  61 - 0x3d
      13'h13B3: dout  = 8'b10000011; // 5043 : 131 - 0x83
      13'h13B4: dout  = 8'b11000111; // 5044 : 199 - 0xc7
      13'h13B5: dout  = 8'b11111111; // 5045 : 255 - 0xff
      13'h13B6: dout  = 8'b11111111; // 5046 : 255 - 0xff
      13'h13B7: dout  = 8'b00111100; // 5047 :  60 - 0x3c
      13'h13B8: dout  = 8'b01000000; // 5048 :  64 - 0x40
      13'h13B9: dout  = 8'b10000000; // 5049 : 128 - 0x80
      13'h13BA: dout  = 8'b11000010; // 5050 : 194 - 0xc2
      13'h13BB: dout  = 8'b01111100; // 5051 : 124 - 0x7c
      13'h13BC: dout  = 8'b00111000; // 5052 :  56 - 0x38
      13'h13BD: dout  = 8'b00000000; // 5053 :   0 - 0x0
      13'h13BE: dout  = 8'b11000011; // 5054 : 195 - 0xc3
      13'h13BF: dout  = 8'b00111100; // 5055 :  60 - 0x3c
      13'h13C0: dout  = 8'b11111100; // 5056 : 252 - 0xfc -- Background 0x3c
      13'h13C1: dout  = 8'b11111110; // 5057 : 254 - 0xfe
      13'h13C2: dout  = 8'b11111111; // 5058 : 255 - 0xff
      13'h13C3: dout  = 8'b11111110; // 5059 : 254 - 0xfe
      13'h13C4: dout  = 8'b11111110; // 5060 : 254 - 0xfe
      13'h13C5: dout  = 8'b11111000; // 5061 : 248 - 0xf8
      13'h13C6: dout  = 8'b01100000; // 5062 :  96 - 0x60
      13'h13C7: dout  = 8'b00000000; // 5063 :   0 - 0x0
      13'h13C8: dout  = 8'b00000100; // 5064 :   4 - 0x4
      13'h13C9: dout  = 8'b00000010; // 5065 :   2 - 0x2
      13'h13CA: dout  = 8'b00000001; // 5066 :   1 - 0x1
      13'h13CB: dout  = 8'b00000000; // 5067 :   0 - 0x0
      13'h13CC: dout  = 8'b00000110; // 5068 :   6 - 0x6
      13'h13CD: dout  = 8'b10011000; // 5069 : 152 - 0x98
      13'h13CE: dout  = 8'b01100000; // 5070 :  96 - 0x60
      13'h13CF: dout  = 8'b00000000; // 5071 :   0 - 0x0
      13'h13D0: dout  = 8'b11000000; // 5072 : 192 - 0xc0 -- Background 0x3d
      13'h13D1: dout  = 8'b00100000; // 5073 :  32 - 0x20
      13'h13D2: dout  = 8'b00010000; // 5074 :  16 - 0x10
      13'h13D3: dout  = 8'b00010000; // 5075 :  16 - 0x10
      13'h13D4: dout  = 8'b00010000; // 5076 :  16 - 0x10
      13'h13D5: dout  = 8'b00010000; // 5077 :  16 - 0x10
      13'h13D6: dout  = 8'b00100000; // 5078 :  32 - 0x20
      13'h13D7: dout  = 8'b11000000; // 5079 : 192 - 0xc0
      13'h13D8: dout  = 8'b11000000; // 5080 : 192 - 0xc0
      13'h13D9: dout  = 8'b11100000; // 5081 : 224 - 0xe0
      13'h13DA: dout  = 8'b11110000; // 5082 : 240 - 0xf0
      13'h13DB: dout  = 8'b11110000; // 5083 : 240 - 0xf0
      13'h13DC: dout  = 8'b11110000; // 5084 : 240 - 0xf0
      13'h13DD: dout  = 8'b11110000; // 5085 : 240 - 0xf0
      13'h13DE: dout  = 8'b11100000; // 5086 : 224 - 0xe0
      13'h13DF: dout  = 8'b11000000; // 5087 : 192 - 0xc0
      13'h13E0: dout  = 8'b00000000; // 5088 :   0 - 0x0 -- Background 0x3e
      13'h13E1: dout  = 8'b00000000; // 5089 :   0 - 0x0
      13'h13E2: dout  = 8'b00000000; // 5090 :   0 - 0x0
      13'h13E3: dout  = 8'b00000000; // 5091 :   0 - 0x0
      13'h13E4: dout  = 8'b00111111; // 5092 :  63 - 0x3f
      13'h13E5: dout  = 8'b01111111; // 5093 : 127 - 0x7f
      13'h13E6: dout  = 8'b11100000; // 5094 : 224 - 0xe0
      13'h13E7: dout  = 8'b11000000; // 5095 : 192 - 0xc0
      13'h13E8: dout  = 8'b00000000; // 5096 :   0 - 0x0
      13'h13E9: dout  = 8'b00000000; // 5097 :   0 - 0x0
      13'h13EA: dout  = 8'b00000000; // 5098 :   0 - 0x0
      13'h13EB: dout  = 8'b00000000; // 5099 :   0 - 0x0
      13'h13EC: dout  = 8'b00000000; // 5100 :   0 - 0x0
      13'h13ED: dout  = 8'b00000000; // 5101 :   0 - 0x0
      13'h13EE: dout  = 8'b00011100; // 5102 :  28 - 0x1c
      13'h13EF: dout  = 8'b00111110; // 5103 :  62 - 0x3e
      13'h13F0: dout  = 8'b10001000; // 5104 : 136 - 0x88 -- Background 0x3f
      13'h13F1: dout  = 8'b10011100; // 5105 : 156 - 0x9c
      13'h13F2: dout  = 8'b10001000; // 5106 : 136 - 0x88
      13'h13F3: dout  = 8'b10000000; // 5107 : 128 - 0x80
      13'h13F4: dout  = 8'b10000000; // 5108 : 128 - 0x80
      13'h13F5: dout  = 8'b10000000; // 5109 : 128 - 0x80
      13'h13F6: dout  = 8'b10000000; // 5110 : 128 - 0x80
      13'h13F7: dout  = 8'b10000000; // 5111 : 128 - 0x80
      13'h13F8: dout  = 8'b01111111; // 5112 : 127 - 0x7f
      13'h13F9: dout  = 8'b01111111; // 5113 : 127 - 0x7f
      13'h13FA: dout  = 8'b01111111; // 5114 : 127 - 0x7f
      13'h13FB: dout  = 8'b00111110; // 5115 :  62 - 0x3e
      13'h13FC: dout  = 8'b00011100; // 5116 :  28 - 0x1c
      13'h13FD: dout  = 8'b00000000; // 5117 :   0 - 0x0
      13'h13FE: dout  = 8'b00000000; // 5118 :   0 - 0x0
      13'h13FF: dout  = 8'b00000000; // 5119 :   0 - 0x0
      13'h1400: dout  = 8'b11111110; // 5120 : 254 - 0xfe -- Background 0x40
      13'h1401: dout  = 8'b11111110; // 5121 : 254 - 0xfe
      13'h1402: dout  = 8'b11111110; // 5122 : 254 - 0xfe
      13'h1403: dout  = 8'b11111110; // 5123 : 254 - 0xfe
      13'h1404: dout  = 8'b11111110; // 5124 : 254 - 0xfe
      13'h1405: dout  = 8'b11111110; // 5125 : 254 - 0xfe
      13'h1406: dout  = 8'b11111110; // 5126 : 254 - 0xfe
      13'h1407: dout  = 8'b11111110; // 5127 : 254 - 0xfe
      13'h1408: dout  = 8'b11111111; // 5128 : 255 - 0xff
      13'h1409: dout  = 8'b11111111; // 5129 : 255 - 0xff
      13'h140A: dout  = 8'b11111111; // 5130 : 255 - 0xff
      13'h140B: dout  = 8'b11111111; // 5131 : 255 - 0xff
      13'h140C: dout  = 8'b11111111; // 5132 : 255 - 0xff
      13'h140D: dout  = 8'b11111111; // 5133 : 255 - 0xff
      13'h140E: dout  = 8'b11111111; // 5134 : 255 - 0xff
      13'h140F: dout  = 8'b11111111; // 5135 : 255 - 0xff
      13'h1410: dout  = 8'b00001000; // 5136 :   8 - 0x8 -- Background 0x41
      13'h1411: dout  = 8'b00010100; // 5137 :  20 - 0x14
      13'h1412: dout  = 8'b00100100; // 5138 :  36 - 0x24
      13'h1413: dout  = 8'b11000100; // 5139 : 196 - 0xc4
      13'h1414: dout  = 8'b00000011; // 5140 :   3 - 0x3
      13'h1415: dout  = 8'b01000000; // 5141 :  64 - 0x40
      13'h1416: dout  = 8'b10100001; // 5142 : 161 - 0xa1
      13'h1417: dout  = 8'b00100110; // 5143 :  38 - 0x26
      13'h1418: dout  = 8'b00000000; // 5144 :   0 - 0x0
      13'h1419: dout  = 8'b00001000; // 5145 :   8 - 0x8
      13'h141A: dout  = 8'b00011000; // 5146 :  24 - 0x18
      13'h141B: dout  = 8'b00111000; // 5147 :  56 - 0x38
      13'h141C: dout  = 8'b11111100; // 5148 : 252 - 0xfc
      13'h141D: dout  = 8'b10111111; // 5149 : 191 - 0xbf
      13'h141E: dout  = 8'b01011110; // 5150 :  94 - 0x5e
      13'h141F: dout  = 8'b11011001; // 5151 : 217 - 0xd9
      13'h1420: dout  = 8'b11111111; // 5152 : 255 - 0xff -- Background 0x42
      13'h1421: dout  = 8'b11111111; // 5153 : 255 - 0xff
      13'h1422: dout  = 8'b11111111; // 5154 : 255 - 0xff
      13'h1423: dout  = 8'b11111111; // 5155 : 255 - 0xff
      13'h1424: dout  = 8'b01111111; // 5156 : 127 - 0x7f
      13'h1425: dout  = 8'b01111111; // 5157 : 127 - 0x7f
      13'h1426: dout  = 8'b01111111; // 5158 : 127 - 0x7f
      13'h1427: dout  = 8'b01111111; // 5159 : 127 - 0x7f
      13'h1428: dout  = 8'b10000001; // 5160 : 129 - 0x81
      13'h1429: dout  = 8'b10000001; // 5161 : 129 - 0x81
      13'h142A: dout  = 8'b10000001; // 5162 : 129 - 0x81
      13'h142B: dout  = 8'b10000001; // 5163 : 129 - 0x81
      13'h142C: dout  = 8'b10000001; // 5164 : 129 - 0x81
      13'h142D: dout  = 8'b10000001; // 5165 : 129 - 0x81
      13'h142E: dout  = 8'b10000001; // 5166 : 129 - 0x81
      13'h142F: dout  = 8'b10000001; // 5167 : 129 - 0x81
      13'h1430: dout  = 8'b11111111; // 5168 : 255 - 0xff -- Background 0x43
      13'h1431: dout  = 8'b11111111; // 5169 : 255 - 0xff
      13'h1432: dout  = 8'b11111111; // 5170 : 255 - 0xff
      13'h1433: dout  = 8'b11111111; // 5171 : 255 - 0xff
      13'h1434: dout  = 8'b11111111; // 5172 : 255 - 0xff
      13'h1435: dout  = 8'b11111111; // 5173 : 255 - 0xff
      13'h1436: dout  = 8'b11111111; // 5174 : 255 - 0xff
      13'h1437: dout  = 8'b11111111; // 5175 : 255 - 0xff
      13'h1438: dout  = 8'b00000001; // 5176 :   1 - 0x1
      13'h1439: dout  = 8'b00000001; // 5177 :   1 - 0x1
      13'h143A: dout  = 8'b00000001; // 5178 :   1 - 0x1
      13'h143B: dout  = 8'b00000001; // 5179 :   1 - 0x1
      13'h143C: dout  = 8'b00000001; // 5180 :   1 - 0x1
      13'h143D: dout  = 8'b00000001; // 5181 :   1 - 0x1
      13'h143E: dout  = 8'b00000001; // 5182 :   1 - 0x1
      13'h143F: dout  = 8'b00000001; // 5183 :   1 - 0x1
      13'h1440: dout  = 8'b01111111; // 5184 : 127 - 0x7f -- Background 0x44
      13'h1441: dout  = 8'b10000000; // 5185 : 128 - 0x80
      13'h1442: dout  = 8'b10000000; // 5186 : 128 - 0x80
      13'h1443: dout  = 8'b10011000; // 5187 : 152 - 0x98
      13'h1444: dout  = 8'b10011100; // 5188 : 156 - 0x9c
      13'h1445: dout  = 8'b10001100; // 5189 : 140 - 0x8c
      13'h1446: dout  = 8'b10000000; // 5190 : 128 - 0x80
      13'h1447: dout  = 8'b10000000; // 5191 : 128 - 0x80
      13'h1448: dout  = 8'b00000000; // 5192 :   0 - 0x0
      13'h1449: dout  = 8'b01111111; // 5193 : 127 - 0x7f
      13'h144A: dout  = 8'b01111111; // 5194 : 127 - 0x7f
      13'h144B: dout  = 8'b01100111; // 5195 : 103 - 0x67
      13'h144C: dout  = 8'b01100111; // 5196 : 103 - 0x67
      13'h144D: dout  = 8'b01111111; // 5197 : 127 - 0x7f
      13'h144E: dout  = 8'b01111111; // 5198 : 127 - 0x7f
      13'h144F: dout  = 8'b01111111; // 5199 : 127 - 0x7f
      13'h1450: dout  = 8'b11111111; // 5200 : 255 - 0xff -- Background 0x45
      13'h1451: dout  = 8'b00000001; // 5201 :   1 - 0x1
      13'h1452: dout  = 8'b00000001; // 5202 :   1 - 0x1
      13'h1453: dout  = 8'b11111111; // 5203 : 255 - 0xff
      13'h1454: dout  = 8'b00010000; // 5204 :  16 - 0x10
      13'h1455: dout  = 8'b00010000; // 5205 :  16 - 0x10
      13'h1456: dout  = 8'b00010000; // 5206 :  16 - 0x10
      13'h1457: dout  = 8'b11111111; // 5207 : 255 - 0xff
      13'h1458: dout  = 8'b00000000; // 5208 :   0 - 0x0
      13'h1459: dout  = 8'b11111111; // 5209 : 255 - 0xff
      13'h145A: dout  = 8'b11111111; // 5210 : 255 - 0xff
      13'h145B: dout  = 8'b11111111; // 5211 : 255 - 0xff
      13'h145C: dout  = 8'b11111111; // 5212 : 255 - 0xff
      13'h145D: dout  = 8'b11111111; // 5213 : 255 - 0xff
      13'h145E: dout  = 8'b11111111; // 5214 : 255 - 0xff
      13'h145F: dout  = 8'b11111111; // 5215 : 255 - 0xff
      13'h1460: dout  = 8'b10000000; // 5216 : 128 - 0x80 -- Background 0x46
      13'h1461: dout  = 8'b10000000; // 5217 : 128 - 0x80
      13'h1462: dout  = 8'b10000000; // 5218 : 128 - 0x80
      13'h1463: dout  = 8'b10000000; // 5219 : 128 - 0x80
      13'h1464: dout  = 8'b10000000; // 5220 : 128 - 0x80
      13'h1465: dout  = 8'b10000000; // 5221 : 128 - 0x80
      13'h1466: dout  = 8'b10000000; // 5222 : 128 - 0x80
      13'h1467: dout  = 8'b10000000; // 5223 : 128 - 0x80
      13'h1468: dout  = 8'b01111111; // 5224 : 127 - 0x7f
      13'h1469: dout  = 8'b01111111; // 5225 : 127 - 0x7f
      13'h146A: dout  = 8'b01111111; // 5226 : 127 - 0x7f
      13'h146B: dout  = 8'b01111111; // 5227 : 127 - 0x7f
      13'h146C: dout  = 8'b01111111; // 5228 : 127 - 0x7f
      13'h146D: dout  = 8'b01111111; // 5229 : 127 - 0x7f
      13'h146E: dout  = 8'b01111111; // 5230 : 127 - 0x7f
      13'h146F: dout  = 8'b01111111; // 5231 : 127 - 0x7f
      13'h1470: dout  = 8'b00000001; // 5232 :   1 - 0x1 -- Background 0x47
      13'h1471: dout  = 8'b00000001; // 5233 :   1 - 0x1
      13'h1472: dout  = 8'b00000001; // 5234 :   1 - 0x1
      13'h1473: dout  = 8'b11111111; // 5235 : 255 - 0xff
      13'h1474: dout  = 8'b00010000; // 5236 :  16 - 0x10
      13'h1475: dout  = 8'b00010000; // 5237 :  16 - 0x10
      13'h1476: dout  = 8'b00010000; // 5238 :  16 - 0x10
      13'h1477: dout  = 8'b11111111; // 5239 : 255 - 0xff
      13'h1478: dout  = 8'b11111111; // 5240 : 255 - 0xff
      13'h1479: dout  = 8'b11111111; // 5241 : 255 - 0xff
      13'h147A: dout  = 8'b11111111; // 5242 : 255 - 0xff
      13'h147B: dout  = 8'b11111111; // 5243 : 255 - 0xff
      13'h147C: dout  = 8'b11111111; // 5244 : 255 - 0xff
      13'h147D: dout  = 8'b11111111; // 5245 : 255 - 0xff
      13'h147E: dout  = 8'b11111111; // 5246 : 255 - 0xff
      13'h147F: dout  = 8'b11111111; // 5247 : 255 - 0xff
      13'h1480: dout  = 8'b11111111; // 5248 : 255 - 0xff -- Background 0x48
      13'h1481: dout  = 8'b00000000; // 5249 :   0 - 0x0
      13'h1482: dout  = 8'b00000000; // 5250 :   0 - 0x0
      13'h1483: dout  = 8'b00000000; // 5251 :   0 - 0x0
      13'h1484: dout  = 8'b00000000; // 5252 :   0 - 0x0
      13'h1485: dout  = 8'b00000000; // 5253 :   0 - 0x0
      13'h1486: dout  = 8'b00000000; // 5254 :   0 - 0x0
      13'h1487: dout  = 8'b00000000; // 5255 :   0 - 0x0
      13'h1488: dout  = 8'b00000000; // 5256 :   0 - 0x0
      13'h1489: dout  = 8'b11111111; // 5257 : 255 - 0xff
      13'h148A: dout  = 8'b11111111; // 5258 : 255 - 0xff
      13'h148B: dout  = 8'b11111111; // 5259 : 255 - 0xff
      13'h148C: dout  = 8'b11111111; // 5260 : 255 - 0xff
      13'h148D: dout  = 8'b11111111; // 5261 : 255 - 0xff
      13'h148E: dout  = 8'b11111111; // 5262 : 255 - 0xff
      13'h148F: dout  = 8'b11111111; // 5263 : 255 - 0xff
      13'h1490: dout  = 8'b11111110; // 5264 : 254 - 0xfe -- Background 0x49
      13'h1491: dout  = 8'b00000001; // 5265 :   1 - 0x1
      13'h1492: dout  = 8'b00000001; // 5266 :   1 - 0x1
      13'h1493: dout  = 8'b00011001; // 5267 :  25 - 0x19
      13'h1494: dout  = 8'b00011101; // 5268 :  29 - 0x1d
      13'h1495: dout  = 8'b00001101; // 5269 :  13 - 0xd
      13'h1496: dout  = 8'b00000001; // 5270 :   1 - 0x1
      13'h1497: dout  = 8'b00000001; // 5271 :   1 - 0x1
      13'h1498: dout  = 8'b00000000; // 5272 :   0 - 0x0
      13'h1499: dout  = 8'b11111111; // 5273 : 255 - 0xff
      13'h149A: dout  = 8'b11111111; // 5274 : 255 - 0xff
      13'h149B: dout  = 8'b11100111; // 5275 : 231 - 0xe7
      13'h149C: dout  = 8'b11100111; // 5276 : 231 - 0xe7
      13'h149D: dout  = 8'b11111111; // 5277 : 255 - 0xff
      13'h149E: dout  = 8'b11111111; // 5278 : 255 - 0xff
      13'h149F: dout  = 8'b11111111; // 5279 : 255 - 0xff
      13'h14A0: dout  = 8'b00000001; // 5280 :   1 - 0x1 -- Background 0x4a
      13'h14A1: dout  = 8'b00000001; // 5281 :   1 - 0x1
      13'h14A2: dout  = 8'b00000001; // 5282 :   1 - 0x1
      13'h14A3: dout  = 8'b00000001; // 5283 :   1 - 0x1
      13'h14A4: dout  = 8'b00000001; // 5284 :   1 - 0x1
      13'h14A5: dout  = 8'b00000001; // 5285 :   1 - 0x1
      13'h14A6: dout  = 8'b00000001; // 5286 :   1 - 0x1
      13'h14A7: dout  = 8'b00000001; // 5287 :   1 - 0x1
      13'h14A8: dout  = 8'b11111111; // 5288 : 255 - 0xff
      13'h14A9: dout  = 8'b11111111; // 5289 : 255 - 0xff
      13'h14AA: dout  = 8'b11111111; // 5290 : 255 - 0xff
      13'h14AB: dout  = 8'b11111111; // 5291 : 255 - 0xff
      13'h14AC: dout  = 8'b11111111; // 5292 : 255 - 0xff
      13'h14AD: dout  = 8'b11111111; // 5293 : 255 - 0xff
      13'h14AE: dout  = 8'b11111111; // 5294 : 255 - 0xff
      13'h14AF: dout  = 8'b11111111; // 5295 : 255 - 0xff
      13'h14B0: dout  = 8'b00111111; // 5296 :  63 - 0x3f -- Background 0x4b
      13'h14B1: dout  = 8'b01111111; // 5297 : 127 - 0x7f
      13'h14B2: dout  = 8'b01111111; // 5298 : 127 - 0x7f
      13'h14B3: dout  = 8'b11111111; // 5299 : 255 - 0xff
      13'h14B4: dout  = 8'b11111111; // 5300 : 255 - 0xff
      13'h14B5: dout  = 8'b11111111; // 5301 : 255 - 0xff
      13'h14B6: dout  = 8'b11111111; // 5302 : 255 - 0xff
      13'h14B7: dout  = 8'b11111111; // 5303 : 255 - 0xff
      13'h14B8: dout  = 8'b00111111; // 5304 :  63 - 0x3f
      13'h14B9: dout  = 8'b01100000; // 5305 :  96 - 0x60
      13'h14BA: dout  = 8'b01000000; // 5306 :  64 - 0x40
      13'h14BB: dout  = 8'b11000000; // 5307 : 192 - 0xc0
      13'h14BC: dout  = 8'b10000000; // 5308 : 128 - 0x80
      13'h14BD: dout  = 8'b10000000; // 5309 : 128 - 0x80
      13'h14BE: dout  = 8'b10000000; // 5310 : 128 - 0x80
      13'h14BF: dout  = 8'b10000000; // 5311 : 128 - 0x80
      13'h14C0: dout  = 8'b11111111; // 5312 : 255 - 0xff -- Background 0x4c
      13'h14C1: dout  = 8'b11111111; // 5313 : 255 - 0xff
      13'h14C2: dout  = 8'b11111111; // 5314 : 255 - 0xff
      13'h14C3: dout  = 8'b11111111; // 5315 : 255 - 0xff
      13'h14C4: dout  = 8'b11111111; // 5316 : 255 - 0xff
      13'h14C5: dout  = 8'b11111111; // 5317 : 255 - 0xff
      13'h14C6: dout  = 8'b01111110; // 5318 : 126 - 0x7e
      13'h14C7: dout  = 8'b00111100; // 5319 :  60 - 0x3c
      13'h14C8: dout  = 8'b10000000; // 5320 : 128 - 0x80
      13'h14C9: dout  = 8'b10000000; // 5321 : 128 - 0x80
      13'h14CA: dout  = 8'b10000000; // 5322 : 128 - 0x80
      13'h14CB: dout  = 8'b10000000; // 5323 : 128 - 0x80
      13'h14CC: dout  = 8'b10000000; // 5324 : 128 - 0x80
      13'h14CD: dout  = 8'b10000001; // 5325 : 129 - 0x81
      13'h14CE: dout  = 8'b01000010; // 5326 :  66 - 0x42
      13'h14CF: dout  = 8'b00111100; // 5327 :  60 - 0x3c
      13'h14D0: dout  = 8'b11111111; // 5328 : 255 - 0xff -- Background 0x4d
      13'h14D1: dout  = 8'b11111111; // 5329 : 255 - 0xff
      13'h14D2: dout  = 8'b11111111; // 5330 : 255 - 0xff
      13'h14D3: dout  = 8'b11111111; // 5331 : 255 - 0xff
      13'h14D4: dout  = 8'b11111111; // 5332 : 255 - 0xff
      13'h14D5: dout  = 8'b11111111; // 5333 : 255 - 0xff
      13'h14D6: dout  = 8'b11111111; // 5334 : 255 - 0xff
      13'h14D7: dout  = 8'b11111111; // 5335 : 255 - 0xff
      13'h14D8: dout  = 8'b11111111; // 5336 : 255 - 0xff
      13'h14D9: dout  = 8'b00000000; // 5337 :   0 - 0x0
      13'h14DA: dout  = 8'b00000000; // 5338 :   0 - 0x0
      13'h14DB: dout  = 8'b00000000; // 5339 :   0 - 0x0
      13'h14DC: dout  = 8'b00000000; // 5340 :   0 - 0x0
      13'h14DD: dout  = 8'b00000000; // 5341 :   0 - 0x0
      13'h14DE: dout  = 8'b00000000; // 5342 :   0 - 0x0
      13'h14DF: dout  = 8'b00000000; // 5343 :   0 - 0x0
      13'h14E0: dout  = 8'b11111111; // 5344 : 255 - 0xff -- Background 0x4e
      13'h14E1: dout  = 8'b11111111; // 5345 : 255 - 0xff
      13'h14E2: dout  = 8'b11111111; // 5346 : 255 - 0xff
      13'h14E3: dout  = 8'b11111111; // 5347 : 255 - 0xff
      13'h14E4: dout  = 8'b11111111; // 5348 : 255 - 0xff
      13'h14E5: dout  = 8'b11111111; // 5349 : 255 - 0xff
      13'h14E6: dout  = 8'b11111110; // 5350 : 254 - 0xfe
      13'h14E7: dout  = 8'b01111100; // 5351 : 124 - 0x7c
      13'h14E8: dout  = 8'b00000000; // 5352 :   0 - 0x0
      13'h14E9: dout  = 8'b00000000; // 5353 :   0 - 0x0
      13'h14EA: dout  = 8'b00000000; // 5354 :   0 - 0x0
      13'h14EB: dout  = 8'b00000000; // 5355 :   0 - 0x0
      13'h14EC: dout  = 8'b00000000; // 5356 :   0 - 0x0
      13'h14ED: dout  = 8'b00000001; // 5357 :   1 - 0x1
      13'h14EE: dout  = 8'b10000010; // 5358 : 130 - 0x82
      13'h14EF: dout  = 8'b01111100; // 5359 : 124 - 0x7c
      13'h14F0: dout  = 8'b11111111; // 5360 : 255 - 0xff -- Background 0x4f
      13'h14F1: dout  = 8'b11111111; // 5361 : 255 - 0xff
      13'h14F2: dout  = 8'b11111111; // 5362 : 255 - 0xff
      13'h14F3: dout  = 8'b11111111; // 5363 : 255 - 0xff
      13'h14F4: dout  = 8'b11111111; // 5364 : 255 - 0xff
      13'h14F5: dout  = 8'b11111111; // 5365 : 255 - 0xff
      13'h14F6: dout  = 8'b11111110; // 5366 : 254 - 0xfe
      13'h14F7: dout  = 8'b01111100; // 5367 : 124 - 0x7c
      13'h14F8: dout  = 8'b00000000; // 5368 :   0 - 0x0
      13'h14F9: dout  = 8'b00000000; // 5369 :   0 - 0x0
      13'h14FA: dout  = 8'b00000000; // 5370 :   0 - 0x0
      13'h14FB: dout  = 8'b00000000; // 5371 :   0 - 0x0
      13'h14FC: dout  = 8'b00000000; // 5372 :   0 - 0x0
      13'h14FD: dout  = 8'b00000001; // 5373 :   1 - 0x1
      13'h14FE: dout  = 8'b10000011; // 5374 : 131 - 0x83
      13'h14FF: dout  = 8'b11111111; // 5375 : 255 - 0xff
      13'h1500: dout  = 8'b11111000; // 5376 : 248 - 0xf8 -- Background 0x50
      13'h1501: dout  = 8'b11111100; // 5377 : 252 - 0xfc
      13'h1502: dout  = 8'b11111110; // 5378 : 254 - 0xfe
      13'h1503: dout  = 8'b11111110; // 5379 : 254 - 0xfe
      13'h1504: dout  = 8'b11111111; // 5380 : 255 - 0xff
      13'h1505: dout  = 8'b11111111; // 5381 : 255 - 0xff
      13'h1506: dout  = 8'b11111111; // 5382 : 255 - 0xff
      13'h1507: dout  = 8'b11111111; // 5383 : 255 - 0xff
      13'h1508: dout  = 8'b11111000; // 5384 : 248 - 0xf8
      13'h1509: dout  = 8'b00000100; // 5385 :   4 - 0x4
      13'h150A: dout  = 8'b00000010; // 5386 :   2 - 0x2
      13'h150B: dout  = 8'b00000010; // 5387 :   2 - 0x2
      13'h150C: dout  = 8'b00000001; // 5388 :   1 - 0x1
      13'h150D: dout  = 8'b00000001; // 5389 :   1 - 0x1
      13'h150E: dout  = 8'b00000001; // 5390 :   1 - 0x1
      13'h150F: dout  = 8'b00000001; // 5391 :   1 - 0x1
      13'h1510: dout  = 8'b11111111; // 5392 : 255 - 0xff -- Background 0x51
      13'h1511: dout  = 8'b11111111; // 5393 : 255 - 0xff
      13'h1512: dout  = 8'b11111111; // 5394 : 255 - 0xff
      13'h1513: dout  = 8'b11111111; // 5395 : 255 - 0xff
      13'h1514: dout  = 8'b11111111; // 5396 : 255 - 0xff
      13'h1515: dout  = 8'b11111111; // 5397 : 255 - 0xff
      13'h1516: dout  = 8'b01111110; // 5398 : 126 - 0x7e
      13'h1517: dout  = 8'b00111100; // 5399 :  60 - 0x3c
      13'h1518: dout  = 8'b00000001; // 5400 :   1 - 0x1
      13'h1519: dout  = 8'b00000001; // 5401 :   1 - 0x1
      13'h151A: dout  = 8'b00000001; // 5402 :   1 - 0x1
      13'h151B: dout  = 8'b00000001; // 5403 :   1 - 0x1
      13'h151C: dout  = 8'b00000001; // 5404 :   1 - 0x1
      13'h151D: dout  = 8'b10000001; // 5405 : 129 - 0x81
      13'h151E: dout  = 8'b01000010; // 5406 :  66 - 0x42
      13'h151F: dout  = 8'b00111100; // 5407 :  60 - 0x3c
      13'h1520: dout  = 8'b00000000; // 5408 :   0 - 0x0 -- Background 0x52
      13'h1521: dout  = 8'b00001000; // 5409 :   8 - 0x8
      13'h1522: dout  = 8'b00001000; // 5410 :   8 - 0x8
      13'h1523: dout  = 8'b00001000; // 5411 :   8 - 0x8
      13'h1524: dout  = 8'b00010000; // 5412 :  16 - 0x10
      13'h1525: dout  = 8'b00010000; // 5413 :  16 - 0x10
      13'h1526: dout  = 8'b00010000; // 5414 :  16 - 0x10
      13'h1527: dout  = 8'b00000000; // 5415 :   0 - 0x0
      13'h1528: dout  = 8'b11111111; // 5416 : 255 - 0xff
      13'h1529: dout  = 8'b11111111; // 5417 : 255 - 0xff
      13'h152A: dout  = 8'b11111111; // 5418 : 255 - 0xff
      13'h152B: dout  = 8'b11111111; // 5419 : 255 - 0xff
      13'h152C: dout  = 8'b11111111; // 5420 : 255 - 0xff
      13'h152D: dout  = 8'b11111111; // 5421 : 255 - 0xff
      13'h152E: dout  = 8'b11111111; // 5422 : 255 - 0xff
      13'h152F: dout  = 8'b11111111; // 5423 : 255 - 0xff
      13'h1530: dout  = 8'b00000000; // 5424 :   0 - 0x0 -- Background 0x53
      13'h1531: dout  = 8'b01111111; // 5425 : 127 - 0x7f
      13'h1532: dout  = 8'b01111111; // 5426 : 127 - 0x7f
      13'h1533: dout  = 8'b01111000; // 5427 : 120 - 0x78
      13'h1534: dout  = 8'b01110011; // 5428 : 115 - 0x73
      13'h1535: dout  = 8'b01110011; // 5429 : 115 - 0x73
      13'h1536: dout  = 8'b01110011; // 5430 : 115 - 0x73
      13'h1537: dout  = 8'b01111111; // 5431 : 127 - 0x7f
      13'h1538: dout  = 8'b01111111; // 5432 : 127 - 0x7f
      13'h1539: dout  = 8'b10000000; // 5433 : 128 - 0x80
      13'h153A: dout  = 8'b10100000; // 5434 : 160 - 0xa0
      13'h153B: dout  = 8'b10000111; // 5435 : 135 - 0x87
      13'h153C: dout  = 8'b10001111; // 5436 : 143 - 0x8f
      13'h153D: dout  = 8'b10001110; // 5437 : 142 - 0x8e
      13'h153E: dout  = 8'b10001110; // 5438 : 142 - 0x8e
      13'h153F: dout  = 8'b10000110; // 5439 : 134 - 0x86
      13'h1540: dout  = 8'b00000000; // 5440 :   0 - 0x0 -- Background 0x54
      13'h1541: dout  = 8'b11111111; // 5441 : 255 - 0xff
      13'h1542: dout  = 8'b11111111; // 5442 : 255 - 0xff
      13'h1543: dout  = 8'b00111111; // 5443 :  63 - 0x3f
      13'h1544: dout  = 8'b10011111; // 5444 : 159 - 0x9f
      13'h1545: dout  = 8'b10011111; // 5445 : 159 - 0x9f
      13'h1546: dout  = 8'b10011111; // 5446 : 159 - 0x9f
      13'h1547: dout  = 8'b00011111; // 5447 :  31 - 0x1f
      13'h1548: dout  = 8'b11111110; // 5448 : 254 - 0xfe
      13'h1549: dout  = 8'b00000001; // 5449 :   1 - 0x1
      13'h154A: dout  = 8'b00000101; // 5450 :   5 - 0x5
      13'h154B: dout  = 8'b11000001; // 5451 : 193 - 0xc1
      13'h154C: dout  = 8'b11100001; // 5452 : 225 - 0xe1
      13'h154D: dout  = 8'b01110001; // 5453 : 113 - 0x71
      13'h154E: dout  = 8'b01110001; // 5454 : 113 - 0x71
      13'h154F: dout  = 8'b11110001; // 5455 : 241 - 0xf1
      13'h1550: dout  = 8'b01111110; // 5456 : 126 - 0x7e -- Background 0x55
      13'h1551: dout  = 8'b01111110; // 5457 : 126 - 0x7e
      13'h1552: dout  = 8'b01111111; // 5458 : 127 - 0x7f
      13'h1553: dout  = 8'b01111110; // 5459 : 126 - 0x7e
      13'h1554: dout  = 8'b01111110; // 5460 : 126 - 0x7e
      13'h1555: dout  = 8'b01111111; // 5461 : 127 - 0x7f
      13'h1556: dout  = 8'b01111111; // 5462 : 127 - 0x7f
      13'h1557: dout  = 8'b11111111; // 5463 : 255 - 0xff
      13'h1558: dout  = 8'b10000001; // 5464 : 129 - 0x81
      13'h1559: dout  = 8'b10000001; // 5465 : 129 - 0x81
      13'h155A: dout  = 8'b10000000; // 5466 : 128 - 0x80
      13'h155B: dout  = 8'b10000001; // 5467 : 129 - 0x81
      13'h155C: dout  = 8'b10000001; // 5468 : 129 - 0x81
      13'h155D: dout  = 8'b10100000; // 5469 : 160 - 0xa0
      13'h155E: dout  = 8'b10000000; // 5470 : 128 - 0x80
      13'h155F: dout  = 8'b11111111; // 5471 : 255 - 0xff
      13'h1560: dout  = 8'b01111111; // 5472 : 127 - 0x7f -- Background 0x56
      13'h1561: dout  = 8'b01111111; // 5473 : 127 - 0x7f
      13'h1562: dout  = 8'b11111111; // 5474 : 255 - 0xff
      13'h1563: dout  = 8'b01111111; // 5475 : 127 - 0x7f
      13'h1564: dout  = 8'b01111111; // 5476 : 127 - 0x7f
      13'h1565: dout  = 8'b11111111; // 5477 : 255 - 0xff
      13'h1566: dout  = 8'b11111111; // 5478 : 255 - 0xff
      13'h1567: dout  = 8'b11111111; // 5479 : 255 - 0xff
      13'h1568: dout  = 8'b11110001; // 5480 : 241 - 0xf1
      13'h1569: dout  = 8'b11000001; // 5481 : 193 - 0xc1
      13'h156A: dout  = 8'b11000001; // 5482 : 193 - 0xc1
      13'h156B: dout  = 8'b10000001; // 5483 : 129 - 0x81
      13'h156C: dout  = 8'b11000001; // 5484 : 193 - 0xc1
      13'h156D: dout  = 8'b11000101; // 5485 : 197 - 0xc5
      13'h156E: dout  = 8'b00000001; // 5486 :   1 - 0x1
      13'h156F: dout  = 8'b11111111; // 5487 : 255 - 0xff
      13'h1570: dout  = 8'b01111111; // 5488 : 127 - 0x7f -- Background 0x57
      13'h1571: dout  = 8'b10000000; // 5489 : 128 - 0x80
      13'h1572: dout  = 8'b10100000; // 5490 : 160 - 0xa0
      13'h1573: dout  = 8'b10000000; // 5491 : 128 - 0x80
      13'h1574: dout  = 8'b10000000; // 5492 : 128 - 0x80
      13'h1575: dout  = 8'b10000000; // 5493 : 128 - 0x80
      13'h1576: dout  = 8'b10000000; // 5494 : 128 - 0x80
      13'h1577: dout  = 8'b10000000; // 5495 : 128 - 0x80
      13'h1578: dout  = 8'b01111111; // 5496 : 127 - 0x7f
      13'h1579: dout  = 8'b11111111; // 5497 : 255 - 0xff
      13'h157A: dout  = 8'b11111111; // 5498 : 255 - 0xff
      13'h157B: dout  = 8'b11111111; // 5499 : 255 - 0xff
      13'h157C: dout  = 8'b11111111; // 5500 : 255 - 0xff
      13'h157D: dout  = 8'b11111111; // 5501 : 255 - 0xff
      13'h157E: dout  = 8'b11111111; // 5502 : 255 - 0xff
      13'h157F: dout  = 8'b11111111; // 5503 : 255 - 0xff
      13'h1580: dout  = 8'b11111110; // 5504 : 254 - 0xfe -- Background 0x58
      13'h1581: dout  = 8'b00000001; // 5505 :   1 - 0x1
      13'h1582: dout  = 8'b00000101; // 5506 :   5 - 0x5
      13'h1583: dout  = 8'b00000001; // 5507 :   1 - 0x1
      13'h1584: dout  = 8'b00000001; // 5508 :   1 - 0x1
      13'h1585: dout  = 8'b00000001; // 5509 :   1 - 0x1
      13'h1586: dout  = 8'b00000001; // 5510 :   1 - 0x1
      13'h1587: dout  = 8'b00000001; // 5511 :   1 - 0x1
      13'h1588: dout  = 8'b11111110; // 5512 : 254 - 0xfe
      13'h1589: dout  = 8'b11111111; // 5513 : 255 - 0xff
      13'h158A: dout  = 8'b11111111; // 5514 : 255 - 0xff
      13'h158B: dout  = 8'b11111111; // 5515 : 255 - 0xff
      13'h158C: dout  = 8'b11111111; // 5516 : 255 - 0xff
      13'h158D: dout  = 8'b11111111; // 5517 : 255 - 0xff
      13'h158E: dout  = 8'b11111111; // 5518 : 255 - 0xff
      13'h158F: dout  = 8'b11111111; // 5519 : 255 - 0xff
      13'h1590: dout  = 8'b10000000; // 5520 : 128 - 0x80 -- Background 0x59
      13'h1591: dout  = 8'b10000000; // 5521 : 128 - 0x80
      13'h1592: dout  = 8'b10000000; // 5522 : 128 - 0x80
      13'h1593: dout  = 8'b10000000; // 5523 : 128 - 0x80
      13'h1594: dout  = 8'b10000000; // 5524 : 128 - 0x80
      13'h1595: dout  = 8'b10100000; // 5525 : 160 - 0xa0
      13'h1596: dout  = 8'b10000000; // 5526 : 128 - 0x80
      13'h1597: dout  = 8'b01111111; // 5527 : 127 - 0x7f
      13'h1598: dout  = 8'b11111111; // 5528 : 255 - 0xff
      13'h1599: dout  = 8'b11111111; // 5529 : 255 - 0xff
      13'h159A: dout  = 8'b11111111; // 5530 : 255 - 0xff
      13'h159B: dout  = 8'b11111111; // 5531 : 255 - 0xff
      13'h159C: dout  = 8'b11111111; // 5532 : 255 - 0xff
      13'h159D: dout  = 8'b11111111; // 5533 : 255 - 0xff
      13'h159E: dout  = 8'b11111111; // 5534 : 255 - 0xff
      13'h159F: dout  = 8'b01111111; // 5535 : 127 - 0x7f
      13'h15A0: dout  = 8'b00000001; // 5536 :   1 - 0x1 -- Background 0x5a
      13'h15A1: dout  = 8'b00000001; // 5537 :   1 - 0x1
      13'h15A2: dout  = 8'b00000001; // 5538 :   1 - 0x1
      13'h15A3: dout  = 8'b00000001; // 5539 :   1 - 0x1
      13'h15A4: dout  = 8'b00000001; // 5540 :   1 - 0x1
      13'h15A5: dout  = 8'b00000101; // 5541 :   5 - 0x5
      13'h15A6: dout  = 8'b00000001; // 5542 :   1 - 0x1
      13'h15A7: dout  = 8'b11111110; // 5543 : 254 - 0xfe
      13'h15A8: dout  = 8'b11111111; // 5544 : 255 - 0xff
      13'h15A9: dout  = 8'b11111111; // 5545 : 255 - 0xff
      13'h15AA: dout  = 8'b11111111; // 5546 : 255 - 0xff
      13'h15AB: dout  = 8'b11111111; // 5547 : 255 - 0xff
      13'h15AC: dout  = 8'b11111111; // 5548 : 255 - 0xff
      13'h15AD: dout  = 8'b11111111; // 5549 : 255 - 0xff
      13'h15AE: dout  = 8'b11111111; // 5550 : 255 - 0xff
      13'h15AF: dout  = 8'b11111110; // 5551 : 254 - 0xfe
      13'h15B0: dout  = 8'b00000000; // 5552 :   0 - 0x0 -- Background 0x5b
      13'h15B1: dout  = 8'b00000000; // 5553 :   0 - 0x0
      13'h15B2: dout  = 8'b00000000; // 5554 :   0 - 0x0
      13'h15B3: dout  = 8'b00000000; // 5555 :   0 - 0x0
      13'h15B4: dout  = 8'b11111100; // 5556 : 252 - 0xfc
      13'h15B5: dout  = 8'b11111110; // 5557 : 254 - 0xfe
      13'h15B6: dout  = 8'b00000111; // 5558 :   7 - 0x7
      13'h15B7: dout  = 8'b00000011; // 5559 :   3 - 0x3
      13'h15B8: dout  = 8'b00000000; // 5560 :   0 - 0x0
      13'h15B9: dout  = 8'b00000000; // 5561 :   0 - 0x0
      13'h15BA: dout  = 8'b00000000; // 5562 :   0 - 0x0
      13'h15BB: dout  = 8'b00000000; // 5563 :   0 - 0x0
      13'h15BC: dout  = 8'b00000000; // 5564 :   0 - 0x0
      13'h15BD: dout  = 8'b00000000; // 5565 :   0 - 0x0
      13'h15BE: dout  = 8'b00111000; // 5566 :  56 - 0x38
      13'h15BF: dout  = 8'b01111100; // 5567 : 124 - 0x7c
      13'h15C0: dout  = 8'b00010001; // 5568 :  17 - 0x11 -- Background 0x5c
      13'h15C1: dout  = 8'b00111001; // 5569 :  57 - 0x39
      13'h15C2: dout  = 8'b00010001; // 5570 :  17 - 0x11
      13'h15C3: dout  = 8'b00000001; // 5571 :   1 - 0x1
      13'h15C4: dout  = 8'b00000001; // 5572 :   1 - 0x1
      13'h15C5: dout  = 8'b00000001; // 5573 :   1 - 0x1
      13'h15C6: dout  = 8'b00000001; // 5574 :   1 - 0x1
      13'h15C7: dout  = 8'b00000001; // 5575 :   1 - 0x1
      13'h15C8: dout  = 8'b11111110; // 5576 : 254 - 0xfe
      13'h15C9: dout  = 8'b11111110; // 5577 : 254 - 0xfe
      13'h15CA: dout  = 8'b11111110; // 5578 : 254 - 0xfe
      13'h15CB: dout  = 8'b01111100; // 5579 : 124 - 0x7c
      13'h15CC: dout  = 8'b00111000; // 5580 :  56 - 0x38
      13'h15CD: dout  = 8'b00000000; // 5581 :   0 - 0x0
      13'h15CE: dout  = 8'b00000000; // 5582 :   0 - 0x0
      13'h15CF: dout  = 8'b00000000; // 5583 :   0 - 0x0
      13'h15D0: dout  = 8'b11101111; // 5584 : 239 - 0xef -- Background 0x5d
      13'h15D1: dout  = 8'b00101000; // 5585 :  40 - 0x28
      13'h15D2: dout  = 8'b00101000; // 5586 :  40 - 0x28
      13'h15D3: dout  = 8'b00101000; // 5587 :  40 - 0x28
      13'h15D4: dout  = 8'b00101000; // 5588 :  40 - 0x28
      13'h15D5: dout  = 8'b00101000; // 5589 :  40 - 0x28
      13'h15D6: dout  = 8'b11101111; // 5590 : 239 - 0xef
      13'h15D7: dout  = 8'b00000000; // 5591 :   0 - 0x0
      13'h15D8: dout  = 8'b00100000; // 5592 :  32 - 0x20
      13'h15D9: dout  = 8'b11100111; // 5593 : 231 - 0xe7
      13'h15DA: dout  = 8'b11100111; // 5594 : 231 - 0xe7
      13'h15DB: dout  = 8'b11100111; // 5595 : 231 - 0xe7
      13'h15DC: dout  = 8'b11100111; // 5596 : 231 - 0xe7
      13'h15DD: dout  = 8'b11100111; // 5597 : 231 - 0xe7
      13'h15DE: dout  = 8'b11101111; // 5598 : 239 - 0xef
      13'h15DF: dout  = 8'b00000000; // 5599 :   0 - 0x0
      13'h15E0: dout  = 8'b11111110; // 5600 : 254 - 0xfe -- Background 0x5e
      13'h15E1: dout  = 8'b10000010; // 5601 : 130 - 0x82
      13'h15E2: dout  = 8'b10000010; // 5602 : 130 - 0x82
      13'h15E3: dout  = 8'b10000010; // 5603 : 130 - 0x82
      13'h15E4: dout  = 8'b10000010; // 5604 : 130 - 0x82
      13'h15E5: dout  = 8'b10000010; // 5605 : 130 - 0x82
      13'h15E6: dout  = 8'b11111110; // 5606 : 254 - 0xfe
      13'h15E7: dout  = 8'b00000000; // 5607 :   0 - 0x0
      13'h15E8: dout  = 8'b00000010; // 5608 :   2 - 0x2
      13'h15E9: dout  = 8'b01111110; // 5609 : 126 - 0x7e
      13'h15EA: dout  = 8'b01111110; // 5610 : 126 - 0x7e
      13'h15EB: dout  = 8'b01111110; // 5611 : 126 - 0x7e
      13'h15EC: dout  = 8'b01111110; // 5612 : 126 - 0x7e
      13'h15ED: dout  = 8'b01111110; // 5613 : 126 - 0x7e
      13'h15EE: dout  = 8'b11111110; // 5614 : 254 - 0xfe
      13'h15EF: dout  = 8'b00000000; // 5615 :   0 - 0x0
      13'h15F0: dout  = 8'b10000000; // 5616 : 128 - 0x80 -- Background 0x5f
      13'h15F1: dout  = 8'b10000000; // 5617 : 128 - 0x80
      13'h15F2: dout  = 8'b10000000; // 5618 : 128 - 0x80
      13'h15F3: dout  = 8'b10011000; // 5619 : 152 - 0x98
      13'h15F4: dout  = 8'b10011100; // 5620 : 156 - 0x9c
      13'h15F5: dout  = 8'b10001100; // 5621 : 140 - 0x8c
      13'h15F6: dout  = 8'b10000000; // 5622 : 128 - 0x80
      13'h15F7: dout  = 8'b01111111; // 5623 : 127 - 0x7f
      13'h15F8: dout  = 8'b01111111; // 5624 : 127 - 0x7f
      13'h15F9: dout  = 8'b01111111; // 5625 : 127 - 0x7f
      13'h15FA: dout  = 8'b01111111; // 5626 : 127 - 0x7f
      13'h15FB: dout  = 8'b01100111; // 5627 : 103 - 0x67
      13'h15FC: dout  = 8'b01100111; // 5628 : 103 - 0x67
      13'h15FD: dout  = 8'b01111111; // 5629 : 127 - 0x7f
      13'h15FE: dout  = 8'b01111111; // 5630 : 127 - 0x7f
      13'h15FF: dout  = 8'b01111111; // 5631 : 127 - 0x7f
      13'h1600: dout  = 8'b11111111; // 5632 : 255 - 0xff -- Background 0x60
      13'h1601: dout  = 8'b11111111; // 5633 : 255 - 0xff
      13'h1602: dout  = 8'b10000011; // 5634 : 131 - 0x83
      13'h1603: dout  = 8'b11110011; // 5635 : 243 - 0xf3
      13'h1604: dout  = 8'b11110011; // 5636 : 243 - 0xf3
      13'h1605: dout  = 8'b11110011; // 5637 : 243 - 0xf3
      13'h1606: dout  = 8'b11110011; // 5638 : 243 - 0xf3
      13'h1607: dout  = 8'b11110011; // 5639 : 243 - 0xf3
      13'h1608: dout  = 8'b11111111; // 5640 : 255 - 0xff
      13'h1609: dout  = 8'b10000000; // 5641 : 128 - 0x80
      13'h160A: dout  = 8'b11111100; // 5642 : 252 - 0xfc
      13'h160B: dout  = 8'b10001100; // 5643 : 140 - 0x8c
      13'h160C: dout  = 8'b10001100; // 5644 : 140 - 0x8c
      13'h160D: dout  = 8'b10001100; // 5645 : 140 - 0x8c
      13'h160E: dout  = 8'b10001100; // 5646 : 140 - 0x8c
      13'h160F: dout  = 8'b10001100; // 5647 : 140 - 0x8c
      13'h1610: dout  = 8'b11111111; // 5648 : 255 - 0xff -- Background 0x61
      13'h1611: dout  = 8'b11111111; // 5649 : 255 - 0xff
      13'h1612: dout  = 8'b11110000; // 5650 : 240 - 0xf0
      13'h1613: dout  = 8'b11110110; // 5651 : 246 - 0xf6
      13'h1614: dout  = 8'b11110110; // 5652 : 246 - 0xf6
      13'h1615: dout  = 8'b11110110; // 5653 : 246 - 0xf6
      13'h1616: dout  = 8'b11110110; // 5654 : 246 - 0xf6
      13'h1617: dout  = 8'b11110110; // 5655 : 246 - 0xf6
      13'h1618: dout  = 8'b11111111; // 5656 : 255 - 0xff
      13'h1619: dout  = 8'b00000000; // 5657 :   0 - 0x0
      13'h161A: dout  = 8'b00001111; // 5658 :  15 - 0xf
      13'h161B: dout  = 8'b00001001; // 5659 :   9 - 0x9
      13'h161C: dout  = 8'b00001001; // 5660 :   9 - 0x9
      13'h161D: dout  = 8'b00001001; // 5661 :   9 - 0x9
      13'h161E: dout  = 8'b00001001; // 5662 :   9 - 0x9
      13'h161F: dout  = 8'b00001001; // 5663 :   9 - 0x9
      13'h1620: dout  = 8'b11111111; // 5664 : 255 - 0xff -- Background 0x62
      13'h1621: dout  = 8'b11111111; // 5665 : 255 - 0xff
      13'h1622: dout  = 8'b00000000; // 5666 :   0 - 0x0
      13'h1623: dout  = 8'b00000000; // 5667 :   0 - 0x0
      13'h1624: dout  = 8'b00000000; // 5668 :   0 - 0x0
      13'h1625: dout  = 8'b00000000; // 5669 :   0 - 0x0
      13'h1626: dout  = 8'b00000000; // 5670 :   0 - 0x0
      13'h1627: dout  = 8'b00000000; // 5671 :   0 - 0x0
      13'h1628: dout  = 8'b11111111; // 5672 : 255 - 0xff
      13'h1629: dout  = 8'b00000000; // 5673 :   0 - 0x0
      13'h162A: dout  = 8'b11111111; // 5674 : 255 - 0xff
      13'h162B: dout  = 8'b11111111; // 5675 : 255 - 0xff
      13'h162C: dout  = 8'b11111111; // 5676 : 255 - 0xff
      13'h162D: dout  = 8'b11111111; // 5677 : 255 - 0xff
      13'h162E: dout  = 8'b11111111; // 5678 : 255 - 0xff
      13'h162F: dout  = 8'b11111111; // 5679 : 255 - 0xff
      13'h1630: dout  = 8'b11111111; // 5680 : 255 - 0xff -- Background 0x63
      13'h1631: dout  = 8'b11111111; // 5681 : 255 - 0xff
      13'h1632: dout  = 8'b00000001; // 5682 :   1 - 0x1
      13'h1633: dout  = 8'b01010111; // 5683 :  87 - 0x57
      13'h1634: dout  = 8'b00101111; // 5684 :  47 - 0x2f
      13'h1635: dout  = 8'b01010111; // 5685 :  87 - 0x57
      13'h1636: dout  = 8'b00101111; // 5686 :  47 - 0x2f
      13'h1637: dout  = 8'b01010111; // 5687 :  87 - 0x57
      13'h1638: dout  = 8'b11111111; // 5688 : 255 - 0xff
      13'h1639: dout  = 8'b00000001; // 5689 :   1 - 0x1
      13'h163A: dout  = 8'b11111111; // 5690 : 255 - 0xff
      13'h163B: dout  = 8'b10101001; // 5691 : 169 - 0xa9
      13'h163C: dout  = 8'b11010001; // 5692 : 209 - 0xd1
      13'h163D: dout  = 8'b10101001; // 5693 : 169 - 0xa9
      13'h163E: dout  = 8'b11010001; // 5694 : 209 - 0xd1
      13'h163F: dout  = 8'b10101001; // 5695 : 169 - 0xa9
      13'h1640: dout  = 8'b11110011; // 5696 : 243 - 0xf3 -- Background 0x64
      13'h1641: dout  = 8'b11110011; // 5697 : 243 - 0xf3
      13'h1642: dout  = 8'b11110011; // 5698 : 243 - 0xf3
      13'h1643: dout  = 8'b11110011; // 5699 : 243 - 0xf3
      13'h1644: dout  = 8'b11110011; // 5700 : 243 - 0xf3
      13'h1645: dout  = 8'b11110011; // 5701 : 243 - 0xf3
      13'h1646: dout  = 8'b11111111; // 5702 : 255 - 0xff
      13'h1647: dout  = 8'b00111111; // 5703 :  63 - 0x3f
      13'h1648: dout  = 8'b10001100; // 5704 : 140 - 0x8c
      13'h1649: dout  = 8'b10001100; // 5705 : 140 - 0x8c
      13'h164A: dout  = 8'b10001100; // 5706 : 140 - 0x8c
      13'h164B: dout  = 8'b10001100; // 5707 : 140 - 0x8c
      13'h164C: dout  = 8'b10001100; // 5708 : 140 - 0x8c
      13'h164D: dout  = 8'b10001100; // 5709 : 140 - 0x8c
      13'h164E: dout  = 8'b11111111; // 5710 : 255 - 0xff
      13'h164F: dout  = 8'b00111111; // 5711 :  63 - 0x3f
      13'h1650: dout  = 8'b11110110; // 5712 : 246 - 0xf6 -- Background 0x65
      13'h1651: dout  = 8'b11110110; // 5713 : 246 - 0xf6
      13'h1652: dout  = 8'b11110110; // 5714 : 246 - 0xf6
      13'h1653: dout  = 8'b11110110; // 5715 : 246 - 0xf6
      13'h1654: dout  = 8'b11110110; // 5716 : 246 - 0xf6
      13'h1655: dout  = 8'b11110110; // 5717 : 246 - 0xf6
      13'h1656: dout  = 8'b11111111; // 5718 : 255 - 0xff
      13'h1657: dout  = 8'b11111111; // 5719 : 255 - 0xff
      13'h1658: dout  = 8'b00001001; // 5720 :   9 - 0x9
      13'h1659: dout  = 8'b00001001; // 5721 :   9 - 0x9
      13'h165A: dout  = 8'b00001001; // 5722 :   9 - 0x9
      13'h165B: dout  = 8'b00001001; // 5723 :   9 - 0x9
      13'h165C: dout  = 8'b00001001; // 5724 :   9 - 0x9
      13'h165D: dout  = 8'b00001001; // 5725 :   9 - 0x9
      13'h165E: dout  = 8'b11111111; // 5726 : 255 - 0xff
      13'h165F: dout  = 8'b11111111; // 5727 : 255 - 0xff
      13'h1660: dout  = 8'b00000000; // 5728 :   0 - 0x0 -- Background 0x66
      13'h1661: dout  = 8'b00000000; // 5729 :   0 - 0x0
      13'h1662: dout  = 8'b00000000; // 5730 :   0 - 0x0
      13'h1663: dout  = 8'b00000000; // 5731 :   0 - 0x0
      13'h1664: dout  = 8'b00000000; // 5732 :   0 - 0x0
      13'h1665: dout  = 8'b00000000; // 5733 :   0 - 0x0
      13'h1666: dout  = 8'b11111111; // 5734 : 255 - 0xff
      13'h1667: dout  = 8'b11111111; // 5735 : 255 - 0xff
      13'h1668: dout  = 8'b11111111; // 5736 : 255 - 0xff
      13'h1669: dout  = 8'b11111111; // 5737 : 255 - 0xff
      13'h166A: dout  = 8'b11111111; // 5738 : 255 - 0xff
      13'h166B: dout  = 8'b11111111; // 5739 : 255 - 0xff
      13'h166C: dout  = 8'b11111111; // 5740 : 255 - 0xff
      13'h166D: dout  = 8'b11111111; // 5741 : 255 - 0xff
      13'h166E: dout  = 8'b11111111; // 5742 : 255 - 0xff
      13'h166F: dout  = 8'b11111111; // 5743 : 255 - 0xff
      13'h1670: dout  = 8'b00101111; // 5744 :  47 - 0x2f -- Background 0x67
      13'h1671: dout  = 8'b01010111; // 5745 :  87 - 0x57
      13'h1672: dout  = 8'b00101111; // 5746 :  47 - 0x2f
      13'h1673: dout  = 8'b01010111; // 5747 :  87 - 0x57
      13'h1674: dout  = 8'b00101111; // 5748 :  47 - 0x2f
      13'h1675: dout  = 8'b01010111; // 5749 :  87 - 0x57
      13'h1676: dout  = 8'b11111111; // 5750 : 255 - 0xff
      13'h1677: dout  = 8'b11111100; // 5751 : 252 - 0xfc
      13'h1678: dout  = 8'b11010001; // 5752 : 209 - 0xd1
      13'h1679: dout  = 8'b10101001; // 5753 : 169 - 0xa9
      13'h167A: dout  = 8'b11010001; // 5754 : 209 - 0xd1
      13'h167B: dout  = 8'b10101001; // 5755 : 169 - 0xa9
      13'h167C: dout  = 8'b11010001; // 5756 : 209 - 0xd1
      13'h167D: dout  = 8'b10101001; // 5757 : 169 - 0xa9
      13'h167E: dout  = 8'b11111111; // 5758 : 255 - 0xff
      13'h167F: dout  = 8'b11111100; // 5759 : 252 - 0xfc
      13'h1680: dout  = 8'b00111100; // 5760 :  60 - 0x3c -- Background 0x68
      13'h1681: dout  = 8'b00111100; // 5761 :  60 - 0x3c
      13'h1682: dout  = 8'b00111100; // 5762 :  60 - 0x3c
      13'h1683: dout  = 8'b00111100; // 5763 :  60 - 0x3c
      13'h1684: dout  = 8'b00111100; // 5764 :  60 - 0x3c
      13'h1685: dout  = 8'b00111100; // 5765 :  60 - 0x3c
      13'h1686: dout  = 8'b00111100; // 5766 :  60 - 0x3c
      13'h1687: dout  = 8'b00111100; // 5767 :  60 - 0x3c
      13'h1688: dout  = 8'b00100011; // 5768 :  35 - 0x23
      13'h1689: dout  = 8'b00100011; // 5769 :  35 - 0x23
      13'h168A: dout  = 8'b00100011; // 5770 :  35 - 0x23
      13'h168B: dout  = 8'b00100011; // 5771 :  35 - 0x23
      13'h168C: dout  = 8'b00100011; // 5772 :  35 - 0x23
      13'h168D: dout  = 8'b00100011; // 5773 :  35 - 0x23
      13'h168E: dout  = 8'b00100011; // 5774 :  35 - 0x23
      13'h168F: dout  = 8'b00100011; // 5775 :  35 - 0x23
      13'h1690: dout  = 8'b11111011; // 5776 : 251 - 0xfb -- Background 0x69
      13'h1691: dout  = 8'b11111011; // 5777 : 251 - 0xfb
      13'h1692: dout  = 8'b11111011; // 5778 : 251 - 0xfb
      13'h1693: dout  = 8'b11111011; // 5779 : 251 - 0xfb
      13'h1694: dout  = 8'b11111011; // 5780 : 251 - 0xfb
      13'h1695: dout  = 8'b11111011; // 5781 : 251 - 0xfb
      13'h1696: dout  = 8'b11111011; // 5782 : 251 - 0xfb
      13'h1697: dout  = 8'b11111011; // 5783 : 251 - 0xfb
      13'h1698: dout  = 8'b00000100; // 5784 :   4 - 0x4
      13'h1699: dout  = 8'b00000100; // 5785 :   4 - 0x4
      13'h169A: dout  = 8'b00000100; // 5786 :   4 - 0x4
      13'h169B: dout  = 8'b00000100; // 5787 :   4 - 0x4
      13'h169C: dout  = 8'b00000100; // 5788 :   4 - 0x4
      13'h169D: dout  = 8'b00000100; // 5789 :   4 - 0x4
      13'h169E: dout  = 8'b00000100; // 5790 :   4 - 0x4
      13'h169F: dout  = 8'b00000100; // 5791 :   4 - 0x4
      13'h16A0: dout  = 8'b10111100; // 5792 : 188 - 0xbc -- Background 0x6a
      13'h16A1: dout  = 8'b01011100; // 5793 :  92 - 0x5c
      13'h16A2: dout  = 8'b10111100; // 5794 : 188 - 0xbc
      13'h16A3: dout  = 8'b01011100; // 5795 :  92 - 0x5c
      13'h16A4: dout  = 8'b10111100; // 5796 : 188 - 0xbc
      13'h16A5: dout  = 8'b01011100; // 5797 :  92 - 0x5c
      13'h16A6: dout  = 8'b10111100; // 5798 : 188 - 0xbc
      13'h16A7: dout  = 8'b01011100; // 5799 :  92 - 0x5c
      13'h16A8: dout  = 8'b01000100; // 5800 :  68 - 0x44
      13'h16A9: dout  = 8'b10100100; // 5801 : 164 - 0xa4
      13'h16AA: dout  = 8'b01000100; // 5802 :  68 - 0x44
      13'h16AB: dout  = 8'b10100100; // 5803 : 164 - 0xa4
      13'h16AC: dout  = 8'b01000100; // 5804 :  68 - 0x44
      13'h16AD: dout  = 8'b10100100; // 5805 : 164 - 0xa4
      13'h16AE: dout  = 8'b01000100; // 5806 :  68 - 0x44
      13'h16AF: dout  = 8'b10100100; // 5807 : 164 - 0xa4
      13'h16B0: dout  = 8'b00011111; // 5808 :  31 - 0x1f -- Background 0x6b
      13'h16B1: dout  = 8'b00100000; // 5809 :  32 - 0x20
      13'h16B2: dout  = 8'b01000000; // 5810 :  64 - 0x40
      13'h16B3: dout  = 8'b01000000; // 5811 :  64 - 0x40
      13'h16B4: dout  = 8'b10000000; // 5812 : 128 - 0x80
      13'h16B5: dout  = 8'b10000000; // 5813 : 128 - 0x80
      13'h16B6: dout  = 8'b10000000; // 5814 : 128 - 0x80
      13'h16B7: dout  = 8'b10000001; // 5815 : 129 - 0x81
      13'h16B8: dout  = 8'b00011111; // 5816 :  31 - 0x1f
      13'h16B9: dout  = 8'b00111111; // 5817 :  63 - 0x3f
      13'h16BA: dout  = 8'b01111111; // 5818 : 127 - 0x7f
      13'h16BB: dout  = 8'b01111111; // 5819 : 127 - 0x7f
      13'h16BC: dout  = 8'b11111111; // 5820 : 255 - 0xff
      13'h16BD: dout  = 8'b11111111; // 5821 : 255 - 0xff
      13'h16BE: dout  = 8'b11111111; // 5822 : 255 - 0xff
      13'h16BF: dout  = 8'b11111110; // 5823 : 254 - 0xfe
      13'h16C0: dout  = 8'b11111111; // 5824 : 255 - 0xff -- Background 0x6c
      13'h16C1: dout  = 8'b10000000; // 5825 : 128 - 0x80
      13'h16C2: dout  = 8'b10000000; // 5826 : 128 - 0x80
      13'h16C3: dout  = 8'b11000000; // 5827 : 192 - 0xc0
      13'h16C4: dout  = 8'b11111111; // 5828 : 255 - 0xff
      13'h16C5: dout  = 8'b11111111; // 5829 : 255 - 0xff
      13'h16C6: dout  = 8'b11111110; // 5830 : 254 - 0xfe
      13'h16C7: dout  = 8'b11111110; // 5831 : 254 - 0xfe
      13'h16C8: dout  = 8'b11111111; // 5832 : 255 - 0xff
      13'h16C9: dout  = 8'b01111111; // 5833 : 127 - 0x7f
      13'h16CA: dout  = 8'b01111111; // 5834 : 127 - 0x7f
      13'h16CB: dout  = 8'b00111111; // 5835 :  63 - 0x3f
      13'h16CC: dout  = 8'b00000000; // 5836 :   0 - 0x0
      13'h16CD: dout  = 8'b00000000; // 5837 :   0 - 0x0
      13'h16CE: dout  = 8'b00000001; // 5838 :   1 - 0x1
      13'h16CF: dout  = 8'b00000001; // 5839 :   1 - 0x1
      13'h16D0: dout  = 8'b11111111; // 5840 : 255 - 0xff -- Background 0x6d
      13'h16D1: dout  = 8'b01111111; // 5841 : 127 - 0x7f
      13'h16D2: dout  = 8'b01111111; // 5842 : 127 - 0x7f
      13'h16D3: dout  = 8'b11111111; // 5843 : 255 - 0xff
      13'h16D4: dout  = 8'b11111111; // 5844 : 255 - 0xff
      13'h16D5: dout  = 8'b00000111; // 5845 :   7 - 0x7
      13'h16D6: dout  = 8'b00000011; // 5846 :   3 - 0x3
      13'h16D7: dout  = 8'b00000011; // 5847 :   3 - 0x3
      13'h16D8: dout  = 8'b11111111; // 5848 : 255 - 0xff
      13'h16D9: dout  = 8'b10000000; // 5849 : 128 - 0x80
      13'h16DA: dout  = 8'b10000000; // 5850 : 128 - 0x80
      13'h16DB: dout  = 8'b00000000; // 5851 :   0 - 0x0
      13'h16DC: dout  = 8'b00000000; // 5852 :   0 - 0x0
      13'h16DD: dout  = 8'b11111000; // 5853 : 248 - 0xf8
      13'h16DE: dout  = 8'b11111100; // 5854 : 252 - 0xfc
      13'h16DF: dout  = 8'b11111100; // 5855 : 252 - 0xfc
      13'h16E0: dout  = 8'b11111111; // 5856 : 255 - 0xff -- Background 0x6e
      13'h16E1: dout  = 8'b00000000; // 5857 :   0 - 0x0
      13'h16E2: dout  = 8'b00000000; // 5858 :   0 - 0x0
      13'h16E3: dout  = 8'b00000000; // 5859 :   0 - 0x0
      13'h16E4: dout  = 8'b00000000; // 5860 :   0 - 0x0
      13'h16E5: dout  = 8'b10000001; // 5861 : 129 - 0x81
      13'h16E6: dout  = 8'b11000011; // 5862 : 195 - 0xc3
      13'h16E7: dout  = 8'b11111111; // 5863 : 255 - 0xff
      13'h16E8: dout  = 8'b11111111; // 5864 : 255 - 0xff
      13'h16E9: dout  = 8'b11111111; // 5865 : 255 - 0xff
      13'h16EA: dout  = 8'b11111111; // 5866 : 255 - 0xff
      13'h16EB: dout  = 8'b11111111; // 5867 : 255 - 0xff
      13'h16EC: dout  = 8'b11111111; // 5868 : 255 - 0xff
      13'h16ED: dout  = 8'b01111110; // 5869 : 126 - 0x7e
      13'h16EE: dout  = 8'b00111100; // 5870 :  60 - 0x3c
      13'h16EF: dout  = 8'b00000000; // 5871 :   0 - 0x0
      13'h16F0: dout  = 8'b11111000; // 5872 : 248 - 0xf8 -- Background 0x6f
      13'h16F1: dout  = 8'b11111100; // 5873 : 252 - 0xfc
      13'h16F2: dout  = 8'b11111110; // 5874 : 254 - 0xfe
      13'h16F3: dout  = 8'b11111110; // 5875 : 254 - 0xfe
      13'h16F4: dout  = 8'b11100011; // 5876 : 227 - 0xe3
      13'h16F5: dout  = 8'b11000001; // 5877 : 193 - 0xc1
      13'h16F6: dout  = 8'b10000001; // 5878 : 129 - 0x81
      13'h16F7: dout  = 8'b10000001; // 5879 : 129 - 0x81
      13'h16F8: dout  = 8'b11111000; // 5880 : 248 - 0xf8
      13'h16F9: dout  = 8'b00000100; // 5881 :   4 - 0x4
      13'h16FA: dout  = 8'b00000010; // 5882 :   2 - 0x2
      13'h16FB: dout  = 8'b00000010; // 5883 :   2 - 0x2
      13'h16FC: dout  = 8'b00011101; // 5884 :  29 - 0x1d
      13'h16FD: dout  = 8'b00111111; // 5885 :  63 - 0x3f
      13'h16FE: dout  = 8'b01111111; // 5886 : 127 - 0x7f
      13'h16FF: dout  = 8'b01111111; // 5887 : 127 - 0x7f
      13'h1700: dout  = 8'b10000011; // 5888 : 131 - 0x83 -- Background 0x70
      13'h1701: dout  = 8'b11111111; // 5889 : 255 - 0xff
      13'h1702: dout  = 8'b11111111; // 5890 : 255 - 0xff
      13'h1703: dout  = 8'b11111111; // 5891 : 255 - 0xff
      13'h1704: dout  = 8'b11111111; // 5892 : 255 - 0xff
      13'h1705: dout  = 8'b11111111; // 5893 : 255 - 0xff
      13'h1706: dout  = 8'b01111111; // 5894 : 127 - 0x7f
      13'h1707: dout  = 8'b00011111; // 5895 :  31 - 0x1f
      13'h1708: dout  = 8'b11111100; // 5896 : 252 - 0xfc
      13'h1709: dout  = 8'b10000000; // 5897 : 128 - 0x80
      13'h170A: dout  = 8'b10000000; // 5898 : 128 - 0x80
      13'h170B: dout  = 8'b10000000; // 5899 : 128 - 0x80
      13'h170C: dout  = 8'b10000000; // 5900 : 128 - 0x80
      13'h170D: dout  = 8'b10000000; // 5901 : 128 - 0x80
      13'h170E: dout  = 8'b01100000; // 5902 :  96 - 0x60
      13'h170F: dout  = 8'b00011111; // 5903 :  31 - 0x1f
      13'h1710: dout  = 8'b11111100; // 5904 : 252 - 0xfc -- Background 0x71
      13'h1711: dout  = 8'b11111100; // 5905 : 252 - 0xfc
      13'h1712: dout  = 8'b11111100; // 5906 : 252 - 0xfc
      13'h1713: dout  = 8'b11111100; // 5907 : 252 - 0xfc
      13'h1714: dout  = 8'b11111110; // 5908 : 254 - 0xfe
      13'h1715: dout  = 8'b11111110; // 5909 : 254 - 0xfe
      13'h1716: dout  = 8'b11111111; // 5910 : 255 - 0xff
      13'h1717: dout  = 8'b11111111; // 5911 : 255 - 0xff
      13'h1718: dout  = 8'b00000011; // 5912 :   3 - 0x3
      13'h1719: dout  = 8'b00000011; // 5913 :   3 - 0x3
      13'h171A: dout  = 8'b00000011; // 5914 :   3 - 0x3
      13'h171B: dout  = 8'b00000011; // 5915 :   3 - 0x3
      13'h171C: dout  = 8'b00000001; // 5916 :   1 - 0x1
      13'h171D: dout  = 8'b00000001; // 5917 :   1 - 0x1
      13'h171E: dout  = 8'b00000000; // 5918 :   0 - 0x0
      13'h171F: dout  = 8'b11111111; // 5919 : 255 - 0xff
      13'h1720: dout  = 8'b00000001; // 5920 :   1 - 0x1 -- Background 0x72
      13'h1721: dout  = 8'b00000001; // 5921 :   1 - 0x1
      13'h1722: dout  = 8'b00000001; // 5922 :   1 - 0x1
      13'h1723: dout  = 8'b00000001; // 5923 :   1 - 0x1
      13'h1724: dout  = 8'b00000011; // 5924 :   3 - 0x3
      13'h1725: dout  = 8'b00000011; // 5925 :   3 - 0x3
      13'h1726: dout  = 8'b00000111; // 5926 :   7 - 0x7
      13'h1727: dout  = 8'b11111111; // 5927 : 255 - 0xff
      13'h1728: dout  = 8'b11111110; // 5928 : 254 - 0xfe
      13'h1729: dout  = 8'b11111110; // 5929 : 254 - 0xfe
      13'h172A: dout  = 8'b11111110; // 5930 : 254 - 0xfe
      13'h172B: dout  = 8'b11111110; // 5931 : 254 - 0xfe
      13'h172C: dout  = 8'b11111100; // 5932 : 252 - 0xfc
      13'h172D: dout  = 8'b11111100; // 5933 : 252 - 0xfc
      13'h172E: dout  = 8'b11111000; // 5934 : 248 - 0xf8
      13'h172F: dout  = 8'b11111111; // 5935 : 255 - 0xff
      13'h1730: dout  = 8'b11111111; // 5936 : 255 - 0xff -- Background 0x73
      13'h1731: dout  = 8'b11111111; // 5937 : 255 - 0xff
      13'h1732: dout  = 8'b11111111; // 5938 : 255 - 0xff
      13'h1733: dout  = 8'b11111111; // 5939 : 255 - 0xff
      13'h1734: dout  = 8'b11111111; // 5940 : 255 - 0xff
      13'h1735: dout  = 8'b11111111; // 5941 : 255 - 0xff
      13'h1736: dout  = 8'b11111111; // 5942 : 255 - 0xff
      13'h1737: dout  = 8'b11111111; // 5943 : 255 - 0xff
      13'h1738: dout  = 8'b00000000; // 5944 :   0 - 0x0
      13'h1739: dout  = 8'b00000000; // 5945 :   0 - 0x0
      13'h173A: dout  = 8'b00000000; // 5946 :   0 - 0x0
      13'h173B: dout  = 8'b00000000; // 5947 :   0 - 0x0
      13'h173C: dout  = 8'b00000000; // 5948 :   0 - 0x0
      13'h173D: dout  = 8'b00000000; // 5949 :   0 - 0x0
      13'h173E: dout  = 8'b00000000; // 5950 :   0 - 0x0
      13'h173F: dout  = 8'b11111111; // 5951 : 255 - 0xff
      13'h1740: dout  = 8'b10000001; // 5952 : 129 - 0x81 -- Background 0x74
      13'h1741: dout  = 8'b11000001; // 5953 : 193 - 0xc1
      13'h1742: dout  = 8'b11100011; // 5954 : 227 - 0xe3
      13'h1743: dout  = 8'b11111111; // 5955 : 255 - 0xff
      13'h1744: dout  = 8'b11111111; // 5956 : 255 - 0xff
      13'h1745: dout  = 8'b11111111; // 5957 : 255 - 0xff
      13'h1746: dout  = 8'b11111111; // 5958 : 255 - 0xff
      13'h1747: dout  = 8'b11111110; // 5959 : 254 - 0xfe
      13'h1748: dout  = 8'b01111111; // 5960 : 127 - 0x7f
      13'h1749: dout  = 8'b00111111; // 5961 :  63 - 0x3f
      13'h174A: dout  = 8'b00011101; // 5962 :  29 - 0x1d
      13'h174B: dout  = 8'b00000001; // 5963 :   1 - 0x1
      13'h174C: dout  = 8'b00000001; // 5964 :   1 - 0x1
      13'h174D: dout  = 8'b00000001; // 5965 :   1 - 0x1
      13'h174E: dout  = 8'b00000011; // 5966 :   3 - 0x3
      13'h174F: dout  = 8'b11111110; // 5967 : 254 - 0xfe
      13'h1750: dout  = 8'b11111111; // 5968 : 255 - 0xff -- Background 0x75
      13'h1751: dout  = 8'b11111111; // 5969 : 255 - 0xff
      13'h1752: dout  = 8'b11111111; // 5970 : 255 - 0xff
      13'h1753: dout  = 8'b11111111; // 5971 : 255 - 0xff
      13'h1754: dout  = 8'b11111111; // 5972 : 255 - 0xff
      13'h1755: dout  = 8'b11111011; // 5973 : 251 - 0xfb
      13'h1756: dout  = 8'b10110101; // 5974 : 181 - 0xb5
      13'h1757: dout  = 8'b11001110; // 5975 : 206 - 0xce
      13'h1758: dout  = 8'b10000000; // 5976 : 128 - 0x80
      13'h1759: dout  = 8'b10000000; // 5977 : 128 - 0x80
      13'h175A: dout  = 8'b10000000; // 5978 : 128 - 0x80
      13'h175B: dout  = 8'b10000000; // 5979 : 128 - 0x80
      13'h175C: dout  = 8'b10000000; // 5980 : 128 - 0x80
      13'h175D: dout  = 8'b10000100; // 5981 : 132 - 0x84
      13'h175E: dout  = 8'b11001010; // 5982 : 202 - 0xca
      13'h175F: dout  = 8'b10110001; // 5983 : 177 - 0xb1
      13'h1760: dout  = 8'b11111111; // 5984 : 255 - 0xff -- Background 0x76
      13'h1761: dout  = 8'b11111111; // 5985 : 255 - 0xff
      13'h1762: dout  = 8'b11111111; // 5986 : 255 - 0xff
      13'h1763: dout  = 8'b11111111; // 5987 : 255 - 0xff
      13'h1764: dout  = 8'b11111111; // 5988 : 255 - 0xff
      13'h1765: dout  = 8'b11011111; // 5989 : 223 - 0xdf
      13'h1766: dout  = 8'b10101101; // 5990 : 173 - 0xad
      13'h1767: dout  = 8'b01110011; // 5991 : 115 - 0x73
      13'h1768: dout  = 8'b00000001; // 5992 :   1 - 0x1
      13'h1769: dout  = 8'b00000001; // 5993 :   1 - 0x1
      13'h176A: dout  = 8'b00000001; // 5994 :   1 - 0x1
      13'h176B: dout  = 8'b00000001; // 5995 :   1 - 0x1
      13'h176C: dout  = 8'b00000001; // 5996 :   1 - 0x1
      13'h176D: dout  = 8'b00100001; // 5997 :  33 - 0x21
      13'h176E: dout  = 8'b01010011; // 5998 :  83 - 0x53
      13'h176F: dout  = 8'b10001101; // 5999 : 141 - 0x8d
      13'h1770: dout  = 8'b01110111; // 6000 : 119 - 0x77 -- Background 0x77
      13'h1771: dout  = 8'b01110111; // 6001 : 119 - 0x77
      13'h1772: dout  = 8'b01110111; // 6002 : 119 - 0x77
      13'h1773: dout  = 8'b01110111; // 6003 : 119 - 0x77
      13'h1774: dout  = 8'b01110111; // 6004 : 119 - 0x77
      13'h1775: dout  = 8'b01110111; // 6005 : 119 - 0x77
      13'h1776: dout  = 8'b01110111; // 6006 : 119 - 0x77
      13'h1777: dout  = 8'b01110111; // 6007 : 119 - 0x77
      13'h1778: dout  = 8'b00000000; // 6008 :   0 - 0x0
      13'h1779: dout  = 8'b00000000; // 6009 :   0 - 0x0
      13'h177A: dout  = 8'b00000000; // 6010 :   0 - 0x0
      13'h177B: dout  = 8'b00000000; // 6011 :   0 - 0x0
      13'h177C: dout  = 8'b01110111; // 6012 : 119 - 0x77
      13'h177D: dout  = 8'b11111111; // 6013 : 255 - 0xff
      13'h177E: dout  = 8'b11111111; // 6014 : 255 - 0xff
      13'h177F: dout  = 8'b11111111; // 6015 : 255 - 0xff
      13'h1780: dout  = 8'b00000000; // 6016 :   0 - 0x0 -- Background 0x78
      13'h1781: dout  = 8'b00000000; // 6017 :   0 - 0x0
      13'h1782: dout  = 8'b00000000; // 6018 :   0 - 0x0
      13'h1783: dout  = 8'b00000000; // 6019 :   0 - 0x0
      13'h1784: dout  = 8'b00000000; // 6020 :   0 - 0x0
      13'h1785: dout  = 8'b00000000; // 6021 :   0 - 0x0
      13'h1786: dout  = 8'b00000000; // 6022 :   0 - 0x0
      13'h1787: dout  = 8'b11111111; // 6023 : 255 - 0xff
      13'h1788: dout  = 8'b11111111; // 6024 : 255 - 0xff
      13'h1789: dout  = 8'b11111111; // 6025 : 255 - 0xff
      13'h178A: dout  = 8'b11111111; // 6026 : 255 - 0xff
      13'h178B: dout  = 8'b11111111; // 6027 : 255 - 0xff
      13'h178C: dout  = 8'b11111111; // 6028 : 255 - 0xff
      13'h178D: dout  = 8'b11111111; // 6029 : 255 - 0xff
      13'h178E: dout  = 8'b11111111; // 6030 : 255 - 0xff
      13'h178F: dout  = 8'b11111111; // 6031 : 255 - 0xff
      13'h1790: dout  = 8'b01110111; // 6032 : 119 - 0x77 -- Background 0x79
      13'h1791: dout  = 8'b01110111; // 6033 : 119 - 0x77
      13'h1792: dout  = 8'b01110111; // 6034 : 119 - 0x77
      13'h1793: dout  = 8'b01110111; // 6035 : 119 - 0x77
      13'h1794: dout  = 8'b00000000; // 6036 :   0 - 0x0
      13'h1795: dout  = 8'b00000000; // 6037 :   0 - 0x0
      13'h1796: dout  = 8'b00000000; // 6038 :   0 - 0x0
      13'h1797: dout  = 8'b00000000; // 6039 :   0 - 0x0
      13'h1798: dout  = 8'b11111111; // 6040 : 255 - 0xff
      13'h1799: dout  = 8'b11111111; // 6041 : 255 - 0xff
      13'h179A: dout  = 8'b11111111; // 6042 : 255 - 0xff
      13'h179B: dout  = 8'b01110111; // 6043 : 119 - 0x77
      13'h179C: dout  = 8'b01110111; // 6044 : 119 - 0x77
      13'h179D: dout  = 8'b01110111; // 6045 : 119 - 0x77
      13'h179E: dout  = 8'b01110111; // 6046 : 119 - 0x77
      13'h179F: dout  = 8'b01110111; // 6047 : 119 - 0x77
      13'h17A0: dout  = 8'b00000001; // 6048 :   1 - 0x1 -- Background 0x7a
      13'h17A1: dout  = 8'b00000001; // 6049 :   1 - 0x1
      13'h17A2: dout  = 8'b00000001; // 6050 :   1 - 0x1
      13'h17A3: dout  = 8'b00011001; // 6051 :  25 - 0x19
      13'h17A4: dout  = 8'b00011101; // 6052 :  29 - 0x1d
      13'h17A5: dout  = 8'b00001101; // 6053 :  13 - 0xd
      13'h17A6: dout  = 8'b00000001; // 6054 :   1 - 0x1
      13'h17A7: dout  = 8'b11111110; // 6055 : 254 - 0xfe
      13'h17A8: dout  = 8'b11111111; // 6056 : 255 - 0xff
      13'h17A9: dout  = 8'b11111111; // 6057 : 255 - 0xff
      13'h17AA: dout  = 8'b11111111; // 6058 : 255 - 0xff
      13'h17AB: dout  = 8'b11100111; // 6059 : 231 - 0xe7
      13'h17AC: dout  = 8'b11100111; // 6060 : 231 - 0xe7
      13'h17AD: dout  = 8'b11111111; // 6061 : 255 - 0xff
      13'h17AE: dout  = 8'b11111111; // 6062 : 255 - 0xff
      13'h17AF: dout  = 8'b11111110; // 6063 : 254 - 0xfe
      13'h17B0: dout  = 8'b00100000; // 6064 :  32 - 0x20 -- Background 0x7b
      13'h17B1: dout  = 8'b01111000; // 6065 : 120 - 0x78
      13'h17B2: dout  = 8'b01111111; // 6066 : 127 - 0x7f
      13'h17B3: dout  = 8'b11111110; // 6067 : 254 - 0xfe
      13'h17B4: dout  = 8'b11111110; // 6068 : 254 - 0xfe
      13'h17B5: dout  = 8'b11111110; // 6069 : 254 - 0xfe
      13'h17B6: dout  = 8'b11111110; // 6070 : 254 - 0xfe
      13'h17B7: dout  = 8'b11111110; // 6071 : 254 - 0xfe
      13'h17B8: dout  = 8'b00000000; // 6072 :   0 - 0x0
      13'h17B9: dout  = 8'b00100001; // 6073 :  33 - 0x21
      13'h17BA: dout  = 8'b00100001; // 6074 :  33 - 0x21
      13'h17BB: dout  = 8'b01000001; // 6075 :  65 - 0x41
      13'h17BC: dout  = 8'b01000001; // 6076 :  65 - 0x41
      13'h17BD: dout  = 8'b01000001; // 6077 :  65 - 0x41
      13'h17BE: dout  = 8'b01000001; // 6078 :  65 - 0x41
      13'h17BF: dout  = 8'b01000001; // 6079 :  65 - 0x41
      13'h17C0: dout  = 8'b00000100; // 6080 :   4 - 0x4 -- Background 0x7c
      13'h17C1: dout  = 8'b10011010; // 6081 : 154 - 0x9a
      13'h17C2: dout  = 8'b11111010; // 6082 : 250 - 0xfa
      13'h17C3: dout  = 8'b11111101; // 6083 : 253 - 0xfd
      13'h17C4: dout  = 8'b11111101; // 6084 : 253 - 0xfd
      13'h17C5: dout  = 8'b11111101; // 6085 : 253 - 0xfd
      13'h17C6: dout  = 8'b11111101; // 6086 : 253 - 0xfd
      13'h17C7: dout  = 8'b11111101; // 6087 : 253 - 0xfd
      13'h17C8: dout  = 8'b00000000; // 6088 :   0 - 0x0
      13'h17C9: dout  = 8'b10000000; // 6089 : 128 - 0x80
      13'h17CA: dout  = 8'b10000000; // 6090 : 128 - 0x80
      13'h17CB: dout  = 8'b10000000; // 6091 : 128 - 0x80
      13'h17CC: dout  = 8'b10000000; // 6092 : 128 - 0x80
      13'h17CD: dout  = 8'b10000000; // 6093 : 128 - 0x80
      13'h17CE: dout  = 8'b10000000; // 6094 : 128 - 0x80
      13'h17CF: dout  = 8'b10000000; // 6095 : 128 - 0x80
      13'h17D0: dout  = 8'b01111110; // 6096 : 126 - 0x7e -- Background 0x7d
      13'h17D1: dout  = 8'b00111000; // 6097 :  56 - 0x38
      13'h17D2: dout  = 8'b00100001; // 6098 :  33 - 0x21
      13'h17D3: dout  = 8'b00000000; // 6099 :   0 - 0x0
      13'h17D4: dout  = 8'b00000001; // 6100 :   1 - 0x1
      13'h17D5: dout  = 8'b00000000; // 6101 :   0 - 0x0
      13'h17D6: dout  = 8'b00000001; // 6102 :   1 - 0x1
      13'h17D7: dout  = 8'b00000000; // 6103 :   0 - 0x0
      13'h17D8: dout  = 8'b00100001; // 6104 :  33 - 0x21
      13'h17D9: dout  = 8'b00100001; // 6105 :  33 - 0x21
      13'h17DA: dout  = 8'b00000001; // 6106 :   1 - 0x1
      13'h17DB: dout  = 8'b00000001; // 6107 :   1 - 0x1
      13'h17DC: dout  = 8'b00000001; // 6108 :   1 - 0x1
      13'h17DD: dout  = 8'b00000001; // 6109 :   1 - 0x1
      13'h17DE: dout  = 8'b00000001; // 6110 :   1 - 0x1
      13'h17DF: dout  = 8'b00000001; // 6111 :   1 - 0x1
      13'h17E0: dout  = 8'b11111010; // 6112 : 250 - 0xfa -- Background 0x7e
      13'h17E1: dout  = 8'b10001010; // 6113 : 138 - 0x8a
      13'h17E2: dout  = 8'b10000100; // 6114 : 132 - 0x84
      13'h17E3: dout  = 8'b10000000; // 6115 : 128 - 0x80
      13'h17E4: dout  = 8'b10000000; // 6116 : 128 - 0x80
      13'h17E5: dout  = 8'b10000000; // 6117 : 128 - 0x80
      13'h17E6: dout  = 8'b10000000; // 6118 : 128 - 0x80
      13'h17E7: dout  = 8'b10000000; // 6119 : 128 - 0x80
      13'h17E8: dout  = 8'b10000000; // 6120 : 128 - 0x80
      13'h17E9: dout  = 8'b10000000; // 6121 : 128 - 0x80
      13'h17EA: dout  = 8'b10000000; // 6122 : 128 - 0x80
      13'h17EB: dout  = 8'b10000000; // 6123 : 128 - 0x80
      13'h17EC: dout  = 8'b10000000; // 6124 : 128 - 0x80
      13'h17ED: dout  = 8'b10000000; // 6125 : 128 - 0x80
      13'h17EE: dout  = 8'b10000000; // 6126 : 128 - 0x80
      13'h17EF: dout  = 8'b10000000; // 6127 : 128 - 0x80
      13'h17F0: dout  = 8'b00000010; // 6128 :   2 - 0x2 -- Background 0x7f
      13'h17F1: dout  = 8'b00000100; // 6129 :   4 - 0x4
      13'h17F2: dout  = 8'b00000000; // 6130 :   0 - 0x0
      13'h17F3: dout  = 8'b00010000; // 6131 :  16 - 0x10
      13'h17F4: dout  = 8'b00000000; // 6132 :   0 - 0x0
      13'h17F5: dout  = 8'b01000000; // 6133 :  64 - 0x40
      13'h17F6: dout  = 8'b10000000; // 6134 : 128 - 0x80
      13'h17F7: dout  = 8'b00000000; // 6135 :   0 - 0x0
      13'h17F8: dout  = 8'b00000001; // 6136 :   1 - 0x1
      13'h17F9: dout  = 8'b00000001; // 6137 :   1 - 0x1
      13'h17FA: dout  = 8'b00000110; // 6138 :   6 - 0x6
      13'h17FB: dout  = 8'b00001000; // 6139 :   8 - 0x8
      13'h17FC: dout  = 8'b00011000; // 6140 :  24 - 0x18
      13'h17FD: dout  = 8'b00100000; // 6141 :  32 - 0x20
      13'h17FE: dout  = 8'b00100000; // 6142 :  32 - 0x20
      13'h17FF: dout  = 8'b11000000; // 6143 : 192 - 0xc0
      13'h1800: dout  = 8'b00001011; // 6144 :  11 - 0xb -- Background 0x80
      13'h1801: dout  = 8'b00001011; // 6145 :  11 - 0xb
      13'h1802: dout  = 8'b00111011; // 6146 :  59 - 0x3b
      13'h1803: dout  = 8'b00001011; // 6147 :  11 - 0xb
      13'h1804: dout  = 8'b11111011; // 6148 : 251 - 0xfb
      13'h1805: dout  = 8'b00001011; // 6149 :  11 - 0xb
      13'h1806: dout  = 8'b00001011; // 6150 :  11 - 0xb
      13'h1807: dout  = 8'b00001010; // 6151 :  10 - 0xa
      13'h1808: dout  = 8'b00000100; // 6152 :   4 - 0x4
      13'h1809: dout  = 8'b00000100; // 6153 :   4 - 0x4
      13'h180A: dout  = 8'b11000100; // 6154 : 196 - 0xc4
      13'h180B: dout  = 8'b11110100; // 6155 : 244 - 0xf4
      13'h180C: dout  = 8'b11110100; // 6156 : 244 - 0xf4
      13'h180D: dout  = 8'b00000100; // 6157 :   4 - 0x4
      13'h180E: dout  = 8'b00000100; // 6158 :   4 - 0x4
      13'h180F: dout  = 8'b00000101; // 6159 :   5 - 0x5
      13'h1810: dout  = 8'b10010000; // 6160 : 144 - 0x90 -- Background 0x81
      13'h1811: dout  = 8'b00010000; // 6161 :  16 - 0x10
      13'h1812: dout  = 8'b00011111; // 6162 :  31 - 0x1f
      13'h1813: dout  = 8'b00010000; // 6163 :  16 - 0x10
      13'h1814: dout  = 8'b00011111; // 6164 :  31 - 0x1f
      13'h1815: dout  = 8'b00010000; // 6165 :  16 - 0x10
      13'h1816: dout  = 8'b00010000; // 6166 :  16 - 0x10
      13'h1817: dout  = 8'b10010000; // 6167 : 144 - 0x90
      13'h1818: dout  = 8'b01110000; // 6168 : 112 - 0x70
      13'h1819: dout  = 8'b11110000; // 6169 : 240 - 0xf0
      13'h181A: dout  = 8'b11110000; // 6170 : 240 - 0xf0
      13'h181B: dout  = 8'b11111111; // 6171 : 255 - 0xff
      13'h181C: dout  = 8'b11111111; // 6172 : 255 - 0xff
      13'h181D: dout  = 8'b11110000; // 6173 : 240 - 0xf0
      13'h181E: dout  = 8'b11110000; // 6174 : 240 - 0xf0
      13'h181F: dout  = 8'b01110000; // 6175 : 112 - 0x70
      13'h1820: dout  = 8'b00111111; // 6176 :  63 - 0x3f -- Background 0x82
      13'h1821: dout  = 8'b01111000; // 6177 : 120 - 0x78
      13'h1822: dout  = 8'b11100111; // 6178 : 231 - 0xe7
      13'h1823: dout  = 8'b11001111; // 6179 : 207 - 0xcf
      13'h1824: dout  = 8'b01011000; // 6180 :  88 - 0x58
      13'h1825: dout  = 8'b01011000; // 6181 :  88 - 0x58
      13'h1826: dout  = 8'b01010000; // 6182 :  80 - 0x50
      13'h1827: dout  = 8'b10010000; // 6183 : 144 - 0x90
      13'h1828: dout  = 8'b11000000; // 6184 : 192 - 0xc0
      13'h1829: dout  = 8'b10000111; // 6185 : 135 - 0x87
      13'h182A: dout  = 8'b00011000; // 6186 :  24 - 0x18
      13'h182B: dout  = 8'b10110000; // 6187 : 176 - 0xb0
      13'h182C: dout  = 8'b11100111; // 6188 : 231 - 0xe7
      13'h182D: dout  = 8'b11100111; // 6189 : 231 - 0xe7
      13'h182E: dout  = 8'b11101111; // 6190 : 239 - 0xef
      13'h182F: dout  = 8'b11101111; // 6191 : 239 - 0xef
      13'h1830: dout  = 8'b10110000; // 6192 : 176 - 0xb0 -- Background 0x83
      13'h1831: dout  = 8'b11111100; // 6193 : 252 - 0xfc
      13'h1832: dout  = 8'b11100010; // 6194 : 226 - 0xe2
      13'h1833: dout  = 8'b11000001; // 6195 : 193 - 0xc1
      13'h1834: dout  = 8'b11000001; // 6196 : 193 - 0xc1
      13'h1835: dout  = 8'b10000011; // 6197 : 131 - 0x83
      13'h1836: dout  = 8'b10001111; // 6198 : 143 - 0x8f
      13'h1837: dout  = 8'b01111110; // 6199 : 126 - 0x7e
      13'h1838: dout  = 8'b01101111; // 6200 : 111 - 0x6f
      13'h1839: dout  = 8'b01000011; // 6201 :  67 - 0x43
      13'h183A: dout  = 8'b01011101; // 6202 :  93 - 0x5d
      13'h183B: dout  = 8'b00111111; // 6203 :  63 - 0x3f
      13'h183C: dout  = 8'b00111111; // 6204 :  63 - 0x3f
      13'h183D: dout  = 8'b01111111; // 6205 : 127 - 0x7f
      13'h183E: dout  = 8'b01111111; // 6206 : 127 - 0x7f
      13'h183F: dout  = 8'b11111111; // 6207 : 255 - 0xff
      13'h1840: dout  = 8'b11111110; // 6208 : 254 - 0xfe -- Background 0x84
      13'h1841: dout  = 8'b00000011; // 6209 :   3 - 0x3
      13'h1842: dout  = 8'b00001111; // 6210 :  15 - 0xf
      13'h1843: dout  = 8'b10010001; // 6211 : 145 - 0x91
      13'h1844: dout  = 8'b01110000; // 6212 : 112 - 0x70
      13'h1845: dout  = 8'b01100000; // 6213 :  96 - 0x60
      13'h1846: dout  = 8'b00100000; // 6214 :  32 - 0x20
      13'h1847: dout  = 8'b00110001; // 6215 :  49 - 0x31
      13'h1848: dout  = 8'b00000011; // 6216 :   3 - 0x3
      13'h1849: dout  = 8'b11111111; // 6217 : 255 - 0xff
      13'h184A: dout  = 8'b11110001; // 6218 : 241 - 0xf1
      13'h184B: dout  = 8'b01101110; // 6219 : 110 - 0x6e
      13'h184C: dout  = 8'b11001111; // 6220 : 207 - 0xcf
      13'h184D: dout  = 8'b11011111; // 6221 : 223 - 0xdf
      13'h184E: dout  = 8'b11111111; // 6222 : 255 - 0xff
      13'h184F: dout  = 8'b11111111; // 6223 : 255 - 0xff
      13'h1850: dout  = 8'b00111111; // 6224 :  63 - 0x3f -- Background 0x85
      13'h1851: dout  = 8'b00111111; // 6225 :  63 - 0x3f
      13'h1852: dout  = 8'b00011101; // 6226 :  29 - 0x1d
      13'h1853: dout  = 8'b00111001; // 6227 :  57 - 0x39
      13'h1854: dout  = 8'b01111011; // 6228 : 123 - 0x7b
      13'h1855: dout  = 8'b11110011; // 6229 : 243 - 0xf3
      13'h1856: dout  = 8'b10000110; // 6230 : 134 - 0x86
      13'h1857: dout  = 8'b11111110; // 6231 : 254 - 0xfe
      13'h1858: dout  = 8'b11111101; // 6232 : 253 - 0xfd
      13'h1859: dout  = 8'b11111011; // 6233 : 251 - 0xfb
      13'h185A: dout  = 8'b11111011; // 6234 : 251 - 0xfb
      13'h185B: dout  = 8'b11110111; // 6235 : 247 - 0xf7
      13'h185C: dout  = 8'b11110111; // 6236 : 247 - 0xf7
      13'h185D: dout  = 8'b00001111; // 6237 :  15 - 0xf
      13'h185E: dout  = 8'b01111111; // 6238 : 127 - 0x7f
      13'h185F: dout  = 8'b11111111; // 6239 : 255 - 0xff
      13'h1860: dout  = 8'b11111111; // 6240 : 255 - 0xff -- Background 0x86
      13'h1861: dout  = 8'b11111111; // 6241 : 255 - 0xff
      13'h1862: dout  = 8'b11111111; // 6242 : 255 - 0xff
      13'h1863: dout  = 8'b11111111; // 6243 : 255 - 0xff
      13'h1864: dout  = 8'b11111111; // 6244 : 255 - 0xff
      13'h1865: dout  = 8'b10000000; // 6245 : 128 - 0x80
      13'h1866: dout  = 8'b10000000; // 6246 : 128 - 0x80
      13'h1867: dout  = 8'b11111111; // 6247 : 255 - 0xff
      13'h1868: dout  = 8'b11111111; // 6248 : 255 - 0xff
      13'h1869: dout  = 8'b10000000; // 6249 : 128 - 0x80
      13'h186A: dout  = 8'b10000000; // 6250 : 128 - 0x80
      13'h186B: dout  = 8'b10000000; // 6251 : 128 - 0x80
      13'h186C: dout  = 8'b10000000; // 6252 : 128 - 0x80
      13'h186D: dout  = 8'b11111111; // 6253 : 255 - 0xff
      13'h186E: dout  = 8'b11111111; // 6254 : 255 - 0xff
      13'h186F: dout  = 8'b10000000; // 6255 : 128 - 0x80
      13'h1870: dout  = 8'b11111110; // 6256 : 254 - 0xfe -- Background 0x87
      13'h1871: dout  = 8'b11111111; // 6257 : 255 - 0xff
      13'h1872: dout  = 8'b11111111; // 6258 : 255 - 0xff
      13'h1873: dout  = 8'b11111111; // 6259 : 255 - 0xff
      13'h1874: dout  = 8'b11111111; // 6260 : 255 - 0xff
      13'h1875: dout  = 8'b00000011; // 6261 :   3 - 0x3
      13'h1876: dout  = 8'b00000011; // 6262 :   3 - 0x3
      13'h1877: dout  = 8'b11111111; // 6263 : 255 - 0xff
      13'h1878: dout  = 8'b11111110; // 6264 : 254 - 0xfe
      13'h1879: dout  = 8'b00000011; // 6265 :   3 - 0x3
      13'h187A: dout  = 8'b00000011; // 6266 :   3 - 0x3
      13'h187B: dout  = 8'b00000011; // 6267 :   3 - 0x3
      13'h187C: dout  = 8'b00000011; // 6268 :   3 - 0x3
      13'h187D: dout  = 8'b11111111; // 6269 : 255 - 0xff
      13'h187E: dout  = 8'b11111111; // 6270 : 255 - 0xff
      13'h187F: dout  = 8'b00000011; // 6271 :   3 - 0x3
      13'h1880: dout  = 8'b00000000; // 6272 :   0 - 0x0 -- Background 0x88
      13'h1881: dout  = 8'b11111111; // 6273 : 255 - 0xff
      13'h1882: dout  = 8'b11111111; // 6274 : 255 - 0xff
      13'h1883: dout  = 8'b11111111; // 6275 : 255 - 0xff
      13'h1884: dout  = 8'b11111111; // 6276 : 255 - 0xff
      13'h1885: dout  = 8'b11111111; // 6277 : 255 - 0xff
      13'h1886: dout  = 8'b00000000; // 6278 :   0 - 0x0
      13'h1887: dout  = 8'b00000000; // 6279 :   0 - 0x0
      13'h1888: dout  = 8'b00000000; // 6280 :   0 - 0x0
      13'h1889: dout  = 8'b11111111; // 6281 : 255 - 0xff
      13'h188A: dout  = 8'b00000000; // 6282 :   0 - 0x0
      13'h188B: dout  = 8'b00000000; // 6283 :   0 - 0x0
      13'h188C: dout  = 8'b00000000; // 6284 :   0 - 0x0
      13'h188D: dout  = 8'b00000000; // 6285 :   0 - 0x0
      13'h188E: dout  = 8'b11111111; // 6286 : 255 - 0xff
      13'h188F: dout  = 8'b11111111; // 6287 : 255 - 0xff
      13'h1890: dout  = 8'b00111100; // 6288 :  60 - 0x3c -- Background 0x89
      13'h1891: dout  = 8'b11111100; // 6289 : 252 - 0xfc
      13'h1892: dout  = 8'b11111100; // 6290 : 252 - 0xfc
      13'h1893: dout  = 8'b11111100; // 6291 : 252 - 0xfc
      13'h1894: dout  = 8'b11111100; // 6292 : 252 - 0xfc
      13'h1895: dout  = 8'b11111100; // 6293 : 252 - 0xfc
      13'h1896: dout  = 8'b00000100; // 6294 :   4 - 0x4
      13'h1897: dout  = 8'b00000100; // 6295 :   4 - 0x4
      13'h1898: dout  = 8'b00100011; // 6296 :  35 - 0x23
      13'h1899: dout  = 8'b11110011; // 6297 : 243 - 0xf3
      13'h189A: dout  = 8'b00001011; // 6298 :  11 - 0xb
      13'h189B: dout  = 8'b00001011; // 6299 :  11 - 0xb
      13'h189C: dout  = 8'b00001011; // 6300 :  11 - 0xb
      13'h189D: dout  = 8'b00000111; // 6301 :   7 - 0x7
      13'h189E: dout  = 8'b11111111; // 6302 : 255 - 0xff
      13'h189F: dout  = 8'b11111111; // 6303 : 255 - 0xff
      13'h18A0: dout  = 8'b11111111; // 6304 : 255 - 0xff -- Background 0x8a
      13'h18A1: dout  = 8'b11111111; // 6305 : 255 - 0xff
      13'h18A2: dout  = 8'b11111111; // 6306 : 255 - 0xff
      13'h18A3: dout  = 8'b11111111; // 6307 : 255 - 0xff
      13'h18A4: dout  = 8'b10000000; // 6308 : 128 - 0x80
      13'h18A5: dout  = 8'b11111111; // 6309 : 255 - 0xff
      13'h18A6: dout  = 8'b11111111; // 6310 : 255 - 0xff
      13'h18A7: dout  = 8'b11111111; // 6311 : 255 - 0xff
      13'h18A8: dout  = 8'b10000000; // 6312 : 128 - 0x80
      13'h18A9: dout  = 8'b10000000; // 6313 : 128 - 0x80
      13'h18AA: dout  = 8'b10000000; // 6314 : 128 - 0x80
      13'h18AB: dout  = 8'b10000000; // 6315 : 128 - 0x80
      13'h18AC: dout  = 8'b11111111; // 6316 : 255 - 0xff
      13'h18AD: dout  = 8'b10000000; // 6317 : 128 - 0x80
      13'h18AE: dout  = 8'b10000000; // 6318 : 128 - 0x80
      13'h18AF: dout  = 8'b10000000; // 6319 : 128 - 0x80
      13'h18B0: dout  = 8'b11111111; // 6320 : 255 - 0xff -- Background 0x8b
      13'h18B1: dout  = 8'b11111111; // 6321 : 255 - 0xff
      13'h18B2: dout  = 8'b11111111; // 6322 : 255 - 0xff
      13'h18B3: dout  = 8'b11111111; // 6323 : 255 - 0xff
      13'h18B4: dout  = 8'b00000011; // 6324 :   3 - 0x3
      13'h18B5: dout  = 8'b11111111; // 6325 : 255 - 0xff
      13'h18B6: dout  = 8'b11111111; // 6326 : 255 - 0xff
      13'h18B7: dout  = 8'b11111111; // 6327 : 255 - 0xff
      13'h18B8: dout  = 8'b00000011; // 6328 :   3 - 0x3
      13'h18B9: dout  = 8'b00000011; // 6329 :   3 - 0x3
      13'h18BA: dout  = 8'b00000011; // 6330 :   3 - 0x3
      13'h18BB: dout  = 8'b00000011; // 6331 :   3 - 0x3
      13'h18BC: dout  = 8'b11111111; // 6332 : 255 - 0xff
      13'h18BD: dout  = 8'b00000011; // 6333 :   3 - 0x3
      13'h18BE: dout  = 8'b00000011; // 6334 :   3 - 0x3
      13'h18BF: dout  = 8'b00000011; // 6335 :   3 - 0x3
      13'h18C0: dout  = 8'b11111111; // 6336 : 255 - 0xff -- Background 0x8c
      13'h18C1: dout  = 8'b11111111; // 6337 : 255 - 0xff
      13'h18C2: dout  = 8'b11111111; // 6338 : 255 - 0xff
      13'h18C3: dout  = 8'b11111111; // 6339 : 255 - 0xff
      13'h18C4: dout  = 8'b11111111; // 6340 : 255 - 0xff
      13'h18C5: dout  = 8'b00000000; // 6341 :   0 - 0x0
      13'h18C6: dout  = 8'b11111111; // 6342 : 255 - 0xff
      13'h18C7: dout  = 8'b11111111; // 6343 : 255 - 0xff
      13'h18C8: dout  = 8'b00000000; // 6344 :   0 - 0x0
      13'h18C9: dout  = 8'b00000000; // 6345 :   0 - 0x0
      13'h18CA: dout  = 8'b00000000; // 6346 :   0 - 0x0
      13'h18CB: dout  = 8'b00000000; // 6347 :   0 - 0x0
      13'h18CC: dout  = 8'b00000000; // 6348 :   0 - 0x0
      13'h18CD: dout  = 8'b11111111; // 6349 : 255 - 0xff
      13'h18CE: dout  = 8'b00000000; // 6350 :   0 - 0x0
      13'h18CF: dout  = 8'b00000000; // 6351 :   0 - 0x0
      13'h18D0: dout  = 8'b11111100; // 6352 : 252 - 0xfc -- Background 0x8d
      13'h18D1: dout  = 8'b11111100; // 6353 : 252 - 0xfc
      13'h18D2: dout  = 8'b11111110; // 6354 : 254 - 0xfe
      13'h18D3: dout  = 8'b11111110; // 6355 : 254 - 0xfe
      13'h18D4: dout  = 8'b11111110; // 6356 : 254 - 0xfe
      13'h18D5: dout  = 8'b00000010; // 6357 :   2 - 0x2
      13'h18D6: dout  = 8'b11111110; // 6358 : 254 - 0xfe
      13'h18D7: dout  = 8'b11111110; // 6359 : 254 - 0xfe
      13'h18D8: dout  = 8'b00000111; // 6360 :   7 - 0x7
      13'h18D9: dout  = 8'b00000111; // 6361 :   7 - 0x7
      13'h18DA: dout  = 8'b00000011; // 6362 :   3 - 0x3
      13'h18DB: dout  = 8'b00000011; // 6363 :   3 - 0x3
      13'h18DC: dout  = 8'b00000011; // 6364 :   3 - 0x3
      13'h18DD: dout  = 8'b11111111; // 6365 : 255 - 0xff
      13'h18DE: dout  = 8'b00000011; // 6366 :   3 - 0x3
      13'h18DF: dout  = 8'b00000011; // 6367 :   3 - 0x3
      13'h18E0: dout  = 8'b11111111; // 6368 : 255 - 0xff -- Background 0x8e
      13'h18E1: dout  = 8'b10000000; // 6369 : 128 - 0x80
      13'h18E2: dout  = 8'b10000000; // 6370 : 128 - 0x80
      13'h18E3: dout  = 8'b10000000; // 6371 : 128 - 0x80
      13'h18E4: dout  = 8'b10000000; // 6372 : 128 - 0x80
      13'h18E5: dout  = 8'b10000000; // 6373 : 128 - 0x80
      13'h18E6: dout  = 8'b10000000; // 6374 : 128 - 0x80
      13'h18E7: dout  = 8'b10000000; // 6375 : 128 - 0x80
      13'h18E8: dout  = 8'b10000000; // 6376 : 128 - 0x80
      13'h18E9: dout  = 8'b11111111; // 6377 : 255 - 0xff
      13'h18EA: dout  = 8'b11111111; // 6378 : 255 - 0xff
      13'h18EB: dout  = 8'b11111111; // 6379 : 255 - 0xff
      13'h18EC: dout  = 8'b11111111; // 6380 : 255 - 0xff
      13'h18ED: dout  = 8'b11111111; // 6381 : 255 - 0xff
      13'h18EE: dout  = 8'b11111111; // 6382 : 255 - 0xff
      13'h18EF: dout  = 8'b11111111; // 6383 : 255 - 0xff
      13'h18F0: dout  = 8'b11111111; // 6384 : 255 - 0xff -- Background 0x8f
      13'h18F1: dout  = 8'b00000011; // 6385 :   3 - 0x3
      13'h18F2: dout  = 8'b00000011; // 6386 :   3 - 0x3
      13'h18F3: dout  = 8'b00000011; // 6387 :   3 - 0x3
      13'h18F4: dout  = 8'b00000011; // 6388 :   3 - 0x3
      13'h18F5: dout  = 8'b00000011; // 6389 :   3 - 0x3
      13'h18F6: dout  = 8'b00000011; // 6390 :   3 - 0x3
      13'h18F7: dout  = 8'b00000011; // 6391 :   3 - 0x3
      13'h18F8: dout  = 8'b00000011; // 6392 :   3 - 0x3
      13'h18F9: dout  = 8'b11111111; // 6393 : 255 - 0xff
      13'h18FA: dout  = 8'b11111111; // 6394 : 255 - 0xff
      13'h18FB: dout  = 8'b11111111; // 6395 : 255 - 0xff
      13'h18FC: dout  = 8'b11111111; // 6396 : 255 - 0xff
      13'h18FD: dout  = 8'b11111111; // 6397 : 255 - 0xff
      13'h18FE: dout  = 8'b11111111; // 6398 : 255 - 0xff
      13'h18FF: dout  = 8'b11111111; // 6399 : 255 - 0xff
      13'h1900: dout  = 8'b00000010; // 6400 :   2 - 0x2 -- Background 0x90
      13'h1901: dout  = 8'b00000010; // 6401 :   2 - 0x2
      13'h1902: dout  = 8'b00000010; // 6402 :   2 - 0x2
      13'h1903: dout  = 8'b00000010; // 6403 :   2 - 0x2
      13'h1904: dout  = 8'b00000010; // 6404 :   2 - 0x2
      13'h1905: dout  = 8'b00000010; // 6405 :   2 - 0x2
      13'h1906: dout  = 8'b00000100; // 6406 :   4 - 0x4
      13'h1907: dout  = 8'b00000100; // 6407 :   4 - 0x4
      13'h1908: dout  = 8'b11111111; // 6408 : 255 - 0xff
      13'h1909: dout  = 8'b11111111; // 6409 : 255 - 0xff
      13'h190A: dout  = 8'b11111111; // 6410 : 255 - 0xff
      13'h190B: dout  = 8'b11111111; // 6411 : 255 - 0xff
      13'h190C: dout  = 8'b11111111; // 6412 : 255 - 0xff
      13'h190D: dout  = 8'b11111111; // 6413 : 255 - 0xff
      13'h190E: dout  = 8'b11111111; // 6414 : 255 - 0xff
      13'h190F: dout  = 8'b11111111; // 6415 : 255 - 0xff
      13'h1910: dout  = 8'b10000000; // 6416 : 128 - 0x80 -- Background 0x91
      13'h1911: dout  = 8'b10000000; // 6417 : 128 - 0x80
      13'h1912: dout  = 8'b10101010; // 6418 : 170 - 0xaa
      13'h1913: dout  = 8'b11010101; // 6419 : 213 - 0xd5
      13'h1914: dout  = 8'b10101010; // 6420 : 170 - 0xaa
      13'h1915: dout  = 8'b11111111; // 6421 : 255 - 0xff
      13'h1916: dout  = 8'b11111111; // 6422 : 255 - 0xff
      13'h1917: dout  = 8'b11111111; // 6423 : 255 - 0xff
      13'h1918: dout  = 8'b11111111; // 6424 : 255 - 0xff
      13'h1919: dout  = 8'b11111111; // 6425 : 255 - 0xff
      13'h191A: dout  = 8'b11010101; // 6426 : 213 - 0xd5
      13'h191B: dout  = 8'b10101010; // 6427 : 170 - 0xaa
      13'h191C: dout  = 8'b11010101; // 6428 : 213 - 0xd5
      13'h191D: dout  = 8'b10000000; // 6429 : 128 - 0x80
      13'h191E: dout  = 8'b10000000; // 6430 : 128 - 0x80
      13'h191F: dout  = 8'b11111111; // 6431 : 255 - 0xff
      13'h1920: dout  = 8'b00000011; // 6432 :   3 - 0x3 -- Background 0x92
      13'h1921: dout  = 8'b00000011; // 6433 :   3 - 0x3
      13'h1922: dout  = 8'b10101011; // 6434 : 171 - 0xab
      13'h1923: dout  = 8'b01010111; // 6435 :  87 - 0x57
      13'h1924: dout  = 8'b10101011; // 6436 : 171 - 0xab
      13'h1925: dout  = 8'b11111111; // 6437 : 255 - 0xff
      13'h1926: dout  = 8'b11111111; // 6438 : 255 - 0xff
      13'h1927: dout  = 8'b11111110; // 6439 : 254 - 0xfe
      13'h1928: dout  = 8'b11111111; // 6440 : 255 - 0xff
      13'h1929: dout  = 8'b11111111; // 6441 : 255 - 0xff
      13'h192A: dout  = 8'b01010111; // 6442 :  87 - 0x57
      13'h192B: dout  = 8'b10101011; // 6443 : 171 - 0xab
      13'h192C: dout  = 8'b01010111; // 6444 :  87 - 0x57
      13'h192D: dout  = 8'b00000011; // 6445 :   3 - 0x3
      13'h192E: dout  = 8'b00000011; // 6446 :   3 - 0x3
      13'h192F: dout  = 8'b11111110; // 6447 : 254 - 0xfe
      13'h1930: dout  = 8'b00000000; // 6448 :   0 - 0x0 -- Background 0x93
      13'h1931: dout  = 8'b01010101; // 6449 :  85 - 0x55
      13'h1932: dout  = 8'b10101010; // 6450 : 170 - 0xaa
      13'h1933: dout  = 8'b01010101; // 6451 :  85 - 0x55
      13'h1934: dout  = 8'b11111111; // 6452 : 255 - 0xff
      13'h1935: dout  = 8'b11111111; // 6453 : 255 - 0xff
      13'h1936: dout  = 8'b11111111; // 6454 : 255 - 0xff
      13'h1937: dout  = 8'b00000000; // 6455 :   0 - 0x0
      13'h1938: dout  = 8'b11111111; // 6456 : 255 - 0xff
      13'h1939: dout  = 8'b10101010; // 6457 : 170 - 0xaa
      13'h193A: dout  = 8'b01010101; // 6458 :  85 - 0x55
      13'h193B: dout  = 8'b10101010; // 6459 : 170 - 0xaa
      13'h193C: dout  = 8'b00000000; // 6460 :   0 - 0x0
      13'h193D: dout  = 8'b00000000; // 6461 :   0 - 0x0
      13'h193E: dout  = 8'b11111111; // 6462 : 255 - 0xff
      13'h193F: dout  = 8'b00000000; // 6463 :   0 - 0x0
      13'h1940: dout  = 8'b00000100; // 6464 :   4 - 0x4 -- Background 0x94
      13'h1941: dout  = 8'b01010100; // 6465 :  84 - 0x54
      13'h1942: dout  = 8'b10101100; // 6466 : 172 - 0xac
      13'h1943: dout  = 8'b01011100; // 6467 :  92 - 0x5c
      13'h1944: dout  = 8'b11111100; // 6468 : 252 - 0xfc
      13'h1945: dout  = 8'b11111100; // 6469 : 252 - 0xfc
      13'h1946: dout  = 8'b11111100; // 6470 : 252 - 0xfc
      13'h1947: dout  = 8'b00111100; // 6471 :  60 - 0x3c
      13'h1948: dout  = 8'b11111111; // 6472 : 255 - 0xff
      13'h1949: dout  = 8'b10101111; // 6473 : 175 - 0xaf
      13'h194A: dout  = 8'b01010111; // 6474 :  87 - 0x57
      13'h194B: dout  = 8'b10101011; // 6475 : 171 - 0xab
      13'h194C: dout  = 8'b00001011; // 6476 :  11 - 0xb
      13'h194D: dout  = 8'b00001011; // 6477 :  11 - 0xb
      13'h194E: dout  = 8'b11110011; // 6478 : 243 - 0xf3
      13'h194F: dout  = 8'b00100011; // 6479 :  35 - 0x23
      13'h1950: dout  = 8'b00111111; // 6480 :  63 - 0x3f -- Background 0x95
      13'h1951: dout  = 8'b00111111; // 6481 :  63 - 0x3f
      13'h1952: dout  = 8'b00111111; // 6482 :  63 - 0x3f
      13'h1953: dout  = 8'b00111111; // 6483 :  63 - 0x3f
      13'h1954: dout  = 8'b00000000; // 6484 :   0 - 0x0
      13'h1955: dout  = 8'b00000000; // 6485 :   0 - 0x0
      13'h1956: dout  = 8'b00000000; // 6486 :   0 - 0x0
      13'h1957: dout  = 8'b11111111; // 6487 : 255 - 0xff
      13'h1958: dout  = 8'b11111111; // 6488 : 255 - 0xff
      13'h1959: dout  = 8'b11111111; // 6489 : 255 - 0xff
      13'h195A: dout  = 8'b11111111; // 6490 : 255 - 0xff
      13'h195B: dout  = 8'b11111111; // 6491 : 255 - 0xff
      13'h195C: dout  = 8'b11111111; // 6492 : 255 - 0xff
      13'h195D: dout  = 8'b11111111; // 6493 : 255 - 0xff
      13'h195E: dout  = 8'b11111111; // 6494 : 255 - 0xff
      13'h195F: dout  = 8'b11111111; // 6495 : 255 - 0xff
      13'h1960: dout  = 8'b01111110; // 6496 : 126 - 0x7e -- Background 0x96
      13'h1961: dout  = 8'b01111100; // 6497 : 124 - 0x7c
      13'h1962: dout  = 8'b01111100; // 6498 : 124 - 0x7c
      13'h1963: dout  = 8'b01111000; // 6499 : 120 - 0x78
      13'h1964: dout  = 8'b00000000; // 6500 :   0 - 0x0
      13'h1965: dout  = 8'b00000000; // 6501 :   0 - 0x0
      13'h1966: dout  = 8'b00000000; // 6502 :   0 - 0x0
      13'h1967: dout  = 8'b11111111; // 6503 : 255 - 0xff
      13'h1968: dout  = 8'b11111111; // 6504 : 255 - 0xff
      13'h1969: dout  = 8'b11111111; // 6505 : 255 - 0xff
      13'h196A: dout  = 8'b11111111; // 6506 : 255 - 0xff
      13'h196B: dout  = 8'b11111111; // 6507 : 255 - 0xff
      13'h196C: dout  = 8'b11111111; // 6508 : 255 - 0xff
      13'h196D: dout  = 8'b11111111; // 6509 : 255 - 0xff
      13'h196E: dout  = 8'b11111111; // 6510 : 255 - 0xff
      13'h196F: dout  = 8'b11111111; // 6511 : 255 - 0xff
      13'h1970: dout  = 8'b00011111; // 6512 :  31 - 0x1f -- Background 0x97
      13'h1971: dout  = 8'b00001111; // 6513 :  15 - 0xf
      13'h1972: dout  = 8'b00001111; // 6514 :  15 - 0xf
      13'h1973: dout  = 8'b00000111; // 6515 :   7 - 0x7
      13'h1974: dout  = 8'b00000000; // 6516 :   0 - 0x0
      13'h1975: dout  = 8'b00000000; // 6517 :   0 - 0x0
      13'h1976: dout  = 8'b00000000; // 6518 :   0 - 0x0
      13'h1977: dout  = 8'b11111111; // 6519 : 255 - 0xff
      13'h1978: dout  = 8'b11111111; // 6520 : 255 - 0xff
      13'h1979: dout  = 8'b11111111; // 6521 : 255 - 0xff
      13'h197A: dout  = 8'b11111111; // 6522 : 255 - 0xff
      13'h197B: dout  = 8'b11111111; // 6523 : 255 - 0xff
      13'h197C: dout  = 8'b11111111; // 6524 : 255 - 0xff
      13'h197D: dout  = 8'b11111111; // 6525 : 255 - 0xff
      13'h197E: dout  = 8'b11111111; // 6526 : 255 - 0xff
      13'h197F: dout  = 8'b11111111; // 6527 : 255 - 0xff
      13'h1980: dout  = 8'b11111110; // 6528 : 254 - 0xfe -- Background 0x98
      13'h1981: dout  = 8'b11111100; // 6529 : 252 - 0xfc
      13'h1982: dout  = 8'b11111100; // 6530 : 252 - 0xfc
      13'h1983: dout  = 8'b11111000; // 6531 : 248 - 0xf8
      13'h1984: dout  = 8'b00000000; // 6532 :   0 - 0x0
      13'h1985: dout  = 8'b00000000; // 6533 :   0 - 0x0
      13'h1986: dout  = 8'b00000000; // 6534 :   0 - 0x0
      13'h1987: dout  = 8'b11111111; // 6535 : 255 - 0xff
      13'h1988: dout  = 8'b11111111; // 6536 : 255 - 0xff
      13'h1989: dout  = 8'b11111111; // 6537 : 255 - 0xff
      13'h198A: dout  = 8'b11111111; // 6538 : 255 - 0xff
      13'h198B: dout  = 8'b11111111; // 6539 : 255 - 0xff
      13'h198C: dout  = 8'b11111111; // 6540 : 255 - 0xff
      13'h198D: dout  = 8'b11111111; // 6541 : 255 - 0xff
      13'h198E: dout  = 8'b11111111; // 6542 : 255 - 0xff
      13'h198F: dout  = 8'b11111111; // 6543 : 255 - 0xff
      13'h1990: dout  = 8'b00000000; // 6544 :   0 - 0x0 -- Background 0x99
      13'h1991: dout  = 8'b00000000; // 6545 :   0 - 0x0
      13'h1992: dout  = 8'b00000000; // 6546 :   0 - 0x0
      13'h1993: dout  = 8'b00000000; // 6547 :   0 - 0x0
      13'h1994: dout  = 8'b11111111; // 6548 : 255 - 0xff
      13'h1995: dout  = 8'b11111111; // 6549 : 255 - 0xff
      13'h1996: dout  = 8'b00000000; // 6550 :   0 - 0x0
      13'h1997: dout  = 8'b00000000; // 6551 :   0 - 0x0
      13'h1998: dout  = 8'b00000000; // 6552 :   0 - 0x0
      13'h1999: dout  = 8'b00000000; // 6553 :   0 - 0x0
      13'h199A: dout  = 8'b00000000; // 6554 :   0 - 0x0
      13'h199B: dout  = 8'b00000000; // 6555 :   0 - 0x0
      13'h199C: dout  = 8'b00000000; // 6556 :   0 - 0x0
      13'h199D: dout  = 8'b00000000; // 6557 :   0 - 0x0
      13'h199E: dout  = 8'b00000000; // 6558 :   0 - 0x0
      13'h199F: dout  = 8'b00000000; // 6559 :   0 - 0x0
      13'h19A0: dout  = 8'b00011000; // 6560 :  24 - 0x18 -- Background 0x9a
      13'h19A1: dout  = 8'b00011000; // 6561 :  24 - 0x18
      13'h19A2: dout  = 8'b00011000; // 6562 :  24 - 0x18
      13'h19A3: dout  = 8'b00011000; // 6563 :  24 - 0x18
      13'h19A4: dout  = 8'b00011000; // 6564 :  24 - 0x18
      13'h19A5: dout  = 8'b00011000; // 6565 :  24 - 0x18
      13'h19A6: dout  = 8'b00011000; // 6566 :  24 - 0x18
      13'h19A7: dout  = 8'b00011000; // 6567 :  24 - 0x18
      13'h19A8: dout  = 8'b00000000; // 6568 :   0 - 0x0
      13'h19A9: dout  = 8'b00000000; // 6569 :   0 - 0x0
      13'h19AA: dout  = 8'b00000000; // 6570 :   0 - 0x0
      13'h19AB: dout  = 8'b00000000; // 6571 :   0 - 0x0
      13'h19AC: dout  = 8'b00000000; // 6572 :   0 - 0x0
      13'h19AD: dout  = 8'b00000000; // 6573 :   0 - 0x0
      13'h19AE: dout  = 8'b00000000; // 6574 :   0 - 0x0
      13'h19AF: dout  = 8'b00000000; // 6575 :   0 - 0x0
      13'h19B0: dout  = 8'b00000111; // 6576 :   7 - 0x7 -- Background 0x9b
      13'h19B1: dout  = 8'b00011111; // 6577 :  31 - 0x1f
      13'h19B2: dout  = 8'b00111111; // 6578 :  63 - 0x3f
      13'h19B3: dout  = 8'b11111111; // 6579 : 255 - 0xff
      13'h19B4: dout  = 8'b01111111; // 6580 : 127 - 0x7f
      13'h19B5: dout  = 8'b01111111; // 6581 : 127 - 0x7f
      13'h19B6: dout  = 8'b11111111; // 6582 : 255 - 0xff
      13'h19B7: dout  = 8'b11111111; // 6583 : 255 - 0xff
      13'h19B8: dout  = 8'b11111111; // 6584 : 255 - 0xff
      13'h19B9: dout  = 8'b11111111; // 6585 : 255 - 0xff
      13'h19BA: dout  = 8'b11111111; // 6586 : 255 - 0xff
      13'h19BB: dout  = 8'b11111111; // 6587 : 255 - 0xff
      13'h19BC: dout  = 8'b11111111; // 6588 : 255 - 0xff
      13'h19BD: dout  = 8'b11111111; // 6589 : 255 - 0xff
      13'h19BE: dout  = 8'b11111111; // 6590 : 255 - 0xff
      13'h19BF: dout  = 8'b11111111; // 6591 : 255 - 0xff
      13'h19C0: dout  = 8'b11100001; // 6592 : 225 - 0xe1 -- Background 0x9c
      13'h19C1: dout  = 8'b11111001; // 6593 : 249 - 0xf9
      13'h19C2: dout  = 8'b11111101; // 6594 : 253 - 0xfd
      13'h19C3: dout  = 8'b11111111; // 6595 : 255 - 0xff
      13'h19C4: dout  = 8'b11111110; // 6596 : 254 - 0xfe
      13'h19C5: dout  = 8'b11111110; // 6597 : 254 - 0xfe
      13'h19C6: dout  = 8'b11111111; // 6598 : 255 - 0xff
      13'h19C7: dout  = 8'b11111111; // 6599 : 255 - 0xff
      13'h19C8: dout  = 8'b11111111; // 6600 : 255 - 0xff
      13'h19C9: dout  = 8'b11111111; // 6601 : 255 - 0xff
      13'h19CA: dout  = 8'b11111111; // 6602 : 255 - 0xff
      13'h19CB: dout  = 8'b11111111; // 6603 : 255 - 0xff
      13'h19CC: dout  = 8'b11111111; // 6604 : 255 - 0xff
      13'h19CD: dout  = 8'b11111111; // 6605 : 255 - 0xff
      13'h19CE: dout  = 8'b11111111; // 6606 : 255 - 0xff
      13'h19CF: dout  = 8'b11111111; // 6607 : 255 - 0xff
      13'h19D0: dout  = 8'b11110000; // 6608 : 240 - 0xf0 -- Background 0x9d
      13'h19D1: dout  = 8'b00010000; // 6609 :  16 - 0x10
      13'h19D2: dout  = 8'b00010000; // 6610 :  16 - 0x10
      13'h19D3: dout  = 8'b00010000; // 6611 :  16 - 0x10
      13'h19D4: dout  = 8'b00010000; // 6612 :  16 - 0x10
      13'h19D5: dout  = 8'b00010000; // 6613 :  16 - 0x10
      13'h19D6: dout  = 8'b00010000; // 6614 :  16 - 0x10
      13'h19D7: dout  = 8'b11111111; // 6615 : 255 - 0xff
      13'h19D8: dout  = 8'b00000000; // 6616 :   0 - 0x0
      13'h19D9: dout  = 8'b11100000; // 6617 : 224 - 0xe0
      13'h19DA: dout  = 8'b11100000; // 6618 : 224 - 0xe0
      13'h19DB: dout  = 8'b11100000; // 6619 : 224 - 0xe0
      13'h19DC: dout  = 8'b11100000; // 6620 : 224 - 0xe0
      13'h19DD: dout  = 8'b11100000; // 6621 : 224 - 0xe0
      13'h19DE: dout  = 8'b11100000; // 6622 : 224 - 0xe0
      13'h19DF: dout  = 8'b11100000; // 6623 : 224 - 0xe0
      13'h19E0: dout  = 8'b00011111; // 6624 :  31 - 0x1f -- Background 0x9e
      13'h19E1: dout  = 8'b00010000; // 6625 :  16 - 0x10
      13'h19E2: dout  = 8'b00010000; // 6626 :  16 - 0x10
      13'h19E3: dout  = 8'b00010000; // 6627 :  16 - 0x10
      13'h19E4: dout  = 8'b00010000; // 6628 :  16 - 0x10
      13'h19E5: dout  = 8'b00010000; // 6629 :  16 - 0x10
      13'h19E6: dout  = 8'b00010000; // 6630 :  16 - 0x10
      13'h19E7: dout  = 8'b11111111; // 6631 : 255 - 0xff
      13'h19E8: dout  = 8'b00000000; // 6632 :   0 - 0x0
      13'h19E9: dout  = 8'b00001111; // 6633 :  15 - 0xf
      13'h19EA: dout  = 8'b00001111; // 6634 :  15 - 0xf
      13'h19EB: dout  = 8'b00001111; // 6635 :  15 - 0xf
      13'h19EC: dout  = 8'b00001111; // 6636 :  15 - 0xf
      13'h19ED: dout  = 8'b00001111; // 6637 :  15 - 0xf
      13'h19EE: dout  = 8'b00001111; // 6638 :  15 - 0xf
      13'h19EF: dout  = 8'b00001111; // 6639 :  15 - 0xf
      13'h19F0: dout  = 8'b10010010; // 6640 : 146 - 0x92 -- Background 0x9f
      13'h19F1: dout  = 8'b10010010; // 6641 : 146 - 0x92
      13'h19F2: dout  = 8'b10010010; // 6642 : 146 - 0x92
      13'h19F3: dout  = 8'b11111110; // 6643 : 254 - 0xfe
      13'h19F4: dout  = 8'b11111110; // 6644 : 254 - 0xfe
      13'h19F5: dout  = 8'b00000000; // 6645 :   0 - 0x0
      13'h19F6: dout  = 8'b00000000; // 6646 :   0 - 0x0
      13'h19F7: dout  = 8'b00000000; // 6647 :   0 - 0x0
      13'h19F8: dout  = 8'b01001000; // 6648 :  72 - 0x48
      13'h19F9: dout  = 8'b01001000; // 6649 :  72 - 0x48
      13'h19FA: dout  = 8'b01101100; // 6650 : 108 - 0x6c
      13'h19FB: dout  = 8'b00000000; // 6651 :   0 - 0x0
      13'h19FC: dout  = 8'b00000000; // 6652 :   0 - 0x0
      13'h19FD: dout  = 8'b00000000; // 6653 :   0 - 0x0
      13'h19FE: dout  = 8'b11111110; // 6654 : 254 - 0xfe
      13'h19FF: dout  = 8'b00000000; // 6655 :   0 - 0x0
      13'h1A00: dout  = 8'b00001010; // 6656 :  10 - 0xa -- Background 0xa0
      13'h1A01: dout  = 8'b00001010; // 6657 :  10 - 0xa
      13'h1A02: dout  = 8'b00111010; // 6658 :  58 - 0x3a
      13'h1A03: dout  = 8'b00001010; // 6659 :  10 - 0xa
      13'h1A04: dout  = 8'b11111011; // 6660 : 251 - 0xfb
      13'h1A05: dout  = 8'b00001011; // 6661 :  11 - 0xb
      13'h1A06: dout  = 8'b00001011; // 6662 :  11 - 0xb
      13'h1A07: dout  = 8'b00001011; // 6663 :  11 - 0xb
      13'h1A08: dout  = 8'b00000101; // 6664 :   5 - 0x5
      13'h1A09: dout  = 8'b00000101; // 6665 :   5 - 0x5
      13'h1A0A: dout  = 8'b11000101; // 6666 : 197 - 0xc5
      13'h1A0B: dout  = 8'b11110101; // 6667 : 245 - 0xf5
      13'h1A0C: dout  = 8'b11110100; // 6668 : 244 - 0xf4
      13'h1A0D: dout  = 8'b00000100; // 6669 :   4 - 0x4
      13'h1A0E: dout  = 8'b00000100; // 6670 :   4 - 0x4
      13'h1A0F: dout  = 8'b00000100; // 6671 :   4 - 0x4
      13'h1A10: dout  = 8'b10010000; // 6672 : 144 - 0x90 -- Background 0xa1
      13'h1A11: dout  = 8'b10010000; // 6673 : 144 - 0x90
      13'h1A12: dout  = 8'b10011111; // 6674 : 159 - 0x9f
      13'h1A13: dout  = 8'b10010000; // 6675 : 144 - 0x90
      13'h1A14: dout  = 8'b10011111; // 6676 : 159 - 0x9f
      13'h1A15: dout  = 8'b10010000; // 6677 : 144 - 0x90
      13'h1A16: dout  = 8'b10010000; // 6678 : 144 - 0x90
      13'h1A17: dout  = 8'b10010000; // 6679 : 144 - 0x90
      13'h1A18: dout  = 8'b01110000; // 6680 : 112 - 0x70
      13'h1A19: dout  = 8'b01110000; // 6681 : 112 - 0x70
      13'h1A1A: dout  = 8'b01110000; // 6682 : 112 - 0x70
      13'h1A1B: dout  = 8'b01111111; // 6683 : 127 - 0x7f
      13'h1A1C: dout  = 8'b01111111; // 6684 : 127 - 0x7f
      13'h1A1D: dout  = 8'b01110000; // 6685 : 112 - 0x70
      13'h1A1E: dout  = 8'b01110000; // 6686 : 112 - 0x70
      13'h1A1F: dout  = 8'b01110000; // 6687 : 112 - 0x70
      13'h1A20: dout  = 8'b00000001; // 6688 :   1 - 0x1 -- Background 0xa2
      13'h1A21: dout  = 8'b00000001; // 6689 :   1 - 0x1
      13'h1A22: dout  = 8'b00000001; // 6690 :   1 - 0x1
      13'h1A23: dout  = 8'b00000001; // 6691 :   1 - 0x1
      13'h1A24: dout  = 8'b00000001; // 6692 :   1 - 0x1
      13'h1A25: dout  = 8'b00000001; // 6693 :   1 - 0x1
      13'h1A26: dout  = 8'b00000001; // 6694 :   1 - 0x1
      13'h1A27: dout  = 8'b00000001; // 6695 :   1 - 0x1
      13'h1A28: dout  = 8'b00000000; // 6696 :   0 - 0x0
      13'h1A29: dout  = 8'b00000000; // 6697 :   0 - 0x0
      13'h1A2A: dout  = 8'b00000000; // 6698 :   0 - 0x0
      13'h1A2B: dout  = 8'b00000000; // 6699 :   0 - 0x0
      13'h1A2C: dout  = 8'b00000000; // 6700 :   0 - 0x0
      13'h1A2D: dout  = 8'b00000000; // 6701 :   0 - 0x0
      13'h1A2E: dout  = 8'b00000000; // 6702 :   0 - 0x0
      13'h1A2F: dout  = 8'b00000000; // 6703 :   0 - 0x0
      13'h1A30: dout  = 8'b10000000; // 6704 : 128 - 0x80 -- Background 0xa3
      13'h1A31: dout  = 8'b10000000; // 6705 : 128 - 0x80
      13'h1A32: dout  = 8'b10000000; // 6706 : 128 - 0x80
      13'h1A33: dout  = 8'b10000000; // 6707 : 128 - 0x80
      13'h1A34: dout  = 8'b10000000; // 6708 : 128 - 0x80
      13'h1A35: dout  = 8'b10000000; // 6709 : 128 - 0x80
      13'h1A36: dout  = 8'b10000000; // 6710 : 128 - 0x80
      13'h1A37: dout  = 8'b10000000; // 6711 : 128 - 0x80
      13'h1A38: dout  = 8'b00000000; // 6712 :   0 - 0x0
      13'h1A39: dout  = 8'b00000000; // 6713 :   0 - 0x0
      13'h1A3A: dout  = 8'b00000000; // 6714 :   0 - 0x0
      13'h1A3B: dout  = 8'b00000000; // 6715 :   0 - 0x0
      13'h1A3C: dout  = 8'b00000000; // 6716 :   0 - 0x0
      13'h1A3D: dout  = 8'b00000000; // 6717 :   0 - 0x0
      13'h1A3E: dout  = 8'b00000000; // 6718 :   0 - 0x0
      13'h1A3F: dout  = 8'b00000000; // 6719 :   0 - 0x0
      13'h1A40: dout  = 8'b00001000; // 6720 :   8 - 0x8 -- Background 0xa4
      13'h1A41: dout  = 8'b10001000; // 6721 : 136 - 0x88
      13'h1A42: dout  = 8'b10010001; // 6722 : 145 - 0x91
      13'h1A43: dout  = 8'b11010001; // 6723 : 209 - 0xd1
      13'h1A44: dout  = 8'b01010011; // 6724 :  83 - 0x53
      13'h1A45: dout  = 8'b01010011; // 6725 :  83 - 0x53
      13'h1A46: dout  = 8'b01110011; // 6726 : 115 - 0x73
      13'h1A47: dout  = 8'b00111111; // 6727 :  63 - 0x3f
      13'h1A48: dout  = 8'b11111111; // 6728 : 255 - 0xff
      13'h1A49: dout  = 8'b11111111; // 6729 : 255 - 0xff
      13'h1A4A: dout  = 8'b11111111; // 6730 : 255 - 0xff
      13'h1A4B: dout  = 8'b11111111; // 6731 : 255 - 0xff
      13'h1A4C: dout  = 8'b11111111; // 6732 : 255 - 0xff
      13'h1A4D: dout  = 8'b11111110; // 6733 : 254 - 0xfe
      13'h1A4E: dout  = 8'b10111110; // 6734 : 190 - 0xbe
      13'h1A4F: dout  = 8'b11001110; // 6735 : 206 - 0xce
      13'h1A50: dout  = 8'b00000000; // 6736 :   0 - 0x0 -- Background 0xa5
      13'h1A51: dout  = 8'b00000000; // 6737 :   0 - 0x0
      13'h1A52: dout  = 8'b00000111; // 6738 :   7 - 0x7
      13'h1A53: dout  = 8'b00001111; // 6739 :  15 - 0xf
      13'h1A54: dout  = 8'b00001100; // 6740 :  12 - 0xc
      13'h1A55: dout  = 8'b00011011; // 6741 :  27 - 0x1b
      13'h1A56: dout  = 8'b00011011; // 6742 :  27 - 0x1b
      13'h1A57: dout  = 8'b00011011; // 6743 :  27 - 0x1b
      13'h1A58: dout  = 8'b00000000; // 6744 :   0 - 0x0
      13'h1A59: dout  = 8'b00000000; // 6745 :   0 - 0x0
      13'h1A5A: dout  = 8'b00000000; // 6746 :   0 - 0x0
      13'h1A5B: dout  = 8'b00000000; // 6747 :   0 - 0x0
      13'h1A5C: dout  = 8'b00000011; // 6748 :   3 - 0x3
      13'h1A5D: dout  = 8'b00000100; // 6749 :   4 - 0x4
      13'h1A5E: dout  = 8'b00000100; // 6750 :   4 - 0x4
      13'h1A5F: dout  = 8'b00000100; // 6751 :   4 - 0x4
      13'h1A60: dout  = 8'b00000000; // 6752 :   0 - 0x0 -- Background 0xa6
      13'h1A61: dout  = 8'b00000000; // 6753 :   0 - 0x0
      13'h1A62: dout  = 8'b11100000; // 6754 : 224 - 0xe0
      13'h1A63: dout  = 8'b11110000; // 6755 : 240 - 0xf0
      13'h1A64: dout  = 8'b11110000; // 6756 : 240 - 0xf0
      13'h1A65: dout  = 8'b11111000; // 6757 : 248 - 0xf8
      13'h1A66: dout  = 8'b11111000; // 6758 : 248 - 0xf8
      13'h1A67: dout  = 8'b11111000; // 6759 : 248 - 0xf8
      13'h1A68: dout  = 8'b00000000; // 6760 :   0 - 0x0
      13'h1A69: dout  = 8'b00000000; // 6761 :   0 - 0x0
      13'h1A6A: dout  = 8'b01100000; // 6762 :  96 - 0x60
      13'h1A6B: dout  = 8'b00110000; // 6763 :  48 - 0x30
      13'h1A6C: dout  = 8'b00110000; // 6764 :  48 - 0x30
      13'h1A6D: dout  = 8'b10011000; // 6765 : 152 - 0x98
      13'h1A6E: dout  = 8'b10011000; // 6766 : 152 - 0x98
      13'h1A6F: dout  = 8'b10011000; // 6767 : 152 - 0x98
      13'h1A70: dout  = 8'b00011011; // 6768 :  27 - 0x1b -- Background 0xa7
      13'h1A71: dout  = 8'b00011011; // 6769 :  27 - 0x1b
      13'h1A72: dout  = 8'b00011011; // 6770 :  27 - 0x1b
      13'h1A73: dout  = 8'b00011011; // 6771 :  27 - 0x1b
      13'h1A74: dout  = 8'b00011011; // 6772 :  27 - 0x1b
      13'h1A75: dout  = 8'b00001111; // 6773 :  15 - 0xf
      13'h1A76: dout  = 8'b00001111; // 6774 :  15 - 0xf
      13'h1A77: dout  = 8'b00000111; // 6775 :   7 - 0x7
      13'h1A78: dout  = 8'b00000100; // 6776 :   4 - 0x4
      13'h1A79: dout  = 8'b00000100; // 6777 :   4 - 0x4
      13'h1A7A: dout  = 8'b00000100; // 6778 :   4 - 0x4
      13'h1A7B: dout  = 8'b00000100; // 6779 :   4 - 0x4
      13'h1A7C: dout  = 8'b00000100; // 6780 :   4 - 0x4
      13'h1A7D: dout  = 8'b00000011; // 6781 :   3 - 0x3
      13'h1A7E: dout  = 8'b00000000; // 6782 :   0 - 0x0
      13'h1A7F: dout  = 8'b00000000; // 6783 :   0 - 0x0
      13'h1A80: dout  = 8'b11111000; // 6784 : 248 - 0xf8 -- Background 0xa8
      13'h1A81: dout  = 8'b11111000; // 6785 : 248 - 0xf8
      13'h1A82: dout  = 8'b11111000; // 6786 : 248 - 0xf8
      13'h1A83: dout  = 8'b11111000; // 6787 : 248 - 0xf8
      13'h1A84: dout  = 8'b11111000; // 6788 : 248 - 0xf8
      13'h1A85: dout  = 8'b11110000; // 6789 : 240 - 0xf0
      13'h1A86: dout  = 8'b11110000; // 6790 : 240 - 0xf0
      13'h1A87: dout  = 8'b11100000; // 6791 : 224 - 0xe0
      13'h1A88: dout  = 8'b10011000; // 6792 : 152 - 0x98
      13'h1A89: dout  = 8'b10011000; // 6793 : 152 - 0x98
      13'h1A8A: dout  = 8'b10011000; // 6794 : 152 - 0x98
      13'h1A8B: dout  = 8'b10011000; // 6795 : 152 - 0x98
      13'h1A8C: dout  = 8'b10011000; // 6796 : 152 - 0x98
      13'h1A8D: dout  = 8'b00110000; // 6797 :  48 - 0x30
      13'h1A8E: dout  = 8'b00110000; // 6798 :  48 - 0x30
      13'h1A8F: dout  = 8'b01100000; // 6799 :  96 - 0x60
      13'h1A90: dout  = 8'b11110001; // 6800 : 241 - 0xf1 -- Background 0xa9
      13'h1A91: dout  = 8'b00010001; // 6801 :  17 - 0x11
      13'h1A92: dout  = 8'b00010001; // 6802 :  17 - 0x11
      13'h1A93: dout  = 8'b00011111; // 6803 :  31 - 0x1f
      13'h1A94: dout  = 8'b00010000; // 6804 :  16 - 0x10
      13'h1A95: dout  = 8'b00010000; // 6805 :  16 - 0x10
      13'h1A96: dout  = 8'b00010000; // 6806 :  16 - 0x10
      13'h1A97: dout  = 8'b11111111; // 6807 : 255 - 0xff
      13'h1A98: dout  = 8'b00001111; // 6808 :  15 - 0xf
      13'h1A99: dout  = 8'b11101111; // 6809 : 239 - 0xef
      13'h1A9A: dout  = 8'b11101111; // 6810 : 239 - 0xef
      13'h1A9B: dout  = 8'b11101111; // 6811 : 239 - 0xef
      13'h1A9C: dout  = 8'b11101111; // 6812 : 239 - 0xef
      13'h1A9D: dout  = 8'b11101111; // 6813 : 239 - 0xef
      13'h1A9E: dout  = 8'b11101111; // 6814 : 239 - 0xef
      13'h1A9F: dout  = 8'b11100000; // 6815 : 224 - 0xe0
      13'h1AA0: dout  = 8'b00011111; // 6816 :  31 - 0x1f -- Background 0xaa
      13'h1AA1: dout  = 8'b00010000; // 6817 :  16 - 0x10
      13'h1AA2: dout  = 8'b00010000; // 6818 :  16 - 0x10
      13'h1AA3: dout  = 8'b11110000; // 6819 : 240 - 0xf0
      13'h1AA4: dout  = 8'b00010000; // 6820 :  16 - 0x10
      13'h1AA5: dout  = 8'b00010000; // 6821 :  16 - 0x10
      13'h1AA6: dout  = 8'b00010000; // 6822 :  16 - 0x10
      13'h1AA7: dout  = 8'b11111111; // 6823 : 255 - 0xff
      13'h1AA8: dout  = 8'b11100000; // 6824 : 224 - 0xe0
      13'h1AA9: dout  = 8'b11101111; // 6825 : 239 - 0xef
      13'h1AAA: dout  = 8'b11101111; // 6826 : 239 - 0xef
      13'h1AAB: dout  = 8'b11101111; // 6827 : 239 - 0xef
      13'h1AAC: dout  = 8'b11101111; // 6828 : 239 - 0xef
      13'h1AAD: dout  = 8'b11101111; // 6829 : 239 - 0xef
      13'h1AAE: dout  = 8'b11101111; // 6830 : 239 - 0xef
      13'h1AAF: dout  = 8'b00001111; // 6831 :  15 - 0xf
      13'h1AB0: dout  = 8'b01111111; // 6832 : 127 - 0x7f -- Background 0xab
      13'h1AB1: dout  = 8'b10111111; // 6833 : 191 - 0xbf
      13'h1AB2: dout  = 8'b11011111; // 6834 : 223 - 0xdf
      13'h1AB3: dout  = 8'b11101111; // 6835 : 239 - 0xef
      13'h1AB4: dout  = 8'b11110000; // 6836 : 240 - 0xf0
      13'h1AB5: dout  = 8'b11110000; // 6837 : 240 - 0xf0
      13'h1AB6: dout  = 8'b11110000; // 6838 : 240 - 0xf0
      13'h1AB7: dout  = 8'b11110000; // 6839 : 240 - 0xf0
      13'h1AB8: dout  = 8'b10000000; // 6840 : 128 - 0x80
      13'h1AB9: dout  = 8'b01000000; // 6841 :  64 - 0x40
      13'h1ABA: dout  = 8'b00100000; // 6842 :  32 - 0x20
      13'h1ABB: dout  = 8'b00010000; // 6843 :  16 - 0x10
      13'h1ABC: dout  = 8'b00001111; // 6844 :  15 - 0xf
      13'h1ABD: dout  = 8'b00001111; // 6845 :  15 - 0xf
      13'h1ABE: dout  = 8'b00001111; // 6846 :  15 - 0xf
      13'h1ABF: dout  = 8'b00001111; // 6847 :  15 - 0xf
      13'h1AC0: dout  = 8'b11110000; // 6848 : 240 - 0xf0 -- Background 0xac
      13'h1AC1: dout  = 8'b11110000; // 6849 : 240 - 0xf0
      13'h1AC2: dout  = 8'b11110000; // 6850 : 240 - 0xf0
      13'h1AC3: dout  = 8'b11110000; // 6851 : 240 - 0xf0
      13'h1AC4: dout  = 8'b11111111; // 6852 : 255 - 0xff
      13'h1AC5: dout  = 8'b11111111; // 6853 : 255 - 0xff
      13'h1AC6: dout  = 8'b11111111; // 6854 : 255 - 0xff
      13'h1AC7: dout  = 8'b11111111; // 6855 : 255 - 0xff
      13'h1AC8: dout  = 8'b00001111; // 6856 :  15 - 0xf
      13'h1AC9: dout  = 8'b00001111; // 6857 :  15 - 0xf
      13'h1ACA: dout  = 8'b00001111; // 6858 :  15 - 0xf
      13'h1ACB: dout  = 8'b00001111; // 6859 :  15 - 0xf
      13'h1ACC: dout  = 8'b00011111; // 6860 :  31 - 0x1f
      13'h1ACD: dout  = 8'b00111111; // 6861 :  63 - 0x3f
      13'h1ACE: dout  = 8'b01111111; // 6862 : 127 - 0x7f
      13'h1ACF: dout  = 8'b11111111; // 6863 : 255 - 0xff
      13'h1AD0: dout  = 8'b11111111; // 6864 : 255 - 0xff -- Background 0xad
      13'h1AD1: dout  = 8'b11111111; // 6865 : 255 - 0xff
      13'h1AD2: dout  = 8'b11111111; // 6866 : 255 - 0xff
      13'h1AD3: dout  = 8'b11111111; // 6867 : 255 - 0xff
      13'h1AD4: dout  = 8'b00001111; // 6868 :  15 - 0xf
      13'h1AD5: dout  = 8'b00001111; // 6869 :  15 - 0xf
      13'h1AD6: dout  = 8'b00001111; // 6870 :  15 - 0xf
      13'h1AD7: dout  = 8'b00001111; // 6871 :  15 - 0xf
      13'h1AD8: dout  = 8'b00000001; // 6872 :   1 - 0x1
      13'h1AD9: dout  = 8'b00000011; // 6873 :   3 - 0x3
      13'h1ADA: dout  = 8'b00000111; // 6874 :   7 - 0x7
      13'h1ADB: dout  = 8'b00001111; // 6875 :  15 - 0xf
      13'h1ADC: dout  = 8'b11111111; // 6876 : 255 - 0xff
      13'h1ADD: dout  = 8'b11111111; // 6877 : 255 - 0xff
      13'h1ADE: dout  = 8'b11111111; // 6878 : 255 - 0xff
      13'h1ADF: dout  = 8'b11111111; // 6879 : 255 - 0xff
      13'h1AE0: dout  = 8'b00001111; // 6880 :  15 - 0xf -- Background 0xae
      13'h1AE1: dout  = 8'b00001111; // 6881 :  15 - 0xf
      13'h1AE2: dout  = 8'b00001111; // 6882 :  15 - 0xf
      13'h1AE3: dout  = 8'b00001111; // 6883 :  15 - 0xf
      13'h1AE4: dout  = 8'b11110111; // 6884 : 247 - 0xf7
      13'h1AE5: dout  = 8'b11111011; // 6885 : 251 - 0xfb
      13'h1AE6: dout  = 8'b11111101; // 6886 : 253 - 0xfd
      13'h1AE7: dout  = 8'b11111110; // 6887 : 254 - 0xfe
      13'h1AE8: dout  = 8'b11111111; // 6888 : 255 - 0xff
      13'h1AE9: dout  = 8'b11111111; // 6889 : 255 - 0xff
      13'h1AEA: dout  = 8'b11111111; // 6890 : 255 - 0xff
      13'h1AEB: dout  = 8'b11111111; // 6891 : 255 - 0xff
      13'h1AEC: dout  = 8'b11111111; // 6892 : 255 - 0xff
      13'h1AED: dout  = 8'b11111111; // 6893 : 255 - 0xff
      13'h1AEE: dout  = 8'b11111111; // 6894 : 255 - 0xff
      13'h1AEF: dout  = 8'b11111111; // 6895 : 255 - 0xff
      13'h1AF0: dout  = 8'b00000000; // 6896 :   0 - 0x0 -- Background 0xaf
      13'h1AF1: dout  = 8'b00000000; // 6897 :   0 - 0x0
      13'h1AF2: dout  = 8'b00000000; // 6898 :   0 - 0x0
      13'h1AF3: dout  = 8'b00000000; // 6899 :   0 - 0x0
      13'h1AF4: dout  = 8'b00000000; // 6900 :   0 - 0x0
      13'h1AF5: dout  = 8'b00000000; // 6901 :   0 - 0x0
      13'h1AF6: dout  = 8'b00011000; // 6902 :  24 - 0x18
      13'h1AF7: dout  = 8'b00011000; // 6903 :  24 - 0x18
      13'h1AF8: dout  = 8'b00000000; // 6904 :   0 - 0x0
      13'h1AF9: dout  = 8'b00000000; // 6905 :   0 - 0x0
      13'h1AFA: dout  = 8'b00000000; // 6906 :   0 - 0x0
      13'h1AFB: dout  = 8'b00000000; // 6907 :   0 - 0x0
      13'h1AFC: dout  = 8'b00000000; // 6908 :   0 - 0x0
      13'h1AFD: dout  = 8'b00000000; // 6909 :   0 - 0x0
      13'h1AFE: dout  = 8'b00000000; // 6910 :   0 - 0x0
      13'h1AFF: dout  = 8'b00000000; // 6911 :   0 - 0x0
      13'h1B00: dout  = 8'b00011111; // 6912 :  31 - 0x1f -- Background 0xb0
      13'h1B01: dout  = 8'b00111111; // 6913 :  63 - 0x3f
      13'h1B02: dout  = 8'b01111111; // 6914 : 127 - 0x7f
      13'h1B03: dout  = 8'b01111111; // 6915 : 127 - 0x7f
      13'h1B04: dout  = 8'b01111111; // 6916 : 127 - 0x7f
      13'h1B05: dout  = 8'b11111111; // 6917 : 255 - 0xff
      13'h1B06: dout  = 8'b11111111; // 6918 : 255 - 0xff
      13'h1B07: dout  = 8'b11111111; // 6919 : 255 - 0xff
      13'h1B08: dout  = 8'b00011111; // 6920 :  31 - 0x1f
      13'h1B09: dout  = 8'b00100000; // 6921 :  32 - 0x20
      13'h1B0A: dout  = 8'b01000000; // 6922 :  64 - 0x40
      13'h1B0B: dout  = 8'b01000000; // 6923 :  64 - 0x40
      13'h1B0C: dout  = 8'b01000000; // 6924 :  64 - 0x40
      13'h1B0D: dout  = 8'b10000000; // 6925 : 128 - 0x80
      13'h1B0E: dout  = 8'b10000010; // 6926 : 130 - 0x82
      13'h1B0F: dout  = 8'b10000010; // 6927 : 130 - 0x82
      13'h1B10: dout  = 8'b11111111; // 6928 : 255 - 0xff -- Background 0xb1
      13'h1B11: dout  = 8'b11111111; // 6929 : 255 - 0xff
      13'h1B12: dout  = 8'b11111111; // 6930 : 255 - 0xff
      13'h1B13: dout  = 8'b01111111; // 6931 : 127 - 0x7f
      13'h1B14: dout  = 8'b01111111; // 6932 : 127 - 0x7f
      13'h1B15: dout  = 8'b01111111; // 6933 : 127 - 0x7f
      13'h1B16: dout  = 8'b00111111; // 6934 :  63 - 0x3f
      13'h1B17: dout  = 8'b00011110; // 6935 :  30 - 0x1e
      13'h1B18: dout  = 8'b10000010; // 6936 : 130 - 0x82
      13'h1B19: dout  = 8'b10000000; // 6937 : 128 - 0x80
      13'h1B1A: dout  = 8'b10100000; // 6938 : 160 - 0xa0
      13'h1B1B: dout  = 8'b01000100; // 6939 :  68 - 0x44
      13'h1B1C: dout  = 8'b01000011; // 6940 :  67 - 0x43
      13'h1B1D: dout  = 8'b01000000; // 6941 :  64 - 0x40
      13'h1B1E: dout  = 8'b00100001; // 6942 :  33 - 0x21
      13'h1B1F: dout  = 8'b00011110; // 6943 :  30 - 0x1e
      13'h1B20: dout  = 8'b11111000; // 6944 : 248 - 0xf8 -- Background 0xb2
      13'h1B21: dout  = 8'b11111100; // 6945 : 252 - 0xfc
      13'h1B22: dout  = 8'b11111110; // 6946 : 254 - 0xfe
      13'h1B23: dout  = 8'b11111110; // 6947 : 254 - 0xfe
      13'h1B24: dout  = 8'b11111110; // 6948 : 254 - 0xfe
      13'h1B25: dout  = 8'b11111111; // 6949 : 255 - 0xff
      13'h1B26: dout  = 8'b11111111; // 6950 : 255 - 0xff
      13'h1B27: dout  = 8'b11111111; // 6951 : 255 - 0xff
      13'h1B28: dout  = 8'b11111000; // 6952 : 248 - 0xf8
      13'h1B29: dout  = 8'b00000100; // 6953 :   4 - 0x4
      13'h1B2A: dout  = 8'b00000010; // 6954 :   2 - 0x2
      13'h1B2B: dout  = 8'b00000010; // 6955 :   2 - 0x2
      13'h1B2C: dout  = 8'b00000010; // 6956 :   2 - 0x2
      13'h1B2D: dout  = 8'b00000001; // 6957 :   1 - 0x1
      13'h1B2E: dout  = 8'b01000001; // 6958 :  65 - 0x41
      13'h1B2F: dout  = 8'b01000001; // 6959 :  65 - 0x41
      13'h1B30: dout  = 8'b11111111; // 6960 : 255 - 0xff -- Background 0xb3
      13'h1B31: dout  = 8'b11111111; // 6961 : 255 - 0xff
      13'h1B32: dout  = 8'b11111111; // 6962 : 255 - 0xff
      13'h1B33: dout  = 8'b11111110; // 6963 : 254 - 0xfe
      13'h1B34: dout  = 8'b11111110; // 6964 : 254 - 0xfe
      13'h1B35: dout  = 8'b11111110; // 6965 : 254 - 0xfe
      13'h1B36: dout  = 8'b11111100; // 6966 : 252 - 0xfc
      13'h1B37: dout  = 8'b01111000; // 6967 : 120 - 0x78
      13'h1B38: dout  = 8'b01000001; // 6968 :  65 - 0x41
      13'h1B39: dout  = 8'b00000001; // 6969 :   1 - 0x1
      13'h1B3A: dout  = 8'b00000101; // 6970 :   5 - 0x5
      13'h1B3B: dout  = 8'b00100010; // 6971 :  34 - 0x22
      13'h1B3C: dout  = 8'b11000010; // 6972 : 194 - 0xc2
      13'h1B3D: dout  = 8'b00000010; // 6973 :   2 - 0x2
      13'h1B3E: dout  = 8'b10000100; // 6974 : 132 - 0x84
      13'h1B3F: dout  = 8'b01111000; // 6975 : 120 - 0x78
      13'h1B40: dout  = 8'b01111111; // 6976 : 127 - 0x7f -- Background 0xb4
      13'h1B41: dout  = 8'b10000000; // 6977 : 128 - 0x80
      13'h1B42: dout  = 8'b10000000; // 6978 : 128 - 0x80
      13'h1B43: dout  = 8'b10000000; // 6979 : 128 - 0x80
      13'h1B44: dout  = 8'b10000000; // 6980 : 128 - 0x80
      13'h1B45: dout  = 8'b10000000; // 6981 : 128 - 0x80
      13'h1B46: dout  = 8'b10000000; // 6982 : 128 - 0x80
      13'h1B47: dout  = 8'b10000000; // 6983 : 128 - 0x80
      13'h1B48: dout  = 8'b10000000; // 6984 : 128 - 0x80
      13'h1B49: dout  = 8'b01111111; // 6985 : 127 - 0x7f
      13'h1B4A: dout  = 8'b01111111; // 6986 : 127 - 0x7f
      13'h1B4B: dout  = 8'b01111111; // 6987 : 127 - 0x7f
      13'h1B4C: dout  = 8'b01111111; // 6988 : 127 - 0x7f
      13'h1B4D: dout  = 8'b01111111; // 6989 : 127 - 0x7f
      13'h1B4E: dout  = 8'b01111111; // 6990 : 127 - 0x7f
      13'h1B4F: dout  = 8'b01111111; // 6991 : 127 - 0x7f
      13'h1B50: dout  = 8'b11011110; // 6992 : 222 - 0xde -- Background 0xb5
      13'h1B51: dout  = 8'b01100001; // 6993 :  97 - 0x61
      13'h1B52: dout  = 8'b01100001; // 6994 :  97 - 0x61
      13'h1B53: dout  = 8'b01100001; // 6995 :  97 - 0x61
      13'h1B54: dout  = 8'b01110001; // 6996 : 113 - 0x71
      13'h1B55: dout  = 8'b01011110; // 6997 :  94 - 0x5e
      13'h1B56: dout  = 8'b01111111; // 6998 : 127 - 0x7f
      13'h1B57: dout  = 8'b01100001; // 6999 :  97 - 0x61
      13'h1B58: dout  = 8'b01100001; // 7000 :  97 - 0x61
      13'h1B59: dout  = 8'b11011111; // 7001 : 223 - 0xdf
      13'h1B5A: dout  = 8'b11011111; // 7002 : 223 - 0xdf
      13'h1B5B: dout  = 8'b11011111; // 7003 : 223 - 0xdf
      13'h1B5C: dout  = 8'b11011111; // 7004 : 223 - 0xdf
      13'h1B5D: dout  = 8'b11111111; // 7005 : 255 - 0xff
      13'h1B5E: dout  = 8'b11000001; // 7006 : 193 - 0xc1
      13'h1B5F: dout  = 8'b11011111; // 7007 : 223 - 0xdf
      13'h1B60: dout  = 8'b10000000; // 7008 : 128 - 0x80 -- Background 0xb6
      13'h1B61: dout  = 8'b10000000; // 7009 : 128 - 0x80
      13'h1B62: dout  = 8'b11000000; // 7010 : 192 - 0xc0
      13'h1B63: dout  = 8'b11110000; // 7011 : 240 - 0xf0
      13'h1B64: dout  = 8'b10111111; // 7012 : 191 - 0xbf
      13'h1B65: dout  = 8'b10001111; // 7013 : 143 - 0x8f
      13'h1B66: dout  = 8'b10000001; // 7014 : 129 - 0x81
      13'h1B67: dout  = 8'b01111110; // 7015 : 126 - 0x7e
      13'h1B68: dout  = 8'b01111111; // 7016 : 127 - 0x7f
      13'h1B69: dout  = 8'b01111111; // 7017 : 127 - 0x7f
      13'h1B6A: dout  = 8'b11111111; // 7018 : 255 - 0xff
      13'h1B6B: dout  = 8'b00111111; // 7019 :  63 - 0x3f
      13'h1B6C: dout  = 8'b01001111; // 7020 :  79 - 0x4f
      13'h1B6D: dout  = 8'b01110001; // 7021 : 113 - 0x71
      13'h1B6E: dout  = 8'b01111111; // 7022 : 127 - 0x7f
      13'h1B6F: dout  = 8'b11111111; // 7023 : 255 - 0xff
      13'h1B70: dout  = 8'b01100001; // 7024 :  97 - 0x61 -- Background 0xb7
      13'h1B71: dout  = 8'b01100001; // 7025 :  97 - 0x61
      13'h1B72: dout  = 8'b11000001; // 7026 : 193 - 0xc1
      13'h1B73: dout  = 8'b11000001; // 7027 : 193 - 0xc1
      13'h1B74: dout  = 8'b10000001; // 7028 : 129 - 0x81
      13'h1B75: dout  = 8'b10000001; // 7029 : 129 - 0x81
      13'h1B76: dout  = 8'b10000011; // 7030 : 131 - 0x83
      13'h1B77: dout  = 8'b11111110; // 7031 : 254 - 0xfe
      13'h1B78: dout  = 8'b11011111; // 7032 : 223 - 0xdf
      13'h1B79: dout  = 8'b11011111; // 7033 : 223 - 0xdf
      13'h1B7A: dout  = 8'b10111111; // 7034 : 191 - 0xbf
      13'h1B7B: dout  = 8'b10111111; // 7035 : 191 - 0xbf
      13'h1B7C: dout  = 8'b01111111; // 7036 : 127 - 0x7f
      13'h1B7D: dout  = 8'b01111111; // 7037 : 127 - 0x7f
      13'h1B7E: dout  = 8'b01111111; // 7038 : 127 - 0x7f
      13'h1B7F: dout  = 8'b01111111; // 7039 : 127 - 0x7f
      13'h1B80: dout  = 8'b00000000; // 7040 :   0 - 0x0 -- Background 0xb8
      13'h1B81: dout  = 8'b00000000; // 7041 :   0 - 0x0
      13'h1B82: dout  = 8'b00000011; // 7042 :   3 - 0x3
      13'h1B83: dout  = 8'b00001111; // 7043 :  15 - 0xf
      13'h1B84: dout  = 8'b00011111; // 7044 :  31 - 0x1f
      13'h1B85: dout  = 8'b00111111; // 7045 :  63 - 0x3f
      13'h1B86: dout  = 8'b01111111; // 7046 : 127 - 0x7f
      13'h1B87: dout  = 8'b01111111; // 7047 : 127 - 0x7f
      13'h1B88: dout  = 8'b00000000; // 7048 :   0 - 0x0
      13'h1B89: dout  = 8'b00000000; // 7049 :   0 - 0x0
      13'h1B8A: dout  = 8'b00000011; // 7050 :   3 - 0x3
      13'h1B8B: dout  = 8'b00001100; // 7051 :  12 - 0xc
      13'h1B8C: dout  = 8'b00010000; // 7052 :  16 - 0x10
      13'h1B8D: dout  = 8'b00100000; // 7053 :  32 - 0x20
      13'h1B8E: dout  = 8'b01000000; // 7054 :  64 - 0x40
      13'h1B8F: dout  = 8'b01000000; // 7055 :  64 - 0x40
      13'h1B90: dout  = 8'b00000000; // 7056 :   0 - 0x0 -- Background 0xb9
      13'h1B91: dout  = 8'b00000000; // 7057 :   0 - 0x0
      13'h1B92: dout  = 8'b11000000; // 7058 : 192 - 0xc0
      13'h1B93: dout  = 8'b11110000; // 7059 : 240 - 0xf0
      13'h1B94: dout  = 8'b11111000; // 7060 : 248 - 0xf8
      13'h1B95: dout  = 8'b11111100; // 7061 : 252 - 0xfc
      13'h1B96: dout  = 8'b11111110; // 7062 : 254 - 0xfe
      13'h1B97: dout  = 8'b11111110; // 7063 : 254 - 0xfe
      13'h1B98: dout  = 8'b00000000; // 7064 :   0 - 0x0
      13'h1B99: dout  = 8'b00000000; // 7065 :   0 - 0x0
      13'h1B9A: dout  = 8'b11000000; // 7066 : 192 - 0xc0
      13'h1B9B: dout  = 8'b00110000; // 7067 :  48 - 0x30
      13'h1B9C: dout  = 8'b00001000; // 7068 :   8 - 0x8
      13'h1B9D: dout  = 8'b00000100; // 7069 :   4 - 0x4
      13'h1B9E: dout  = 8'b00000010; // 7070 :   2 - 0x2
      13'h1B9F: dout  = 8'b00000010; // 7071 :   2 - 0x2
      13'h1BA0: dout  = 8'b11111111; // 7072 : 255 - 0xff -- Background 0xba
      13'h1BA1: dout  = 8'b11111111; // 7073 : 255 - 0xff
      13'h1BA2: dout  = 8'b11111111; // 7074 : 255 - 0xff
      13'h1BA3: dout  = 8'b11111111; // 7075 : 255 - 0xff
      13'h1BA4: dout  = 8'b11111111; // 7076 : 255 - 0xff
      13'h1BA5: dout  = 8'b11111111; // 7077 : 255 - 0xff
      13'h1BA6: dout  = 8'b11111111; // 7078 : 255 - 0xff
      13'h1BA7: dout  = 8'b11111111; // 7079 : 255 - 0xff
      13'h1BA8: dout  = 8'b10000000; // 7080 : 128 - 0x80
      13'h1BA9: dout  = 8'b10000000; // 7081 : 128 - 0x80
      13'h1BAA: dout  = 8'b10000000; // 7082 : 128 - 0x80
      13'h1BAB: dout  = 8'b10000000; // 7083 : 128 - 0x80
      13'h1BAC: dout  = 8'b10000000; // 7084 : 128 - 0x80
      13'h1BAD: dout  = 8'b10000000; // 7085 : 128 - 0x80
      13'h1BAE: dout  = 8'b10000000; // 7086 : 128 - 0x80
      13'h1BAF: dout  = 8'b10000000; // 7087 : 128 - 0x80
      13'h1BB0: dout  = 8'b11111111; // 7088 : 255 - 0xff -- Background 0xbb
      13'h1BB1: dout  = 8'b11111111; // 7089 : 255 - 0xff
      13'h1BB2: dout  = 8'b11111111; // 7090 : 255 - 0xff
      13'h1BB3: dout  = 8'b11111111; // 7091 : 255 - 0xff
      13'h1BB4: dout  = 8'b11111111; // 7092 : 255 - 0xff
      13'h1BB5: dout  = 8'b11111111; // 7093 : 255 - 0xff
      13'h1BB6: dout  = 8'b11111111; // 7094 : 255 - 0xff
      13'h1BB7: dout  = 8'b11111111; // 7095 : 255 - 0xff
      13'h1BB8: dout  = 8'b00000001; // 7096 :   1 - 0x1
      13'h1BB9: dout  = 8'b00000001; // 7097 :   1 - 0x1
      13'h1BBA: dout  = 8'b00000001; // 7098 :   1 - 0x1
      13'h1BBB: dout  = 8'b00000001; // 7099 :   1 - 0x1
      13'h1BBC: dout  = 8'b00000001; // 7100 :   1 - 0x1
      13'h1BBD: dout  = 8'b00000001; // 7101 :   1 - 0x1
      13'h1BBE: dout  = 8'b00000001; // 7102 :   1 - 0x1
      13'h1BBF: dout  = 8'b00000001; // 7103 :   1 - 0x1
      13'h1BC0: dout  = 8'b01111111; // 7104 : 127 - 0x7f -- Background 0xbc
      13'h1BC1: dout  = 8'b01111111; // 7105 : 127 - 0x7f
      13'h1BC2: dout  = 8'b01111111; // 7106 : 127 - 0x7f
      13'h1BC3: dout  = 8'b00111111; // 7107 :  63 - 0x3f
      13'h1BC4: dout  = 8'b00111111; // 7108 :  63 - 0x3f
      13'h1BC5: dout  = 8'b00011111; // 7109 :  31 - 0x1f
      13'h1BC6: dout  = 8'b00001111; // 7110 :  15 - 0xf
      13'h1BC7: dout  = 8'b00000111; // 7111 :   7 - 0x7
      13'h1BC8: dout  = 8'b01000000; // 7112 :  64 - 0x40
      13'h1BC9: dout  = 8'b01000000; // 7113 :  64 - 0x40
      13'h1BCA: dout  = 8'b01000000; // 7114 :  64 - 0x40
      13'h1BCB: dout  = 8'b00100000; // 7115 :  32 - 0x20
      13'h1BCC: dout  = 8'b00110000; // 7116 :  48 - 0x30
      13'h1BCD: dout  = 8'b00011100; // 7117 :  28 - 0x1c
      13'h1BCE: dout  = 8'b00001111; // 7118 :  15 - 0xf
      13'h1BCF: dout  = 8'b00000111; // 7119 :   7 - 0x7
      13'h1BD0: dout  = 8'b11111110; // 7120 : 254 - 0xfe -- Background 0xbd
      13'h1BD1: dout  = 8'b11111110; // 7121 : 254 - 0xfe
      13'h1BD2: dout  = 8'b11111110; // 7122 : 254 - 0xfe
      13'h1BD3: dout  = 8'b11111100; // 7123 : 252 - 0xfc
      13'h1BD4: dout  = 8'b11111100; // 7124 : 252 - 0xfc
      13'h1BD5: dout  = 8'b11111000; // 7125 : 248 - 0xf8
      13'h1BD6: dout  = 8'b11110000; // 7126 : 240 - 0xf0
      13'h1BD7: dout  = 8'b11110000; // 7127 : 240 - 0xf0
      13'h1BD8: dout  = 8'b00000010; // 7128 :   2 - 0x2
      13'h1BD9: dout  = 8'b00000010; // 7129 :   2 - 0x2
      13'h1BDA: dout  = 8'b00000010; // 7130 :   2 - 0x2
      13'h1BDB: dout  = 8'b00000100; // 7131 :   4 - 0x4
      13'h1BDC: dout  = 8'b00001100; // 7132 :  12 - 0xc
      13'h1BDD: dout  = 8'b00111000; // 7133 :  56 - 0x38
      13'h1BDE: dout  = 8'b11110000; // 7134 : 240 - 0xf0
      13'h1BDF: dout  = 8'b11110000; // 7135 : 240 - 0xf0
      13'h1BE0: dout  = 8'b00001111; // 7136 :  15 - 0xf -- Background 0xbe
      13'h1BE1: dout  = 8'b00001111; // 7137 :  15 - 0xf
      13'h1BE2: dout  = 8'b00001111; // 7138 :  15 - 0xf
      13'h1BE3: dout  = 8'b00001111; // 7139 :  15 - 0xf
      13'h1BE4: dout  = 8'b00001111; // 7140 :  15 - 0xf
      13'h1BE5: dout  = 8'b00001111; // 7141 :  15 - 0xf
      13'h1BE6: dout  = 8'b00000111; // 7142 :   7 - 0x7
      13'h1BE7: dout  = 8'b00001111; // 7143 :  15 - 0xf
      13'h1BE8: dout  = 8'b00001000; // 7144 :   8 - 0x8
      13'h1BE9: dout  = 8'b00001000; // 7145 :   8 - 0x8
      13'h1BEA: dout  = 8'b00001000; // 7146 :   8 - 0x8
      13'h1BEB: dout  = 8'b00001000; // 7147 :   8 - 0x8
      13'h1BEC: dout  = 8'b00001000; // 7148 :   8 - 0x8
      13'h1BED: dout  = 8'b00001100; // 7149 :  12 - 0xc
      13'h1BEE: dout  = 8'b00000101; // 7150 :   5 - 0x5
      13'h1BEF: dout  = 8'b00001010; // 7151 :  10 - 0xa
      13'h1BF0: dout  = 8'b11110000; // 7152 : 240 - 0xf0 -- Background 0xbf
      13'h1BF1: dout  = 8'b11110000; // 7153 : 240 - 0xf0
      13'h1BF2: dout  = 8'b11110000; // 7154 : 240 - 0xf0
      13'h1BF3: dout  = 8'b11110000; // 7155 : 240 - 0xf0
      13'h1BF4: dout  = 8'b11110000; // 7156 : 240 - 0xf0
      13'h1BF5: dout  = 8'b11110000; // 7157 : 240 - 0xf0
      13'h1BF6: dout  = 8'b11100000; // 7158 : 224 - 0xe0
      13'h1BF7: dout  = 8'b11110000; // 7159 : 240 - 0xf0
      13'h1BF8: dout  = 8'b00010000; // 7160 :  16 - 0x10
      13'h1BF9: dout  = 8'b01010000; // 7161 :  80 - 0x50
      13'h1BFA: dout  = 8'b01010000; // 7162 :  80 - 0x50
      13'h1BFB: dout  = 8'b01010000; // 7163 :  80 - 0x50
      13'h1BFC: dout  = 8'b01010000; // 7164 :  80 - 0x50
      13'h1BFD: dout  = 8'b00110000; // 7165 :  48 - 0x30
      13'h1BFE: dout  = 8'b10100000; // 7166 : 160 - 0xa0
      13'h1BFF: dout  = 8'b01010000; // 7167 :  80 - 0x50
      13'h1C00: dout  = 8'b10000001; // 7168 : 129 - 0x81 -- Background 0xc0
      13'h1C01: dout  = 8'b11000001; // 7169 : 193 - 0xc1
      13'h1C02: dout  = 8'b10100011; // 7170 : 163 - 0xa3
      13'h1C03: dout  = 8'b10100011; // 7171 : 163 - 0xa3
      13'h1C04: dout  = 8'b10011101; // 7172 : 157 - 0x9d
      13'h1C05: dout  = 8'b10000001; // 7173 : 129 - 0x81
      13'h1C06: dout  = 8'b10000001; // 7174 : 129 - 0x81
      13'h1C07: dout  = 8'b10000001; // 7175 : 129 - 0x81
      13'h1C08: dout  = 8'b00000000; // 7176 :   0 - 0x0
      13'h1C09: dout  = 8'b01000001; // 7177 :  65 - 0x41
      13'h1C0A: dout  = 8'b00100010; // 7178 :  34 - 0x22
      13'h1C0B: dout  = 8'b00100010; // 7179 :  34 - 0x22
      13'h1C0C: dout  = 8'b00011100; // 7180 :  28 - 0x1c
      13'h1C0D: dout  = 8'b00000000; // 7181 :   0 - 0x0
      13'h1C0E: dout  = 8'b00000000; // 7182 :   0 - 0x0
      13'h1C0F: dout  = 8'b00000000; // 7183 :   0 - 0x0
      13'h1C10: dout  = 8'b11100011; // 7184 : 227 - 0xe3 -- Background 0xc1
      13'h1C11: dout  = 8'b11110111; // 7185 : 247 - 0xf7
      13'h1C12: dout  = 8'b11000001; // 7186 : 193 - 0xc1
      13'h1C13: dout  = 8'b11000001; // 7187 : 193 - 0xc1
      13'h1C14: dout  = 8'b11000001; // 7188 : 193 - 0xc1
      13'h1C15: dout  = 8'b11000001; // 7189 : 193 - 0xc1
      13'h1C16: dout  = 8'b11110111; // 7190 : 247 - 0xf7
      13'h1C17: dout  = 8'b11100011; // 7191 : 227 - 0xe3
      13'h1C18: dout  = 8'b11100011; // 7192 : 227 - 0xe3
      13'h1C19: dout  = 8'b00010100; // 7193 :  20 - 0x14
      13'h1C1A: dout  = 8'b00111110; // 7194 :  62 - 0x3e
      13'h1C1B: dout  = 8'b00111110; // 7195 :  62 - 0x3e
      13'h1C1C: dout  = 8'b00111110; // 7196 :  62 - 0x3e
      13'h1C1D: dout  = 8'b00111110; // 7197 :  62 - 0x3e
      13'h1C1E: dout  = 8'b00010100; // 7198 :  20 - 0x14
      13'h1C1F: dout  = 8'b11100011; // 7199 : 227 - 0xe3
      13'h1C20: dout  = 8'b00000000; // 7200 :   0 - 0x0 -- Background 0xc2
      13'h1C21: dout  = 8'b00000000; // 7201 :   0 - 0x0
      13'h1C22: dout  = 8'b00000111; // 7202 :   7 - 0x7
      13'h1C23: dout  = 8'b00001111; // 7203 :  15 - 0xf
      13'h1C24: dout  = 8'b00001100; // 7204 :  12 - 0xc
      13'h1C25: dout  = 8'b00011011; // 7205 :  27 - 0x1b
      13'h1C26: dout  = 8'b00011011; // 7206 :  27 - 0x1b
      13'h1C27: dout  = 8'b00011011; // 7207 :  27 - 0x1b
      13'h1C28: dout  = 8'b11111111; // 7208 : 255 - 0xff
      13'h1C29: dout  = 8'b11111111; // 7209 : 255 - 0xff
      13'h1C2A: dout  = 8'b11111000; // 7210 : 248 - 0xf8
      13'h1C2B: dout  = 8'b11110000; // 7211 : 240 - 0xf0
      13'h1C2C: dout  = 8'b11110000; // 7212 : 240 - 0xf0
      13'h1C2D: dout  = 8'b11100000; // 7213 : 224 - 0xe0
      13'h1C2E: dout  = 8'b11100000; // 7214 : 224 - 0xe0
      13'h1C2F: dout  = 8'b11100000; // 7215 : 224 - 0xe0
      13'h1C30: dout  = 8'b00000000; // 7216 :   0 - 0x0 -- Background 0xc3
      13'h1C31: dout  = 8'b00000000; // 7217 :   0 - 0x0
      13'h1C32: dout  = 8'b11100000; // 7218 : 224 - 0xe0
      13'h1C33: dout  = 8'b11110000; // 7219 : 240 - 0xf0
      13'h1C34: dout  = 8'b11110000; // 7220 : 240 - 0xf0
      13'h1C35: dout  = 8'b11111000; // 7221 : 248 - 0xf8
      13'h1C36: dout  = 8'b11111000; // 7222 : 248 - 0xf8
      13'h1C37: dout  = 8'b11111000; // 7223 : 248 - 0xf8
      13'h1C38: dout  = 8'b11111111; // 7224 : 255 - 0xff
      13'h1C39: dout  = 8'b11111111; // 7225 : 255 - 0xff
      13'h1C3A: dout  = 8'b01111111; // 7226 : 127 - 0x7f
      13'h1C3B: dout  = 8'b00111111; // 7227 :  63 - 0x3f
      13'h1C3C: dout  = 8'b00111111; // 7228 :  63 - 0x3f
      13'h1C3D: dout  = 8'b10011111; // 7229 : 159 - 0x9f
      13'h1C3E: dout  = 8'b10011111; // 7230 : 159 - 0x9f
      13'h1C3F: dout  = 8'b10011111; // 7231 : 159 - 0x9f
      13'h1C40: dout  = 8'b00011011; // 7232 :  27 - 0x1b -- Background 0xc4
      13'h1C41: dout  = 8'b00011011; // 7233 :  27 - 0x1b
      13'h1C42: dout  = 8'b00011011; // 7234 :  27 - 0x1b
      13'h1C43: dout  = 8'b00011011; // 7235 :  27 - 0x1b
      13'h1C44: dout  = 8'b00011011; // 7236 :  27 - 0x1b
      13'h1C45: dout  = 8'b00001111; // 7237 :  15 - 0xf
      13'h1C46: dout  = 8'b00001111; // 7238 :  15 - 0xf
      13'h1C47: dout  = 8'b00000111; // 7239 :   7 - 0x7
      13'h1C48: dout  = 8'b11100000; // 7240 : 224 - 0xe0
      13'h1C49: dout  = 8'b11100000; // 7241 : 224 - 0xe0
      13'h1C4A: dout  = 8'b11100000; // 7242 : 224 - 0xe0
      13'h1C4B: dout  = 8'b11100000; // 7243 : 224 - 0xe0
      13'h1C4C: dout  = 8'b11100000; // 7244 : 224 - 0xe0
      13'h1C4D: dout  = 8'b11110011; // 7245 : 243 - 0xf3
      13'h1C4E: dout  = 8'b11110000; // 7246 : 240 - 0xf0
      13'h1C4F: dout  = 8'b11111000; // 7247 : 248 - 0xf8
      13'h1C50: dout  = 8'b11111000; // 7248 : 248 - 0xf8 -- Background 0xc5
      13'h1C51: dout  = 8'b11111000; // 7249 : 248 - 0xf8
      13'h1C52: dout  = 8'b11111000; // 7250 : 248 - 0xf8
      13'h1C53: dout  = 8'b11111000; // 7251 : 248 - 0xf8
      13'h1C54: dout  = 8'b11111000; // 7252 : 248 - 0xf8
      13'h1C55: dout  = 8'b11110000; // 7253 : 240 - 0xf0
      13'h1C56: dout  = 8'b11110000; // 7254 : 240 - 0xf0
      13'h1C57: dout  = 8'b11100000; // 7255 : 224 - 0xe0
      13'h1C58: dout  = 8'b10011111; // 7256 : 159 - 0x9f
      13'h1C59: dout  = 8'b10011111; // 7257 : 159 - 0x9f
      13'h1C5A: dout  = 8'b10011111; // 7258 : 159 - 0x9f
      13'h1C5B: dout  = 8'b10011111; // 7259 : 159 - 0x9f
      13'h1C5C: dout  = 8'b10011111; // 7260 : 159 - 0x9f
      13'h1C5D: dout  = 8'b00111111; // 7261 :  63 - 0x3f
      13'h1C5E: dout  = 8'b00111111; // 7262 :  63 - 0x3f
      13'h1C5F: dout  = 8'b01111111; // 7263 : 127 - 0x7f
      13'h1C60: dout  = 8'b11100000; // 7264 : 224 - 0xe0 -- Background 0xc6
      13'h1C61: dout  = 8'b11111111; // 7265 : 255 - 0xff
      13'h1C62: dout  = 8'b11111111; // 7266 : 255 - 0xff
      13'h1C63: dout  = 8'b11111111; // 7267 : 255 - 0xff
      13'h1C64: dout  = 8'b11111111; // 7268 : 255 - 0xff
      13'h1C65: dout  = 8'b11111111; // 7269 : 255 - 0xff
      13'h1C66: dout  = 8'b11111111; // 7270 : 255 - 0xff
      13'h1C67: dout  = 8'b11111111; // 7271 : 255 - 0xff
      13'h1C68: dout  = 8'b00000000; // 7272 :   0 - 0x0
      13'h1C69: dout  = 8'b01110000; // 7273 : 112 - 0x70
      13'h1C6A: dout  = 8'b00011111; // 7274 :  31 - 0x1f
      13'h1C6B: dout  = 8'b00010000; // 7275 :  16 - 0x10
      13'h1C6C: dout  = 8'b01110000; // 7276 : 112 - 0x70
      13'h1C6D: dout  = 8'b01111111; // 7277 : 127 - 0x7f
      13'h1C6E: dout  = 8'b01111111; // 7278 : 127 - 0x7f
      13'h1C6F: dout  = 8'b01111111; // 7279 : 127 - 0x7f
      13'h1C70: dout  = 8'b00000111; // 7280 :   7 - 0x7 -- Background 0xc7
      13'h1C71: dout  = 8'b11111111; // 7281 : 255 - 0xff
      13'h1C72: dout  = 8'b11111111; // 7282 : 255 - 0xff
      13'h1C73: dout  = 8'b11111111; // 7283 : 255 - 0xff
      13'h1C74: dout  = 8'b11111111; // 7284 : 255 - 0xff
      13'h1C75: dout  = 8'b11111111; // 7285 : 255 - 0xff
      13'h1C76: dout  = 8'b11111111; // 7286 : 255 - 0xff
      13'h1C77: dout  = 8'b11111111; // 7287 : 255 - 0xff
      13'h1C78: dout  = 8'b00000000; // 7288 :   0 - 0x0
      13'h1C79: dout  = 8'b00000011; // 7289 :   3 - 0x3
      13'h1C7A: dout  = 8'b11111000; // 7290 : 248 - 0xf8
      13'h1C7B: dout  = 8'b00000000; // 7291 :   0 - 0x0
      13'h1C7C: dout  = 8'b00000011; // 7292 :   3 - 0x3
      13'h1C7D: dout  = 8'b11111011; // 7293 : 251 - 0xfb
      13'h1C7E: dout  = 8'b11111011; // 7294 : 251 - 0xfb
      13'h1C7F: dout  = 8'b11111011; // 7295 : 251 - 0xfb
      13'h1C80: dout  = 8'b11111111; // 7296 : 255 - 0xff -- Background 0xc8
      13'h1C81: dout  = 8'b11111111; // 7297 : 255 - 0xff
      13'h1C82: dout  = 8'b11111111; // 7298 : 255 - 0xff
      13'h1C83: dout  = 8'b11111111; // 7299 : 255 - 0xff
      13'h1C84: dout  = 8'b11111111; // 7300 : 255 - 0xff
      13'h1C85: dout  = 8'b11111110; // 7301 : 254 - 0xfe
      13'h1C86: dout  = 8'b11111111; // 7302 : 255 - 0xff
      13'h1C87: dout  = 8'b11101111; // 7303 : 239 - 0xef
      13'h1C88: dout  = 8'b01111100; // 7304 : 124 - 0x7c
      13'h1C89: dout  = 8'b01111011; // 7305 : 123 - 0x7b
      13'h1C8A: dout  = 8'b01110110; // 7306 : 118 - 0x76
      13'h1C8B: dout  = 8'b01110101; // 7307 : 117 - 0x75
      13'h1C8C: dout  = 8'b01110101; // 7308 : 117 - 0x75
      13'h1C8D: dout  = 8'b01110111; // 7309 : 119 - 0x77
      13'h1C8E: dout  = 8'b00010111; // 7310 :  23 - 0x17
      13'h1C8F: dout  = 8'b01100111; // 7311 : 103 - 0x67
      13'h1C90: dout  = 8'b11111111; // 7312 : 255 - 0xff -- Background 0xc9
      13'h1C91: dout  = 8'b11011111; // 7313 : 223 - 0xdf
      13'h1C92: dout  = 8'b11101111; // 7314 : 239 - 0xef
      13'h1C93: dout  = 8'b10101111; // 7315 : 175 - 0xaf
      13'h1C94: dout  = 8'b10101111; // 7316 : 175 - 0xaf
      13'h1C95: dout  = 8'b01101111; // 7317 : 111 - 0x6f
      13'h1C96: dout  = 8'b11101111; // 7318 : 239 - 0xef
      13'h1C97: dout  = 8'b11100111; // 7319 : 231 - 0xe7
      13'h1C98: dout  = 8'b00111011; // 7320 :  59 - 0x3b
      13'h1C99: dout  = 8'b11111011; // 7321 : 251 - 0xfb
      13'h1C9A: dout  = 8'b01111011; // 7322 : 123 - 0x7b
      13'h1C9B: dout  = 8'b11111011; // 7323 : 251 - 0xfb
      13'h1C9C: dout  = 8'b11111011; // 7324 : 251 - 0xfb
      13'h1C9D: dout  = 8'b11110011; // 7325 : 243 - 0xf3
      13'h1C9E: dout  = 8'b11111000; // 7326 : 248 - 0xf8
      13'h1C9F: dout  = 8'b11110011; // 7327 : 243 - 0xf3
      13'h1CA0: dout  = 8'b00011111; // 7328 :  31 - 0x1f -- Background 0xca
      13'h1CA1: dout  = 8'b00011111; // 7329 :  31 - 0x1f
      13'h1CA2: dout  = 8'b00111111; // 7330 :  63 - 0x3f
      13'h1CA3: dout  = 8'b00111111; // 7331 :  63 - 0x3f
      13'h1CA4: dout  = 8'b01110000; // 7332 : 112 - 0x70
      13'h1CA5: dout  = 8'b01100011; // 7333 :  99 - 0x63
      13'h1CA6: dout  = 8'b11100111; // 7334 : 231 - 0xe7
      13'h1CA7: dout  = 8'b11100101; // 7335 : 229 - 0xe5
      13'h1CA8: dout  = 8'b00001111; // 7336 :  15 - 0xf
      13'h1CA9: dout  = 8'b00001111; // 7337 :  15 - 0xf
      13'h1CAA: dout  = 8'b00011111; // 7338 :  31 - 0x1f
      13'h1CAB: dout  = 8'b00011111; // 7339 :  31 - 0x1f
      13'h1CAC: dout  = 8'b00111111; // 7340 :  63 - 0x3f
      13'h1CAD: dout  = 8'b00111100; // 7341 :  60 - 0x3c
      13'h1CAE: dout  = 8'b01111000; // 7342 : 120 - 0x78
      13'h1CAF: dout  = 8'b01111010; // 7343 : 122 - 0x7a
      13'h1CB0: dout  = 8'b11110000; // 7344 : 240 - 0xf0 -- Background 0xcb
      13'h1CB1: dout  = 8'b11110000; // 7345 : 240 - 0xf0
      13'h1CB2: dout  = 8'b11111000; // 7346 : 248 - 0xf8
      13'h1CB3: dout  = 8'b11111000; // 7347 : 248 - 0xf8
      13'h1CB4: dout  = 8'b00001100; // 7348 :  12 - 0xc
      13'h1CB5: dout  = 8'b11000100; // 7349 : 196 - 0xc4
      13'h1CB6: dout  = 8'b11100100; // 7350 : 228 - 0xe4
      13'h1CB7: dout  = 8'b10100110; // 7351 : 166 - 0xa6
      13'h1CB8: dout  = 8'b11111000; // 7352 : 248 - 0xf8
      13'h1CB9: dout  = 8'b11111000; // 7353 : 248 - 0xf8
      13'h1CBA: dout  = 8'b11111100; // 7354 : 252 - 0xfc
      13'h1CBB: dout  = 8'b11111100; // 7355 : 252 - 0xfc
      13'h1CBC: dout  = 8'b11111110; // 7356 : 254 - 0xfe
      13'h1CBD: dout  = 8'b00111110; // 7357 :  62 - 0x3e
      13'h1CBE: dout  = 8'b00011110; // 7358 :  30 - 0x1e
      13'h1CBF: dout  = 8'b01011111; // 7359 :  95 - 0x5f
      13'h1CC0: dout  = 8'b11101001; // 7360 : 233 - 0xe9 -- Background 0xcc
      13'h1CC1: dout  = 8'b11101001; // 7361 : 233 - 0xe9
      13'h1CC2: dout  = 8'b11101001; // 7362 : 233 - 0xe9
      13'h1CC3: dout  = 8'b11101111; // 7363 : 239 - 0xef
      13'h1CC4: dout  = 8'b11100010; // 7364 : 226 - 0xe2
      13'h1CC5: dout  = 8'b11100011; // 7365 : 227 - 0xe3
      13'h1CC6: dout  = 8'b11110000; // 7366 : 240 - 0xf0
      13'h1CC7: dout  = 8'b11111111; // 7367 : 255 - 0xff
      13'h1CC8: dout  = 8'b01110110; // 7368 : 118 - 0x76
      13'h1CC9: dout  = 8'b01110110; // 7369 : 118 - 0x76
      13'h1CCA: dout  = 8'b01110110; // 7370 : 118 - 0x76
      13'h1CCB: dout  = 8'b01110000; // 7371 : 112 - 0x70
      13'h1CCC: dout  = 8'b01111101; // 7372 : 125 - 0x7d
      13'h1CCD: dout  = 8'b01111100; // 7373 : 124 - 0x7c
      13'h1CCE: dout  = 8'b01111111; // 7374 : 127 - 0x7f
      13'h1CCF: dout  = 8'b01111111; // 7375 : 127 - 0x7f
      13'h1CD0: dout  = 8'b10010110; // 7376 : 150 - 0x96 -- Background 0xcd
      13'h1CD1: dout  = 8'b10010110; // 7377 : 150 - 0x96
      13'h1CD2: dout  = 8'b10010110; // 7378 : 150 - 0x96
      13'h1CD3: dout  = 8'b11110110; // 7379 : 246 - 0xf6
      13'h1CD4: dout  = 8'b01000110; // 7380 :  70 - 0x46
      13'h1CD5: dout  = 8'b11000110; // 7381 : 198 - 0xc6
      13'h1CD6: dout  = 8'b00001110; // 7382 :  14 - 0xe
      13'h1CD7: dout  = 8'b11111110; // 7383 : 254 - 0xfe
      13'h1CD8: dout  = 8'b01101111; // 7384 : 111 - 0x6f
      13'h1CD9: dout  = 8'b01101111; // 7385 : 111 - 0x6f
      13'h1CDA: dout  = 8'b01101111; // 7386 : 111 - 0x6f
      13'h1CDB: dout  = 8'b00001111; // 7387 :  15 - 0xf
      13'h1CDC: dout  = 8'b10111111; // 7388 : 191 - 0xbf
      13'h1CDD: dout  = 8'b00111111; // 7389 :  63 - 0x3f
      13'h1CDE: dout  = 8'b11111111; // 7390 : 255 - 0xff
      13'h1CDF: dout  = 8'b11111111; // 7391 : 255 - 0xff
      13'h1CE0: dout  = 8'b00000000; // 7392 :   0 - 0x0 -- Background 0xce
      13'h1CE1: dout  = 8'b00000000; // 7393 :   0 - 0x0
      13'h1CE2: dout  = 8'b00000000; // 7394 :   0 - 0x0
      13'h1CE3: dout  = 8'b00000000; // 7395 :   0 - 0x0
      13'h1CE4: dout  = 8'b00000000; // 7396 :   0 - 0x0
      13'h1CE5: dout  = 8'b00000000; // 7397 :   0 - 0x0
      13'h1CE6: dout  = 8'b01111110; // 7398 : 126 - 0x7e
      13'h1CE7: dout  = 8'b00111100; // 7399 :  60 - 0x3c
      13'h1CE8: dout  = 8'b00111100; // 7400 :  60 - 0x3c
      13'h1CE9: dout  = 8'b01111110; // 7401 : 126 - 0x7e
      13'h1CEA: dout  = 8'b01111110; // 7402 : 126 - 0x7e
      13'h1CEB: dout  = 8'b11111111; // 7403 : 255 - 0xff
      13'h1CEC: dout  = 8'b11111111; // 7404 : 255 - 0xff
      13'h1CED: dout  = 8'b11111111; // 7405 : 255 - 0xff
      13'h1CEE: dout  = 8'b01000010; // 7406 :  66 - 0x42
      13'h1CEF: dout  = 8'b00000000; // 7407 :   0 - 0x0
      13'h1CF0: dout  = 8'b00111100; // 7408 :  60 - 0x3c -- Background 0xcf
      13'h1CF1: dout  = 8'b01000010; // 7409 :  66 - 0x42
      13'h1CF2: dout  = 8'b10011001; // 7410 : 153 - 0x99
      13'h1CF3: dout  = 8'b10100001; // 7411 : 161 - 0xa1
      13'h1CF4: dout  = 8'b10100001; // 7412 : 161 - 0xa1
      13'h1CF5: dout  = 8'b10011001; // 7413 : 153 - 0x99
      13'h1CF6: dout  = 8'b01000010; // 7414 :  66 - 0x42
      13'h1CF7: dout  = 8'b00111100; // 7415 :  60 - 0x3c
      13'h1CF8: dout  = 8'b00000000; // 7416 :   0 - 0x0
      13'h1CF9: dout  = 8'b00000000; // 7417 :   0 - 0x0
      13'h1CFA: dout  = 8'b00000000; // 7418 :   0 - 0x0
      13'h1CFB: dout  = 8'b00000000; // 7419 :   0 - 0x0
      13'h1CFC: dout  = 8'b00000000; // 7420 :   0 - 0x0
      13'h1CFD: dout  = 8'b00000000; // 7421 :   0 - 0x0
      13'h1CFE: dout  = 8'b00000000; // 7422 :   0 - 0x0
      13'h1CFF: dout  = 8'b00000000; // 7423 :   0 - 0x0
      13'h1D00: dout  = 8'b00001111; // 7424 :  15 - 0xf -- Background 0xd0
      13'h1D01: dout  = 8'b00011111; // 7425 :  31 - 0x1f
      13'h1D02: dout  = 8'b00011111; // 7426 :  31 - 0x1f
      13'h1D03: dout  = 8'b00111111; // 7427 :  63 - 0x3f
      13'h1D04: dout  = 8'b00111111; // 7428 :  63 - 0x3f
      13'h1D05: dout  = 8'b01111111; // 7429 : 127 - 0x7f
      13'h1D06: dout  = 8'b01111111; // 7430 : 127 - 0x7f
      13'h1D07: dout  = 8'b01111111; // 7431 : 127 - 0x7f
      13'h1D08: dout  = 8'b11110000; // 7432 : 240 - 0xf0
      13'h1D09: dout  = 8'b11100000; // 7433 : 224 - 0xe0
      13'h1D0A: dout  = 8'b11100000; // 7434 : 224 - 0xe0
      13'h1D0B: dout  = 8'b11000000; // 7435 : 192 - 0xc0
      13'h1D0C: dout  = 8'b11000000; // 7436 : 192 - 0xc0
      13'h1D0D: dout  = 8'b10000000; // 7437 : 128 - 0x80
      13'h1D0E: dout  = 8'b10000000; // 7438 : 128 - 0x80
      13'h1D0F: dout  = 8'b10000000; // 7439 : 128 - 0x80
      13'h1D10: dout  = 8'b11110000; // 7440 : 240 - 0xf0 -- Background 0xd1
      13'h1D11: dout  = 8'b11111000; // 7441 : 248 - 0xf8
      13'h1D12: dout  = 8'b11111000; // 7442 : 248 - 0xf8
      13'h1D13: dout  = 8'b11111100; // 7443 : 252 - 0xfc
      13'h1D14: dout  = 8'b11111100; // 7444 : 252 - 0xfc
      13'h1D15: dout  = 8'b11111110; // 7445 : 254 - 0xfe
      13'h1D16: dout  = 8'b11111110; // 7446 : 254 - 0xfe
      13'h1D17: dout  = 8'b11111110; // 7447 : 254 - 0xfe
      13'h1D18: dout  = 8'b00001111; // 7448 :  15 - 0xf
      13'h1D19: dout  = 8'b00000111; // 7449 :   7 - 0x7
      13'h1D1A: dout  = 8'b00000111; // 7450 :   7 - 0x7
      13'h1D1B: dout  = 8'b00000011; // 7451 :   3 - 0x3
      13'h1D1C: dout  = 8'b00000011; // 7452 :   3 - 0x3
      13'h1D1D: dout  = 8'b00000001; // 7453 :   1 - 0x1
      13'h1D1E: dout  = 8'b00000001; // 7454 :   1 - 0x1
      13'h1D1F: dout  = 8'b00000001; // 7455 :   1 - 0x1
      13'h1D20: dout  = 8'b01111111; // 7456 : 127 - 0x7f -- Background 0xd2
      13'h1D21: dout  = 8'b01111111; // 7457 : 127 - 0x7f
      13'h1D22: dout  = 8'b00111111; // 7458 :  63 - 0x3f
      13'h1D23: dout  = 8'b00111111; // 7459 :  63 - 0x3f
      13'h1D24: dout  = 8'b00111111; // 7460 :  63 - 0x3f
      13'h1D25: dout  = 8'b00111111; // 7461 :  63 - 0x3f
      13'h1D26: dout  = 8'b00011111; // 7462 :  31 - 0x1f
      13'h1D27: dout  = 8'b00011111; // 7463 :  31 - 0x1f
      13'h1D28: dout  = 8'b10000000; // 7464 : 128 - 0x80
      13'h1D29: dout  = 8'b10000000; // 7465 : 128 - 0x80
      13'h1D2A: dout  = 8'b11000000; // 7466 : 192 - 0xc0
      13'h1D2B: dout  = 8'b11000000; // 7467 : 192 - 0xc0
      13'h1D2C: dout  = 8'b11100000; // 7468 : 224 - 0xe0
      13'h1D2D: dout  = 8'b11111000; // 7469 : 248 - 0xf8
      13'h1D2E: dout  = 8'b11111110; // 7470 : 254 - 0xfe
      13'h1D2F: dout  = 8'b11111111; // 7471 : 255 - 0xff
      13'h1D30: dout  = 8'b11111110; // 7472 : 254 - 0xfe -- Background 0xd3
      13'h1D31: dout  = 8'b11111111; // 7473 : 255 - 0xff
      13'h1D32: dout  = 8'b11111111; // 7474 : 255 - 0xff
      13'h1D33: dout  = 8'b11111111; // 7475 : 255 - 0xff
      13'h1D34: dout  = 8'b11111100; // 7476 : 252 - 0xfc
      13'h1D35: dout  = 8'b11111100; // 7477 : 252 - 0xfc
      13'h1D36: dout  = 8'b11111110; // 7478 : 254 - 0xfe
      13'h1D37: dout  = 8'b11111110; // 7479 : 254 - 0xfe
      13'h1D38: dout  = 8'b11111111; // 7480 : 255 - 0xff
      13'h1D39: dout  = 8'b01111111; // 7481 : 127 - 0x7f
      13'h1D3A: dout  = 8'b00011111; // 7482 :  31 - 0x1f
      13'h1D3B: dout  = 8'b00000111; // 7483 :   7 - 0x7
      13'h1D3C: dout  = 8'b00000011; // 7484 :   3 - 0x3
      13'h1D3D: dout  = 8'b00000011; // 7485 :   3 - 0x3
      13'h1D3E: dout  = 8'b00000001; // 7486 :   1 - 0x1
      13'h1D3F: dout  = 8'b10000001; // 7487 : 129 - 0x81
      13'h1D40: dout  = 8'b01111111; // 7488 : 127 - 0x7f -- Background 0xd4
      13'h1D41: dout  = 8'b01111111; // 7489 : 127 - 0x7f
      13'h1D42: dout  = 8'b01111111; // 7490 : 127 - 0x7f
      13'h1D43: dout  = 8'b00111111; // 7491 :  63 - 0x3f
      13'h1D44: dout  = 8'b00111111; // 7492 :  63 - 0x3f
      13'h1D45: dout  = 8'b00111111; // 7493 :  63 - 0x3f
      13'h1D46: dout  = 8'b00111111; // 7494 :  63 - 0x3f
      13'h1D47: dout  = 8'b00011111; // 7495 :  31 - 0x1f
      13'h1D48: dout  = 8'b10000000; // 7496 : 128 - 0x80
      13'h1D49: dout  = 8'b10000000; // 7497 : 128 - 0x80
      13'h1D4A: dout  = 8'b10000000; // 7498 : 128 - 0x80
      13'h1D4B: dout  = 8'b11000000; // 7499 : 192 - 0xc0
      13'h1D4C: dout  = 8'b11000000; // 7500 : 192 - 0xc0
      13'h1D4D: dout  = 8'b11100000; // 7501 : 224 - 0xe0
      13'h1D4E: dout  = 8'b11100000; // 7502 : 224 - 0xe0
      13'h1D4F: dout  = 8'b11110000; // 7503 : 240 - 0xf0
      13'h1D50: dout  = 8'b11111110; // 7504 : 254 - 0xfe -- Background 0xd5
      13'h1D51: dout  = 8'b11111110; // 7505 : 254 - 0xfe
      13'h1D52: dout  = 8'b11111111; // 7506 : 255 - 0xff
      13'h1D53: dout  = 8'b11111111; // 7507 : 255 - 0xff
      13'h1D54: dout  = 8'b11111111; // 7508 : 255 - 0xff
      13'h1D55: dout  = 8'b11111111; // 7509 : 255 - 0xff
      13'h1D56: dout  = 8'b11111111; // 7510 : 255 - 0xff
      13'h1D57: dout  = 8'b11111110; // 7511 : 254 - 0xfe
      13'h1D58: dout  = 8'b00000001; // 7512 :   1 - 0x1
      13'h1D59: dout  = 8'b00000001; // 7513 :   1 - 0x1
      13'h1D5A: dout  = 8'b00000001; // 7514 :   1 - 0x1
      13'h1D5B: dout  = 8'b00000011; // 7515 :   3 - 0x3
      13'h1D5C: dout  = 8'b00000011; // 7516 :   3 - 0x3
      13'h1D5D: dout  = 8'b00000111; // 7517 :   7 - 0x7
      13'h1D5E: dout  = 8'b00000111; // 7518 :   7 - 0x7
      13'h1D5F: dout  = 8'b00001111; // 7519 :  15 - 0xf
      13'h1D60: dout  = 8'b00011111; // 7520 :  31 - 0x1f -- Background 0xd6
      13'h1D61: dout  = 8'b00001111; // 7521 :  15 - 0xf
      13'h1D62: dout  = 8'b00001111; // 7522 :  15 - 0xf
      13'h1D63: dout  = 8'b00000111; // 7523 :   7 - 0x7
      13'h1D64: dout  = 8'b00000000; // 7524 :   0 - 0x0
      13'h1D65: dout  = 8'b00000000; // 7525 :   0 - 0x0
      13'h1D66: dout  = 8'b00000000; // 7526 :   0 - 0x0
      13'h1D67: dout  = 8'b00000000; // 7527 :   0 - 0x0
      13'h1D68: dout  = 8'b11111111; // 7528 : 255 - 0xff
      13'h1D69: dout  = 8'b11111111; // 7529 : 255 - 0xff
      13'h1D6A: dout  = 8'b11111111; // 7530 : 255 - 0xff
      13'h1D6B: dout  = 8'b11111111; // 7531 : 255 - 0xff
      13'h1D6C: dout  = 8'b11111111; // 7532 : 255 - 0xff
      13'h1D6D: dout  = 8'b11111111; // 7533 : 255 - 0xff
      13'h1D6E: dout  = 8'b11111111; // 7534 : 255 - 0xff
      13'h1D6F: dout  = 8'b11111111; // 7535 : 255 - 0xff
      13'h1D70: dout  = 8'b11111110; // 7536 : 254 - 0xfe -- Background 0xd7
      13'h1D71: dout  = 8'b11111100; // 7537 : 252 - 0xfc
      13'h1D72: dout  = 8'b11111100; // 7538 : 252 - 0xfc
      13'h1D73: dout  = 8'b11111000; // 7539 : 248 - 0xf8
      13'h1D74: dout  = 8'b00000000; // 7540 :   0 - 0x0
      13'h1D75: dout  = 8'b00000000; // 7541 :   0 - 0x0
      13'h1D76: dout  = 8'b00000000; // 7542 :   0 - 0x0
      13'h1D77: dout  = 8'b00000000; // 7543 :   0 - 0x0
      13'h1D78: dout  = 8'b11111111; // 7544 : 255 - 0xff
      13'h1D79: dout  = 8'b11111111; // 7545 : 255 - 0xff
      13'h1D7A: dout  = 8'b11111111; // 7546 : 255 - 0xff
      13'h1D7B: dout  = 8'b11111111; // 7547 : 255 - 0xff
      13'h1D7C: dout  = 8'b11111111; // 7548 : 255 - 0xff
      13'h1D7D: dout  = 8'b11111111; // 7549 : 255 - 0xff
      13'h1D7E: dout  = 8'b11111111; // 7550 : 255 - 0xff
      13'h1D7F: dout  = 8'b11111111; // 7551 : 255 - 0xff
      13'h1D80: dout  = 8'b01111110; // 7552 : 126 - 0x7e -- Background 0xd8
      13'h1D81: dout  = 8'b01111110; // 7553 : 126 - 0x7e
      13'h1D82: dout  = 8'b01111110; // 7554 : 126 - 0x7e
      13'h1D83: dout  = 8'b01111110; // 7555 : 126 - 0x7e
      13'h1D84: dout  = 8'b01111111; // 7556 : 127 - 0x7f
      13'h1D85: dout  = 8'b01111111; // 7557 : 127 - 0x7f
      13'h1D86: dout  = 8'b01111111; // 7558 : 127 - 0x7f
      13'h1D87: dout  = 8'b01111111; // 7559 : 127 - 0x7f
      13'h1D88: dout  = 8'b10000001; // 7560 : 129 - 0x81
      13'h1D89: dout  = 8'b10000001; // 7561 : 129 - 0x81
      13'h1D8A: dout  = 8'b10000001; // 7562 : 129 - 0x81
      13'h1D8B: dout  = 8'b10000001; // 7563 : 129 - 0x81
      13'h1D8C: dout  = 8'b10000001; // 7564 : 129 - 0x81
      13'h1D8D: dout  = 8'b10000001; // 7565 : 129 - 0x81
      13'h1D8E: dout  = 8'b10000001; // 7566 : 129 - 0x81
      13'h1D8F: dout  = 8'b10000001; // 7567 : 129 - 0x81
      13'h1D90: dout  = 8'b11111111; // 7568 : 255 - 0xff -- Background 0xd9
      13'h1D91: dout  = 8'b11111111; // 7569 : 255 - 0xff
      13'h1D92: dout  = 8'b11111111; // 7570 : 255 - 0xff
      13'h1D93: dout  = 8'b11111111; // 7571 : 255 - 0xff
      13'h1D94: dout  = 8'b11111111; // 7572 : 255 - 0xff
      13'h1D95: dout  = 8'b11111111; // 7573 : 255 - 0xff
      13'h1D96: dout  = 8'b11111111; // 7574 : 255 - 0xff
      13'h1D97: dout  = 8'b11111110; // 7575 : 254 - 0xfe
      13'h1D98: dout  = 8'b00000001; // 7576 :   1 - 0x1
      13'h1D99: dout  = 8'b00000001; // 7577 :   1 - 0x1
      13'h1D9A: dout  = 8'b00000001; // 7578 :   1 - 0x1
      13'h1D9B: dout  = 8'b00000011; // 7579 :   3 - 0x3
      13'h1D9C: dout  = 8'b00000011; // 7580 :   3 - 0x3
      13'h1D9D: dout  = 8'b00000111; // 7581 :   7 - 0x7
      13'h1D9E: dout  = 8'b00000111; // 7582 :   7 - 0x7
      13'h1D9F: dout  = 8'b00001111; // 7583 :  15 - 0xf
      13'h1DA0: dout  = 8'b11111110; // 7584 : 254 - 0xfe -- Background 0xda
      13'h1DA1: dout  = 8'b11111110; // 7585 : 254 - 0xfe
      13'h1DA2: dout  = 8'b11111110; // 7586 : 254 - 0xfe
      13'h1DA3: dout  = 8'b11111110; // 7587 : 254 - 0xfe
      13'h1DA4: dout  = 8'b11111111; // 7588 : 255 - 0xff
      13'h1DA5: dout  = 8'b11111111; // 7589 : 255 - 0xff
      13'h1DA6: dout  = 8'b11111111; // 7590 : 255 - 0xff
      13'h1DA7: dout  = 8'b11111111; // 7591 : 255 - 0xff
      13'h1DA8: dout  = 8'b00000001; // 7592 :   1 - 0x1
      13'h1DA9: dout  = 8'b00000001; // 7593 :   1 - 0x1
      13'h1DAA: dout  = 8'b00000001; // 7594 :   1 - 0x1
      13'h1DAB: dout  = 8'b00000001; // 7595 :   1 - 0x1
      13'h1DAC: dout  = 8'b00000001; // 7596 :   1 - 0x1
      13'h1DAD: dout  = 8'b00000001; // 7597 :   1 - 0x1
      13'h1DAE: dout  = 8'b00000001; // 7598 :   1 - 0x1
      13'h1DAF: dout  = 8'b00000001; // 7599 :   1 - 0x1
      13'h1DB0: dout  = 8'b01111111; // 7600 : 127 - 0x7f -- Background 0xdb
      13'h1DB1: dout  = 8'b01111111; // 7601 : 127 - 0x7f
      13'h1DB2: dout  = 8'b01111111; // 7602 : 127 - 0x7f
      13'h1DB3: dout  = 8'b01111111; // 7603 : 127 - 0x7f
      13'h1DB4: dout  = 8'b01111111; // 7604 : 127 - 0x7f
      13'h1DB5: dout  = 8'b01111111; // 7605 : 127 - 0x7f
      13'h1DB6: dout  = 8'b01111111; // 7606 : 127 - 0x7f
      13'h1DB7: dout  = 8'b01111111; // 7607 : 127 - 0x7f
      13'h1DB8: dout  = 8'b10000001; // 7608 : 129 - 0x81
      13'h1DB9: dout  = 8'b10000001; // 7609 : 129 - 0x81
      13'h1DBA: dout  = 8'b10000001; // 7610 : 129 - 0x81
      13'h1DBB: dout  = 8'b10000001; // 7611 : 129 - 0x81
      13'h1DBC: dout  = 8'b10000001; // 7612 : 129 - 0x81
      13'h1DBD: dout  = 8'b10000001; // 7613 : 129 - 0x81
      13'h1DBE: dout  = 8'b10000001; // 7614 : 129 - 0x81
      13'h1DBF: dout  = 8'b10000001; // 7615 : 129 - 0x81
      13'h1DC0: dout  = 8'b11111111; // 7616 : 255 - 0xff -- Background 0xdc
      13'h1DC1: dout  = 8'b11111111; // 7617 : 255 - 0xff
      13'h1DC2: dout  = 8'b11111111; // 7618 : 255 - 0xff
      13'h1DC3: dout  = 8'b11111111; // 7619 : 255 - 0xff
      13'h1DC4: dout  = 8'b11111100; // 7620 : 252 - 0xfc
      13'h1DC5: dout  = 8'b11111110; // 7621 : 254 - 0xfe
      13'h1DC6: dout  = 8'b11111110; // 7622 : 254 - 0xfe
      13'h1DC7: dout  = 8'b01111110; // 7623 : 126 - 0x7e
      13'h1DC8: dout  = 8'b11111111; // 7624 : 255 - 0xff
      13'h1DC9: dout  = 8'b00000011; // 7625 :   3 - 0x3
      13'h1DCA: dout  = 8'b00000011; // 7626 :   3 - 0x3
      13'h1DCB: dout  = 8'b00000011; // 7627 :   3 - 0x3
      13'h1DCC: dout  = 8'b00000011; // 7628 :   3 - 0x3
      13'h1DCD: dout  = 8'b00000011; // 7629 :   3 - 0x3
      13'h1DCE: dout  = 8'b00000011; // 7630 :   3 - 0x3
      13'h1DCF: dout  = 8'b11111111; // 7631 : 255 - 0xff
      13'h1DD0: dout  = 8'b11111111; // 7632 : 255 - 0xff -- Background 0xdd
      13'h1DD1: dout  = 8'b11111111; // 7633 : 255 - 0xff
      13'h1DD2: dout  = 8'b11111111; // 7634 : 255 - 0xff
      13'h1DD3: dout  = 8'b11111111; // 7635 : 255 - 0xff
      13'h1DD4: dout  = 8'b00000000; // 7636 :   0 - 0x0
      13'h1DD5: dout  = 8'b00000000; // 7637 :   0 - 0x0
      13'h1DD6: dout  = 8'b00000000; // 7638 :   0 - 0x0
      13'h1DD7: dout  = 8'b00000000; // 7639 :   0 - 0x0
      13'h1DD8: dout  = 8'b11111111; // 7640 : 255 - 0xff
      13'h1DD9: dout  = 8'b11111111; // 7641 : 255 - 0xff
      13'h1DDA: dout  = 8'b11111111; // 7642 : 255 - 0xff
      13'h1DDB: dout  = 8'b11111111; // 7643 : 255 - 0xff
      13'h1DDC: dout  = 8'b11111111; // 7644 : 255 - 0xff
      13'h1DDD: dout  = 8'b11111111; // 7645 : 255 - 0xff
      13'h1DDE: dout  = 8'b11111111; // 7646 : 255 - 0xff
      13'h1DDF: dout  = 8'b11111111; // 7647 : 255 - 0xff
      13'h1DE0: dout  = 8'b01111111; // 7648 : 127 - 0x7f -- Background 0xde
      13'h1DE1: dout  = 8'b01111111; // 7649 : 127 - 0x7f
      13'h1DE2: dout  = 8'b01111111; // 7650 : 127 - 0x7f
      13'h1DE3: dout  = 8'b01111111; // 7651 : 127 - 0x7f
      13'h1DE4: dout  = 8'b01111111; // 7652 : 127 - 0x7f
      13'h1DE5: dout  = 8'b01111111; // 7653 : 127 - 0x7f
      13'h1DE6: dout  = 8'b01111111; // 7654 : 127 - 0x7f
      13'h1DE7: dout  = 8'b01111111; // 7655 : 127 - 0x7f
      13'h1DE8: dout  = 8'b10000000; // 7656 : 128 - 0x80
      13'h1DE9: dout  = 8'b10000000; // 7657 : 128 - 0x80
      13'h1DEA: dout  = 8'b10000000; // 7658 : 128 - 0x80
      13'h1DEB: dout  = 8'b10000000; // 7659 : 128 - 0x80
      13'h1DEC: dout  = 8'b10000000; // 7660 : 128 - 0x80
      13'h1DED: dout  = 8'b10000000; // 7661 : 128 - 0x80
      13'h1DEE: dout  = 8'b10000000; // 7662 : 128 - 0x80
      13'h1DEF: dout  = 8'b10000000; // 7663 : 128 - 0x80
      13'h1DF0: dout  = 8'b11111111; // 7664 : 255 - 0xff -- Background 0xdf
      13'h1DF1: dout  = 8'b11111111; // 7665 : 255 - 0xff
      13'h1DF2: dout  = 8'b11111111; // 7666 : 255 - 0xff
      13'h1DF3: dout  = 8'b11111111; // 7667 : 255 - 0xff
      13'h1DF4: dout  = 8'b11111111; // 7668 : 255 - 0xff
      13'h1DF5: dout  = 8'b11111111; // 7669 : 255 - 0xff
      13'h1DF6: dout  = 8'b11111111; // 7670 : 255 - 0xff
      13'h1DF7: dout  = 8'b11111110; // 7671 : 254 - 0xfe
      13'h1DF8: dout  = 8'b00000001; // 7672 :   1 - 0x1
      13'h1DF9: dout  = 8'b00000001; // 7673 :   1 - 0x1
      13'h1DFA: dout  = 8'b00000001; // 7674 :   1 - 0x1
      13'h1DFB: dout  = 8'b00000011; // 7675 :   3 - 0x3
      13'h1DFC: dout  = 8'b00000111; // 7676 :   7 - 0x7
      13'h1DFD: dout  = 8'b00000011; // 7677 :   3 - 0x3
      13'h1DFE: dout  = 8'b00000001; // 7678 :   1 - 0x1
      13'h1DFF: dout  = 8'b00000001; // 7679 :   1 - 0x1
      13'h1E00: dout  = 8'b01111110; // 7680 : 126 - 0x7e -- Background 0xe0
      13'h1E01: dout  = 8'b01111110; // 7681 : 126 - 0x7e
      13'h1E02: dout  = 8'b01111111; // 7682 : 127 - 0x7f
      13'h1E03: dout  = 8'b01111111; // 7683 : 127 - 0x7f
      13'h1E04: dout  = 8'b01111111; // 7684 : 127 - 0x7f
      13'h1E05: dout  = 8'b01111111; // 7685 : 127 - 0x7f
      13'h1E06: dout  = 8'b01111111; // 7686 : 127 - 0x7f
      13'h1E07: dout  = 8'b01111111; // 7687 : 127 - 0x7f
      13'h1E08: dout  = 8'b10000001; // 7688 : 129 - 0x81
      13'h1E09: dout  = 8'b10000001; // 7689 : 129 - 0x81
      13'h1E0A: dout  = 8'b10000001; // 7690 : 129 - 0x81
      13'h1E0B: dout  = 8'b10000001; // 7691 : 129 - 0x81
      13'h1E0C: dout  = 8'b10000001; // 7692 : 129 - 0x81
      13'h1E0D: dout  = 8'b10000001; // 7693 : 129 - 0x81
      13'h1E0E: dout  = 8'b10000001; // 7694 : 129 - 0x81
      13'h1E0F: dout  = 8'b10000001; // 7695 : 129 - 0x81
      13'h1E10: dout  = 8'b00111111; // 7696 :  63 - 0x3f -- Background 0xe1
      13'h1E11: dout  = 8'b00111111; // 7697 :  63 - 0x3f
      13'h1E12: dout  = 8'b00111111; // 7698 :  63 - 0x3f
      13'h1E13: dout  = 8'b00111111; // 7699 :  63 - 0x3f
      13'h1E14: dout  = 8'b00000000; // 7700 :   0 - 0x0
      13'h1E15: dout  = 8'b00000000; // 7701 :   0 - 0x0
      13'h1E16: dout  = 8'b00000000; // 7702 :   0 - 0x0
      13'h1E17: dout  = 8'b00000000; // 7703 :   0 - 0x0
      13'h1E18: dout  = 8'b11111111; // 7704 : 255 - 0xff
      13'h1E19: dout  = 8'b11111111; // 7705 : 255 - 0xff
      13'h1E1A: dout  = 8'b11111111; // 7706 : 255 - 0xff
      13'h1E1B: dout  = 8'b11111111; // 7707 : 255 - 0xff
      13'h1E1C: dout  = 8'b11111111; // 7708 : 255 - 0xff
      13'h1E1D: dout  = 8'b11111111; // 7709 : 255 - 0xff
      13'h1E1E: dout  = 8'b11111111; // 7710 : 255 - 0xff
      13'h1E1F: dout  = 8'b11111111; // 7711 : 255 - 0xff
      13'h1E20: dout  = 8'b01111110; // 7712 : 126 - 0x7e -- Background 0xe2
      13'h1E21: dout  = 8'b01111100; // 7713 : 124 - 0x7c
      13'h1E22: dout  = 8'b01111100; // 7714 : 124 - 0x7c
      13'h1E23: dout  = 8'b01111000; // 7715 : 120 - 0x78
      13'h1E24: dout  = 8'b00000000; // 7716 :   0 - 0x0
      13'h1E25: dout  = 8'b00000000; // 7717 :   0 - 0x0
      13'h1E26: dout  = 8'b00000000; // 7718 :   0 - 0x0
      13'h1E27: dout  = 8'b00000000; // 7719 :   0 - 0x0
      13'h1E28: dout  = 8'b11111111; // 7720 : 255 - 0xff
      13'h1E29: dout  = 8'b11111111; // 7721 : 255 - 0xff
      13'h1E2A: dout  = 8'b11111111; // 7722 : 255 - 0xff
      13'h1E2B: dout  = 8'b11111111; // 7723 : 255 - 0xff
      13'h1E2C: dout  = 8'b11111111; // 7724 : 255 - 0xff
      13'h1E2D: dout  = 8'b11111111; // 7725 : 255 - 0xff
      13'h1E2E: dout  = 8'b11111111; // 7726 : 255 - 0xff
      13'h1E2F: dout  = 8'b11111111; // 7727 : 255 - 0xff
      13'h1E30: dout  = 8'b11111110; // 7728 : 254 - 0xfe -- Background 0xe3
      13'h1E31: dout  = 8'b11111110; // 7729 : 254 - 0xfe
      13'h1E32: dout  = 8'b11111111; // 7730 : 255 - 0xff
      13'h1E33: dout  = 8'b11111111; // 7731 : 255 - 0xff
      13'h1E34: dout  = 8'b01111111; // 7732 : 127 - 0x7f
      13'h1E35: dout  = 8'b01111111; // 7733 : 127 - 0x7f
      13'h1E36: dout  = 8'b01111111; // 7734 : 127 - 0x7f
      13'h1E37: dout  = 8'b01111111; // 7735 : 127 - 0x7f
      13'h1E38: dout  = 8'b10000001; // 7736 : 129 - 0x81
      13'h1E39: dout  = 8'b10000001; // 7737 : 129 - 0x81
      13'h1E3A: dout  = 8'b10000001; // 7738 : 129 - 0x81
      13'h1E3B: dout  = 8'b10000001; // 7739 : 129 - 0x81
      13'h1E3C: dout  = 8'b10000001; // 7740 : 129 - 0x81
      13'h1E3D: dout  = 8'b10000001; // 7741 : 129 - 0x81
      13'h1E3E: dout  = 8'b10000001; // 7742 : 129 - 0x81
      13'h1E3F: dout  = 8'b10000001; // 7743 : 129 - 0x81
      13'h1E40: dout  = 8'b01111111; // 7744 : 127 - 0x7f -- Background 0xe4
      13'h1E41: dout  = 8'b01111111; // 7745 : 127 - 0x7f
      13'h1E42: dout  = 8'b00111111; // 7746 :  63 - 0x3f
      13'h1E43: dout  = 8'b00111111; // 7747 :  63 - 0x3f
      13'h1E44: dout  = 8'b00111111; // 7748 :  63 - 0x3f
      13'h1E45: dout  = 8'b00111111; // 7749 :  63 - 0x3f
      13'h1E46: dout  = 8'b00011111; // 7750 :  31 - 0x1f
      13'h1E47: dout  = 8'b00011111; // 7751 :  31 - 0x1f
      13'h1E48: dout  = 8'b10000000; // 7752 : 128 - 0x80
      13'h1E49: dout  = 8'b10000000; // 7753 : 128 - 0x80
      13'h1E4A: dout  = 8'b11000000; // 7754 : 192 - 0xc0
      13'h1E4B: dout  = 8'b11000000; // 7755 : 192 - 0xc0
      13'h1E4C: dout  = 8'b11100000; // 7756 : 224 - 0xe0
      13'h1E4D: dout  = 8'b11111000; // 7757 : 248 - 0xf8
      13'h1E4E: dout  = 8'b11111110; // 7758 : 254 - 0xfe
      13'h1E4F: dout  = 8'b11111111; // 7759 : 255 - 0xff
      13'h1E50: dout  = 8'b00111111; // 7760 :  63 - 0x3f -- Background 0xe5
      13'h1E51: dout  = 8'b10111111; // 7761 : 191 - 0xbf
      13'h1E52: dout  = 8'b11111111; // 7762 : 255 - 0xff
      13'h1E53: dout  = 8'b11111111; // 7763 : 255 - 0xff
      13'h1E54: dout  = 8'b11111100; // 7764 : 252 - 0xfc
      13'h1E55: dout  = 8'b11111100; // 7765 : 252 - 0xfc
      13'h1E56: dout  = 8'b11111110; // 7766 : 254 - 0xfe
      13'h1E57: dout  = 8'b11111110; // 7767 : 254 - 0xfe
      13'h1E58: dout  = 8'b11111111; // 7768 : 255 - 0xff
      13'h1E59: dout  = 8'b01111111; // 7769 : 127 - 0x7f
      13'h1E5A: dout  = 8'b00011111; // 7770 :  31 - 0x1f
      13'h1E5B: dout  = 8'b00000111; // 7771 :   7 - 0x7
      13'h1E5C: dout  = 8'b00000011; // 7772 :   3 - 0x3
      13'h1E5D: dout  = 8'b00000011; // 7773 :   3 - 0x3
      13'h1E5E: dout  = 8'b00000001; // 7774 :   1 - 0x1
      13'h1E5F: dout  = 8'b10000001; // 7775 : 129 - 0x81
      13'h1E60: dout  = 8'b01111111; // 7776 : 127 - 0x7f -- Background 0xe6
      13'h1E61: dout  = 8'b01111111; // 7777 : 127 - 0x7f
      13'h1E62: dout  = 8'b01111110; // 7778 : 126 - 0x7e
      13'h1E63: dout  = 8'b01111110; // 7779 : 126 - 0x7e
      13'h1E64: dout  = 8'b01111111; // 7780 : 127 - 0x7f
      13'h1E65: dout  = 8'b01111111; // 7781 : 127 - 0x7f
      13'h1E66: dout  = 8'b01111111; // 7782 : 127 - 0x7f
      13'h1E67: dout  = 8'b01111111; // 7783 : 127 - 0x7f
      13'h1E68: dout  = 8'b10000001; // 7784 : 129 - 0x81
      13'h1E69: dout  = 8'b10000001; // 7785 : 129 - 0x81
      13'h1E6A: dout  = 8'b10000001; // 7786 : 129 - 0x81
      13'h1E6B: dout  = 8'b10000001; // 7787 : 129 - 0x81
      13'h1E6C: dout  = 8'b10000001; // 7788 : 129 - 0x81
      13'h1E6D: dout  = 8'b10000001; // 7789 : 129 - 0x81
      13'h1E6E: dout  = 8'b10000001; // 7790 : 129 - 0x81
      13'h1E6F: dout  = 8'b10000001; // 7791 : 129 - 0x81
      13'h1E70: dout  = 8'b01111110; // 7792 : 126 - 0x7e -- Background 0xe7
      13'h1E71: dout  = 8'b01111110; // 7793 : 126 - 0x7e
      13'h1E72: dout  = 8'b01111110; // 7794 : 126 - 0x7e
      13'h1E73: dout  = 8'b01111110; // 7795 : 126 - 0x7e
      13'h1E74: dout  = 8'b01111111; // 7796 : 127 - 0x7f
      13'h1E75: dout  = 8'b01111111; // 7797 : 127 - 0x7f
      13'h1E76: dout  = 8'b01111111; // 7798 : 127 - 0x7f
      13'h1E77: dout  = 8'b01111111; // 7799 : 127 - 0x7f
      13'h1E78: dout  = 8'b10000001; // 7800 : 129 - 0x81
      13'h1E79: dout  = 8'b10000001; // 7801 : 129 - 0x81
      13'h1E7A: dout  = 8'b10000001; // 7802 : 129 - 0x81
      13'h1E7B: dout  = 8'b10000001; // 7803 : 129 - 0x81
      13'h1E7C: dout  = 8'b10000001; // 7804 : 129 - 0x81
      13'h1E7D: dout  = 8'b10000001; // 7805 : 129 - 0x81
      13'h1E7E: dout  = 8'b10000001; // 7806 : 129 - 0x81
      13'h1E7F: dout  = 8'b10000001; // 7807 : 129 - 0x81
      13'h1E80: dout  = 8'b10000001; // 7808 : 129 - 0x81 -- Background 0xe8
      13'h1E81: dout  = 8'b11000011; // 7809 : 195 - 0xc3
      13'h1E82: dout  = 8'b11000011; // 7810 : 195 - 0xc3
      13'h1E83: dout  = 8'b11100111; // 7811 : 231 - 0xe7
      13'h1E84: dout  = 8'b11100111; // 7812 : 231 - 0xe7
      13'h1E85: dout  = 8'b11111111; // 7813 : 255 - 0xff
      13'h1E86: dout  = 8'b11111111; // 7814 : 255 - 0xff
      13'h1E87: dout  = 8'b11111111; // 7815 : 255 - 0xff
      13'h1E88: dout  = 8'b01111110; // 7816 : 126 - 0x7e
      13'h1E89: dout  = 8'b00111100; // 7817 :  60 - 0x3c
      13'h1E8A: dout  = 8'b00111100; // 7818 :  60 - 0x3c
      13'h1E8B: dout  = 8'b00011000; // 7819 :  24 - 0x18
      13'h1E8C: dout  = 8'b00011000; // 7820 :  24 - 0x18
      13'h1E8D: dout  = 8'b00000000; // 7821 :   0 - 0x0
      13'h1E8E: dout  = 8'b00000000; // 7822 :   0 - 0x0
      13'h1E8F: dout  = 8'b00000000; // 7823 :   0 - 0x0
      13'h1E90: dout  = 8'b00001111; // 7824 :  15 - 0xf -- Background 0xe9
      13'h1E91: dout  = 8'b01000011; // 7825 :  67 - 0x43
      13'h1E92: dout  = 8'b01011011; // 7826 :  91 - 0x5b
      13'h1E93: dout  = 8'b01010011; // 7827 :  83 - 0x53
      13'h1E94: dout  = 8'b00110001; // 7828 :  49 - 0x31
      13'h1E95: dout  = 8'b00011001; // 7829 :  25 - 0x19
      13'h1E96: dout  = 8'b00001111; // 7830 :  15 - 0xf
      13'h1E97: dout  = 8'b00000111; // 7831 :   7 - 0x7
      13'h1E98: dout  = 8'b11110010; // 7832 : 242 - 0xf2
      13'h1E99: dout  = 8'b11111110; // 7833 : 254 - 0xfe
      13'h1E9A: dout  = 8'b11111110; // 7834 : 254 - 0xfe
      13'h1E9B: dout  = 8'b11111111; // 7835 : 255 - 0xff
      13'h1E9C: dout  = 8'b11111111; // 7836 : 255 - 0xff
      13'h1E9D: dout  = 8'b11101111; // 7837 : 239 - 0xef
      13'h1E9E: dout  = 8'b11110111; // 7838 : 247 - 0xf7
      13'h1E9F: dout  = 8'b11111000; // 7839 : 248 - 0xf8
      13'h1EA0: dout  = 8'b11000001; // 7840 : 193 - 0xc1 -- Background 0xea
      13'h1EA1: dout  = 8'b11000011; // 7841 : 195 - 0xc3
      13'h1EA2: dout  = 8'b11000110; // 7842 : 198 - 0xc6
      13'h1EA3: dout  = 8'b10000100; // 7843 : 132 - 0x84
      13'h1EA4: dout  = 8'b11111100; // 7844 : 252 - 0xfc
      13'h1EA5: dout  = 8'b11111100; // 7845 : 252 - 0xfc
      13'h1EA6: dout  = 8'b00001110; // 7846 :  14 - 0xe
      13'h1EA7: dout  = 8'b00000010; // 7847 :   2 - 0x2
      13'h1EA8: dout  = 8'b10111111; // 7848 : 191 - 0xbf
      13'h1EA9: dout  = 8'b10111110; // 7849 : 190 - 0xbe
      13'h1EAA: dout  = 8'b10111101; // 7850 : 189 - 0xbd
      13'h1EAB: dout  = 8'b01111011; // 7851 : 123 - 0x7b
      13'h1EAC: dout  = 8'b01111011; // 7852 : 123 - 0x7b
      13'h1EAD: dout  = 8'b00000111; // 7853 :   7 - 0x7
      13'h1EAE: dout  = 8'b11110011; // 7854 : 243 - 0xf3
      13'h1EAF: dout  = 8'b11111101; // 7855 : 253 - 0xfd
      13'h1EB0: dout  = 8'b00010000; // 7856 :  16 - 0x10 -- Background 0xeb
      13'h1EB1: dout  = 8'b00100000; // 7857 :  32 - 0x20
      13'h1EB2: dout  = 8'b00100010; // 7858 :  34 - 0x22
      13'h1EB3: dout  = 8'b10111010; // 7859 : 186 - 0xba
      13'h1EB4: dout  = 8'b11100110; // 7860 : 230 - 0xe6
      13'h1EB5: dout  = 8'b11100001; // 7861 : 225 - 0xe1
      13'h1EB6: dout  = 8'b11000000; // 7862 : 192 - 0xc0
      13'h1EB7: dout  = 8'b11000000; // 7863 : 192 - 0xc0
      13'h1EB8: dout  = 8'b11111111; // 7864 : 255 - 0xff
      13'h1EB9: dout  = 8'b11111111; // 7865 : 255 - 0xff
      13'h1EBA: dout  = 8'b11111111; // 7866 : 255 - 0xff
      13'h1EBB: dout  = 8'b01100111; // 7867 : 103 - 0x67
      13'h1EBC: dout  = 8'b01011001; // 7868 :  89 - 0x59
      13'h1EBD: dout  = 8'b10011110; // 7869 : 158 - 0x9e
      13'h1EBE: dout  = 8'b10111111; // 7870 : 191 - 0xbf
      13'h1EBF: dout  = 8'b10111111; // 7871 : 191 - 0xbf
      13'h1EC0: dout  = 8'b00100000; // 7872 :  32 - 0x20 -- Background 0xec
      13'h1EC1: dout  = 8'b10100110; // 7873 : 166 - 0xa6
      13'h1EC2: dout  = 8'b01010100; // 7874 :  84 - 0x54
      13'h1EC3: dout  = 8'b00100110; // 7875 :  38 - 0x26
      13'h1EC4: dout  = 8'b00100000; // 7876 :  32 - 0x20
      13'h1EC5: dout  = 8'b11000110; // 7877 : 198 - 0xc6
      13'h1EC6: dout  = 8'b01010100; // 7878 :  84 - 0x54
      13'h1EC7: dout  = 8'b00100110; // 7879 :  38 - 0x26
      13'h1EC8: dout  = 8'b00100000; // 7880 :  32 - 0x20
      13'h1EC9: dout  = 8'b11100110; // 7881 : 230 - 0xe6
      13'h1ECA: dout  = 8'b01010100; // 7882 :  84 - 0x54
      13'h1ECB: dout  = 8'b00100110; // 7883 :  38 - 0x26
      13'h1ECC: dout  = 8'b00100001; // 7884 :  33 - 0x21
      13'h1ECD: dout  = 8'b00000110; // 7885 :   6 - 0x6
      13'h1ECE: dout  = 8'b01010100; // 7886 :  84 - 0x54
      13'h1ECF: dout  = 8'b00100110; // 7887 :  38 - 0x26
      13'h1ED0: dout  = 8'b00100000; // 7888 :  32 - 0x20 -- Background 0xed
      13'h1ED1: dout  = 8'b10000101; // 7889 : 133 - 0x85
      13'h1ED2: dout  = 8'b00000001; // 7890 :   1 - 0x1
      13'h1ED3: dout  = 8'b01000100; // 7891 :  68 - 0x44
      13'h1ED4: dout  = 8'b00100000; // 7892 :  32 - 0x20
      13'h1ED5: dout  = 8'b10000110; // 7893 : 134 - 0x86
      13'h1ED6: dout  = 8'b01010100; // 7894 :  84 - 0x54
      13'h1ED7: dout  = 8'b01001000; // 7895 :  72 - 0x48
      13'h1ED8: dout  = 8'b00100000; // 7896 :  32 - 0x20
      13'h1ED9: dout  = 8'b10011010; // 7897 : 154 - 0x9a
      13'h1EDA: dout  = 8'b00000001; // 7898 :   1 - 0x1
      13'h1EDB: dout  = 8'b01001001; // 7899 :  73 - 0x49
      13'h1EDC: dout  = 8'b00100000; // 7900 :  32 - 0x20
      13'h1EDD: dout  = 8'b10100101; // 7901 : 165 - 0xa5
      13'h1EDE: dout  = 8'b11001001; // 7902 : 201 - 0xc9
      13'h1EDF: dout  = 8'b01000110; // 7903 :  70 - 0x46
      13'h1EE0: dout  = 8'b00100000; // 7904 :  32 - 0x20 -- Background 0xee
      13'h1EE1: dout  = 8'b10111010; // 7905 : 186 - 0xba
      13'h1EE2: dout  = 8'b11001001; // 7906 : 201 - 0xc9
      13'h1EE3: dout  = 8'b01001010; // 7907 :  74 - 0x4a
      13'h1EE4: dout  = 8'b00100000; // 7908 :  32 - 0x20
      13'h1EE5: dout  = 8'b10100110; // 7909 : 166 - 0xa6
      13'h1EE6: dout  = 8'b00001010; // 7910 :  10 - 0xa
      13'h1EE7: dout  = 8'b11010000; // 7911 : 208 - 0xd0
      13'h1EE8: dout  = 8'b11010001; // 7912 : 209 - 0xd1
      13'h1EE9: dout  = 8'b11011000; // 7913 : 216 - 0xd8
      13'h1EEA: dout  = 8'b11011000; // 7914 : 216 - 0xd8
      13'h1EEB: dout  = 8'b11011110; // 7915 : 222 - 0xde
      13'h1EEC: dout  = 8'b11010001; // 7916 : 209 - 0xd1
      13'h1EED: dout  = 8'b11010000; // 7917 : 208 - 0xd0
      13'h1EEE: dout  = 8'b11011010; // 7918 : 218 - 0xda
      13'h1EEF: dout  = 8'b11011110; // 7919 : 222 - 0xde
      13'h1EF0: dout  = 8'b11010001; // 7920 : 209 - 0xd1 -- Background 0xef
      13'h1EF1: dout  = 8'b00100000; // 7921 :  32 - 0x20
      13'h1EF2: dout  = 8'b11000110; // 7922 : 198 - 0xc6
      13'h1EF3: dout  = 8'b00001010; // 7923 :  10 - 0xa
      13'h1EF4: dout  = 8'b11010010; // 7924 : 210 - 0xd2
      13'h1EF5: dout  = 8'b11010011; // 7925 : 211 - 0xd3
      13'h1EF6: dout  = 8'b11011011; // 7926 : 219 - 0xdb
      13'h1EF7: dout  = 8'b11011011; // 7927 : 219 - 0xdb
      13'h1EF8: dout  = 8'b11011011; // 7928 : 219 - 0xdb
      13'h1EF9: dout  = 8'b11011001; // 7929 : 217 - 0xd9
      13'h1EFA: dout  = 8'b11011011; // 7930 : 219 - 0xdb
      13'h1EFB: dout  = 8'b11011100; // 7931 : 220 - 0xdc
      13'h1EFC: dout  = 8'b11011011; // 7932 : 219 - 0xdb
      13'h1EFD: dout  = 8'b11011111; // 7933 : 223 - 0xdf
      13'h1EFE: dout  = 8'b00100000; // 7934 :  32 - 0x20
      13'h1EFF: dout  = 8'b11100110; // 7935 : 230 - 0xe6
      13'h1F00: dout  = 8'b00001010; // 7936 :  10 - 0xa -- Background 0xf0
      13'h1F01: dout  = 8'b11010100; // 7937 : 212 - 0xd4
      13'h1F02: dout  = 8'b11010101; // 7938 : 213 - 0xd5
      13'h1F03: dout  = 8'b11010100; // 7939 : 212 - 0xd4
      13'h1F04: dout  = 8'b11011001; // 7940 : 217 - 0xd9
      13'h1F05: dout  = 8'b11011011; // 7941 : 219 - 0xdb
      13'h1F06: dout  = 8'b11100010; // 7942 : 226 - 0xe2
      13'h1F07: dout  = 8'b11010100; // 7943 : 212 - 0xd4
      13'h1F08: dout  = 8'b11011010; // 7944 : 218 - 0xda
      13'h1F09: dout  = 8'b11011011; // 7945 : 219 - 0xdb
      13'h1F0A: dout  = 8'b11100000; // 7946 : 224 - 0xe0
      13'h1F0B: dout  = 8'b00100001; // 7947 :  33 - 0x21
      13'h1F0C: dout  = 8'b00000110; // 7948 :   6 - 0x6
      13'h1F0D: dout  = 8'b00001010; // 7949 :  10 - 0xa
      13'h1F0E: dout  = 8'b11010110; // 7950 : 214 - 0xd6
      13'h1F0F: dout  = 8'b11010111; // 7951 : 215 - 0xd7
      13'h1F10: dout  = 8'b11010110; // 7952 : 214 - 0xd6 -- Background 0xf1
      13'h1F11: dout  = 8'b11010111; // 7953 : 215 - 0xd7
      13'h1F12: dout  = 8'b11100001; // 7954 : 225 - 0xe1
      13'h1F13: dout  = 8'b00100110; // 7955 :  38 - 0x26
      13'h1F14: dout  = 8'b11010110; // 7956 : 214 - 0xd6
      13'h1F15: dout  = 8'b11011101; // 7957 : 221 - 0xdd
      13'h1F16: dout  = 8'b11100001; // 7958 : 225 - 0xe1
      13'h1F17: dout  = 8'b11100001; // 7959 : 225 - 0xe1
      13'h1F18: dout  = 8'b00100001; // 7960 :  33 - 0x21
      13'h1F19: dout  = 8'b00100110; // 7961 :  38 - 0x26
      13'h1F1A: dout  = 8'b00010100; // 7962 :  20 - 0x14
      13'h1F1B: dout  = 8'b11010000; // 7963 : 208 - 0xd0
      13'h1F1C: dout  = 8'b11101000; // 7964 : 232 - 0xe8
      13'h1F1D: dout  = 8'b11010001; // 7965 : 209 - 0xd1
      13'h1F1E: dout  = 8'b11010000; // 7966 : 208 - 0xd0
      13'h1F1F: dout  = 8'b11010001; // 7967 : 209 - 0xd1
      13'h1F20: dout  = 8'b11011110; // 7968 : 222 - 0xde -- Background 0xf2
      13'h1F21: dout  = 8'b11010001; // 7969 : 209 - 0xd1
      13'h1F22: dout  = 8'b11011000; // 7970 : 216 - 0xd8
      13'h1F23: dout  = 8'b11010000; // 7971 : 208 - 0xd0
      13'h1F24: dout  = 8'b11010001; // 7972 : 209 - 0xd1
      13'h1F25: dout  = 8'b00100110; // 7973 :  38 - 0x26
      13'h1F26: dout  = 8'b11011110; // 7974 : 222 - 0xde
      13'h1F27: dout  = 8'b11010001; // 7975 : 209 - 0xd1
      13'h1F28: dout  = 8'b11011110; // 7976 : 222 - 0xde
      13'h1F29: dout  = 8'b11010001; // 7977 : 209 - 0xd1
      13'h1F2A: dout  = 8'b11010000; // 7978 : 208 - 0xd0
      13'h1F2B: dout  = 8'b11010001; // 7979 : 209 - 0xd1
      13'h1F2C: dout  = 8'b11010000; // 7980 : 208 - 0xd0
      13'h1F2D: dout  = 8'b11010001; // 7981 : 209 - 0xd1
      13'h1F2E: dout  = 8'b00100110; // 7982 :  38 - 0x26
      13'h1F2F: dout  = 8'b00100001; // 7983 :  33 - 0x21
      13'h1F30: dout  = 8'b01000110; // 7984 :  70 - 0x46 -- Background 0xf3
      13'h1F31: dout  = 8'b00010100; // 7985 :  20 - 0x14
      13'h1F32: dout  = 8'b11011011; // 7986 : 219 - 0xdb
      13'h1F33: dout  = 8'b01000010; // 7987 :  66 - 0x42
      13'h1F34: dout  = 8'b01000010; // 7988 :  66 - 0x42
      13'h1F35: dout  = 8'b11011011; // 7989 : 219 - 0xdb
      13'h1F36: dout  = 8'b01000010; // 7990 :  66 - 0x42
      13'h1F37: dout  = 8'b11011011; // 7991 : 219 - 0xdb
      13'h1F38: dout  = 8'b01000010; // 7992 :  66 - 0x42
      13'h1F39: dout  = 8'b11011011; // 7993 : 219 - 0xdb
      13'h1F3A: dout  = 8'b11011011; // 7994 : 219 - 0xdb
      13'h1F3B: dout  = 8'b01000010; // 7995 :  66 - 0x42
      13'h1F3C: dout  = 8'b00100110; // 7996 :  38 - 0x26
      13'h1F3D: dout  = 8'b11011011; // 7997 : 219 - 0xdb
      13'h1F3E: dout  = 8'b01000010; // 7998 :  66 - 0x42
      13'h1F3F: dout  = 8'b11011011; // 7999 : 219 - 0xdb
      13'h1F40: dout  = 8'b01000010; // 8000 :  66 - 0x42 -- Background 0xf4
      13'h1F41: dout  = 8'b11011011; // 8001 : 219 - 0xdb
      13'h1F42: dout  = 8'b01000010; // 8002 :  66 - 0x42
      13'h1F43: dout  = 8'b11011011; // 8003 : 219 - 0xdb
      13'h1F44: dout  = 8'b01000010; // 8004 :  66 - 0x42
      13'h1F45: dout  = 8'b00100110; // 8005 :  38 - 0x26
      13'h1F46: dout  = 8'b00100001; // 8006 :  33 - 0x21
      13'h1F47: dout  = 8'b01100110; // 8007 : 102 - 0x66
      13'h1F48: dout  = 8'b01000110; // 8008 :  70 - 0x46
      13'h1F49: dout  = 8'b11011011; // 8009 : 219 - 0xdb
      13'h1F4A: dout  = 8'b00100001; // 8010 :  33 - 0x21
      13'h1F4B: dout  = 8'b01101100; // 8011 : 108 - 0x6c
      13'h1F4C: dout  = 8'b00001110; // 8012 :  14 - 0xe
      13'h1F4D: dout  = 8'b11011111; // 8013 : 223 - 0xdf
      13'h1F4E: dout  = 8'b11011011; // 8014 : 219 - 0xdb
      13'h1F4F: dout  = 8'b11011011; // 8015 : 219 - 0xdb
      13'h1F50: dout  = 8'b11011011; // 8016 : 219 - 0xdb -- Background 0xf5
      13'h1F51: dout  = 8'b00100110; // 8017 :  38 - 0x26
      13'h1F52: dout  = 8'b11011011; // 8018 : 219 - 0xdb
      13'h1F53: dout  = 8'b11011111; // 8019 : 223 - 0xdf
      13'h1F54: dout  = 8'b11011011; // 8020 : 219 - 0xdb
      13'h1F55: dout  = 8'b11011111; // 8021 : 223 - 0xdf
      13'h1F56: dout  = 8'b11011011; // 8022 : 219 - 0xdb
      13'h1F57: dout  = 8'b11011011; // 8023 : 219 - 0xdb
      13'h1F58: dout  = 8'b11100100; // 8024 : 228 - 0xe4
      13'h1F59: dout  = 8'b11100101; // 8025 : 229 - 0xe5
      13'h1F5A: dout  = 8'b00100110; // 8026 :  38 - 0x26
      13'h1F5B: dout  = 8'b00100001; // 8027 :  33 - 0x21
      13'h1F5C: dout  = 8'b10000110; // 8028 : 134 - 0x86
      13'h1F5D: dout  = 8'b00010100; // 8029 :  20 - 0x14
      13'h1F5E: dout  = 8'b11011011; // 8030 : 219 - 0xdb
      13'h1F5F: dout  = 8'b11011011; // 8031 : 219 - 0xdb
      13'h1F60: dout  = 8'b11011011; // 8032 : 219 - 0xdb -- Background 0xf6
      13'h1F61: dout  = 8'b11011110; // 8033 : 222 - 0xde
      13'h1F62: dout  = 8'b01000011; // 8034 :  67 - 0x43
      13'h1F63: dout  = 8'b11011011; // 8035 : 219 - 0xdb
      13'h1F64: dout  = 8'b11100000; // 8036 : 224 - 0xe0
      13'h1F65: dout  = 8'b11011011; // 8037 : 219 - 0xdb
      13'h1F66: dout  = 8'b11011011; // 8038 : 219 - 0xdb
      13'h1F67: dout  = 8'b11011011; // 8039 : 219 - 0xdb
      13'h1F68: dout  = 8'b00100110; // 8040 :  38 - 0x26
      13'h1F69: dout  = 8'b11011011; // 8041 : 219 - 0xdb
      13'h1F6A: dout  = 8'b11100011; // 8042 : 227 - 0xe3
      13'h1F6B: dout  = 8'b11011011; // 8043 : 219 - 0xdb
      13'h1F6C: dout  = 8'b11100000; // 8044 : 224 - 0xe0
      13'h1F6D: dout  = 8'b11011011; // 8045 : 219 - 0xdb
      13'h1F6E: dout  = 8'b11011011; // 8046 : 219 - 0xdb
      13'h1F6F: dout  = 8'b11100110; // 8047 : 230 - 0xe6
      13'h1F70: dout  = 8'b11100011; // 8048 : 227 - 0xe3 -- Background 0xf7
      13'h1F71: dout  = 8'b00100110; // 8049 :  38 - 0x26
      13'h1F72: dout  = 8'b00100001; // 8050 :  33 - 0x21
      13'h1F73: dout  = 8'b10100110; // 8051 : 166 - 0xa6
      13'h1F74: dout  = 8'b00010100; // 8052 :  20 - 0x14
      13'h1F75: dout  = 8'b11011011; // 8053 : 219 - 0xdb
      13'h1F76: dout  = 8'b11011011; // 8054 : 219 - 0xdb
      13'h1F77: dout  = 8'b11011011; // 8055 : 219 - 0xdb
      13'h1F78: dout  = 8'b11011011; // 8056 : 219 - 0xdb
      13'h1F79: dout  = 8'b01000010; // 8057 :  66 - 0x42
      13'h1F7A: dout  = 8'b11011011; // 8058 : 219 - 0xdb
      13'h1F7B: dout  = 8'b11011011; // 8059 : 219 - 0xdb
      13'h1F7C: dout  = 8'b11011011; // 8060 : 219 - 0xdb
      13'h1F7D: dout  = 8'b11010100; // 8061 : 212 - 0xd4
      13'h1F7E: dout  = 8'b11011001; // 8062 : 217 - 0xd9
      13'h1F7F: dout  = 8'b00100110; // 8063 :  38 - 0x26
      13'h1F80: dout  = 8'b11011011; // 8064 : 219 - 0xdb -- Background 0xf8
      13'h1F81: dout  = 8'b11011001; // 8065 : 217 - 0xd9
      13'h1F82: dout  = 8'b11011011; // 8066 : 219 - 0xdb
      13'h1F83: dout  = 8'b11011011; // 8067 : 219 - 0xdb
      13'h1F84: dout  = 8'b11010100; // 8068 : 212 - 0xd4
      13'h1F85: dout  = 8'b11011001; // 8069 : 217 - 0xd9
      13'h1F86: dout  = 8'b11010100; // 8070 : 212 - 0xd4
      13'h1F87: dout  = 8'b11011001; // 8071 : 217 - 0xd9
      13'h1F88: dout  = 8'b11100111; // 8072 : 231 - 0xe7
      13'h1F89: dout  = 8'b00100001; // 8073 :  33 - 0x21
      13'h1F8A: dout  = 8'b11000101; // 8074 : 197 - 0xc5
      13'h1F8B: dout  = 8'b00010110; // 8075 :  22 - 0x16
      13'h1F8C: dout  = 8'b01011111; // 8076 :  95 - 0x5f
      13'h1F8D: dout  = 8'b10010101; // 8077 : 149 - 0x95
      13'h1F8E: dout  = 8'b10010101; // 8078 : 149 - 0x95
      13'h1F8F: dout  = 8'b10010101; // 8079 : 149 - 0x95
      13'h1F90: dout  = 8'b10010101; // 8080 : 149 - 0x95 -- Background 0xf9
      13'h1F91: dout  = 8'b10010101; // 8081 : 149 - 0x95
      13'h1F92: dout  = 8'b10010101; // 8082 : 149 - 0x95
      13'h1F93: dout  = 8'b10010101; // 8083 : 149 - 0x95
      13'h1F94: dout  = 8'b10010101; // 8084 : 149 - 0x95
      13'h1F95: dout  = 8'b10010111; // 8085 : 151 - 0x97
      13'h1F96: dout  = 8'b10011000; // 8086 : 152 - 0x98
      13'h1F97: dout  = 8'b01111000; // 8087 : 120 - 0x78
      13'h1F98: dout  = 8'b10010101; // 8088 : 149 - 0x95
      13'h1F99: dout  = 8'b10010110; // 8089 : 150 - 0x96
      13'h1F9A: dout  = 8'b10010101; // 8090 : 149 - 0x95
      13'h1F9B: dout  = 8'b10010101; // 8091 : 149 - 0x95
      13'h1F9C: dout  = 8'b10010111; // 8092 : 151 - 0x97
      13'h1F9D: dout  = 8'b10011000; // 8093 : 152 - 0x98
      13'h1F9E: dout  = 8'b10010111; // 8094 : 151 - 0x97
      13'h1F9F: dout  = 8'b10011000; // 8095 : 152 - 0x98
      13'h1FA0: dout  = 8'b10010101; // 8096 : 149 - 0x95 -- Background 0xfa
      13'h1FA1: dout  = 8'b01111010; // 8097 : 122 - 0x7a
      13'h1FA2: dout  = 8'b00100001; // 8098 :  33 - 0x21
      13'h1FA3: dout  = 8'b11101101; // 8099 : 237 - 0xed
      13'h1FA4: dout  = 8'b00001110; // 8100 :  14 - 0xe
      13'h1FA5: dout  = 8'b11001111; // 8101 : 207 - 0xcf
      13'h1FA6: dout  = 8'b00000001; // 8102 :   1 - 0x1
      13'h1FA7: dout  = 8'b00001001; // 8103 :   9 - 0x9
      13'h1FA8: dout  = 8'b00001000; // 8104 :   8 - 0x8
      13'h1FA9: dout  = 8'b00000101; // 8105 :   5 - 0x5
      13'h1FAA: dout  = 8'b00100100; // 8106 :  36 - 0x24
      13'h1FAB: dout  = 8'b00010111; // 8107 :  23 - 0x17
      13'h1FAC: dout  = 8'b00010010; // 8108 :  18 - 0x12
      13'h1FAD: dout  = 8'b00010111; // 8109 :  23 - 0x17
      13'h1FAE: dout  = 8'b00011101; // 8110 :  29 - 0x1d
      13'h1FAF: dout  = 8'b00001110; // 8111 :  14 - 0xe
      13'h1FB0: dout  = 8'b00010111; // 8112 :  23 - 0x17 -- Background 0xfb
      13'h1FB1: dout  = 8'b00001101; // 8113 :  13 - 0xd
      13'h1FB2: dout  = 8'b00011000; // 8114 :  24 - 0x18
      13'h1FB3: dout  = 8'b00100010; // 8115 :  34 - 0x22
      13'h1FB4: dout  = 8'b01001011; // 8116 :  75 - 0x4b
      13'h1FB5: dout  = 8'b00001101; // 8117 :  13 - 0xd
      13'h1FB6: dout  = 8'b00000001; // 8118 :   1 - 0x1
      13'h1FB7: dout  = 8'b00100100; // 8119 :  36 - 0x24
      13'h1FB8: dout  = 8'b00011001; // 8120 :  25 - 0x19
      13'h1FB9: dout  = 8'b00010101; // 8121 :  21 - 0x15
      13'h1FBA: dout  = 8'b00001010; // 8122 :  10 - 0xa
      13'h1FBB: dout  = 8'b00100010; // 8123 :  34 - 0x22
      13'h1FBC: dout  = 8'b00001110; // 8124 :  14 - 0xe
      13'h1FBD: dout  = 8'b00011011; // 8125 :  27 - 0x1b
      13'h1FBE: dout  = 8'b00100100; // 8126 :  36 - 0x24
      13'h1FBF: dout  = 8'b00010000; // 8127 :  16 - 0x10
      13'h1FC0: dout  = 8'b00001010; // 8128 :  10 - 0xa -- Background 0xfc
      13'h1FC1: dout  = 8'b00010110; // 8129 :  22 - 0x16
      13'h1FC2: dout  = 8'b00001110; // 8130 :  14 - 0xe
      13'h1FC3: dout  = 8'b00100010; // 8131 :  34 - 0x22
      13'h1FC4: dout  = 8'b10001011; // 8132 : 139 - 0x8b
      13'h1FC5: dout  = 8'b00001101; // 8133 :  13 - 0xd
      13'h1FC6: dout  = 8'b00000010; // 8134 :   2 - 0x2
      13'h1FC7: dout  = 8'b00100100; // 8135 :  36 - 0x24
      13'h1FC8: dout  = 8'b00011001; // 8136 :  25 - 0x19
      13'h1FC9: dout  = 8'b00010101; // 8137 :  21 - 0x15
      13'h1FCA: dout  = 8'b00001010; // 8138 :  10 - 0xa
      13'h1FCB: dout  = 8'b00100010; // 8139 :  34 - 0x22
      13'h1FCC: dout  = 8'b00001110; // 8140 :  14 - 0xe
      13'h1FCD: dout  = 8'b00011011; // 8141 :  27 - 0x1b
      13'h1FCE: dout  = 8'b00100100; // 8142 :  36 - 0x24
      13'h1FCF: dout  = 8'b00010000; // 8143 :  16 - 0x10
      13'h1FD0: dout  = 8'b00001010; // 8144 :  10 - 0xa -- Background 0xfd
      13'h1FD1: dout  = 8'b00010110; // 8145 :  22 - 0x16
      13'h1FD2: dout  = 8'b00001110; // 8146 :  14 - 0xe
      13'h1FD3: dout  = 8'b00100010; // 8147 :  34 - 0x22
      13'h1FD4: dout  = 8'b11101100; // 8148 : 236 - 0xec
      13'h1FD5: dout  = 8'b00000100; // 8149 :   4 - 0x4
      13'h1FD6: dout  = 8'b00011101; // 8150 :  29 - 0x1d
      13'h1FD7: dout  = 8'b00011000; // 8151 :  24 - 0x18
      13'h1FD8: dout  = 8'b00011001; // 8152 :  25 - 0x19
      13'h1FD9: dout  = 8'b00101000; // 8153 :  40 - 0x28
      13'h1FDA: dout  = 8'b00100010; // 8154 :  34 - 0x22
      13'h1FDB: dout  = 8'b11110110; // 8155 : 246 - 0xf6
      13'h1FDC: dout  = 8'b00000001; // 8156 :   1 - 0x1
      13'h1FDD: dout  = 8'b00000000; // 8157 :   0 - 0x0
      13'h1FDE: dout  = 8'b00100011; // 8158 :  35 - 0x23
      13'h1FDF: dout  = 8'b11001001; // 8159 : 201 - 0xc9
      13'h1FE0: dout  = 8'b01010110; // 8160 :  86 - 0x56 -- Background 0xfe
      13'h1FE1: dout  = 8'b01010101; // 8161 :  85 - 0x55
      13'h1FE2: dout  = 8'b00100011; // 8162 :  35 - 0x23
      13'h1FE3: dout  = 8'b11100010; // 8163 : 226 - 0xe2
      13'h1FE4: dout  = 8'b00000100; // 8164 :   4 - 0x4
      13'h1FE5: dout  = 8'b10011001; // 8165 : 153 - 0x99
      13'h1FE6: dout  = 8'b10101010; // 8166 : 170 - 0xaa
      13'h1FE7: dout  = 8'b10101010; // 8167 : 170 - 0xaa
      13'h1FE8: dout  = 8'b10101010; // 8168 : 170 - 0xaa
      13'h1FE9: dout  = 8'b00100011; // 8169 :  35 - 0x23
      13'h1FEA: dout  = 8'b11101010; // 8170 : 234 - 0xea
      13'h1FEB: dout  = 8'b00000100; // 8171 :   4 - 0x4
      13'h1FEC: dout  = 8'b10011001; // 8172 : 153 - 0x99
      13'h1FED: dout  = 8'b10101010; // 8173 : 170 - 0xaa
      13'h1FEE: dout  = 8'b10101010; // 8174 : 170 - 0xaa
      13'h1FEF: dout  = 8'b10101010; // 8175 : 170 - 0xaa
      13'h1FF0: dout  = 8'b00000000; // 8176 :   0 - 0x0 -- Background 0xff
      13'h1FF1: dout  = 8'b11111111; // 8177 : 255 - 0xff
      13'h1FF2: dout  = 8'b11111111; // 8178 : 255 - 0xff
      13'h1FF3: dout  = 8'b11111111; // 8179 : 255 - 0xff
      13'h1FF4: dout  = 8'b11111111; // 8180 : 255 - 0xff
      13'h1FF5: dout  = 8'b11111111; // 8181 : 255 - 0xff
      13'h1FF6: dout  = 8'b11111111; // 8182 : 255 - 0xff
      13'h1FF7: dout  = 8'b11111111; // 8183 : 255 - 0xff
      13'h1FF8: dout  = 8'b11111111; // 8184 : 255 - 0xff
      13'h1FF9: dout  = 8'b11111111; // 8185 : 255 - 0xff
      13'h1FFA: dout  = 8'b11111111; // 8186 : 255 - 0xff
      13'h1FFB: dout  = 8'b11111111; // 8187 : 255 - 0xff
      13'h1FFC: dout  = 8'b11111111; // 8188 : 255 - 0xff
      13'h1FFD: dout  = 8'b11111111; // 8189 : 255 - 0xff
      13'h1FFE: dout  = 8'b11111111; // 8190 : 255 - 0xff
      13'h1FFF: dout  = 8'b11111111; // 8191 : 255 - 0xff
    endcase
  end

endmodule
