--- Autcmatically generated VHDL ROM from a NES memory file----
---   NAME TABLE
-- https://wiki.nesdev.com/w/index.php/PPU_nametables
--- Only the first Name Table: 1KiB


---  Original memory dump file name: donkeykong_ntable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory with clock ------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_NTABLE_DONKEYKONG is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(10-1 downto 0);  --1024 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_NTABLE_DONKEYKONG;

architecture BEHAVIORAL of ROM_NTABLE_DONKEYKONG is
  signal addr_int  : natural range 0 to 2**10-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
     ------- Name Table 0---------
    "00100100", --    0 -  0x0  :   36 - 0x24 -- line 0x0
    "00100100", --    1 -  0x1  :   36 - 0x24
    "00100100", --    2 -  0x2  :   36 - 0x24
    "00100100", --    3 -  0x3  :   36 - 0x24
    "00100100", --    4 -  0x4  :   36 - 0x24
    "00100100", --    5 -  0x5  :   36 - 0x24
    "00100100", --    6 -  0x6  :   36 - 0x24
    "00100100", --    7 -  0x7  :   36 - 0x24
    "00100100", --    8 -  0x8  :   36 - 0x24
    "00100100", --    9 -  0x9  :   36 - 0x24
    "00100100", --   10 -  0xa  :   36 - 0x24
    "00100100", --   11 -  0xb  :   36 - 0x24
    "00100100", --   12 -  0xc  :   36 - 0x24
    "00100100", --   13 -  0xd  :   36 - 0x24
    "00100100", --   14 -  0xe  :   36 - 0x24
    "00100100", --   15 -  0xf  :   36 - 0x24
    "00100100", --   16 - 0x10  :   36 - 0x24
    "00100100", --   17 - 0x11  :   36 - 0x24
    "00100100", --   18 - 0x12  :   36 - 0x24
    "00100100", --   19 - 0x13  :   36 - 0x24
    "00100100", --   20 - 0x14  :   36 - 0x24
    "00100100", --   21 - 0x15  :   36 - 0x24
    "00100100", --   22 - 0x16  :   36 - 0x24
    "00100100", --   23 - 0x17  :   36 - 0x24
    "00100100", --   24 - 0x18  :   36 - 0x24
    "00100100", --   25 - 0x19  :   36 - 0x24
    "00100100", --   26 - 0x1a  :   36 - 0x24
    "00100100", --   27 - 0x1b  :   36 - 0x24
    "00100100", --   28 - 0x1c  :   36 - 0x24
    "00100100", --   29 - 0x1d  :   36 - 0x24
    "00100100", --   30 - 0x1e  :   36 - 0x24
    "00100100", --   31 - 0x1f  :   36 - 0x24
    "00100100", --   32 - 0x20  :   36 - 0x24 -- line 0x1
    "00100100", --   33 - 0x21  :   36 - 0x24
    "00100100", --   34 - 0x22  :   36 - 0x24
    "00100100", --   35 - 0x23  :   36 - 0x24
    "00100100", --   36 - 0x24  :   36 - 0x24
    "00100100", --   37 - 0x25  :   36 - 0x24
    "00100100", --   38 - 0x26  :   36 - 0x24
    "00100100", --   39 - 0x27  :   36 - 0x24
    "00100100", --   40 - 0x28  :   36 - 0x24
    "00100100", --   41 - 0x29  :   36 - 0x24
    "00111111", --   42 - 0x2a  :   63 - 0x3f
    "00100100", --   43 - 0x2b  :   36 - 0x24
    "00111111", --   44 - 0x2c  :   63 - 0x3f
    "00100100", --   45 - 0x2d  :   36 - 0x24
    "00100100", --   46 - 0x2e  :   36 - 0x24
    "00100100", --   47 - 0x2f  :   36 - 0x24
    "00100100", --   48 - 0x30  :   36 - 0x24
    "00100100", --   49 - 0x31  :   36 - 0x24
    "00100100", --   50 - 0x32  :   36 - 0x24
    "00100100", --   51 - 0x33  :   36 - 0x24
    "00100100", --   52 - 0x34  :   36 - 0x24
    "00100100", --   53 - 0x35  :   36 - 0x24
    "00100100", --   54 - 0x36  :   36 - 0x24
    "00100100", --   55 - 0x37  :   36 - 0x24
    "00100100", --   56 - 0x38  :   36 - 0x24
    "00100100", --   57 - 0x39  :   36 - 0x24
    "00100100", --   58 - 0x3a  :   36 - 0x24
    "00100100", --   59 - 0x3b  :   36 - 0x24
    "00100100", --   60 - 0x3c  :   36 - 0x24
    "00100100", --   61 - 0x3d  :   36 - 0x24
    "00100100", --   62 - 0x3e  :   36 - 0x24
    "00100100", --   63 - 0x3f  :   36 - 0x24
    "00100100", --   64 - 0x40  :   36 - 0x24 -- line 0x2
    "00100100", --   65 - 0x41  :   36 - 0x24
    "00100100", --   66 - 0x42  :   36 - 0x24
    "00100100", --   67 - 0x43  :   36 - 0x24
    "00100100", --   68 - 0x44  :   36 - 0x24
    "00100100", --   69 - 0x45  :   36 - 0x24
    "00100100", --   70 - 0x46  :   36 - 0x24
    "00100100", --   71 - 0x47  :   36 - 0x24
    "00100100", --   72 - 0x48  :   36 - 0x24
    "00100100", --   73 - 0x49  :   36 - 0x24
    "00111111", --   74 - 0x4a  :   63 - 0x3f
    "00100100", --   75 - 0x4b  :   36 - 0x24
    "00111111", --   76 - 0x4c  :   63 - 0x3f
    "00100100", --   77 - 0x4d  :   36 - 0x24
    "00100100", --   78 - 0x4e  :   36 - 0x24
    "00100100", --   79 - 0x4f  :   36 - 0x24
    "00100100", --   80 - 0x50  :   36 - 0x24
    "00100100", --   81 - 0x51  :   36 - 0x24
    "00100100", --   82 - 0x52  :   36 - 0x24
    "00100100", --   83 - 0x53  :   36 - 0x24
    "00100100", --   84 - 0x54  :   36 - 0x24
    "00100100", --   85 - 0x55  :   36 - 0x24
    "00100100", --   86 - 0x56  :   36 - 0x24
    "00100100", --   87 - 0x57  :   36 - 0x24
    "00100100", --   88 - 0x58  :   36 - 0x24
    "00100100", --   89 - 0x59  :   36 - 0x24
    "00100100", --   90 - 0x5a  :   36 - 0x24
    "00100100", --   91 - 0x5b  :   36 - 0x24
    "00100100", --   92 - 0x5c  :   36 - 0x24
    "00100100", --   93 - 0x5d  :   36 - 0x24
    "00100100", --   94 - 0x5e  :   36 - 0x24
    "00100100", --   95 - 0x5f  :   36 - 0x24
    "00100100", --   96 - 0x60  :   36 - 0x24 -- line 0x3
    "00100100", --   97 - 0x61  :   36 - 0x24
    "00100100", --   98 - 0x62  :   36 - 0x24
    "11111111", --   99 - 0x63  :  255 - 0xff
    "00000000", --  100 - 0x64  :    0 - 0x0
    "00000000", --  101 - 0x65  :    0 - 0x0
    "00000010", --  102 - 0x66  :    2 - 0x2
    "00000010", --  103 - 0x67  :    2 - 0x2
    "00000000", --  104 - 0x68  :    0 - 0x0
    "00000000", --  105 - 0x69  :    0 - 0x0
    "00111111", --  106 - 0x6a  :   63 - 0x3f
    "00100100", --  107 - 0x6b  :   36 - 0x24
    "00111111", --  108 - 0x6c  :   63 - 0x3f
    "11010000", --  109 - 0x6d  :  208 - 0xd0
    "11010001", --  110 - 0x6e  :  209 - 0xd1
    "11010010", --  111 - 0x6f  :  210 - 0xd2
    "00000000", --  112 - 0x70  :    0 - 0x0
    "00000000", --  113 - 0x71  :    0 - 0x0
    "00000010", --  114 - 0x72  :    2 - 0x2
    "00000010", --  115 - 0x73  :    2 - 0x2
    "00000000", --  116 - 0x74  :    0 - 0x0
    "00000000", --  117 - 0x75  :    0 - 0x0
    "00100100", --  118 - 0x76  :   36 - 0x24
    "00100100", --  119 - 0x77  :   36 - 0x24
    "00100100", --  120 - 0x78  :   36 - 0x24
    "00100100", --  121 - 0x79  :   36 - 0x24
    "00100100", --  122 - 0x7a  :   36 - 0x24
    "00100100", --  123 - 0x7b  :   36 - 0x24
    "00100100", --  124 - 0x7c  :   36 - 0x24
    "00100100", --  125 - 0x7d  :   36 - 0x24
    "00100100", --  126 - 0x7e  :   36 - 0x24
    "00100100", --  127 - 0x7f  :   36 - 0x24
    "00100100", --  128 - 0x80  :   36 - 0x24 -- line 0x4
    "01010000", --  129 - 0x81  :   80 - 0x50
    "01010100", --  130 - 0x82  :   84 - 0x54
    "01011000", --  131 - 0x83  :   88 - 0x58
    "00100100", --  132 - 0x84  :   36 - 0x24
    "00100100", --  133 - 0x85  :   36 - 0x24
    "10001100", --  134 - 0x86  :  140 - 0x8c
    "10010000", --  135 - 0x87  :  144 - 0x90
    "10010100", --  136 - 0x88  :  148 - 0x94
    "10011000", --  137 - 0x89  :  152 - 0x98
    "00111111", --  138 - 0x8a  :   63 - 0x3f
    "00100100", --  139 - 0x8b  :   36 - 0x24
    "00111111", --  140 - 0x8c  :   63 - 0x3f
    "00100100", --  141 - 0x8d  :   36 - 0x24
    "00100100", --  142 - 0x8e  :   36 - 0x24
    "00100100", --  143 - 0x8f  :   36 - 0x24
    "00100100", --  144 - 0x90  :   36 - 0x24
    "00100100", --  145 - 0x91  :   36 - 0x24
    "00100100", --  146 - 0x92  :   36 - 0x24
    "00100100", --  147 - 0x93  :   36 - 0x24
    "00100101", --  148 - 0x94  :   37 - 0x25
    "00010110", --  149 - 0x95  :   22 - 0x16
    "00101010", --  150 - 0x96  :   42 - 0x2a
    "00100110", --  151 - 0x97  :   38 - 0x26
    "00100111", --  152 - 0x98  :   39 - 0x27
    "00101000", --  153 - 0x99  :   40 - 0x28
    "00101001", --  154 - 0x9a  :   41 - 0x29
    "00101010", --  155 - 0x9b  :   42 - 0x2a
    "00010101", --  156 - 0x9c  :   21 - 0x15
    "00101101", --  157 - 0x9d  :   45 - 0x2d
    "00100100", --  158 - 0x9e  :   36 - 0x24
    "00100100", --  159 - 0x9f  :   36 - 0x24
    "00100100", --  160 - 0xa0  :   36 - 0x24 -- line 0x5
    "01010001", --  161 - 0xa1  :   81 - 0x51
    "01010101", --  162 - 0xa2  :   85 - 0x55
    "01011001", --  163 - 0xa3  :   89 - 0x59
    "00100100", --  164 - 0xa4  :   36 - 0x24
    "00100100", --  165 - 0xa5  :   36 - 0x24
    "10001101", --  166 - 0xa6  :  141 - 0x8d
    "10010001", --  167 - 0xa7  :  145 - 0x91
    "10010101", --  168 - 0xa8  :  149 - 0x95
    "10011001", --  169 - 0xa9  :  153 - 0x99
    "00111111", --  170 - 0xaa  :   63 - 0x3f
    "00100100", --  171 - 0xab  :   36 - 0x24
    "00111111", --  172 - 0xac  :   63 - 0x3f
    "00110000", --  173 - 0xad  :   48 - 0x30
    "00110000", --  174 - 0xae  :   48 - 0x30
    "00110000", --  175 - 0xaf  :   48 - 0x30
    "00110000", --  176 - 0xb0  :   48 - 0x30
    "00110000", --  177 - 0xb1  :   48 - 0x30
    "00110000", --  178 - 0xb2  :   48 - 0x30
    "00100100", --  179 - 0xb3  :   36 - 0x24
    "00101011", --  180 - 0xb4  :   43 - 0x2b
    "00000010", --  181 - 0xb5  :    2 - 0x2
    "00101100", --  182 - 0xb6  :   44 - 0x2c
    "00000011", --  183 - 0xb7  :    3 - 0x3
    "00000000", --  184 - 0xb8  :    0 - 0x0
    "00000000", --  185 - 0xb9  :    0 - 0x0
    "00000000", --  186 - 0xba  :    0 - 0x0
    "00101100", --  187 - 0xbb  :   44 - 0x2c
    "00000001", --  188 - 0xbc  :    1 - 0x1
    "00101111", --  189 - 0xbd  :   47 - 0x2f
    "00100100", --  190 - 0xbe  :   36 - 0x24
    "00100100", --  191 - 0xbf  :   36 - 0x24
    "00100100", --  192 - 0xc0  :   36 - 0x24 -- line 0x6
    "01010010", --  193 - 0xc1  :   82 - 0x52
    "01010110", --  194 - 0xc2  :   86 - 0x56
    "01011010", --  195 - 0xc3  :   90 - 0x5a
    "00100100", --  196 - 0xc4  :   36 - 0x24
    "10001010", --  197 - 0xc5  :  138 - 0x8a
    "10001110", --  198 - 0xc6  :  142 - 0x8e
    "10010010", --  199 - 0xc7  :  146 - 0x92
    "10010110", --  200 - 0xc8  :  150 - 0x96
    "10011010", --  201 - 0xc9  :  154 - 0x9a
    "00110000", --  202 - 0xca  :   48 - 0x30
    "00110000", --  203 - 0xcb  :   48 - 0x30
    "00110000", --  204 - 0xcc  :   48 - 0x30
    "00100100", --  205 - 0xcd  :   36 - 0x24
    "00100100", --  206 - 0xce  :   36 - 0x24
    "00100100", --  207 - 0xcf  :   36 - 0x24
    "00100100", --  208 - 0xd0  :   36 - 0x24
    "00100100", --  209 - 0xd1  :   36 - 0x24
    "00111111", --  210 - 0xd2  :   63 - 0x3f
    "00100100", --  211 - 0xd3  :   36 - 0x24
    "00100100", --  212 - 0xd4  :   36 - 0x24
    "00100100", --  213 - 0xd5  :   36 - 0x24
    "00100100", --  214 - 0xd6  :   36 - 0x24
    "00100100", --  215 - 0xd7  :   36 - 0x24
    "00100100", --  216 - 0xd8  :   36 - 0x24
    "00100100", --  217 - 0xd9  :   36 - 0x24
    "00100100", --  218 - 0xda  :   36 - 0x24
    "00100100", --  219 - 0xdb  :   36 - 0x24
    "00100100", --  220 - 0xdc  :   36 - 0x24
    "00100100", --  221 - 0xdd  :   36 - 0x24
    "00100100", --  222 - 0xde  :   36 - 0x24
    "00100100", --  223 - 0xdf  :   36 - 0x24
    "00100100", --  224 - 0xe0  :   36 - 0x24 -- line 0x7
    "01010011", --  225 - 0xe1  :   83 - 0x53
    "01010111", --  226 - 0xe2  :   87 - 0x57
    "01011011", --  227 - 0xe3  :   91 - 0x5b
    "10001001", --  228 - 0xe4  :  137 - 0x89
    "10001011", --  229 - 0xe5  :  139 - 0x8b
    "10001111", --  230 - 0xe6  :  143 - 0x8f
    "10010011", --  231 - 0xe7  :  147 - 0x93
    "10010111", --  232 - 0xe8  :  151 - 0x97
    "10011011", --  233 - 0xe9  :  155 - 0x9b
    "00111111", --  234 - 0xea  :   63 - 0x3f
    "00100100", --  235 - 0xeb  :   36 - 0x24
    "00111111", --  236 - 0xec  :   63 - 0x3f
    "00100100", --  237 - 0xed  :   36 - 0x24
    "00100100", --  238 - 0xee  :   36 - 0x24
    "00100100", --  239 - 0xef  :   36 - 0x24
    "00100100", --  240 - 0xf0  :   36 - 0x24
    "00100100", --  241 - 0xf1  :   36 - 0x24
    "00111111", --  242 - 0xf2  :   63 - 0x3f
    "00100100", --  243 - 0xf3  :   36 - 0x24
    "00100100", --  244 - 0xf4  :   36 - 0x24
    "00100100", --  245 - 0xf5  :   36 - 0x24
    "00100100", --  246 - 0xf6  :   36 - 0x24
    "00100100", --  247 - 0xf7  :   36 - 0x24
    "00100100", --  248 - 0xf8  :   36 - 0x24
    "00100100", --  249 - 0xf9  :   36 - 0x24
    "00100100", --  250 - 0xfa  :   36 - 0x24
    "00100100", --  251 - 0xfb  :   36 - 0x24
    "00100100", --  252 - 0xfc  :   36 - 0x24
    "00100100", --  253 - 0xfd  :   36 - 0x24
    "00100100", --  254 - 0xfe  :   36 - 0x24
    "00100100", --  255 - 0xff  :   36 - 0x24
    "00100100", --  256 - 0x100  :   36 - 0x24 -- line 0x8
    "00100100", --  257 - 0x101  :   36 - 0x24
    "00110000", --  258 - 0x102  :   48 - 0x30
    "00110000", --  259 - 0x103  :   48 - 0x30
    "00110000", --  260 - 0x104  :   48 - 0x30
    "00110000", --  261 - 0x105  :   48 - 0x30
    "00110000", --  262 - 0x106  :   48 - 0x30
    "00110000", --  263 - 0x107  :   48 - 0x30
    "00110000", --  264 - 0x108  :   48 - 0x30
    "00110000", --  265 - 0x109  :   48 - 0x30
    "00110000", --  266 - 0x10a  :   48 - 0x30
    "00110000", --  267 - 0x10b  :   48 - 0x30
    "00110000", --  268 - 0x10c  :   48 - 0x30
    "00110000", --  269 - 0x10d  :   48 - 0x30
    "00110000", --  270 - 0x10e  :   48 - 0x30
    "00110000", --  271 - 0x10f  :   48 - 0x30
    "00111110", --  272 - 0x110  :   62 - 0x3e
    "00111110", --  273 - 0x111  :   62 - 0x3e
    "01000101", --  274 - 0x112  :   69 - 0x45
    "00111101", --  275 - 0x113  :   61 - 0x3d
    "00111101", --  276 - 0x114  :   61 - 0x3d
    "00111101", --  277 - 0x115  :   61 - 0x3d
    "00111100", --  278 - 0x116  :   60 - 0x3c
    "00111100", --  279 - 0x117  :   60 - 0x3c
    "00111100", --  280 - 0x118  :   60 - 0x3c
    "00111011", --  281 - 0x119  :   59 - 0x3b
    "00111011", --  282 - 0x11a  :   59 - 0x3b
    "00111011", --  283 - 0x11b  :   59 - 0x3b
    "00100100", --  284 - 0x11c  :   36 - 0x24
    "00100100", --  285 - 0x11d  :   36 - 0x24
    "00100100", --  286 - 0x11e  :   36 - 0x24
    "00100100", --  287 - 0x11f  :   36 - 0x24
    "00100100", --  288 - 0x120  :   36 - 0x24 -- line 0x9
    "00100100", --  289 - 0x121  :   36 - 0x24
    "00100100", --  290 - 0x122  :   36 - 0x24
    "00100100", --  291 - 0x123  :   36 - 0x24
    "00100100", --  292 - 0x124  :   36 - 0x24
    "00100100", --  293 - 0x125  :   36 - 0x24
    "00100100", --  294 - 0x126  :   36 - 0x24
    "00100100", --  295 - 0x127  :   36 - 0x24
    "00100100", --  296 - 0x128  :   36 - 0x24
    "00100100", --  297 - 0x129  :   36 - 0x24
    "00100100", --  298 - 0x12a  :   36 - 0x24
    "00100100", --  299 - 0x12b  :   36 - 0x24
    "00100100", --  300 - 0x12c  :   36 - 0x24
    "00111111", --  301 - 0x12d  :   63 - 0x3f
    "00100100", --  302 - 0x12e  :   36 - 0x24
    "00100100", --  303 - 0x12f  :   36 - 0x24
    "00110111", --  304 - 0x130  :   55 - 0x37
    "00110111", --  305 - 0x131  :   55 - 0x37
    "00110111", --  306 - 0x132  :   55 - 0x37
    "00110110", --  307 - 0x133  :   54 - 0x36
    "00110110", --  308 - 0x134  :   54 - 0x36
    "00110110", --  309 - 0x135  :   54 - 0x36
    "00110101", --  310 - 0x136  :   53 - 0x35
    "00110101", --  311 - 0x137  :   53 - 0x35
    "00110101", --  312 - 0x138  :   53 - 0x35
    "01001001", --  313 - 0x139  :   73 - 0x49
    "00110100", --  314 - 0x13a  :   52 - 0x34
    "00110100", --  315 - 0x13b  :   52 - 0x34
    "00100100", --  316 - 0x13c  :   36 - 0x24
    "00100100", --  317 - 0x13d  :   36 - 0x24
    "00100100", --  318 - 0x13e  :   36 - 0x24
    "00100100", --  319 - 0x13f  :   36 - 0x24
    "00100100", --  320 - 0x140  :   36 - 0x24 -- line 0xa
    "00100100", --  321 - 0x141  :   36 - 0x24
    "00100100", --  322 - 0x142  :   36 - 0x24
    "00100100", --  323 - 0x143  :   36 - 0x24
    "00100100", --  324 - 0x144  :   36 - 0x24
    "00100100", --  325 - 0x145  :   36 - 0x24
    "00100100", --  326 - 0x146  :   36 - 0x24
    "00100100", --  327 - 0x147  :   36 - 0x24
    "00100100", --  328 - 0x148  :   36 - 0x24
    "00100100", --  329 - 0x149  :   36 - 0x24
    "00100100", --  330 - 0x14a  :   36 - 0x24
    "00100100", --  331 - 0x14b  :   36 - 0x24
    "00100100", --  332 - 0x14c  :   36 - 0x24
    "00100100", --  333 - 0x14d  :   36 - 0x24
    "00100100", --  334 - 0x14e  :   36 - 0x24
    "00100100", --  335 - 0x14f  :   36 - 0x24
    "00100100", --  336 - 0x150  :   36 - 0x24
    "00100100", --  337 - 0x151  :   36 - 0x24
    "00100100", --  338 - 0x152  :   36 - 0x24
    "00100100", --  339 - 0x153  :   36 - 0x24
    "00100100", --  340 - 0x154  :   36 - 0x24
    "00100100", --  341 - 0x155  :   36 - 0x24
    "00100100", --  342 - 0x156  :   36 - 0x24
    "00100100", --  343 - 0x157  :   36 - 0x24
    "00100100", --  344 - 0x158  :   36 - 0x24
    "00111111", --  345 - 0x159  :   63 - 0x3f
    "00100100", --  346 - 0x15a  :   36 - 0x24
    "00100100", --  347 - 0x15b  :   36 - 0x24
    "00100100", --  348 - 0x15c  :   36 - 0x24
    "00100100", --  349 - 0x15d  :   36 - 0x24
    "00100100", --  350 - 0x15e  :   36 - 0x24
    "00100100", --  351 - 0x15f  :   36 - 0x24
    "00100100", --  352 - 0x160  :   36 - 0x24 -- line 0xb
    "00100100", --  353 - 0x161  :   36 - 0x24
    "00100100", --  354 - 0x162  :   36 - 0x24
    "00100100", --  355 - 0x163  :   36 - 0x24
    "00100100", --  356 - 0x164  :   36 - 0x24
    "00100100", --  357 - 0x165  :   36 - 0x24
    "00100100", --  358 - 0x166  :   36 - 0x24
    "00100100", --  359 - 0x167  :   36 - 0x24
    "00100100", --  360 - 0x168  :   36 - 0x24
    "00100100", --  361 - 0x169  :   36 - 0x24
    "00100100", --  362 - 0x16a  :   36 - 0x24
    "00100100", --  363 - 0x16b  :   36 - 0x24
    "00100100", --  364 - 0x16c  :   36 - 0x24
    "01000000", --  365 - 0x16d  :   64 - 0x40
    "00111000", --  366 - 0x16e  :   56 - 0x38
    "00111000", --  367 - 0x16f  :   56 - 0x38
    "00111001", --  368 - 0x170  :   57 - 0x39
    "00111001", --  369 - 0x171  :   57 - 0x39
    "00111001", --  370 - 0x172  :   57 - 0x39
    "00111010", --  371 - 0x173  :   58 - 0x3a
    "00111010", --  372 - 0x174  :   58 - 0x3a
    "00111010", --  373 - 0x175  :   58 - 0x3a
    "00111011", --  374 - 0x176  :   59 - 0x3b
    "00111011", --  375 - 0x177  :   59 - 0x3b
    "00111011", --  376 - 0x178  :   59 - 0x3b
    "01000011", --  377 - 0x179  :   67 - 0x43
    "00111100", --  378 - 0x17a  :   60 - 0x3c
    "00111100", --  379 - 0x17b  :   60 - 0x3c
    "00111101", --  380 - 0x17c  :   61 - 0x3d
    "00111101", --  381 - 0x17d  :   61 - 0x3d
    "00100100", --  382 - 0x17e  :   36 - 0x24
    "00100100", --  383 - 0x17f  :   36 - 0x24
    "00100100", --  384 - 0x180  :   36 - 0x24 -- line 0xc
    "00100100", --  385 - 0x181  :   36 - 0x24
    "00100100", --  386 - 0x182  :   36 - 0x24
    "00100100", --  387 - 0x183  :   36 - 0x24
    "00111101", --  388 - 0x184  :   61 - 0x3d
    "00111101", --  389 - 0x185  :   61 - 0x3d
    "00111101", --  390 - 0x186  :   61 - 0x3d
    "00111110", --  391 - 0x187  :   62 - 0x3e
    "00111110", --  392 - 0x188  :   62 - 0x3e
    "00111110", --  393 - 0x189  :   62 - 0x3e
    "00110000", --  394 - 0x18a  :   48 - 0x30
    "00110000", --  395 - 0x18b  :   48 - 0x30
    "00110000", --  396 - 0x18c  :   48 - 0x30
    "00110001", --  397 - 0x18d  :   49 - 0x31
    "00110001", --  398 - 0x18e  :   49 - 0x31
    "00110001", --  399 - 0x18f  :   49 - 0x31
    "00110010", --  400 - 0x190  :   50 - 0x32
    "00110010", --  401 - 0x191  :   50 - 0x32
    "00110010", --  402 - 0x192  :   50 - 0x32
    "00110011", --  403 - 0x193  :   51 - 0x33
    "00110011", --  404 - 0x194  :   51 - 0x33
    "00110011", --  405 - 0x195  :   51 - 0x33
    "00110100", --  406 - 0x196  :   52 - 0x34
    "01001001", --  407 - 0x197  :   73 - 0x49
    "00110100", --  408 - 0x198  :   52 - 0x34
    "00110101", --  409 - 0x199  :   53 - 0x35
    "00110101", --  410 - 0x19a  :   53 - 0x35
    "00110101", --  411 - 0x19b  :   53 - 0x35
    "00110110", --  412 - 0x19c  :   54 - 0x36
    "00110110", --  413 - 0x19d  :   54 - 0x36
    "00100100", --  414 - 0x19e  :   36 - 0x24
    "00100100", --  415 - 0x19f  :   36 - 0x24
    "00100100", --  416 - 0x1a0  :   36 - 0x24 -- line 0xd
    "00100100", --  417 - 0x1a1  :   36 - 0x24
    "00100100", --  418 - 0x1a2  :   36 - 0x24
    "00100100", --  419 - 0x1a3  :   36 - 0x24
    "00110110", --  420 - 0x1a4  :   54 - 0x36
    "00110110", --  421 - 0x1a5  :   54 - 0x36
    "01001011", --  422 - 0x1a6  :   75 - 0x4b
    "00110111", --  423 - 0x1a7  :   55 - 0x37
    "00110111", --  424 - 0x1a8  :   55 - 0x37
    "00110111", --  425 - 0x1a9  :   55 - 0x37
    "00100100", --  426 - 0x1aa  :   36 - 0x24
    "00111111", --  427 - 0x1ab  :   63 - 0x3f
    "00100100", --  428 - 0x1ac  :   36 - 0x24
    "00100100", --  429 - 0x1ad  :   36 - 0x24
    "00100100", --  430 - 0x1ae  :   36 - 0x24
    "00100100", --  431 - 0x1af  :   36 - 0x24
    "00100100", --  432 - 0x1b0  :   36 - 0x24
    "00100100", --  433 - 0x1b1  :   36 - 0x24
    "00100100", --  434 - 0x1b2  :   36 - 0x24
    "00100100", --  435 - 0x1b3  :   36 - 0x24
    "00100100", --  436 - 0x1b4  :   36 - 0x24
    "00100100", --  437 - 0x1b5  :   36 - 0x24
    "00100100", --  438 - 0x1b6  :   36 - 0x24
    "00100100", --  439 - 0x1b7  :   36 - 0x24
    "00100100", --  440 - 0x1b8  :   36 - 0x24
    "00100100", --  441 - 0x1b9  :   36 - 0x24
    "00100100", --  442 - 0x1ba  :   36 - 0x24
    "00100100", --  443 - 0x1bb  :   36 - 0x24
    "00100100", --  444 - 0x1bc  :   36 - 0x24
    "00100100", --  445 - 0x1bd  :   36 - 0x24
    "00100100", --  446 - 0x1be  :   36 - 0x24
    "00100100", --  447 - 0x1bf  :   36 - 0x24
    "00100100", --  448 - 0x1c0  :   36 - 0x24 -- line 0xe
    "00100100", --  449 - 0x1c1  :   36 - 0x24
    "00100100", --  450 - 0x1c2  :   36 - 0x24
    "00100100", --  451 - 0x1c3  :   36 - 0x24
    "00100100", --  452 - 0x1c4  :   36 - 0x24
    "00100100", --  453 - 0x1c5  :   36 - 0x24
    "00111111", --  454 - 0x1c6  :   63 - 0x3f
    "00100100", --  455 - 0x1c7  :   36 - 0x24
    "00100100", --  456 - 0x1c8  :   36 - 0x24
    "00100100", --  457 - 0x1c9  :   36 - 0x24
    "00100100", --  458 - 0x1ca  :   36 - 0x24
    "00111111", --  459 - 0x1cb  :   63 - 0x3f
    "00100100", --  460 - 0x1cc  :   36 - 0x24
    "00100100", --  461 - 0x1cd  :   36 - 0x24
    "00100100", --  462 - 0x1ce  :   36 - 0x24
    "00100100", --  463 - 0x1cf  :   36 - 0x24
    "00100100", --  464 - 0x1d0  :   36 - 0x24
    "00100100", --  465 - 0x1d1  :   36 - 0x24
    "00100100", --  466 - 0x1d2  :   36 - 0x24
    "00100100", --  467 - 0x1d3  :   36 - 0x24
    "00100100", --  468 - 0x1d4  :   36 - 0x24
    "00100100", --  469 - 0x1d5  :   36 - 0x24
    "00100100", --  470 - 0x1d6  :   36 - 0x24
    "00100100", --  471 - 0x1d7  :   36 - 0x24
    "00100100", --  472 - 0x1d8  :   36 - 0x24
    "00100100", --  473 - 0x1d9  :   36 - 0x24
    "00100100", --  474 - 0x1da  :   36 - 0x24
    "00100100", --  475 - 0x1db  :   36 - 0x24
    "00100100", --  476 - 0x1dc  :   36 - 0x24
    "00100100", --  477 - 0x1dd  :   36 - 0x24
    "00100100", --  478 - 0x1de  :   36 - 0x24
    "00100100", --  479 - 0x1df  :   36 - 0x24
    "00100100", --  480 - 0x1e0  :   36 - 0x24 -- line 0xf
    "00100100", --  481 - 0x1e1  :   36 - 0x24
    "00110000", --  482 - 0x1e2  :   48 - 0x30
    "00110000", --  483 - 0x1e3  :   48 - 0x30
    "00111110", --  484 - 0x1e4  :   62 - 0x3e
    "00111110", --  485 - 0x1e5  :   62 - 0x3e
    "01000101", --  486 - 0x1e6  :   69 - 0x45
    "00111101", --  487 - 0x1e7  :   61 - 0x3d
    "00111101", --  488 - 0x1e8  :   61 - 0x3d
    "00111101", --  489 - 0x1e9  :   61 - 0x3d
    "00111100", --  490 - 0x1ea  :   60 - 0x3c
    "01000011", --  491 - 0x1eb  :   67 - 0x43
    "00111100", --  492 - 0x1ec  :   60 - 0x3c
    "00111011", --  493 - 0x1ed  :   59 - 0x3b
    "00111011", --  494 - 0x1ee  :   59 - 0x3b
    "00111011", --  495 - 0x1ef  :   59 - 0x3b
    "00111010", --  496 - 0x1f0  :   58 - 0x3a
    "00111010", --  497 - 0x1f1  :   58 - 0x3a
    "00111010", --  498 - 0x1f2  :   58 - 0x3a
    "00111001", --  499 - 0x1f3  :   57 - 0x39
    "00111001", --  500 - 0x1f4  :   57 - 0x39
    "00111001", --  501 - 0x1f5  :   57 - 0x39
    "00111000", --  502 - 0x1f6  :   56 - 0x38
    "01000000", --  503 - 0x1f7  :   64 - 0x40
    "00111000", --  504 - 0x1f8  :   56 - 0x38
    "00100100", --  505 - 0x1f9  :   36 - 0x24
    "00100100", --  506 - 0x1fa  :   36 - 0x24
    "00100100", --  507 - 0x1fb  :   36 - 0x24
    "00100100", --  508 - 0x1fc  :   36 - 0x24
    "00100100", --  509 - 0x1fd  :   36 - 0x24
    "00100100", --  510 - 0x1fe  :   36 - 0x24
    "00100100", --  511 - 0x1ff  :   36 - 0x24
    "00100100", --  512 - 0x200  :   36 - 0x24 -- line 0x10
    "00100100", --  513 - 0x201  :   36 - 0x24
    "00100100", --  514 - 0x202  :   36 - 0x24
    "00100100", --  515 - 0x203  :   36 - 0x24
    "00110111", --  516 - 0x204  :   55 - 0x37
    "00110111", --  517 - 0x205  :   55 - 0x37
    "00110111", --  518 - 0x206  :   55 - 0x37
    "00110110", --  519 - 0x207  :   54 - 0x36
    "00110110", --  520 - 0x208  :   54 - 0x36
    "00110110", --  521 - 0x209  :   54 - 0x36
    "01001010", --  522 - 0x20a  :   74 - 0x4a
    "00110101", --  523 - 0x20b  :   53 - 0x35
    "00110101", --  524 - 0x20c  :   53 - 0x35
    "00110100", --  525 - 0x20d  :   52 - 0x34
    "00110100", --  526 - 0x20e  :   52 - 0x34
    "00110100", --  527 - 0x20f  :   52 - 0x34
    "01001000", --  528 - 0x210  :   72 - 0x48
    "00110011", --  529 - 0x211  :   51 - 0x33
    "00110011", --  530 - 0x212  :   51 - 0x33
    "00110010", --  531 - 0x213  :   50 - 0x32
    "00110010", --  532 - 0x214  :   50 - 0x32
    "00110010", --  533 - 0x215  :   50 - 0x32
    "00110001", --  534 - 0x216  :   49 - 0x31
    "00110001", --  535 - 0x217  :   49 - 0x31
    "00110001", --  536 - 0x218  :   49 - 0x31
    "00110000", --  537 - 0x219  :   48 - 0x30
    "00110000", --  538 - 0x21a  :   48 - 0x30
    "00110000", --  539 - 0x21b  :   48 - 0x30
    "00100100", --  540 - 0x21c  :   36 - 0x24
    "00100100", --  541 - 0x21d  :   36 - 0x24
    "00100100", --  542 - 0x21e  :   36 - 0x24
    "00100100", --  543 - 0x21f  :   36 - 0x24
    "00100100", --  544 - 0x220  :   36 - 0x24 -- line 0x11
    "00100100", --  545 - 0x221  :   36 - 0x24
    "00100100", --  546 - 0x222  :   36 - 0x24
    "00100100", --  547 - 0x223  :   36 - 0x24
    "00100100", --  548 - 0x224  :   36 - 0x24
    "00100100", --  549 - 0x225  :   36 - 0x24
    "00100100", --  550 - 0x226  :   36 - 0x24
    "00100100", --  551 - 0x227  :   36 - 0x24
    "00100100", --  552 - 0x228  :   36 - 0x24
    "00100100", --  553 - 0x229  :   36 - 0x24
    "00100100", --  554 - 0x22a  :   36 - 0x24
    "00100100", --  555 - 0x22b  :   36 - 0x24
    "00100100", --  556 - 0x22c  :   36 - 0x24
    "00100100", --  557 - 0x22d  :   36 - 0x24
    "00100100", --  558 - 0x22e  :   36 - 0x24
    "00100100", --  559 - 0x22f  :   36 - 0x24
    "00111111", --  560 - 0x230  :   63 - 0x3f
    "00100100", --  561 - 0x231  :   36 - 0x24
    "00100100", --  562 - 0x232  :   36 - 0x24
    "00100100", --  563 - 0x233  :   36 - 0x24
    "00100100", --  564 - 0x234  :   36 - 0x24
    "00100100", --  565 - 0x235  :   36 - 0x24
    "00100100", --  566 - 0x236  :   36 - 0x24
    "00100100", --  567 - 0x237  :   36 - 0x24
    "00100100", --  568 - 0x238  :   36 - 0x24
    "00111111", --  569 - 0x239  :   63 - 0x3f
    "00100100", --  570 - 0x23a  :   36 - 0x24
    "00100100", --  571 - 0x23b  :   36 - 0x24
    "00100100", --  572 - 0x23c  :   36 - 0x24
    "00100100", --  573 - 0x23d  :   36 - 0x24
    "00100100", --  574 - 0x23e  :   36 - 0x24
    "00100100", --  575 - 0x23f  :   36 - 0x24
    "00100100", --  576 - 0x240  :   36 - 0x24 -- line 0x12
    "00100100", --  577 - 0x241  :   36 - 0x24
    "00100100", --  578 - 0x242  :   36 - 0x24
    "00100100", --  579 - 0x243  :   36 - 0x24
    "00100100", --  580 - 0x244  :   36 - 0x24
    "00100100", --  581 - 0x245  :   36 - 0x24
    "00100100", --  582 - 0x246  :   36 - 0x24
    "00100100", --  583 - 0x247  :   36 - 0x24
    "00100100", --  584 - 0x248  :   36 - 0x24
    "00100100", --  585 - 0x249  :   36 - 0x24
    "00111111", --  586 - 0x24a  :   63 - 0x3f
    "00100100", --  587 - 0x24b  :   36 - 0x24
    "00100100", --  588 - 0x24c  :   36 - 0x24
    "00100100", --  589 - 0x24d  :   36 - 0x24
    "00100100", --  590 - 0x24e  :   36 - 0x24
    "00100100", --  591 - 0x24f  :   36 - 0x24
    "00111111", --  592 - 0x250  :   63 - 0x3f
    "00100100", --  593 - 0x251  :   36 - 0x24
    "00100100", --  594 - 0x252  :   36 - 0x24
    "00100100", --  595 - 0x253  :   36 - 0x24
    "00100100", --  596 - 0x254  :   36 - 0x24
    "00100100", --  597 - 0x255  :   36 - 0x24
    "00100100", --  598 - 0x256  :   36 - 0x24
    "00100100", --  599 - 0x257  :   36 - 0x24
    "00100100", --  600 - 0x258  :   36 - 0x24
    "01000000", --  601 - 0x259  :   64 - 0x40
    "00111000", --  602 - 0x25a  :   56 - 0x38
    "00111000", --  603 - 0x25b  :   56 - 0x38
    "00111001", --  604 - 0x25c  :   57 - 0x39
    "00111001", --  605 - 0x25d  :   57 - 0x39
    "00100100", --  606 - 0x25e  :   36 - 0x24
    "00100100", --  607 - 0x25f  :   36 - 0x24
    "00100100", --  608 - 0x260  :   36 - 0x24 -- line 0x13
    "00100100", --  609 - 0x261  :   36 - 0x24
    "00100100", --  610 - 0x262  :   36 - 0x24
    "00100100", --  611 - 0x263  :   36 - 0x24
    "00111001", --  612 - 0x264  :   57 - 0x39
    "00111001", --  613 - 0x265  :   57 - 0x39
    "00111001", --  614 - 0x266  :   57 - 0x39
    "00111010", --  615 - 0x267  :   58 - 0x3a
    "00111010", --  616 - 0x268  :   58 - 0x3a
    "00111010", --  617 - 0x269  :   58 - 0x3a
    "01000010", --  618 - 0x26a  :   66 - 0x42
    "00111011", --  619 - 0x26b  :   59 - 0x3b
    "00111011", --  620 - 0x26c  :   59 - 0x3b
    "00111100", --  621 - 0x26d  :   60 - 0x3c
    "00111100", --  622 - 0x26e  :   60 - 0x3c
    "00111100", --  623 - 0x26f  :   60 - 0x3c
    "01000100", --  624 - 0x270  :   68 - 0x44
    "00111101", --  625 - 0x271  :   61 - 0x3d
    "00111101", --  626 - 0x272  :   61 - 0x3d
    "00111110", --  627 - 0x273  :   62 - 0x3e
    "00111110", --  628 - 0x274  :   62 - 0x3e
    "00111110", --  629 - 0x275  :   62 - 0x3e
    "00110000", --  630 - 0x276  :   48 - 0x30
    "00110000", --  631 - 0x277  :   48 - 0x30
    "00110000", --  632 - 0x278  :   48 - 0x30
    "00110001", --  633 - 0x279  :   49 - 0x31
    "00110001", --  634 - 0x27a  :   49 - 0x31
    "00110001", --  635 - 0x27b  :   49 - 0x31
    "00110010", --  636 - 0x27c  :   50 - 0x32
    "00110010", --  637 - 0x27d  :   50 - 0x32
    "00100100", --  638 - 0x27e  :   36 - 0x24
    "00100100", --  639 - 0x27f  :   36 - 0x24
    "00100100", --  640 - 0x280  :   36 - 0x24 -- line 0x14
    "00100100", --  641 - 0x281  :   36 - 0x24
    "00100100", --  642 - 0x282  :   36 - 0x24
    "00100100", --  643 - 0x283  :   36 - 0x24
    "00110010", --  644 - 0x284  :   50 - 0x32
    "00110010", --  645 - 0x285  :   50 - 0x32
    "01000111", --  646 - 0x286  :   71 - 0x47
    "00110011", --  647 - 0x287  :   51 - 0x33
    "00110011", --  648 - 0x288  :   51 - 0x33
    "00110011", --  649 - 0x289  :   51 - 0x33
    "00110100", --  650 - 0x28a  :   52 - 0x34
    "00110100", --  651 - 0x28b  :   52 - 0x34
    "00110100", --  652 - 0x28c  :   52 - 0x34
    "00110101", --  653 - 0x28d  :   53 - 0x35
    "01001010", --  654 - 0x28e  :   74 - 0x4a
    "00110101", --  655 - 0x28f  :   53 - 0x35
    "00110110", --  656 - 0x290  :   54 - 0x36
    "00110110", --  657 - 0x291  :   54 - 0x36
    "00110110", --  658 - 0x292  :   54 - 0x36
    "00110111", --  659 - 0x293  :   55 - 0x37
    "00110111", --  660 - 0x294  :   55 - 0x37
    "00110111", --  661 - 0x295  :   55 - 0x37
    "00100100", --  662 - 0x296  :   36 - 0x24
    "00100100", --  663 - 0x297  :   36 - 0x24
    "00100100", --  664 - 0x298  :   36 - 0x24
    "00100100", --  665 - 0x299  :   36 - 0x24
    "00100100", --  666 - 0x29a  :   36 - 0x24
    "00100100", --  667 - 0x29b  :   36 - 0x24
    "00100100", --  668 - 0x29c  :   36 - 0x24
    "00100100", --  669 - 0x29d  :   36 - 0x24
    "00100100", --  670 - 0x29e  :   36 - 0x24
    "00100100", --  671 - 0x29f  :   36 - 0x24
    "00100100", --  672 - 0x2a0  :   36 - 0x24 -- line 0x15
    "00100100", --  673 - 0x2a1  :   36 - 0x24
    "00100100", --  674 - 0x2a2  :   36 - 0x24
    "00100100", --  675 - 0x2a3  :   36 - 0x24
    "00100100", --  676 - 0x2a4  :   36 - 0x24
    "00100100", --  677 - 0x2a5  :   36 - 0x24
    "00111111", --  678 - 0x2a6  :   63 - 0x3f
    "00100100", --  679 - 0x2a7  :   36 - 0x24
    "00100100", --  680 - 0x2a8  :   36 - 0x24
    "00100100", --  681 - 0x2a9  :   36 - 0x24
    "00100100", --  682 - 0x2aa  :   36 - 0x24
    "00100100", --  683 - 0x2ab  :   36 - 0x24
    "00100100", --  684 - 0x2ac  :   36 - 0x24
    "00100100", --  685 - 0x2ad  :   36 - 0x24
    "00111111", --  686 - 0x2ae  :   63 - 0x3f
    "00100100", --  687 - 0x2af  :   36 - 0x24
    "00100100", --  688 - 0x2b0  :   36 - 0x24
    "00100100", --  689 - 0x2b1  :   36 - 0x24
    "00100100", --  690 - 0x2b2  :   36 - 0x24
    "00100100", --  691 - 0x2b3  :   36 - 0x24
    "00100100", --  692 - 0x2b4  :   36 - 0x24
    "00100100", --  693 - 0x2b5  :   36 - 0x24
    "00100100", --  694 - 0x2b6  :   36 - 0x24
    "00100100", --  695 - 0x2b7  :   36 - 0x24
    "00100100", --  696 - 0x2b8  :   36 - 0x24
    "00100100", --  697 - 0x2b9  :   36 - 0x24
    "00100100", --  698 - 0x2ba  :   36 - 0x24
    "00100100", --  699 - 0x2bb  :   36 - 0x24
    "00100100", --  700 - 0x2bc  :   36 - 0x24
    "00100100", --  701 - 0x2bd  :   36 - 0x24
    "00100100", --  702 - 0x2be  :   36 - 0x24
    "00100100", --  703 - 0x2bf  :   36 - 0x24
    "00100100", --  704 - 0x2c0  :   36 - 0x24 -- line 0x16
    "00100100", --  705 - 0x2c1  :   36 - 0x24
    "00111011", --  706 - 0x2c2  :   59 - 0x3b
    "00111011", --  707 - 0x2c3  :   59 - 0x3b
    "00111010", --  708 - 0x2c4  :   58 - 0x3a
    "00111010", --  709 - 0x2c5  :   58 - 0x3a
    "01000001", --  710 - 0x2c6  :   65 - 0x41
    "00111001", --  711 - 0x2c7  :   57 - 0x39
    "00111001", --  712 - 0x2c8  :   57 - 0x39
    "00111001", --  713 - 0x2c9  :   57 - 0x39
    "00111000", --  714 - 0x2ca  :   56 - 0x38
    "00111000", --  715 - 0x2cb  :   56 - 0x38
    "00111000", --  716 - 0x2cc  :   56 - 0x38
    "00100100", --  717 - 0x2cd  :   36 - 0x24
    "00111111", --  718 - 0x2ce  :   63 - 0x3f
    "00100100", --  719 - 0x2cf  :   36 - 0x24
    "00100100", --  720 - 0x2d0  :   36 - 0x24
    "00100100", --  721 - 0x2d1  :   36 - 0x24
    "00100100", --  722 - 0x2d2  :   36 - 0x24
    "00100100", --  723 - 0x2d3  :   36 - 0x24
    "00100100", --  724 - 0x2d4  :   36 - 0x24
    "00100100", --  725 - 0x2d5  :   36 - 0x24
    "00100100", --  726 - 0x2d6  :   36 - 0x24
    "00100100", --  727 - 0x2d7  :   36 - 0x24
    "00100100", --  728 - 0x2d8  :   36 - 0x24
    "00100100", --  729 - 0x2d9  :   36 - 0x24
    "00100100", --  730 - 0x2da  :   36 - 0x24
    "00100100", --  731 - 0x2db  :   36 - 0x24
    "00100100", --  732 - 0x2dc  :   36 - 0x24
    "00100100", --  733 - 0x2dd  :   36 - 0x24
    "00100100", --  734 - 0x2de  :   36 - 0x24
    "00100100", --  735 - 0x2df  :   36 - 0x24
    "00100100", --  736 - 0x2e0  :   36 - 0x24 -- line 0x17
    "00100100", --  737 - 0x2e1  :   36 - 0x24
    "00110100", --  738 - 0x2e2  :   52 - 0x34
    "00110100", --  739 - 0x2e3  :   52 - 0x34
    "00110011", --  740 - 0x2e4  :   51 - 0x33
    "00110011", --  741 - 0x2e5  :   51 - 0x33
    "00110011", --  742 - 0x2e6  :   51 - 0x33
    "00110010", --  743 - 0x2e7  :   50 - 0x32
    "00110010", --  744 - 0x2e8  :   50 - 0x32
    "00110010", --  745 - 0x2e9  :   50 - 0x32
    "00110001", --  746 - 0x2ea  :   49 - 0x31
    "00110001", --  747 - 0x2eb  :   49 - 0x31
    "01000110", --  748 - 0x2ec  :   70 - 0x46
    "00110000", --  749 - 0x2ed  :   48 - 0x30
    "00110000", --  750 - 0x2ee  :   48 - 0x30
    "00110000", --  751 - 0x2ef  :   48 - 0x30
    "00111110", --  752 - 0x2f0  :   62 - 0x3e
    "00111110", --  753 - 0x2f1  :   62 - 0x3e
    "00111110", --  754 - 0x2f2  :   62 - 0x3e
    "00111101", --  755 - 0x2f3  :   61 - 0x3d
    "00111101", --  756 - 0x2f4  :   61 - 0x3d
    "00111101", --  757 - 0x2f5  :   61 - 0x3d
    "00111100", --  758 - 0x2f6  :   60 - 0x3c
    "00111100", --  759 - 0x2f7  :   60 - 0x3c
    "00111100", --  760 - 0x2f8  :   60 - 0x3c
    "00111011", --  761 - 0x2f9  :   59 - 0x3b
    "00111011", --  762 - 0x2fa  :   59 - 0x3b
    "00111011", --  763 - 0x2fb  :   59 - 0x3b
    "00100100", --  764 - 0x2fc  :   36 - 0x24
    "00100100", --  765 - 0x2fd  :   36 - 0x24
    "00100100", --  766 - 0x2fe  :   36 - 0x24
    "00100100", --  767 - 0x2ff  :   36 - 0x24
    "00100100", --  768 - 0x300  :   36 - 0x24 -- line 0x18
    "00100100", --  769 - 0x301  :   36 - 0x24
    "00100100", --  770 - 0x302  :   36 - 0x24
    "00100100", --  771 - 0x303  :   36 - 0x24
    "00100100", --  772 - 0x304  :   36 - 0x24
    "00100100", --  773 - 0x305  :   36 - 0x24
    "00100100", --  774 - 0x306  :   36 - 0x24
    "00100100", --  775 - 0x307  :   36 - 0x24
    "00100100", --  776 - 0x308  :   36 - 0x24
    "00100100", --  777 - 0x309  :   36 - 0x24
    "00100100", --  778 - 0x30a  :   36 - 0x24
    "00100100", --  779 - 0x30b  :   36 - 0x24
    "00111111", --  780 - 0x30c  :   63 - 0x3f
    "00100100", --  781 - 0x30d  :   36 - 0x24
    "00100100", --  782 - 0x30e  :   36 - 0x24
    "00100100", --  783 - 0x30f  :   36 - 0x24
    "00110111", --  784 - 0x310  :   55 - 0x37
    "00110111", --  785 - 0x311  :   55 - 0x37
    "00110111", --  786 - 0x312  :   55 - 0x37
    "00110110", --  787 - 0x313  :   54 - 0x36
    "00110110", --  788 - 0x314  :   54 - 0x36
    "00110110", --  789 - 0x315  :   54 - 0x36
    "00110101", --  790 - 0x316  :   53 - 0x35
    "00110101", --  791 - 0x317  :   53 - 0x35
    "00110101", --  792 - 0x318  :   53 - 0x35
    "01001001", --  793 - 0x319  :   73 - 0x49
    "00110100", --  794 - 0x31a  :   52 - 0x34
    "00110100", --  795 - 0x31b  :   52 - 0x34
    "00100100", --  796 - 0x31c  :   36 - 0x24
    "00100100", --  797 - 0x31d  :   36 - 0x24
    "00100100", --  798 - 0x31e  :   36 - 0x24
    "00100100", --  799 - 0x31f  :   36 - 0x24
    "00100100", --  800 - 0x320  :   36 - 0x24 -- line 0x19
    "00100100", --  801 - 0x321  :   36 - 0x24
    "00100100", --  802 - 0x322  :   36 - 0x24
    "00100100", --  803 - 0x323  :   36 - 0x24
    "01001100", --  804 - 0x324  :   76 - 0x4c
    "01001110", --  805 - 0x325  :   78 - 0x4e
    "00100100", --  806 - 0x326  :   36 - 0x24
    "00100100", --  807 - 0x327  :   36 - 0x24
    "00100100", --  808 - 0x328  :   36 - 0x24
    "00100100", --  809 - 0x329  :   36 - 0x24
    "00100100", --  810 - 0x32a  :   36 - 0x24
    "00100100", --  811 - 0x32b  :   36 - 0x24
    "00100100", --  812 - 0x32c  :   36 - 0x24
    "00100100", --  813 - 0x32d  :   36 - 0x24
    "00100100", --  814 - 0x32e  :   36 - 0x24
    "00100100", --  815 - 0x32f  :   36 - 0x24
    "00100100", --  816 - 0x330  :   36 - 0x24
    "00100100", --  817 - 0x331  :   36 - 0x24
    "00100100", --  818 - 0x332  :   36 - 0x24
    "00100100", --  819 - 0x333  :   36 - 0x24
    "00100100", --  820 - 0x334  :   36 - 0x24
    "00100100", --  821 - 0x335  :   36 - 0x24
    "00100100", --  822 - 0x336  :   36 - 0x24
    "00100100", --  823 - 0x337  :   36 - 0x24
    "00100100", --  824 - 0x338  :   36 - 0x24
    "00111111", --  825 - 0x339  :   63 - 0x3f
    "00100100", --  826 - 0x33a  :   36 - 0x24
    "00100100", --  827 - 0x33b  :   36 - 0x24
    "00100100", --  828 - 0x33c  :   36 - 0x24
    "00100100", --  829 - 0x33d  :   36 - 0x24
    "00100100", --  830 - 0x33e  :   36 - 0x24
    "00100100", --  831 - 0x33f  :   36 - 0x24
    "00100100", --  832 - 0x340  :   36 - 0x24 -- line 0x1a
    "00100100", --  833 - 0x341  :   36 - 0x24
    "00100100", --  834 - 0x342  :   36 - 0x24
    "00100100", --  835 - 0x343  :   36 - 0x24
    "01001101", --  836 - 0x344  :   77 - 0x4d
    "01001111", --  837 - 0x345  :   79 - 0x4f
    "00100100", --  838 - 0x346  :   36 - 0x24
    "00100100", --  839 - 0x347  :   36 - 0x24
    "00100100", --  840 - 0x348  :   36 - 0x24
    "00100100", --  841 - 0x349  :   36 - 0x24
    "00100100", --  842 - 0x34a  :   36 - 0x24
    "00100100", --  843 - 0x34b  :   36 - 0x24
    "00111111", --  844 - 0x34c  :   63 - 0x3f
    "00100100", --  845 - 0x34d  :   36 - 0x24
    "00100100", --  846 - 0x34e  :   36 - 0x24
    "00100100", --  847 - 0x34f  :   36 - 0x24
    "00111000", --  848 - 0x350  :   56 - 0x38
    "00111000", --  849 - 0x351  :   56 - 0x38
    "00111000", --  850 - 0x352  :   56 - 0x38
    "00111001", --  851 - 0x353  :   57 - 0x39
    "00111001", --  852 - 0x354  :   57 - 0x39
    "00111001", --  853 - 0x355  :   57 - 0x39
    "00111010", --  854 - 0x356  :   58 - 0x3a
    "00111010", --  855 - 0x357  :   58 - 0x3a
    "00111010", --  856 - 0x358  :   58 - 0x3a
    "01000010", --  857 - 0x359  :   66 - 0x42
    "00111011", --  858 - 0x35a  :   59 - 0x3b
    "00111011", --  859 - 0x35b  :   59 - 0x3b
    "00111100", --  860 - 0x35c  :   60 - 0x3c
    "00111100", --  861 - 0x35d  :   60 - 0x3c
    "00111100", --  862 - 0x35e  :   60 - 0x3c
    "00100100", --  863 - 0x35f  :   36 - 0x24
    "00100100", --  864 - 0x360  :   36 - 0x24 -- line 0x1b
    "00110000", --  865 - 0x361  :   48 - 0x30
    "00110000", --  866 - 0x362  :   48 - 0x30
    "00110000", --  867 - 0x363  :   48 - 0x30
    "00110000", --  868 - 0x364  :   48 - 0x30
    "00110000", --  869 - 0x365  :   48 - 0x30
    "00110000", --  870 - 0x366  :   48 - 0x30
    "00110000", --  871 - 0x367  :   48 - 0x30
    "00110000", --  872 - 0x368  :   48 - 0x30
    "00110000", --  873 - 0x369  :   48 - 0x30
    "00110000", --  874 - 0x36a  :   48 - 0x30
    "00110000", --  875 - 0x36b  :   48 - 0x30
    "00110000", --  876 - 0x36c  :   48 - 0x30
    "00110000", --  877 - 0x36d  :   48 - 0x30
    "00110000", --  878 - 0x36e  :   48 - 0x30
    "00110000", --  879 - 0x36f  :   48 - 0x30
    "00110001", --  880 - 0x370  :   49 - 0x31
    "00110001", --  881 - 0x371  :   49 - 0x31
    "00110001", --  882 - 0x372  :   49 - 0x31
    "00110010", --  883 - 0x373  :   50 - 0x32
    "00110010", --  884 - 0x374  :   50 - 0x32
    "00110010", --  885 - 0x375  :   50 - 0x32
    "00110011", --  886 - 0x376  :   51 - 0x33
    "00110011", --  887 - 0x377  :   51 - 0x33
    "00110011", --  888 - 0x378  :   51 - 0x33
    "00110100", --  889 - 0x379  :   52 - 0x34
    "00110100", --  890 - 0x37a  :   52 - 0x34
    "00110100", --  891 - 0x37b  :   52 - 0x34
    "00110101", --  892 - 0x37c  :   53 - 0x35
    "00110101", --  893 - 0x37d  :   53 - 0x35
    "00110101", --  894 - 0x37e  :   53 - 0x35
    "00100100", --  895 - 0x37f  :   36 - 0x24
    "00100100", --  896 - 0x380  :   36 - 0x24 -- line 0x1c
    "00100100", --  897 - 0x381  :   36 - 0x24
    "00100100", --  898 - 0x382  :   36 - 0x24
    "00100100", --  899 - 0x383  :   36 - 0x24
    "00100100", --  900 - 0x384  :   36 - 0x24
    "00100100", --  901 - 0x385  :   36 - 0x24
    "00100100", --  902 - 0x386  :   36 - 0x24
    "00100100", --  903 - 0x387  :   36 - 0x24
    "00100100", --  904 - 0x388  :   36 - 0x24
    "00100100", --  905 - 0x389  :   36 - 0x24
    "00100100", --  906 - 0x38a  :   36 - 0x24
    "00100100", --  907 - 0x38b  :   36 - 0x24
    "00100100", --  908 - 0x38c  :   36 - 0x24
    "00100100", --  909 - 0x38d  :   36 - 0x24
    "00100100", --  910 - 0x38e  :   36 - 0x24
    "00100100", --  911 - 0x38f  :   36 - 0x24
    "00100100", --  912 - 0x390  :   36 - 0x24
    "00100100", --  913 - 0x391  :   36 - 0x24
    "00100100", --  914 - 0x392  :   36 - 0x24
    "00100100", --  915 - 0x393  :   36 - 0x24
    "00100100", --  916 - 0x394  :   36 - 0x24
    "00100100", --  917 - 0x395  :   36 - 0x24
    "00100100", --  918 - 0x396  :   36 - 0x24
    "00100100", --  919 - 0x397  :   36 - 0x24
    "00100100", --  920 - 0x398  :   36 - 0x24
    "00100100", --  921 - 0x399  :   36 - 0x24
    "00100100", --  922 - 0x39a  :   36 - 0x24
    "00100100", --  923 - 0x39b  :   36 - 0x24
    "00100100", --  924 - 0x39c  :   36 - 0x24
    "00100100", --  925 - 0x39d  :   36 - 0x24
    "00100100", --  926 - 0x39e  :   36 - 0x24
    "00100100", --  927 - 0x39f  :   36 - 0x24
    "00100100", --  928 - 0x3a0  :   36 - 0x24 -- line 0x1d
    "00100100", --  929 - 0x3a1  :   36 - 0x24
    "00100100", --  930 - 0x3a2  :   36 - 0x24
    "00100100", --  931 - 0x3a3  :   36 - 0x24
    "00100100", --  932 - 0x3a4  :   36 - 0x24
    "00100100", --  933 - 0x3a5  :   36 - 0x24
    "00100100", --  934 - 0x3a6  :   36 - 0x24
    "00100100", --  935 - 0x3a7  :   36 - 0x24
    "00100100", --  936 - 0x3a8  :   36 - 0x24
    "00100100", --  937 - 0x3a9  :   36 - 0x24
    "00100100", --  938 - 0x3aa  :   36 - 0x24
    "00100100", --  939 - 0x3ab  :   36 - 0x24
    "00100100", --  940 - 0x3ac  :   36 - 0x24
    "00100100", --  941 - 0x3ad  :   36 - 0x24
    "00100100", --  942 - 0x3ae  :   36 - 0x24
    "00100100", --  943 - 0x3af  :   36 - 0x24
    "00100100", --  944 - 0x3b0  :   36 - 0x24
    "00100100", --  945 - 0x3b1  :   36 - 0x24
    "00100100", --  946 - 0x3b2  :   36 - 0x24
    "00100100", --  947 - 0x3b3  :   36 - 0x24
    "00100100", --  948 - 0x3b4  :   36 - 0x24
    "00100100", --  949 - 0x3b5  :   36 - 0x24
    "00100100", --  950 - 0x3b6  :   36 - 0x24
    "00100100", --  951 - 0x3b7  :   36 - 0x24
    "00100100", --  952 - 0x3b8  :   36 - 0x24
    "00100100", --  953 - 0x3b9  :   36 - 0x24
    "00100100", --  954 - 0x3ba  :   36 - 0x24
    "00100100", --  955 - 0x3bb  :   36 - 0x24
    "00100100", --  956 - 0x3bc  :   36 - 0x24
    "00100100", --  957 - 0x3bd  :   36 - 0x24
    "00100100", --  958 - 0x3be  :   36 - 0x24
    "00100100", --  959 - 0x3bf  :   36 - 0x24
        ---- Attribute Table 0----
    "11111111", --  960 - 0x3c0  :  255 - 0xff
    "11111111", --  961 - 0x3c1  :  255 - 0xff
    "11111111", --  962 - 0x3c2  :  255 - 0xff
    "11111111", --  963 - 0x3c3  :  255 - 0xff
    "11111111", --  964 - 0x3c4  :  255 - 0xff
    "11111111", --  965 - 0x3c5  :  255 - 0xff
    "11111111", --  966 - 0x3c6  :  255 - 0xff
    "11111111", --  967 - 0x3c7  :  255 - 0xff
    "01010101", --  968 - 0x3c8  :   85 - 0x55
    "10101010", --  969 - 0x3c9  :  170 - 0xaa
    "00100010", --  970 - 0x3ca  :   34 - 0x22
    "00000000", --  971 - 0x3cb  :    0 - 0x0
    "00000000", --  972 - 0x3cc  :    0 - 0x0
    "00001111", --  973 - 0x3cd  :   15 - 0xf
    "00001111", --  974 - 0x3ce  :   15 - 0xf
    "00001111", --  975 - 0x3cf  :   15 - 0xf
    "00000000", --  976 - 0x3d0  :    0 - 0x0
    "00000000", --  977 - 0x3d1  :    0 - 0x0
    "00000000", --  978 - 0x3d2  :    0 - 0x0
    "00000000", --  979 - 0x3d3  :    0 - 0x0
    "00000000", --  980 - 0x3d4  :    0 - 0x0
    "00000000", --  981 - 0x3d5  :    0 - 0x0
    "00000000", --  982 - 0x3d6  :    0 - 0x0
    "00000000", --  983 - 0x3d7  :    0 - 0x0
    "00000000", --  984 - 0x3d8  :    0 - 0x0
    "00000000", --  985 - 0x3d9  :    0 - 0x0
    "00000000", --  986 - 0x3da  :    0 - 0x0
    "00000000", --  987 - 0x3db  :    0 - 0x0
    "00000000", --  988 - 0x3dc  :    0 - 0x0
    "00000000", --  989 - 0x3dd  :    0 - 0x0
    "00000000", --  990 - 0x3de  :    0 - 0x0
    "00000000", --  991 - 0x3df  :    0 - 0x0
    "00000000", --  992 - 0x3e0  :    0 - 0x0
    "00000000", --  993 - 0x3e1  :    0 - 0x0
    "00000000", --  994 - 0x3e2  :    0 - 0x0
    "00000000", --  995 - 0x3e3  :    0 - 0x0
    "00000000", --  996 - 0x3e4  :    0 - 0x0
    "00000000", --  997 - 0x3e5  :    0 - 0x0
    "00000000", --  998 - 0x3e6  :    0 - 0x0
    "00000000", --  999 - 0x3e7  :    0 - 0x0
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0
    "00000000", -- 1001 - 0x3e9  :    0 - 0x0
    "00000000", -- 1002 - 0x3ea  :    0 - 0x0
    "00000000", -- 1003 - 0x3eb  :    0 - 0x0
    "00000000", -- 1004 - 0x3ec  :    0 - 0x0
    "00000000", -- 1005 - 0x3ed  :    0 - 0x0
    "00000000", -- 1006 - 0x3ee  :    0 - 0x0
    "00000000", -- 1007 - 0x3ef  :    0 - 0x0
    "00000000", -- 1008 - 0x3f0  :    0 - 0x0
    "00000000", -- 1009 - 0x3f1  :    0 - 0x0
    "00000000", -- 1010 - 0x3f2  :    0 - 0x0
    "00000000", -- 1011 - 0x3f3  :    0 - 0x0
    "00000000", -- 1012 - 0x3f4  :    0 - 0x0
    "00000000", -- 1013 - 0x3f5  :    0 - 0x0
    "00000000", -- 1014 - 0x3f6  :    0 - 0x0
    "00000000", -- 1015 - 0x3f7  :    0 - 0x0
    "00000000", -- 1016 - 0x3f8  :    0 - 0x0
    "00000000", -- 1017 - 0x3f9  :    0 - 0x0
    "00000000", -- 1018 - 0x3fa  :    0 - 0x0
    "00000000", -- 1019 - 0x3fb  :    0 - 0x0
    "00000000", -- 1020 - 0x3fc  :    0 - 0x0
    "00000000", -- 1021 - 0x3fd  :    0 - 0x0
    "00000000", -- 1022 - 0x3fe  :    0 - 0x0
    "00000000"  -- 1023 - 0x3ff  :    0 - 0x0
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
