//- Autcmatically generated verilog ROM from a NES memory file----
//-   SPRITEs MEMORY (OAM)
// https://wiki.nesdev.com/w/index.php/PPU_OAM


//-  Original memory dump file name: pacman_oam_00.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_OAM_PACMAN_00
  (
     input     clk,   // clock
     input      [8-1:0] addr,  //256 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
      8'h0: dout <= 8'b10101011; //    0 : 171 - 0xab -- Sprite 0x0
      8'h1: dout <= 8'b00000010; //    1 :   2 - 0x2
      8'h2: dout <= 8'b00000000; //    2 :   0 - 0x0
      8'h3: dout <= 8'b01001111; //    3 :  79 - 0x4f
      8'h4: dout <= 8'b10101011; //    4 : 171 - 0xab -- Sprite 0x1
      8'h5: dout <= 8'b00000001; //    5 :   1 - 0x1
      8'h6: dout <= 8'b00000000; //    6 :   0 - 0x0
      8'h7: dout <= 8'b01010111; //    7 :  87 - 0x57
      8'h8: dout <= 8'b10110011; //    8 : 179 - 0xb3 -- Sprite 0x2
      8'h9: dout <= 8'b00000010; //    9 :   2 - 0x2
      8'hA: dout <= 8'b10000000; //   10 : 128 - 0x80
      8'hB: dout <= 8'b01001111; //   11 :  79 - 0x4f
      8'hC: dout <= 8'b10110011; //   12 : 179 - 0xb3 -- Sprite 0x3
      8'hD: dout <= 8'b00000001; //   13 :   1 - 0x1
      8'hE: dout <= 8'b10000000; //   14 : 128 - 0x80
      8'hF: dout <= 8'b01010111; //   15 :  87 - 0x57
      8'h10: dout <= 8'b01011011; //   16 :  91 - 0x5b -- Sprite 0x4
      8'h11: dout <= 8'b00011011; //   17 :  27 - 0x1b
      8'h12: dout <= 8'b00000000; //   18 :   0 - 0x0
      8'h13: dout <= 8'b01010000; //   19 :  80 - 0x50
      8'h14: dout <= 8'b01011011; //   20 :  91 - 0x5b -- Sprite 0x5
      8'h15: dout <= 8'b00011100; //   21 :  28 - 0x1c
      8'h16: dout <= 8'b00000000; //   22 :   0 - 0x0
      8'h17: dout <= 8'b01011000; //   23 :  88 - 0x58
      8'h18: dout <= 8'b01100011; //   24 :  99 - 0x63 -- Sprite 0x6
      8'h19: dout <= 8'b00011101; //   25 :  29 - 0x1d
      8'h1A: dout <= 8'b00000000; //   26 :   0 - 0x0
      8'h1B: dout <= 8'b01010000; //   27 :  80 - 0x50
      8'h1C: dout <= 8'b01100011; //   28 :  99 - 0x63 -- Sprite 0x7
      8'h1D: dout <= 8'b00011111; //   29 :  31 - 0x1f
      8'h1E: dout <= 8'b00000000; //   30 :   0 - 0x0
      8'h1F: dout <= 8'b01011000; //   31 :  88 - 0x58
      8'h20: dout <= 8'b01101111; //   32 : 111 - 0x6f -- Sprite 0x8
      8'h21: dout <= 8'b00011000; //   33 :  24 - 0x18
      8'h22: dout <= 8'b00000001; //   34 :   1 - 0x1
      8'h23: dout <= 8'b01010100; //   35 :  84 - 0x54
      8'h24: dout <= 8'b01101111; //   36 : 111 - 0x6f -- Sprite 0x9
      8'h25: dout <= 8'b00011000; //   37 :  24 - 0x18
      8'h26: dout <= 8'b01000001; //   38 :  65 - 0x41
      8'h27: dout <= 8'b01011100; //   39 :  92 - 0x5c
      8'h28: dout <= 8'b01110111; //   40 : 119 - 0x77 -- Sprite 0xa
      8'h29: dout <= 8'b00011001; //   41 :  25 - 0x19
      8'h2A: dout <= 8'b00000001; //   42 :   1 - 0x1
      8'h2B: dout <= 8'b01010100; //   43 :  84 - 0x54
      8'h2C: dout <= 8'b01110111; //   44 : 119 - 0x77 -- Sprite 0xb
      8'h2D: dout <= 8'b00011001; //   45 :  25 - 0x19
      8'h2E: dout <= 8'b01000001; //   46 :  65 - 0x41
      8'h2F: dout <= 8'b01011100; //   47 :  92 - 0x5c
      8'h30: dout <= 8'b01101111; //   48 : 111 - 0x6f -- Sprite 0xc
      8'h31: dout <= 8'b00011000; //   49 :  24 - 0x18
      8'h32: dout <= 8'b00000010; //   50 :   2 - 0x2
      8'h33: dout <= 8'b01001100; //   51 :  76 - 0x4c
      8'h34: dout <= 8'b01101111; //   52 : 111 - 0x6f -- Sprite 0xd
      8'h35: dout <= 8'b00011000; //   53 :  24 - 0x18
      8'h36: dout <= 8'b01000010; //   54 :  66 - 0x42
      8'h37: dout <= 8'b01010100; //   55 :  84 - 0x54
      8'h38: dout <= 8'b01110111; //   56 : 119 - 0x77 -- Sprite 0xe
      8'h39: dout <= 8'b00011001; //   57 :  25 - 0x19
      8'h3A: dout <= 8'b00000010; //   58 :   2 - 0x2
      8'h3B: dout <= 8'b01001100; //   59 :  76 - 0x4c
      8'h3C: dout <= 8'b01110111; //   60 : 119 - 0x77 -- Sprite 0xf
      8'h3D: dout <= 8'b00011001; //   61 :  25 - 0x19
      8'h3E: dout <= 8'b01000010; //   62 :  66 - 0x42
      8'h3F: dout <= 8'b01010100; //   63 :  84 - 0x54
      8'h40: dout <= 8'b01101111; //   64 : 111 - 0x6f -- Sprite 0x10
      8'h41: dout <= 8'b00011000; //   65 :  24 - 0x18
      8'h42: dout <= 8'b00000011; //   66 :   3 - 0x3
      8'h43: dout <= 8'b01011100; //   67 :  92 - 0x5c
      8'h44: dout <= 8'b01101111; //   68 : 111 - 0x6f -- Sprite 0x11
      8'h45: dout <= 8'b00011000; //   69 :  24 - 0x18
      8'h46: dout <= 8'b01000011; //   70 :  67 - 0x43
      8'h47: dout <= 8'b01100100; //   71 : 100 - 0x64
      8'h48: dout <= 8'b01110111; //   72 : 119 - 0x77 -- Sprite 0x12
      8'h49: dout <= 8'b00011001; //   73 :  25 - 0x19
      8'h4A: dout <= 8'b00000011; //   74 :   3 - 0x3
      8'h4B: dout <= 8'b01011100; //   75 :  92 - 0x5c
      8'h4C: dout <= 8'b01110111; //   76 : 119 - 0x77 -- Sprite 0x13
      8'h4D: dout <= 8'b00011001; //   77 :  25 - 0x19
      8'h4E: dout <= 8'b01000011; //   78 :  67 - 0x43
      8'h4F: dout <= 8'b01100100; //   79 : 100 - 0x64
      8'h50: dout <= 8'b11111111; //   80 : 255 - 0xff -- Sprite 0x14
      8'h51: dout <= 8'b01001100; //   81 :  76 - 0x4c
      8'h52: dout <= 8'b00000000; //   82 :   0 - 0x0
      8'h53: dout <= 8'b11111111; //   83 : 255 - 0xff
      8'h54: dout <= 8'b11111111; //   84 : 255 - 0xff -- Sprite 0x15
      8'h55: dout <= 8'b01001100; //   85 :  76 - 0x4c
      8'h56: dout <= 8'b00000000; //   86 :   0 - 0x0
      8'h57: dout <= 8'b11111111; //   87 : 255 - 0xff
      8'h58: dout <= 8'b11111111; //   88 : 255 - 0xff -- Sprite 0x16
      8'h59: dout <= 8'b01001100; //   89 :  76 - 0x4c
      8'h5A: dout <= 8'b00000000; //   90 :   0 - 0x0
      8'h5B: dout <= 8'b11111111; //   91 : 255 - 0xff
      8'h5C: dout <= 8'b11111111; //   92 : 255 - 0xff -- Sprite 0x17
      8'h5D: dout <= 8'b01001100; //   93 :  76 - 0x4c
      8'h5E: dout <= 8'b00000000; //   94 :   0 - 0x0
      8'h5F: dout <= 8'b11111111; //   95 : 255 - 0xff
      8'h60: dout <= 8'b00000000; //   96 :   0 - 0x0 -- Sprite 0x18
      8'h61: dout <= 8'b00000000; //   97 :   0 - 0x0
      8'h62: dout <= 8'b00000000; //   98 :   0 - 0x0
      8'h63: dout <= 8'b00000000; //   99 :   0 - 0x0
      8'h64: dout <= 8'b00000000; //  100 :   0 - 0x0 -- Sprite 0x19
      8'h65: dout <= 8'b00000000; //  101 :   0 - 0x0
      8'h66: dout <= 8'b00000000; //  102 :   0 - 0x0
      8'h67: dout <= 8'b00000000; //  103 :   0 - 0x0
      8'h68: dout <= 8'b00000000; //  104 :   0 - 0x0 -- Sprite 0x1a
      8'h69: dout <= 8'b00000000; //  105 :   0 - 0x0
      8'h6A: dout <= 8'b00000000; //  106 :   0 - 0x0
      8'h6B: dout <= 8'b00000000; //  107 :   0 - 0x0
      8'h6C: dout <= 8'b00000000; //  108 :   0 - 0x0 -- Sprite 0x1b
      8'h6D: dout <= 8'b00000000; //  109 :   0 - 0x0
      8'h6E: dout <= 8'b00000000; //  110 :   0 - 0x0
      8'h6F: dout <= 8'b00000000; //  111 :   0 - 0x0
      8'h70: dout <= 8'b00000000; //  112 :   0 - 0x0 -- Sprite 0x1c
      8'h71: dout <= 8'b00000000; //  113 :   0 - 0x0
      8'h72: dout <= 8'b00000000; //  114 :   0 - 0x0
      8'h73: dout <= 8'b00000000; //  115 :   0 - 0x0
      8'h74: dout <= 8'b00000000; //  116 :   0 - 0x0 -- Sprite 0x1d
      8'h75: dout <= 8'b00000000; //  117 :   0 - 0x0
      8'h76: dout <= 8'b00000000; //  118 :   0 - 0x0
      8'h77: dout <= 8'b00000000; //  119 :   0 - 0x0
      8'h78: dout <= 8'b00000000; //  120 :   0 - 0x0 -- Sprite 0x1e
      8'h79: dout <= 8'b00000000; //  121 :   0 - 0x0
      8'h7A: dout <= 8'b00000000; //  122 :   0 - 0x0
      8'h7B: dout <= 8'b00000000; //  123 :   0 - 0x0
      8'h7C: dout <= 8'b00000000; //  124 :   0 - 0x0 -- Sprite 0x1f
      8'h7D: dout <= 8'b00000000; //  125 :   0 - 0x0
      8'h7E: dout <= 8'b00000000; //  126 :   0 - 0x0
      8'h7F: dout <= 8'b00000000; //  127 :   0 - 0x0
      8'h80: dout <= 8'b00000000; //  128 :   0 - 0x0 -- Sprite 0x20
      8'h81: dout <= 8'b00000000; //  129 :   0 - 0x0
      8'h82: dout <= 8'b00000000; //  130 :   0 - 0x0
      8'h83: dout <= 8'b00000000; //  131 :   0 - 0x0
      8'h84: dout <= 8'b00000000; //  132 :   0 - 0x0 -- Sprite 0x21
      8'h85: dout <= 8'b00000000; //  133 :   0 - 0x0
      8'h86: dout <= 8'b00000000; //  134 :   0 - 0x0
      8'h87: dout <= 8'b00000000; //  135 :   0 - 0x0
      8'h88: dout <= 8'b00000000; //  136 :   0 - 0x0 -- Sprite 0x22
      8'h89: dout <= 8'b00000000; //  137 :   0 - 0x0
      8'h8A: dout <= 8'b00000000; //  138 :   0 - 0x0
      8'h8B: dout <= 8'b00000000; //  139 :   0 - 0x0
      8'h8C: dout <= 8'b00000000; //  140 :   0 - 0x0 -- Sprite 0x23
      8'h8D: dout <= 8'b00000000; //  141 :   0 - 0x0
      8'h8E: dout <= 8'b00000000; //  142 :   0 - 0x0
      8'h8F: dout <= 8'b00000000; //  143 :   0 - 0x0
      8'h90: dout <= 8'b00000000; //  144 :   0 - 0x0 -- Sprite 0x24
      8'h91: dout <= 8'b00000000; //  145 :   0 - 0x0
      8'h92: dout <= 8'b00000000; //  146 :   0 - 0x0
      8'h93: dout <= 8'b00000000; //  147 :   0 - 0x0
      8'h94: dout <= 8'b00000000; //  148 :   0 - 0x0 -- Sprite 0x25
      8'h95: dout <= 8'b00000000; //  149 :   0 - 0x0
      8'h96: dout <= 8'b00000000; //  150 :   0 - 0x0
      8'h97: dout <= 8'b00000000; //  151 :   0 - 0x0
      8'h98: dout <= 8'b00000000; //  152 :   0 - 0x0 -- Sprite 0x26
      8'h99: dout <= 8'b00000000; //  153 :   0 - 0x0
      8'h9A: dout <= 8'b00000000; //  154 :   0 - 0x0
      8'h9B: dout <= 8'b00000000; //  155 :   0 - 0x0
      8'h9C: dout <= 8'b00000000; //  156 :   0 - 0x0 -- Sprite 0x27
      8'h9D: dout <= 8'b00000000; //  157 :   0 - 0x0
      8'h9E: dout <= 8'b00000000; //  158 :   0 - 0x0
      8'h9F: dout <= 8'b00000000; //  159 :   0 - 0x0
      8'hA0: dout <= 8'b00000000; //  160 :   0 - 0x0 -- Sprite 0x28
      8'hA1: dout <= 8'b00000000; //  161 :   0 - 0x0
      8'hA2: dout <= 8'b00000000; //  162 :   0 - 0x0
      8'hA3: dout <= 8'b00000000; //  163 :   0 - 0x0
      8'hA4: dout <= 8'b00000000; //  164 :   0 - 0x0 -- Sprite 0x29
      8'hA5: dout <= 8'b00000000; //  165 :   0 - 0x0
      8'hA6: dout <= 8'b00000000; //  166 :   0 - 0x0
      8'hA7: dout <= 8'b00000000; //  167 :   0 - 0x0
      8'hA8: dout <= 8'b00000000; //  168 :   0 - 0x0 -- Sprite 0x2a
      8'hA9: dout <= 8'b00000000; //  169 :   0 - 0x0
      8'hAA: dout <= 8'b00000000; //  170 :   0 - 0x0
      8'hAB: dout <= 8'b00000000; //  171 :   0 - 0x0
      8'hAC: dout <= 8'b00000000; //  172 :   0 - 0x0 -- Sprite 0x2b
      8'hAD: dout <= 8'b00000000; //  173 :   0 - 0x0
      8'hAE: dout <= 8'b00000000; //  174 :   0 - 0x0
      8'hAF: dout <= 8'b00000000; //  175 :   0 - 0x0
      8'hB0: dout <= 8'b00000000; //  176 :   0 - 0x0 -- Sprite 0x2c
      8'hB1: dout <= 8'b00000000; //  177 :   0 - 0x0
      8'hB2: dout <= 8'b00000000; //  178 :   0 - 0x0
      8'hB3: dout <= 8'b00000000; //  179 :   0 - 0x0
      8'hB4: dout <= 8'b00000000; //  180 :   0 - 0x0 -- Sprite 0x2d
      8'hB5: dout <= 8'b00000000; //  181 :   0 - 0x0
      8'hB6: dout <= 8'b00000000; //  182 :   0 - 0x0
      8'hB7: dout <= 8'b00000000; //  183 :   0 - 0x0
      8'hB8: dout <= 8'b00000000; //  184 :   0 - 0x0 -- Sprite 0x2e
      8'hB9: dout <= 8'b00000000; //  185 :   0 - 0x0
      8'hBA: dout <= 8'b00000000; //  186 :   0 - 0x0
      8'hBB: dout <= 8'b00000000; //  187 :   0 - 0x0
      8'hBC: dout <= 8'b00000000; //  188 :   0 - 0x0 -- Sprite 0x2f
      8'hBD: dout <= 8'b00000000; //  189 :   0 - 0x0
      8'hBE: dout <= 8'b00000000; //  190 :   0 - 0x0
      8'hBF: dout <= 8'b00000000; //  191 :   0 - 0x0
      8'hC0: dout <= 8'b00000000; //  192 :   0 - 0x0 -- Sprite 0x30
      8'hC1: dout <= 8'b00000000; //  193 :   0 - 0x0
      8'hC2: dout <= 8'b00000000; //  194 :   0 - 0x0
      8'hC3: dout <= 8'b00000000; //  195 :   0 - 0x0
      8'hC4: dout <= 8'b00000000; //  196 :   0 - 0x0 -- Sprite 0x31
      8'hC5: dout <= 8'b00000000; //  197 :   0 - 0x0
      8'hC6: dout <= 8'b00000000; //  198 :   0 - 0x0
      8'hC7: dout <= 8'b00000000; //  199 :   0 - 0x0
      8'hC8: dout <= 8'b00000000; //  200 :   0 - 0x0 -- Sprite 0x32
      8'hC9: dout <= 8'b00000000; //  201 :   0 - 0x0
      8'hCA: dout <= 8'b00000000; //  202 :   0 - 0x0
      8'hCB: dout <= 8'b00000000; //  203 :   0 - 0x0
      8'hCC: dout <= 8'b00000000; //  204 :   0 - 0x0 -- Sprite 0x33
      8'hCD: dout <= 8'b00000000; //  205 :   0 - 0x0
      8'hCE: dout <= 8'b00000000; //  206 :   0 - 0x0
      8'hCF: dout <= 8'b00000000; //  207 :   0 - 0x0
      8'hD0: dout <= 8'b00000000; //  208 :   0 - 0x0 -- Sprite 0x34
      8'hD1: dout <= 8'b00000000; //  209 :   0 - 0x0
      8'hD2: dout <= 8'b00000000; //  210 :   0 - 0x0
      8'hD3: dout <= 8'b00000000; //  211 :   0 - 0x0
      8'hD4: dout <= 8'b00000000; //  212 :   0 - 0x0 -- Sprite 0x35
      8'hD5: dout <= 8'b00000000; //  213 :   0 - 0x0
      8'hD6: dout <= 8'b00000000; //  214 :   0 - 0x0
      8'hD7: dout <= 8'b00000000; //  215 :   0 - 0x0
      8'hD8: dout <= 8'b00000000; //  216 :   0 - 0x0 -- Sprite 0x36
      8'hD9: dout <= 8'b00000000; //  217 :   0 - 0x0
      8'hDA: dout <= 8'b00000000; //  218 :   0 - 0x0
      8'hDB: dout <= 8'b00000000; //  219 :   0 - 0x0
      8'hDC: dout <= 8'b00000000; //  220 :   0 - 0x0 -- Sprite 0x37
      8'hDD: dout <= 8'b00000000; //  221 :   0 - 0x0
      8'hDE: dout <= 8'b00000000; //  222 :   0 - 0x0
      8'hDF: dout <= 8'b00000000; //  223 :   0 - 0x0
      8'hE0: dout <= 8'b00000000; //  224 :   0 - 0x0 -- Sprite 0x38
      8'hE1: dout <= 8'b00000000; //  225 :   0 - 0x0
      8'hE2: dout <= 8'b00000000; //  226 :   0 - 0x0
      8'hE3: dout <= 8'b00000000; //  227 :   0 - 0x0
      8'hE4: dout <= 8'b00000000; //  228 :   0 - 0x0 -- Sprite 0x39
      8'hE5: dout <= 8'b00000000; //  229 :   0 - 0x0
      8'hE6: dout <= 8'b00000000; //  230 :   0 - 0x0
      8'hE7: dout <= 8'b00000000; //  231 :   0 - 0x0
      8'hE8: dout <= 8'b00000000; //  232 :   0 - 0x0 -- Sprite 0x3a
      8'hE9: dout <= 8'b00000000; //  233 :   0 - 0x0
      8'hEA: dout <= 8'b00000000; //  234 :   0 - 0x0
      8'hEB: dout <= 8'b00000000; //  235 :   0 - 0x0
      8'hEC: dout <= 8'b00000000; //  236 :   0 - 0x0 -- Sprite 0x3b
      8'hED: dout <= 8'b00000000; //  237 :   0 - 0x0
      8'hEE: dout <= 8'b00000000; //  238 :   0 - 0x0
      8'hEF: dout <= 8'b00000000; //  239 :   0 - 0x0
      8'hF0: dout <= 8'b00000000; //  240 :   0 - 0x0 -- Sprite 0x3c
      8'hF1: dout <= 8'b00000000; //  241 :   0 - 0x0
      8'hF2: dout <= 8'b00000000; //  242 :   0 - 0x0
      8'hF3: dout <= 8'b00000000; //  243 :   0 - 0x0
      8'hF4: dout <= 8'b00000000; //  244 :   0 - 0x0 -- Sprite 0x3d
      8'hF5: dout <= 8'b00000000; //  245 :   0 - 0x0
      8'hF6: dout <= 8'b00000000; //  246 :   0 - 0x0
      8'hF7: dout <= 8'b00000000; //  247 :   0 - 0x0
      8'hF8: dout <= 8'b00000000; //  248 :   0 - 0x0 -- Sprite 0x3e
      8'hF9: dout <= 8'b00000000; //  249 :   0 - 0x0
      8'hFA: dout <= 8'b00000000; //  250 :   0 - 0x0
      8'hFB: dout <= 8'b00000000; //  251 :   0 - 0x0
      8'hFC: dout <= 8'b00000000; //  252 :   0 - 0x0 -- Sprite 0x3f
      8'hFD: dout <= 8'b00000000; //  253 :   0 - 0x0
      8'hFE: dout <= 8'b00000000; //  254 :   0 - 0x0
      8'hFF: dout <= 8'b00000000; //  255 :   0 - 0x0
    endcase
  end

endmodule
