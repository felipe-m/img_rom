--- Autcmatically generated VHDL ROM from a NES memory file----
---   SPRITEs MEMORY (OAM)
-- https://wiki.nesdev.com/w/index.php/PPU_OAM


---  Original memory dump file name: sprilo_oam_00.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_OAM_SPRILO_00 is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(8-1 downto 0);  --256 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_OAM_SPRILO_00;

architecture BEHAVIORAL of ROM_OAM_SPRILO_00 is
  signal addr_int  : natural range 0 to 2**8-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
    "00110000", --    0 -  0x0  :   48 - 0x30 -- Sprite 0x0
    "00001001", --    1 -  0x1  :    9 - 0x9
    "00000001", --    2 -  0x2  :    1 - 0x1
    "10010001", --    3 -  0x3  :  145 - 0x91
    "11111110", --    4 -  0x4  :  254 - 0xfe -- Sprite 0x1
    "11111110", --    5 -  0x5  :  254 - 0xfe
    "11100010", --    6 -  0x6  :  226 - 0xe2
    "11111110", --    7 -  0x7  :  254 - 0xfe
    "11111110", --    8 -  0x8  :  254 - 0xfe -- Sprite 0x2
    "11111110", --    9 -  0x9  :  254 - 0xfe
    "11100010", --   10 -  0xa  :  226 - 0xe2
    "11111110", --   11 -  0xb  :  254 - 0xfe
    "11111110", --   12 -  0xc  :  254 - 0xfe -- Sprite 0x3
    "11111110", --   13 -  0xd  :  254 - 0xfe
    "11100010", --   14 -  0xe  :  226 - 0xe2
    "11111110", --   15 -  0xf  :  254 - 0xfe
    "11111110", --   16 - 0x10  :  254 - 0xfe -- Sprite 0x4
    "11111110", --   17 - 0x11  :  254 - 0xfe
    "11100010", --   18 - 0x12  :  226 - 0xe2
    "11111110", --   19 - 0x13  :  254 - 0xfe
    "11111110", --   20 - 0x14  :  254 - 0xfe -- Sprite 0x5
    "11111110", --   21 - 0x15  :  254 - 0xfe
    "11100010", --   22 - 0x16  :  226 - 0xe2
    "11111110", --   23 - 0x17  :  254 - 0xfe
    "11111110", --   24 - 0x18  :  254 - 0xfe -- Sprite 0x6
    "11111110", --   25 - 0x19  :  254 - 0xfe
    "11100010", --   26 - 0x1a  :  226 - 0xe2
    "11111110", --   27 - 0x1b  :  254 - 0xfe
    "11111110", --   28 - 0x1c  :  254 - 0xfe -- Sprite 0x7
    "11111110", --   29 - 0x1d  :  254 - 0xfe
    "11100010", --   30 - 0x1e  :  226 - 0xe2
    "11111110", --   31 - 0x1f  :  254 - 0xfe
    "11111110", --   32 - 0x20  :  254 - 0xfe -- Sprite 0x8
    "11111110", --   33 - 0x21  :  254 - 0xfe
    "11100010", --   34 - 0x22  :  226 - 0xe2
    "11111110", --   35 - 0x23  :  254 - 0xfe
    "11111110", --   36 - 0x24  :  254 - 0xfe -- Sprite 0x9
    "11111110", --   37 - 0x25  :  254 - 0xfe
    "11100010", --   38 - 0x26  :  226 - 0xe2
    "11111110", --   39 - 0x27  :  254 - 0xfe
    "11111110", --   40 - 0x28  :  254 - 0xfe -- Sprite 0xa
    "11111110", --   41 - 0x29  :  254 - 0xfe
    "11100010", --   42 - 0x2a  :  226 - 0xe2
    "11111110", --   43 - 0x2b  :  254 - 0xfe
    "11111110", --   44 - 0x2c  :  254 - 0xfe -- Sprite 0xb
    "11111110", --   45 - 0x2d  :  254 - 0xfe
    "11100010", --   46 - 0x2e  :  226 - 0xe2
    "11111110", --   47 - 0x2f  :  254 - 0xfe
    "11111110", --   48 - 0x30  :  254 - 0xfe -- Sprite 0xc
    "11111110", --   49 - 0x31  :  254 - 0xfe
    "11100010", --   50 - 0x32  :  226 - 0xe2
    "11111110", --   51 - 0x33  :  254 - 0xfe
    "11111110", --   52 - 0x34  :  254 - 0xfe -- Sprite 0xd
    "11111110", --   53 - 0x35  :  254 - 0xfe
    "11100010", --   54 - 0x36  :  226 - 0xe2
    "11111110", --   55 - 0x37  :  254 - 0xfe
    "11111110", --   56 - 0x38  :  254 - 0xfe -- Sprite 0xe
    "11111110", --   57 - 0x39  :  254 - 0xfe
    "11100010", --   58 - 0x3a  :  226 - 0xe2
    "11111110", --   59 - 0x3b  :  254 - 0xfe
    "11111110", --   60 - 0x3c  :  254 - 0xfe -- Sprite 0xf
    "11111110", --   61 - 0x3d  :  254 - 0xfe
    "11100010", --   62 - 0x3e  :  226 - 0xe2
    "11111110", --   63 - 0x3f  :  254 - 0xfe
    "11111110", --   64 - 0x40  :  254 - 0xfe -- Sprite 0x10
    "11111110", --   65 - 0x41  :  254 - 0xfe
    "11100010", --   66 - 0x42  :  226 - 0xe2
    "11111110", --   67 - 0x43  :  254 - 0xfe
    "11111110", --   68 - 0x44  :  254 - 0xfe -- Sprite 0x11
    "11111110", --   69 - 0x45  :  254 - 0xfe
    "11100010", --   70 - 0x46  :  226 - 0xe2
    "11111110", --   71 - 0x47  :  254 - 0xfe
    "11111110", --   72 - 0x48  :  254 - 0xfe -- Sprite 0x12
    "11111110", --   73 - 0x49  :  254 - 0xfe
    "11100010", --   74 - 0x4a  :  226 - 0xe2
    "11111110", --   75 - 0x4b  :  254 - 0xfe
    "11111110", --   76 - 0x4c  :  254 - 0xfe -- Sprite 0x13
    "11111110", --   77 - 0x4d  :  254 - 0xfe
    "11100010", --   78 - 0x4e  :  226 - 0xe2
    "11111110", --   79 - 0x4f  :  254 - 0xfe
    "11111110", --   80 - 0x50  :  254 - 0xfe -- Sprite 0x14
    "11111110", --   81 - 0x51  :  254 - 0xfe
    "11100010", --   82 - 0x52  :  226 - 0xe2
    "11111110", --   83 - 0x53  :  254 - 0xfe
    "11111110", --   84 - 0x54  :  254 - 0xfe -- Sprite 0x15
    "11111110", --   85 - 0x55  :  254 - 0xfe
    "11100010", --   86 - 0x56  :  226 - 0xe2
    "11111110", --   87 - 0x57  :  254 - 0xfe
    "11111110", --   88 - 0x58  :  254 - 0xfe -- Sprite 0x16
    "11111110", --   89 - 0x59  :  254 - 0xfe
    "11100010", --   90 - 0x5a  :  226 - 0xe2
    "11111110", --   91 - 0x5b  :  254 - 0xfe
    "11111110", --   92 - 0x5c  :  254 - 0xfe -- Sprite 0x17
    "11111110", --   93 - 0x5d  :  254 - 0xfe
    "11100010", --   94 - 0x5e  :  226 - 0xe2
    "11111110", --   95 - 0x5f  :  254 - 0xfe
    "11111110", --   96 - 0x60  :  254 - 0xfe -- Sprite 0x18
    "11111110", --   97 - 0x61  :  254 - 0xfe
    "11100010", --   98 - 0x62  :  226 - 0xe2
    "11111110", --   99 - 0x63  :  254 - 0xfe
    "11111110", --  100 - 0x64  :  254 - 0xfe -- Sprite 0x19
    "11111110", --  101 - 0x65  :  254 - 0xfe
    "11100010", --  102 - 0x66  :  226 - 0xe2
    "11111110", --  103 - 0x67  :  254 - 0xfe
    "11111110", --  104 - 0x68  :  254 - 0xfe -- Sprite 0x1a
    "11111110", --  105 - 0x69  :  254 - 0xfe
    "11100010", --  106 - 0x6a  :  226 - 0xe2
    "11111110", --  107 - 0x6b  :  254 - 0xfe
    "11111110", --  108 - 0x6c  :  254 - 0xfe -- Sprite 0x1b
    "11111110", --  109 - 0x6d  :  254 - 0xfe
    "11100010", --  110 - 0x6e  :  226 - 0xe2
    "11111110", --  111 - 0x6f  :  254 - 0xfe
    "11111110", --  112 - 0x70  :  254 - 0xfe -- Sprite 0x1c
    "11111110", --  113 - 0x71  :  254 - 0xfe
    "11100010", --  114 - 0x72  :  226 - 0xe2
    "11111110", --  115 - 0x73  :  254 - 0xfe
    "11111110", --  116 - 0x74  :  254 - 0xfe -- Sprite 0x1d
    "11111110", --  117 - 0x75  :  254 - 0xfe
    "11100010", --  118 - 0x76  :  226 - 0xe2
    "11111110", --  119 - 0x77  :  254 - 0xfe
    "11111110", --  120 - 0x78  :  254 - 0xfe -- Sprite 0x1e
    "11111110", --  121 - 0x79  :  254 - 0xfe
    "11100010", --  122 - 0x7a  :  226 - 0xe2
    "11111110", --  123 - 0x7b  :  254 - 0xfe
    "11111110", --  124 - 0x7c  :  254 - 0xfe -- Sprite 0x1f
    "11111110", --  125 - 0x7d  :  254 - 0xfe
    "11100010", --  126 - 0x7e  :  226 - 0xe2
    "11111110", --  127 - 0x7f  :  254 - 0xfe
    "11111110", --  128 - 0x80  :  254 - 0xfe -- Sprite 0x20
    "11111110", --  129 - 0x81  :  254 - 0xfe
    "11100010", --  130 - 0x82  :  226 - 0xe2
    "11111110", --  131 - 0x83  :  254 - 0xfe
    "11111110", --  132 - 0x84  :  254 - 0xfe -- Sprite 0x21
    "11111110", --  133 - 0x85  :  254 - 0xfe
    "11100010", --  134 - 0x86  :  226 - 0xe2
    "11111110", --  135 - 0x87  :  254 - 0xfe
    "11111110", --  136 - 0x88  :  254 - 0xfe -- Sprite 0x22
    "11111110", --  137 - 0x89  :  254 - 0xfe
    "11100010", --  138 - 0x8a  :  226 - 0xe2
    "11111110", --  139 - 0x8b  :  254 - 0xfe
    "11111110", --  140 - 0x8c  :  254 - 0xfe -- Sprite 0x23
    "11111110", --  141 - 0x8d  :  254 - 0xfe
    "11100010", --  142 - 0x8e  :  226 - 0xe2
    "11111110", --  143 - 0x8f  :  254 - 0xfe
    "11111110", --  144 - 0x90  :  254 - 0xfe -- Sprite 0x24
    "11111110", --  145 - 0x91  :  254 - 0xfe
    "11100010", --  146 - 0x92  :  226 - 0xe2
    "11111110", --  147 - 0x93  :  254 - 0xfe
    "11111110", --  148 - 0x94  :  254 - 0xfe -- Sprite 0x25
    "11111110", --  149 - 0x95  :  254 - 0xfe
    "11100010", --  150 - 0x96  :  226 - 0xe2
    "11111110", --  151 - 0x97  :  254 - 0xfe
    "11111110", --  152 - 0x98  :  254 - 0xfe -- Sprite 0x26
    "11111110", --  153 - 0x99  :  254 - 0xfe
    "11100010", --  154 - 0x9a  :  226 - 0xe2
    "11111110", --  155 - 0x9b  :  254 - 0xfe
    "11111110", --  156 - 0x9c  :  254 - 0xfe -- Sprite 0x27
    "11111110", --  157 - 0x9d  :  254 - 0xfe
    "11100010", --  158 - 0x9e  :  226 - 0xe2
    "11111110", --  159 - 0x9f  :  254 - 0xfe
    "11111110", --  160 - 0xa0  :  254 - 0xfe -- Sprite 0x28
    "11111110", --  161 - 0xa1  :  254 - 0xfe
    "11100010", --  162 - 0xa2  :  226 - 0xe2
    "11111110", --  163 - 0xa3  :  254 - 0xfe
    "11111110", --  164 - 0xa4  :  254 - 0xfe -- Sprite 0x29
    "11111110", --  165 - 0xa5  :  254 - 0xfe
    "11100010", --  166 - 0xa6  :  226 - 0xe2
    "11111110", --  167 - 0xa7  :  254 - 0xfe
    "11111110", --  168 - 0xa8  :  254 - 0xfe -- Sprite 0x2a
    "11111110", --  169 - 0xa9  :  254 - 0xfe
    "11100010", --  170 - 0xaa  :  226 - 0xe2
    "11111110", --  171 - 0xab  :  254 - 0xfe
    "11111110", --  172 - 0xac  :  254 - 0xfe -- Sprite 0x2b
    "11111110", --  173 - 0xad  :  254 - 0xfe
    "11100010", --  174 - 0xae  :  226 - 0xe2
    "11111110", --  175 - 0xaf  :  254 - 0xfe
    "11111110", --  176 - 0xb0  :  254 - 0xfe -- Sprite 0x2c
    "11111110", --  177 - 0xb1  :  254 - 0xfe
    "11100010", --  178 - 0xb2  :  226 - 0xe2
    "11111110", --  179 - 0xb3  :  254 - 0xfe
    "11111110", --  180 - 0xb4  :  254 - 0xfe -- Sprite 0x2d
    "11111110", --  181 - 0xb5  :  254 - 0xfe
    "11100010", --  182 - 0xb6  :  226 - 0xe2
    "11111110", --  183 - 0xb7  :  254 - 0xfe
    "11111110", --  184 - 0xb8  :  254 - 0xfe -- Sprite 0x2e
    "11111110", --  185 - 0xb9  :  254 - 0xfe
    "11100010", --  186 - 0xba  :  226 - 0xe2
    "11111110", --  187 - 0xbb  :  254 - 0xfe
    "11111110", --  188 - 0xbc  :  254 - 0xfe -- Sprite 0x2f
    "11111110", --  189 - 0xbd  :  254 - 0xfe
    "11100010", --  190 - 0xbe  :  226 - 0xe2
    "11111110", --  191 - 0xbf  :  254 - 0xfe
    "11111110", --  192 - 0xc0  :  254 - 0xfe -- Sprite 0x30
    "11111110", --  193 - 0xc1  :  254 - 0xfe
    "11100010", --  194 - 0xc2  :  226 - 0xe2
    "11111110", --  195 - 0xc3  :  254 - 0xfe
    "11111110", --  196 - 0xc4  :  254 - 0xfe -- Sprite 0x31
    "11111110", --  197 - 0xc5  :  254 - 0xfe
    "11100010", --  198 - 0xc6  :  226 - 0xe2
    "11111110", --  199 - 0xc7  :  254 - 0xfe
    "11111110", --  200 - 0xc8  :  254 - 0xfe -- Sprite 0x32
    "11111110", --  201 - 0xc9  :  254 - 0xfe
    "11100010", --  202 - 0xca  :  226 - 0xe2
    "11111110", --  203 - 0xcb  :  254 - 0xfe
    "11111110", --  204 - 0xcc  :  254 - 0xfe -- Sprite 0x33
    "11111110", --  205 - 0xcd  :  254 - 0xfe
    "11100010", --  206 - 0xce  :  226 - 0xe2
    "11111110", --  207 - 0xcf  :  254 - 0xfe
    "11111110", --  208 - 0xd0  :  254 - 0xfe -- Sprite 0x34
    "11111110", --  209 - 0xd1  :  254 - 0xfe
    "11100010", --  210 - 0xd2  :  226 - 0xe2
    "11111110", --  211 - 0xd3  :  254 - 0xfe
    "11111110", --  212 - 0xd4  :  254 - 0xfe -- Sprite 0x35
    "11111110", --  213 - 0xd5  :  254 - 0xfe
    "11100010", --  214 - 0xd6  :  226 - 0xe2
    "11111110", --  215 - 0xd7  :  254 - 0xfe
    "11111110", --  216 - 0xd8  :  254 - 0xfe -- Sprite 0x36
    "11111110", --  217 - 0xd9  :  254 - 0xfe
    "11100010", --  218 - 0xda  :  226 - 0xe2
    "11111110", --  219 - 0xdb  :  254 - 0xfe
    "11111110", --  220 - 0xdc  :  254 - 0xfe -- Sprite 0x37
    "11111110", --  221 - 0xdd  :  254 - 0xfe
    "11100010", --  222 - 0xde  :  226 - 0xe2
    "11111110", --  223 - 0xdf  :  254 - 0xfe
    "11111110", --  224 - 0xe0  :  254 - 0xfe -- Sprite 0x38
    "11111110", --  225 - 0xe1  :  254 - 0xfe
    "11100010", --  226 - 0xe2  :  226 - 0xe2
    "11111110", --  227 - 0xe3  :  254 - 0xfe
    "11111110", --  228 - 0xe4  :  254 - 0xfe -- Sprite 0x39
    "11111110", --  229 - 0xe5  :  254 - 0xfe
    "11100010", --  230 - 0xe6  :  226 - 0xe2
    "11111110", --  231 - 0xe7  :  254 - 0xfe
    "11111110", --  232 - 0xe8  :  254 - 0xfe -- Sprite 0x3a
    "11111110", --  233 - 0xe9  :  254 - 0xfe
    "11100010", --  234 - 0xea  :  226 - 0xe2
    "11111110", --  235 - 0xeb  :  254 - 0xfe
    "11111110", --  236 - 0xec  :  254 - 0xfe -- Sprite 0x3b
    "11111110", --  237 - 0xed  :  254 - 0xfe
    "11100010", --  238 - 0xee  :  226 - 0xe2
    "11111110", --  239 - 0xef  :  254 - 0xfe
    "11111110", --  240 - 0xf0  :  254 - 0xfe -- Sprite 0x3c
    "11111110", --  241 - 0xf1  :  254 - 0xfe
    "11100010", --  242 - 0xf2  :  226 - 0xe2
    "11111110", --  243 - 0xf3  :  254 - 0xfe
    "11111110", --  244 - 0xf4  :  254 - 0xfe -- Sprite 0x3d
    "11111110", --  245 - 0xf5  :  254 - 0xfe
    "11100010", --  246 - 0xf6  :  226 - 0xe2
    "11111110", --  247 - 0xf7  :  254 - 0xfe
    "11111110", --  248 - 0xf8  :  254 - 0xfe -- Sprite 0x3e
    "11111110", --  249 - 0xf9  :  254 - 0xfe
    "11100010", --  250 - 0xfa  :  226 - 0xe2
    "11111110", --  251 - 0xfb  :  254 - 0xfe
    "11111110", --  252 - 0xfc  :  254 - 0xfe -- Sprite 0x3f
    "11111110", --  253 - 0xfd  :  254 - 0xfe
    "11100010", --  254 - 0xfe  :  226 - 0xe2
    "11111110"  --  255 - 0xff  :  254 - 0xfe
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
