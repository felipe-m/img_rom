--- Autcmatically generated VHDL ROM from a NES memory file----
---   PATTERN TABLE WITH ONLY ONE COLOR PLANE
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


---  Original memory dump file name: nova_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_NOVA_color0 is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(12-1 downto 0);  --4096 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_NOVA_color0;

architecture BEHAVIORAL of ROM_PTABLE_NOVA_color0 is
  signal addr_int  : natural range 0 to 2**12-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Sprite pattern Table
    "11111111", --    0 -  0x0  :  255 - 0xff -- Sprite 0x0
    "11111111", --    1 -  0x1  :  255 - 0xff
    "11000000", --    2 -  0x2  :  192 - 0xc0
    "11000000", --    3 -  0x3  :  192 - 0xc0
    "11000000", --    4 -  0x4  :  192 - 0xc0
    "11000000", --    5 -  0x5  :  192 - 0xc0
    "11010101", --    6 -  0x6  :  213 - 0xd5
    "11111111", --    7 -  0x7  :  255 - 0xff
    "11111111", --    8 -  0x8  :  255 - 0xff -- Sprite 0x1
    "11111111", --    9 -  0x9  :  255 - 0xff
    "11001110", --   10 -  0xa  :  206 - 0xce
    "11000110", --   11 -  0xb  :  198 - 0xc6
    "11001110", --   12 -  0xc  :  206 - 0xce
    "11000110", --   13 -  0xd  :  198 - 0xc6
    "11101110", --   14 -  0xe  :  238 - 0xee
    "11111111", --   15 -  0xf  :  255 - 0xff
    "11111111", --   16 - 0x10  :  255 - 0xff -- Sprite 0x2
    "11111111", --   17 - 0x11  :  255 - 0xff
    "01110001", --   18 - 0x12  :  113 - 0x71
    "00110011", --   19 - 0x13  :   51 - 0x33
    "01110001", --   20 - 0x14  :  113 - 0x71
    "00110011", --   21 - 0x15  :   51 - 0x33
    "01110101", --   22 - 0x16  :  117 - 0x75
    "11111111", --   23 - 0x17  :  255 - 0xff
    "11111111", --   24 - 0x18  :  255 - 0xff -- Sprite 0x3
    "11111111", --   25 - 0x19  :  255 - 0xff
    "00000011", --   26 - 0x1a  :    3 - 0x3
    "00000001", --   27 - 0x1b  :    1 - 0x1
    "00000011", --   28 - 0x1c  :    3 - 0x3
    "00000001", --   29 - 0x1d  :    1 - 0x1
    "10101011", --   30 - 0x1e  :  171 - 0xab
    "11111111", --   31 - 0x1f  :  255 - 0xff
    "11111111", --   32 - 0x20  :  255 - 0xff -- Sprite 0x4
    "11111111", --   33 - 0x21  :  255 - 0xff
    "11100000", --   34 - 0x22  :  224 - 0xe0
    "11000110", --   35 - 0x23  :  198 - 0xc6
    "11000110", --   36 - 0x24  :  198 - 0xc6
    "11110110", --   37 - 0x25  :  246 - 0xf6
    "11110000", --   38 - 0x26  :  240 - 0xf0
    "11110001", --   39 - 0x27  :  241 - 0xf1
    "11000111", --   40 - 0x28  :  199 - 0xc7 -- Sprite 0x5
    "11001111", --   41 - 0x29  :  207 - 0xcf
    "11011111", --   42 - 0x2a  :  223 - 0xdf
    "11011111", --   43 - 0x2b  :  223 - 0xdf
    "11001110", --   44 - 0x2c  :  206 - 0xce
    "11100000", --   45 - 0x2d  :  224 - 0xe0
    "11111111", --   46 - 0x2e  :  255 - 0xff
    "11111111", --   47 - 0x2f  :  255 - 0xff
    "11111111", --   48 - 0x30  :  255 - 0xff -- Sprite 0x6
    "11111111", --   49 - 0x31  :  255 - 0xff
    "00000111", --   50 - 0x32  :    7 - 0x7
    "01100011", --   51 - 0x33  :   99 - 0x63
    "01100011", --   52 - 0x34  :   99 - 0x63
    "01101111", --   53 - 0x35  :  111 - 0x6f
    "00001111", --   54 - 0x36  :   15 - 0xf
    "10001111", --   55 - 0x37  :  143 - 0x8f
    "11100011", --   56 - 0x38  :  227 - 0xe3 -- Sprite 0x7
    "11110011", --   57 - 0x39  :  243 - 0xf3
    "11111011", --   58 - 0x3a  :  251 - 0xfb
    "11111011", --   59 - 0x3b  :  251 - 0xfb
    "01110011", --   60 - 0x3c  :  115 - 0x73
    "00000111", --   61 - 0x3d  :    7 - 0x7
    "11111111", --   62 - 0x3e  :  255 - 0xff
    "11111111", --   63 - 0x3f  :  255 - 0xff
    "11111111", --   64 - 0x40  :  255 - 0xff -- Sprite 0x8
    "11010101", --   65 - 0x41  :  213 - 0xd5
    "10101010", --   66 - 0x42  :  170 - 0xaa
    "11010101", --   67 - 0x43  :  213 - 0xd5
    "10101010", --   68 - 0x44  :  170 - 0xaa
    "11010101", --   69 - 0x45  :  213 - 0xd5
    "10101010", --   70 - 0x46  :  170 - 0xaa
    "11010101", --   71 - 0x47  :  213 - 0xd5
    "10101010", --   72 - 0x48  :  170 - 0xaa -- Sprite 0x9
    "11010101", --   73 - 0x49  :  213 - 0xd5
    "10101010", --   74 - 0x4a  :  170 - 0xaa
    "11010101", --   75 - 0x4b  :  213 - 0xd5
    "10101010", --   76 - 0x4c  :  170 - 0xaa
    "11110101", --   77 - 0x4d  :  245 - 0xf5
    "10101010", --   78 - 0x4e  :  170 - 0xaa
    "11111111", --   79 - 0x4f  :  255 - 0xff
    "11111111", --   80 - 0x50  :  255 - 0xff -- Sprite 0xa
    "01010101", --   81 - 0x51  :   85 - 0x55
    "10101111", --   82 - 0x52  :  175 - 0xaf
    "01010101", --   83 - 0x53  :   85 - 0x55
    "10101011", --   84 - 0x54  :  171 - 0xab
    "01010101", --   85 - 0x55  :   85 - 0x55
    "10101011", --   86 - 0x56  :  171 - 0xab
    "01010101", --   87 - 0x57  :   85 - 0x55
    "10101011", --   88 - 0x58  :  171 - 0xab -- Sprite 0xb
    "01010101", --   89 - 0x59  :   85 - 0x55
    "10101011", --   90 - 0x5a  :  171 - 0xab
    "01010101", --   91 - 0x5b  :   85 - 0x55
    "10101011", --   92 - 0x5c  :  171 - 0xab
    "01010101", --   93 - 0x5d  :   85 - 0x55
    "10101011", --   94 - 0x5e  :  171 - 0xab
    "11111111", --   95 - 0x5f  :  255 - 0xff
    "11111111", --   96 - 0x60  :  255 - 0xff -- Sprite 0xc
    "11010101", --   97 - 0x61  :  213 - 0xd5
    "10100000", --   98 - 0x62  :  160 - 0xa0
    "11010000", --   99 - 0x63  :  208 - 0xd0
    "10001111", --  100 - 0x64  :  143 - 0x8f
    "11001000", --  101 - 0x65  :  200 - 0xc8
    "10001000", --  102 - 0x66  :  136 - 0x88
    "11001000", --  103 - 0x67  :  200 - 0xc8
    "10001000", --  104 - 0x68  :  136 - 0x88 -- Sprite 0xd
    "11001000", --  105 - 0x69  :  200 - 0xc8
    "10001000", --  106 - 0x6a  :  136 - 0x88
    "11001111", --  107 - 0x6b  :  207 - 0xcf
    "10010000", --  108 - 0x6c  :  144 - 0x90
    "11100000", --  109 - 0x6d  :  224 - 0xe0
    "11101010", --  110 - 0x6e  :  234 - 0xea
    "11111111", --  111 - 0x6f  :  255 - 0xff
    "11111111", --  112 - 0x70  :  255 - 0xff -- Sprite 0xe
    "01011011", --  113 - 0x71  :   91 - 0x5b
    "00000111", --  114 - 0x72  :    7 - 0x7
    "00001001", --  115 - 0x73  :    9 - 0x9
    "11110011", --  116 - 0x74  :  243 - 0xf3
    "00010001", --  117 - 0x75  :   17 - 0x11
    "00010011", --  118 - 0x76  :   19 - 0x13
    "00010001", --  119 - 0x77  :   17 - 0x11
    "00010011", --  120 - 0x78  :   19 - 0x13 -- Sprite 0xf
    "00010001", --  121 - 0x79  :   17 - 0x11
    "00010011", --  122 - 0x7a  :   19 - 0x13
    "11110001", --  123 - 0x7b  :  241 - 0xf1
    "00001011", --  124 - 0x7c  :   11 - 0xb
    "00000101", --  125 - 0x7d  :    5 - 0x5
    "10101011", --  126 - 0x7e  :  171 - 0xab
    "11111111", --  127 - 0x7f  :  255 - 0xff
    "11010000", --  128 - 0x80  :  208 - 0xd0 -- Sprite 0x10
    "10010000", --  129 - 0x81  :  144 - 0x90
    "11011111", --  130 - 0x82  :  223 - 0xdf
    "10011010", --  131 - 0x83  :  154 - 0x9a
    "11010101", --  132 - 0x84  :  213 - 0xd5
    "10011111", --  133 - 0x85  :  159 - 0x9f
    "11010000", --  134 - 0x86  :  208 - 0xd0
    "10010000", --  135 - 0x87  :  144 - 0x90
    "00001001", --  136 - 0x88  :    9 - 0x9 -- Sprite 0x11
    "00001011", --  137 - 0x89  :   11 - 0xb
    "11111001", --  138 - 0x8a  :  249 - 0xf9
    "10101011", --  139 - 0x8b  :  171 - 0xab
    "01011001", --  140 - 0x8c  :   89 - 0x59
    "11111011", --  141 - 0x8d  :  251 - 0xfb
    "00001001", --  142 - 0x8e  :    9 - 0x9
    "00001011", --  143 - 0x8f  :   11 - 0xb
    "00011000", --  144 - 0x90  :   24 - 0x18 -- Sprite 0x12
    "00010100", --  145 - 0x91  :   20 - 0x14
    "00010100", --  146 - 0x92  :   20 - 0x14
    "00111010", --  147 - 0x93  :   58 - 0x3a
    "00111010", --  148 - 0x94  :   58 - 0x3a
    "01111010", --  149 - 0x95  :  122 - 0x7a
    "01111010", --  150 - 0x96  :  122 - 0x7a
    "01111010", --  151 - 0x97  :  122 - 0x7a
    "11111011", --  152 - 0x98  :  251 - 0xfb -- Sprite 0x13
    "11111101", --  153 - 0x99  :  253 - 0xfd
    "11111101", --  154 - 0x9a  :  253 - 0xfd
    "11111101", --  155 - 0x9b  :  253 - 0xfd
    "11111101", --  156 - 0x9c  :  253 - 0xfd
    "11111101", --  157 - 0x9d  :  253 - 0xfd
    "10000001", --  158 - 0x9e  :  129 - 0x81
    "11111111", --  159 - 0x9f  :  255 - 0xff
    "00000000", --  160 - 0xa0  :    0 - 0x0 -- Sprite 0x14
    "00000111", --  161 - 0xa1  :    7 - 0x7
    "00000010", --  162 - 0xa2  :    2 - 0x2
    "00000100", --  163 - 0xa3  :    4 - 0x4
    "00000011", --  164 - 0xa4  :    3 - 0x3
    "00000011", --  165 - 0xa5  :    3 - 0x3
    "00001101", --  166 - 0xa6  :   13 - 0xd
    "00010111", --  167 - 0xa7  :   23 - 0x17
    "00101111", --  168 - 0xa8  :   47 - 0x2f -- Sprite 0x15
    "01001111", --  169 - 0xa9  :   79 - 0x4f
    "01001111", --  170 - 0xaa  :   79 - 0x4f
    "01001111", --  171 - 0xab  :   79 - 0x4f
    "01001111", --  172 - 0xac  :   79 - 0x4f
    "00100111", --  173 - 0xad  :   39 - 0x27
    "00010000", --  174 - 0xae  :   16 - 0x10
    "00001111", --  175 - 0xaf  :   15 - 0xf
    "00000000", --  176 - 0xb0  :    0 - 0x0 -- Sprite 0x16
    "11100000", --  177 - 0xb1  :  224 - 0xe0
    "10100000", --  178 - 0xb2  :  160 - 0xa0
    "00100000", --  179 - 0xb3  :   32 - 0x20
    "11000000", --  180 - 0xb4  :  192 - 0xc0
    "01000000", --  181 - 0xb5  :   64 - 0x40
    "00110000", --  182 - 0xb6  :   48 - 0x30
    "11101000", --  183 - 0xb7  :  232 - 0xe8
    "11110100", --  184 - 0xb8  :  244 - 0xf4 -- Sprite 0x17
    "11110010", --  185 - 0xb9  :  242 - 0xf2
    "11110010", --  186 - 0xba  :  242 - 0xf2
    "11110010", --  187 - 0xbb  :  242 - 0xf2
    "11110010", --  188 - 0xbc  :  242 - 0xf2
    "11100100", --  189 - 0xbd  :  228 - 0xe4
    "00001000", --  190 - 0xbe  :    8 - 0x8
    "11110000", --  191 - 0xbf  :  240 - 0xf0
    "00111111", --  192 - 0xc0  :   63 - 0x3f -- Sprite 0x18
    "01000000", --  193 - 0xc1  :   64 - 0x40
    "01000000", --  194 - 0xc2  :   64 - 0x40
    "10000000", --  195 - 0xc3  :  128 - 0x80
    "10000000", --  196 - 0xc4  :  128 - 0x80
    "01111111", --  197 - 0xc5  :  127 - 0x7f
    "00000001", --  198 - 0xc6  :    1 - 0x1
    "01111111", --  199 - 0xc7  :  127 - 0x7f
    "11111100", --  200 - 0xc8  :  252 - 0xfc -- Sprite 0x19
    "00000010", --  201 - 0xc9  :    2 - 0x2
    "00000010", --  202 - 0xca  :    2 - 0x2
    "00000001", --  203 - 0xcb  :    1 - 0x1
    "00000001", --  204 - 0xcc  :    1 - 0x1
    "11111110", --  205 - 0xcd  :  254 - 0xfe
    "10000000", --  206 - 0xce  :  128 - 0x80
    "11111110", --  207 - 0xcf  :  254 - 0xfe
    "00000000", --  208 - 0xd0  :    0 - 0x0 -- Sprite 0x1a
    "00000000", --  209 - 0xd1  :    0 - 0x0
    "00111111", --  210 - 0xd2  :   63 - 0x3f
    "01000000", --  211 - 0xd3  :   64 - 0x40
    "01000000", --  212 - 0xd4  :   64 - 0x40
    "10000000", --  213 - 0xd5  :  128 - 0x80
    "10000000", --  214 - 0xd6  :  128 - 0x80
    "01111111", --  215 - 0xd7  :  127 - 0x7f
    "00000000", --  216 - 0xd8  :    0 - 0x0 -- Sprite 0x1b
    "00000000", --  217 - 0xd9  :    0 - 0x0
    "11111100", --  218 - 0xda  :  252 - 0xfc
    "00000010", --  219 - 0xdb  :    2 - 0x2
    "00000010", --  220 - 0xdc  :    2 - 0x2
    "00000001", --  221 - 0xdd  :    1 - 0x1
    "00000001", --  222 - 0xde  :    1 - 0x1
    "11111110", --  223 - 0xdf  :  254 - 0xfe
    "01111111", --  224 - 0xe0  :  127 - 0x7f -- Sprite 0x1c
    "10000000", --  225 - 0xe1  :  128 - 0x80
    "10000000", --  226 - 0xe2  :  128 - 0x80
    "10000000", --  227 - 0xe3  :  128 - 0x80
    "10011011", --  228 - 0xe4  :  155 - 0x9b
    "10100100", --  229 - 0xe5  :  164 - 0xa4
    "10100110", --  230 - 0xe6  :  166 - 0xa6
    "10000000", --  231 - 0xe7  :  128 - 0x80
    "10000000", --  232 - 0xe8  :  128 - 0x80 -- Sprite 0x1d
    "01111111", --  233 - 0xe9  :  127 - 0x7f
    "00000010", --  234 - 0xea  :    2 - 0x2
    "00000010", --  235 - 0xeb  :    2 - 0x2
    "00000010", --  236 - 0xec  :    2 - 0x2
    "00000010", --  237 - 0xed  :    2 - 0x2
    "00000010", --  238 - 0xee  :    2 - 0x2
    "00001111", --  239 - 0xef  :   15 - 0xf
    "11111110", --  240 - 0xf0  :  254 - 0xfe -- Sprite 0x1e
    "00000001", --  241 - 0xf1  :    1 - 0x1
    "00000001", --  242 - 0xf2  :    1 - 0x1
    "00000001", --  243 - 0xf3  :    1 - 0x1
    "01000001", --  244 - 0xf4  :   65 - 0x41
    "11110101", --  245 - 0xf5  :  245 - 0xf5
    "00011101", --  246 - 0xf6  :   29 - 0x1d
    "00000001", --  247 - 0xf7  :    1 - 0x1
    "00000001", --  248 - 0xf8  :    1 - 0x1 -- Sprite 0x1f
    "11111110", --  249 - 0xf9  :  254 - 0xfe
    "01000000", --  250 - 0xfa  :   64 - 0x40
    "01000000", --  251 - 0xfb  :   64 - 0x40
    "01000000", --  252 - 0xfc  :   64 - 0x40
    "01000000", --  253 - 0xfd  :   64 - 0x40
    "01000000", --  254 - 0xfe  :   64 - 0x40
    "11110000", --  255 - 0xff  :  240 - 0xf0
    "00000111", --  256 - 0x100  :    7 - 0x7 -- Sprite 0x20
    "00011111", --  257 - 0x101  :   31 - 0x1f
    "00111111", --  258 - 0x102  :   63 - 0x3f
    "01111111", --  259 - 0x103  :  127 - 0x7f
    "01111111", --  260 - 0x104  :  127 - 0x7f
    "11111111", --  261 - 0x105  :  255 - 0xff
    "11111111", --  262 - 0x106  :  255 - 0xff
    "11111111", --  263 - 0x107  :  255 - 0xff
    "11100000", --  264 - 0x108  :  224 - 0xe0 -- Sprite 0x21
    "11111000", --  265 - 0x109  :  248 - 0xf8
    "11111100", --  266 - 0x10a  :  252 - 0xfc
    "11111110", --  267 - 0x10b  :  254 - 0xfe
    "11111110", --  268 - 0x10c  :  254 - 0xfe
    "11111111", --  269 - 0x10d  :  255 - 0xff
    "11111111", --  270 - 0x10e  :  255 - 0xff
    "11111111", --  271 - 0x10f  :  255 - 0xff
    "00000111", --  272 - 0x110  :    7 - 0x7 -- Sprite 0x22
    "00011111", --  273 - 0x111  :   31 - 0x1f
    "00111111", --  274 - 0x112  :   63 - 0x3f
    "01111111", --  275 - 0x113  :  127 - 0x7f
    "01111111", --  276 - 0x114  :  127 - 0x7f
    "11111111", --  277 - 0x115  :  255 - 0xff
    "11111111", --  278 - 0x116  :  255 - 0xff
    "11111111", --  279 - 0x117  :  255 - 0xff
    "11100000", --  280 - 0x118  :  224 - 0xe0 -- Sprite 0x23
    "11111000", --  281 - 0x119  :  248 - 0xf8
    "11111100", --  282 - 0x11a  :  252 - 0xfc
    "11111110", --  283 - 0x11b  :  254 - 0xfe
    "11111110", --  284 - 0x11c  :  254 - 0xfe
    "11111111", --  285 - 0x11d  :  255 - 0xff
    "11111111", --  286 - 0x11e  :  255 - 0xff
    "11111111", --  287 - 0x11f  :  255 - 0xff
    "00000000", --  288 - 0x120  :    0 - 0x0 -- Sprite 0x24
    "00000000", --  289 - 0x121  :    0 - 0x0
    "00000000", --  290 - 0x122  :    0 - 0x0
    "00000000", --  291 - 0x123  :    0 - 0x0
    "00000000", --  292 - 0x124  :    0 - 0x0
    "00000000", --  293 - 0x125  :    0 - 0x0
    "00000000", --  294 - 0x126  :    0 - 0x0
    "00000000", --  295 - 0x127  :    0 - 0x0
    "00101111", --  296 - 0x128  :   47 - 0x2f -- Sprite 0x25
    "01001111", --  297 - 0x129  :   79 - 0x4f
    "01001111", --  298 - 0x12a  :   79 - 0x4f
    "01001111", --  299 - 0x12b  :   79 - 0x4f
    "01001111", --  300 - 0x12c  :   79 - 0x4f
    "00100111", --  301 - 0x12d  :   39 - 0x27
    "00010000", --  302 - 0x12e  :   16 - 0x10
    "00001111", --  303 - 0x12f  :   15 - 0xf
    "00000000", --  304 - 0x130  :    0 - 0x0 -- Sprite 0x26
    "11100000", --  305 - 0x131  :  224 - 0xe0
    "10100000", --  306 - 0x132  :  160 - 0xa0
    "00100000", --  307 - 0x133  :   32 - 0x20
    "11000000", --  308 - 0x134  :  192 - 0xc0
    "01000000", --  309 - 0x135  :   64 - 0x40
    "00110000", --  310 - 0x136  :   48 - 0x30
    "11101000", --  311 - 0x137  :  232 - 0xe8
    "11110100", --  312 - 0x138  :  244 - 0xf4 -- Sprite 0x27
    "11110010", --  313 - 0x139  :  242 - 0xf2
    "11110010", --  314 - 0x13a  :  242 - 0xf2
    "11110010", --  315 - 0x13b  :  242 - 0xf2
    "11110010", --  316 - 0x13c  :  242 - 0xf2
    "11100100", --  317 - 0x13d  :  228 - 0xe4
    "00001000", --  318 - 0x13e  :    8 - 0x8
    "11110000", --  319 - 0x13f  :  240 - 0xf0
    "11111111", --  320 - 0x140  :  255 - 0xff -- Sprite 0x28
    "11010101", --  321 - 0x141  :  213 - 0xd5
    "10100011", --  322 - 0x142  :  163 - 0xa3
    "11010111", --  323 - 0x143  :  215 - 0xd7
    "10001111", --  324 - 0x144  :  143 - 0x8f
    "11001111", --  325 - 0x145  :  207 - 0xcf
    "10001011", --  326 - 0x146  :  139 - 0x8b
    "11001011", --  327 - 0x147  :  203 - 0xcb
    "10001111", --  328 - 0x148  :  143 - 0x8f -- Sprite 0x29
    "11001111", --  329 - 0x149  :  207 - 0xcf
    "10001111", --  330 - 0x14a  :  143 - 0x8f
    "11001111", --  331 - 0x14b  :  207 - 0xcf
    "10010000", --  332 - 0x14c  :  144 - 0x90
    "11100000", --  333 - 0x14d  :  224 - 0xe0
    "11101010", --  334 - 0x14e  :  234 - 0xea
    "11111111", --  335 - 0x14f  :  255 - 0xff
    "11111111", --  336 - 0x150  :  255 - 0xff -- Sprite 0x2a
    "11011011", --  337 - 0x151  :  219 - 0xdb
    "11000111", --  338 - 0x152  :  199 - 0xc7
    "11101001", --  339 - 0x153  :  233 - 0xe9
    "11110011", --  340 - 0x154  :  243 - 0xf3
    "11110001", --  341 - 0x155  :  241 - 0xf1
    "11010011", --  342 - 0x156  :  211 - 0xd3
    "11010001", --  343 - 0x157  :  209 - 0xd1
    "11110011", --  344 - 0x158  :  243 - 0xf3 -- Sprite 0x2b
    "11110001", --  345 - 0x159  :  241 - 0xf1
    "11110011", --  346 - 0x15a  :  243 - 0xf3
    "11110001", --  347 - 0x15b  :  241 - 0xf1
    "00001011", --  348 - 0x15c  :   11 - 0xb
    "00000101", --  349 - 0x15d  :    5 - 0x5
    "10101011", --  350 - 0x15e  :  171 - 0xab
    "11111111", --  351 - 0x15f  :  255 - 0xff
    "00000000", --  352 - 0x160  :    0 - 0x0 -- Sprite 0x2c
    "00000000", --  353 - 0x161  :    0 - 0x0
    "00000000", --  354 - 0x162  :    0 - 0x0
    "00000000", --  355 - 0x163  :    0 - 0x0
    "00000000", --  356 - 0x164  :    0 - 0x0
    "00000000", --  357 - 0x165  :    0 - 0x0
    "00000000", --  358 - 0x166  :    0 - 0x0
    "00000000", --  359 - 0x167  :    0 - 0x0
    "00101111", --  360 - 0x168  :   47 - 0x2f -- Sprite 0x2d
    "01001111", --  361 - 0x169  :   79 - 0x4f
    "01001111", --  362 - 0x16a  :   79 - 0x4f
    "01001111", --  363 - 0x16b  :   79 - 0x4f
    "01001111", --  364 - 0x16c  :   79 - 0x4f
    "00100111", --  365 - 0x16d  :   39 - 0x27
    "00010000", --  366 - 0x16e  :   16 - 0x10
    "00001111", --  367 - 0x16f  :   15 - 0xf
    "00000000", --  368 - 0x170  :    0 - 0x0 -- Sprite 0x2e
    "00000000", --  369 - 0x171  :    0 - 0x0
    "00000000", --  370 - 0x172  :    0 - 0x0
    "00000000", --  371 - 0x173  :    0 - 0x0
    "00000000", --  372 - 0x174  :    0 - 0x0
    "00000000", --  373 - 0x175  :    0 - 0x0
    "00000000", --  374 - 0x176  :    0 - 0x0
    "00000000", --  375 - 0x177  :    0 - 0x0
    "11110100", --  376 - 0x178  :  244 - 0xf4 -- Sprite 0x2f
    "11110010", --  377 - 0x179  :  242 - 0xf2
    "11110010", --  378 - 0x17a  :  242 - 0xf2
    "11110010", --  379 - 0x17b  :  242 - 0xf2
    "11110010", --  380 - 0x17c  :  242 - 0xf2
    "11100100", --  381 - 0x17d  :  228 - 0xe4
    "00001000", --  382 - 0x17e  :    8 - 0x8
    "11110000", --  383 - 0x17f  :  240 - 0xf0
    "00011000", --  384 - 0x180  :   24 - 0x18 -- Sprite 0x30
    "00100100", --  385 - 0x181  :   36 - 0x24
    "01000010", --  386 - 0x182  :   66 - 0x42
    "10100101", --  387 - 0x183  :  165 - 0xa5
    "11100111", --  388 - 0x184  :  231 - 0xe7
    "00100100", --  389 - 0x185  :   36 - 0x24
    "00100100", --  390 - 0x186  :   36 - 0x24
    "00111100", --  391 - 0x187  :   60 - 0x3c
    "00111100", --  392 - 0x188  :   60 - 0x3c -- Sprite 0x31
    "00100100", --  393 - 0x189  :   36 - 0x24
    "00100100", --  394 - 0x18a  :   36 - 0x24
    "01100110", --  395 - 0x18b  :  102 - 0x66
    "10100101", --  396 - 0x18c  :  165 - 0xa5
    "01000010", --  397 - 0x18d  :   66 - 0x42
    "00100100", --  398 - 0x18e  :   36 - 0x24
    "00011000", --  399 - 0x18f  :   24 - 0x18
    "00000010", --  400 - 0x190  :    2 - 0x2 -- Sprite 0x32
    "00000010", --  401 - 0x191  :    2 - 0x2
    "00000011", --  402 - 0x192  :    3 - 0x3
    "00000010", --  403 - 0x193  :    2 - 0x2
    "00000010", --  404 - 0x194  :    2 - 0x2
    "00000010", --  405 - 0x195  :    2 - 0x2
    "00000011", --  406 - 0x196  :    3 - 0x3
    "00000010", --  407 - 0x197  :    2 - 0x2
    "01000000", --  408 - 0x198  :   64 - 0x40 -- Sprite 0x33
    "11000000", --  409 - 0x199  :  192 - 0xc0
    "01000000", --  410 - 0x19a  :   64 - 0x40
    "01000000", --  411 - 0x19b  :   64 - 0x40
    "01000000", --  412 - 0x19c  :   64 - 0x40
    "11000000", --  413 - 0x19d  :  192 - 0xc0
    "01000000", --  414 - 0x19e  :   64 - 0x40
    "01000000", --  415 - 0x19f  :   64 - 0x40
    "00000000", --  416 - 0x1a0  :    0 - 0x0 -- Sprite 0x34
    "00011000", --  417 - 0x1a1  :   24 - 0x18
    "00111100", --  418 - 0x1a2  :   60 - 0x3c
    "01100010", --  419 - 0x1a3  :   98 - 0x62
    "01100001", --  420 - 0x1a4  :   97 - 0x61
    "11000000", --  421 - 0x1a5  :  192 - 0xc0
    "11000000", --  422 - 0x1a6  :  192 - 0xc0
    "11000000", --  423 - 0x1a7  :  192 - 0xc0
    "01100000", --  424 - 0x1a8  :   96 - 0x60 -- Sprite 0x35
    "01100000", --  425 - 0x1a9  :   96 - 0x60
    "00110000", --  426 - 0x1aa  :   48 - 0x30
    "00011000", --  427 - 0x1ab  :   24 - 0x18
    "00001100", --  428 - 0x1ac  :   12 - 0xc
    "00000110", --  429 - 0x1ad  :    6 - 0x6
    "00000010", --  430 - 0x1ae  :    2 - 0x2
    "00000001", --  431 - 0x1af  :    1 - 0x1
    "00000000", --  432 - 0x1b0  :    0 - 0x0 -- Sprite 0x36
    "00011000", --  433 - 0x1b1  :   24 - 0x18
    "00100100", --  434 - 0x1b2  :   36 - 0x24
    "01000010", --  435 - 0x1b3  :   66 - 0x42
    "10000010", --  436 - 0x1b4  :  130 - 0x82
    "00000001", --  437 - 0x1b5  :    1 - 0x1
    "00000001", --  438 - 0x1b6  :    1 - 0x1
    "00000001", --  439 - 0x1b7  :    1 - 0x1
    "00000010", --  440 - 0x1b8  :    2 - 0x2 -- Sprite 0x37
    "00000010", --  441 - 0x1b9  :    2 - 0x2
    "00000100", --  442 - 0x1ba  :    4 - 0x4
    "00001000", --  443 - 0x1bb  :    8 - 0x8
    "00010000", --  444 - 0x1bc  :   16 - 0x10
    "00100000", --  445 - 0x1bd  :   32 - 0x20
    "01000000", --  446 - 0x1be  :   64 - 0x40
    "10000000", --  447 - 0x1bf  :  128 - 0x80
    "00000000", --  448 - 0x1c0  :    0 - 0x0 -- Sprite 0x38
    "00000110", --  449 - 0x1c1  :    6 - 0x6
    "00001101", --  450 - 0x1c2  :   13 - 0xd
    "00001100", --  451 - 0x1c3  :   12 - 0xc
    "00001100", --  452 - 0x1c4  :   12 - 0xc
    "00000110", --  453 - 0x1c5  :    6 - 0x6
    "00000010", --  454 - 0x1c6  :    2 - 0x2
    "00000001", --  455 - 0x1c7  :    1 - 0x1
    "11111111", --  456 - 0x1c8  :  255 - 0xff -- Sprite 0x39
    "00000000", --  457 - 0x1c9  :    0 - 0x0
    "00000000", --  458 - 0x1ca  :    0 - 0x0
    "00000000", --  459 - 0x1cb  :    0 - 0x0
    "00000000", --  460 - 0x1cc  :    0 - 0x0
    "00000000", --  461 - 0x1cd  :    0 - 0x0
    "00000000", --  462 - 0x1ce  :    0 - 0x0
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "00000000", --  464 - 0x1d0  :    0 - 0x0 -- Sprite 0x3a
    "01100000", --  465 - 0x1d1  :   96 - 0x60
    "10010000", --  466 - 0x1d2  :  144 - 0x90
    "00010000", --  467 - 0x1d3  :   16 - 0x10
    "00010000", --  468 - 0x1d4  :   16 - 0x10
    "00100000", --  469 - 0x1d5  :   32 - 0x20
    "01000000", --  470 - 0x1d6  :   64 - 0x40
    "10000000", --  471 - 0x1d7  :  128 - 0x80
    "00000000", --  472 - 0x1d8  :    0 - 0x0 -- Sprite 0x3b
    "01010100", --  473 - 0x1d9  :   84 - 0x54
    "00000010", --  474 - 0x1da  :    2 - 0x2
    "01000000", --  475 - 0x1db  :   64 - 0x40
    "00000010", --  476 - 0x1dc  :    2 - 0x2
    "01000000", --  477 - 0x1dd  :   64 - 0x40
    "00101010", --  478 - 0x1de  :   42 - 0x2a
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "11111111", --  480 - 0x1e0  :  255 - 0xff -- Sprite 0x3c
    "11111111", --  481 - 0x1e1  :  255 - 0xff
    "11111111", --  482 - 0x1e2  :  255 - 0xff
    "11111111", --  483 - 0x1e3  :  255 - 0xff
    "11111111", --  484 - 0x1e4  :  255 - 0xff
    "11111111", --  485 - 0x1e5  :  255 - 0xff
    "11111111", --  486 - 0x1e6  :  255 - 0xff
    "11111111", --  487 - 0x1e7  :  255 - 0xff
    "00000000", --  488 - 0x1e8  :    0 - 0x0 -- Sprite 0x3d
    "00000000", --  489 - 0x1e9  :    0 - 0x0
    "00000000", --  490 - 0x1ea  :    0 - 0x0
    "00000000", --  491 - 0x1eb  :    0 - 0x0
    "00000000", --  492 - 0x1ec  :    0 - 0x0
    "00000000", --  493 - 0x1ed  :    0 - 0x0
    "00000000", --  494 - 0x1ee  :    0 - 0x0
    "00000000", --  495 - 0x1ef  :    0 - 0x0
    "11111111", --  496 - 0x1f0  :  255 - 0xff -- Sprite 0x3e
    "11111111", --  497 - 0x1f1  :  255 - 0xff
    "11111111", --  498 - 0x1f2  :  255 - 0xff
    "11111111", --  499 - 0x1f3  :  255 - 0xff
    "11111111", --  500 - 0x1f4  :  255 - 0xff
    "11111111", --  501 - 0x1f5  :  255 - 0xff
    "11111111", --  502 - 0x1f6  :  255 - 0xff
    "11111111", --  503 - 0x1f7  :  255 - 0xff
    "00000000", --  504 - 0x1f8  :    0 - 0x0 -- Sprite 0x3f
    "00000000", --  505 - 0x1f9  :    0 - 0x0
    "00000000", --  506 - 0x1fa  :    0 - 0x0
    "00000000", --  507 - 0x1fb  :    0 - 0x0
    "00000000", --  508 - 0x1fc  :    0 - 0x0
    "00000000", --  509 - 0x1fd  :    0 - 0x0
    "00000000", --  510 - 0x1fe  :    0 - 0x0
    "00000000", --  511 - 0x1ff  :    0 - 0x0
    "00111100", --  512 - 0x200  :   60 - 0x3c -- Sprite 0x40
    "01000010", --  513 - 0x201  :   66 - 0x42
    "10011001", --  514 - 0x202  :  153 - 0x99
    "10100101", --  515 - 0x203  :  165 - 0xa5
    "10100101", --  516 - 0x204  :  165 - 0xa5
    "10011010", --  517 - 0x205  :  154 - 0x9a
    "01000000", --  518 - 0x206  :   64 - 0x40
    "00111100", --  519 - 0x207  :   60 - 0x3c
    "00001100", --  520 - 0x208  :   12 - 0xc -- Sprite 0x41
    "00010010", --  521 - 0x209  :   18 - 0x12
    "00100010", --  522 - 0x20a  :   34 - 0x22
    "00100010", --  523 - 0x20b  :   34 - 0x22
    "01111110", --  524 - 0x20c  :  126 - 0x7e
    "00100010", --  525 - 0x20d  :   34 - 0x22
    "00100100", --  526 - 0x20e  :   36 - 0x24
    "00000000", --  527 - 0x20f  :    0 - 0x0
    "00111100", --  528 - 0x210  :   60 - 0x3c -- Sprite 0x42
    "01000010", --  529 - 0x211  :   66 - 0x42
    "01010010", --  530 - 0x212  :   82 - 0x52
    "00011100", --  531 - 0x213  :   28 - 0x1c
    "00010010", --  532 - 0x214  :   18 - 0x12
    "00110010", --  533 - 0x215  :   50 - 0x32
    "00011100", --  534 - 0x216  :   28 - 0x1c
    "00000000", --  535 - 0x217  :    0 - 0x0
    "00011000", --  536 - 0x218  :   24 - 0x18 -- Sprite 0x43
    "00100100", --  537 - 0x219  :   36 - 0x24
    "01010100", --  538 - 0x21a  :   84 - 0x54
    "01001000", --  539 - 0x21b  :   72 - 0x48
    "01000010", --  540 - 0x21c  :   66 - 0x42
    "00100100", --  541 - 0x21d  :   36 - 0x24
    "00011000", --  542 - 0x21e  :   24 - 0x18
    "00000000", --  543 - 0x21f  :    0 - 0x0
    "01011000", --  544 - 0x220  :   88 - 0x58 -- Sprite 0x44
    "11100100", --  545 - 0x221  :  228 - 0xe4
    "01000010", --  546 - 0x222  :   66 - 0x42
    "01000010", --  547 - 0x223  :   66 - 0x42
    "00100010", --  548 - 0x224  :   34 - 0x22
    "01100100", --  549 - 0x225  :  100 - 0x64
    "00111000", --  550 - 0x226  :   56 - 0x38
    "00000000", --  551 - 0x227  :    0 - 0x0
    "00011100", --  552 - 0x228  :   28 - 0x1c -- Sprite 0x45
    "00100000", --  553 - 0x229  :   32 - 0x20
    "00100000", --  554 - 0x22a  :   32 - 0x20
    "00101100", --  555 - 0x22b  :   44 - 0x2c
    "01110000", --  556 - 0x22c  :  112 - 0x70
    "00100010", --  557 - 0x22d  :   34 - 0x22
    "00011100", --  558 - 0x22e  :   28 - 0x1c
    "00000000", --  559 - 0x22f  :    0 - 0x0
    "00011100", --  560 - 0x230  :   28 - 0x1c -- Sprite 0x46
    "00100000", --  561 - 0x231  :   32 - 0x20
    "00100000", --  562 - 0x232  :   32 - 0x20
    "00101100", --  563 - 0x233  :   44 - 0x2c
    "01110000", --  564 - 0x234  :  112 - 0x70
    "00010000", --  565 - 0x235  :   16 - 0x10
    "00010000", --  566 - 0x236  :   16 - 0x10
    "00000000", --  567 - 0x237  :    0 - 0x0
    "00011000", --  568 - 0x238  :   24 - 0x18 -- Sprite 0x47
    "00100100", --  569 - 0x239  :   36 - 0x24
    "01000000", --  570 - 0x23a  :   64 - 0x40
    "01001110", --  571 - 0x23b  :   78 - 0x4e
    "01000010", --  572 - 0x23c  :   66 - 0x42
    "00100100", --  573 - 0x23d  :   36 - 0x24
    "00011000", --  574 - 0x23e  :   24 - 0x18
    "00000000", --  575 - 0x23f  :    0 - 0x0
    "00100000", --  576 - 0x240  :   32 - 0x20 -- Sprite 0x48
    "01000100", --  577 - 0x241  :   68 - 0x44
    "01000100", --  578 - 0x242  :   68 - 0x44
    "01000100", --  579 - 0x243  :   68 - 0x44
    "11111100", --  580 - 0x244  :  252 - 0xfc
    "01000100", --  581 - 0x245  :   68 - 0x44
    "01001000", --  582 - 0x246  :   72 - 0x48
    "00000000", --  583 - 0x247  :    0 - 0x0
    "00010000", --  584 - 0x248  :   16 - 0x10 -- Sprite 0x49
    "00010000", --  585 - 0x249  :   16 - 0x10
    "00010000", --  586 - 0x24a  :   16 - 0x10
    "00010000", --  587 - 0x24b  :   16 - 0x10
    "00010000", --  588 - 0x24c  :   16 - 0x10
    "00001000", --  589 - 0x24d  :    8 - 0x8
    "00001000", --  590 - 0x24e  :    8 - 0x8
    "00000000", --  591 - 0x24f  :    0 - 0x0
    "00001000", --  592 - 0x250  :    8 - 0x8 -- Sprite 0x4a
    "00001000", --  593 - 0x251  :    8 - 0x8
    "00000100", --  594 - 0x252  :    4 - 0x4
    "00000100", --  595 - 0x253  :    4 - 0x4
    "01000100", --  596 - 0x254  :   68 - 0x44
    "01001000", --  597 - 0x255  :   72 - 0x48
    "00110000", --  598 - 0x256  :   48 - 0x30
    "00000000", --  599 - 0x257  :    0 - 0x0
    "01000100", --  600 - 0x258  :   68 - 0x44 -- Sprite 0x4b
    "01000100", --  601 - 0x259  :   68 - 0x44
    "01001000", --  602 - 0x25a  :   72 - 0x48
    "01110000", --  603 - 0x25b  :  112 - 0x70
    "01001000", --  604 - 0x25c  :   72 - 0x48
    "00100100", --  605 - 0x25d  :   36 - 0x24
    "00100010", --  606 - 0x25e  :   34 - 0x22
    "00000000", --  607 - 0x25f  :    0 - 0x0
    "00010000", --  608 - 0x260  :   16 - 0x10 -- Sprite 0x4c
    "00100000", --  609 - 0x261  :   32 - 0x20
    "00100000", --  610 - 0x262  :   32 - 0x20
    "00100000", --  611 - 0x263  :   32 - 0x20
    "01000000", --  612 - 0x264  :   64 - 0x40
    "01000000", --  613 - 0x265  :   64 - 0x40
    "01000110", --  614 - 0x266  :   70 - 0x46
    "00111000", --  615 - 0x267  :   56 - 0x38
    "00100100", --  616 - 0x268  :   36 - 0x24 -- Sprite 0x4d
    "01011010", --  617 - 0x269  :   90 - 0x5a
    "01011010", --  618 - 0x26a  :   90 - 0x5a
    "01011010", --  619 - 0x26b  :   90 - 0x5a
    "01000010", --  620 - 0x26c  :   66 - 0x42
    "01000010", --  621 - 0x26d  :   66 - 0x42
    "00100010", --  622 - 0x26e  :   34 - 0x22
    "00000000", --  623 - 0x26f  :    0 - 0x0
    "00100100", --  624 - 0x270  :   36 - 0x24 -- Sprite 0x4e
    "01010010", --  625 - 0x271  :   82 - 0x52
    "01010010", --  626 - 0x272  :   82 - 0x52
    "01010010", --  627 - 0x273  :   82 - 0x52
    "01010010", --  628 - 0x274  :   82 - 0x52
    "01010010", --  629 - 0x275  :   82 - 0x52
    "01001100", --  630 - 0x276  :   76 - 0x4c
    "00000000", --  631 - 0x277  :    0 - 0x0
    "00111000", --  632 - 0x278  :   56 - 0x38 -- Sprite 0x4f
    "01000100", --  633 - 0x279  :   68 - 0x44
    "10000010", --  634 - 0x27a  :  130 - 0x82
    "10000010", --  635 - 0x27b  :  130 - 0x82
    "10000010", --  636 - 0x27c  :  130 - 0x82
    "01000100", --  637 - 0x27d  :   68 - 0x44
    "00111000", --  638 - 0x27e  :   56 - 0x38
    "00000000", --  639 - 0x27f  :    0 - 0x0
    "01111111", --  640 - 0x280  :  127 - 0x7f -- Sprite 0x50
    "11000000", --  641 - 0x281  :  192 - 0xc0
    "10000000", --  642 - 0x282  :  128 - 0x80
    "10000000", --  643 - 0x283  :  128 - 0x80
    "10000000", --  644 - 0x284  :  128 - 0x80
    "11000011", --  645 - 0x285  :  195 - 0xc3
    "11111111", --  646 - 0x286  :  255 - 0xff
    "11111111", --  647 - 0x287  :  255 - 0xff
    "11111110", --  648 - 0x288  :  254 - 0xfe -- Sprite 0x51
    "00000011", --  649 - 0x289  :    3 - 0x3
    "00000001", --  650 - 0x28a  :    1 - 0x1
    "00000001", --  651 - 0x28b  :    1 - 0x1
    "00000001", --  652 - 0x28c  :    1 - 0x1
    "11000011", --  653 - 0x28d  :  195 - 0xc3
    "11111111", --  654 - 0x28e  :  255 - 0xff
    "11111111", --  655 - 0x28f  :  255 - 0xff
    "00000000", --  656 - 0x290  :    0 - 0x0 -- Sprite 0x52
    "00000111", --  657 - 0x291  :    7 - 0x7
    "00001100", --  658 - 0x292  :   12 - 0xc
    "00011000", --  659 - 0x293  :   24 - 0x18
    "00110000", --  660 - 0x294  :   48 - 0x30
    "01100000", --  661 - 0x295  :   96 - 0x60
    "01000000", --  662 - 0x296  :   64 - 0x40
    "01001111", --  663 - 0x297  :   79 - 0x4f
    "00000000", --  664 - 0x298  :    0 - 0x0 -- Sprite 0x53
    "11110000", --  665 - 0x299  :  240 - 0xf0
    "01010000", --  666 - 0x29a  :   80 - 0x50
    "01001000", --  667 - 0x29b  :   72 - 0x48
    "01001100", --  668 - 0x29c  :   76 - 0x4c
    "01000100", --  669 - 0x29d  :   68 - 0x44
    "10000010", --  670 - 0x29e  :  130 - 0x82
    "10000011", --  671 - 0x29f  :  131 - 0x83
    "01111111", --  672 - 0x2a0  :  127 - 0x7f -- Sprite 0x54
    "11011110", --  673 - 0x2a1  :  222 - 0xde
    "10001110", --  674 - 0x2a2  :  142 - 0x8e
    "11000101", --  675 - 0x2a3  :  197 - 0xc5
    "10010010", --  676 - 0x2a4  :  146 - 0x92
    "11000111", --  677 - 0x2a5  :  199 - 0xc7
    "11100010", --  678 - 0x2a6  :  226 - 0xe2
    "11010000", --  679 - 0x2a7  :  208 - 0xd0
    "11111111", --  680 - 0x2a8  :  255 - 0xff -- Sprite 0x55
    "11011110", --  681 - 0x2a9  :  222 - 0xde
    "10001110", --  682 - 0x2aa  :  142 - 0x8e
    "11000101", --  683 - 0x2ab  :  197 - 0xc5
    "10010010", --  684 - 0x2ac  :  146 - 0x92
    "01000111", --  685 - 0x2ad  :   71 - 0x47
    "11100010", --  686 - 0x2ae  :  226 - 0xe2
    "01010000", --  687 - 0x2af  :   80 - 0x50
    "11111110", --  688 - 0x2b0  :  254 - 0xfe -- Sprite 0x56
    "11011111", --  689 - 0x2b1  :  223 - 0xdf
    "10001111", --  690 - 0x2b2  :  143 - 0x8f
    "11000101", --  691 - 0x2b3  :  197 - 0xc5
    "10010011", --  692 - 0x2b4  :  147 - 0x93
    "01000111", --  693 - 0x2b5  :   71 - 0x47
    "11100011", --  694 - 0x2b6  :  227 - 0xe3
    "01010001", --  695 - 0x2b7  :   81 - 0x51
    "01111111", --  696 - 0x2b8  :  127 - 0x7f -- Sprite 0x57
    "10000000", --  697 - 0x2b9  :  128 - 0x80
    "10110011", --  698 - 0x2ba  :  179 - 0xb3
    "01001100", --  699 - 0x2bb  :   76 - 0x4c
    "00111111", --  700 - 0x2bc  :   63 - 0x3f
    "00000011", --  701 - 0x2bd  :    3 - 0x3
    "00000000", --  702 - 0x2be  :    0 - 0x0
    "00000000", --  703 - 0x2bf  :    0 - 0x0
    "11111111", --  704 - 0x2c0  :  255 - 0xff -- Sprite 0x58
    "00000000", --  705 - 0x2c1  :    0 - 0x0
    "00110011", --  706 - 0x2c2  :   51 - 0x33
    "11001100", --  707 - 0x2c3  :  204 - 0xcc
    "00110011", --  708 - 0x2c4  :   51 - 0x33
    "11111111", --  709 - 0x2c5  :  255 - 0xff
    "00000000", --  710 - 0x2c6  :    0 - 0x0
    "00000000", --  711 - 0x2c7  :    0 - 0x0
    "11111110", --  712 - 0x2c8  :  254 - 0xfe -- Sprite 0x59
    "00000001", --  713 - 0x2c9  :    1 - 0x1
    "00110011", --  714 - 0x2ca  :   51 - 0x33
    "11001110", --  715 - 0x2cb  :  206 - 0xce
    "00111100", --  716 - 0x2cc  :   60 - 0x3c
    "11000000", --  717 - 0x2cd  :  192 - 0xc0
    "00000000", --  718 - 0x2ce  :    0 - 0x0
    "00000000", --  719 - 0x2cf  :    0 - 0x0
    "00000000", --  720 - 0x2d0  :    0 - 0x0 -- Sprite 0x5a
    "00000000", --  721 - 0x2d1  :    0 - 0x0
    "00000000", --  722 - 0x2d2  :    0 - 0x0
    "00000000", --  723 - 0x2d3  :    0 - 0x0
    "00000000", --  724 - 0x2d4  :    0 - 0x0
    "00000000", --  725 - 0x2d5  :    0 - 0x0
    "00000000", --  726 - 0x2d6  :    0 - 0x0
    "00000000", --  727 - 0x2d7  :    0 - 0x0
    "00000000", --  728 - 0x2d8  :    0 - 0x0 -- Sprite 0x5b
    "00000000", --  729 - 0x2d9  :    0 - 0x0
    "00000000", --  730 - 0x2da  :    0 - 0x0
    "00000001", --  731 - 0x2db  :    1 - 0x1
    "00000011", --  732 - 0x2dc  :    3 - 0x3
    "00000011", --  733 - 0x2dd  :    3 - 0x3
    "00000111", --  734 - 0x2de  :    7 - 0x7
    "00111111", --  735 - 0x2df  :   63 - 0x3f
    "00000000", --  736 - 0x2e0  :    0 - 0x0 -- Sprite 0x5c
    "00000001", --  737 - 0x2e1  :    1 - 0x1
    "01111111", --  738 - 0x2e2  :  127 - 0x7f
    "11111111", --  739 - 0x2e3  :  255 - 0xff
    "11111111", --  740 - 0x2e4  :  255 - 0xff
    "11111111", --  741 - 0x2e5  :  255 - 0xff
    "11111111", --  742 - 0x2e6  :  255 - 0xff
    "11111111", --  743 - 0x2e7  :  255 - 0xff
    "11111111", --  744 - 0x2e8  :  255 - 0xff -- Sprite 0x5d
    "11111111", --  745 - 0x2e9  :  255 - 0xff
    "11111111", --  746 - 0x2ea  :  255 - 0xff
    "11111111", --  747 - 0x2eb  :  255 - 0xff
    "11111111", --  748 - 0x2ec  :  255 - 0xff
    "11111111", --  749 - 0x2ed  :  255 - 0xff
    "11111111", --  750 - 0x2ee  :  255 - 0xff
    "11111111", --  751 - 0x2ef  :  255 - 0xff
    "00000000", --  752 - 0x2f0  :    0 - 0x0 -- Sprite 0x5e
    "10000000", --  753 - 0x2f1  :  128 - 0x80
    "11111110", --  754 - 0x2f2  :  254 - 0xfe
    "11111111", --  755 - 0x2f3  :  255 - 0xff
    "11111111", --  756 - 0x2f4  :  255 - 0xff
    "11111111", --  757 - 0x2f5  :  255 - 0xff
    "11111111", --  758 - 0x2f6  :  255 - 0xff
    "11111111", --  759 - 0x2f7  :  255 - 0xff
    "00000000", --  760 - 0x2f8  :    0 - 0x0 -- Sprite 0x5f
    "00000000", --  761 - 0x2f9  :    0 - 0x0
    "00000000", --  762 - 0x2fa  :    0 - 0x0
    "10000000", --  763 - 0x2fb  :  128 - 0x80
    "11000000", --  764 - 0x2fc  :  192 - 0xc0
    "11000000", --  765 - 0x2fd  :  192 - 0xc0
    "11100000", --  766 - 0x2fe  :  224 - 0xe0
    "11111000", --  767 - 0x2ff  :  248 - 0xf8
    "11111111", --  768 - 0x300  :  255 - 0xff -- Sprite 0x60
    "11111111", --  769 - 0x301  :  255 - 0xff
    "11111111", --  770 - 0x302  :  255 - 0xff
    "11111111", --  771 - 0x303  :  255 - 0xff
    "11111111", --  772 - 0x304  :  255 - 0xff
    "11111111", --  773 - 0x305  :  255 - 0xff
    "11111111", --  774 - 0x306  :  255 - 0xff
    "11111111", --  775 - 0x307  :  255 - 0xff
    "11111111", --  776 - 0x308  :  255 - 0xff -- Sprite 0x61
    "11111111", --  777 - 0x309  :  255 - 0xff
    "11111111", --  778 - 0x30a  :  255 - 0xff
    "11111111", --  779 - 0x30b  :  255 - 0xff
    "11111111", --  780 - 0x30c  :  255 - 0xff
    "11111111", --  781 - 0x30d  :  255 - 0xff
    "11111111", --  782 - 0x30e  :  255 - 0xff
    "11111111", --  783 - 0x30f  :  255 - 0xff
    "01111000", --  784 - 0x310  :  120 - 0x78 -- Sprite 0x62
    "01100000", --  785 - 0x311  :   96 - 0x60
    "01000000", --  786 - 0x312  :   64 - 0x40
    "01000000", --  787 - 0x313  :   64 - 0x40
    "01000000", --  788 - 0x314  :   64 - 0x40
    "01100000", --  789 - 0x315  :   96 - 0x60
    "00110000", --  790 - 0x316  :   48 - 0x30
    "00011111", --  791 - 0x317  :   31 - 0x1f
    "10000001", --  792 - 0x318  :  129 - 0x81 -- Sprite 0x63
    "10000011", --  793 - 0x319  :  131 - 0x83
    "11000001", --  794 - 0x31a  :  193 - 0xc1
    "01000011", --  795 - 0x31b  :   67 - 0x43
    "01000001", --  796 - 0x31c  :   65 - 0x41
    "01100011", --  797 - 0x31d  :   99 - 0x63
    "00100110", --  798 - 0x31e  :   38 - 0x26
    "11111000", --  799 - 0x31f  :  248 - 0xf8
    "10111001", --  800 - 0x320  :  185 - 0xb9 -- Sprite 0x64
    "10010100", --  801 - 0x321  :  148 - 0x94
    "10001110", --  802 - 0x322  :  142 - 0x8e
    "11000101", --  803 - 0x323  :  197 - 0xc5
    "10010010", --  804 - 0x324  :  146 - 0x92
    "11000111", --  805 - 0x325  :  199 - 0xc7
    "11100010", --  806 - 0x326  :  226 - 0xe2
    "11010000", --  807 - 0x327  :  208 - 0xd0
    "10111001", --  808 - 0x328  :  185 - 0xb9 -- Sprite 0x65
    "00010100", --  809 - 0x329  :   20 - 0x14
    "10001110", --  810 - 0x32a  :  142 - 0x8e
    "11000101", --  811 - 0x32b  :  197 - 0xc5
    "10010010", --  812 - 0x32c  :  146 - 0x92
    "01000111", --  813 - 0x32d  :   71 - 0x47
    "11100010", --  814 - 0x32e  :  226 - 0xe2
    "01010000", --  815 - 0x32f  :   80 - 0x50
    "10111001", --  816 - 0x330  :  185 - 0xb9 -- Sprite 0x66
    "00010101", --  817 - 0x331  :   21 - 0x15
    "10001111", --  818 - 0x332  :  143 - 0x8f
    "11000101", --  819 - 0x333  :  197 - 0xc5
    "10010011", --  820 - 0x334  :  147 - 0x93
    "01000111", --  821 - 0x335  :   71 - 0x47
    "11100011", --  822 - 0x336  :  227 - 0xe3
    "01010001", --  823 - 0x337  :   81 - 0x51
    "01111111", --  824 - 0x338  :  127 - 0x7f -- Sprite 0x67
    "10000000", --  825 - 0x339  :  128 - 0x80
    "11001100", --  826 - 0x33a  :  204 - 0xcc
    "01111111", --  827 - 0x33b  :  127 - 0x7f
    "00111111", --  828 - 0x33c  :   63 - 0x3f
    "00000011", --  829 - 0x33d  :    3 - 0x3
    "00000000", --  830 - 0x33e  :    0 - 0x0
    "00000000", --  831 - 0x33f  :    0 - 0x0
    "11111111", --  832 - 0x340  :  255 - 0xff -- Sprite 0x68
    "00000000", --  833 - 0x341  :    0 - 0x0
    "11001100", --  834 - 0x342  :  204 - 0xcc
    "00110011", --  835 - 0x343  :   51 - 0x33
    "11111111", --  836 - 0x344  :  255 - 0xff
    "11111111", --  837 - 0x345  :  255 - 0xff
    "00000000", --  838 - 0x346  :    0 - 0x0
    "00000000", --  839 - 0x347  :    0 - 0x0
    "11111110", --  840 - 0x348  :  254 - 0xfe -- Sprite 0x69
    "00000001", --  841 - 0x349  :    1 - 0x1
    "11001101", --  842 - 0x34a  :  205 - 0xcd
    "00111110", --  843 - 0x34b  :   62 - 0x3e
    "11111100", --  844 - 0x34c  :  252 - 0xfc
    "11000000", --  845 - 0x34d  :  192 - 0xc0
    "00000000", --  846 - 0x34e  :    0 - 0x0
    "00000000", --  847 - 0x34f  :    0 - 0x0
    "00000000", --  848 - 0x350  :    0 - 0x0 -- Sprite 0x6a
    "00000000", --  849 - 0x351  :    0 - 0x0
    "00000000", --  850 - 0x352  :    0 - 0x0
    "00000000", --  851 - 0x353  :    0 - 0x0
    "00000000", --  852 - 0x354  :    0 - 0x0
    "00000000", --  853 - 0x355  :    0 - 0x0
    "00000000", --  854 - 0x356  :    0 - 0x0
    "00000000", --  855 - 0x357  :    0 - 0x0
    "01111111", --  856 - 0x358  :  127 - 0x7f -- Sprite 0x6b
    "11111111", --  857 - 0x359  :  255 - 0xff
    "11111111", --  858 - 0x35a  :  255 - 0xff
    "11111111", --  859 - 0x35b  :  255 - 0xff
    "01111111", --  860 - 0x35c  :  127 - 0x7f
    "00110000", --  861 - 0x35d  :   48 - 0x30
    "00001111", --  862 - 0x35e  :   15 - 0xf
    "00000000", --  863 - 0x35f  :    0 - 0x0
    "11111111", --  864 - 0x360  :  255 - 0xff -- Sprite 0x6c
    "11111111", --  865 - 0x361  :  255 - 0xff
    "11111111", --  866 - 0x362  :  255 - 0xff
    "11111111", --  867 - 0x363  :  255 - 0xff
    "11111111", --  868 - 0x364  :  255 - 0xff
    "11111110", --  869 - 0x365  :  254 - 0xfe
    "00000001", --  870 - 0x366  :    1 - 0x1
    "11111110", --  871 - 0x367  :  254 - 0xfe
    "00000000", --  872 - 0x368  :    0 - 0x0 -- Sprite 0x6d
    "00000000", --  873 - 0x369  :    0 - 0x0
    "00000000", --  874 - 0x36a  :    0 - 0x0
    "00000000", --  875 - 0x36b  :    0 - 0x0
    "00000000", --  876 - 0x36c  :    0 - 0x0
    "00000000", --  877 - 0x36d  :    0 - 0x0
    "00000000", --  878 - 0x36e  :    0 - 0x0
    "00000000", --  879 - 0x36f  :    0 - 0x0
    "00000000", --  880 - 0x370  :    0 - 0x0 -- Sprite 0x6e
    "00000000", --  881 - 0x371  :    0 - 0x0
    "00000000", --  882 - 0x372  :    0 - 0x0
    "00000000", --  883 - 0x373  :    0 - 0x0
    "00000000", --  884 - 0x374  :    0 - 0x0
    "00000000", --  885 - 0x375  :    0 - 0x0
    "00000000", --  886 - 0x376  :    0 - 0x0
    "00000000", --  887 - 0x377  :    0 - 0x0
    "11111100", --  888 - 0x378  :  252 - 0xfc -- Sprite 0x6f
    "11111110", --  889 - 0x379  :  254 - 0xfe
    "11111111", --  890 - 0x37a  :  255 - 0xff
    "11111111", --  891 - 0x37b  :  255 - 0xff
    "11110010", --  892 - 0x37c  :  242 - 0xf2
    "00001100", --  893 - 0x37d  :   12 - 0xc
    "11110000", --  894 - 0x37e  :  240 - 0xf0
    "00000000", --  895 - 0x37f  :    0 - 0x0
    "01111111", --  896 - 0x380  :  127 - 0x7f -- Sprite 0x70
    "11000000", --  897 - 0x381  :  192 - 0xc0
    "10000000", --  898 - 0x382  :  128 - 0x80
    "10000000", --  899 - 0x383  :  128 - 0x80
    "11100011", --  900 - 0x384  :  227 - 0xe3
    "11111111", --  901 - 0x385  :  255 - 0xff
    "11111111", --  902 - 0x386  :  255 - 0xff
    "11111111", --  903 - 0x387  :  255 - 0xff
    "11111111", --  904 - 0x388  :  255 - 0xff -- Sprite 0x71
    "00000000", --  905 - 0x389  :    0 - 0x0
    "00000000", --  906 - 0x38a  :    0 - 0x0
    "00000000", --  907 - 0x38b  :    0 - 0x0
    "00000000", --  908 - 0x38c  :    0 - 0x0
    "11000011", --  909 - 0x38d  :  195 - 0xc3
    "11111111", --  910 - 0x38e  :  255 - 0xff
    "11111111", --  911 - 0x38f  :  255 - 0xff
    "11111110", --  912 - 0x390  :  254 - 0xfe -- Sprite 0x72
    "00000011", --  913 - 0x391  :    3 - 0x3
    "00000001", --  914 - 0x392  :    1 - 0x1
    "00000001", --  915 - 0x393  :    1 - 0x1
    "11000111", --  916 - 0x394  :  199 - 0xc7
    "11111111", --  917 - 0x395  :  255 - 0xff
    "11111111", --  918 - 0x396  :  255 - 0xff
    "11111111", --  919 - 0x397  :  255 - 0xff
    "11111111", --  920 - 0x398  :  255 - 0xff -- Sprite 0x73
    "11111111", --  921 - 0x399  :  255 - 0xff
    "11111111", --  922 - 0x39a  :  255 - 0xff
    "11111111", --  923 - 0x39b  :  255 - 0xff
    "11111111", --  924 - 0x39c  :  255 - 0xff
    "11111111", --  925 - 0x39d  :  255 - 0xff
    "11111111", --  926 - 0x39e  :  255 - 0xff
    "11111111", --  927 - 0x39f  :  255 - 0xff
    "10111001", --  928 - 0x3a0  :  185 - 0xb9 -- Sprite 0x74
    "10010100", --  929 - 0x3a1  :  148 - 0x94
    "10001110", --  930 - 0x3a2  :  142 - 0x8e
    "11000101", --  931 - 0x3a3  :  197 - 0xc5
    "10010010", --  932 - 0x3a4  :  146 - 0x92
    "11000111", --  933 - 0x3a5  :  199 - 0xc7
    "11100010", --  934 - 0x3a6  :  226 - 0xe2
    "01111111", --  935 - 0x3a7  :  127 - 0x7f
    "10111001", --  936 - 0x3a8  :  185 - 0xb9 -- Sprite 0x75
    "00010100", --  937 - 0x3a9  :   20 - 0x14
    "10001110", --  938 - 0x3aa  :  142 - 0x8e
    "11000101", --  939 - 0x3ab  :  197 - 0xc5
    "10010010", --  940 - 0x3ac  :  146 - 0x92
    "01000111", --  941 - 0x3ad  :   71 - 0x47
    "11100010", --  942 - 0x3ae  :  226 - 0xe2
    "11111111", --  943 - 0x3af  :  255 - 0xff
    "10111001", --  944 - 0x3b0  :  185 - 0xb9 -- Sprite 0x76
    "00010101", --  945 - 0x3b1  :   21 - 0x15
    "10001111", --  946 - 0x3b2  :  143 - 0x8f
    "11000101", --  947 - 0x3b3  :  197 - 0xc5
    "10010011", --  948 - 0x3b4  :  147 - 0x93
    "01000111", --  949 - 0x3b5  :   71 - 0x47
    "11100011", --  950 - 0x3b6  :  227 - 0xe3
    "11111110", --  951 - 0x3b7  :  254 - 0xfe
    "11111111", --  952 - 0x3b8  :  255 - 0xff -- Sprite 0x77
    "11111111", --  953 - 0x3b9  :  255 - 0xff
    "11111111", --  954 - 0x3ba  :  255 - 0xff
    "11111111", --  955 - 0x3bb  :  255 - 0xff
    "11111111", --  956 - 0x3bc  :  255 - 0xff
    "11111111", --  957 - 0x3bd  :  255 - 0xff
    "11111111", --  958 - 0x3be  :  255 - 0xff
    "11111111", --  959 - 0x3bf  :  255 - 0xff
    "00000000", --  960 - 0x3c0  :    0 - 0x0 -- Sprite 0x78
    "00000000", --  961 - 0x3c1  :    0 - 0x0
    "00000000", --  962 - 0x3c2  :    0 - 0x0
    "00000000", --  963 - 0x3c3  :    0 - 0x0
    "00000000", --  964 - 0x3c4  :    0 - 0x0
    "00000000", --  965 - 0x3c5  :    0 - 0x0
    "00000000", --  966 - 0x3c6  :    0 - 0x0
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "00000000", --  968 - 0x3c8  :    0 - 0x0 -- Sprite 0x79
    "00000000", --  969 - 0x3c9  :    0 - 0x0
    "00000000", --  970 - 0x3ca  :    0 - 0x0
    "00000000", --  971 - 0x3cb  :    0 - 0x0
    "00000000", --  972 - 0x3cc  :    0 - 0x0
    "00000000", --  973 - 0x3cd  :    0 - 0x0
    "00000000", --  974 - 0x3ce  :    0 - 0x0
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "00000000", --  976 - 0x3d0  :    0 - 0x0 -- Sprite 0x7a
    "00000000", --  977 - 0x3d1  :    0 - 0x0
    "00000000", --  978 - 0x3d2  :    0 - 0x0
    "00000000", --  979 - 0x3d3  :    0 - 0x0
    "00000000", --  980 - 0x3d4  :    0 - 0x0
    "00000000", --  981 - 0x3d5  :    0 - 0x0
    "00000000", --  982 - 0x3d6  :    0 - 0x0
    "00000000", --  983 - 0x3d7  :    0 - 0x0
    "00000000", --  984 - 0x3d8  :    0 - 0x0 -- Sprite 0x7b
    "00000000", --  985 - 0x3d9  :    0 - 0x0
    "00000000", --  986 - 0x3da  :    0 - 0x0
    "00000000", --  987 - 0x3db  :    0 - 0x0
    "00000000", --  988 - 0x3dc  :    0 - 0x0
    "00000000", --  989 - 0x3dd  :    0 - 0x0
    "00000000", --  990 - 0x3de  :    0 - 0x0
    "00000000", --  991 - 0x3df  :    0 - 0x0
    "00100010", --  992 - 0x3e0  :   34 - 0x22 -- Sprite 0x7c
    "01010101", --  993 - 0x3e1  :   85 - 0x55
    "10101010", --  994 - 0x3e2  :  170 - 0xaa
    "00000101", --  995 - 0x3e3  :    5 - 0x5
    "00000100", --  996 - 0x3e4  :    4 - 0x4
    "00001010", --  997 - 0x3e5  :   10 - 0xa
    "01010000", --  998 - 0x3e6  :   80 - 0x50
    "00000010", --  999 - 0x3e7  :    2 - 0x2
    "01110011", -- 1000 - 0x3e8  :  115 - 0x73 -- Sprite 0x7d
    "11111111", -- 1001 - 0x3e9  :  255 - 0xff
    "11111111", -- 1002 - 0x3ea  :  255 - 0xff
    "10111101", -- 1003 - 0x3eb  :  189 - 0xbd
    "01101110", -- 1004 - 0x3ec  :  110 - 0x6e
    "00001010", -- 1005 - 0x3ed  :   10 - 0xa
    "01010000", -- 1006 - 0x3ee  :   80 - 0x50
    "00000010", -- 1007 - 0x3ef  :    2 - 0x2
    "00100000", -- 1008 - 0x3f0  :   32 - 0x20 -- Sprite 0x7e
    "01010000", -- 1009 - 0x3f1  :   80 - 0x50
    "10000100", -- 1010 - 0x3f2  :  132 - 0x84
    "00000000", -- 1011 - 0x3f3  :    0 - 0x0
    "00100100", -- 1012 - 0x3f4  :   36 - 0x24
    "01011010", -- 1013 - 0x3f5  :   90 - 0x5a
    "00010000", -- 1014 - 0x3f6  :   16 - 0x10
    "00000000", -- 1015 - 0x3f7  :    0 - 0x0
    "11111111", -- 1016 - 0x3f8  :  255 - 0xff -- Sprite 0x7f
    "01010000", -- 1017 - 0x3f9  :   80 - 0x50
    "10000100", -- 1018 - 0x3fa  :  132 - 0x84
    "00000000", -- 1019 - 0x3fb  :    0 - 0x0
    "00100100", -- 1020 - 0x3fc  :   36 - 0x24
    "01011010", -- 1021 - 0x3fd  :   90 - 0x5a
    "00010000", -- 1022 - 0x3fe  :   16 - 0x10
    "00000000", -- 1023 - 0x3ff  :    0 - 0x0
    "11111111", -- 1024 - 0x400  :  255 - 0xff -- Sprite 0x80
    "10000000", -- 1025 - 0x401  :  128 - 0x80
    "11001111", -- 1026 - 0x402  :  207 - 0xcf
    "01001000", -- 1027 - 0x403  :   72 - 0x48
    "11001111", -- 1028 - 0x404  :  207 - 0xcf
    "10000000", -- 1029 - 0x405  :  128 - 0x80
    "11001111", -- 1030 - 0x406  :  207 - 0xcf
    "01001000", -- 1031 - 0x407  :   72 - 0x48
    "11111111", -- 1032 - 0x408  :  255 - 0xff -- Sprite 0x81
    "10000000", -- 1033 - 0x409  :  128 - 0x80
    "11111111", -- 1034 - 0x40a  :  255 - 0xff
    "10000000", -- 1035 - 0x40b  :  128 - 0x80
    "10000000", -- 1036 - 0x40c  :  128 - 0x80
    "11011111", -- 1037 - 0x40d  :  223 - 0xdf
    "10110000", -- 1038 - 0x40e  :  176 - 0xb0
    "11000000", -- 1039 - 0x40f  :  192 - 0xc0
    "11111111", -- 1040 - 0x410  :  255 - 0xff -- Sprite 0x82
    "00000001", -- 1041 - 0x411  :    1 - 0x1
    "11110011", -- 1042 - 0x412  :  243 - 0xf3
    "00010010", -- 1043 - 0x413  :   18 - 0x12
    "11110011", -- 1044 - 0x414  :  243 - 0xf3
    "00000001", -- 1045 - 0x415  :    1 - 0x1
    "11110011", -- 1046 - 0x416  :  243 - 0xf3
    "00010010", -- 1047 - 0x417  :   18 - 0x12
    "11111111", -- 1048 - 0x418  :  255 - 0xff -- Sprite 0x83
    "00000000", -- 1049 - 0x419  :    0 - 0x0
    "11111111", -- 1050 - 0x41a  :  255 - 0xff
    "00000000", -- 1051 - 0x41b  :    0 - 0x0
    "00000000", -- 1052 - 0x41c  :    0 - 0x0
    "11111111", -- 1053 - 0x41d  :  255 - 0xff
    "00000000", -- 1054 - 0x41e  :    0 - 0x0
    "00000000", -- 1055 - 0x41f  :    0 - 0x0
    "11111111", -- 1056 - 0x420  :  255 - 0xff -- Sprite 0x84
    "10000010", -- 1057 - 0x421  :  130 - 0x82
    "00010000", -- 1058 - 0x422  :   16 - 0x10
    "00000000", -- 1059 - 0x423  :    0 - 0x0
    "00000000", -- 1060 - 0x424  :    0 - 0x0
    "00010000", -- 1061 - 0x425  :   16 - 0x10
    "01000100", -- 1062 - 0x426  :   68 - 0x44
    "11111111", -- 1063 - 0x427  :  255 - 0xff
    "11111111", -- 1064 - 0x428  :  255 - 0xff -- Sprite 0x85
    "00000001", -- 1065 - 0x429  :    1 - 0x1
    "11111111", -- 1066 - 0x42a  :  255 - 0xff
    "00000001", -- 1067 - 0x42b  :    1 - 0x1
    "00000001", -- 1068 - 0x42c  :    1 - 0x1
    "11110011", -- 1069 - 0x42d  :  243 - 0xf3
    "00001101", -- 1070 - 0x42e  :   13 - 0xd
    "00000011", -- 1071 - 0x42f  :    3 - 0x3
    "00000000", -- 1072 - 0x430  :    0 - 0x0 -- Sprite 0x86
    "00000000", -- 1073 - 0x431  :    0 - 0x0
    "00000000", -- 1074 - 0x432  :    0 - 0x0
    "00000000", -- 1075 - 0x433  :    0 - 0x0
    "00000000", -- 1076 - 0x434  :    0 - 0x0
    "00000000", -- 1077 - 0x435  :    0 - 0x0
    "00000000", -- 1078 - 0x436  :    0 - 0x0
    "00000000", -- 1079 - 0x437  :    0 - 0x0
    "00000000", -- 1080 - 0x438  :    0 - 0x0 -- Sprite 0x87
    "00000000", -- 1081 - 0x439  :    0 - 0x0
    "00000000", -- 1082 - 0x43a  :    0 - 0x0
    "00000000", -- 1083 - 0x43b  :    0 - 0x0
    "00000000", -- 1084 - 0x43c  :    0 - 0x0
    "00000000", -- 1085 - 0x43d  :    0 - 0x0
    "00000000", -- 1086 - 0x43e  :    0 - 0x0
    "00000000", -- 1087 - 0x43f  :    0 - 0x0
    "00000111", -- 1088 - 0x440  :    7 - 0x7 -- Sprite 0x88
    "00011110", -- 1089 - 0x441  :   30 - 0x1e
    "00101111", -- 1090 - 0x442  :   47 - 0x2f
    "01010011", -- 1091 - 0x443  :   83 - 0x53
    "01101110", -- 1092 - 0x444  :  110 - 0x6e
    "11011011", -- 1093 - 0x445  :  219 - 0xdb
    "11111010", -- 1094 - 0x446  :  250 - 0xfa
    "11010101", -- 1095 - 0x447  :  213 - 0xd5
    "10111011", -- 1096 - 0x448  :  187 - 0xbb -- Sprite 0x89
    "11110010", -- 1097 - 0x449  :  242 - 0xf2
    "11011101", -- 1098 - 0x44a  :  221 - 0xdd
    "01001111", -- 1099 - 0x44b  :   79 - 0x4f
    "01111011", -- 1100 - 0x44c  :  123 - 0x7b
    "00110010", -- 1101 - 0x44d  :   50 - 0x32
    "00011111", -- 1102 - 0x44e  :   31 - 0x1f
    "00000111", -- 1103 - 0x44f  :    7 - 0x7
    "11100000", -- 1104 - 0x450  :  224 - 0xe0 -- Sprite 0x8a
    "11011000", -- 1105 - 0x451  :  216 - 0xd8
    "01010100", -- 1106 - 0x452  :   84 - 0x54
    "11101010", -- 1107 - 0x453  :  234 - 0xea
    "10111010", -- 1108 - 0x454  :  186 - 0xba
    "10010011", -- 1109 - 0x455  :  147 - 0x93
    "11011111", -- 1110 - 0x456  :  223 - 0xdf
    "10111101", -- 1111 - 0x457  :  189 - 0xbd
    "01101011", -- 1112 - 0x458  :  107 - 0x6b -- Sprite 0x8b
    "10011111", -- 1113 - 0x459  :  159 - 0x9f
    "01011101", -- 1114 - 0x45a  :   93 - 0x5d
    "10110110", -- 1115 - 0x45b  :  182 - 0xb6
    "11101010", -- 1116 - 0x45c  :  234 - 0xea
    "11001100", -- 1117 - 0x45d  :  204 - 0xcc
    "01111000", -- 1118 - 0x45e  :  120 - 0x78
    "11100000", -- 1119 - 0x45f  :  224 - 0xe0
    "00000111", -- 1120 - 0x460  :    7 - 0x7 -- Sprite 0x8c
    "00011000", -- 1121 - 0x461  :   24 - 0x18
    "00100011", -- 1122 - 0x462  :   35 - 0x23
    "01001100", -- 1123 - 0x463  :   76 - 0x4c
    "01110000", -- 1124 - 0x464  :  112 - 0x70
    "10100001", -- 1125 - 0x465  :  161 - 0xa1
    "10100110", -- 1126 - 0x466  :  166 - 0xa6
    "10101000", -- 1127 - 0x467  :  168 - 0xa8
    "10100101", -- 1128 - 0x468  :  165 - 0xa5 -- Sprite 0x8d
    "10100010", -- 1129 - 0x469  :  162 - 0xa2
    "10010000", -- 1130 - 0x46a  :  144 - 0x90
    "01001000", -- 1131 - 0x46b  :   72 - 0x48
    "01000111", -- 1132 - 0x46c  :   71 - 0x47
    "00100000", -- 1133 - 0x46d  :   32 - 0x20
    "00011001", -- 1134 - 0x46e  :   25 - 0x19
    "00000111", -- 1135 - 0x46f  :    7 - 0x7
    "11100000", -- 1136 - 0x470  :  224 - 0xe0 -- Sprite 0x8e
    "00011000", -- 1137 - 0x471  :   24 - 0x18
    "00000100", -- 1138 - 0x472  :    4 - 0x4
    "11000010", -- 1139 - 0x473  :  194 - 0xc2
    "00110010", -- 1140 - 0x474  :   50 - 0x32
    "00001001", -- 1141 - 0x475  :    9 - 0x9
    "11000101", -- 1142 - 0x476  :  197 - 0xc5
    "00100101", -- 1143 - 0x477  :   37 - 0x25
    "10100101", -- 1144 - 0x478  :  165 - 0xa5 -- Sprite 0x8f
    "01100101", -- 1145 - 0x479  :  101 - 0x65
    "01000101", -- 1146 - 0x47a  :   69 - 0x45
    "10001010", -- 1147 - 0x47b  :  138 - 0x8a
    "10010010", -- 1148 - 0x47c  :  146 - 0x92
    "00100100", -- 1149 - 0x47d  :   36 - 0x24
    "11011000", -- 1150 - 0x47e  :  216 - 0xd8
    "11100000", -- 1151 - 0x47f  :  224 - 0xe0
    "00000000", -- 1152 - 0x480  :    0 - 0x0 -- Sprite 0x90
    "00000000", -- 1153 - 0x481  :    0 - 0x0
    "00100000", -- 1154 - 0x482  :   32 - 0x20
    "00110000", -- 1155 - 0x483  :   48 - 0x30
    "00101100", -- 1156 - 0x484  :   44 - 0x2c
    "00100010", -- 1157 - 0x485  :   34 - 0x22
    "00010001", -- 1158 - 0x486  :   17 - 0x11
    "00001000", -- 1159 - 0x487  :    8 - 0x8
    "00000100", -- 1160 - 0x488  :    4 - 0x4 -- Sprite 0x91
    "11110010", -- 1161 - 0x489  :  242 - 0xf2
    "11001111", -- 1162 - 0x48a  :  207 - 0xcf
    "00110000", -- 1163 - 0x48b  :   48 - 0x30
    "00001100", -- 1164 - 0x48c  :   12 - 0xc
    "11111111", -- 1165 - 0x48d  :  255 - 0xff
    "10000000", -- 1166 - 0x48e  :  128 - 0x80
    "11111111", -- 1167 - 0x48f  :  255 - 0xff
    "01000010", -- 1168 - 0x490  :   66 - 0x42 -- Sprite 0x92
    "10100101", -- 1169 - 0x491  :  165 - 0xa5
    "10100101", -- 1170 - 0x492  :  165 - 0xa5
    "10011001", -- 1171 - 0x493  :  153 - 0x99
    "10011001", -- 1172 - 0x494  :  153 - 0x99
    "10011001", -- 1173 - 0x495  :  153 - 0x99
    "00000001", -- 1174 - 0x496  :    1 - 0x1
    "00000000", -- 1175 - 0x497  :    0 - 0x0
    "11111111", -- 1176 - 0x498  :  255 - 0xff -- Sprite 0x93
    "11111111", -- 1177 - 0x499  :  255 - 0xff
    "11111111", -- 1178 - 0x49a  :  255 - 0xff
    "10000001", -- 1179 - 0x49b  :  129 - 0x81
    "11111111", -- 1180 - 0x49c  :  255 - 0xff
    "11111111", -- 1181 - 0x49d  :  255 - 0xff
    "11111111", -- 1182 - 0x49e  :  255 - 0xff
    "10000001", -- 1183 - 0x49f  :  129 - 0x81
    "00000000", -- 1184 - 0x4a0  :    0 - 0x0 -- Sprite 0x94
    "00000000", -- 1185 - 0x4a1  :    0 - 0x0
    "00000100", -- 1186 - 0x4a2  :    4 - 0x4
    "00001100", -- 1187 - 0x4a3  :   12 - 0xc
    "00110100", -- 1188 - 0x4a4  :   52 - 0x34
    "01000100", -- 1189 - 0x4a5  :   68 - 0x44
    "10001000", -- 1190 - 0x4a6  :  136 - 0x88
    "00010000", -- 1191 - 0x4a7  :   16 - 0x10
    "00100000", -- 1192 - 0x4a8  :   32 - 0x20 -- Sprite 0x95
    "01001111", -- 1193 - 0x4a9  :   79 - 0x4f
    "11110011", -- 1194 - 0x4aa  :  243 - 0xf3
    "00001100", -- 1195 - 0x4ab  :   12 - 0xc
    "00110000", -- 1196 - 0x4ac  :   48 - 0x30
    "11111111", -- 1197 - 0x4ad  :  255 - 0xff
    "00000001", -- 1198 - 0x4ae  :    1 - 0x1
    "11111111", -- 1199 - 0x4af  :  255 - 0xff
    "01111111", -- 1200 - 0x4b0  :  127 - 0x7f -- Sprite 0x96
    "11111111", -- 1201 - 0x4b1  :  255 - 0xff
    "11111111", -- 1202 - 0x4b2  :  255 - 0xff
    "11111111", -- 1203 - 0x4b3  :  255 - 0xff
    "11111011", -- 1204 - 0x4b4  :  251 - 0xfb
    "11111111", -- 1205 - 0x4b5  :  255 - 0xff
    "11111111", -- 1206 - 0x4b6  :  255 - 0xff
    "11111111", -- 1207 - 0x4b7  :  255 - 0xff
    "11111111", -- 1208 - 0x4b8  :  255 - 0xff -- Sprite 0x97
    "11111111", -- 1209 - 0x4b9  :  255 - 0xff
    "11111111", -- 1210 - 0x4ba  :  255 - 0xff
    "11111111", -- 1211 - 0x4bb  :  255 - 0xff
    "11111111", -- 1212 - 0x4bc  :  255 - 0xff
    "11111111", -- 1213 - 0x4bd  :  255 - 0xff
    "11111110", -- 1214 - 0x4be  :  254 - 0xfe
    "11111111", -- 1215 - 0x4bf  :  255 - 0xff
    "11111111", -- 1216 - 0x4c0  :  255 - 0xff -- Sprite 0x98
    "10111111", -- 1217 - 0x4c1  :  191 - 0xbf
    "11111111", -- 1218 - 0x4c2  :  255 - 0xff
    "11111111", -- 1219 - 0x4c3  :  255 - 0xff
    "11111011", -- 1220 - 0x4c4  :  251 - 0xfb
    "11111111", -- 1221 - 0x4c5  :  255 - 0xff
    "11111111", -- 1222 - 0x4c6  :  255 - 0xff
    "11111111", -- 1223 - 0x4c7  :  255 - 0xff
    "11111111", -- 1224 - 0x4c8  :  255 - 0xff -- Sprite 0x99
    "11111111", -- 1225 - 0x4c9  :  255 - 0xff
    "11111111", -- 1226 - 0x4ca  :  255 - 0xff
    "11111111", -- 1227 - 0x4cb  :  255 - 0xff
    "11111111", -- 1228 - 0x4cc  :  255 - 0xff
    "11111111", -- 1229 - 0x4cd  :  255 - 0xff
    "11111110", -- 1230 - 0x4ce  :  254 - 0xfe
    "11111111", -- 1231 - 0x4cf  :  255 - 0xff
    "11111110", -- 1232 - 0x4d0  :  254 - 0xfe -- Sprite 0x9a
    "11111111", -- 1233 - 0x4d1  :  255 - 0xff
    "11111111", -- 1234 - 0x4d2  :  255 - 0xff
    "11111111", -- 1235 - 0x4d3  :  255 - 0xff
    "11111011", -- 1236 - 0x4d4  :  251 - 0xfb
    "11111111", -- 1237 - 0x4d5  :  255 - 0xff
    "11111111", -- 1238 - 0x4d6  :  255 - 0xff
    "11111111", -- 1239 - 0x4d7  :  255 - 0xff
    "11111111", -- 1240 - 0x4d8  :  255 - 0xff -- Sprite 0x9b
    "11111111", -- 1241 - 0x4d9  :  255 - 0xff
    "11111111", -- 1242 - 0x4da  :  255 - 0xff
    "11111111", -- 1243 - 0x4db  :  255 - 0xff
    "11111111", -- 1244 - 0x4dc  :  255 - 0xff
    "11111111", -- 1245 - 0x4dd  :  255 - 0xff
    "11111111", -- 1246 - 0x4de  :  255 - 0xff
    "11111111", -- 1247 - 0x4df  :  255 - 0xff
    "11111111", -- 1248 - 0x4e0  :  255 - 0xff -- Sprite 0x9c
    "11111111", -- 1249 - 0x4e1  :  255 - 0xff
    "10100000", -- 1250 - 0x4e2  :  160 - 0xa0
    "10010000", -- 1251 - 0x4e3  :  144 - 0x90
    "10001000", -- 1252 - 0x4e4  :  136 - 0x88
    "10000100", -- 1253 - 0x4e5  :  132 - 0x84
    "01101010", -- 1254 - 0x4e6  :  106 - 0x6a
    "00111111", -- 1255 - 0x4e7  :   63 - 0x3f
    "11111111", -- 1256 - 0x4e8  :  255 - 0xff -- Sprite 0x9d
    "11111111", -- 1257 - 0x4e9  :  255 - 0xff
    "00100001", -- 1258 - 0x4ea  :   33 - 0x21
    "00010001", -- 1259 - 0x4eb  :   17 - 0x11
    "00001001", -- 1260 - 0x4ec  :    9 - 0x9
    "00000101", -- 1261 - 0x4ed  :    5 - 0x5
    "10101010", -- 1262 - 0x4ee  :  170 - 0xaa
    "11111100", -- 1263 - 0x4ef  :  252 - 0xfc
    "11111111", -- 1264 - 0x4f0  :  255 - 0xff -- Sprite 0x9e
    "11111111", -- 1265 - 0x4f1  :  255 - 0xff
    "00100000", -- 1266 - 0x4f2  :   32 - 0x20
    "00010000", -- 1267 - 0x4f3  :   16 - 0x10
    "00001000", -- 1268 - 0x4f4  :    8 - 0x8
    "00000100", -- 1269 - 0x4f5  :    4 - 0x4
    "10101010", -- 1270 - 0x4f6  :  170 - 0xaa
    "11111111", -- 1271 - 0x4f7  :  255 - 0xff
    "00000000", -- 1272 - 0x4f8  :    0 - 0x0 -- Sprite 0x9f
    "00000000", -- 1273 - 0x4f9  :    0 - 0x0
    "00000000", -- 1274 - 0x4fa  :    0 - 0x0
    "00000000", -- 1275 - 0x4fb  :    0 - 0x0
    "00000000", -- 1276 - 0x4fc  :    0 - 0x0
    "00000000", -- 1277 - 0x4fd  :    0 - 0x0
    "00000000", -- 1278 - 0x4fe  :    0 - 0x0
    "00000000", -- 1279 - 0x4ff  :    0 - 0x0
    "11111111", -- 1280 - 0x500  :  255 - 0xff -- Sprite 0xa0
    "11010101", -- 1281 - 0x501  :  213 - 0xd5
    "11111111", -- 1282 - 0x502  :  255 - 0xff
    "00000010", -- 1283 - 0x503  :    2 - 0x2
    "00000010", -- 1284 - 0x504  :    2 - 0x2
    "00000010", -- 1285 - 0x505  :    2 - 0x2
    "00000010", -- 1286 - 0x506  :    2 - 0x2
    "00000010", -- 1287 - 0x507  :    2 - 0x2
    "00000010", -- 1288 - 0x508  :    2 - 0x2 -- Sprite 0xa1
    "00000010", -- 1289 - 0x509  :    2 - 0x2
    "00000010", -- 1290 - 0x50a  :    2 - 0x2
    "00000010", -- 1291 - 0x50b  :    2 - 0x2
    "00000010", -- 1292 - 0x50c  :    2 - 0x2
    "00000010", -- 1293 - 0x50d  :    2 - 0x2
    "00000010", -- 1294 - 0x50e  :    2 - 0x2
    "00000010", -- 1295 - 0x50f  :    2 - 0x2
    "11111111", -- 1296 - 0x510  :  255 - 0xff -- Sprite 0xa2
    "01010101", -- 1297 - 0x511  :   85 - 0x55
    "11111111", -- 1298 - 0x512  :  255 - 0xff
    "01000000", -- 1299 - 0x513  :   64 - 0x40
    "01000000", -- 1300 - 0x514  :   64 - 0x40
    "01000000", -- 1301 - 0x515  :   64 - 0x40
    "01000000", -- 1302 - 0x516  :   64 - 0x40
    "01000000", -- 1303 - 0x517  :   64 - 0x40
    "01000000", -- 1304 - 0x518  :   64 - 0x40 -- Sprite 0xa3
    "01000000", -- 1305 - 0x519  :   64 - 0x40
    "01000000", -- 1306 - 0x51a  :   64 - 0x40
    "01000000", -- 1307 - 0x51b  :   64 - 0x40
    "01000000", -- 1308 - 0x51c  :   64 - 0x40
    "01000000", -- 1309 - 0x51d  :   64 - 0x40
    "01000000", -- 1310 - 0x51e  :   64 - 0x40
    "01000000", -- 1311 - 0x51f  :   64 - 0x40
    "00110001", -- 1312 - 0x520  :   49 - 0x31 -- Sprite 0xa4
    "01001000", -- 1313 - 0x521  :   72 - 0x48
    "01000101", -- 1314 - 0x522  :   69 - 0x45
    "10000101", -- 1315 - 0x523  :  133 - 0x85
    "10000011", -- 1316 - 0x524  :  131 - 0x83
    "10000010", -- 1317 - 0x525  :  130 - 0x82
    "01100010", -- 1318 - 0x526  :   98 - 0x62
    "00010010", -- 1319 - 0x527  :   18 - 0x12
    "00110010", -- 1320 - 0x528  :   50 - 0x32 -- Sprite 0xa5
    "00100010", -- 1321 - 0x529  :   34 - 0x22
    "01000010", -- 1322 - 0x52a  :   66 - 0x42
    "01000000", -- 1323 - 0x52b  :   64 - 0x40
    "01000000", -- 1324 - 0x52c  :   64 - 0x40
    "00100000", -- 1325 - 0x52d  :   32 - 0x20
    "00011110", -- 1326 - 0x52e  :   30 - 0x1e
    "00000111", -- 1327 - 0x52f  :    7 - 0x7
    "10000000", -- 1328 - 0x530  :  128 - 0x80 -- Sprite 0xa6
    "11100000", -- 1329 - 0x531  :  224 - 0xe0
    "00111000", -- 1330 - 0x532  :   56 - 0x38
    "00100100", -- 1331 - 0x533  :   36 - 0x24
    "00000100", -- 1332 - 0x534  :    4 - 0x4
    "00001000", -- 1333 - 0x535  :    8 - 0x8
    "00110000", -- 1334 - 0x536  :   48 - 0x30
    "00100000", -- 1335 - 0x537  :   32 - 0x20
    "00110000", -- 1336 - 0x538  :   48 - 0x30 -- Sprite 0xa7
    "00001000", -- 1337 - 0x539  :    8 - 0x8
    "00001000", -- 1338 - 0x53a  :    8 - 0x8
    "00110000", -- 1339 - 0x53b  :   48 - 0x30
    "00100000", -- 1340 - 0x53c  :   32 - 0x20
    "00100000", -- 1341 - 0x53d  :   32 - 0x20
    "00110000", -- 1342 - 0x53e  :   48 - 0x30
    "11110000", -- 1343 - 0x53f  :  240 - 0xf0
    "11111111", -- 1344 - 0x540  :  255 - 0xff -- Sprite 0xa8
    "11010010", -- 1345 - 0x541  :  210 - 0xd2
    "11110100", -- 1346 - 0x542  :  244 - 0xf4
    "11011000", -- 1347 - 0x543  :  216 - 0xd8
    "11111000", -- 1348 - 0x544  :  248 - 0xf8
    "11010100", -- 1349 - 0x545  :  212 - 0xd4
    "11110010", -- 1350 - 0x546  :  242 - 0xf2
    "11010001", -- 1351 - 0x547  :  209 - 0xd1
    "11110001", -- 1352 - 0x548  :  241 - 0xf1 -- Sprite 0xa9
    "11010010", -- 1353 - 0x549  :  210 - 0xd2
    "11110100", -- 1354 - 0x54a  :  244 - 0xf4
    "11011000", -- 1355 - 0x54b  :  216 - 0xd8
    "11111000", -- 1356 - 0x54c  :  248 - 0xf8
    "11010100", -- 1357 - 0x54d  :  212 - 0xd4
    "11110010", -- 1358 - 0x54e  :  242 - 0xf2
    "11111111", -- 1359 - 0x54f  :  255 - 0xff
    "11111111", -- 1360 - 0x550  :  255 - 0xff -- Sprite 0xaa
    "01000010", -- 1361 - 0x551  :   66 - 0x42
    "00100100", -- 1362 - 0x552  :   36 - 0x24
    "00011000", -- 1363 - 0x553  :   24 - 0x18
    "00011000", -- 1364 - 0x554  :   24 - 0x18
    "00100100", -- 1365 - 0x555  :   36 - 0x24
    "01000010", -- 1366 - 0x556  :   66 - 0x42
    "10000001", -- 1367 - 0x557  :  129 - 0x81
    "10000001", -- 1368 - 0x558  :  129 - 0x81 -- Sprite 0xab
    "01000010", -- 1369 - 0x559  :   66 - 0x42
    "00100100", -- 1370 - 0x55a  :   36 - 0x24
    "00011000", -- 1371 - 0x55b  :   24 - 0x18
    "00011000", -- 1372 - 0x55c  :   24 - 0x18
    "00100100", -- 1373 - 0x55d  :   36 - 0x24
    "01000010", -- 1374 - 0x55e  :   66 - 0x42
    "11111111", -- 1375 - 0x55f  :  255 - 0xff
    "11111111", -- 1376 - 0x560  :  255 - 0xff -- Sprite 0xac
    "01001101", -- 1377 - 0x561  :   77 - 0x4d
    "00101111", -- 1378 - 0x562  :   47 - 0x2f
    "00011101", -- 1379 - 0x563  :   29 - 0x1d
    "00011111", -- 1380 - 0x564  :   31 - 0x1f
    "00101101", -- 1381 - 0x565  :   45 - 0x2d
    "01001111", -- 1382 - 0x566  :   79 - 0x4f
    "10001101", -- 1383 - 0x567  :  141 - 0x8d
    "10001111", -- 1384 - 0x568  :  143 - 0x8f -- Sprite 0xad
    "01001101", -- 1385 - 0x569  :   77 - 0x4d
    "00101111", -- 1386 - 0x56a  :   47 - 0x2f
    "00011101", -- 1387 - 0x56b  :   29 - 0x1d
    "00011111", -- 1388 - 0x56c  :   31 - 0x1f
    "00101101", -- 1389 - 0x56d  :   45 - 0x2d
    "01001111", -- 1390 - 0x56e  :   79 - 0x4f
    "11111111", -- 1391 - 0x56f  :  255 - 0xff
    "00000001", -- 1392 - 0x570  :    1 - 0x1 -- Sprite 0xae
    "00000011", -- 1393 - 0x571  :    3 - 0x3
    "00000110", -- 1394 - 0x572  :    6 - 0x6
    "00000111", -- 1395 - 0x573  :    7 - 0x7
    "00000111", -- 1396 - 0x574  :    7 - 0x7
    "00000111", -- 1397 - 0x575  :    7 - 0x7
    "00000110", -- 1398 - 0x576  :    6 - 0x6
    "00000111", -- 1399 - 0x577  :    7 - 0x7
    "00000110", -- 1400 - 0x578  :    6 - 0x6 -- Sprite 0xaf
    "00000110", -- 1401 - 0x579  :    6 - 0x6
    "00001110", -- 1402 - 0x57a  :   14 - 0xe
    "00001111", -- 1403 - 0x57b  :   15 - 0xf
    "00001110", -- 1404 - 0x57c  :   14 - 0xe
    "00011010", -- 1405 - 0x57d  :   26 - 0x1a
    "00011011", -- 1406 - 0x57e  :   27 - 0x1b
    "00001111", -- 1407 - 0x57f  :   15 - 0xf
    "00000000", -- 1408 - 0x580  :    0 - 0x0 -- Sprite 0xb0
    "11000000", -- 1409 - 0x581  :  192 - 0xc0
    "11110000", -- 1410 - 0x582  :  240 - 0xf0
    "10001000", -- 1411 - 0x583  :  136 - 0x88
    "00010100", -- 1412 - 0x584  :   20 - 0x14
    "01101000", -- 1413 - 0x585  :  104 - 0x68
    "10101000", -- 1414 - 0x586  :  168 - 0xa8
    "00101100", -- 1415 - 0x587  :   44 - 0x2c
    "00000100", -- 1416 - 0x588  :    4 - 0x4 -- Sprite 0xb1
    "00111000", -- 1417 - 0x589  :   56 - 0x38
    "00010000", -- 1418 - 0x58a  :   16 - 0x10
    "10100000", -- 1419 - 0x58b  :  160 - 0xa0
    "01100000", -- 1420 - 0x58c  :   96 - 0x60
    "00100000", -- 1421 - 0x58d  :   32 - 0x20
    "00010000", -- 1422 - 0x58e  :   16 - 0x10
    "10001000", -- 1423 - 0x58f  :  136 - 0x88
    "00001111", -- 1424 - 0x590  :   15 - 0xf -- Sprite 0xb2
    "00011011", -- 1425 - 0x591  :   27 - 0x1b
    "00011011", -- 1426 - 0x592  :   27 - 0x1b
    "00001110", -- 1427 - 0x593  :   14 - 0xe
    "00000110", -- 1428 - 0x594  :    6 - 0x6
    "00001100", -- 1429 - 0x595  :   12 - 0xc
    "00001100", -- 1430 - 0x596  :   12 - 0xc
    "00111111", -- 1431 - 0x597  :   63 - 0x3f
    "01111111", -- 1432 - 0x598  :  127 - 0x7f -- Sprite 0xb3
    "01100000", -- 1433 - 0x599  :   96 - 0x60
    "01100000", -- 1434 - 0x59a  :   96 - 0x60
    "01100000", -- 1435 - 0x59b  :   96 - 0x60
    "01100000", -- 1436 - 0x59c  :   96 - 0x60
    "01100000", -- 1437 - 0x59d  :   96 - 0x60
    "01101010", -- 1438 - 0x59e  :  106 - 0x6a
    "01111111", -- 1439 - 0x59f  :  127 - 0x7f
    "01001000", -- 1440 - 0x5a0  :   72 - 0x48 -- Sprite 0xb4
    "00110000", -- 1441 - 0x5a1  :   48 - 0x30
    "00010000", -- 1442 - 0x5a2  :   16 - 0x10
    "00010000", -- 1443 - 0x5a3  :   16 - 0x10
    "00001000", -- 1444 - 0x5a4  :    8 - 0x8
    "00001000", -- 1445 - 0x5a5  :    8 - 0x8
    "00001000", -- 1446 - 0x5a6  :    8 - 0x8
    "11111100", -- 1447 - 0x5a7  :  252 - 0xfc
    "11111110", -- 1448 - 0x5a8  :  254 - 0xfe -- Sprite 0xb5
    "00000110", -- 1449 - 0x5a9  :    6 - 0x6
    "00000010", -- 1450 - 0x5aa  :    2 - 0x2
    "00000110", -- 1451 - 0x5ab  :    6 - 0x6
    "00000010", -- 1452 - 0x5ac  :    2 - 0x2
    "00000110", -- 1453 - 0x5ad  :    6 - 0x6
    "10101010", -- 1454 - 0x5ae  :  170 - 0xaa
    "11111110", -- 1455 - 0x5af  :  254 - 0xfe
    "11111111", -- 1456 - 0x5b0  :  255 - 0xff -- Sprite 0xb6
    "10000000", -- 1457 - 0x5b1  :  128 - 0x80
    "10000000", -- 1458 - 0x5b2  :  128 - 0x80
    "10000000", -- 1459 - 0x5b3  :  128 - 0x80
    "10000000", -- 1460 - 0x5b4  :  128 - 0x80
    "10000000", -- 1461 - 0x5b5  :  128 - 0x80
    "10010101", -- 1462 - 0x5b6  :  149 - 0x95
    "11111111", -- 1463 - 0x5b7  :  255 - 0xff
    "11111111", -- 1464 - 0x5b8  :  255 - 0xff -- Sprite 0xb7
    "10000100", -- 1465 - 0x5b9  :  132 - 0x84
    "10001100", -- 1466 - 0x5ba  :  140 - 0x8c
    "10000100", -- 1467 - 0x5bb  :  132 - 0x84
    "10001100", -- 1468 - 0x5bc  :  140 - 0x8c
    "10000100", -- 1469 - 0x5bd  :  132 - 0x84
    "10101100", -- 1470 - 0x5be  :  172 - 0xac
    "11111111", -- 1471 - 0x5bf  :  255 - 0xff
    "11111111", -- 1472 - 0x5c0  :  255 - 0xff -- Sprite 0xb8
    "00100001", -- 1473 - 0x5c1  :   33 - 0x21
    "01100001", -- 1474 - 0x5c2  :   97 - 0x61
    "00100011", -- 1475 - 0x5c3  :   35 - 0x23
    "01100001", -- 1476 - 0x5c4  :   97 - 0x61
    "00100011", -- 1477 - 0x5c5  :   35 - 0x23
    "01100101", -- 1478 - 0x5c6  :  101 - 0x65
    "11111111", -- 1479 - 0x5c7  :  255 - 0xff
    "11111111", -- 1480 - 0x5c8  :  255 - 0xff -- Sprite 0xb9
    "00000001", -- 1481 - 0x5c9  :    1 - 0x1
    "00000011", -- 1482 - 0x5ca  :    3 - 0x3
    "00000001", -- 1483 - 0x5cb  :    1 - 0x1
    "00000011", -- 1484 - 0x5cc  :    3 - 0x3
    "00000001", -- 1485 - 0x5cd  :    1 - 0x1
    "10101011", -- 1486 - 0x5ce  :  171 - 0xab
    "11111111", -- 1487 - 0x5cf  :  255 - 0xff
    "11111111", -- 1488 - 0x5d0  :  255 - 0xff -- Sprite 0xba
    "11010101", -- 1489 - 0x5d1  :  213 - 0xd5
    "10101010", -- 1490 - 0x5d2  :  170 - 0xaa
    "11111111", -- 1491 - 0x5d3  :  255 - 0xff
    "10000000", -- 1492 - 0x5d4  :  128 - 0x80
    "10000000", -- 1493 - 0x5d5  :  128 - 0x80
    "10010101", -- 1494 - 0x5d6  :  149 - 0x95
    "11111111", -- 1495 - 0x5d7  :  255 - 0xff
    "00000000", -- 1496 - 0x5d8  :    0 - 0x0 -- Sprite 0xbb
    "00000000", -- 1497 - 0x5d9  :    0 - 0x0
    "00000000", -- 1498 - 0x5da  :    0 - 0x0
    "00000000", -- 1499 - 0x5db  :    0 - 0x0
    "00000000", -- 1500 - 0x5dc  :    0 - 0x0
    "00000000", -- 1501 - 0x5dd  :    0 - 0x0
    "00000000", -- 1502 - 0x5de  :    0 - 0x0
    "00000000", -- 1503 - 0x5df  :    0 - 0x0
    "11111111", -- 1504 - 0x5e0  :  255 - 0xff -- Sprite 0xbc
    "01010101", -- 1505 - 0x5e1  :   85 - 0x55
    "10101011", -- 1506 - 0x5e2  :  171 - 0xab
    "11111111", -- 1507 - 0x5e3  :  255 - 0xff
    "01100001", -- 1508 - 0x5e4  :   97 - 0x61
    "00100011", -- 1509 - 0x5e5  :   35 - 0x23
    "01100101", -- 1510 - 0x5e6  :  101 - 0x65
    "11111111", -- 1511 - 0x5e7  :  255 - 0xff
    "00000000", -- 1512 - 0x5e8  :    0 - 0x0 -- Sprite 0xbd
    "00000000", -- 1513 - 0x5e9  :    0 - 0x0
    "00000000", -- 1514 - 0x5ea  :    0 - 0x0
    "00000000", -- 1515 - 0x5eb  :    0 - 0x0
    "00000000", -- 1516 - 0x5ec  :    0 - 0x0
    "00000000", -- 1517 - 0x5ed  :    0 - 0x0
    "00000000", -- 1518 - 0x5ee  :    0 - 0x0
    "00000000", -- 1519 - 0x5ef  :    0 - 0x0
    "00000000", -- 1520 - 0x5f0  :    0 - 0x0 -- Sprite 0xbe
    "00000000", -- 1521 - 0x5f1  :    0 - 0x0
    "00000000", -- 1522 - 0x5f2  :    0 - 0x0
    "00000000", -- 1523 - 0x5f3  :    0 - 0x0
    "00000000", -- 1524 - 0x5f4  :    0 - 0x0
    "00000000", -- 1525 - 0x5f5  :    0 - 0x0
    "00000000", -- 1526 - 0x5f6  :    0 - 0x0
    "00000000", -- 1527 - 0x5f7  :    0 - 0x0
    "00000000", -- 1528 - 0x5f8  :    0 - 0x0 -- Sprite 0xbf
    "00000000", -- 1529 - 0x5f9  :    0 - 0x0
    "00000000", -- 1530 - 0x5fa  :    0 - 0x0
    "00000000", -- 1531 - 0x5fb  :    0 - 0x0
    "00000000", -- 1532 - 0x5fc  :    0 - 0x0
    "00000000", -- 1533 - 0x5fd  :    0 - 0x0
    "00000000", -- 1534 - 0x5fe  :    0 - 0x0
    "00000000", -- 1535 - 0x5ff  :    0 - 0x0
    "00000000", -- 1536 - 0x600  :    0 - 0x0 -- Sprite 0xc0
    "00000000", -- 1537 - 0x601  :    0 - 0x0
    "00000000", -- 1538 - 0x602  :    0 - 0x0
    "00000000", -- 1539 - 0x603  :    0 - 0x0
    "00000000", -- 1540 - 0x604  :    0 - 0x0
    "00000000", -- 1541 - 0x605  :    0 - 0x0
    "00000000", -- 1542 - 0x606  :    0 - 0x0
    "00000000", -- 1543 - 0x607  :    0 - 0x0
    "00000000", -- 1544 - 0x608  :    0 - 0x0 -- Sprite 0xc1
    "00000000", -- 1545 - 0x609  :    0 - 0x0
    "00000000", -- 1546 - 0x60a  :    0 - 0x0
    "00000000", -- 1547 - 0x60b  :    0 - 0x0
    "00000000", -- 1548 - 0x60c  :    0 - 0x0
    "00000000", -- 1549 - 0x60d  :    0 - 0x0
    "00000000", -- 1550 - 0x60e  :    0 - 0x0
    "00000000", -- 1551 - 0x60f  :    0 - 0x0
    "00000000", -- 1552 - 0x610  :    0 - 0x0 -- Sprite 0xc2
    "00000000", -- 1553 - 0x611  :    0 - 0x0
    "00000000", -- 1554 - 0x612  :    0 - 0x0
    "00000000", -- 1555 - 0x613  :    0 - 0x0
    "00000000", -- 1556 - 0x614  :    0 - 0x0
    "00000000", -- 1557 - 0x615  :    0 - 0x0
    "00000000", -- 1558 - 0x616  :    0 - 0x0
    "00000000", -- 1559 - 0x617  :    0 - 0x0
    "00000000", -- 1560 - 0x618  :    0 - 0x0 -- Sprite 0xc3
    "00000000", -- 1561 - 0x619  :    0 - 0x0
    "00000000", -- 1562 - 0x61a  :    0 - 0x0
    "00000000", -- 1563 - 0x61b  :    0 - 0x0
    "00000000", -- 1564 - 0x61c  :    0 - 0x0
    "00000000", -- 1565 - 0x61d  :    0 - 0x0
    "00000000", -- 1566 - 0x61e  :    0 - 0x0
    "00000000", -- 1567 - 0x61f  :    0 - 0x0
    "00000000", -- 1568 - 0x620  :    0 - 0x0 -- Sprite 0xc4
    "00000000", -- 1569 - 0x621  :    0 - 0x0
    "00000000", -- 1570 - 0x622  :    0 - 0x0
    "00000000", -- 1571 - 0x623  :    0 - 0x0
    "00000000", -- 1572 - 0x624  :    0 - 0x0
    "00000000", -- 1573 - 0x625  :    0 - 0x0
    "00000000", -- 1574 - 0x626  :    0 - 0x0
    "00000000", -- 1575 - 0x627  :    0 - 0x0
    "00000000", -- 1576 - 0x628  :    0 - 0x0 -- Sprite 0xc5
    "00000000", -- 1577 - 0x629  :    0 - 0x0
    "00000001", -- 1578 - 0x62a  :    1 - 0x1
    "00000110", -- 1579 - 0x62b  :    6 - 0x6
    "00001010", -- 1580 - 0x62c  :   10 - 0xa
    "00010100", -- 1581 - 0x62d  :   20 - 0x14
    "00010000", -- 1582 - 0x62e  :   16 - 0x10
    "00101000", -- 1583 - 0x62f  :   40 - 0x28
    "00011111", -- 1584 - 0x630  :   31 - 0x1f -- Sprite 0xc6
    "01100000", -- 1585 - 0x631  :   96 - 0x60
    "10100000", -- 1586 - 0x632  :  160 - 0xa0
    "01000000", -- 1587 - 0x633  :   64 - 0x40
    "00000000", -- 1588 - 0x634  :    0 - 0x0
    "00000000", -- 1589 - 0x635  :    0 - 0x0
    "00000000", -- 1590 - 0x636  :    0 - 0x0
    "00000000", -- 1591 - 0x637  :    0 - 0x0
    "00110000", -- 1592 - 0x638  :   48 - 0x30 -- Sprite 0xc7
    "01000000", -- 1593 - 0x639  :   64 - 0x40
    "01100000", -- 1594 - 0x63a  :   96 - 0x60
    "11000000", -- 1595 - 0x63b  :  192 - 0xc0
    "10000000", -- 1596 - 0x63c  :  128 - 0x80
    "10100000", -- 1597 - 0x63d  :  160 - 0xa0
    "11000000", -- 1598 - 0x63e  :  192 - 0xc0
    "10000000", -- 1599 - 0x63f  :  128 - 0x80
    "11111111", -- 1600 - 0x640  :  255 - 0xff -- Sprite 0xc8
    "00000000", -- 1601 - 0x641  :    0 - 0x0
    "00000000", -- 1602 - 0x642  :    0 - 0x0
    "00000000", -- 1603 - 0x643  :    0 - 0x0
    "00000000", -- 1604 - 0x644  :    0 - 0x0
    "00000000", -- 1605 - 0x645  :    0 - 0x0
    "00000000", -- 1606 - 0x646  :    0 - 0x0
    "00000000", -- 1607 - 0x647  :    0 - 0x0
    "00010100", -- 1608 - 0x648  :   20 - 0x14 -- Sprite 0xc9
    "00101010", -- 1609 - 0x649  :   42 - 0x2a
    "00010110", -- 1610 - 0x64a  :   22 - 0x16
    "00101011", -- 1611 - 0x64b  :   43 - 0x2b
    "00010101", -- 1612 - 0x64c  :   21 - 0x15
    "00101011", -- 1613 - 0x64d  :   43 - 0x2b
    "00010101", -- 1614 - 0x64e  :   21 - 0x15
    "00101011", -- 1615 - 0x64f  :   43 - 0x2b
    "00000000", -- 1616 - 0x650  :    0 - 0x0 -- Sprite 0xca
    "00000100", -- 1617 - 0x651  :    4 - 0x4
    "00000100", -- 1618 - 0x652  :    4 - 0x4
    "00000101", -- 1619 - 0x653  :    5 - 0x5
    "00010101", -- 1620 - 0x654  :   21 - 0x15
    "00010101", -- 1621 - 0x655  :   21 - 0x15
    "01010101", -- 1622 - 0x656  :   85 - 0x55
    "01010101", -- 1623 - 0x657  :   85 - 0x55
    "00000000", -- 1624 - 0x658  :    0 - 0x0 -- Sprite 0xcb
    "00000000", -- 1625 - 0x659  :    0 - 0x0
    "00010000", -- 1626 - 0x65a  :   16 - 0x10
    "00010000", -- 1627 - 0x65b  :   16 - 0x10
    "01010001", -- 1628 - 0x65c  :   81 - 0x51
    "01010101", -- 1629 - 0x65d  :   85 - 0x55
    "01010101", -- 1630 - 0x65e  :   85 - 0x55
    "01010101", -- 1631 - 0x65f  :   85 - 0x55
    "00000000", -- 1632 - 0x660  :    0 - 0x0 -- Sprite 0xcc
    "00000000", -- 1633 - 0x661  :    0 - 0x0
    "00000000", -- 1634 - 0x662  :    0 - 0x0
    "00000101", -- 1635 - 0x663  :    5 - 0x5
    "00001111", -- 1636 - 0x664  :   15 - 0xf
    "00000111", -- 1637 - 0x665  :    7 - 0x7
    "00000011", -- 1638 - 0x666  :    3 - 0x3
    "00000001", -- 1639 - 0x667  :    1 - 0x1
    "00000000", -- 1640 - 0x668  :    0 - 0x0 -- Sprite 0xcd
    "00000000", -- 1641 - 0x669  :    0 - 0x0
    "10000000", -- 1642 - 0x66a  :  128 - 0x80
    "11010000", -- 1643 - 0x66b  :  208 - 0xd0
    "11111000", -- 1644 - 0x66c  :  248 - 0xf8
    "11110000", -- 1645 - 0x66d  :  240 - 0xf0
    "11100000", -- 1646 - 0x66e  :  224 - 0xe0
    "11000000", -- 1647 - 0x66f  :  192 - 0xc0
    "00000000", -- 1648 - 0x670  :    0 - 0x0 -- Sprite 0xce
    "00000000", -- 1649 - 0x671  :    0 - 0x0
    "00000000", -- 1650 - 0x672  :    0 - 0x0
    "01111000", -- 1651 - 0x673  :  120 - 0x78
    "11001111", -- 1652 - 0x674  :  207 - 0xcf
    "10000000", -- 1653 - 0x675  :  128 - 0x80
    "11001111", -- 1654 - 0x676  :  207 - 0xcf
    "01001000", -- 1655 - 0x677  :   72 - 0x48
    "00000000", -- 1656 - 0x678  :    0 - 0x0 -- Sprite 0xcf
    "00000000", -- 1657 - 0x679  :    0 - 0x0
    "00000000", -- 1658 - 0x67a  :    0 - 0x0
    "00011110", -- 1659 - 0x67b  :   30 - 0x1e
    "11110011", -- 1660 - 0x67c  :  243 - 0xf3
    "00000001", -- 1661 - 0x67d  :    1 - 0x1
    "11110011", -- 1662 - 0x67e  :  243 - 0xf3
    "00010010", -- 1663 - 0x67f  :   18 - 0x12
    "00000000", -- 1664 - 0x680  :    0 - 0x0 -- Sprite 0xd0
    "00000000", -- 1665 - 0x681  :    0 - 0x0
    "00000000", -- 1666 - 0x682  :    0 - 0x0
    "00000000", -- 1667 - 0x683  :    0 - 0x0
    "00000000", -- 1668 - 0x684  :    0 - 0x0
    "00000000", -- 1669 - 0x685  :    0 - 0x0
    "00000000", -- 1670 - 0x686  :    0 - 0x0
    "00000000", -- 1671 - 0x687  :    0 - 0x0
    "00000000", -- 1672 - 0x688  :    0 - 0x0 -- Sprite 0xd1
    "00000000", -- 1673 - 0x689  :    0 - 0x0
    "00000000", -- 1674 - 0x68a  :    0 - 0x0
    "00000000", -- 1675 - 0x68b  :    0 - 0x0
    "00000000", -- 1676 - 0x68c  :    0 - 0x0
    "00000000", -- 1677 - 0x68d  :    0 - 0x0
    "00000000", -- 1678 - 0x68e  :    0 - 0x0
    "00000000", -- 1679 - 0x68f  :    0 - 0x0
    "00001000", -- 1680 - 0x690  :    8 - 0x8 -- Sprite 0xd2
    "00001100", -- 1681 - 0x691  :   12 - 0xc
    "00001000", -- 1682 - 0x692  :    8 - 0x8
    "00001000", -- 1683 - 0x693  :    8 - 0x8
    "00001010", -- 1684 - 0x694  :   10 - 0xa
    "00001000", -- 1685 - 0x695  :    8 - 0x8
    "00001000", -- 1686 - 0x696  :    8 - 0x8
    "00001100", -- 1687 - 0x697  :   12 - 0xc
    "00010000", -- 1688 - 0x698  :   16 - 0x10 -- Sprite 0xd3
    "00010000", -- 1689 - 0x699  :   16 - 0x10
    "00110000", -- 1690 - 0x69a  :   48 - 0x30
    "00010000", -- 1691 - 0x69b  :   16 - 0x10
    "01010000", -- 1692 - 0x69c  :   80 - 0x50
    "00010000", -- 1693 - 0x69d  :   16 - 0x10
    "00110000", -- 1694 - 0x69e  :   48 - 0x30
    "00010000", -- 1695 - 0x69f  :   16 - 0x10
    "00000000", -- 1696 - 0x6a0  :    0 - 0x0 -- Sprite 0xd4
    "00000000", -- 1697 - 0x6a1  :    0 - 0x0
    "00000000", -- 1698 - 0x6a2  :    0 - 0x0
    "00000000", -- 1699 - 0x6a3  :    0 - 0x0
    "00000000", -- 1700 - 0x6a4  :    0 - 0x0
    "00000000", -- 1701 - 0x6a5  :    0 - 0x0
    "00000000", -- 1702 - 0x6a6  :    0 - 0x0
    "00000000", -- 1703 - 0x6a7  :    0 - 0x0
    "11111000", -- 1704 - 0x6a8  :  248 - 0xf8 -- Sprite 0xd5
    "00000110", -- 1705 - 0x6a9  :    6 - 0x6
    "00000001", -- 1706 - 0x6aa  :    1 - 0x1
    "00000000", -- 1707 - 0x6ab  :    0 - 0x0
    "00000000", -- 1708 - 0x6ac  :    0 - 0x0
    "00000000", -- 1709 - 0x6ad  :    0 - 0x0
    "00000000", -- 1710 - 0x6ae  :    0 - 0x0
    "00000000", -- 1711 - 0x6af  :    0 - 0x0
    "00000000", -- 1712 - 0x6b0  :    0 - 0x0 -- Sprite 0xd6
    "00000000", -- 1713 - 0x6b1  :    0 - 0x0
    "10000000", -- 1714 - 0x6b2  :  128 - 0x80
    "01100000", -- 1715 - 0x6b3  :   96 - 0x60
    "01010000", -- 1716 - 0x6b4  :   80 - 0x50
    "10101000", -- 1717 - 0x6b5  :  168 - 0xa8
    "01011000", -- 1718 - 0x6b6  :   88 - 0x58
    "00101100", -- 1719 - 0x6b7  :   44 - 0x2c
    "10100000", -- 1720 - 0x6b8  :  160 - 0xa0 -- Sprite 0xd7
    "11000000", -- 1721 - 0x6b9  :  192 - 0xc0
    "10000000", -- 1722 - 0x6ba  :  128 - 0x80
    "01010000", -- 1723 - 0x6bb  :   80 - 0x50
    "01100000", -- 1724 - 0x6bc  :   96 - 0x60
    "00111000", -- 1725 - 0x6bd  :   56 - 0x38
    "00001000", -- 1726 - 0x6be  :    8 - 0x8
    "00000111", -- 1727 - 0x6bf  :    7 - 0x7
    "00000000", -- 1728 - 0x6c0  :    0 - 0x0 -- Sprite 0xd8
    "00000000", -- 1729 - 0x6c1  :    0 - 0x0
    "00000000", -- 1730 - 0x6c2  :    0 - 0x0
    "00000000", -- 1731 - 0x6c3  :    0 - 0x0
    "00000000", -- 1732 - 0x6c4  :    0 - 0x0
    "00000000", -- 1733 - 0x6c5  :    0 - 0x0
    "00000000", -- 1734 - 0x6c6  :    0 - 0x0
    "11111111", -- 1735 - 0x6c7  :  255 - 0xff
    "00010101", -- 1736 - 0x6c8  :   21 - 0x15 -- Sprite 0xd9
    "00101011", -- 1737 - 0x6c9  :   43 - 0x2b
    "00010101", -- 1738 - 0x6ca  :   21 - 0x15
    "00101010", -- 1739 - 0x6cb  :   42 - 0x2a
    "01010110", -- 1740 - 0x6cc  :   86 - 0x56
    "10101100", -- 1741 - 0x6cd  :  172 - 0xac
    "01010000", -- 1742 - 0x6ce  :   80 - 0x50
    "11100000", -- 1743 - 0x6cf  :  224 - 0xe0
    "00000001", -- 1744 - 0x6d0  :    1 - 0x1 -- Sprite 0xda
    "00001101", -- 1745 - 0x6d1  :   13 - 0xd
    "00010011", -- 1746 - 0x6d2  :   19 - 0x13
    "00001101", -- 1747 - 0x6d3  :   13 - 0xd
    "00000001", -- 1748 - 0x6d4  :    1 - 0x1
    "00000001", -- 1749 - 0x6d5  :    1 - 0x1
    "00000001", -- 1750 - 0x6d6  :    1 - 0x1
    "00000001", -- 1751 - 0x6d7  :    1 - 0x1
    "11000000", -- 1752 - 0x6d8  :  192 - 0xc0 -- Sprite 0xdb
    "01000000", -- 1753 - 0x6d9  :   64 - 0x40
    "01000000", -- 1754 - 0x6da  :   64 - 0x40
    "01011000", -- 1755 - 0x6db  :   88 - 0x58
    "01100100", -- 1756 - 0x6dc  :  100 - 0x64
    "01011000", -- 1757 - 0x6dd  :   88 - 0x58
    "01000000", -- 1758 - 0x6de  :   64 - 0x40
    "01000000", -- 1759 - 0x6df  :   64 - 0x40
    "00000000", -- 1760 - 0x6e0  :    0 - 0x0 -- Sprite 0xdc
    "00000000", -- 1761 - 0x6e1  :    0 - 0x0
    "00000000", -- 1762 - 0x6e2  :    0 - 0x0
    "00000110", -- 1763 - 0x6e3  :    6 - 0x6
    "00000111", -- 1764 - 0x6e4  :    7 - 0x7
    "00000111", -- 1765 - 0x6e5  :    7 - 0x7
    "00000111", -- 1766 - 0x6e6  :    7 - 0x7
    "00000011", -- 1767 - 0x6e7  :    3 - 0x3
    "00000000", -- 1768 - 0x6e8  :    0 - 0x0 -- Sprite 0xdd
    "00000000", -- 1769 - 0x6e9  :    0 - 0x0
    "00000000", -- 1770 - 0x6ea  :    0 - 0x0
    "10110000", -- 1771 - 0x6eb  :  176 - 0xb0
    "11110000", -- 1772 - 0x6ec  :  240 - 0xf0
    "11110000", -- 1773 - 0x6ed  :  240 - 0xf0
    "11110000", -- 1774 - 0x6ee  :  240 - 0xf0
    "11100000", -- 1775 - 0x6ef  :  224 - 0xe0
    "11001111", -- 1776 - 0x6f0  :  207 - 0xcf -- Sprite 0xde
    "10000000", -- 1777 - 0x6f1  :  128 - 0x80
    "11001111", -- 1778 - 0x6f2  :  207 - 0xcf
    "01001000", -- 1779 - 0x6f3  :   72 - 0x48
    "01001000", -- 1780 - 0x6f4  :   72 - 0x48
    "01001000", -- 1781 - 0x6f5  :   72 - 0x48
    "01001000", -- 1782 - 0x6f6  :   72 - 0x48
    "01001000", -- 1783 - 0x6f7  :   72 - 0x48
    "11110011", -- 1784 - 0x6f8  :  243 - 0xf3 -- Sprite 0xdf
    "00000001", -- 1785 - 0x6f9  :    1 - 0x1
    "11110011", -- 1786 - 0x6fa  :  243 - 0xf3
    "00010010", -- 1787 - 0x6fb  :   18 - 0x12
    "00010010", -- 1788 - 0x6fc  :   18 - 0x12
    "00010010", -- 1789 - 0x6fd  :   18 - 0x12
    "00010010", -- 1790 - 0x6fe  :   18 - 0x12
    "00010010", -- 1791 - 0x6ff  :   18 - 0x12
    "00000000", -- 1792 - 0x700  :    0 - 0x0 -- Sprite 0xe0
    "00000000", -- 1793 - 0x701  :    0 - 0x0
    "00000000", -- 1794 - 0x702  :    0 - 0x0
    "00000000", -- 1795 - 0x703  :    0 - 0x0
    "00000000", -- 1796 - 0x704  :    0 - 0x0
    "00000000", -- 1797 - 0x705  :    0 - 0x0
    "00000000", -- 1798 - 0x706  :    0 - 0x0
    "00000000", -- 1799 - 0x707  :    0 - 0x0
    "00000000", -- 1800 - 0x708  :    0 - 0x0 -- Sprite 0xe1
    "00000000", -- 1801 - 0x709  :    0 - 0x0
    "00000000", -- 1802 - 0x70a  :    0 - 0x0
    "00000000", -- 1803 - 0x70b  :    0 - 0x0
    "00000000", -- 1804 - 0x70c  :    0 - 0x0
    "00000000", -- 1805 - 0x70d  :    0 - 0x0
    "00000000", -- 1806 - 0x70e  :    0 - 0x0
    "00000000", -- 1807 - 0x70f  :    0 - 0x0
    "00000000", -- 1808 - 0x710  :    0 - 0x0 -- Sprite 0xe2
    "00000000", -- 1809 - 0x711  :    0 - 0x0
    "00000000", -- 1810 - 0x712  :    0 - 0x0
    "00000000", -- 1811 - 0x713  :    0 - 0x0
    "00000000", -- 1812 - 0x714  :    0 - 0x0
    "00000000", -- 1813 - 0x715  :    0 - 0x0
    "00000000", -- 1814 - 0x716  :    0 - 0x0
    "00000000", -- 1815 - 0x717  :    0 - 0x0
    "00000000", -- 1816 - 0x718  :    0 - 0x0 -- Sprite 0xe3
    "00000000", -- 1817 - 0x719  :    0 - 0x0
    "00000000", -- 1818 - 0x71a  :    0 - 0x0
    "00000000", -- 1819 - 0x71b  :    0 - 0x0
    "00000000", -- 1820 - 0x71c  :    0 - 0x0
    "00000000", -- 1821 - 0x71d  :    0 - 0x0
    "00000000", -- 1822 - 0x71e  :    0 - 0x0
    "00000000", -- 1823 - 0x71f  :    0 - 0x0
    "00000000", -- 1824 - 0x720  :    0 - 0x0 -- Sprite 0xe4
    "00000000", -- 1825 - 0x721  :    0 - 0x0
    "00000000", -- 1826 - 0x722  :    0 - 0x0
    "00000000", -- 1827 - 0x723  :    0 - 0x0
    "00000000", -- 1828 - 0x724  :    0 - 0x0
    "00000000", -- 1829 - 0x725  :    0 - 0x0
    "00000000", -- 1830 - 0x726  :    0 - 0x0
    "00000000", -- 1831 - 0x727  :    0 - 0x0
    "00000000", -- 1832 - 0x728  :    0 - 0x0 -- Sprite 0xe5
    "00000000", -- 1833 - 0x729  :    0 - 0x0
    "00000000", -- 1834 - 0x72a  :    0 - 0x0
    "00000000", -- 1835 - 0x72b  :    0 - 0x0
    "00000000", -- 1836 - 0x72c  :    0 - 0x0
    "00000000", -- 1837 - 0x72d  :    0 - 0x0
    "00000000", -- 1838 - 0x72e  :    0 - 0x0
    "00000000", -- 1839 - 0x72f  :    0 - 0x0
    "00000000", -- 1840 - 0x730  :    0 - 0x0 -- Sprite 0xe6
    "00000000", -- 1841 - 0x731  :    0 - 0x0
    "00000000", -- 1842 - 0x732  :    0 - 0x0
    "00000000", -- 1843 - 0x733  :    0 - 0x0
    "00000000", -- 1844 - 0x734  :    0 - 0x0
    "00000000", -- 1845 - 0x735  :    0 - 0x0
    "00000000", -- 1846 - 0x736  :    0 - 0x0
    "00000000", -- 1847 - 0x737  :    0 - 0x0
    "00000000", -- 1848 - 0x738  :    0 - 0x0 -- Sprite 0xe7
    "00000000", -- 1849 - 0x739  :    0 - 0x0
    "00000000", -- 1850 - 0x73a  :    0 - 0x0
    "00000000", -- 1851 - 0x73b  :    0 - 0x0
    "00000000", -- 1852 - 0x73c  :    0 - 0x0
    "00000000", -- 1853 - 0x73d  :    0 - 0x0
    "00000000", -- 1854 - 0x73e  :    0 - 0x0
    "00000000", -- 1855 - 0x73f  :    0 - 0x0
    "00000000", -- 1856 - 0x740  :    0 - 0x0 -- Sprite 0xe8
    "00000000", -- 1857 - 0x741  :    0 - 0x0
    "00000000", -- 1858 - 0x742  :    0 - 0x0
    "00000000", -- 1859 - 0x743  :    0 - 0x0
    "00000000", -- 1860 - 0x744  :    0 - 0x0
    "00000000", -- 1861 - 0x745  :    0 - 0x0
    "00000000", -- 1862 - 0x746  :    0 - 0x0
    "00000000", -- 1863 - 0x747  :    0 - 0x0
    "00000000", -- 1864 - 0x748  :    0 - 0x0 -- Sprite 0xe9
    "00000000", -- 1865 - 0x749  :    0 - 0x0
    "00000000", -- 1866 - 0x74a  :    0 - 0x0
    "00000000", -- 1867 - 0x74b  :    0 - 0x0
    "00000000", -- 1868 - 0x74c  :    0 - 0x0
    "00000000", -- 1869 - 0x74d  :    0 - 0x0
    "00000000", -- 1870 - 0x74e  :    0 - 0x0
    "00000000", -- 1871 - 0x74f  :    0 - 0x0
    "00000000", -- 1872 - 0x750  :    0 - 0x0 -- Sprite 0xea
    "00000000", -- 1873 - 0x751  :    0 - 0x0
    "00000000", -- 1874 - 0x752  :    0 - 0x0
    "00000000", -- 1875 - 0x753  :    0 - 0x0
    "00000000", -- 1876 - 0x754  :    0 - 0x0
    "00000000", -- 1877 - 0x755  :    0 - 0x0
    "00000000", -- 1878 - 0x756  :    0 - 0x0
    "00000000", -- 1879 - 0x757  :    0 - 0x0
    "00000000", -- 1880 - 0x758  :    0 - 0x0 -- Sprite 0xeb
    "00000000", -- 1881 - 0x759  :    0 - 0x0
    "00000000", -- 1882 - 0x75a  :    0 - 0x0
    "00000000", -- 1883 - 0x75b  :    0 - 0x0
    "00000000", -- 1884 - 0x75c  :    0 - 0x0
    "00000000", -- 1885 - 0x75d  :    0 - 0x0
    "00000000", -- 1886 - 0x75e  :    0 - 0x0
    "00000000", -- 1887 - 0x75f  :    0 - 0x0
    "00000000", -- 1888 - 0x760  :    0 - 0x0 -- Sprite 0xec
    "00000000", -- 1889 - 0x761  :    0 - 0x0
    "00000000", -- 1890 - 0x762  :    0 - 0x0
    "00000000", -- 1891 - 0x763  :    0 - 0x0
    "00000000", -- 1892 - 0x764  :    0 - 0x0
    "00000000", -- 1893 - 0x765  :    0 - 0x0
    "00000000", -- 1894 - 0x766  :    0 - 0x0
    "00000000", -- 1895 - 0x767  :    0 - 0x0
    "00000000", -- 1896 - 0x768  :    0 - 0x0 -- Sprite 0xed
    "00000000", -- 1897 - 0x769  :    0 - 0x0
    "00000000", -- 1898 - 0x76a  :    0 - 0x0
    "00000000", -- 1899 - 0x76b  :    0 - 0x0
    "00000000", -- 1900 - 0x76c  :    0 - 0x0
    "00000000", -- 1901 - 0x76d  :    0 - 0x0
    "00000000", -- 1902 - 0x76e  :    0 - 0x0
    "00000000", -- 1903 - 0x76f  :    0 - 0x0
    "00000000", -- 1904 - 0x770  :    0 - 0x0 -- Sprite 0xee
    "00000000", -- 1905 - 0x771  :    0 - 0x0
    "00000000", -- 1906 - 0x772  :    0 - 0x0
    "00000000", -- 1907 - 0x773  :    0 - 0x0
    "00000000", -- 1908 - 0x774  :    0 - 0x0
    "00000000", -- 1909 - 0x775  :    0 - 0x0
    "00000000", -- 1910 - 0x776  :    0 - 0x0
    "00000000", -- 1911 - 0x777  :    0 - 0x0
    "00000000", -- 1912 - 0x778  :    0 - 0x0 -- Sprite 0xef
    "00000000", -- 1913 - 0x779  :    0 - 0x0
    "00000000", -- 1914 - 0x77a  :    0 - 0x0
    "00000000", -- 1915 - 0x77b  :    0 - 0x0
    "00000000", -- 1916 - 0x77c  :    0 - 0x0
    "00000000", -- 1917 - 0x77d  :    0 - 0x0
    "00000000", -- 1918 - 0x77e  :    0 - 0x0
    "00000000", -- 1919 - 0x77f  :    0 - 0x0
    "00000000", -- 1920 - 0x780  :    0 - 0x0 -- Sprite 0xf0
    "00000000", -- 1921 - 0x781  :    0 - 0x0
    "00000000", -- 1922 - 0x782  :    0 - 0x0
    "00000000", -- 1923 - 0x783  :    0 - 0x0
    "00000000", -- 1924 - 0x784  :    0 - 0x0
    "00000000", -- 1925 - 0x785  :    0 - 0x0
    "00000000", -- 1926 - 0x786  :    0 - 0x0
    "00000000", -- 1927 - 0x787  :    0 - 0x0
    "00000000", -- 1928 - 0x788  :    0 - 0x0 -- Sprite 0xf1
    "00000000", -- 1929 - 0x789  :    0 - 0x0
    "00000000", -- 1930 - 0x78a  :    0 - 0x0
    "00000000", -- 1931 - 0x78b  :    0 - 0x0
    "00000000", -- 1932 - 0x78c  :    0 - 0x0
    "00000000", -- 1933 - 0x78d  :    0 - 0x0
    "00000000", -- 1934 - 0x78e  :    0 - 0x0
    "00000000", -- 1935 - 0x78f  :    0 - 0x0
    "00000000", -- 1936 - 0x790  :    0 - 0x0 -- Sprite 0xf2
    "00000000", -- 1937 - 0x791  :    0 - 0x0
    "00000000", -- 1938 - 0x792  :    0 - 0x0
    "00000000", -- 1939 - 0x793  :    0 - 0x0
    "00000000", -- 1940 - 0x794  :    0 - 0x0
    "00000000", -- 1941 - 0x795  :    0 - 0x0
    "00000000", -- 1942 - 0x796  :    0 - 0x0
    "00000000", -- 1943 - 0x797  :    0 - 0x0
    "00000000", -- 1944 - 0x798  :    0 - 0x0 -- Sprite 0xf3
    "00000000", -- 1945 - 0x799  :    0 - 0x0
    "00000000", -- 1946 - 0x79a  :    0 - 0x0
    "00000000", -- 1947 - 0x79b  :    0 - 0x0
    "00000000", -- 1948 - 0x79c  :    0 - 0x0
    "00000000", -- 1949 - 0x79d  :    0 - 0x0
    "00000000", -- 1950 - 0x79e  :    0 - 0x0
    "00000000", -- 1951 - 0x79f  :    0 - 0x0
    "00000000", -- 1952 - 0x7a0  :    0 - 0x0 -- Sprite 0xf4
    "00000000", -- 1953 - 0x7a1  :    0 - 0x0
    "00000000", -- 1954 - 0x7a2  :    0 - 0x0
    "00000000", -- 1955 - 0x7a3  :    0 - 0x0
    "00000000", -- 1956 - 0x7a4  :    0 - 0x0
    "00000000", -- 1957 - 0x7a5  :    0 - 0x0
    "00000000", -- 1958 - 0x7a6  :    0 - 0x0
    "00000000", -- 1959 - 0x7a7  :    0 - 0x0
    "00000000", -- 1960 - 0x7a8  :    0 - 0x0 -- Sprite 0xf5
    "00000000", -- 1961 - 0x7a9  :    0 - 0x0
    "00000000", -- 1962 - 0x7aa  :    0 - 0x0
    "00000000", -- 1963 - 0x7ab  :    0 - 0x0
    "00000000", -- 1964 - 0x7ac  :    0 - 0x0
    "00000000", -- 1965 - 0x7ad  :    0 - 0x0
    "00000000", -- 1966 - 0x7ae  :    0 - 0x0
    "00000000", -- 1967 - 0x7af  :    0 - 0x0
    "00000000", -- 1968 - 0x7b0  :    0 - 0x0 -- Sprite 0xf6
    "00000000", -- 1969 - 0x7b1  :    0 - 0x0
    "00000000", -- 1970 - 0x7b2  :    0 - 0x0
    "00000000", -- 1971 - 0x7b3  :    0 - 0x0
    "00000000", -- 1972 - 0x7b4  :    0 - 0x0
    "00000000", -- 1973 - 0x7b5  :    0 - 0x0
    "00000000", -- 1974 - 0x7b6  :    0 - 0x0
    "00000000", -- 1975 - 0x7b7  :    0 - 0x0
    "00000000", -- 1976 - 0x7b8  :    0 - 0x0 -- Sprite 0xf7
    "00000000", -- 1977 - 0x7b9  :    0 - 0x0
    "00000000", -- 1978 - 0x7ba  :    0 - 0x0
    "00000000", -- 1979 - 0x7bb  :    0 - 0x0
    "00000000", -- 1980 - 0x7bc  :    0 - 0x0
    "00000000", -- 1981 - 0x7bd  :    0 - 0x0
    "00000000", -- 1982 - 0x7be  :    0 - 0x0
    "00000000", -- 1983 - 0x7bf  :    0 - 0x0
    "00000000", -- 1984 - 0x7c0  :    0 - 0x0 -- Sprite 0xf8
    "00000000", -- 1985 - 0x7c1  :    0 - 0x0
    "00000000", -- 1986 - 0x7c2  :    0 - 0x0
    "00000000", -- 1987 - 0x7c3  :    0 - 0x0
    "00000000", -- 1988 - 0x7c4  :    0 - 0x0
    "00000000", -- 1989 - 0x7c5  :    0 - 0x0
    "00000000", -- 1990 - 0x7c6  :    0 - 0x0
    "00000000", -- 1991 - 0x7c7  :    0 - 0x0
    "00000000", -- 1992 - 0x7c8  :    0 - 0x0 -- Sprite 0xf9
    "00000000", -- 1993 - 0x7c9  :    0 - 0x0
    "00000000", -- 1994 - 0x7ca  :    0 - 0x0
    "00000000", -- 1995 - 0x7cb  :    0 - 0x0
    "00000000", -- 1996 - 0x7cc  :    0 - 0x0
    "00000000", -- 1997 - 0x7cd  :    0 - 0x0
    "00000000", -- 1998 - 0x7ce  :    0 - 0x0
    "00000000", -- 1999 - 0x7cf  :    0 - 0x0
    "00000000", -- 2000 - 0x7d0  :    0 - 0x0 -- Sprite 0xfa
    "00000000", -- 2001 - 0x7d1  :    0 - 0x0
    "00000000", -- 2002 - 0x7d2  :    0 - 0x0
    "00000000", -- 2003 - 0x7d3  :    0 - 0x0
    "00000000", -- 2004 - 0x7d4  :    0 - 0x0
    "00000000", -- 2005 - 0x7d5  :    0 - 0x0
    "00000000", -- 2006 - 0x7d6  :    0 - 0x0
    "00000000", -- 2007 - 0x7d7  :    0 - 0x0
    "00000000", -- 2008 - 0x7d8  :    0 - 0x0 -- Sprite 0xfb
    "00000000", -- 2009 - 0x7d9  :    0 - 0x0
    "00000000", -- 2010 - 0x7da  :    0 - 0x0
    "00000000", -- 2011 - 0x7db  :    0 - 0x0
    "00000000", -- 2012 - 0x7dc  :    0 - 0x0
    "00000000", -- 2013 - 0x7dd  :    0 - 0x0
    "00000000", -- 2014 - 0x7de  :    0 - 0x0
    "00000000", -- 2015 - 0x7df  :    0 - 0x0
    "00000000", -- 2016 - 0x7e0  :    0 - 0x0 -- Sprite 0xfc
    "00000000", -- 2017 - 0x7e1  :    0 - 0x0
    "10001110", -- 2018 - 0x7e2  :  142 - 0x8e
    "10001010", -- 2019 - 0x7e3  :  138 - 0x8a
    "10001010", -- 2020 - 0x7e4  :  138 - 0x8a
    "10001010", -- 2021 - 0x7e5  :  138 - 0x8a
    "10001010", -- 2022 - 0x7e6  :  138 - 0x8a
    "11101110", -- 2023 - 0x7e7  :  238 - 0xee
    "00000000", -- 2024 - 0x7e8  :    0 - 0x0 -- Sprite 0xfd
    "00000000", -- 2025 - 0x7e9  :    0 - 0x0
    "01001100", -- 2026 - 0x7ea  :   76 - 0x4c
    "10101010", -- 2027 - 0x7eb  :  170 - 0xaa
    "10101010", -- 2028 - 0x7ec  :  170 - 0xaa
    "11101010", -- 2029 - 0x7ed  :  234 - 0xea
    "10101010", -- 2030 - 0x7ee  :  170 - 0xaa
    "10101100", -- 2031 - 0x7ef  :  172 - 0xac
    "00000000", -- 2032 - 0x7f0  :    0 - 0x0 -- Sprite 0xfe
    "00000000", -- 2033 - 0x7f1  :    0 - 0x0
    "11101100", -- 2034 - 0x7f2  :  236 - 0xec
    "01001010", -- 2035 - 0x7f3  :   74 - 0x4a
    "01001010", -- 2036 - 0x7f4  :   74 - 0x4a
    "01001010", -- 2037 - 0x7f5  :   74 - 0x4a
    "01001010", -- 2038 - 0x7f6  :   74 - 0x4a
    "11101010", -- 2039 - 0x7f7  :  234 - 0xea
    "00000000", -- 2040 - 0x7f8  :    0 - 0x0 -- Sprite 0xff
    "00000000", -- 2041 - 0x7f9  :    0 - 0x0
    "01100000", -- 2042 - 0x7fa  :   96 - 0x60
    "10001000", -- 2043 - 0x7fb  :  136 - 0x88
    "10100000", -- 2044 - 0x7fc  :  160 - 0xa0
    "10100000", -- 2045 - 0x7fd  :  160 - 0xa0
    "10101000", -- 2046 - 0x7fe  :  168 - 0xa8
    "01000000", -- 2047 - 0x7ff  :   64 - 0x40
          -- Background pattern Table
    "00000000", -- 2048 - 0x800  :    0 - 0x0 -- Background 0x0
    "00001111", -- 2049 - 0x801  :   15 - 0xf
    "00000100", -- 2050 - 0x802  :    4 - 0x4
    "00000011", -- 2051 - 0x803  :    3 - 0x3
    "00000011", -- 2052 - 0x804  :    3 - 0x3
    "00000011", -- 2053 - 0x805  :    3 - 0x3
    "00000100", -- 2054 - 0x806  :    4 - 0x4
    "00111010", -- 2055 - 0x807  :   58 - 0x3a
    "00000000", -- 2056 - 0x808  :    0 - 0x0 -- Background 0x1
    "00111000", -- 2057 - 0x809  :   56 - 0x38
    "11000110", -- 2058 - 0x80a  :  198 - 0xc6
    "11001011", -- 2059 - 0x80b  :  203 - 0xcb
    "11011100", -- 2060 - 0x80c  :  220 - 0xdc
    "00111010", -- 2061 - 0x80d  :   58 - 0x3a
    "10011010", -- 2062 - 0x80e  :  154 - 0x9a
    "10000001", -- 2063 - 0x80f  :  129 - 0x81
    "01000101", -- 2064 - 0x810  :   69 - 0x45 -- Background 0x2
    "10000111", -- 2065 - 0x811  :  135 - 0x87
    "10000011", -- 2066 - 0x812  :  131 - 0x83
    "10000001", -- 2067 - 0x813  :  129 - 0x81
    "10000001", -- 2068 - 0x814  :  129 - 0x81
    "10000001", -- 2069 - 0x815  :  129 - 0x81
    "01000001", -- 2070 - 0x816  :   65 - 0x41
    "00100001", -- 2071 - 0x817  :   33 - 0x21
    "01111111", -- 2072 - 0x818  :  127 - 0x7f -- Background 0x3
    "01111110", -- 2073 - 0x819  :  126 - 0x7e
    "11111100", -- 2074 - 0x81a  :  252 - 0xfc
    "00111000", -- 2075 - 0x81b  :   56 - 0x38
    "00011000", -- 2076 - 0x81c  :   24 - 0x18
    "10001100", -- 2077 - 0x81d  :  140 - 0x8c
    "11000100", -- 2078 - 0x81e  :  196 - 0xc4
    "11111100", -- 2079 - 0x81f  :  252 - 0xfc
    "00100011", -- 2080 - 0x820  :   35 - 0x23 -- Background 0x4
    "00100011", -- 2081 - 0x821  :   35 - 0x23
    "00100001", -- 2082 - 0x822  :   33 - 0x21
    "00100000", -- 2083 - 0x823  :   32 - 0x20
    "00010011", -- 2084 - 0x824  :   19 - 0x13
    "00001100", -- 2085 - 0x825  :   12 - 0xc
    "00000000", -- 2086 - 0x826  :    0 - 0x0
    "00000000", -- 2087 - 0x827  :    0 - 0x0
    "11111100", -- 2088 - 0x828  :  252 - 0xfc -- Background 0x5
    "11111100", -- 2089 - 0x829  :  252 - 0xfc
    "11111100", -- 2090 - 0x82a  :  252 - 0xfc
    "11111100", -- 2091 - 0x82b  :  252 - 0xfc
    "10010000", -- 2092 - 0x82c  :  144 - 0x90
    "10010000", -- 2093 - 0x82d  :  144 - 0x90
    "10001000", -- 2094 - 0x82e  :  136 - 0x88
    "11111000", -- 2095 - 0x82f  :  248 - 0xf8
    "00100011", -- 2096 - 0x830  :   35 - 0x23 -- Background 0x6
    "00100011", -- 2097 - 0x831  :   35 - 0x23
    "00100001", -- 2098 - 0x832  :   33 - 0x21
    "00100000", -- 2099 - 0x833  :   32 - 0x20
    "00010011", -- 2100 - 0x834  :   19 - 0x13
    "00001101", -- 2101 - 0x835  :   13 - 0xd
    "00000010", -- 2102 - 0x836  :    2 - 0x2
    "00000001", -- 2103 - 0x837  :    1 - 0x1
    "11111100", -- 2104 - 0x838  :  252 - 0xfc -- Background 0x7
    "11111100", -- 2105 - 0x839  :  252 - 0xfc
    "11111100", -- 2106 - 0x83a  :  252 - 0xfc
    "11111100", -- 2107 - 0x83b  :  252 - 0xfc
    "10100100", -- 2108 - 0x83c  :  164 - 0xa4
    "00100100", -- 2109 - 0x83d  :   36 - 0x24
    "01010010", -- 2110 - 0x83e  :   82 - 0x52
    "11101110", -- 2111 - 0x83f  :  238 - 0xee
    "00100011", -- 2112 - 0x840  :   35 - 0x23 -- Background 0x8
    "00100011", -- 2113 - 0x841  :   35 - 0x23
    "00100001", -- 2114 - 0x842  :   33 - 0x21
    "00100000", -- 2115 - 0x843  :   32 - 0x20
    "00010011", -- 2116 - 0x844  :   19 - 0x13
    "00001101", -- 2117 - 0x845  :   13 - 0xd
    "00000001", -- 2118 - 0x846  :    1 - 0x1
    "00000001", -- 2119 - 0x847  :    1 - 0x1
    "11111110", -- 2120 - 0x848  :  254 - 0xfe -- Background 0x9
    "11111110", -- 2121 - 0x849  :  254 - 0xfe
    "11111110", -- 2122 - 0x84a  :  254 - 0xfe
    "11111111", -- 2123 - 0x84b  :  255 - 0xff
    "10010001", -- 2124 - 0x84c  :  145 - 0x91
    "00101111", -- 2125 - 0x84d  :   47 - 0x2f
    "01000000", -- 2126 - 0x84e  :   64 - 0x40
    "11100000", -- 2127 - 0x84f  :  224 - 0xe0
    "00100011", -- 2128 - 0x850  :   35 - 0x23 -- Background 0xa
    "00100011", -- 2129 - 0x851  :   35 - 0x23
    "00100001", -- 2130 - 0x852  :   33 - 0x21
    "00100000", -- 2131 - 0x853  :   32 - 0x20
    "00010011", -- 2132 - 0x854  :   19 - 0x13
    "00001110", -- 2133 - 0x855  :   14 - 0xe
    "00000001", -- 2134 - 0x856  :    1 - 0x1
    "00000000", -- 2135 - 0x857  :    0 - 0x0
    "11111110", -- 2136 - 0x858  :  254 - 0xfe -- Background 0xb
    "11111110", -- 2137 - 0x859  :  254 - 0xfe
    "11111110", -- 2138 - 0x85a  :  254 - 0xfe
    "11111100", -- 2139 - 0x85b  :  252 - 0xfc
    "00100100", -- 2140 - 0x85c  :   36 - 0x24
    "00100010", -- 2141 - 0x85d  :   34 - 0x22
    "11010010", -- 2142 - 0x85e  :  210 - 0xd2
    "00001111", -- 2143 - 0x85f  :   15 - 0xf
    "01111111", -- 2144 - 0x860  :  127 - 0x7f -- Background 0xc
    "01111110", -- 2145 - 0x861  :  126 - 0x7e
    "11111100", -- 2146 - 0x862  :  252 - 0xfc
    "00000010", -- 2147 - 0x863  :    2 - 0x2
    "00000100", -- 2148 - 0x864  :    4 - 0x4
    "11111100", -- 2149 - 0x865  :  252 - 0xfc
    "11111100", -- 2150 - 0x866  :  252 - 0xfc
    "11111110", -- 2151 - 0x867  :  254 - 0xfe
    "01000101", -- 2152 - 0x868  :   69 - 0x45 -- Background 0xd
    "10000111", -- 2153 - 0x869  :  135 - 0x87
    "10000011", -- 2154 - 0x86a  :  131 - 0x83
    "10000010", -- 2155 - 0x86b  :  130 - 0x82
    "10000010", -- 2156 - 0x86c  :  130 - 0x82
    "10000100", -- 2157 - 0x86d  :  132 - 0x84
    "01000100", -- 2158 - 0x86e  :   68 - 0x44
    "00100100", -- 2159 - 0x86f  :   36 - 0x24
    "01111111", -- 2160 - 0x870  :  127 - 0x7f -- Background 0xe
    "01111110", -- 2161 - 0x871  :  126 - 0x7e
    "11111100", -- 2162 - 0x872  :  252 - 0xfc
    "11111000", -- 2163 - 0x873  :  248 - 0xf8
    "01111000", -- 2164 - 0x874  :  120 - 0x78
    "01111100", -- 2165 - 0x875  :  124 - 0x7c
    "11111100", -- 2166 - 0x876  :  252 - 0xfc
    "11111110", -- 2167 - 0x877  :  254 - 0xfe
    "00000000", -- 2168 - 0x878  :    0 - 0x0 -- Background 0xf
    "00001111", -- 2169 - 0x879  :   15 - 0xf
    "00000100", -- 2170 - 0x87a  :    4 - 0x4
    "00000011", -- 2171 - 0x87b  :    3 - 0x3
    "00000011", -- 2172 - 0x87c  :    3 - 0x3
    "00000011", -- 2173 - 0x87d  :    3 - 0x3
    "00000100", -- 2174 - 0x87e  :    4 - 0x4
    "00000010", -- 2175 - 0x87f  :    2 - 0x2
    "00000111", -- 2176 - 0x880  :    7 - 0x7 -- Background 0x10
    "00001100", -- 2177 - 0x881  :   12 - 0xc
    "00010000", -- 2178 - 0x882  :   16 - 0x10
    "00010000", -- 2179 - 0x883  :   16 - 0x10
    "00010000", -- 2180 - 0x884  :   16 - 0x10
    "00100000", -- 2181 - 0x885  :   32 - 0x20
    "00100000", -- 2182 - 0x886  :   32 - 0x20
    "00100001", -- 2183 - 0x887  :   33 - 0x21
    "11111111", -- 2184 - 0x888  :  255 - 0xff -- Background 0x11
    "01111110", -- 2185 - 0x889  :  126 - 0x7e
    "01111100", -- 2186 - 0x88a  :  124 - 0x7c
    "01111000", -- 2187 - 0x88b  :  120 - 0x78
    "01011000", -- 2188 - 0x88c  :   88 - 0x58
    "10001100", -- 2189 - 0x88d  :  140 - 0x8c
    "11000100", -- 2190 - 0x88e  :  196 - 0xc4
    "11111100", -- 2191 - 0x88f  :  252 - 0xfc
    "00100011", -- 2192 - 0x890  :   35 - 0x23 -- Background 0x12
    "00100011", -- 2193 - 0x891  :   35 - 0x23
    "00100001", -- 2194 - 0x892  :   33 - 0x21
    "00100000", -- 2195 - 0x893  :   32 - 0x20
    "00010011", -- 2196 - 0x894  :   19 - 0x13
    "00001100", -- 2197 - 0x895  :   12 - 0xc
    "00000000", -- 2198 - 0x896  :    0 - 0x0
    "00000000", -- 2199 - 0x897  :    0 - 0x0
    "00000001", -- 2200 - 0x898  :    1 - 0x1 -- Background 0x13
    "00000001", -- 2201 - 0x899  :    1 - 0x1
    "00000011", -- 2202 - 0x89a  :    3 - 0x3
    "00000100", -- 2203 - 0x89b  :    4 - 0x4
    "00001000", -- 2204 - 0x89c  :    8 - 0x8
    "00010000", -- 2205 - 0x89d  :   16 - 0x10
    "00010000", -- 2206 - 0x89e  :   16 - 0x10
    "00100000", -- 2207 - 0x89f  :   32 - 0x20
    "01111111", -- 2208 - 0x8a0  :  127 - 0x7f -- Background 0x14
    "11111110", -- 2209 - 0x8a1  :  254 - 0xfe
    "00000110", -- 2210 - 0x8a2  :    6 - 0x6
    "00000001", -- 2211 - 0x8a3  :    1 - 0x1
    "00000001", -- 2212 - 0x8a4  :    1 - 0x1
    "00000001", -- 2213 - 0x8a5  :    1 - 0x1
    "00000111", -- 2214 - 0x8a6  :    7 - 0x7
    "11111110", -- 2215 - 0x8a7  :  254 - 0xfe
    "00000101", -- 2216 - 0x8a8  :    5 - 0x5 -- Background 0x15
    "00000101", -- 2217 - 0x8a9  :    5 - 0x5
    "00000111", -- 2218 - 0x8aa  :    7 - 0x7
    "00000100", -- 2219 - 0x8ab  :    4 - 0x4
    "00000100", -- 2220 - 0x8ac  :    4 - 0x4
    "00001111", -- 2221 - 0x8ad  :   15 - 0xf
    "00110000", -- 2222 - 0x8ae  :   48 - 0x30
    "01000000", -- 2223 - 0x8af  :   64 - 0x40
    "11111100", -- 2224 - 0x8b0  :  252 - 0xfc -- Background 0x16
    "11111000", -- 2225 - 0x8b1  :  248 - 0xf8
    "11110000", -- 2226 - 0x8b2  :  240 - 0xf0
    "11100000", -- 2227 - 0x8b3  :  224 - 0xe0
    "01100000", -- 2228 - 0x8b4  :   96 - 0x60
    "11110000", -- 2229 - 0x8b5  :  240 - 0xf0
    "00011100", -- 2230 - 0x8b6  :   28 - 0x1c
    "00000010", -- 2231 - 0x8b7  :    2 - 0x2
    "10000000", -- 2232 - 0x8b8  :  128 - 0x80 -- Background 0x17
    "10000000", -- 2233 - 0x8b9  :  128 - 0x80
    "10000000", -- 2234 - 0x8ba  :  128 - 0x80
    "10000011", -- 2235 - 0x8bb  :  131 - 0x83
    "01001111", -- 2236 - 0x8bc  :   79 - 0x4f
    "00110010", -- 2237 - 0x8bd  :   50 - 0x32
    "00000010", -- 2238 - 0x8be  :    2 - 0x2
    "00000011", -- 2239 - 0x8bf  :    3 - 0x3
    "00000010", -- 2240 - 0x8c0  :    2 - 0x2 -- Background 0x18
    "00000001", -- 2241 - 0x8c1  :    1 - 0x1
    "00000010", -- 2242 - 0x8c2  :    2 - 0x2
    "11111100", -- 2243 - 0x8c3  :  252 - 0xfc
    "11000000", -- 2244 - 0x8c4  :  192 - 0xc0
    "01000000", -- 2245 - 0x8c5  :   64 - 0x40
    "00100000", -- 2246 - 0x8c6  :   32 - 0x20
    "11100000", -- 2247 - 0x8c7  :  224 - 0xe0
    "00001011", -- 2248 - 0x8c8  :   11 - 0xb -- Background 0x19
    "00001011", -- 2249 - 0x8c9  :   11 - 0xb
    "00001111", -- 2250 - 0x8ca  :   15 - 0xf
    "00001001", -- 2251 - 0x8cb  :    9 - 0x9
    "00001000", -- 2252 - 0x8cc  :    8 - 0x8
    "00001001", -- 2253 - 0x8cd  :    9 - 0x9
    "00001111", -- 2254 - 0x8ce  :   15 - 0xf
    "00110000", -- 2255 - 0x8cf  :   48 - 0x30
    "11111000", -- 2256 - 0x8d0  :  248 - 0xf8 -- Background 0x1a
    "11110000", -- 2257 - 0x8d1  :  240 - 0xf0
    "11100000", -- 2258 - 0x8d2  :  224 - 0xe0
    "11000000", -- 2259 - 0x8d3  :  192 - 0xc0
    "11000000", -- 2260 - 0x8d4  :  192 - 0xc0
    "11000000", -- 2261 - 0x8d5  :  192 - 0xc0
    "11111000", -- 2262 - 0x8d6  :  248 - 0xf8
    "00011111", -- 2263 - 0x8d7  :   31 - 0x1f
    "01000000", -- 2264 - 0x8d8  :   64 - 0x40 -- Background 0x1b
    "01000000", -- 2265 - 0x8d9  :   64 - 0x40
    "10000000", -- 2266 - 0x8da  :  128 - 0x80
    "10000000", -- 2267 - 0x8db  :  128 - 0x80
    "01000000", -- 2268 - 0x8dc  :   64 - 0x40
    "00111111", -- 2269 - 0x8dd  :   63 - 0x3f
    "00000100", -- 2270 - 0x8de  :    4 - 0x4
    "00000111", -- 2271 - 0x8df  :    7 - 0x7
    "00000000", -- 2272 - 0x8e0  :    0 - 0x0 -- Background 0x1c
    "00000000", -- 2273 - 0x8e1  :    0 - 0x0
    "00000000", -- 2274 - 0x8e2  :    0 - 0x0
    "00000000", -- 2275 - 0x8e3  :    0 - 0x0
    "00000000", -- 2276 - 0x8e4  :    0 - 0x0
    "11111111", -- 2277 - 0x8e5  :  255 - 0xff
    "01000000", -- 2278 - 0x8e6  :   64 - 0x40
    "11000000", -- 2279 - 0x8e7  :  192 - 0xc0
    "11000000", -- 2280 - 0x8e8  :  192 - 0xc0 -- Background 0x1d
    "00100000", -- 2281 - 0x8e9  :   32 - 0x20
    "00100000", -- 2282 - 0x8ea  :   32 - 0x20
    "00100000", -- 2283 - 0x8eb  :   32 - 0x20
    "01000000", -- 2284 - 0x8ec  :   64 - 0x40
    "10000000", -- 2285 - 0x8ed  :  128 - 0x80
    "00000000", -- 2286 - 0x8ee  :    0 - 0x0
    "00000000", -- 2287 - 0x8ef  :    0 - 0x0
    "01111111", -- 2288 - 0x8f0  :  127 - 0x7f -- Background 0x1e
    "01100010", -- 2289 - 0x8f1  :   98 - 0x62
    "11000100", -- 2290 - 0x8f2  :  196 - 0xc4
    "00011000", -- 2291 - 0x8f3  :   24 - 0x18
    "00111100", -- 2292 - 0x8f4  :   60 - 0x3c
    "11111110", -- 2293 - 0x8f5  :  254 - 0xfe
    "11111110", -- 2294 - 0x8f6  :  254 - 0xfe
    "11111110", -- 2295 - 0x8f7  :  254 - 0xfe
    "00000000", -- 2296 - 0x8f8  :    0 - 0x0 -- Background 0x1f
    "00111000", -- 2297 - 0x8f9  :   56 - 0x38
    "11000110", -- 2298 - 0x8fa  :  198 - 0xc6
    "11001011", -- 2299 - 0x8fb  :  203 - 0xcb
    "11011100", -- 2300 - 0x8fc  :  220 - 0xdc
    "00111010", -- 2301 - 0x8fd  :   58 - 0x3a
    "10011010", -- 2302 - 0x8fe  :  154 - 0x9a
    "11100001", -- 2303 - 0x8ff  :  225 - 0xe1
    "00000000", -- 2304 - 0x900  :    0 - 0x0 -- Background 0x20
    "00011100", -- 2305 - 0x901  :   28 - 0x1c
    "00010011", -- 2306 - 0x902  :   19 - 0x13
    "00001000", -- 2307 - 0x903  :    8 - 0x8
    "00010000", -- 2308 - 0x904  :   16 - 0x10
    "00001000", -- 2309 - 0x905  :    8 - 0x8
    "00010000", -- 2310 - 0x906  :   16 - 0x10
    "00010000", -- 2311 - 0x907  :   16 - 0x10
    "00000000", -- 2312 - 0x908  :    0 - 0x0 -- Background 0x21
    "00111000", -- 2313 - 0x909  :   56 - 0x38
    "11001000", -- 2314 - 0x90a  :  200 - 0xc8
    "00010000", -- 2315 - 0x90b  :   16 - 0x10
    "00001000", -- 2316 - 0x90c  :    8 - 0x8
    "00010000", -- 2317 - 0x90d  :   16 - 0x10
    "00001000", -- 2318 - 0x90e  :    8 - 0x8
    "00001000", -- 2319 - 0x90f  :    8 - 0x8
    "00001000", -- 2320 - 0x910  :    8 - 0x8 -- Background 0x22
    "00011100", -- 2321 - 0x911  :   28 - 0x1c
    "00100111", -- 2322 - 0x912  :   39 - 0x27
    "00101111", -- 2323 - 0x913  :   47 - 0x2f
    "00011111", -- 2324 - 0x914  :   31 - 0x1f
    "00001111", -- 2325 - 0x915  :   15 - 0xf
    "00001111", -- 2326 - 0x916  :   15 - 0xf
    "00001111", -- 2327 - 0x917  :   15 - 0xf
    "00010000", -- 2328 - 0x918  :   16 - 0x10 -- Background 0x23
    "00111100", -- 2329 - 0x919  :   60 - 0x3c
    "11000010", -- 2330 - 0x91a  :  194 - 0xc2
    "10000010", -- 2331 - 0x91b  :  130 - 0x82
    "10000010", -- 2332 - 0x91c  :  130 - 0x82
    "10000010", -- 2333 - 0x91d  :  130 - 0x82
    "00010010", -- 2334 - 0x91e  :   18 - 0x12
    "00011100", -- 2335 - 0x91f  :   28 - 0x1c
    "00001111", -- 2336 - 0x920  :   15 - 0xf -- Background 0x24
    "00001110", -- 2337 - 0x921  :   14 - 0xe
    "00010100", -- 2338 - 0x922  :   20 - 0x14
    "00010100", -- 2339 - 0x923  :   20 - 0x14
    "00010010", -- 2340 - 0x924  :   18 - 0x12
    "00100101", -- 2341 - 0x925  :   37 - 0x25
    "01000100", -- 2342 - 0x926  :   68 - 0x44
    "00111000", -- 2343 - 0x927  :   56 - 0x38
    "00010000", -- 2344 - 0x928  :   16 - 0x10 -- Background 0x25
    "00010000", -- 2345 - 0x929  :   16 - 0x10
    "00010000", -- 2346 - 0x92a  :   16 - 0x10
    "00101100", -- 2347 - 0x92b  :   44 - 0x2c
    "01000100", -- 2348 - 0x92c  :   68 - 0x44
    "11000100", -- 2349 - 0x92d  :  196 - 0xc4
    "00111000", -- 2350 - 0x92e  :   56 - 0x38
    "00000000", -- 2351 - 0x92f  :    0 - 0x0
    "00000000", -- 2352 - 0x930  :    0 - 0x0 -- Background 0x26
    "00000000", -- 2353 - 0x931  :    0 - 0x0
    "00000000", -- 2354 - 0x932  :    0 - 0x0
    "00000000", -- 2355 - 0x933  :    0 - 0x0
    "00000000", -- 2356 - 0x934  :    0 - 0x0
    "00000000", -- 2357 - 0x935  :    0 - 0x0
    "00000000", -- 2358 - 0x936  :    0 - 0x0
    "00000000", -- 2359 - 0x937  :    0 - 0x0
    "00000000", -- 2360 - 0x938  :    0 - 0x0 -- Background 0x27
    "00000000", -- 2361 - 0x939  :    0 - 0x0
    "00000000", -- 2362 - 0x93a  :    0 - 0x0
    "00000000", -- 2363 - 0x93b  :    0 - 0x0
    "00000000", -- 2364 - 0x93c  :    0 - 0x0
    "00000000", -- 2365 - 0x93d  :    0 - 0x0
    "00000000", -- 2366 - 0x93e  :    0 - 0x0
    "00000000", -- 2367 - 0x93f  :    0 - 0x0
    "00000000", -- 2368 - 0x940  :    0 - 0x0 -- Background 0x28
    "00000000", -- 2369 - 0x941  :    0 - 0x0
    "00000000", -- 2370 - 0x942  :    0 - 0x0
    "00000000", -- 2371 - 0x943  :    0 - 0x0
    "00000000", -- 2372 - 0x944  :    0 - 0x0
    "00000000", -- 2373 - 0x945  :    0 - 0x0
    "00000000", -- 2374 - 0x946  :    0 - 0x0
    "00000000", -- 2375 - 0x947  :    0 - 0x0
    "00100000", -- 2376 - 0x948  :   32 - 0x20 -- Background 0x29
    "00100000", -- 2377 - 0x949  :   32 - 0x20
    "00100000", -- 2378 - 0x94a  :   32 - 0x20
    "00100000", -- 2379 - 0x94b  :   32 - 0x20
    "00010011", -- 2380 - 0x94c  :   19 - 0x13
    "00001101", -- 2381 - 0x94d  :   13 - 0xd
    "00000010", -- 2382 - 0x94e  :    2 - 0x2
    "00000001", -- 2383 - 0x94f  :    1 - 0x1
    "00100000", -- 2384 - 0x950  :   32 - 0x20 -- Background 0x2a
    "00100000", -- 2385 - 0x951  :   32 - 0x20
    "00100000", -- 2386 - 0x952  :   32 - 0x20
    "00100000", -- 2387 - 0x953  :   32 - 0x20
    "00010011", -- 2388 - 0x954  :   19 - 0x13
    "00001101", -- 2389 - 0x955  :   13 - 0xd
    "00000001", -- 2390 - 0x956  :    1 - 0x1
    "00000001", -- 2391 - 0x957  :    1 - 0x1
    "00000000", -- 2392 - 0x958  :    0 - 0x0 -- Background 0x2b
    "00000000", -- 2393 - 0x959  :    0 - 0x0
    "00000000", -- 2394 - 0x95a  :    0 - 0x0
    "00000000", -- 2395 - 0x95b  :    0 - 0x0
    "00000000", -- 2396 - 0x95c  :    0 - 0x0
    "00000000", -- 2397 - 0x95d  :    0 - 0x0
    "00000000", -- 2398 - 0x95e  :    0 - 0x0
    "00000000", -- 2399 - 0x95f  :    0 - 0x0
    "00000000", -- 2400 - 0x960  :    0 - 0x0 -- Background 0x2c
    "00000000", -- 2401 - 0x961  :    0 - 0x0
    "00000000", -- 2402 - 0x962  :    0 - 0x0
    "00000000", -- 2403 - 0x963  :    0 - 0x0
    "00000000", -- 2404 - 0x964  :    0 - 0x0
    "00000000", -- 2405 - 0x965  :    0 - 0x0
    "00000000", -- 2406 - 0x966  :    0 - 0x0
    "00000000", -- 2407 - 0x967  :    0 - 0x0
    "00111100", -- 2408 - 0x968  :   60 - 0x3c -- Background 0x2d
    "00000000", -- 2409 - 0x969  :    0 - 0x0
    "10000001", -- 2410 - 0x96a  :  129 - 0x81
    "10011001", -- 2411 - 0x96b  :  153 - 0x99
    "10011001", -- 2412 - 0x96c  :  153 - 0x99
    "10000001", -- 2413 - 0x96d  :  129 - 0x81
    "00000000", -- 2414 - 0x96e  :    0 - 0x0
    "00111100", -- 2415 - 0x96f  :   60 - 0x3c
    "00000000", -- 2416 - 0x970  :    0 - 0x0 -- Background 0x2e
    "00000000", -- 2417 - 0x971  :    0 - 0x0
    "00000000", -- 2418 - 0x972  :    0 - 0x0
    "00000000", -- 2419 - 0x973  :    0 - 0x0
    "00000000", -- 2420 - 0x974  :    0 - 0x0
    "00000000", -- 2421 - 0x975  :    0 - 0x0
    "00000000", -- 2422 - 0x976  :    0 - 0x0
    "00000000", -- 2423 - 0x977  :    0 - 0x0
    "10011111", -- 2424 - 0x978  :  159 - 0x9f -- Background 0x2f
    "10011110", -- 2425 - 0x979  :  158 - 0x9e
    "10011100", -- 2426 - 0x97a  :  156 - 0x9c
    "00011000", -- 2427 - 0x97b  :   24 - 0x18
    "00111000", -- 2428 - 0x97c  :   56 - 0x38
    "11111100", -- 2429 - 0x97d  :  252 - 0xfc
    "11111100", -- 2430 - 0x97e  :  252 - 0xfc
    "11111100", -- 2431 - 0x97f  :  252 - 0xfc
    "01111111", -- 2432 - 0x980  :  127 - 0x7f -- Background 0x30
    "01111110", -- 2433 - 0x981  :  126 - 0x7e
    "11111100", -- 2434 - 0x982  :  252 - 0xfc
    "00111000", -- 2435 - 0x983  :   56 - 0x38
    "00111000", -- 2436 - 0x984  :   56 - 0x38
    "00000100", -- 2437 - 0x985  :    4 - 0x4
    "10000100", -- 2438 - 0x986  :  132 - 0x84
    "11111100", -- 2439 - 0x987  :  252 - 0xfc
    "01111111", -- 2440 - 0x988  :  127 - 0x7f -- Background 0x31
    "01111110", -- 2441 - 0x989  :  126 - 0x7e
    "11111100", -- 2442 - 0x98a  :  252 - 0xfc
    "00111000", -- 2443 - 0x98b  :   56 - 0x38
    "00111000", -- 2444 - 0x98c  :   56 - 0x38
    "00011100", -- 2445 - 0x98d  :   28 - 0x1c
    "10000100", -- 2446 - 0x98e  :  132 - 0x84
    "11000100", -- 2447 - 0x98f  :  196 - 0xc4
    "01111111", -- 2448 - 0x990  :  127 - 0x7f -- Background 0x32
    "01111110", -- 2449 - 0x991  :  126 - 0x7e
    "11111100", -- 2450 - 0x992  :  252 - 0xfc
    "00111000", -- 2451 - 0x993  :   56 - 0x38
    "00100100", -- 2452 - 0x994  :   36 - 0x24
    "00000100", -- 2453 - 0x995  :    4 - 0x4
    "10011100", -- 2454 - 0x996  :  156 - 0x9c
    "11111100", -- 2455 - 0x997  :  252 - 0xfc
    "00100011", -- 2456 - 0x998  :   35 - 0x23 -- Background 0x33
    "00100011", -- 2457 - 0x999  :   35 - 0x23
    "00100001", -- 2458 - 0x99a  :   33 - 0x21
    "00100000", -- 2459 - 0x99b  :   32 - 0x20
    "00010011", -- 2460 - 0x99c  :   19 - 0x13
    "00001101", -- 2461 - 0x99d  :   13 - 0xd
    "00000001", -- 2462 - 0x99e  :    1 - 0x1
    "00000001", -- 2463 - 0x99f  :    1 - 0x1
    "11111100", -- 2464 - 0x9a0  :  252 - 0xfc -- Background 0x34
    "11111100", -- 2465 - 0x9a1  :  252 - 0xfc
    "11111100", -- 2466 - 0x9a2  :  252 - 0xfc
    "11111100", -- 2467 - 0x9a3  :  252 - 0xfc
    "10100100", -- 2468 - 0x9a4  :  164 - 0xa4
    "00100100", -- 2469 - 0x9a5  :   36 - 0x24
    "00010010", -- 2470 - 0x9a6  :   18 - 0x12
    "11101110", -- 2471 - 0x9a7  :  238 - 0xee
    "00100011", -- 2472 - 0x9a8  :   35 - 0x23 -- Background 0x35
    "00100011", -- 2473 - 0x9a9  :   35 - 0x23
    "00100001", -- 2474 - 0x9aa  :   33 - 0x21
    "00100000", -- 2475 - 0x9ab  :   32 - 0x20
    "00010011", -- 2476 - 0x9ac  :   19 - 0x13
    "00001110", -- 2477 - 0x9ad  :   14 - 0xe
    "00000010", -- 2478 - 0x9ae  :    2 - 0x2
    "00000001", -- 2479 - 0x9af  :    1 - 0x1
    "11111100", -- 2480 - 0x9b0  :  252 - 0xfc -- Background 0x36
    "11111100", -- 2481 - 0x9b1  :  252 - 0xfc
    "11111100", -- 2482 - 0x9b2  :  252 - 0xfc
    "11111100", -- 2483 - 0x9b3  :  252 - 0xfc
    "10100110", -- 2484 - 0x9b4  :  166 - 0xa6
    "00110001", -- 2485 - 0x9b5  :   49 - 0x31
    "01001001", -- 2486 - 0x9b6  :   73 - 0x49
    "11000110", -- 2487 - 0x9b7  :  198 - 0xc6
    "11111100", -- 2488 - 0x9b8  :  252 - 0xfc -- Background 0x37
    "11111100", -- 2489 - 0x9b9  :  252 - 0xfc
    "11111100", -- 2490 - 0x9ba  :  252 - 0xfc
    "11111100", -- 2491 - 0x9bb  :  252 - 0xfc
    "10100100", -- 2492 - 0x9bc  :  164 - 0xa4
    "00100100", -- 2493 - 0x9bd  :   36 - 0x24
    "00010010", -- 2494 - 0x9be  :   18 - 0x12
    "11101110", -- 2495 - 0x9bf  :  238 - 0xee
    "00000000", -- 2496 - 0x9c0  :    0 - 0x0 -- Background 0x38
    "00000000", -- 2497 - 0x9c1  :    0 - 0x0
    "00000000", -- 2498 - 0x9c2  :    0 - 0x0
    "00000000", -- 2499 - 0x9c3  :    0 - 0x0
    "00000000", -- 2500 - 0x9c4  :    0 - 0x0
    "00000000", -- 2501 - 0x9c5  :    0 - 0x0
    "00000000", -- 2502 - 0x9c6  :    0 - 0x0
    "00000000", -- 2503 - 0x9c7  :    0 - 0x0
    "00000000", -- 2504 - 0x9c8  :    0 - 0x0 -- Background 0x39
    "00000000", -- 2505 - 0x9c9  :    0 - 0x0
    "00000000", -- 2506 - 0x9ca  :    0 - 0x0
    "00000000", -- 2507 - 0x9cb  :    0 - 0x0
    "00000000", -- 2508 - 0x9cc  :    0 - 0x0
    "00000000", -- 2509 - 0x9cd  :    0 - 0x0
    "00000000", -- 2510 - 0x9ce  :    0 - 0x0
    "00000000", -- 2511 - 0x9cf  :    0 - 0x0
    "00000000", -- 2512 - 0x9d0  :    0 - 0x0 -- Background 0x3a
    "00000000", -- 2513 - 0x9d1  :    0 - 0x0
    "00000000", -- 2514 - 0x9d2  :    0 - 0x0
    "00000000", -- 2515 - 0x9d3  :    0 - 0x0
    "00000000", -- 2516 - 0x9d4  :    0 - 0x0
    "00000000", -- 2517 - 0x9d5  :    0 - 0x0
    "00000000", -- 2518 - 0x9d6  :    0 - 0x0
    "00000000", -- 2519 - 0x9d7  :    0 - 0x0
    "00000000", -- 2520 - 0x9d8  :    0 - 0x0 -- Background 0x3b
    "00000000", -- 2521 - 0x9d9  :    0 - 0x0
    "00000000", -- 2522 - 0x9da  :    0 - 0x0
    "00000000", -- 2523 - 0x9db  :    0 - 0x0
    "00000000", -- 2524 - 0x9dc  :    0 - 0x0
    "00000000", -- 2525 - 0x9dd  :    0 - 0x0
    "00000000", -- 2526 - 0x9de  :    0 - 0x0
    "00000000", -- 2527 - 0x9df  :    0 - 0x0
    "00000000", -- 2528 - 0x9e0  :    0 - 0x0 -- Background 0x3c
    "00000000", -- 2529 - 0x9e1  :    0 - 0x0
    "00000000", -- 2530 - 0x9e2  :    0 - 0x0
    "00000000", -- 2531 - 0x9e3  :    0 - 0x0
    "00000000", -- 2532 - 0x9e4  :    0 - 0x0
    "00000000", -- 2533 - 0x9e5  :    0 - 0x0
    "00000000", -- 2534 - 0x9e6  :    0 - 0x0
    "00000000", -- 2535 - 0x9e7  :    0 - 0x0
    "00000000", -- 2536 - 0x9e8  :    0 - 0x0 -- Background 0x3d
    "00000000", -- 2537 - 0x9e9  :    0 - 0x0
    "00000000", -- 2538 - 0x9ea  :    0 - 0x0
    "00000000", -- 2539 - 0x9eb  :    0 - 0x0
    "00000000", -- 2540 - 0x9ec  :    0 - 0x0
    "00000000", -- 2541 - 0x9ed  :    0 - 0x0
    "00000000", -- 2542 - 0x9ee  :    0 - 0x0
    "00000000", -- 2543 - 0x9ef  :    0 - 0x0
    "00000000", -- 2544 - 0x9f0  :    0 - 0x0 -- Background 0x3e
    "00000000", -- 2545 - 0x9f1  :    0 - 0x0
    "00000000", -- 2546 - 0x9f2  :    0 - 0x0
    "00000000", -- 2547 - 0x9f3  :    0 - 0x0
    "00000000", -- 2548 - 0x9f4  :    0 - 0x0
    "00000000", -- 2549 - 0x9f5  :    0 - 0x0
    "00000000", -- 2550 - 0x9f6  :    0 - 0x0
    "00000000", -- 2551 - 0x9f7  :    0 - 0x0
    "00000000", -- 2552 - 0x9f8  :    0 - 0x0 -- Background 0x3f
    "00000000", -- 2553 - 0x9f9  :    0 - 0x0
    "00000000", -- 2554 - 0x9fa  :    0 - 0x0
    "00000000", -- 2555 - 0x9fb  :    0 - 0x0
    "00000000", -- 2556 - 0x9fc  :    0 - 0x0
    "00000000", -- 2557 - 0x9fd  :    0 - 0x0
    "00000000", -- 2558 - 0x9fe  :    0 - 0x0
    "00000000", -- 2559 - 0x9ff  :    0 - 0x0
    "00000000", -- 2560 - 0xa00  :    0 - 0x0 -- Background 0x40
    "00111110", -- 2561 - 0xa01  :   62 - 0x3e
    "01111111", -- 2562 - 0xa02  :  127 - 0x7f
    "01111111", -- 2563 - 0xa03  :  127 - 0x7f
    "01111111", -- 2564 - 0xa04  :  127 - 0x7f
    "01111111", -- 2565 - 0xa05  :  127 - 0x7f
    "01111111", -- 2566 - 0xa06  :  127 - 0x7f
    "00111110", -- 2567 - 0xa07  :   62 - 0x3e
    "00000000", -- 2568 - 0xa08  :    0 - 0x0 -- Background 0x41
    "00111100", -- 2569 - 0xa09  :   60 - 0x3c
    "00011100", -- 2570 - 0xa0a  :   28 - 0x1c
    "00011100", -- 2571 - 0xa0b  :   28 - 0x1c
    "00011100", -- 2572 - 0xa0c  :   28 - 0x1c
    "00011100", -- 2573 - 0xa0d  :   28 - 0x1c
    "00011100", -- 2574 - 0xa0e  :   28 - 0x1c
    "00011100", -- 2575 - 0xa0f  :   28 - 0x1c
    "00000000", -- 2576 - 0xa10  :    0 - 0x0 -- Background 0x42
    "01111100", -- 2577 - 0xa11  :  124 - 0x7c
    "01111111", -- 2578 - 0xa12  :  127 - 0x7f
    "01100111", -- 2579 - 0xa13  :  103 - 0x67
    "00111111", -- 2580 - 0xa14  :   63 - 0x3f
    "01111110", -- 2581 - 0xa15  :  126 - 0x7e
    "01111111", -- 2582 - 0xa16  :  127 - 0x7f
    "01111111", -- 2583 - 0xa17  :  127 - 0x7f
    "00000000", -- 2584 - 0xa18  :    0 - 0x0 -- Background 0x43
    "01111110", -- 2585 - 0xa19  :  126 - 0x7e
    "01111111", -- 2586 - 0xa1a  :  127 - 0x7f
    "01111111", -- 2587 - 0xa1b  :  127 - 0x7f
    "00011111", -- 2588 - 0xa1c  :   31 - 0x1f
    "01110111", -- 2589 - 0xa1d  :  119 - 0x77
    "01111111", -- 2590 - 0xa1e  :  127 - 0x7f
    "01111110", -- 2591 - 0xa1f  :  126 - 0x7e
    "00000000", -- 2592 - 0xa20  :    0 - 0x0 -- Background 0x44
    "00001110", -- 2593 - 0xa21  :   14 - 0xe
    "00011110", -- 2594 - 0xa22  :   30 - 0x1e
    "00111110", -- 2595 - 0xa23  :   62 - 0x3e
    "01111110", -- 2596 - 0xa24  :  126 - 0x7e
    "01111111", -- 2597 - 0xa25  :  127 - 0x7f
    "01111110", -- 2598 - 0xa26  :  126 - 0x7e
    "00001100", -- 2599 - 0xa27  :   12 - 0xc
    "00000000", -- 2600 - 0xa28  :    0 - 0x0 -- Background 0x45
    "01111111", -- 2601 - 0xa29  :  127 - 0x7f
    "01111111", -- 2602 - 0xa2a  :  127 - 0x7f
    "01111111", -- 2603 - 0xa2b  :  127 - 0x7f
    "01111111", -- 2604 - 0xa2c  :  127 - 0x7f
    "01110111", -- 2605 - 0xa2d  :  119 - 0x77
    "01111111", -- 2606 - 0xa2e  :  127 - 0x7f
    "01111110", -- 2607 - 0xa2f  :  126 - 0x7e
    "00000000", -- 2608 - 0xa30  :    0 - 0x0 -- Background 0x46
    "00111110", -- 2609 - 0xa31  :   62 - 0x3e
    "01111110", -- 2610 - 0xa32  :  126 - 0x7e
    "01111111", -- 2611 - 0xa33  :  127 - 0x7f
    "01111111", -- 2612 - 0xa34  :  127 - 0x7f
    "01110111", -- 2613 - 0xa35  :  119 - 0x77
    "01111111", -- 2614 - 0xa36  :  127 - 0x7f
    "00111110", -- 2615 - 0xa37  :   62 - 0x3e
    "00000000", -- 2616 - 0xa38  :    0 - 0x0 -- Background 0x47
    "01111110", -- 2617 - 0xa39  :  126 - 0x7e
    "01111110", -- 2618 - 0xa3a  :  126 - 0x7e
    "00011110", -- 2619 - 0xa3b  :   30 - 0x1e
    "00011100", -- 2620 - 0xa3c  :   28 - 0x1c
    "00111100", -- 2621 - 0xa3d  :   60 - 0x3c
    "00111000", -- 2622 - 0xa3e  :   56 - 0x38
    "00111000", -- 2623 - 0xa3f  :   56 - 0x38
    "00000000", -- 2624 - 0xa40  :    0 - 0x0 -- Background 0x48
    "00111110", -- 2625 - 0xa41  :   62 - 0x3e
    "01111111", -- 2626 - 0xa42  :  127 - 0x7f
    "01111111", -- 2627 - 0xa43  :  127 - 0x7f
    "01111111", -- 2628 - 0xa44  :  127 - 0x7f
    "01111111", -- 2629 - 0xa45  :  127 - 0x7f
    "01111111", -- 2630 - 0xa46  :  127 - 0x7f
    "00111110", -- 2631 - 0xa47  :   62 - 0x3e
    "00000000", -- 2632 - 0xa48  :    0 - 0x0 -- Background 0x49
    "00111110", -- 2633 - 0xa49  :   62 - 0x3e
    "01111111", -- 2634 - 0xa4a  :  127 - 0x7f
    "01110111", -- 2635 - 0xa4b  :  119 - 0x77
    "01111111", -- 2636 - 0xa4c  :  127 - 0x7f
    "01111111", -- 2637 - 0xa4d  :  127 - 0x7f
    "00111111", -- 2638 - 0xa4e  :   63 - 0x3f
    "00111110", -- 2639 - 0xa4f  :   62 - 0x3e
    "11111111", -- 2640 - 0xa50  :  255 - 0xff -- Background 0x4a
    "10011001", -- 2641 - 0xa51  :  153 - 0x99
    "10011001", -- 2642 - 0xa52  :  153 - 0x99
    "10011001", -- 2643 - 0xa53  :  153 - 0x99
    "10011001", -- 2644 - 0xa54  :  153 - 0x99
    "10011001", -- 2645 - 0xa55  :  153 - 0x99
    "10011001", -- 2646 - 0xa56  :  153 - 0x99
    "11111111", -- 2647 - 0xa57  :  255 - 0xff
    "11110000", -- 2648 - 0xa58  :  240 - 0xf0 -- Background 0x4b
    "10010000", -- 2649 - 0xa59  :  144 - 0x90
    "10010000", -- 2650 - 0xa5a  :  144 - 0x90
    "10010000", -- 2651 - 0xa5b  :  144 - 0x90
    "10010000", -- 2652 - 0xa5c  :  144 - 0x90
    "10010000", -- 2653 - 0xa5d  :  144 - 0x90
    "10010000", -- 2654 - 0xa5e  :  144 - 0x90
    "11110000", -- 2655 - 0xa5f  :  240 - 0xf0
    "11111111", -- 2656 - 0xa60  :  255 - 0xff -- Background 0x4c
    "11111111", -- 2657 - 0xa61  :  255 - 0xff
    "11111111", -- 2658 - 0xa62  :  255 - 0xff
    "11111111", -- 2659 - 0xa63  :  255 - 0xff
    "11111111", -- 2660 - 0xa64  :  255 - 0xff
    "11111111", -- 2661 - 0xa65  :  255 - 0xff
    "11111111", -- 2662 - 0xa66  :  255 - 0xff
    "11111111", -- 2663 - 0xa67  :  255 - 0xff
    "11111111", -- 2664 - 0xa68  :  255 - 0xff -- Background 0x4d
    "11111111", -- 2665 - 0xa69  :  255 - 0xff
    "11111111", -- 2666 - 0xa6a  :  255 - 0xff
    "11111111", -- 2667 - 0xa6b  :  255 - 0xff
    "11111111", -- 2668 - 0xa6c  :  255 - 0xff
    "11111111", -- 2669 - 0xa6d  :  255 - 0xff
    "11111111", -- 2670 - 0xa6e  :  255 - 0xff
    "11111111", -- 2671 - 0xa6f  :  255 - 0xff
    "11111111", -- 2672 - 0xa70  :  255 - 0xff -- Background 0x4e
    "11111111", -- 2673 - 0xa71  :  255 - 0xff
    "11111111", -- 2674 - 0xa72  :  255 - 0xff
    "11111111", -- 2675 - 0xa73  :  255 - 0xff
    "11111111", -- 2676 - 0xa74  :  255 - 0xff
    "11111111", -- 2677 - 0xa75  :  255 - 0xff
    "11111111", -- 2678 - 0xa76  :  255 - 0xff
    "11111111", -- 2679 - 0xa77  :  255 - 0xff
    "11111111", -- 2680 - 0xa78  :  255 - 0xff -- Background 0x4f
    "11111111", -- 2681 - 0xa79  :  255 - 0xff
    "11111111", -- 2682 - 0xa7a  :  255 - 0xff
    "11111111", -- 2683 - 0xa7b  :  255 - 0xff
    "11111111", -- 2684 - 0xa7c  :  255 - 0xff
    "11111111", -- 2685 - 0xa7d  :  255 - 0xff
    "11111111", -- 2686 - 0xa7e  :  255 - 0xff
    "11111111", -- 2687 - 0xa7f  :  255 - 0xff
    "00010000", -- 2688 - 0xa80  :   16 - 0x10 -- Background 0x50
    "00101000", -- 2689 - 0xa81  :   40 - 0x28
    "11101110", -- 2690 - 0xa82  :  238 - 0xee
    "10000010", -- 2691 - 0xa83  :  130 - 0x82
    "01000100", -- 2692 - 0xa84  :   68 - 0x44
    "01000100", -- 2693 - 0xa85  :   68 - 0x44
    "10010010", -- 2694 - 0xa86  :  146 - 0x92
    "11101110", -- 2695 - 0xa87  :  238 - 0xee
    "00010000", -- 2696 - 0xa88  :   16 - 0x10 -- Background 0x51
    "00101000", -- 2697 - 0xa89  :   40 - 0x28
    "11101110", -- 2698 - 0xa8a  :  238 - 0xee
    "10000010", -- 2699 - 0xa8b  :  130 - 0x82
    "01000100", -- 2700 - 0xa8c  :   68 - 0x44
    "01000100", -- 2701 - 0xa8d  :   68 - 0x44
    "10010010", -- 2702 - 0xa8e  :  146 - 0x92
    "11101110", -- 2703 - 0xa8f  :  238 - 0xee
    "00010000", -- 2704 - 0xa90  :   16 - 0x10 -- Background 0x52
    "00111000", -- 2705 - 0xa91  :   56 - 0x38
    "11111110", -- 2706 - 0xa92  :  254 - 0xfe
    "11111110", -- 2707 - 0xa93  :  254 - 0xfe
    "01111100", -- 2708 - 0xa94  :  124 - 0x7c
    "01111100", -- 2709 - 0xa95  :  124 - 0x7c
    "11111110", -- 2710 - 0xa96  :  254 - 0xfe
    "11101110", -- 2711 - 0xa97  :  238 - 0xee
    "11111111", -- 2712 - 0xa98  :  255 - 0xff -- Background 0x53
    "11111111", -- 2713 - 0xa99  :  255 - 0xff
    "11111111", -- 2714 - 0xa9a  :  255 - 0xff
    "11111111", -- 2715 - 0xa9b  :  255 - 0xff
    "11111111", -- 2716 - 0xa9c  :  255 - 0xff
    "11111111", -- 2717 - 0xa9d  :  255 - 0xff
    "11111111", -- 2718 - 0xa9e  :  255 - 0xff
    "11111111", -- 2719 - 0xa9f  :  255 - 0xff
    "00000000", -- 2720 - 0xaa0  :    0 - 0x0 -- Background 0x54
    "00000000", -- 2721 - 0xaa1  :    0 - 0x0
    "00000000", -- 2722 - 0xaa2  :    0 - 0x0
    "00000000", -- 2723 - 0xaa3  :    0 - 0x0
    "00000000", -- 2724 - 0xaa4  :    0 - 0x0
    "00000000", -- 2725 - 0xaa5  :    0 - 0x0
    "00000000", -- 2726 - 0xaa6  :    0 - 0x0
    "00000000", -- 2727 - 0xaa7  :    0 - 0x0
    "11111111", -- 2728 - 0xaa8  :  255 - 0xff -- Background 0x55
    "11111111", -- 2729 - 0xaa9  :  255 - 0xff
    "11111111", -- 2730 - 0xaaa  :  255 - 0xff
    "11111111", -- 2731 - 0xaab  :  255 - 0xff
    "11111111", -- 2732 - 0xaac  :  255 - 0xff
    "11111111", -- 2733 - 0xaad  :  255 - 0xff
    "11111111", -- 2734 - 0xaae  :  255 - 0xff
    "11111111", -- 2735 - 0xaaf  :  255 - 0xff
    "00101010", -- 2736 - 0xab0  :   42 - 0x2a -- Background 0x56
    "01000101", -- 2737 - 0xab1  :   69 - 0x45
    "00001000", -- 2738 - 0xab2  :    8 - 0x8
    "00010101", -- 2739 - 0xab3  :   21 - 0x15
    "00100000", -- 2740 - 0xab4  :   32 - 0x20
    "01000101", -- 2741 - 0xab5  :   69 - 0x45
    "10101000", -- 2742 - 0xab6  :  168 - 0xa8
    "00000000", -- 2743 - 0xab7  :    0 - 0x0
    "00001000", -- 2744 - 0xab8  :    8 - 0x8 -- Background 0x57
    "01010101", -- 2745 - 0xab9  :   85 - 0x55
    "10100000", -- 2746 - 0xaba  :  160 - 0xa0
    "00010000", -- 2747 - 0xabb  :   16 - 0x10
    "10000000", -- 2748 - 0xabc  :  128 - 0x80
    "00010100", -- 2749 - 0xabd  :   20 - 0x14
    "00100010", -- 2750 - 0xabe  :   34 - 0x22
    "00000000", -- 2751 - 0xabf  :    0 - 0x0
    "11111111", -- 2752 - 0xac0  :  255 - 0xff -- Background 0x58
    "11010101", -- 2753 - 0xac1  :  213 - 0xd5
    "10100000", -- 2754 - 0xac2  :  160 - 0xa0
    "11010000", -- 2755 - 0xac3  :  208 - 0xd0
    "10001111", -- 2756 - 0xac4  :  143 - 0x8f
    "11001000", -- 2757 - 0xac5  :  200 - 0xc8
    "10001000", -- 2758 - 0xac6  :  136 - 0x88
    "11001000", -- 2759 - 0xac7  :  200 - 0xc8
    "10001000", -- 2760 - 0xac8  :  136 - 0x88 -- Background 0x59
    "11001000", -- 2761 - 0xac9  :  200 - 0xc8
    "10001000", -- 2762 - 0xaca  :  136 - 0x88
    "11001111", -- 2763 - 0xacb  :  207 - 0xcf
    "10010000", -- 2764 - 0xacc  :  144 - 0x90
    "11100000", -- 2765 - 0xacd  :  224 - 0xe0
    "11101010", -- 2766 - 0xace  :  234 - 0xea
    "11111111", -- 2767 - 0xacf  :  255 - 0xff
    "11111111", -- 2768 - 0xad0  :  255 - 0xff -- Background 0x5a
    "01011011", -- 2769 - 0xad1  :   91 - 0x5b
    "00000111", -- 2770 - 0xad2  :    7 - 0x7
    "00001001", -- 2771 - 0xad3  :    9 - 0x9
    "11110011", -- 2772 - 0xad4  :  243 - 0xf3
    "00010001", -- 2773 - 0xad5  :   17 - 0x11
    "00010011", -- 2774 - 0xad6  :   19 - 0x13
    "00010001", -- 2775 - 0xad7  :   17 - 0x11
    "00010011", -- 2776 - 0xad8  :   19 - 0x13 -- Background 0x5b
    "00010001", -- 2777 - 0xad9  :   17 - 0x11
    "00010011", -- 2778 - 0xada  :   19 - 0x13
    "11110001", -- 2779 - 0xadb  :  241 - 0xf1
    "00001011", -- 2780 - 0xadc  :   11 - 0xb
    "00000101", -- 2781 - 0xadd  :    5 - 0x5
    "10101011", -- 2782 - 0xade  :  171 - 0xab
    "11111111", -- 2783 - 0xadf  :  255 - 0xff
    "00011100", -- 2784 - 0xae0  :   28 - 0x1c -- Background 0x5c
    "00100010", -- 2785 - 0xae1  :   34 - 0x22
    "01000001", -- 2786 - 0xae2  :   65 - 0x41
    "01000001", -- 2787 - 0xae3  :   65 - 0x41
    "01000001", -- 2788 - 0xae4  :   65 - 0x41
    "00100010", -- 2789 - 0xae5  :   34 - 0x22
    "00100010", -- 2790 - 0xae6  :   34 - 0x22
    "00011100", -- 2791 - 0xae7  :   28 - 0x1c
    "00001000", -- 2792 - 0xae8  :    8 - 0x8 -- Background 0x5d
    "00010000", -- 2793 - 0xae9  :   16 - 0x10
    "00010000", -- 2794 - 0xaea  :   16 - 0x10
    "00001000", -- 2795 - 0xaeb  :    8 - 0x8
    "00000100", -- 2796 - 0xaec  :    4 - 0x4
    "00000100", -- 2797 - 0xaed  :    4 - 0x4
    "00001000", -- 2798 - 0xaee  :    8 - 0x8
    "00010000", -- 2799 - 0xaef  :   16 - 0x10
    "00110110", -- 2800 - 0xaf0  :   54 - 0x36 -- Background 0x5e
    "01101011", -- 2801 - 0xaf1  :  107 - 0x6b
    "01001001", -- 2802 - 0xaf2  :   73 - 0x49
    "01000001", -- 2803 - 0xaf3  :   65 - 0x41
    "01000001", -- 2804 - 0xaf4  :   65 - 0x41
    "00100010", -- 2805 - 0xaf5  :   34 - 0x22
    "00010100", -- 2806 - 0xaf6  :   20 - 0x14
    "00001000", -- 2807 - 0xaf7  :    8 - 0x8
    "00111110", -- 2808 - 0xaf8  :   62 - 0x3e -- Background 0x5f
    "01101011", -- 2809 - 0xaf9  :  107 - 0x6b
    "00100010", -- 2810 - 0xafa  :   34 - 0x22
    "01100011", -- 2811 - 0xafb  :   99 - 0x63
    "00100010", -- 2812 - 0xafc  :   34 - 0x22
    "01100011", -- 2813 - 0xafd  :   99 - 0x63
    "00100010", -- 2814 - 0xafe  :   34 - 0x22
    "01111111", -- 2815 - 0xaff  :  127 - 0x7f
    "11111111", -- 2816 - 0xb00  :  255 - 0xff -- Background 0x60
    "11111111", -- 2817 - 0xb01  :  255 - 0xff
    "11111111", -- 2818 - 0xb02  :  255 - 0xff
    "11111111", -- 2819 - 0xb03  :  255 - 0xff
    "11010101", -- 2820 - 0xb04  :  213 - 0xd5
    "10101010", -- 2821 - 0xb05  :  170 - 0xaa
    "11010101", -- 2822 - 0xb06  :  213 - 0xd5
    "11111111", -- 2823 - 0xb07  :  255 - 0xff
    "11111111", -- 2824 - 0xb08  :  255 - 0xff -- Background 0x61
    "11111111", -- 2825 - 0xb09  :  255 - 0xff
    "11111111", -- 2826 - 0xb0a  :  255 - 0xff
    "11111111", -- 2827 - 0xb0b  :  255 - 0xff
    "01010101", -- 2828 - 0xb0c  :   85 - 0x55
    "10101010", -- 2829 - 0xb0d  :  170 - 0xaa
    "01010101", -- 2830 - 0xb0e  :   85 - 0x55
    "11111111", -- 2831 - 0xb0f  :  255 - 0xff
    "11111111", -- 2832 - 0xb10  :  255 - 0xff -- Background 0x62
    "11111111", -- 2833 - 0xb11  :  255 - 0xff
    "11111111", -- 2834 - 0xb12  :  255 - 0xff
    "11111111", -- 2835 - 0xb13  :  255 - 0xff
    "01010101", -- 2836 - 0xb14  :   85 - 0x55
    "10101011", -- 2837 - 0xb15  :  171 - 0xab
    "01010101", -- 2838 - 0xb16  :   85 - 0x55
    "11111111", -- 2839 - 0xb17  :  255 - 0xff
    "00000000", -- 2840 - 0xb18  :    0 - 0x0 -- Background 0x63
    "00000000", -- 2841 - 0xb19  :    0 - 0x0
    "00000000", -- 2842 - 0xb1a  :    0 - 0x0
    "00000000", -- 2843 - 0xb1b  :    0 - 0x0
    "00000000", -- 2844 - 0xb1c  :    0 - 0x0
    "00000000", -- 2845 - 0xb1d  :    0 - 0x0
    "00000000", -- 2846 - 0xb1e  :    0 - 0x0
    "00000000", -- 2847 - 0xb1f  :    0 - 0x0
    "00000001", -- 2848 - 0xb20  :    1 - 0x1 -- Background 0x64
    "00000001", -- 2849 - 0xb21  :    1 - 0x1
    "00000011", -- 2850 - 0xb22  :    3 - 0x3
    "00000011", -- 2851 - 0xb23  :    3 - 0x3
    "00000110", -- 2852 - 0xb24  :    6 - 0x6
    "00000110", -- 2853 - 0xb25  :    6 - 0x6
    "00001100", -- 2854 - 0xb26  :   12 - 0xc
    "00001100", -- 2855 - 0xb27  :   12 - 0xc
    "00011000", -- 2856 - 0xb28  :   24 - 0x18 -- Background 0x65
    "00011000", -- 2857 - 0xb29  :   24 - 0x18
    "00110000", -- 2858 - 0xb2a  :   48 - 0x30
    "00110000", -- 2859 - 0xb2b  :   48 - 0x30
    "01100000", -- 2860 - 0xb2c  :   96 - 0x60
    "01100000", -- 2861 - 0xb2d  :   96 - 0x60
    "11101010", -- 2862 - 0xb2e  :  234 - 0xea
    "11111111", -- 2863 - 0xb2f  :  255 - 0xff
    "10000000", -- 2864 - 0xb30  :  128 - 0x80 -- Background 0x66
    "10000000", -- 2865 - 0xb31  :  128 - 0x80
    "11000000", -- 2866 - 0xb32  :  192 - 0xc0
    "01000000", -- 2867 - 0xb33  :   64 - 0x40
    "10100000", -- 2868 - 0xb34  :  160 - 0xa0
    "01100000", -- 2869 - 0xb35  :   96 - 0x60
    "00110000", -- 2870 - 0xb36  :   48 - 0x30
    "00010000", -- 2871 - 0xb37  :   16 - 0x10
    "00101000", -- 2872 - 0xb38  :   40 - 0x28 -- Background 0x67
    "00011000", -- 2873 - 0xb39  :   24 - 0x18
    "00001100", -- 2874 - 0xb3a  :   12 - 0xc
    "00010100", -- 2875 - 0xb3b  :   20 - 0x14
    "00001010", -- 2876 - 0xb3c  :   10 - 0xa
    "00000110", -- 2877 - 0xb3d  :    6 - 0x6
    "10101011", -- 2878 - 0xb3e  :  171 - 0xab
    "11111111", -- 2879 - 0xb3f  :  255 - 0xff
    "00000000", -- 2880 - 0xb40  :    0 - 0x0 -- Background 0x68
    "00000000", -- 2881 - 0xb41  :    0 - 0x0
    "00000000", -- 2882 - 0xb42  :    0 - 0x0
    "00000000", -- 2883 - 0xb43  :    0 - 0x0
    "00000000", -- 2884 - 0xb44  :    0 - 0x0
    "00000000", -- 2885 - 0xb45  :    0 - 0x0
    "00000000", -- 2886 - 0xb46  :    0 - 0x0
    "00000000", -- 2887 - 0xb47  :    0 - 0x0
    "00000000", -- 2888 - 0xb48  :    0 - 0x0 -- Background 0x69
    "00000000", -- 2889 - 0xb49  :    0 - 0x0
    "00000000", -- 2890 - 0xb4a  :    0 - 0x0
    "00000000", -- 2891 - 0xb4b  :    0 - 0x0
    "00000000", -- 2892 - 0xb4c  :    0 - 0x0
    "00000000", -- 2893 - 0xb4d  :    0 - 0x0
    "00000000", -- 2894 - 0xb4e  :    0 - 0x0
    "00000000", -- 2895 - 0xb4f  :    0 - 0x0
    "00000000", -- 2896 - 0xb50  :    0 - 0x0 -- Background 0x6a
    "00000000", -- 2897 - 0xb51  :    0 - 0x0
    "00000000", -- 2898 - 0xb52  :    0 - 0x0
    "00000000", -- 2899 - 0xb53  :    0 - 0x0
    "00000000", -- 2900 - 0xb54  :    0 - 0x0
    "00000000", -- 2901 - 0xb55  :    0 - 0x0
    "00000000", -- 2902 - 0xb56  :    0 - 0x0
    "00000000", -- 2903 - 0xb57  :    0 - 0x0
    "00000000", -- 2904 - 0xb58  :    0 - 0x0 -- Background 0x6b
    "00000000", -- 2905 - 0xb59  :    0 - 0x0
    "00000000", -- 2906 - 0xb5a  :    0 - 0x0
    "00000000", -- 2907 - 0xb5b  :    0 - 0x0
    "00000000", -- 2908 - 0xb5c  :    0 - 0x0
    "00000000", -- 2909 - 0xb5d  :    0 - 0x0
    "00000000", -- 2910 - 0xb5e  :    0 - 0x0
    "00000000", -- 2911 - 0xb5f  :    0 - 0x0
    "00000000", -- 2912 - 0xb60  :    0 - 0x0 -- Background 0x6c
    "00000000", -- 2913 - 0xb61  :    0 - 0x0
    "00000000", -- 2914 - 0xb62  :    0 - 0x0
    "00000000", -- 2915 - 0xb63  :    0 - 0x0
    "00000000", -- 2916 - 0xb64  :    0 - 0x0
    "00000000", -- 2917 - 0xb65  :    0 - 0x0
    "00000000", -- 2918 - 0xb66  :    0 - 0x0
    "00000000", -- 2919 - 0xb67  :    0 - 0x0
    "00000000", -- 2920 - 0xb68  :    0 - 0x0 -- Background 0x6d
    "00000000", -- 2921 - 0xb69  :    0 - 0x0
    "00000000", -- 2922 - 0xb6a  :    0 - 0x0
    "00000000", -- 2923 - 0xb6b  :    0 - 0x0
    "00000000", -- 2924 - 0xb6c  :    0 - 0x0
    "00000000", -- 2925 - 0xb6d  :    0 - 0x0
    "00000000", -- 2926 - 0xb6e  :    0 - 0x0
    "00000000", -- 2927 - 0xb6f  :    0 - 0x0
    "00000000", -- 2928 - 0xb70  :    0 - 0x0 -- Background 0x6e
    "00000000", -- 2929 - 0xb71  :    0 - 0x0
    "00000000", -- 2930 - 0xb72  :    0 - 0x0
    "00000000", -- 2931 - 0xb73  :    0 - 0x0
    "00000000", -- 2932 - 0xb74  :    0 - 0x0
    "00000000", -- 2933 - 0xb75  :    0 - 0x0
    "00000000", -- 2934 - 0xb76  :    0 - 0x0
    "00000000", -- 2935 - 0xb77  :    0 - 0x0
    "00000000", -- 2936 - 0xb78  :    0 - 0x0 -- Background 0x6f
    "00000000", -- 2937 - 0xb79  :    0 - 0x0
    "00000000", -- 2938 - 0xb7a  :    0 - 0x0
    "00000000", -- 2939 - 0xb7b  :    0 - 0x0
    "00000000", -- 2940 - 0xb7c  :    0 - 0x0
    "00000000", -- 2941 - 0xb7d  :    0 - 0x0
    "00000000", -- 2942 - 0xb7e  :    0 - 0x0
    "00000000", -- 2943 - 0xb7f  :    0 - 0x0
    "00000000", -- 2944 - 0xb80  :    0 - 0x0 -- Background 0x70
    "00000000", -- 2945 - 0xb81  :    0 - 0x0
    "00000000", -- 2946 - 0xb82  :    0 - 0x0
    "00000000", -- 2947 - 0xb83  :    0 - 0x0
    "00000000", -- 2948 - 0xb84  :    0 - 0x0
    "00000000", -- 2949 - 0xb85  :    0 - 0x0
    "00000000", -- 2950 - 0xb86  :    0 - 0x0
    "00000000", -- 2951 - 0xb87  :    0 - 0x0
    "00000000", -- 2952 - 0xb88  :    0 - 0x0 -- Background 0x71
    "00000000", -- 2953 - 0xb89  :    0 - 0x0
    "00000000", -- 2954 - 0xb8a  :    0 - 0x0
    "00000000", -- 2955 - 0xb8b  :    0 - 0x0
    "00000000", -- 2956 - 0xb8c  :    0 - 0x0
    "00000000", -- 2957 - 0xb8d  :    0 - 0x0
    "00000000", -- 2958 - 0xb8e  :    0 - 0x0
    "00000000", -- 2959 - 0xb8f  :    0 - 0x0
    "00000000", -- 2960 - 0xb90  :    0 - 0x0 -- Background 0x72
    "00000000", -- 2961 - 0xb91  :    0 - 0x0
    "00000000", -- 2962 - 0xb92  :    0 - 0x0
    "00000000", -- 2963 - 0xb93  :    0 - 0x0
    "00000000", -- 2964 - 0xb94  :    0 - 0x0
    "00000000", -- 2965 - 0xb95  :    0 - 0x0
    "00000000", -- 2966 - 0xb96  :    0 - 0x0
    "00000000", -- 2967 - 0xb97  :    0 - 0x0
    "00000000", -- 2968 - 0xb98  :    0 - 0x0 -- Background 0x73
    "00000000", -- 2969 - 0xb99  :    0 - 0x0
    "00000000", -- 2970 - 0xb9a  :    0 - 0x0
    "00000000", -- 2971 - 0xb9b  :    0 - 0x0
    "00000000", -- 2972 - 0xb9c  :    0 - 0x0
    "00000000", -- 2973 - 0xb9d  :    0 - 0x0
    "00000000", -- 2974 - 0xb9e  :    0 - 0x0
    "00000000", -- 2975 - 0xb9f  :    0 - 0x0
    "00000000", -- 2976 - 0xba0  :    0 - 0x0 -- Background 0x74
    "00000000", -- 2977 - 0xba1  :    0 - 0x0
    "00000000", -- 2978 - 0xba2  :    0 - 0x0
    "00000000", -- 2979 - 0xba3  :    0 - 0x0
    "00000000", -- 2980 - 0xba4  :    0 - 0x0
    "00000000", -- 2981 - 0xba5  :    0 - 0x0
    "00000000", -- 2982 - 0xba6  :    0 - 0x0
    "00000000", -- 2983 - 0xba7  :    0 - 0x0
    "00000000", -- 2984 - 0xba8  :    0 - 0x0 -- Background 0x75
    "00000000", -- 2985 - 0xba9  :    0 - 0x0
    "00000000", -- 2986 - 0xbaa  :    0 - 0x0
    "00000000", -- 2987 - 0xbab  :    0 - 0x0
    "00000000", -- 2988 - 0xbac  :    0 - 0x0
    "00000000", -- 2989 - 0xbad  :    0 - 0x0
    "00000000", -- 2990 - 0xbae  :    0 - 0x0
    "00000000", -- 2991 - 0xbaf  :    0 - 0x0
    "00000000", -- 2992 - 0xbb0  :    0 - 0x0 -- Background 0x76
    "00000000", -- 2993 - 0xbb1  :    0 - 0x0
    "00000000", -- 2994 - 0xbb2  :    0 - 0x0
    "00000000", -- 2995 - 0xbb3  :    0 - 0x0
    "00000000", -- 2996 - 0xbb4  :    0 - 0x0
    "00000000", -- 2997 - 0xbb5  :    0 - 0x0
    "00000000", -- 2998 - 0xbb6  :    0 - 0x0
    "00000000", -- 2999 - 0xbb7  :    0 - 0x0
    "00000000", -- 3000 - 0xbb8  :    0 - 0x0 -- Background 0x77
    "00000000", -- 3001 - 0xbb9  :    0 - 0x0
    "00000000", -- 3002 - 0xbba  :    0 - 0x0
    "00000000", -- 3003 - 0xbbb  :    0 - 0x0
    "00000000", -- 3004 - 0xbbc  :    0 - 0x0
    "00000000", -- 3005 - 0xbbd  :    0 - 0x0
    "00000000", -- 3006 - 0xbbe  :    0 - 0x0
    "00000000", -- 3007 - 0xbbf  :    0 - 0x0
    "00000000", -- 3008 - 0xbc0  :    0 - 0x0 -- Background 0x78
    "00000000", -- 3009 - 0xbc1  :    0 - 0x0
    "00000000", -- 3010 - 0xbc2  :    0 - 0x0
    "00000000", -- 3011 - 0xbc3  :    0 - 0x0
    "00000000", -- 3012 - 0xbc4  :    0 - 0x0
    "00000000", -- 3013 - 0xbc5  :    0 - 0x0
    "00000000", -- 3014 - 0xbc6  :    0 - 0x0
    "00000000", -- 3015 - 0xbc7  :    0 - 0x0
    "00000000", -- 3016 - 0xbc8  :    0 - 0x0 -- Background 0x79
    "00000000", -- 3017 - 0xbc9  :    0 - 0x0
    "00000000", -- 3018 - 0xbca  :    0 - 0x0
    "00000000", -- 3019 - 0xbcb  :    0 - 0x0
    "00000000", -- 3020 - 0xbcc  :    0 - 0x0
    "00000000", -- 3021 - 0xbcd  :    0 - 0x0
    "00000000", -- 3022 - 0xbce  :    0 - 0x0
    "00000000", -- 3023 - 0xbcf  :    0 - 0x0
    "00000000", -- 3024 - 0xbd0  :    0 - 0x0 -- Background 0x7a
    "00000000", -- 3025 - 0xbd1  :    0 - 0x0
    "00000000", -- 3026 - 0xbd2  :    0 - 0x0
    "00000000", -- 3027 - 0xbd3  :    0 - 0x0
    "00000000", -- 3028 - 0xbd4  :    0 - 0x0
    "00000000", -- 3029 - 0xbd5  :    0 - 0x0
    "00000000", -- 3030 - 0xbd6  :    0 - 0x0
    "00000000", -- 3031 - 0xbd7  :    0 - 0x0
    "00000000", -- 3032 - 0xbd8  :    0 - 0x0 -- Background 0x7b
    "00000000", -- 3033 - 0xbd9  :    0 - 0x0
    "00000000", -- 3034 - 0xbda  :    0 - 0x0
    "00000000", -- 3035 - 0xbdb  :    0 - 0x0
    "00000000", -- 3036 - 0xbdc  :    0 - 0x0
    "00000000", -- 3037 - 0xbdd  :    0 - 0x0
    "00000000", -- 3038 - 0xbde  :    0 - 0x0
    "00000000", -- 3039 - 0xbdf  :    0 - 0x0
    "00000000", -- 3040 - 0xbe0  :    0 - 0x0 -- Background 0x7c
    "00000000", -- 3041 - 0xbe1  :    0 - 0x0
    "00000000", -- 3042 - 0xbe2  :    0 - 0x0
    "00000000", -- 3043 - 0xbe3  :    0 - 0x0
    "00000000", -- 3044 - 0xbe4  :    0 - 0x0
    "00000000", -- 3045 - 0xbe5  :    0 - 0x0
    "00000000", -- 3046 - 0xbe6  :    0 - 0x0
    "00000000", -- 3047 - 0xbe7  :    0 - 0x0
    "00000000", -- 3048 - 0xbe8  :    0 - 0x0 -- Background 0x7d
    "00000000", -- 3049 - 0xbe9  :    0 - 0x0
    "00000000", -- 3050 - 0xbea  :    0 - 0x0
    "00000000", -- 3051 - 0xbeb  :    0 - 0x0
    "00000000", -- 3052 - 0xbec  :    0 - 0x0
    "00000000", -- 3053 - 0xbed  :    0 - 0x0
    "00000000", -- 3054 - 0xbee  :    0 - 0x0
    "00000000", -- 3055 - 0xbef  :    0 - 0x0
    "00000000", -- 3056 - 0xbf0  :    0 - 0x0 -- Background 0x7e
    "00000000", -- 3057 - 0xbf1  :    0 - 0x0
    "00000000", -- 3058 - 0xbf2  :    0 - 0x0
    "00000000", -- 3059 - 0xbf3  :    0 - 0x0
    "00000000", -- 3060 - 0xbf4  :    0 - 0x0
    "00000000", -- 3061 - 0xbf5  :    0 - 0x0
    "00000000", -- 3062 - 0xbf6  :    0 - 0x0
    "00000000", -- 3063 - 0xbf7  :    0 - 0x0
    "00000000", -- 3064 - 0xbf8  :    0 - 0x0 -- Background 0x7f
    "00000000", -- 3065 - 0xbf9  :    0 - 0x0
    "00000000", -- 3066 - 0xbfa  :    0 - 0x0
    "00000000", -- 3067 - 0xbfb  :    0 - 0x0
    "00000000", -- 3068 - 0xbfc  :    0 - 0x0
    "00000000", -- 3069 - 0xbfd  :    0 - 0x0
    "00000000", -- 3070 - 0xbfe  :    0 - 0x0
    "00000000", -- 3071 - 0xbff  :    0 - 0x0
    "00000011", -- 3072 - 0xc00  :    3 - 0x3 -- Background 0x80
    "00001111", -- 3073 - 0xc01  :   15 - 0xf
    "00011100", -- 3074 - 0xc02  :   28 - 0x1c
    "00110000", -- 3075 - 0xc03  :   48 - 0x30
    "00100000", -- 3076 - 0xc04  :   32 - 0x20
    "01000000", -- 3077 - 0xc05  :   64 - 0x40
    "01000000", -- 3078 - 0xc06  :   64 - 0x40
    "01111111", -- 3079 - 0xc07  :  127 - 0x7f
    "00000001", -- 3080 - 0xc08  :    1 - 0x1 -- Background 0x81
    "00000001", -- 3081 - 0xc09  :    1 - 0x1
    "00000001", -- 3082 - 0xc0a  :    1 - 0x1
    "00000001", -- 3083 - 0xc0b  :    1 - 0x1
    "00000001", -- 3084 - 0xc0c  :    1 - 0x1
    "00000001", -- 3085 - 0xc0d  :    1 - 0x1
    "00000011", -- 3086 - 0xc0e  :    3 - 0x3
    "00000011", -- 3087 - 0xc0f  :    3 - 0x3
    "11000000", -- 3088 - 0xc10  :  192 - 0xc0 -- Background 0x82
    "11110000", -- 3089 - 0xc11  :  240 - 0xf0
    "00111000", -- 3090 - 0xc12  :   56 - 0x38
    "00001110", -- 3091 - 0xc13  :   14 - 0xe
    "00011110", -- 3092 - 0xc14  :   30 - 0x1e
    "00011110", -- 3093 - 0xc15  :   30 - 0x1e
    "00000010", -- 3094 - 0xc16  :    2 - 0x2
    "11111110", -- 3095 - 0xc17  :  254 - 0xfe
    "10000000", -- 3096 - 0xc18  :  128 - 0x80 -- Background 0x83
    "10000000", -- 3097 - 0xc19  :  128 - 0x80
    "10000000", -- 3098 - 0xc1a  :  128 - 0x80
    "10000000", -- 3099 - 0xc1b  :  128 - 0x80
    "10000000", -- 3100 - 0xc1c  :  128 - 0x80
    "11100000", -- 3101 - 0xc1d  :  224 - 0xe0
    "00010000", -- 3102 - 0xc1e  :   16 - 0x10
    "11110000", -- 3103 - 0xc1f  :  240 - 0xf0
    "00000011", -- 3104 - 0xc20  :    3 - 0x3 -- Background 0x84
    "00001111", -- 3105 - 0xc21  :   15 - 0xf
    "00011100", -- 3106 - 0xc22  :   28 - 0x1c
    "00110000", -- 3107 - 0xc23  :   48 - 0x30
    "00100000", -- 3108 - 0xc24  :   32 - 0x20
    "01000000", -- 3109 - 0xc25  :   64 - 0x40
    "01000000", -- 3110 - 0xc26  :   64 - 0x40
    "01111111", -- 3111 - 0xc27  :  127 - 0x7f
    "00000011", -- 3112 - 0xc28  :    3 - 0x3 -- Background 0x85
    "00000110", -- 3113 - 0xc29  :    6 - 0x6
    "00000110", -- 3114 - 0xc2a  :    6 - 0x6
    "00011100", -- 3115 - 0xc2b  :   28 - 0x1c
    "00011000", -- 3116 - 0xc2c  :   24 - 0x18
    "00110110", -- 3117 - 0xc2d  :   54 - 0x36
    "00110001", -- 3118 - 0xc2e  :   49 - 0x31
    "00001111", -- 3119 - 0xc2f  :   15 - 0xf
    "11000000", -- 3120 - 0xc30  :  192 - 0xc0 -- Background 0x86
    "11110000", -- 3121 - 0xc31  :  240 - 0xf0
    "00111000", -- 3122 - 0xc32  :   56 - 0x38
    "00001110", -- 3123 - 0xc33  :   14 - 0xe
    "00011110", -- 3124 - 0xc34  :   30 - 0x1e
    "00011110", -- 3125 - 0xc35  :   30 - 0x1e
    "00000010", -- 3126 - 0xc36  :    2 - 0x2
    "11111110", -- 3127 - 0xc37  :  254 - 0xfe
    "11000000", -- 3128 - 0xc38  :  192 - 0xc0 -- Background 0x87
    "01100000", -- 3129 - 0xc39  :   96 - 0x60
    "01100000", -- 3130 - 0xc3a  :   96 - 0x60
    "00110000", -- 3131 - 0xc3b  :   48 - 0x30
    "00111110", -- 3132 - 0xc3c  :   62 - 0x3e
    "00011001", -- 3133 - 0xc3d  :   25 - 0x19
    "00110011", -- 3134 - 0xc3e  :   51 - 0x33
    "00111100", -- 3135 - 0xc3f  :   60 - 0x3c
    "00000011", -- 3136 - 0xc40  :    3 - 0x3 -- Background 0x88
    "00000111", -- 3137 - 0xc41  :    7 - 0x7
    "00000111", -- 3138 - 0xc42  :    7 - 0x7
    "00001011", -- 3139 - 0xc43  :   11 - 0xb
    "00010000", -- 3140 - 0xc44  :   16 - 0x10
    "01100000", -- 3141 - 0xc45  :   96 - 0x60
    "11110000", -- 3142 - 0xc46  :  240 - 0xf0
    "11110000", -- 3143 - 0xc47  :  240 - 0xf0
    "11110000", -- 3144 - 0xc48  :  240 - 0xf0 -- Background 0x89
    "11110000", -- 3145 - 0xc49  :  240 - 0xf0
    "01100000", -- 3146 - 0xc4a  :   96 - 0x60
    "00010000", -- 3147 - 0xc4b  :   16 - 0x10
    "00001011", -- 3148 - 0xc4c  :   11 - 0xb
    "00000111", -- 3149 - 0xc4d  :    7 - 0x7
    "00000111", -- 3150 - 0xc4e  :    7 - 0x7
    "00000011", -- 3151 - 0xc4f  :    3 - 0x3
    "00000000", -- 3152 - 0xc50  :    0 - 0x0 -- Background 0x8a
    "00011100", -- 3153 - 0xc51  :   28 - 0x1c
    "00111111", -- 3154 - 0xc52  :   63 - 0x3f
    "01111000", -- 3155 - 0xc53  :  120 - 0x78
    "01110000", -- 3156 - 0xc54  :  112 - 0x70
    "01100000", -- 3157 - 0xc55  :   96 - 0x60
    "00100000", -- 3158 - 0xc56  :   32 - 0x20
    "00100000", -- 3159 - 0xc57  :   32 - 0x20
    "00100000", -- 3160 - 0xc58  :   32 - 0x20 -- Background 0x8b
    "00100000", -- 3161 - 0xc59  :   32 - 0x20
    "01100000", -- 3162 - 0xc5a  :   96 - 0x60
    "01110000", -- 3163 - 0xc5b  :  112 - 0x70
    "01111000", -- 3164 - 0xc5c  :  120 - 0x78
    "00111111", -- 3165 - 0xc5d  :   63 - 0x3f
    "00011100", -- 3166 - 0xc5e  :   28 - 0x1c
    "00000000", -- 3167 - 0xc5f  :    0 - 0x0
    "00000011", -- 3168 - 0xc60  :    3 - 0x3 -- Background 0x8c
    "00001100", -- 3169 - 0xc61  :   12 - 0xc
    "00011110", -- 3170 - 0xc62  :   30 - 0x1e
    "00100110", -- 3171 - 0xc63  :   38 - 0x26
    "01000110", -- 3172 - 0xc64  :   70 - 0x46
    "01100100", -- 3173 - 0xc65  :  100 - 0x64
    "01110000", -- 3174 - 0xc66  :  112 - 0x70
    "11110000", -- 3175 - 0xc67  :  240 - 0xf0
    "10101010", -- 3176 - 0xc68  :  170 - 0xaa -- Background 0x8d
    "11111111", -- 3177 - 0xc69  :  255 - 0xff
    "01111111", -- 3178 - 0xc6a  :  127 - 0x7f
    "00111001", -- 3179 - 0xc6b  :   57 - 0x39
    "00011001", -- 3180 - 0xc6c  :   25 - 0x19
    "00001011", -- 3181 - 0xc6d  :   11 - 0xb
    "00001000", -- 3182 - 0xc6e  :    8 - 0x8
    "00000111", -- 3183 - 0xc6f  :    7 - 0x7
    "11000000", -- 3184 - 0xc70  :  192 - 0xc0 -- Background 0x8e
    "00110000", -- 3185 - 0xc71  :   48 - 0x30
    "00001000", -- 3186 - 0xc72  :    8 - 0x8
    "01000100", -- 3187 - 0xc73  :   68 - 0x44
    "01100010", -- 3188 - 0xc74  :   98 - 0x62
    "01100010", -- 3189 - 0xc75  :   98 - 0x62
    "00000001", -- 3190 - 0xc76  :    1 - 0x1
    "00111111", -- 3191 - 0xc77  :   63 - 0x3f
    "10001011", -- 3192 - 0xc78  :  139 - 0x8b -- Background 0x8f
    "11000001", -- 3193 - 0xc79  :  193 - 0xc1
    "11111110", -- 3194 - 0xc7a  :  254 - 0xfe
    "11111100", -- 3195 - 0xc7b  :  252 - 0xfc
    "11110000", -- 3196 - 0xc7c  :  240 - 0xf0
    "11110000", -- 3197 - 0xc7d  :  240 - 0xf0
    "11111000", -- 3198 - 0xc7e  :  248 - 0xf8
    "11110000", -- 3199 - 0xc7f  :  240 - 0xf0
    "00000011", -- 3200 - 0xc80  :    3 - 0x3 -- Background 0x90
    "00001110", -- 3201 - 0xc81  :   14 - 0xe
    "00010110", -- 3202 - 0xc82  :   22 - 0x16
    "00100110", -- 3203 - 0xc83  :   38 - 0x26
    "01100011", -- 3204 - 0xc84  :   99 - 0x63
    "01110010", -- 3205 - 0xc85  :  114 - 0x72
    "01110000", -- 3206 - 0xc86  :  112 - 0x70
    "11010000", -- 3207 - 0xc87  :  208 - 0xd0
    "10101010", -- 3208 - 0xc88  :  170 - 0xaa -- Background 0x91
    "11111111", -- 3209 - 0xc89  :  255 - 0xff
    "01111111", -- 3210 - 0xc8a  :  127 - 0x7f
    "00111100", -- 3211 - 0xc8b  :   60 - 0x3c
    "00011100", -- 3212 - 0xc8c  :   28 - 0x1c
    "00000100", -- 3213 - 0xc8d  :    4 - 0x4
    "00000010", -- 3214 - 0xc8e  :    2 - 0x2
    "00000001", -- 3215 - 0xc8f  :    1 - 0x1
    "11000000", -- 3216 - 0xc90  :  192 - 0xc0 -- Background 0x92
    "00110000", -- 3217 - 0xc91  :   48 - 0x30
    "00001000", -- 3218 - 0xc92  :    8 - 0x8
    "00100100", -- 3219 - 0xc93  :   36 - 0x24
    "00110010", -- 3220 - 0xc94  :   50 - 0x32
    "00110010", -- 3221 - 0xc95  :   50 - 0x32
    "00000001", -- 3222 - 0xc96  :    1 - 0x1
    "00011111", -- 3223 - 0xc97  :   31 - 0x1f
    "10001011", -- 3224 - 0xc98  :  139 - 0x8b -- Background 0x93
    "11000001", -- 3225 - 0xc99  :  193 - 0xc1
    "11111110", -- 3226 - 0xc9a  :  254 - 0xfe
    "11111100", -- 3227 - 0xc9b  :  252 - 0xfc
    "11110000", -- 3228 - 0xc9c  :  240 - 0xf0
    "11000000", -- 3229 - 0xc9d  :  192 - 0xc0
    "00100000", -- 3230 - 0xc9e  :   32 - 0x20
    "11100000", -- 3231 - 0xc9f  :  224 - 0xe0
    "00000011", -- 3232 - 0xca0  :    3 - 0x3 -- Background 0x94
    "00001111", -- 3233 - 0xca1  :   15 - 0xf
    "00010011", -- 3234 - 0xca2  :   19 - 0x13
    "00110001", -- 3235 - 0xca3  :   49 - 0x31
    "01111001", -- 3236 - 0xca4  :  121 - 0x79
    "01011001", -- 3237 - 0xca5  :   89 - 0x59
    "01001000", -- 3238 - 0xca6  :   72 - 0x48
    "11001100", -- 3239 - 0xca7  :  204 - 0xcc
    "10010101", -- 3240 - 0xca8  :  149 - 0x95 -- Background 0x95
    "11111111", -- 3241 - 0xca9  :  255 - 0xff
    "01111111", -- 3242 - 0xcaa  :  127 - 0x7f
    "00111110", -- 3243 - 0xcab  :   62 - 0x3e
    "00011111", -- 3244 - 0xcac  :   31 - 0x1f
    "00001111", -- 3245 - 0xcad  :   15 - 0xf
    "00001111", -- 3246 - 0xcae  :   15 - 0xf
    "00000111", -- 3247 - 0xcaf  :    7 - 0x7
    "11000000", -- 3248 - 0xcb0  :  192 - 0xc0 -- Background 0x96
    "00110000", -- 3249 - 0xcb1  :   48 - 0x30
    "00001000", -- 3250 - 0xcb2  :    8 - 0x8
    "10010100", -- 3251 - 0xcb3  :  148 - 0x94
    "10011010", -- 3252 - 0xcb4  :  154 - 0x9a
    "00011010", -- 3253 - 0xcb5  :   26 - 0x1a
    "00000001", -- 3254 - 0xcb6  :    1 - 0x1
    "00001111", -- 3255 - 0xcb7  :   15 - 0xf
    "01000101", -- 3256 - 0xcb8  :   69 - 0x45 -- Background 0x97
    "11100001", -- 3257 - 0xcb9  :  225 - 0xe1
    "11111110", -- 3258 - 0xcba  :  254 - 0xfe
    "01111100", -- 3259 - 0xcbb  :  124 - 0x7c
    "00110000", -- 3260 - 0xcbc  :   48 - 0x30
    "00110000", -- 3261 - 0xcbd  :   48 - 0x30
    "10001000", -- 3262 - 0xcbe  :  136 - 0x88
    "01111000", -- 3263 - 0xcbf  :  120 - 0x78
    "00000001", -- 3264 - 0xcc0  :    1 - 0x1 -- Background 0x98
    "00000000", -- 3265 - 0xcc1  :    0 - 0x0
    "00000000", -- 3266 - 0xcc2  :    0 - 0x0
    "00000000", -- 3267 - 0xcc3  :    0 - 0x0
    "00000001", -- 3268 - 0xcc4  :    1 - 0x1
    "00000001", -- 3269 - 0xcc5  :    1 - 0x1
    "00000010", -- 3270 - 0xcc6  :    2 - 0x2
    "00000110", -- 3271 - 0xcc7  :    6 - 0x6
    "01111000", -- 3272 - 0xcc8  :  120 - 0x78 -- Background 0x99
    "00101010", -- 3273 - 0xcc9  :   42 - 0x2a
    "01010100", -- 3274 - 0xcca  :   84 - 0x54
    "00101001", -- 3275 - 0xccb  :   41 - 0x29
    "00101111", -- 3276 - 0xccc  :   47 - 0x2f
    "00110111", -- 3277 - 0xccd  :   55 - 0x37
    "00000011", -- 3278 - 0xcce  :    3 - 0x3
    "00000111", -- 3279 - 0xccf  :    7 - 0x7
    "10110000", -- 3280 - 0xcd0  :  176 - 0xb0 -- Background 0x9a
    "11101000", -- 3281 - 0xcd1  :  232 - 0xe8
    "10001100", -- 3282 - 0xcd2  :  140 - 0x8c
    "10011110", -- 3283 - 0xcd3  :  158 - 0x9e
    "00011111", -- 3284 - 0xcd4  :   31 - 0x1f
    "00001111", -- 3285 - 0xcd5  :   15 - 0xf
    "10010110", -- 3286 - 0xcd6  :  150 - 0x96
    "00011100", -- 3287 - 0xcd7  :   28 - 0x1c
    "00001100", -- 3288 - 0xcd8  :   12 - 0xc -- Background 0x9b
    "00111000", -- 3289 - 0xcd9  :   56 - 0x38
    "11101000", -- 3290 - 0xcda  :  232 - 0xe8
    "11010000", -- 3291 - 0xcdb  :  208 - 0xd0
    "11100000", -- 3292 - 0xcdc  :  224 - 0xe0
    "10000000", -- 3293 - 0xcdd  :  128 - 0x80
    "00000000", -- 3294 - 0xcde  :    0 - 0x0
    "10000000", -- 3295 - 0xcdf  :  128 - 0x80
    "00000001", -- 3296 - 0xce0  :    1 - 0x1 -- Background 0x9c
    "00000000", -- 3297 - 0xce1  :    0 - 0x0
    "00000000", -- 3298 - 0xce2  :    0 - 0x0
    "00000000", -- 3299 - 0xce3  :    0 - 0x0
    "00000001", -- 3300 - 0xce4  :    1 - 0x1
    "00000001", -- 3301 - 0xce5  :    1 - 0x1
    "00000010", -- 3302 - 0xce6  :    2 - 0x2
    "00000110", -- 3303 - 0xce7  :    6 - 0x6
    "01111000", -- 3304 - 0xce8  :  120 - 0x78 -- Background 0x9d
    "00101010", -- 3305 - 0xce9  :   42 - 0x2a
    "01010100", -- 3306 - 0xcea  :   84 - 0x54
    "00101001", -- 3307 - 0xceb  :   41 - 0x29
    "00101111", -- 3308 - 0xcec  :   47 - 0x2f
    "00111100", -- 3309 - 0xced  :   60 - 0x3c
    "00011110", -- 3310 - 0xcee  :   30 - 0x1e
    "00000000", -- 3311 - 0xcef  :    0 - 0x0
    "10110000", -- 3312 - 0xcf0  :  176 - 0xb0 -- Background 0x9e
    "11101000", -- 3313 - 0xcf1  :  232 - 0xe8
    "10001100", -- 3314 - 0xcf2  :  140 - 0x8c
    "10011110", -- 3315 - 0xcf3  :  158 - 0x9e
    "00011111", -- 3316 - 0xcf4  :   31 - 0x1f
    "00001111", -- 3317 - 0xcf5  :   15 - 0xf
    "10010110", -- 3318 - 0xcf6  :  150 - 0x96
    "00011100", -- 3319 - 0xcf7  :   28 - 0x1c
    "00001100", -- 3320 - 0xcf8  :   12 - 0xc -- Background 0x9f
    "00111000", -- 3321 - 0xcf9  :   56 - 0x38
    "11101000", -- 3322 - 0xcfa  :  232 - 0xe8
    "11110000", -- 3323 - 0xcfb  :  240 - 0xf0
    "11000000", -- 3324 - 0xcfc  :  192 - 0xc0
    "01110000", -- 3325 - 0xcfd  :  112 - 0x70
    "11000000", -- 3326 - 0xcfe  :  192 - 0xc0
    "00000000", -- 3327 - 0xcff  :    0 - 0x0
    "00000011", -- 3328 - 0xd00  :    3 - 0x3 -- Background 0xa0
    "00001111", -- 3329 - 0xd01  :   15 - 0xf
    "00011100", -- 3330 - 0xd02  :   28 - 0x1c
    "00110000", -- 3331 - 0xd03  :   48 - 0x30
    "01100000", -- 3332 - 0xd04  :   96 - 0x60
    "01100000", -- 3333 - 0xd05  :   96 - 0x60
    "11000000", -- 3334 - 0xd06  :  192 - 0xc0
    "11000000", -- 3335 - 0xd07  :  192 - 0xc0
    "11000000", -- 3336 - 0xd08  :  192 - 0xc0 -- Background 0xa1
    "11000000", -- 3337 - 0xd09  :  192 - 0xc0
    "01100000", -- 3338 - 0xd0a  :   96 - 0x60
    "01100000", -- 3339 - 0xd0b  :   96 - 0x60
    "00110000", -- 3340 - 0xd0c  :   48 - 0x30
    "00011010", -- 3341 - 0xd0d  :   26 - 0x1a
    "00001101", -- 3342 - 0xd0e  :   13 - 0xd
    "00000011", -- 3343 - 0xd0f  :    3 - 0x3
    "11000000", -- 3344 - 0xd10  :  192 - 0xc0 -- Background 0xa2
    "11110000", -- 3345 - 0xd11  :  240 - 0xf0
    "00111000", -- 3346 - 0xd12  :   56 - 0x38
    "00001100", -- 3347 - 0xd13  :   12 - 0xc
    "00000110", -- 3348 - 0xd14  :    6 - 0x6
    "00000010", -- 3349 - 0xd15  :    2 - 0x2
    "00000101", -- 3350 - 0xd16  :    5 - 0x5
    "00000011", -- 3351 - 0xd17  :    3 - 0x3
    "00000101", -- 3352 - 0xd18  :    5 - 0x5 -- Background 0xa3
    "00001011", -- 3353 - 0xd19  :   11 - 0xb
    "00010110", -- 3354 - 0xd1a  :   22 - 0x16
    "00101010", -- 3355 - 0xd1b  :   42 - 0x2a
    "01010100", -- 3356 - 0xd1c  :   84 - 0x54
    "10101000", -- 3357 - 0xd1d  :  168 - 0xa8
    "01110000", -- 3358 - 0xd1e  :  112 - 0x70
    "11000000", -- 3359 - 0xd1f  :  192 - 0xc0
    "00000000", -- 3360 - 0xd20  :    0 - 0x0 -- Background 0xa4
    "00001111", -- 3361 - 0xd21  :   15 - 0xf
    "00011111", -- 3362 - 0xd22  :   31 - 0x1f
    "00110001", -- 3363 - 0xd23  :   49 - 0x31
    "00111111", -- 3364 - 0xd24  :   63 - 0x3f
    "01111111", -- 3365 - 0xd25  :  127 - 0x7f
    "11111111", -- 3366 - 0xd26  :  255 - 0xff
    "11011111", -- 3367 - 0xd27  :  223 - 0xdf
    "11000000", -- 3368 - 0xd28  :  192 - 0xc0 -- Background 0xa5
    "11000111", -- 3369 - 0xd29  :  199 - 0xc7
    "01101111", -- 3370 - 0xd2a  :  111 - 0x6f
    "01100111", -- 3371 - 0xd2b  :  103 - 0x67
    "01100011", -- 3372 - 0xd2c  :   99 - 0x63
    "00110000", -- 3373 - 0xd2d  :   48 - 0x30
    "00011000", -- 3374 - 0xd2e  :   24 - 0x18
    "00000111", -- 3375 - 0xd2f  :    7 - 0x7
    "00000000", -- 3376 - 0xd30  :    0 - 0x0 -- Background 0xa6
    "11110000", -- 3377 - 0xd31  :  240 - 0xf0
    "11111000", -- 3378 - 0xd32  :  248 - 0xf8
    "10001100", -- 3379 - 0xd33  :  140 - 0x8c
    "11111100", -- 3380 - 0xd34  :  252 - 0xfc
    "11111110", -- 3381 - 0xd35  :  254 - 0xfe
    "11111101", -- 3382 - 0xd36  :  253 - 0xfd
    "11111001", -- 3383 - 0xd37  :  249 - 0xf9
    "00000011", -- 3384 - 0xd38  :    3 - 0x3 -- Background 0xa7
    "11100101", -- 3385 - 0xd39  :  229 - 0xe5
    "11110010", -- 3386 - 0xd3a  :  242 - 0xf2
    "11100110", -- 3387 - 0xd3b  :  230 - 0xe6
    "11001010", -- 3388 - 0xd3c  :  202 - 0xca
    "00010100", -- 3389 - 0xd3d  :   20 - 0x14
    "00111000", -- 3390 - 0xd3e  :   56 - 0x38
    "11100000", -- 3391 - 0xd3f  :  224 - 0xe0
    "00000000", -- 3392 - 0xd40  :    0 - 0x0 -- Background 0xa8
    "00001111", -- 3393 - 0xd41  :   15 - 0xf
    "00011111", -- 3394 - 0xd42  :   31 - 0x1f
    "00110001", -- 3395 - 0xd43  :   49 - 0x31
    "00111111", -- 3396 - 0xd44  :   63 - 0x3f
    "01111111", -- 3397 - 0xd45  :  127 - 0x7f
    "11111111", -- 3398 - 0xd46  :  255 - 0xff
    "11011111", -- 3399 - 0xd47  :  223 - 0xdf
    "11000000", -- 3400 - 0xd48  :  192 - 0xc0 -- Background 0xa9
    "11000011", -- 3401 - 0xd49  :  195 - 0xc3
    "11000111", -- 3402 - 0xd4a  :  199 - 0xc7
    "11001111", -- 3403 - 0xd4b  :  207 - 0xcf
    "11000111", -- 3404 - 0xd4c  :  199 - 0xc7
    "11000000", -- 3405 - 0xd4d  :  192 - 0xc0
    "11100000", -- 3406 - 0xd4e  :  224 - 0xe0
    "11111111", -- 3407 - 0xd4f  :  255 - 0xff
    "00000000", -- 3408 - 0xd50  :    0 - 0x0 -- Background 0xaa
    "11110000", -- 3409 - 0xd51  :  240 - 0xf0
    "11111000", -- 3410 - 0xd52  :  248 - 0xf8
    "10001100", -- 3411 - 0xd53  :  140 - 0x8c
    "11111100", -- 3412 - 0xd54  :  252 - 0xfc
    "11111110", -- 3413 - 0xd55  :  254 - 0xfe
    "11111101", -- 3414 - 0xd56  :  253 - 0xfd
    "11111001", -- 3415 - 0xd57  :  249 - 0xf9
    "00000011", -- 3416 - 0xd58  :    3 - 0x3 -- Background 0xab
    "11000101", -- 3417 - 0xd59  :  197 - 0xc5
    "11100011", -- 3418 - 0xd5a  :  227 - 0xe3
    "11110101", -- 3419 - 0xd5b  :  245 - 0xf5
    "11100011", -- 3420 - 0xd5c  :  227 - 0xe3
    "00000101", -- 3421 - 0xd5d  :    5 - 0x5
    "00001011", -- 3422 - 0xd5e  :   11 - 0xb
    "11111111", -- 3423 - 0xd5f  :  255 - 0xff
    "10000011", -- 3424 - 0xd60  :  131 - 0x83 -- Background 0xac
    "10001100", -- 3425 - 0xd61  :  140 - 0x8c
    "10010000", -- 3426 - 0xd62  :  144 - 0x90
    "10010000", -- 3427 - 0xd63  :  144 - 0x90
    "11100000", -- 3428 - 0xd64  :  224 - 0xe0
    "10100000", -- 3429 - 0xd65  :  160 - 0xa0
    "10101111", -- 3430 - 0xd66  :  175 - 0xaf
    "01101111", -- 3431 - 0xd67  :  111 - 0x6f
    "11111011", -- 3432 - 0xd68  :  251 - 0xfb -- Background 0xad
    "00000101", -- 3433 - 0xd69  :    5 - 0x5
    "00000101", -- 3434 - 0xd6a  :    5 - 0x5
    "00000101", -- 3435 - 0xd6b  :    5 - 0x5
    "01000101", -- 3436 - 0xd6c  :   69 - 0x45
    "01100101", -- 3437 - 0xd6d  :  101 - 0x65
    "11110101", -- 3438 - 0xd6e  :  245 - 0xf5
    "11111101", -- 3439 - 0xd6f  :  253 - 0xfd
    "10000011", -- 3440 - 0xd70  :  131 - 0x83 -- Background 0xae
    "10001100", -- 3441 - 0xd71  :  140 - 0x8c
    "10010000", -- 3442 - 0xd72  :  144 - 0x90
    "10010000", -- 3443 - 0xd73  :  144 - 0x90
    "11100000", -- 3444 - 0xd74  :  224 - 0xe0
    "10100000", -- 3445 - 0xd75  :  160 - 0xa0
    "10101111", -- 3446 - 0xd76  :  175 - 0xaf
    "01101111", -- 3447 - 0xd77  :  111 - 0x6f
    "11111011", -- 3448 - 0xd78  :  251 - 0xfb -- Background 0xaf
    "00000101", -- 3449 - 0xd79  :    5 - 0x5
    "00000101", -- 3450 - 0xd7a  :    5 - 0x5
    "00000101", -- 3451 - 0xd7b  :    5 - 0x5
    "11000101", -- 3452 - 0xd7c  :  197 - 0xc5
    "11100101", -- 3453 - 0xd7d  :  229 - 0xe5
    "11110101", -- 3454 - 0xd7e  :  245 - 0xf5
    "11111101", -- 3455 - 0xd7f  :  253 - 0xfd
    "00000000", -- 3456 - 0xd80  :    0 - 0x0 -- Background 0xb0
    "00000011", -- 3457 - 0xd81  :    3 - 0x3
    "00001111", -- 3458 - 0xd82  :   15 - 0xf
    "00111111", -- 3459 - 0xd83  :   63 - 0x3f
    "01111111", -- 3460 - 0xd84  :  127 - 0x7f
    "01111111", -- 3461 - 0xd85  :  127 - 0x7f
    "11111111", -- 3462 - 0xd86  :  255 - 0xff
    "11111111", -- 3463 - 0xd87  :  255 - 0xff
    "11111111", -- 3464 - 0xd88  :  255 - 0xff -- Background 0xb1
    "10001111", -- 3465 - 0xd89  :  143 - 0x8f
    "10000000", -- 3466 - 0xd8a  :  128 - 0x80
    "11110000", -- 3467 - 0xd8b  :  240 - 0xf0
    "11111111", -- 3468 - 0xd8c  :  255 - 0xff
    "11111111", -- 3469 - 0xd8d  :  255 - 0xff
    "01111111", -- 3470 - 0xd8e  :  127 - 0x7f
    "00001111", -- 3471 - 0xd8f  :   15 - 0xf
    "00000000", -- 3472 - 0xd90  :    0 - 0x0 -- Background 0xb2
    "11000000", -- 3473 - 0xd91  :  192 - 0xc0
    "11110000", -- 3474 - 0xd92  :  240 - 0xf0
    "11111100", -- 3475 - 0xd93  :  252 - 0xfc
    "11111110", -- 3476 - 0xd94  :  254 - 0xfe
    "11111110", -- 3477 - 0xd95  :  254 - 0xfe
    "11111111", -- 3478 - 0xd96  :  255 - 0xff
    "11111111", -- 3479 - 0xd97  :  255 - 0xff
    "11111111", -- 3480 - 0xd98  :  255 - 0xff -- Background 0xb3
    "11110001", -- 3481 - 0xd99  :  241 - 0xf1
    "00000001", -- 3482 - 0xd9a  :    1 - 0x1
    "00001111", -- 3483 - 0xd9b  :   15 - 0xf
    "11111111", -- 3484 - 0xd9c  :  255 - 0xff
    "11111111", -- 3485 - 0xd9d  :  255 - 0xff
    "11111110", -- 3486 - 0xd9e  :  254 - 0xfe
    "11110000", -- 3487 - 0xd9f  :  240 - 0xf0
    "00000000", -- 3488 - 0xda0  :    0 - 0x0 -- Background 0xb4
    "00000011", -- 3489 - 0xda1  :    3 - 0x3
    "00001110", -- 3490 - 0xda2  :   14 - 0xe
    "00110101", -- 3491 - 0xda3  :   53 - 0x35
    "01101110", -- 3492 - 0xda4  :  110 - 0x6e
    "01010101", -- 3493 - 0xda5  :   85 - 0x55
    "10111010", -- 3494 - 0xda6  :  186 - 0xba
    "11010111", -- 3495 - 0xda7  :  215 - 0xd7
    "11111010", -- 3496 - 0xda8  :  250 - 0xfa -- Background 0xb5
    "10001111", -- 3497 - 0xda9  :  143 - 0x8f
    "10000000", -- 3498 - 0xdaa  :  128 - 0x80
    "11110000", -- 3499 - 0xdab  :  240 - 0xf0
    "10101111", -- 3500 - 0xdac  :  175 - 0xaf
    "11010101", -- 3501 - 0xdad  :  213 - 0xd5
    "01111010", -- 3502 - 0xdae  :  122 - 0x7a
    "00001111", -- 3503 - 0xdaf  :   15 - 0xf
    "00000000", -- 3504 - 0xdb0  :    0 - 0x0 -- Background 0xb6
    "11000000", -- 3505 - 0xdb1  :  192 - 0xc0
    "10110000", -- 3506 - 0xdb2  :  176 - 0xb0
    "01011100", -- 3507 - 0xdb3  :   92 - 0x5c
    "11101010", -- 3508 - 0xdb4  :  234 - 0xea
    "01011110", -- 3509 - 0xdb5  :   94 - 0x5e
    "10101011", -- 3510 - 0xdb6  :  171 - 0xab
    "01110101", -- 3511 - 0xdb7  :  117 - 0x75
    "10101111", -- 3512 - 0xdb8  :  175 - 0xaf -- Background 0xb7
    "11110001", -- 3513 - 0xdb9  :  241 - 0xf1
    "00000001", -- 3514 - 0xdba  :    1 - 0x1
    "00001111", -- 3515 - 0xdbb  :   15 - 0xf
    "11111011", -- 3516 - 0xdbc  :  251 - 0xfb
    "01010101", -- 3517 - 0xdbd  :   85 - 0x55
    "10101110", -- 3518 - 0xdbe  :  174 - 0xae
    "11110000", -- 3519 - 0xdbf  :  240 - 0xf0
    "00000000", -- 3520 - 0xdc0  :    0 - 0x0 -- Background 0xb8
    "00000011", -- 3521 - 0xdc1  :    3 - 0x3
    "00001100", -- 3522 - 0xdc2  :   12 - 0xc
    "00110000", -- 3523 - 0xdc3  :   48 - 0x30
    "01000100", -- 3524 - 0xdc4  :   68 - 0x44
    "01000000", -- 3525 - 0xdc5  :   64 - 0x40
    "10010000", -- 3526 - 0xdc6  :  144 - 0x90
    "10000010", -- 3527 - 0xdc7  :  130 - 0x82
    "11110000", -- 3528 - 0xdc8  :  240 - 0xf0 -- Background 0xb9
    "11111111", -- 3529 - 0xdc9  :  255 - 0xff
    "11111111", -- 3530 - 0xdca  :  255 - 0xff
    "11111111", -- 3531 - 0xdcb  :  255 - 0xff
    "10001111", -- 3532 - 0xdcc  :  143 - 0x8f
    "10000000", -- 3533 - 0xdcd  :  128 - 0x80
    "01110000", -- 3534 - 0xdce  :  112 - 0x70
    "00001111", -- 3535 - 0xdcf  :   15 - 0xf
    "00000000", -- 3536 - 0xdd0  :    0 - 0x0 -- Background 0xba
    "11000000", -- 3537 - 0xdd1  :  192 - 0xc0
    "00110000", -- 3538 - 0xdd2  :   48 - 0x30
    "00001100", -- 3539 - 0xdd3  :   12 - 0xc
    "01000010", -- 3540 - 0xdd4  :   66 - 0x42
    "00001010", -- 3541 - 0xdd5  :   10 - 0xa
    "00000001", -- 3542 - 0xdd6  :    1 - 0x1
    "00100001", -- 3543 - 0xdd7  :   33 - 0x21
    "00001111", -- 3544 - 0xdd8  :   15 - 0xf -- Background 0xbb
    "11111111", -- 3545 - 0xdd9  :  255 - 0xff
    "11111111", -- 3546 - 0xdda  :  255 - 0xff
    "11111111", -- 3547 - 0xddb  :  255 - 0xff
    "11110001", -- 3548 - 0xddc  :  241 - 0xf1
    "00000001", -- 3549 - 0xddd  :    1 - 0x1
    "00001110", -- 3550 - 0xdde  :   14 - 0xe
    "11110000", -- 3551 - 0xddf  :  240 - 0xf0
    "11110011", -- 3552 - 0xde0  :  243 - 0xf3 -- Background 0xbc
    "11111111", -- 3553 - 0xde1  :  255 - 0xff
    "11000100", -- 3554 - 0xde2  :  196 - 0xc4
    "11000000", -- 3555 - 0xde3  :  192 - 0xc0
    "01000000", -- 3556 - 0xde4  :   64 - 0x40
    "01100011", -- 3557 - 0xde5  :   99 - 0x63
    "11000111", -- 3558 - 0xde6  :  199 - 0xc7
    "11000110", -- 3559 - 0xde7  :  198 - 0xc6
    "11000110", -- 3560 - 0xde8  :  198 - 0xc6 -- Background 0xbd
    "11000110", -- 3561 - 0xde9  :  198 - 0xc6
    "01100011", -- 3562 - 0xdea  :   99 - 0x63
    "01000000", -- 3563 - 0xdeb  :   64 - 0x40
    "11000000", -- 3564 - 0xdec  :  192 - 0xc0
    "11000100", -- 3565 - 0xded  :  196 - 0xc4
    "11001100", -- 3566 - 0xdee  :  204 - 0xcc
    "11110011", -- 3567 - 0xdef  :  243 - 0xf3
    "11001111", -- 3568 - 0xdf0  :  207 - 0xcf -- Background 0xbe
    "11111111", -- 3569 - 0xdf1  :  255 - 0xff
    "00100001", -- 3570 - 0xdf2  :   33 - 0x21
    "00000001", -- 3571 - 0xdf3  :    1 - 0x1
    "00000010", -- 3572 - 0xdf4  :    2 - 0x2
    "11000110", -- 3573 - 0xdf5  :  198 - 0xc6
    "11100001", -- 3574 - 0xdf6  :  225 - 0xe1
    "00100001", -- 3575 - 0xdf7  :   33 - 0x21
    "00100001", -- 3576 - 0xdf8  :   33 - 0x21 -- Background 0xbf
    "00100001", -- 3577 - 0xdf9  :   33 - 0x21
    "11000110", -- 3578 - 0xdfa  :  198 - 0xc6
    "00000010", -- 3579 - 0xdfb  :    2 - 0x2
    "00000001", -- 3580 - 0xdfc  :    1 - 0x1
    "00100001", -- 3581 - 0xdfd  :   33 - 0x21
    "00110001", -- 3582 - 0xdfe  :   49 - 0x31
    "11001111", -- 3583 - 0xdff  :  207 - 0xcf
    "00000000", -- 3584 - 0xe00  :    0 - 0x0 -- Background 0xc0
    "01010000", -- 3585 - 0xe01  :   80 - 0x50
    "10110011", -- 3586 - 0xe02  :  179 - 0xb3
    "10010111", -- 3587 - 0xe03  :  151 - 0x97
    "10011111", -- 3588 - 0xe04  :  159 - 0x9f
    "01101111", -- 3589 - 0xe05  :  111 - 0x6f
    "00011111", -- 3590 - 0xe06  :   31 - 0x1f
    "00011111", -- 3591 - 0xe07  :   31 - 0x1f
    "00011111", -- 3592 - 0xe08  :   31 - 0x1f -- Background 0xc1
    "00011111", -- 3593 - 0xe09  :   31 - 0x1f
    "00001111", -- 3594 - 0xe0a  :   15 - 0xf
    "00000111", -- 3595 - 0xe0b  :    7 - 0x7
    "00011101", -- 3596 - 0xe0c  :   29 - 0x1d
    "00101100", -- 3597 - 0xe0d  :   44 - 0x2c
    "01010100", -- 3598 - 0xe0e  :   84 - 0x54
    "01111100", -- 3599 - 0xe0f  :  124 - 0x7c
    "00000000", -- 3600 - 0xe10  :    0 - 0x0 -- Background 0xc2
    "00001010", -- 3601 - 0xe11  :   10 - 0xa
    "11001101", -- 3602 - 0xe12  :  205 - 0xcd
    "11101001", -- 3603 - 0xe13  :  233 - 0xe9
    "11111001", -- 3604 - 0xe14  :  249 - 0xf9
    "11110110", -- 3605 - 0xe15  :  246 - 0xf6
    "11110000", -- 3606 - 0xe16  :  240 - 0xf0
    "11111000", -- 3607 - 0xe17  :  248 - 0xf8
    "11111000", -- 3608 - 0xe18  :  248 - 0xf8 -- Background 0xc3
    "11111000", -- 3609 - 0xe19  :  248 - 0xf8
    "11110000", -- 3610 - 0xe1a  :  240 - 0xf0
    "11000000", -- 3611 - 0xe1b  :  192 - 0xc0
    "10111000", -- 3612 - 0xe1c  :  184 - 0xb8
    "00110100", -- 3613 - 0xe1d  :   52 - 0x34
    "00101010", -- 3614 - 0xe1e  :   42 - 0x2a
    "00111110", -- 3615 - 0xe1f  :   62 - 0x3e
    "00000101", -- 3616 - 0xe20  :    5 - 0x5 -- Background 0xc4
    "00001010", -- 3617 - 0xe21  :   10 - 0xa
    "00001000", -- 3618 - 0xe22  :    8 - 0x8
    "00001111", -- 3619 - 0xe23  :   15 - 0xf
    "00000001", -- 3620 - 0xe24  :    1 - 0x1
    "00000011", -- 3621 - 0xe25  :    3 - 0x3
    "00000111", -- 3622 - 0xe26  :    7 - 0x7
    "00001111", -- 3623 - 0xe27  :   15 - 0xf
    "00001111", -- 3624 - 0xe28  :   15 - 0xf -- Background 0xc5
    "11101111", -- 3625 - 0xe29  :  239 - 0xef
    "11011111", -- 3626 - 0xe2a  :  223 - 0xdf
    "10101111", -- 3627 - 0xe2b  :  175 - 0xaf
    "01100111", -- 3628 - 0xe2c  :  103 - 0x67
    "00001101", -- 3629 - 0xe2d  :   13 - 0xd
    "00001010", -- 3630 - 0xe2e  :   10 - 0xa
    "00000111", -- 3631 - 0xe2f  :    7 - 0x7
    "00000000", -- 3632 - 0xe30  :    0 - 0x0 -- Background 0xc6
    "10000000", -- 3633 - 0xe31  :  128 - 0x80
    "10000000", -- 3634 - 0xe32  :  128 - 0x80
    "11110000", -- 3635 - 0xe33  :  240 - 0xf0
    "11111000", -- 3636 - 0xe34  :  248 - 0xf8
    "11111100", -- 3637 - 0xe35  :  252 - 0xfc
    "11111100", -- 3638 - 0xe36  :  252 - 0xfc
    "11111100", -- 3639 - 0xe37  :  252 - 0xfc
    "11111100", -- 3640 - 0xe38  :  252 - 0xfc -- Background 0xc7
    "11111110", -- 3641 - 0xe39  :  254 - 0xfe
    "11111001", -- 3642 - 0xe3a  :  249 - 0xf9
    "11111010", -- 3643 - 0xe3b  :  250 - 0xfa
    "11101001", -- 3644 - 0xe3c  :  233 - 0xe9
    "00001110", -- 3645 - 0xe3d  :   14 - 0xe
    "10000000", -- 3646 - 0xe3e  :  128 - 0x80
    "00000000", -- 3647 - 0xe3f  :    0 - 0x0
    "00000000", -- 3648 - 0xe40  :    0 - 0x0 -- Background 0xc8
    "11000000", -- 3649 - 0xe41  :  192 - 0xc0
    "10100000", -- 3650 - 0xe42  :  160 - 0xa0
    "11010011", -- 3651 - 0xe43  :  211 - 0xd3
    "10110111", -- 3652 - 0xe44  :  183 - 0xb7
    "11111111", -- 3653 - 0xe45  :  255 - 0xff
    "00001111", -- 3654 - 0xe46  :   15 - 0xf
    "00011111", -- 3655 - 0xe47  :   31 - 0x1f
    "00011111", -- 3656 - 0xe48  :   31 - 0x1f -- Background 0xc9
    "00001111", -- 3657 - 0xe49  :   15 - 0xf
    "11110111", -- 3658 - 0xe4a  :  247 - 0xf7
    "10110111", -- 3659 - 0xe4b  :  183 - 0xb7
    "11010011", -- 3660 - 0xe4c  :  211 - 0xd3
    "10100000", -- 3661 - 0xe4d  :  160 - 0xa0
    "11000000", -- 3662 - 0xe4e  :  192 - 0xc0
    "00000000", -- 3663 - 0xe4f  :    0 - 0x0
    "00011100", -- 3664 - 0xe50  :   28 - 0x1c -- Background 0xca
    "00100010", -- 3665 - 0xe51  :   34 - 0x22
    "00100100", -- 3666 - 0xe52  :   36 - 0x24
    "11011110", -- 3667 - 0xe53  :  222 - 0xde
    "11110000", -- 3668 - 0xe54  :  240 - 0xf0
    "11111000", -- 3669 - 0xe55  :  248 - 0xf8
    "11111100", -- 3670 - 0xe56  :  252 - 0xfc
    "11111100", -- 3671 - 0xe57  :  252 - 0xfc
    "11111100", -- 3672 - 0xe58  :  252 - 0xfc -- Background 0xcb
    "11111100", -- 3673 - 0xe59  :  252 - 0xfc
    "11111000", -- 3674 - 0xe5a  :  248 - 0xf8
    "11110000", -- 3675 - 0xe5b  :  240 - 0xf0
    "10011110", -- 3676 - 0xe5c  :  158 - 0x9e
    "00100100", -- 3677 - 0xe5d  :   36 - 0x24
    "00100010", -- 3678 - 0xe5e  :   34 - 0x22
    "00011100", -- 3679 - 0xe5f  :   28 - 0x1c
    "00001110", -- 3680 - 0xe60  :   14 - 0xe -- Background 0xcc
    "00010110", -- 3681 - 0xe61  :   22 - 0x16
    "00011010", -- 3682 - 0xe62  :   26 - 0x1a
    "00000100", -- 3683 - 0xe63  :    4 - 0x4
    "01101111", -- 3684 - 0xe64  :  111 - 0x6f
    "10111111", -- 3685 - 0xe65  :  191 - 0xbf
    "11011111", -- 3686 - 0xe66  :  223 - 0xdf
    "10111111", -- 3687 - 0xe67  :  191 - 0xbf
    "01011111", -- 3688 - 0xe68  :   95 - 0x5f -- Background 0xcd
    "00011111", -- 3689 - 0xe69  :   31 - 0x1f
    "00011111", -- 3690 - 0xe6a  :   31 - 0x1f
    "00001111", -- 3691 - 0xe6b  :   15 - 0xf
    "00111111", -- 3692 - 0xe6c  :   63 - 0x3f
    "00100011", -- 3693 - 0xe6d  :   35 - 0x23
    "00101010", -- 3694 - 0xe6e  :   42 - 0x2a
    "00010100", -- 3695 - 0xe6f  :   20 - 0x14
    "00000000", -- 3696 - 0xe70  :    0 - 0x0 -- Background 0xce
    "00000000", -- 3697 - 0xe71  :    0 - 0x0
    "00000000", -- 3698 - 0xe72  :    0 - 0x0
    "00000000", -- 3699 - 0xe73  :    0 - 0x0
    "10001110", -- 3700 - 0xe74  :  142 - 0x8e
    "11001001", -- 3701 - 0xe75  :  201 - 0xc9
    "11101010", -- 3702 - 0xe76  :  234 - 0xea
    "11111001", -- 3703 - 0xe77  :  249 - 0xf9
    "11111110", -- 3704 - 0xe78  :  254 - 0xfe -- Background 0xcf
    "11111000", -- 3705 - 0xe79  :  248 - 0xf8
    "11111000", -- 3706 - 0xe7a  :  248 - 0xf8
    "11111000", -- 3707 - 0xe7b  :  248 - 0xf8
    "11110000", -- 3708 - 0xe7c  :  240 - 0xf0
    "11100000", -- 3709 - 0xe7d  :  224 - 0xe0
    "00000000", -- 3710 - 0xe7e  :    0 - 0x0
    "00000000", -- 3711 - 0xe7f  :    0 - 0x0
    "00000000", -- 3712 - 0xe80  :    0 - 0x0 -- Background 0xd0
    "00000000", -- 3713 - 0xe81  :    0 - 0x0
    "00000100", -- 3714 - 0xe82  :    4 - 0x4
    "00100110", -- 3715 - 0xe83  :   38 - 0x26
    "00101011", -- 3716 - 0xe84  :   43 - 0x2b
    "01110001", -- 3717 - 0xe85  :  113 - 0x71
    "01000000", -- 3718 - 0xe86  :   64 - 0x40
    "01000111", -- 3719 - 0xe87  :   71 - 0x47
    "10001111", -- 3720 - 0xe88  :  143 - 0x8f -- Background 0xd1
    "10001111", -- 3721 - 0xe89  :  143 - 0x8f
    "01001111", -- 3722 - 0xe8a  :   79 - 0x4f
    "01001111", -- 3723 - 0xe8b  :   79 - 0x4f
    "00111111", -- 3724 - 0xe8c  :   63 - 0x3f
    "00010011", -- 3725 - 0xe8d  :   19 - 0x13
    "00010001", -- 3726 - 0xe8e  :   17 - 0x11
    "00011111", -- 3727 - 0xe8f  :   31 - 0x1f
    "00000000", -- 3728 - 0xe90  :    0 - 0x0 -- Background 0xd2
    "10000000", -- 3729 - 0xe91  :  128 - 0x80
    "11001000", -- 3730 - 0xe92  :  200 - 0xc8
    "11010100", -- 3731 - 0xe93  :  212 - 0xd4
    "00100100", -- 3732 - 0xe94  :   36 - 0x24
    "00000010", -- 3733 - 0xe95  :    2 - 0x2
    "00000010", -- 3734 - 0xe96  :    2 - 0x2
    "11110010", -- 3735 - 0xe97  :  242 - 0xf2
    "11110010", -- 3736 - 0xe98  :  242 - 0xf2 -- Background 0xd3
    "11110010", -- 3737 - 0xe99  :  242 - 0xf2
    "11110100", -- 3738 - 0xe9a  :  244 - 0xf4
    "11110100", -- 3739 - 0xe9b  :  244 - 0xf4
    "11110100", -- 3740 - 0xe9c  :  244 - 0xf4
    "11001000", -- 3741 - 0xe9d  :  200 - 0xc8
    "01000100", -- 3742 - 0xe9e  :   68 - 0x44
    "01111100", -- 3743 - 0xe9f  :  124 - 0x7c
    "00000000", -- 3744 - 0xea0  :    0 - 0x0 -- Background 0xd4
    "00000000", -- 3745 - 0xea1  :    0 - 0x0
    "00000000", -- 3746 - 0xea2  :    0 - 0x0
    "00001001", -- 3747 - 0xea3  :    9 - 0x9
    "00011010", -- 3748 - 0xea4  :   26 - 0x1a
    "00010100", -- 3749 - 0xea5  :   20 - 0x14
    "00100000", -- 3750 - 0xea6  :   32 - 0x20
    "01000111", -- 3751 - 0xea7  :   71 - 0x47
    "10001111", -- 3752 - 0xea8  :  143 - 0x8f -- Background 0xd5
    "10001111", -- 3753 - 0xea9  :  143 - 0x8f
    "01001111", -- 3754 - 0xeaa  :   79 - 0x4f
    "01001111", -- 3755 - 0xeab  :   79 - 0x4f
    "00111111", -- 3756 - 0xeac  :   63 - 0x3f
    "01000111", -- 3757 - 0xead  :   71 - 0x47
    "00100010", -- 3758 - 0xeae  :   34 - 0x22
    "00011100", -- 3759 - 0xeaf  :   28 - 0x1c
    "00000000", -- 3760 - 0xeb0  :    0 - 0x0 -- Background 0xd6
    "01000000", -- 3761 - 0xeb1  :   64 - 0x40
    "11000000", -- 3762 - 0xeb2  :  192 - 0xc0
    "00101100", -- 3763 - 0xeb3  :   44 - 0x2c
    "00110100", -- 3764 - 0xeb4  :   52 - 0x34
    "00000100", -- 3765 - 0xeb5  :    4 - 0x4
    "00000010", -- 3766 - 0xeb6  :    2 - 0x2
    "11110010", -- 3767 - 0xeb7  :  242 - 0xf2
    "11110010", -- 3768 - 0xeb8  :  242 - 0xf2 -- Background 0xd7
    "11110010", -- 3769 - 0xeb9  :  242 - 0xf2
    "11110100", -- 3770 - 0xeba  :  244 - 0xf4
    "11110111", -- 3771 - 0xebb  :  247 - 0xf7
    "11111101", -- 3772 - 0xebc  :  253 - 0xfd
    "11100001", -- 3773 - 0xebd  :  225 - 0xe1
    "00010010", -- 3774 - 0xebe  :   18 - 0x12
    "00001100", -- 3775 - 0xebf  :   12 - 0xc
    "01111000", -- 3776 - 0xec0  :  120 - 0x78 -- Background 0xd8
    "01001110", -- 3777 - 0xec1  :   78 - 0x4e
    "11000010", -- 3778 - 0xec2  :  194 - 0xc2
    "10011010", -- 3779 - 0xec3  :  154 - 0x9a
    "10011011", -- 3780 - 0xec4  :  155 - 0x9b
    "11011001", -- 3781 - 0xec5  :  217 - 0xd9
    "01100011", -- 3782 - 0xec6  :   99 - 0x63
    "00111110", -- 3783 - 0xec7  :   62 - 0x3e
    "00011110", -- 3784 - 0xec8  :   30 - 0x1e -- Background 0xd9
    "01110001", -- 3785 - 0xec9  :  113 - 0x71
    "01001001", -- 3786 - 0xeca  :   73 - 0x49
    "10111001", -- 3787 - 0xecb  :  185 - 0xb9
    "10011101", -- 3788 - 0xecc  :  157 - 0x9d
    "01010010", -- 3789 - 0xecd  :   82 - 0x52
    "01110010", -- 3790 - 0xece  :  114 - 0x72
    "00011110", -- 3791 - 0xecf  :   30 - 0x1e
    "01100000", -- 3792 - 0xed0  :   96 - 0x60 -- Background 0xda
    "01011110", -- 3793 - 0xed1  :   94 - 0x5e
    "10001001", -- 3794 - 0xed2  :  137 - 0x89
    "10111101", -- 3795 - 0xed3  :  189 - 0xbd
    "10011101", -- 3796 - 0xed4  :  157 - 0x9d
    "11010011", -- 3797 - 0xed5  :  211 - 0xd3
    "01000110", -- 3798 - 0xed6  :   70 - 0x46
    "01111100", -- 3799 - 0xed7  :  124 - 0x7c
    "00011110", -- 3800 - 0xed8  :   30 - 0x1e -- Background 0xdb
    "00100011", -- 3801 - 0xed9  :   35 - 0x23
    "01001001", -- 3802 - 0xeda  :   73 - 0x49
    "10111101", -- 3803 - 0xedb  :  189 - 0xbd
    "10011001", -- 3804 - 0xedc  :  153 - 0x99
    "01000011", -- 3805 - 0xedd  :   67 - 0x43
    "01101110", -- 3806 - 0xede  :  110 - 0x6e
    "00011000", -- 3807 - 0xedf  :   24 - 0x18
    "00000000", -- 3808 - 0xee0  :    0 - 0x0 -- Background 0xdc
    "00000000", -- 3809 - 0xee1  :    0 - 0x0
    "00000001", -- 3810 - 0xee2  :    1 - 0x1
    "00000010", -- 3811 - 0xee3  :    2 - 0x2
    "00000100", -- 3812 - 0xee4  :    4 - 0x4
    "00000010", -- 3813 - 0xee5  :    2 - 0x2
    "00011110", -- 3814 - 0xee6  :   30 - 0x1e
    "00010000", -- 3815 - 0xee7  :   16 - 0x10
    "00001000", -- 3816 - 0xee8  :    8 - 0x8 -- Background 0xdd
    "00001101", -- 3817 - 0xee9  :   13 - 0xd
    "00111010", -- 3818 - 0xeea  :   58 - 0x3a
    "00100101", -- 3819 - 0xeeb  :   37 - 0x25
    "00011011", -- 3820 - 0xeec  :   27 - 0x1b
    "00001111", -- 3821 - 0xeed  :   15 - 0xf
    "00000111", -- 3822 - 0xeee  :    7 - 0x7
    "00000011", -- 3823 - 0xeef  :    3 - 0x3
    "00000000", -- 3824 - 0xef0  :    0 - 0x0 -- Background 0xde
    "00000000", -- 3825 - 0xef1  :    0 - 0x0
    "00000000", -- 3826 - 0xef2  :    0 - 0x0
    "11000000", -- 3827 - 0xef3  :  192 - 0xc0
    "01000000", -- 3828 - 0xef4  :   64 - 0x40
    "01011000", -- 3829 - 0xef5  :   88 - 0x58
    "01101000", -- 3830 - 0xef6  :  104 - 0x68
    "00001000", -- 3831 - 0xef7  :    8 - 0x8
    "00010000", -- 3832 - 0xef8  :   16 - 0x10 -- Background 0xdf
    "01011100", -- 3833 - 0xef9  :   92 - 0x5c
    "10101000", -- 3834 - 0xefa  :  168 - 0xa8
    "11011000", -- 3835 - 0xefb  :  216 - 0xd8
    "10111000", -- 3836 - 0xefc  :  184 - 0xb8
    "11110000", -- 3837 - 0xefd  :  240 - 0xf0
    "11100000", -- 3838 - 0xefe  :  224 - 0xe0
    "11000000", -- 3839 - 0xeff  :  192 - 0xc0
    "00000000", -- 3840 - 0xf00  :    0 - 0x0 -- Background 0xe0
    "00000000", -- 3841 - 0xf01  :    0 - 0x0
    "00000000", -- 3842 - 0xf02  :    0 - 0x0
    "00010011", -- 3843 - 0xf03  :   19 - 0x13
    "00010011", -- 3844 - 0xf04  :   19 - 0x13
    "00110111", -- 3845 - 0xf05  :   55 - 0x37
    "00110111", -- 3846 - 0xf06  :   55 - 0x37
    "00000111", -- 3847 - 0xf07  :    7 - 0x7
    "00000111", -- 3848 - 0xf08  :    7 - 0x7 -- Background 0xe1
    "00000100", -- 3849 - 0xf09  :    4 - 0x4
    "00000000", -- 3850 - 0xf0a  :    0 - 0x0
    "00000000", -- 3851 - 0xf0b  :    0 - 0x0
    "00000000", -- 3852 - 0xf0c  :    0 - 0x0
    "00100000", -- 3853 - 0xf0d  :   32 - 0x20
    "01110000", -- 3854 - 0xf0e  :  112 - 0x70
    "11111000", -- 3855 - 0xf0f  :  248 - 0xf8
    "00000000", -- 3856 - 0xf10  :    0 - 0x0 -- Background 0xe2
    "00000000", -- 3857 - 0xf11  :    0 - 0x0
    "00000000", -- 3858 - 0xf12  :    0 - 0x0
    "11111000", -- 3859 - 0xf13  :  248 - 0xf8
    "11111100", -- 3860 - 0xf14  :  252 - 0xfc
    "11111100", -- 3861 - 0xf15  :  252 - 0xfc
    "11111100", -- 3862 - 0xf16  :  252 - 0xfc
    "11111101", -- 3863 - 0xf17  :  253 - 0xfd
    "11111100", -- 3864 - 0xf18  :  252 - 0xfc -- Background 0xe3
    "00011100", -- 3865 - 0xf19  :   28 - 0x1c
    "11000000", -- 3866 - 0xf1a  :  192 - 0xc0
    "11100000", -- 3867 - 0xf1b  :  224 - 0xe0
    "00000000", -- 3868 - 0xf1c  :    0 - 0x0
    "00000000", -- 3869 - 0xf1d  :    0 - 0x0
    "00000110", -- 3870 - 0xf1e  :    6 - 0x6
    "00001111", -- 3871 - 0xf1f  :   15 - 0xf
    "00000000", -- 3872 - 0xf20  :    0 - 0x0 -- Background 0xe4
    "00000000", -- 3873 - 0xf21  :    0 - 0x0
    "00000000", -- 3874 - 0xf22  :    0 - 0x0
    "00010011", -- 3875 - 0xf23  :   19 - 0x13
    "00010011", -- 3876 - 0xf24  :   19 - 0x13
    "00110111", -- 3877 - 0xf25  :   55 - 0x37
    "00110111", -- 3878 - 0xf26  :   55 - 0x37
    "00000111", -- 3879 - 0xf27  :    7 - 0x7
    "00000111", -- 3880 - 0xf28  :    7 - 0x7 -- Background 0xe5
    "00000100", -- 3881 - 0xf29  :    4 - 0x4
    "00000001", -- 3882 - 0xf2a  :    1 - 0x1
    "00000000", -- 3883 - 0xf2b  :    0 - 0x0
    "00000000", -- 3884 - 0xf2c  :    0 - 0x0
    "00100000", -- 3885 - 0xf2d  :   32 - 0x20
    "01110000", -- 3886 - 0xf2e  :  112 - 0x70
    "11111000", -- 3887 - 0xf2f  :  248 - 0xf8
    "00000000", -- 3888 - 0xf30  :    0 - 0x0 -- Background 0xe6
    "00000000", -- 3889 - 0xf31  :    0 - 0x0
    "00000000", -- 3890 - 0xf32  :    0 - 0x0
    "11111100", -- 3891 - 0xf33  :  252 - 0xfc
    "11111100", -- 3892 - 0xf34  :  252 - 0xfc
    "11111100", -- 3893 - 0xf35  :  252 - 0xfc
    "11111100", -- 3894 - 0xf36  :  252 - 0xfc
    "11111101", -- 3895 - 0xf37  :  253 - 0xfd
    "11111100", -- 3896 - 0xf38  :  252 - 0xfc -- Background 0xe7
    "00001100", -- 3897 - 0xf39  :   12 - 0xc
    "11000000", -- 3898 - 0xf3a  :  192 - 0xc0
    "11110000", -- 3899 - 0xf3b  :  240 - 0xf0
    "11110000", -- 3900 - 0xf3c  :  240 - 0xf0
    "00000000", -- 3901 - 0xf3d  :    0 - 0x0
    "00000110", -- 3902 - 0xf3e  :    6 - 0x6
    "00001111", -- 3903 - 0xf3f  :   15 - 0xf
    "11111111", -- 3904 - 0xf40  :  255 - 0xff -- Background 0xe8
    "11111111", -- 3905 - 0xf41  :  255 - 0xff
    "01111111", -- 3906 - 0xf42  :  127 - 0x7f
    "01111111", -- 3907 - 0xf43  :  127 - 0x7f
    "01111111", -- 3908 - 0xf44  :  127 - 0x7f
    "00111111", -- 3909 - 0xf45  :   63 - 0x3f
    "00111111", -- 3910 - 0xf46  :   63 - 0x3f
    "00111111", -- 3911 - 0xf47  :   63 - 0x3f
    "00111100", -- 3912 - 0xf48  :   60 - 0x3c -- Background 0xe9
    "00111110", -- 3913 - 0xf49  :   62 - 0x3e
    "00011111", -- 3914 - 0xf4a  :   31 - 0x1f
    "00001111", -- 3915 - 0xf4b  :   15 - 0xf
    "00000111", -- 3916 - 0xf4c  :    7 - 0x7
    "00000000", -- 3917 - 0xf4d  :    0 - 0x0
    "00000000", -- 3918 - 0xf4e  :    0 - 0x0
    "00000000", -- 3919 - 0xf4f  :    0 - 0x0
    "11111111", -- 3920 - 0xf50  :  255 - 0xff -- Background 0xea
    "11111110", -- 3921 - 0xf51  :  254 - 0xfe
    "11111110", -- 3922 - 0xf52  :  254 - 0xfe
    "11111100", -- 3923 - 0xf53  :  252 - 0xfc
    "11111000", -- 3924 - 0xf54  :  248 - 0xf8
    "11110000", -- 3925 - 0xf55  :  240 - 0xf0
    "10110000", -- 3926 - 0xf56  :  176 - 0xb0
    "00111001", -- 3927 - 0xf57  :   57 - 0x39
    "00011111", -- 3928 - 0xf58  :   31 - 0x1f -- Background 0xeb
    "11001111", -- 3929 - 0xf59  :  207 - 0xcf
    "11000110", -- 3930 - 0xf5a  :  198 - 0xc6
    "10000000", -- 3931 - 0xf5b  :  128 - 0x80
    "00000000", -- 3932 - 0xf5c  :    0 - 0x0
    "00000000", -- 3933 - 0xf5d  :    0 - 0x0
    "00000000", -- 3934 - 0xf5e  :    0 - 0x0
    "00000000", -- 3935 - 0xf5f  :    0 - 0x0
    "00000000", -- 3936 - 0xf60  :    0 - 0x0 -- Background 0xec
    "00000000", -- 3937 - 0xf61  :    0 - 0x0
    "00000000", -- 3938 - 0xf62  :    0 - 0x0
    "00000000", -- 3939 - 0xf63  :    0 - 0x0
    "00000000", -- 3940 - 0xf64  :    0 - 0x0
    "00000000", -- 3941 - 0xf65  :    0 - 0x0
    "00001100", -- 3942 - 0xf66  :   12 - 0xc
    "00001100", -- 3943 - 0xf67  :   12 - 0xc
    "00110000", -- 3944 - 0xf68  :   48 - 0x30 -- Background 0xed
    "01000011", -- 3945 - 0xf69  :   67 - 0x43
    "01000000", -- 3946 - 0xf6a  :   64 - 0x40
    "01100000", -- 3947 - 0xf6b  :   96 - 0x60
    "00000011", -- 3948 - 0xf6c  :    3 - 0x3
    "00000000", -- 3949 - 0xf6d  :    0 - 0x0
    "01111111", -- 3950 - 0xf6e  :  127 - 0x7f
    "00000000", -- 3951 - 0xf6f  :    0 - 0x0
    "00000000", -- 3952 - 0xf70  :    0 - 0x0 -- Background 0xee
    "00000000", -- 3953 - 0xf71  :    0 - 0x0
    "00000000", -- 3954 - 0xf72  :    0 - 0x0
    "00000000", -- 3955 - 0xf73  :    0 - 0x0
    "00000000", -- 3956 - 0xf74  :    0 - 0x0
    "00000000", -- 3957 - 0xf75  :    0 - 0x0
    "00110000", -- 3958 - 0xf76  :   48 - 0x30
    "00110000", -- 3959 - 0xf77  :   48 - 0x30
    "00001110", -- 3960 - 0xf78  :   14 - 0xe -- Background 0xef
    "11001011", -- 3961 - 0xf79  :  203 - 0xcb
    "00000000", -- 3962 - 0xf7a  :    0 - 0x0
    "00000000", -- 3963 - 0xf7b  :    0 - 0x0
    "11000000", -- 3964 - 0xf7c  :  192 - 0xc0
    "00000000", -- 3965 - 0xf7d  :    0 - 0x0
    "11111110", -- 3966 - 0xf7e  :  254 - 0xfe
    "00000000", -- 3967 - 0xf7f  :    0 - 0x0
    "00000000", -- 3968 - 0xf80  :    0 - 0x0 -- Background 0xf0
    "00000000", -- 3969 - 0xf81  :    0 - 0x0
    "00000000", -- 3970 - 0xf82  :    0 - 0x0
    "00000000", -- 3971 - 0xf83  :    0 - 0x0
    "00000000", -- 3972 - 0xf84  :    0 - 0x0
    "00000000", -- 3973 - 0xf85  :    0 - 0x0
    "00001100", -- 3974 - 0xf86  :   12 - 0xc
    "00001100", -- 3975 - 0xf87  :   12 - 0xc
    "00110000", -- 3976 - 0xf88  :   48 - 0x30 -- Background 0xf1
    "00100011", -- 3977 - 0xf89  :   35 - 0x23
    "00100000", -- 3978 - 0xf8a  :   32 - 0x20
    "01100000", -- 3979 - 0xf8b  :   96 - 0x60
    "00000011", -- 3980 - 0xf8c  :    3 - 0x3
    "00000000", -- 3981 - 0xf8d  :    0 - 0x0
    "01111111", -- 3982 - 0xf8e  :  127 - 0x7f
    "00000000", -- 3983 - 0xf8f  :    0 - 0x0
    "00000000", -- 3984 - 0xf90  :    0 - 0x0 -- Background 0xf2
    "00000000", -- 3985 - 0xf91  :    0 - 0x0
    "00000000", -- 3986 - 0xf92  :    0 - 0x0
    "00000000", -- 3987 - 0xf93  :    0 - 0x0
    "00000000", -- 3988 - 0xf94  :    0 - 0x0
    "00000000", -- 3989 - 0xf95  :    0 - 0x0
    "00110000", -- 3990 - 0xf96  :   48 - 0x30
    "00110000", -- 3991 - 0xf97  :   48 - 0x30
    "00001001", -- 3992 - 0xf98  :    9 - 0x9 -- Background 0xf3
    "11001111", -- 3993 - 0xf99  :  207 - 0xcf
    "00000000", -- 3994 - 0xf9a  :    0 - 0x0
    "00000000", -- 3995 - 0xf9b  :    0 - 0x0
    "11000000", -- 3996 - 0xf9c  :  192 - 0xc0
    "00000000", -- 3997 - 0xf9d  :    0 - 0x0
    "11111110", -- 3998 - 0xf9e  :  254 - 0xfe
    "00000000", -- 3999 - 0xf9f  :    0 - 0x0
    "00111111", -- 4000 - 0xfa0  :   63 - 0x3f -- Background 0xf4
    "00110101", -- 4001 - 0xfa1  :   53 - 0x35
    "00011010", -- 4002 - 0xfa2  :   26 - 0x1a
    "00001101", -- 4003 - 0xfa3  :   13 - 0xd
    "00001010", -- 4004 - 0xfa4  :   10 - 0xa
    "00001101", -- 4005 - 0xfa5  :   13 - 0xd
    "00001000", -- 4006 - 0xfa6  :    8 - 0x8
    "00111000", -- 4007 - 0xfa7  :   56 - 0x38
    "01110011", -- 4008 - 0xfa8  :  115 - 0x73 -- Background 0xf5
    "11000100", -- 4009 - 0xfa9  :  196 - 0xc4
    "11000100", -- 4010 - 0xfaa  :  196 - 0xc4
    "11000000", -- 4011 - 0xfab  :  192 - 0xc0
    "11000001", -- 4012 - 0xfac  :  193 - 0xc1
    "11000000", -- 4013 - 0xfad  :  192 - 0xc0
    "01100001", -- 4014 - 0xfae  :   97 - 0x61
    "00111111", -- 4015 - 0xfaf  :   63 - 0x3f
    "11111100", -- 4016 - 0xfb0  :  252 - 0xfc -- Background 0xf6
    "01010100", -- 4017 - 0xfb1  :   84 - 0x54
    "10101000", -- 4018 - 0xfb2  :  168 - 0xa8
    "01010000", -- 4019 - 0xfb3  :   80 - 0x50
    "10110000", -- 4020 - 0xfb4  :  176 - 0xb0
    "01010000", -- 4021 - 0xfb5  :   80 - 0x50
    "10010000", -- 4022 - 0xfb6  :  144 - 0x90
    "00011100", -- 4023 - 0xfb7  :   28 - 0x1c
    "10000110", -- 4024 - 0xfb8  :  134 - 0x86 -- Background 0xf7
    "01000010", -- 4025 - 0xfb9  :   66 - 0x42
    "01000111", -- 4026 - 0xfba  :   71 - 0x47
    "01000001", -- 4027 - 0xfbb  :   65 - 0x41
    "10000011", -- 4028 - 0xfbc  :  131 - 0x83
    "00000001", -- 4029 - 0xfbd  :    1 - 0x1
    "10000110", -- 4030 - 0xfbe  :  134 - 0x86
    "11111100", -- 4031 - 0xfbf  :  252 - 0xfc
    "11100100", -- 4032 - 0xfc0  :  228 - 0xe4 -- Background 0xf8
    "11100100", -- 4033 - 0xfc1  :  228 - 0xe4
    "11101111", -- 4034 - 0xfc2  :  239 - 0xef
    "11101111", -- 4035 - 0xfc3  :  239 - 0xef
    "11111111", -- 4036 - 0xfc4  :  255 - 0xff
    "11111111", -- 4037 - 0xfc5  :  255 - 0xff
    "01111111", -- 4038 - 0xfc6  :  127 - 0x7f
    "01111111", -- 4039 - 0xfc7  :  127 - 0x7f
    "00111111", -- 4040 - 0xfc8  :   63 - 0x3f -- Background 0xf9
    "01111111", -- 4041 - 0xfc9  :  127 - 0x7f
    "01111111", -- 4042 - 0xfca  :  127 - 0x7f
    "11111111", -- 4043 - 0xfcb  :  255 - 0xff
    "11111111", -- 4044 - 0xfcc  :  255 - 0xff
    "11111111", -- 4045 - 0xfcd  :  255 - 0xff
    "11111111", -- 4046 - 0xfce  :  255 - 0xff
    "11111111", -- 4047 - 0xfcf  :  255 - 0xff
    "00010011", -- 4048 - 0xfd0  :   19 - 0x13 -- Background 0xfa
    "00010011", -- 4049 - 0xfd1  :   19 - 0x13
    "11111011", -- 4050 - 0xfd2  :  251 - 0xfb
    "11111011", -- 4051 - 0xfd3  :  251 - 0xfb
    "11111111", -- 4052 - 0xfd4  :  255 - 0xff
    "11111111", -- 4053 - 0xfd5  :  255 - 0xff
    "11111110", -- 4054 - 0xfd6  :  254 - 0xfe
    "11111110", -- 4055 - 0xfd7  :  254 - 0xfe
    "11111110", -- 4056 - 0xfd8  :  254 - 0xfe -- Background 0xfb
    "11111111", -- 4057 - 0xfd9  :  255 - 0xff
    "11111111", -- 4058 - 0xfda  :  255 - 0xff
    "11111111", -- 4059 - 0xfdb  :  255 - 0xff
    "11111111", -- 4060 - 0xfdc  :  255 - 0xff
    "11111111", -- 4061 - 0xfdd  :  255 - 0xff
    "11111111", -- 4062 - 0xfde  :  255 - 0xff
    "11111111", -- 4063 - 0xfdf  :  255 - 0xff
    "00000000", -- 4064 - 0xfe0  :    0 - 0x0 -- Background 0xfc
    "00000000", -- 4065 - 0xfe1  :    0 - 0x0
    "01111100", -- 4066 - 0xfe2  :  124 - 0x7c
    "11111110", -- 4067 - 0xfe3  :  254 - 0xfe
    "11111110", -- 4068 - 0xfe4  :  254 - 0xfe
    "01111100", -- 4069 - 0xfe5  :  124 - 0x7c
    "01000100", -- 4070 - 0xfe6  :   68 - 0x44
    "10000010", -- 4071 - 0xfe7  :  130 - 0x82
    "10000010", -- 4072 - 0xfe8  :  130 - 0x82 -- Background 0xfd
    "10000010", -- 4073 - 0xfe9  :  130 - 0x82
    "10000010", -- 4074 - 0xfea  :  130 - 0x82
    "11000110", -- 4075 - 0xfeb  :  198 - 0xc6
    "11111110", -- 4076 - 0xfec  :  254 - 0xfe
    "11111110", -- 4077 - 0xfed  :  254 - 0xfe
    "10111010", -- 4078 - 0xfee  :  186 - 0xba
    "01111100", -- 4079 - 0xfef  :  124 - 0x7c
    "00000000", -- 4080 - 0xff0  :    0 - 0x0 -- Background 0xfe
    "00011001", -- 4081 - 0xff1  :   25 - 0x19
    "00111110", -- 4082 - 0xff2  :   62 - 0x3e
    "00111100", -- 4083 - 0xff3  :   60 - 0x3c
    "00111100", -- 4084 - 0xff4  :   60 - 0x3c
    "00111100", -- 4085 - 0xff5  :   60 - 0x3c
    "00111110", -- 4086 - 0xff6  :   62 - 0x3e
    "00011001", -- 4087 - 0xff7  :   25 - 0x19
    "00000000", -- 4088 - 0xff8  :    0 - 0x0 -- Background 0xff
    "11111110", -- 4089 - 0xff9  :  254 - 0xfe
    "00011101", -- 4090 - 0xffa  :   29 - 0x1d
    "00001111", -- 4091 - 0xffb  :   15 - 0xf
    "00001111", -- 4092 - 0xffc  :   15 - 0xf
    "00001111", -- 4093 - 0xffd  :   15 - 0xf
    "00011101", -- 4094 - 0xffe  :   29 - 0x1d
    "11111110"  -- 4095 - 0xfff  :  254 - 0xfe
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
