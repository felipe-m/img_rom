--- Autcmatically generated VHDL ROM from a NES memory file----
---   NAME TABLE
-- https://wiki.nesdev.com/w/index.php/PPU_nametables
--- Only the first Name Table: 1KiB


---  Original memory dump file name: sprilo_racet4.bin --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory with clock ------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_NTABLE_SPRILO_RACE4 is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(10-1 downto 0);  --1024 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_NTABLE_SPRILO_RACE4;

architecture BEHAVIORAL of ROM_NTABLE_SPRILO_RACE4 is
  signal addr_int  : natural range 0 to 2**10-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
     ------- Name Table 0---------
    "11111010", --    0 -  0x0  :  250 - 0xfa -- line 0x0
    "11111010", --    1 -  0x1  :  250 - 0xfa
    "11101010", --    2 -  0x2  :  234 - 0xea
    "11111010", --    3 -  0x3  :  250 - 0xfa
    "11111010", --    4 -  0x4  :  250 - 0xfa
    "11111010", --    5 -  0x5  :  250 - 0xfa
    "11111010", --    6 -  0x6  :  250 - 0xfa
    "11111010", --    7 -  0x7  :  250 - 0xfa
    "11111001", --    8 -  0x8  :  249 - 0xf9
    "11111010", --    9 -  0x9  :  250 - 0xfa
    "11111010", --   10 -  0xa  :  250 - 0xfa
    "11111010", --   11 -  0xb  :  250 - 0xfa
    "11111010", --   12 -  0xc  :  250 - 0xfa
    "11111010", --   13 -  0xd  :  250 - 0xfa
    "11111010", --   14 -  0xe  :  250 - 0xfa
    "11111010", --   15 -  0xf  :  250 - 0xfa
    "11101001", --   16 - 0x10  :  233 - 0xe9
    "11111010", --   17 - 0x11  :  250 - 0xfa
    "11111010", --   18 - 0x12  :  250 - 0xfa
    "11111010", --   19 - 0x13  :  250 - 0xfa
    "11111010", --   20 - 0x14  :  250 - 0xfa
    "11111010", --   21 - 0x15  :  250 - 0xfa
    "11111010", --   22 - 0x16  :  250 - 0xfa
    "11111010", --   23 - 0x17  :  250 - 0xfa
    "11111010", --   24 - 0x18  :  250 - 0xfa
    "11111010", --   25 - 0x19  :  250 - 0xfa
    "11111010", --   26 - 0x1a  :  250 - 0xfa
    "11111010", --   27 - 0x1b  :  250 - 0xfa
    "11111010", --   28 - 0x1c  :  250 - 0xfa
    "11111010", --   29 - 0x1d  :  250 - 0xfa
    "11111010", --   30 - 0x1e  :  250 - 0xfa
    "11111010", --   31 - 0x1f  :  250 - 0xfa
    "11111010", --   32 - 0x20  :  250 - 0xfa -- line 0x1
    "11111010", --   33 - 0x21  :  250 - 0xfa
    "11111010", --   34 - 0x22  :  250 - 0xfa
    "11100111", --   35 - 0x23  :  231 - 0xe7
    "11111011", --   36 - 0x24  :  251 - 0xfb
    "11111011", --   37 - 0x25  :  251 - 0xfb
    "11111011", --   38 - 0x26  :  251 - 0xfb
    "11111011", --   39 - 0x27  :  251 - 0xfb
    "11111011", --   40 - 0x28  :  251 - 0xfb
    "11111011", --   41 - 0x29  :  251 - 0xfb
    "11111011", --   42 - 0x2a  :  251 - 0xfb
    "11111011", --   43 - 0x2b  :  251 - 0xfb
    "11111011", --   44 - 0x2c  :  251 - 0xfb
    "11111011", --   45 - 0x2d  :  251 - 0xfb
    "11111011", --   46 - 0x2e  :  251 - 0xfb
    "11111011", --   47 - 0x2f  :  251 - 0xfb
    "11111011", --   48 - 0x30  :  251 - 0xfb
    "11111011", --   49 - 0x31  :  251 - 0xfb
    "11111011", --   50 - 0x32  :  251 - 0xfb
    "11111011", --   51 - 0x33  :  251 - 0xfb
    "11111011", --   52 - 0x34  :  251 - 0xfb
    "11111011", --   53 - 0x35  :  251 - 0xfb
    "11101000", --   54 - 0x36  :  232 - 0xe8
    "11111010", --   55 - 0x37  :  250 - 0xfa
    "11111001", --   56 - 0x38  :  249 - 0xf9
    "11111010", --   57 - 0x39  :  250 - 0xfa
    "11111010", --   58 - 0x3a  :  250 - 0xfa
    "11111010", --   59 - 0x3b  :  250 - 0xfa
    "11111010", --   60 - 0x3c  :  250 - 0xfa
    "11111010", --   61 - 0x3d  :  250 - 0xfa
    "11111010", --   62 - 0x3e  :  250 - 0xfa
    "11111010", --   63 - 0x3f  :  250 - 0xfa
    "11111001", --   64 - 0x40  :  249 - 0xf9 -- line 0x2
    "11111010", --   65 - 0x41  :  250 - 0xfa
    "11111010", --   66 - 0x42  :  250 - 0xfa
    "11111100", --   67 - 0x43  :  252 - 0xfc
    "11111111", --   68 - 0x44  :  255 - 0xff
    "11111111", --   69 - 0x45  :  255 - 0xff
    "11111111", --   70 - 0x46  :  255 - 0xff
    "11111111", --   71 - 0x47  :  255 - 0xff
    "11111111", --   72 - 0x48  :  255 - 0xff
    "11111111", --   73 - 0x49  :  255 - 0xff
    "11111111", --   74 - 0x4a  :  255 - 0xff
    "11111111", --   75 - 0x4b  :  255 - 0xff
    "11111111", --   76 - 0x4c  :  255 - 0xff
    "11111111", --   77 - 0x4d  :  255 - 0xff
    "11111111", --   78 - 0x4e  :  255 - 0xff
    "11101111", --   79 - 0x4f  :  239 - 0xef
    "11111111", --   80 - 0x50  :  255 - 0xff
    "11111111", --   81 - 0x51  :  255 - 0xff
    "11111111", --   82 - 0x52  :  255 - 0xff
    "11111111", --   83 - 0x53  :  255 - 0xff
    "11111111", --   84 - 0x54  :  255 - 0xff
    "11111111", --   85 - 0x55  :  255 - 0xff
    "11101100", --   86 - 0x56  :  236 - 0xec
    "11111010", --   87 - 0x57  :  250 - 0xfa
    "11111010", --   88 - 0x58  :  250 - 0xfa
    "11111010", --   89 - 0x59  :  250 - 0xfa
    "11111010", --   90 - 0x5a  :  250 - 0xfa
    "11101010", --   91 - 0x5b  :  234 - 0xea
    "11111010", --   92 - 0x5c  :  250 - 0xfa
    "11111010", --   93 - 0x5d  :  250 - 0xfa
    "11111010", --   94 - 0x5e  :  250 - 0xfa
    "11111010", --   95 - 0x5f  :  250 - 0xfa
    "11111010", --   96 - 0x60  :  250 - 0xfa -- line 0x3
    "11111010", --   97 - 0x61  :  250 - 0xfa
    "11101001", --   98 - 0x62  :  233 - 0xe9
    "11111100", --   99 - 0x63  :  252 - 0xfc
    "11111111", --  100 - 0x64  :  255 - 0xff
    "11111111", --  101 - 0x65  :  255 - 0xff
    "11111111", --  102 - 0x66  :  255 - 0xff
    "11111101", --  103 - 0x67  :  253 - 0xfd
    "11111111", --  104 - 0x68  :  255 - 0xff
    "11111101", --  105 - 0x69  :  253 - 0xfd
    "11111111", --  106 - 0x6a  :  255 - 0xff
    "11111101", --  107 - 0x6b  :  253 - 0xfd
    "11111111", --  108 - 0x6c  :  255 - 0xff
    "11111101", --  109 - 0x6d  :  253 - 0xfd
    "11111111", --  110 - 0x6e  :  255 - 0xff
    "11101111", --  111 - 0x6f  :  239 - 0xef
    "11111111", --  112 - 0x70  :  255 - 0xff
    "11111101", --  113 - 0x71  :  253 - 0xfd
    "11111111", --  114 - 0x72  :  255 - 0xff
    "11111101", --  115 - 0x73  :  253 - 0xfd
    "11111111", --  116 - 0x74  :  255 - 0xff
    "11111111", --  117 - 0x75  :  255 - 0xff
    "11110101", --  118 - 0x76  :  245 - 0xf5
    "11111011", --  119 - 0x77  :  251 - 0xfb
    "11101000", --  120 - 0x78  :  232 - 0xe8
    "11111010", --  121 - 0x79  :  250 - 0xfa
    "11111010", --  122 - 0x7a  :  250 - 0xfa
    "11111010", --  123 - 0x7b  :  250 - 0xfa
    "11111010", --  124 - 0x7c  :  250 - 0xfa
    "11111001", --  125 - 0x7d  :  249 - 0xf9
    "11111010", --  126 - 0x7e  :  250 - 0xfa
    "11111010", --  127 - 0x7f  :  250 - 0xfa
    "11111010", --  128 - 0x80  :  250 - 0xfa -- line 0x4
    "11111010", --  129 - 0x81  :  250 - 0xfa
    "11111010", --  130 - 0x82  :  250 - 0xfa
    "11111100", --  131 - 0x83  :  252 - 0xfc
    "11111111", --  132 - 0x84  :  255 - 0xff
    "11111111", --  133 - 0x85  :  255 - 0xff
    "11111111", --  134 - 0x86  :  255 - 0xff
    "11111101", --  135 - 0x87  :  253 - 0xfd
    "11111111", --  136 - 0x88  :  255 - 0xff
    "11111101", --  137 - 0x89  :  253 - 0xfd
    "11111111", --  138 - 0x8a  :  255 - 0xff
    "11111101", --  139 - 0x8b  :  253 - 0xfd
    "11111111", --  140 - 0x8c  :  255 - 0xff
    "11111101", --  141 - 0x8d  :  253 - 0xfd
    "11111111", --  142 - 0x8e  :  255 - 0xff
    "11101111", --  143 - 0x8f  :  239 - 0xef
    "11111111", --  144 - 0x90  :  255 - 0xff
    "11111101", --  145 - 0x91  :  253 - 0xfd
    "11111111", --  146 - 0x92  :  255 - 0xff
    "11111101", --  147 - 0x93  :  253 - 0xfd
    "11111111", --  148 - 0x94  :  255 - 0xff
    "11111111", --  149 - 0x95  :  255 - 0xff
    "11111111", --  150 - 0x96  :  255 - 0xff
    "11111111", --  151 - 0x97  :  255 - 0xff
    "11101100", --  152 - 0x98  :  236 - 0xec
    "11111010", --  153 - 0x99  :  250 - 0xfa
    "11111010", --  154 - 0x9a  :  250 - 0xfa
    "11111010", --  155 - 0x9b  :  250 - 0xfa
    "11111010", --  156 - 0x9c  :  250 - 0xfa
    "11111001", --  157 - 0x9d  :  249 - 0xf9
    "11111010", --  158 - 0x9e  :  250 - 0xfa
    "11111010", --  159 - 0x9f  :  250 - 0xfa
    "11111010", --  160 - 0xa0  :  250 - 0xfa -- line 0x5
    "11111010", --  161 - 0xa1  :  250 - 0xfa
    "11111010", --  162 - 0xa2  :  250 - 0xfa
    "11111100", --  163 - 0xa3  :  252 - 0xfc
    "11111111", --  164 - 0xa4  :  255 - 0xff
    "11111111", --  165 - 0xa5  :  255 - 0xff
    "11111111", --  166 - 0xa6  :  255 - 0xff
    "11111111", --  167 - 0xa7  :  255 - 0xff
    "11111111", --  168 - 0xa8  :  255 - 0xff
    "11111111", --  169 - 0xa9  :  255 - 0xff
    "11111111", --  170 - 0xaa  :  255 - 0xff
    "11111111", --  171 - 0xab  :  255 - 0xff
    "11111111", --  172 - 0xac  :  255 - 0xff
    "11111111", --  173 - 0xad  :  255 - 0xff
    "11111111", --  174 - 0xae  :  255 - 0xff
    "11101111", --  175 - 0xaf  :  239 - 0xef
    "11111111", --  176 - 0xb0  :  255 - 0xff
    "11111111", --  177 - 0xb1  :  255 - 0xff
    "11111111", --  178 - 0xb2  :  255 - 0xff
    "11111111", --  179 - 0xb3  :  255 - 0xff
    "11111111", --  180 - 0xb4  :  255 - 0xff
    "11111111", --  181 - 0xb5  :  255 - 0xff
    "11111111", --  182 - 0xb6  :  255 - 0xff
    "11111111", --  183 - 0xb7  :  255 - 0xff
    "11101100", --  184 - 0xb8  :  236 - 0xec
    "11111010", --  185 - 0xb9  :  250 - 0xfa
    "11111010", --  186 - 0xba  :  250 - 0xfa
    "11101001", --  187 - 0xbb  :  233 - 0xe9
    "11111010", --  188 - 0xbc  :  250 - 0xfa
    "11111010", --  189 - 0xbd  :  250 - 0xfa
    "11111010", --  190 - 0xbe  :  250 - 0xfa
    "11111010", --  191 - 0xbf  :  250 - 0xfa
    "11111010", --  192 - 0xc0  :  250 - 0xfa -- line 0x6
    "11111001", --  193 - 0xc1  :  249 - 0xf9
    "11111010", --  194 - 0xc2  :  250 - 0xfa
    "11111100", --  195 - 0xc3  :  252 - 0xfc
    "11111111", --  196 - 0xc4  :  255 - 0xff
    "11111110", --  197 - 0xc5  :  254 - 0xfe
    "11111110", --  198 - 0xc6  :  254 - 0xfe
    "11111111", --  199 - 0xc7  :  255 - 0xff
    "11100101", --  200 - 0xc8  :  229 - 0xe5
    "11101011", --  201 - 0xc9  :  235 - 0xeb
    "11101011", --  202 - 0xca  :  235 - 0xeb
    "11101011", --  203 - 0xcb  :  235 - 0xeb
    "11101011", --  204 - 0xcc  :  235 - 0xeb
    "11101011", --  205 - 0xcd  :  235 - 0xeb
    "11101011", --  206 - 0xce  :  235 - 0xeb
    "11101011", --  207 - 0xcf  :  235 - 0xeb
    "11101011", --  208 - 0xd0  :  235 - 0xeb
    "11101011", --  209 - 0xd1  :  235 - 0xeb
    "11101011", --  210 - 0xd2  :  235 - 0xeb
    "11100110", --  211 - 0xd3  :  230 - 0xe6
    "11111111", --  212 - 0xd4  :  255 - 0xff
    "11111110", --  213 - 0xd5  :  254 - 0xfe
    "11111110", --  214 - 0xd6  :  254 - 0xfe
    "11111111", --  215 - 0xd7  :  255 - 0xff
    "11101100", --  216 - 0xd8  :  236 - 0xec
    "11111001", --  217 - 0xd9  :  249 - 0xf9
    "11111010", --  218 - 0xda  :  250 - 0xfa
    "11111010", --  219 - 0xdb  :  250 - 0xfa
    "11111010", --  220 - 0xdc  :  250 - 0xfa
    "11111010", --  221 - 0xdd  :  250 - 0xfa
    "11111010", --  222 - 0xde  :  250 - 0xfa
    "11111010", --  223 - 0xdf  :  250 - 0xfa
    "11111010", --  224 - 0xe0  :  250 - 0xfa -- line 0x7
    "11111010", --  225 - 0xe1  :  250 - 0xfa
    "11111010", --  226 - 0xe2  :  250 - 0xfa
    "11111100", --  227 - 0xe3  :  252 - 0xfc
    "11111111", --  228 - 0xe4  :  255 - 0xff
    "11111111", --  229 - 0xe5  :  255 - 0xff
    "11111111", --  230 - 0xe6  :  255 - 0xff
    "11111111", --  231 - 0xe7  :  255 - 0xff
    "11110101", --  232 - 0xe8  :  245 - 0xf5
    "11111011", --  233 - 0xe9  :  251 - 0xfb
    "11111011", --  234 - 0xea  :  251 - 0xfb
    "11111011", --  235 - 0xeb  :  251 - 0xfb
    "11111011", --  236 - 0xec  :  251 - 0xfb
    "11111011", --  237 - 0xed  :  251 - 0xfb
    "11111011", --  238 - 0xee  :  251 - 0xfb
    "11111011", --  239 - 0xef  :  251 - 0xfb
    "11111011", --  240 - 0xf0  :  251 - 0xfb
    "11111011", --  241 - 0xf1  :  251 - 0xfb
    "11101000", --  242 - 0xf2  :  232 - 0xe8
    "11111100", --  243 - 0xf3  :  252 - 0xfc
    "11111111", --  244 - 0xf4  :  255 - 0xff
    "11111111", --  245 - 0xf5  :  255 - 0xff
    "11111111", --  246 - 0xf6  :  255 - 0xff
    "11111111", --  247 - 0xf7  :  255 - 0xff
    "11110101", --  248 - 0xf8  :  245 - 0xf5
    "11111011", --  249 - 0xf9  :  251 - 0xfb
    "11111011", --  250 - 0xfa  :  251 - 0xfb
    "11111011", --  251 - 0xfb  :  251 - 0xfb
    "11101000", --  252 - 0xfc  :  232 - 0xe8
    "11101010", --  253 - 0xfd  :  234 - 0xea
    "11111010", --  254 - 0xfe  :  250 - 0xfa
    "11111010", --  255 - 0xff  :  250 - 0xfa
    "11111010", --  256 - 0x100  :  250 - 0xfa -- line 0x8
    "11111010", --  257 - 0x101  :  250 - 0xfa
    "11111010", --  258 - 0x102  :  250 - 0xfa
    "11111100", --  259 - 0x103  :  252 - 0xfc
    "11111111", --  260 - 0x104  :  255 - 0xff
    "11111110", --  261 - 0x105  :  254 - 0xfe
    "11111110", --  262 - 0x106  :  254 - 0xfe
    "11111111", --  263 - 0x107  :  255 - 0xff
    "11111111", --  264 - 0x108  :  255 - 0xff
    "11111111", --  265 - 0x109  :  255 - 0xff
    "11111111", --  266 - 0x10a  :  255 - 0xff
    "11111111", --  267 - 0x10b  :  255 - 0xff
    "11111111", --  268 - 0x10c  :  255 - 0xff
    "11111111", --  269 - 0x10d  :  255 - 0xff
    "11111111", --  270 - 0x10e  :  255 - 0xff
    "11111111", --  271 - 0x10f  :  255 - 0xff
    "11111111", --  272 - 0x110  :  255 - 0xff
    "11111111", --  273 - 0x111  :  255 - 0xff
    "11101100", --  274 - 0x112  :  236 - 0xec
    "11111100", --  275 - 0x113  :  252 - 0xfc
    "11111111", --  276 - 0x114  :  255 - 0xff
    "11111110", --  277 - 0x115  :  254 - 0xfe
    "11111110", --  278 - 0x116  :  254 - 0xfe
    "11111111", --  279 - 0x117  :  255 - 0xff
    "11111111", --  280 - 0x118  :  255 - 0xff
    "11111111", --  281 - 0x119  :  255 - 0xff
    "11111111", --  282 - 0x11a  :  255 - 0xff
    "11111111", --  283 - 0x11b  :  255 - 0xff
    "11101100", --  284 - 0x11c  :  236 - 0xec
    "11111010", --  285 - 0x11d  :  250 - 0xfa
    "11111010", --  286 - 0x11e  :  250 - 0xfa
    "11111010", --  287 - 0x11f  :  250 - 0xfa
    "11111010", --  288 - 0x120  :  250 - 0xfa -- line 0x9
    "11111010", --  289 - 0x121  :  250 - 0xfa
    "11101001", --  290 - 0x122  :  233 - 0xe9
    "11111100", --  291 - 0x123  :  252 - 0xfc
    "11111111", --  292 - 0x124  :  255 - 0xff
    "11111111", --  293 - 0x125  :  255 - 0xff
    "11111111", --  294 - 0x126  :  255 - 0xff
    "11111111", --  295 - 0x127  :  255 - 0xff
    "11111101", --  296 - 0x128  :  253 - 0xfd
    "11111111", --  297 - 0x129  :  255 - 0xff
    "11111101", --  298 - 0x12a  :  253 - 0xfd
    "11111111", --  299 - 0x12b  :  255 - 0xff
    "11111101", --  300 - 0x12c  :  253 - 0xfd
    "11111111", --  301 - 0x12d  :  255 - 0xff
    "11111101", --  302 - 0x12e  :  253 - 0xfd
    "11111111", --  303 - 0x12f  :  255 - 0xff
    "11111111", --  304 - 0x130  :  255 - 0xff
    "11111111", --  305 - 0x131  :  255 - 0xff
    "11101100", --  306 - 0x132  :  236 - 0xec
    "11111100", --  307 - 0x133  :  252 - 0xfc
    "11111111", --  308 - 0x134  :  255 - 0xff
    "11111111", --  309 - 0x135  :  255 - 0xff
    "11111111", --  310 - 0x136  :  255 - 0xff
    "11111111", --  311 - 0x137  :  255 - 0xff
    "11111111", --  312 - 0x138  :  255 - 0xff
    "11111101", --  313 - 0x139  :  253 - 0xfd
    "11111111", --  314 - 0x13a  :  255 - 0xff
    "11111111", --  315 - 0x13b  :  255 - 0xff
    "11101100", --  316 - 0x13c  :  236 - 0xec
    "11111010", --  317 - 0x13d  :  250 - 0xfa
    "11111010", --  318 - 0x13e  :  250 - 0xfa
    "11111001", --  319 - 0x13f  :  249 - 0xf9
    "11111010", --  320 - 0x140  :  250 - 0xfa -- line 0xa
    "11111010", --  321 - 0x141  :  250 - 0xfa
    "11111010", --  322 - 0x142  :  250 - 0xfa
    "11111100", --  323 - 0x143  :  252 - 0xfc
    "11111111", --  324 - 0x144  :  255 - 0xff
    "11111111", --  325 - 0x145  :  255 - 0xff
    "11111111", --  326 - 0x146  :  255 - 0xff
    "11111111", --  327 - 0x147  :  255 - 0xff
    "11111101", --  328 - 0x148  :  253 - 0xfd
    "11111111", --  329 - 0x149  :  255 - 0xff
    "11111101", --  330 - 0x14a  :  253 - 0xfd
    "11111111", --  331 - 0x14b  :  255 - 0xff
    "11111101", --  332 - 0x14c  :  253 - 0xfd
    "11111111", --  333 - 0x14d  :  255 - 0xff
    "11111101", --  334 - 0x14e  :  253 - 0xfd
    "11111111", --  335 - 0x14f  :  255 - 0xff
    "11111111", --  336 - 0x150  :  255 - 0xff
    "11111111", --  337 - 0x151  :  255 - 0xff
    "11101100", --  338 - 0x152  :  236 - 0xec
    "11111100", --  339 - 0x153  :  252 - 0xfc
    "11111111", --  340 - 0x154  :  255 - 0xff
    "11111111", --  341 - 0x155  :  255 - 0xff
    "11111111", --  342 - 0x156  :  255 - 0xff
    "11111111", --  343 - 0x157  :  255 - 0xff
    "11111111", --  344 - 0x158  :  255 - 0xff
    "11111101", --  345 - 0x159  :  253 - 0xfd
    "11111111", --  346 - 0x15a  :  255 - 0xff
    "11111111", --  347 - 0x15b  :  255 - 0xff
    "11101100", --  348 - 0x15c  :  236 - 0xec
    "11111010", --  349 - 0x15d  :  250 - 0xfa
    "11111010", --  350 - 0x15e  :  250 - 0xfa
    "11111010", --  351 - 0x15f  :  250 - 0xfa
    "11111010", --  352 - 0x160  :  250 - 0xfa -- line 0xb
    "11111010", --  353 - 0x161  :  250 - 0xfa
    "11111010", --  354 - 0x162  :  250 - 0xfa
    "11111100", --  355 - 0x163  :  252 - 0xfc
    "11111111", --  356 - 0x164  :  255 - 0xff
    "11111111", --  357 - 0x165  :  255 - 0xff
    "11111111", --  358 - 0x166  :  255 - 0xff
    "11111111", --  359 - 0x167  :  255 - 0xff
    "11111111", --  360 - 0x168  :  255 - 0xff
    "11111111", --  361 - 0x169  :  255 - 0xff
    "11111111", --  362 - 0x16a  :  255 - 0xff
    "11111111", --  363 - 0x16b  :  255 - 0xff
    "11111111", --  364 - 0x16c  :  255 - 0xff
    "11111111", --  365 - 0x16d  :  255 - 0xff
    "11111111", --  366 - 0x16e  :  255 - 0xff
    "11111111", --  367 - 0x16f  :  255 - 0xff
    "11111111", --  368 - 0x170  :  255 - 0xff
    "11111111", --  369 - 0x171  :  255 - 0xff
    "11101100", --  370 - 0x172  :  236 - 0xec
    "11111100", --  371 - 0x173  :  252 - 0xfc
    "11111111", --  372 - 0x174  :  255 - 0xff
    "11111111", --  373 - 0x175  :  255 - 0xff
    "11111111", --  374 - 0x176  :  255 - 0xff
    "11111111", --  375 - 0x177  :  255 - 0xff
    "11111111", --  376 - 0x178  :  255 - 0xff
    "11111111", --  377 - 0x179  :  255 - 0xff
    "11111111", --  378 - 0x17a  :  255 - 0xff
    "11111111", --  379 - 0x17b  :  255 - 0xff
    "11110101", --  380 - 0x17c  :  245 - 0xf5
    "11111011", --  381 - 0x17d  :  251 - 0xfb
    "11101000", --  382 - 0x17e  :  232 - 0xe8
    "11111010", --  383 - 0x17f  :  250 - 0xfa
    "11111010", --  384 - 0x180  :  250 - 0xfa -- line 0xc
    "11111010", --  385 - 0x181  :  250 - 0xfa
    "11111010", --  386 - 0x182  :  250 - 0xfa
    "11110111", --  387 - 0x183  :  247 - 0xf7
    "11101011", --  388 - 0x184  :  235 - 0xeb
    "11101011", --  389 - 0x185  :  235 - 0xeb
    "11101011", --  390 - 0x186  :  235 - 0xeb
    "11101011", --  391 - 0x187  :  235 - 0xeb
    "11101011", --  392 - 0x188  :  235 - 0xeb
    "11101011", --  393 - 0x189  :  235 - 0xeb
    "11101011", --  394 - 0x18a  :  235 - 0xeb
    "11101011", --  395 - 0x18b  :  235 - 0xeb
    "11101011", --  396 - 0x18c  :  235 - 0xeb
    "11100110", --  397 - 0x18d  :  230 - 0xe6
    "11111111", --  398 - 0x18e  :  255 - 0xff
    "11111111", --  399 - 0x18f  :  255 - 0xff
    "11111111", --  400 - 0x190  :  255 - 0xff
    "11111111", --  401 - 0x191  :  255 - 0xff
    "11101100", --  402 - 0x192  :  236 - 0xec
    "11110111", --  403 - 0x193  :  247 - 0xf7
    "11101011", --  404 - 0x194  :  235 - 0xeb
    "11101011", --  405 - 0x195  :  235 - 0xeb
    "11101011", --  406 - 0x196  :  235 - 0xeb
    "11100110", --  407 - 0x197  :  230 - 0xe6
    "11111111", --  408 - 0x198  :  255 - 0xff
    "11111111", --  409 - 0x199  :  255 - 0xff
    "11111111", --  410 - 0x19a  :  255 - 0xff
    "11111111", --  411 - 0x19b  :  255 - 0xff
    "11111111", --  412 - 0x19c  :  255 - 0xff
    "11111111", --  413 - 0x19d  :  255 - 0xff
    "11101100", --  414 - 0x19e  :  236 - 0xec
    "11111010", --  415 - 0x19f  :  250 - 0xfa
    "11101010", --  416 - 0x1a0  :  234 - 0xea -- line 0xd
    "11111010", --  417 - 0x1a1  :  250 - 0xfa
    "11111010", --  418 - 0x1a2  :  250 - 0xfa
    "11100111", --  419 - 0x1a3  :  231 - 0xe7
    "11111011", --  420 - 0x1a4  :  251 - 0xfb
    "11111011", --  421 - 0x1a5  :  251 - 0xfb
    "11111011", --  422 - 0x1a6  :  251 - 0xfb
    "11111011", --  423 - 0x1a7  :  251 - 0xfb
    "11111011", --  424 - 0x1a8  :  251 - 0xfb
    "11111011", --  425 - 0x1a9  :  251 - 0xfb
    "11111011", --  426 - 0x1aa  :  251 - 0xfb
    "11111011", --  427 - 0x1ab  :  251 - 0xfb
    "11111011", --  428 - 0x1ac  :  251 - 0xfb
    "11110110", --  429 - 0x1ad  :  246 - 0xf6
    "11111111", --  430 - 0x1ae  :  255 - 0xff
    "11111110", --  431 - 0x1af  :  254 - 0xfe
    "11111110", --  432 - 0x1b0  :  254 - 0xfe
    "11111111", --  433 - 0x1b1  :  255 - 0xff
    "11101100", --  434 - 0x1b2  :  236 - 0xec
    "11101001", --  435 - 0x1b3  :  233 - 0xe9
    "11111010", --  436 - 0x1b4  :  250 - 0xfa
    "11111010", --  437 - 0x1b5  :  250 - 0xfa
    "11111010", --  438 - 0x1b6  :  250 - 0xfa
    "11111100", --  439 - 0x1b7  :  252 - 0xfc
    "11111111", --  440 - 0x1b8  :  255 - 0xff
    "11111111", --  441 - 0x1b9  :  255 - 0xff
    "11111111", --  442 - 0x1ba  :  255 - 0xff
    "11111110", --  443 - 0x1bb  :  254 - 0xfe
    "11111110", --  444 - 0x1bc  :  254 - 0xfe
    "11111111", --  445 - 0x1bd  :  255 - 0xff
    "11101100", --  446 - 0x1be  :  236 - 0xec
    "11101010", --  447 - 0x1bf  :  234 - 0xea
    "11111010", --  448 - 0x1c0  :  250 - 0xfa -- line 0xe
    "11111010", --  449 - 0x1c1  :  250 - 0xfa
    "11111010", --  450 - 0x1c2  :  250 - 0xfa
    "11111100", --  451 - 0x1c3  :  252 - 0xfc
    "11111111", --  452 - 0x1c4  :  255 - 0xff
    "11111111", --  453 - 0x1c5  :  255 - 0xff
    "11111111", --  454 - 0x1c6  :  255 - 0xff
    "11111111", --  455 - 0x1c7  :  255 - 0xff
    "11111111", --  456 - 0x1c8  :  255 - 0xff
    "11111111", --  457 - 0x1c9  :  255 - 0xff
    "11111111", --  458 - 0x1ca  :  255 - 0xff
    "11111111", --  459 - 0x1cb  :  255 - 0xff
    "11111111", --  460 - 0x1cc  :  255 - 0xff
    "11111111", --  461 - 0x1cd  :  255 - 0xff
    "11111111", --  462 - 0x1ce  :  255 - 0xff
    "11111111", --  463 - 0x1cf  :  255 - 0xff
    "11111111", --  464 - 0x1d0  :  255 - 0xff
    "11111111", --  465 - 0x1d1  :  255 - 0xff
    "11101100", --  466 - 0x1d2  :  236 - 0xec
    "11111010", --  467 - 0x1d3  :  250 - 0xfa
    "11111010", --  468 - 0x1d4  :  250 - 0xfa
    "11111010", --  469 - 0x1d5  :  250 - 0xfa
    "11111010", --  470 - 0x1d6  :  250 - 0xfa
    "11110111", --  471 - 0x1d7  :  247 - 0xf7
    "11101011", --  472 - 0x1d8  :  235 - 0xeb
    "11100110", --  473 - 0x1d9  :  230 - 0xe6
    "11111111", --  474 - 0x1da  :  255 - 0xff
    "11111111", --  475 - 0x1db  :  255 - 0xff
    "11111111", --  476 - 0x1dc  :  255 - 0xff
    "11111111", --  477 - 0x1dd  :  255 - 0xff
    "11101100", --  478 - 0x1de  :  236 - 0xec
    "11111010", --  479 - 0x1df  :  250 - 0xfa
    "11111010", --  480 - 0x1e0  :  250 - 0xfa -- line 0xf
    "11111010", --  481 - 0x1e1  :  250 - 0xfa
    "11101001", --  482 - 0x1e2  :  233 - 0xe9
    "11111100", --  483 - 0x1e3  :  252 - 0xfc
    "11111111", --  484 - 0x1e4  :  255 - 0xff
    "11111111", --  485 - 0x1e5  :  255 - 0xff
    "11111111", --  486 - 0x1e6  :  255 - 0xff
    "11111111", --  487 - 0x1e7  :  255 - 0xff
    "11111101", --  488 - 0x1e8  :  253 - 0xfd
    "11111111", --  489 - 0x1e9  :  255 - 0xff
    "11111101", --  490 - 0x1ea  :  253 - 0xfd
    "11111111", --  491 - 0x1eb  :  255 - 0xff
    "11111101", --  492 - 0x1ec  :  253 - 0xfd
    "11111111", --  493 - 0x1ed  :  255 - 0xff
    "11111101", --  494 - 0x1ee  :  253 - 0xfd
    "11111111", --  495 - 0x1ef  :  255 - 0xff
    "11111111", --  496 - 0x1f0  :  255 - 0xff
    "11111111", --  497 - 0x1f1  :  255 - 0xff
    "11101100", --  498 - 0x1f2  :  236 - 0xec
    "11111010", --  499 - 0x1f3  :  250 - 0xfa
    "11111010", --  500 - 0x1f4  :  250 - 0xfa
    "11111010", --  501 - 0x1f5  :  250 - 0xfa
    "11101010", --  502 - 0x1f6  :  234 - 0xea
    "11111010", --  503 - 0x1f7  :  250 - 0xfa
    "11111010", --  504 - 0x1f8  :  250 - 0xfa
    "11111100", --  505 - 0x1f9  :  252 - 0xfc
    "11111111", --  506 - 0x1fa  :  255 - 0xff
    "11111110", --  507 - 0x1fb  :  254 - 0xfe
    "11111110", --  508 - 0x1fc  :  254 - 0xfe
    "11111111", --  509 - 0x1fd  :  255 - 0xff
    "11101100", --  510 - 0x1fe  :  236 - 0xec
    "11111010", --  511 - 0x1ff  :  250 - 0xfa
    "11111010", --  512 - 0x200  :  250 - 0xfa -- line 0x10
    "11111010", --  513 - 0x201  :  250 - 0xfa
    "11111010", --  514 - 0x202  :  250 - 0xfa
    "11111100", --  515 - 0x203  :  252 - 0xfc
    "11111111", --  516 - 0x204  :  255 - 0xff
    "11111111", --  517 - 0x205  :  255 - 0xff
    "11111111", --  518 - 0x206  :  255 - 0xff
    "11111111", --  519 - 0x207  :  255 - 0xff
    "11111101", --  520 - 0x208  :  253 - 0xfd
    "11111111", --  521 - 0x209  :  255 - 0xff
    "11111101", --  522 - 0x20a  :  253 - 0xfd
    "11111111", --  523 - 0x20b  :  255 - 0xff
    "11111101", --  524 - 0x20c  :  253 - 0xfd
    "11111111", --  525 - 0x20d  :  255 - 0xff
    "11111101", --  526 - 0x20e  :  253 - 0xfd
    "11111111", --  527 - 0x20f  :  255 - 0xff
    "11111111", --  528 - 0x210  :  255 - 0xff
    "11111111", --  529 - 0x211  :  255 - 0xff
    "11101100", --  530 - 0x212  :  236 - 0xec
    "11111010", --  531 - 0x213  :  250 - 0xfa
    "11101001", --  532 - 0x214  :  233 - 0xe9
    "11111010", --  533 - 0x215  :  250 - 0xfa
    "11111010", --  534 - 0x216  :  250 - 0xfa
    "11111010", --  535 - 0x217  :  250 - 0xfa
    "11111010", --  536 - 0x218  :  250 - 0xfa
    "11111100", --  537 - 0x219  :  252 - 0xfc
    "11111111", --  538 - 0x21a  :  255 - 0xff
    "11111111", --  539 - 0x21b  :  255 - 0xff
    "11111111", --  540 - 0x21c  :  255 - 0xff
    "11111111", --  541 - 0x21d  :  255 - 0xff
    "11101100", --  542 - 0x21e  :  236 - 0xec
    "11111001", --  543 - 0x21f  :  249 - 0xf9
    "11111010", --  544 - 0x220  :  250 - 0xfa -- line 0x11
    "11111001", --  545 - 0x221  :  249 - 0xf9
    "11111010", --  546 - 0x222  :  250 - 0xfa
    "11111100", --  547 - 0x223  :  252 - 0xfc
    "11111111", --  548 - 0x224  :  255 - 0xff
    "11111110", --  549 - 0x225  :  254 - 0xfe
    "11111110", --  550 - 0x226  :  254 - 0xfe
    "11111111", --  551 - 0x227  :  255 - 0xff
    "11111111", --  552 - 0x228  :  255 - 0xff
    "11111111", --  553 - 0x229  :  255 - 0xff
    "11111111", --  554 - 0x22a  :  255 - 0xff
    "11111111", --  555 - 0x22b  :  255 - 0xff
    "11111111", --  556 - 0x22c  :  255 - 0xff
    "11111111", --  557 - 0x22d  :  255 - 0xff
    "11111111", --  558 - 0x22e  :  255 - 0xff
    "11111111", --  559 - 0x22f  :  255 - 0xff
    "11111111", --  560 - 0x230  :  255 - 0xff
    "11111111", --  561 - 0x231  :  255 - 0xff
    "11101100", --  562 - 0x232  :  236 - 0xec
    "11111010", --  563 - 0x233  :  250 - 0xfa
    "11111010", --  564 - 0x234  :  250 - 0xfa
    "11100111", --  565 - 0x235  :  231 - 0xe7
    "11111011", --  566 - 0x236  :  251 - 0xfb
    "11111011", --  567 - 0x237  :  251 - 0xfb
    "11111011", --  568 - 0x238  :  251 - 0xfb
    "11110110", --  569 - 0x239  :  246 - 0xf6
    "11111111", --  570 - 0x23a  :  255 - 0xff
    "11111110", --  571 - 0x23b  :  254 - 0xfe
    "11111110", --  572 - 0x23c  :  254 - 0xfe
    "11111111", --  573 - 0x23d  :  255 - 0xff
    "11101100", --  574 - 0x23e  :  236 - 0xec
    "11111010", --  575 - 0x23f  :  250 - 0xfa
    "11111010", --  576 - 0x240  :  250 - 0xfa -- line 0x12
    "11111010", --  577 - 0x241  :  250 - 0xfa
    "11111010", --  578 - 0x242  :  250 - 0xfa
    "11111100", --  579 - 0x243  :  252 - 0xfc
    "11111111", --  580 - 0x244  :  255 - 0xff
    "11111111", --  581 - 0x245  :  255 - 0xff
    "11111111", --  582 - 0x246  :  255 - 0xff
    "11111111", --  583 - 0x247  :  255 - 0xff
    "11100101", --  584 - 0x248  :  229 - 0xe5
    "11101011", --  585 - 0x249  :  235 - 0xeb
    "11101011", --  586 - 0x24a  :  235 - 0xeb
    "11101011", --  587 - 0x24b  :  235 - 0xeb
    "11101011", --  588 - 0x24c  :  235 - 0xeb
    "11101011", --  589 - 0x24d  :  235 - 0xeb
    "11101011", --  590 - 0x24e  :  235 - 0xeb
    "11100110", --  591 - 0x24f  :  230 - 0xe6
    "11110100", --  592 - 0x250  :  244 - 0xf4
    "11111110", --  593 - 0x251  :  254 - 0xfe
    "11101100", --  594 - 0x252  :  236 - 0xec
    "11111010", --  595 - 0x253  :  250 - 0xfa
    "11111010", --  596 - 0x254  :  250 - 0xfa
    "11111100", --  597 - 0x255  :  252 - 0xfc
    "11111111", --  598 - 0x256  :  255 - 0xff
    "11111111", --  599 - 0x257  :  255 - 0xff
    "11111111", --  600 - 0x258  :  255 - 0xff
    "11111111", --  601 - 0x259  :  255 - 0xff
    "11111111", --  602 - 0x25a  :  255 - 0xff
    "11111111", --  603 - 0x25b  :  255 - 0xff
    "11111111", --  604 - 0x25c  :  255 - 0xff
    "11111111", --  605 - 0x25d  :  255 - 0xff
    "11101100", --  606 - 0x25e  :  236 - 0xec
    "11111010", --  607 - 0x25f  :  250 - 0xfa
    "11111010", --  608 - 0x260  :  250 - 0xfa -- line 0x13
    "11100111", --  609 - 0x261  :  231 - 0xe7
    "11111011", --  610 - 0x262  :  251 - 0xfb
    "11110110", --  611 - 0x263  :  246 - 0xf6
    "11111111", --  612 - 0x264  :  255 - 0xff
    "11111110", --  613 - 0x265  :  254 - 0xfe
    "11111110", --  614 - 0x266  :  254 - 0xfe
    "11111111", --  615 - 0x267  :  255 - 0xff
    "11101100", --  616 - 0x268  :  236 - 0xec
    "11111010", --  617 - 0x269  :  250 - 0xfa
    "11101010", --  618 - 0x26a  :  234 - 0xea
    "11111010", --  619 - 0x26b  :  250 - 0xfa
    "11111010", --  620 - 0x26c  :  250 - 0xfa
    "11111010", --  621 - 0x26d  :  250 - 0xfa
    "11111010", --  622 - 0x26e  :  250 - 0xfa
    "11111100", --  623 - 0x26f  :  252 - 0xfc
    "11111111", --  624 - 0x270  :  255 - 0xff
    "11111111", --  625 - 0x271  :  255 - 0xff
    "11101100", --  626 - 0x272  :  236 - 0xec
    "11111010", --  627 - 0x273  :  250 - 0xfa
    "11111010", --  628 - 0x274  :  250 - 0xfa
    "11111100", --  629 - 0x275  :  252 - 0xfc
    "11111111", --  630 - 0x276  :  255 - 0xff
    "11111111", --  631 - 0x277  :  255 - 0xff
    "11111111", --  632 - 0x278  :  255 - 0xff
    "11111111", --  633 - 0x279  :  255 - 0xff
    "11111101", --  634 - 0x27a  :  253 - 0xfd
    "11111111", --  635 - 0x27b  :  255 - 0xff
    "11111111", --  636 - 0x27c  :  255 - 0xff
    "11111111", --  637 - 0x27d  :  255 - 0xff
    "11101100", --  638 - 0x27e  :  236 - 0xec
    "11111010", --  639 - 0x27f  :  250 - 0xfa
    "11111010", --  640 - 0x280  :  250 - 0xfa -- line 0x14
    "11111100", --  641 - 0x281  :  252 - 0xfc
    "11111111", --  642 - 0x282  :  255 - 0xff
    "11111111", --  643 - 0x283  :  255 - 0xff
    "11111111", --  644 - 0x284  :  255 - 0xff
    "11111111", --  645 - 0x285  :  255 - 0xff
    "11111111", --  646 - 0x286  :  255 - 0xff
    "11111111", --  647 - 0x287  :  255 - 0xff
    "11101100", --  648 - 0x288  :  236 - 0xec
    "11111010", --  649 - 0x289  :  250 - 0xfa
    "11111010", --  650 - 0x28a  :  250 - 0xfa
    "11111010", --  651 - 0x28b  :  250 - 0xfa
    "11111010", --  652 - 0x28c  :  250 - 0xfa
    "11111010", --  653 - 0x28d  :  250 - 0xfa
    "11111010", --  654 - 0x28e  :  250 - 0xfa
    "11111100", --  655 - 0x28f  :  252 - 0xfc
    "11111110", --  656 - 0x290  :  254 - 0xfe
    "11110100", --  657 - 0x291  :  244 - 0xf4
    "11101100", --  658 - 0x292  :  236 - 0xec
    "11111010", --  659 - 0x293  :  250 - 0xfa
    "11111010", --  660 - 0x294  :  250 - 0xfa
    "11111100", --  661 - 0x295  :  252 - 0xfc
    "11111111", --  662 - 0x296  :  255 - 0xff
    "11111111", --  663 - 0x297  :  255 - 0xff
    "11111111", --  664 - 0x298  :  255 - 0xff
    "11111111", --  665 - 0x299  :  255 - 0xff
    "11111101", --  666 - 0x29a  :  253 - 0xfd
    "11111111", --  667 - 0x29b  :  255 - 0xff
    "11111111", --  668 - 0x29c  :  255 - 0xff
    "11111111", --  669 - 0x29d  :  255 - 0xff
    "11101100", --  670 - 0x29e  :  236 - 0xec
    "11111010", --  671 - 0x29f  :  250 - 0xfa
    "11111010", --  672 - 0x2a0  :  250 - 0xfa -- line 0x15
    "11111100", --  673 - 0x2a1  :  252 - 0xfc
    "11111111", --  674 - 0x2a2  :  255 - 0xff
    "11111111", --  675 - 0x2a3  :  255 - 0xff
    "11111111", --  676 - 0x2a4  :  255 - 0xff
    "11111111", --  677 - 0x2a5  :  255 - 0xff
    "11111111", --  678 - 0x2a6  :  255 - 0xff
    "11111111", --  679 - 0x2a7  :  255 - 0xff
    "11101100", --  680 - 0x2a8  :  236 - 0xec
    "11111010", --  681 - 0x2a9  :  250 - 0xfa
    "11111010", --  682 - 0x2aa  :  250 - 0xfa
    "11101001", --  683 - 0x2ab  :  233 - 0xe9
    "11111010", --  684 - 0x2ac  :  250 - 0xfa
    "11101010", --  685 - 0x2ad  :  234 - 0xea
    "11111010", --  686 - 0x2ae  :  250 - 0xfa
    "11111100", --  687 - 0x2af  :  252 - 0xfc
    "11111111", --  688 - 0x2b0  :  255 - 0xff
    "11111111", --  689 - 0x2b1  :  255 - 0xff
    "11101100", --  690 - 0x2b2  :  236 - 0xec
    "11111010", --  691 - 0x2b3  :  250 - 0xfa
    "11111010", --  692 - 0x2b4  :  250 - 0xfa
    "11111100", --  693 - 0x2b5  :  252 - 0xfc
    "11111111", --  694 - 0x2b6  :  255 - 0xff
    "11111110", --  695 - 0x2b7  :  254 - 0xfe
    "11111110", --  696 - 0x2b8  :  254 - 0xfe
    "11111111", --  697 - 0x2b9  :  255 - 0xff
    "11111111", --  698 - 0x2ba  :  255 - 0xff
    "11111111", --  699 - 0x2bb  :  255 - 0xff
    "11111111", --  700 - 0x2bc  :  255 - 0xff
    "11111111", --  701 - 0x2bd  :  255 - 0xff
    "11101100", --  702 - 0x2be  :  236 - 0xec
    "11111010", --  703 - 0x2bf  :  250 - 0xfa
    "11111010", --  704 - 0x2c0  :  250 - 0xfa -- line 0x16
    "11111100", --  705 - 0x2c1  :  252 - 0xfc
    "11111111", --  706 - 0x2c2  :  255 - 0xff
    "11111111", --  707 - 0x2c3  :  255 - 0xff
    "11111111", --  708 - 0x2c4  :  255 - 0xff
    "11111111", --  709 - 0x2c5  :  255 - 0xff
    "11100101", --  710 - 0x2c6  :  229 - 0xe5
    "11101011", --  711 - 0x2c7  :  235 - 0xeb
    "11111000", --  712 - 0x2c8  :  248 - 0xf8
    "11111010", --  713 - 0x2c9  :  250 - 0xfa
    "11101001", --  714 - 0x2ca  :  233 - 0xe9
    "11111010", --  715 - 0x2cb  :  250 - 0xfa
    "11111010", --  716 - 0x2cc  :  250 - 0xfa
    "11111010", --  717 - 0x2cd  :  250 - 0xfa
    "11111010", --  718 - 0x2ce  :  250 - 0xfa
    "11111100", --  719 - 0x2cf  :  252 - 0xfc
    "11110100", --  720 - 0x2d0  :  244 - 0xf4
    "11111110", --  721 - 0x2d1  :  254 - 0xfe
    "11101100", --  722 - 0x2d2  :  236 - 0xec
    "11111010", --  723 - 0x2d3  :  250 - 0xfa
    "11101010", --  724 - 0x2d4  :  234 - 0xea
    "11111100", --  725 - 0x2d5  :  252 - 0xfc
    "11111111", --  726 - 0x2d6  :  255 - 0xff
    "11111111", --  727 - 0x2d7  :  255 - 0xff
    "11111111", --  728 - 0x2d8  :  255 - 0xff
    "11111111", --  729 - 0x2d9  :  255 - 0xff
    "11100101", --  730 - 0x2da  :  229 - 0xe5
    "11101011", --  731 - 0x2db  :  235 - 0xeb
    "11101011", --  732 - 0x2dc  :  235 - 0xeb
    "11101011", --  733 - 0x2dd  :  235 - 0xeb
    "11111000", --  734 - 0x2de  :  248 - 0xf8
    "11111010", --  735 - 0x2df  :  250 - 0xfa
    "11111001", --  736 - 0x2e0  :  249 - 0xf9 -- line 0x17
    "11111100", --  737 - 0x2e1  :  252 - 0xfc
    "11111111", --  738 - 0x2e2  :  255 - 0xff
    "11111110", --  739 - 0x2e3  :  254 - 0xfe
    "11111110", --  740 - 0x2e4  :  254 - 0xfe
    "11111111", --  741 - 0x2e5  :  255 - 0xff
    "11110101", --  742 - 0x2e6  :  245 - 0xf5
    "11111011", --  743 - 0x2e7  :  251 - 0xfb
    "11111011", --  744 - 0x2e8  :  251 - 0xfb
    "11111011", --  745 - 0x2e9  :  251 - 0xfb
    "11111011", --  746 - 0x2ea  :  251 - 0xfb
    "11111011", --  747 - 0x2eb  :  251 - 0xfb
    "11111011", --  748 - 0x2ec  :  251 - 0xfb
    "11111011", --  749 - 0x2ed  :  251 - 0xfb
    "11111011", --  750 - 0x2ee  :  251 - 0xfb
    "11110110", --  751 - 0x2ef  :  246 - 0xf6
    "11110100", --  752 - 0x2f0  :  244 - 0xf4
    "11111111", --  753 - 0x2f1  :  255 - 0xff
    "11110101", --  754 - 0x2f2  :  245 - 0xf5
    "11111011", --  755 - 0x2f3  :  251 - 0xfb
    "11111011", --  756 - 0x2f4  :  251 - 0xfb
    "11110110", --  757 - 0x2f5  :  246 - 0xf6
    "11111111", --  758 - 0x2f6  :  255 - 0xff
    "11111110", --  759 - 0x2f7  :  254 - 0xfe
    "11111110", --  760 - 0x2f8  :  254 - 0xfe
    "11111111", --  761 - 0x2f9  :  255 - 0xff
    "11101100", --  762 - 0x2fa  :  236 - 0xec
    "11111010", --  763 - 0x2fb  :  250 - 0xfa
    "11111010", --  764 - 0x2fc  :  250 - 0xfa
    "11101010", --  765 - 0x2fd  :  234 - 0xea
    "11111010", --  766 - 0x2fe  :  250 - 0xfa
    "11111010", --  767 - 0x2ff  :  250 - 0xfa
    "11111001", --  768 - 0x300  :  249 - 0xf9 -- line 0x18
    "11111100", --  769 - 0x301  :  252 - 0xfc
    "11111111", --  770 - 0x302  :  255 - 0xff
    "11111111", --  771 - 0x303  :  255 - 0xff
    "11111111", --  772 - 0x304  :  255 - 0xff
    "11111111", --  773 - 0x305  :  255 - 0xff
    "11111111", --  774 - 0x306  :  255 - 0xff
    "11111111", --  775 - 0x307  :  255 - 0xff
    "11111111", --  776 - 0x308  :  255 - 0xff
    "11111111", --  777 - 0x309  :  255 - 0xff
    "11111111", --  778 - 0x30a  :  255 - 0xff
    "11111111", --  779 - 0x30b  :  255 - 0xff
    "11111111", --  780 - 0x30c  :  255 - 0xff
    "11111111", --  781 - 0x30d  :  255 - 0xff
    "11111111", --  782 - 0x30e  :  255 - 0xff
    "11111111", --  783 - 0x30f  :  255 - 0xff
    "11111111", --  784 - 0x310  :  255 - 0xff
    "11111111", --  785 - 0x311  :  255 - 0xff
    "11111111", --  786 - 0x312  :  255 - 0xff
    "11111111", --  787 - 0x313  :  255 - 0xff
    "11111111", --  788 - 0x314  :  255 - 0xff
    "11111111", --  789 - 0x315  :  255 - 0xff
    "11111111", --  790 - 0x316  :  255 - 0xff
    "11111111", --  791 - 0x317  :  255 - 0xff
    "11111111", --  792 - 0x318  :  255 - 0xff
    "11111111", --  793 - 0x319  :  255 - 0xff
    "11101100", --  794 - 0x31a  :  236 - 0xec
    "11111001", --  795 - 0x31b  :  249 - 0xf9
    "11111010", --  796 - 0x31c  :  250 - 0xfa
    "11111010", --  797 - 0x31d  :  250 - 0xfa
    "11111010", --  798 - 0x31e  :  250 - 0xfa
    "11111010", --  799 - 0x31f  :  250 - 0xfa
    "11111010", --  800 - 0x320  :  250 - 0xfa -- line 0x19
    "11111100", --  801 - 0x321  :  252 - 0xfc
    "11111111", --  802 - 0x322  :  255 - 0xff
    "11111111", --  803 - 0x323  :  255 - 0xff
    "11111111", --  804 - 0x324  :  255 - 0xff
    "11111101", --  805 - 0x325  :  253 - 0xfd
    "11111111", --  806 - 0x326  :  255 - 0xff
    "11111101", --  807 - 0x327  :  253 - 0xfd
    "11111111", --  808 - 0x328  :  255 - 0xff
    "11111101", --  809 - 0x329  :  253 - 0xfd
    "11111111", --  810 - 0x32a  :  255 - 0xff
    "11111101", --  811 - 0x32b  :  253 - 0xfd
    "11111111", --  812 - 0x32c  :  255 - 0xff
    "11111101", --  813 - 0x32d  :  253 - 0xfd
    "11111111", --  814 - 0x32e  :  255 - 0xff
    "11111111", --  815 - 0x32f  :  255 - 0xff
    "11111111", --  816 - 0x330  :  255 - 0xff
    "11111101", --  817 - 0x331  :  253 - 0xfd
    "11111111", --  818 - 0x332  :  255 - 0xff
    "11111101", --  819 - 0x333  :  253 - 0xfd
    "11111111", --  820 - 0x334  :  255 - 0xff
    "11111101", --  821 - 0x335  :  253 - 0xfd
    "11111111", --  822 - 0x336  :  255 - 0xff
    "11111110", --  823 - 0x337  :  254 - 0xfe
    "11111110", --  824 - 0x338  :  254 - 0xfe
    "11111111", --  825 - 0x339  :  255 - 0xff
    "11101100", --  826 - 0x33a  :  236 - 0xec
    "11111010", --  827 - 0x33b  :  250 - 0xfa
    "11111010", --  828 - 0x33c  :  250 - 0xfa
    "11111010", --  829 - 0x33d  :  250 - 0xfa
    "11101001", --  830 - 0x33e  :  233 - 0xe9
    "11111010", --  831 - 0x33f  :  250 - 0xfa
    "11111010", --  832 - 0x340  :  250 - 0xfa -- line 0x1a
    "11111100", --  833 - 0x341  :  252 - 0xfc
    "11111111", --  834 - 0x342  :  255 - 0xff
    "11111111", --  835 - 0x343  :  255 - 0xff
    "11111111", --  836 - 0x344  :  255 - 0xff
    "11111101", --  837 - 0x345  :  253 - 0xfd
    "11111111", --  838 - 0x346  :  255 - 0xff
    "11111101", --  839 - 0x347  :  253 - 0xfd
    "11111111", --  840 - 0x348  :  255 - 0xff
    "11111101", --  841 - 0x349  :  253 - 0xfd
    "11111111", --  842 - 0x34a  :  255 - 0xff
    "11111101", --  843 - 0x34b  :  253 - 0xfd
    "11111111", --  844 - 0x34c  :  255 - 0xff
    "11111101", --  845 - 0x34d  :  253 - 0xfd
    "11111111", --  846 - 0x34e  :  255 - 0xff
    "11111101", --  847 - 0x34f  :  253 - 0xfd
    "11111111", --  848 - 0x350  :  255 - 0xff
    "11111101", --  849 - 0x351  :  253 - 0xfd
    "11111111", --  850 - 0x352  :  255 - 0xff
    "11111101", --  851 - 0x353  :  253 - 0xfd
    "11111111", --  852 - 0x354  :  255 - 0xff
    "11111101", --  853 - 0x355  :  253 - 0xfd
    "11111111", --  854 - 0x356  :  255 - 0xff
    "11111111", --  855 - 0x357  :  255 - 0xff
    "11111111", --  856 - 0x358  :  255 - 0xff
    "11111111", --  857 - 0x359  :  255 - 0xff
    "11101100", --  858 - 0x35a  :  236 - 0xec
    "11111010", --  859 - 0x35b  :  250 - 0xfa
    "11101010", --  860 - 0x35c  :  234 - 0xea
    "11111010", --  861 - 0x35d  :  250 - 0xfa
    "11111001", --  862 - 0x35e  :  249 - 0xf9
    "11111010", --  863 - 0x35f  :  250 - 0xfa
    "11111010", --  864 - 0x360  :  250 - 0xfa -- line 0x1b
    "11111100", --  865 - 0x361  :  252 - 0xfc
    "11111111", --  866 - 0x362  :  255 - 0xff
    "11111111", --  867 - 0x363  :  255 - 0xff
    "11111111", --  868 - 0x364  :  255 - 0xff
    "11111111", --  869 - 0x365  :  255 - 0xff
    "11111111", --  870 - 0x366  :  255 - 0xff
    "11111111", --  871 - 0x367  :  255 - 0xff
    "11111111", --  872 - 0x368  :  255 - 0xff
    "11111111", --  873 - 0x369  :  255 - 0xff
    "11111111", --  874 - 0x36a  :  255 - 0xff
    "11111111", --  875 - 0x36b  :  255 - 0xff
    "11111111", --  876 - 0x36c  :  255 - 0xff
    "11111111", --  877 - 0x36d  :  255 - 0xff
    "11111111", --  878 - 0x36e  :  255 - 0xff
    "11111111", --  879 - 0x36f  :  255 - 0xff
    "11111111", --  880 - 0x370  :  255 - 0xff
    "11111111", --  881 - 0x371  :  255 - 0xff
    "11111111", --  882 - 0x372  :  255 - 0xff
    "11111111", --  883 - 0x373  :  255 - 0xff
    "11111111", --  884 - 0x374  :  255 - 0xff
    "11111111", --  885 - 0x375  :  255 - 0xff
    "11111111", --  886 - 0x376  :  255 - 0xff
    "11111111", --  887 - 0x377  :  255 - 0xff
    "11111111", --  888 - 0x378  :  255 - 0xff
    "11111111", --  889 - 0x379  :  255 - 0xff
    "11101100", --  890 - 0x37a  :  236 - 0xec
    "11111010", --  891 - 0x37b  :  250 - 0xfa
    "11111010", --  892 - 0x37c  :  250 - 0xfa
    "11111010", --  893 - 0x37d  :  250 - 0xfa
    "11111010", --  894 - 0x37e  :  250 - 0xfa
    "11111010", --  895 - 0x37f  :  250 - 0xfa
    "11111010", --  896 - 0x380  :  250 - 0xfa -- line 0x1c
    "11110111", --  897 - 0x381  :  247 - 0xf7
    "11101011", --  898 - 0x382  :  235 - 0xeb
    "11101011", --  899 - 0x383  :  235 - 0xeb
    "11101011", --  900 - 0x384  :  235 - 0xeb
    "11101011", --  901 - 0x385  :  235 - 0xeb
    "11101011", --  902 - 0x386  :  235 - 0xeb
    "11101011", --  903 - 0x387  :  235 - 0xeb
    "11101011", --  904 - 0x388  :  235 - 0xeb
    "11101011", --  905 - 0x389  :  235 - 0xeb
    "11101011", --  906 - 0x38a  :  235 - 0xeb
    "11101011", --  907 - 0x38b  :  235 - 0xeb
    "11101011", --  908 - 0x38c  :  235 - 0xeb
    "11101011", --  909 - 0x38d  :  235 - 0xeb
    "11101011", --  910 - 0x38e  :  235 - 0xeb
    "11101011", --  911 - 0x38f  :  235 - 0xeb
    "11101011", --  912 - 0x390  :  235 - 0xeb
    "11101011", --  913 - 0x391  :  235 - 0xeb
    "11101011", --  914 - 0x392  :  235 - 0xeb
    "11101011", --  915 - 0x393  :  235 - 0xeb
    "11101011", --  916 - 0x394  :  235 - 0xeb
    "11101011", --  917 - 0x395  :  235 - 0xeb
    "11101011", --  918 - 0x396  :  235 - 0xeb
    "11101011", --  919 - 0x397  :  235 - 0xeb
    "11101011", --  920 - 0x398  :  235 - 0xeb
    "11101011", --  921 - 0x399  :  235 - 0xeb
    "11111000", --  922 - 0x39a  :  248 - 0xf8
    "11111010", --  923 - 0x39b  :  250 - 0xfa
    "11111010", --  924 - 0x39c  :  250 - 0xfa
    "11101010", --  925 - 0x39d  :  234 - 0xea
    "11111010", --  926 - 0x39e  :  250 - 0xfa
    "11111001", --  927 - 0x39f  :  249 - 0xf9
    "11111010", --  928 - 0x3a0  :  250 - 0xfa -- line 0x1d
    "11111010", --  929 - 0x3a1  :  250 - 0xfa
    "11101001", --  930 - 0x3a2  :  233 - 0xe9
    "11111010", --  931 - 0x3a3  :  250 - 0xfa
    "11111010", --  932 - 0x3a4  :  250 - 0xfa
    "11111010", --  933 - 0x3a5  :  250 - 0xfa
    "11111001", --  934 - 0x3a6  :  249 - 0xf9
    "11111010", --  935 - 0x3a7  :  250 - 0xfa
    "11111010", --  936 - 0x3a8  :  250 - 0xfa
    "11111010", --  937 - 0x3a9  :  250 - 0xfa
    "11111010", --  938 - 0x3aa  :  250 - 0xfa
    "11111010", --  939 - 0x3ab  :  250 - 0xfa
    "11111010", --  940 - 0x3ac  :  250 - 0xfa
    "11111010", --  941 - 0x3ad  :  250 - 0xfa
    "11111010", --  942 - 0x3ae  :  250 - 0xfa
    "11111010", --  943 - 0x3af  :  250 - 0xfa
    "11101010", --  944 - 0x3b0  :  234 - 0xea
    "11111010", --  945 - 0x3b1  :  250 - 0xfa
    "11111010", --  946 - 0x3b2  :  250 - 0xfa
    "11111010", --  947 - 0x3b3  :  250 - 0xfa
    "11111010", --  948 - 0x3b4  :  250 - 0xfa
    "11111001", --  949 - 0x3b5  :  249 - 0xf9
    "11111010", --  950 - 0x3b6  :  250 - 0xfa
    "11111010", --  951 - 0x3b7  :  250 - 0xfa
    "11111010", --  952 - 0x3b8  :  250 - 0xfa
    "11111010", --  953 - 0x3b9  :  250 - 0xfa
    "11111010", --  954 - 0x3ba  :  250 - 0xfa
    "11111001", --  955 - 0x3bb  :  249 - 0xf9
    "11111010", --  956 - 0x3bc  :  250 - 0xfa
    "11111010", --  957 - 0x3bd  :  250 - 0xfa
    "11111010", --  958 - 0x3be  :  250 - 0xfa
    "11111010", --  959 - 0x3bf  :  250 - 0xfa
        ---- Attribute Table 0----
    "01010101", --  960 - 0x3c0  :   85 - 0x55
    "00000101", --  961 - 0x3c1  :    5 - 0x5
    "00000101", --  962 - 0x3c2  :    5 - 0x5
    "00000101", --  963 - 0x3c3  :    5 - 0x5
    "00000101", --  964 - 0x3c4  :    5 - 0x5
    "01000101", --  965 - 0x3c5  :   69 - 0x45
    "01010101", --  966 - 0x3c6  :   85 - 0x55
    "01010101", --  967 - 0x3c7  :   85 - 0x55
    "01010101", --  968 - 0x3c8  :   85 - 0x55
    "00000000", --  969 - 0x3c9  :    0 - 0x0
    "01010000", --  970 - 0x3ca  :   80 - 0x50
    "01010000", --  971 - 0x3cb  :   80 - 0x50
    "01010000", --  972 - 0x3cc  :   80 - 0x50
    "00000000", --  973 - 0x3cd  :    0 - 0x0
    "01010101", --  974 - 0x3ce  :   85 - 0x55
    "01010101", --  975 - 0x3cf  :   85 - 0x55
    "01010101", --  976 - 0x3d0  :   85 - 0x55
    "00000000", --  977 - 0x3d1  :    0 - 0x0
    "00000000", --  978 - 0x3d2  :    0 - 0x0
    "00000000", --  979 - 0x3d3  :    0 - 0x0
    "01000100", --  980 - 0x3d4  :   68 - 0x44
    "00000000", --  981 - 0x3d5  :    0 - 0x0
    "00000000", --  982 - 0x3d6  :    0 - 0x0
    "01010101", --  983 - 0x3d7  :   85 - 0x55
    "01010101", --  984 - 0x3d8  :   85 - 0x55
    "00000101", --  985 - 0x3d9  :    5 - 0x5
    "00000101", --  986 - 0x3da  :    5 - 0x5
    "00000001", --  987 - 0x3db  :    1 - 0x1
    "01000100", --  988 - 0x3dc  :   68 - 0x44
    "01010101", --  989 - 0x3dd  :   85 - 0x55
    "00010000", --  990 - 0x3de  :   16 - 0x10
    "01000100", --  991 - 0x3df  :   68 - 0x44
    "01010101", --  992 - 0x3e0  :   85 - 0x55
    "00000000", --  993 - 0x3e1  :    0 - 0x0
    "01010000", --  994 - 0x3e2  :   80 - 0x50
    "01010000", --  995 - 0x3e3  :   80 - 0x50
    "01000100", --  996 - 0x3e4  :   68 - 0x44
    "00010101", --  997 - 0x3e5  :   21 - 0x15
    "00000001", --  998 - 0x3e6  :    1 - 0x1
    "01000100", --  999 - 0x3e7  :   68 - 0x44
    "00010001", -- 1000 - 0x3e8  :   17 - 0x11
    "01000000", -- 1001 - 0x3e9  :   64 - 0x40
    "01010101", -- 1002 - 0x3ea  :   85 - 0x55
    "01010101", -- 1003 - 0x3eb  :   85 - 0x55
    "01000100", -- 1004 - 0x3ec  :   68 - 0x44
    "00010001", -- 1005 - 0x3ed  :   17 - 0x11
    "01000000", -- 1006 - 0x3ee  :   64 - 0x40
    "01010100", -- 1007 - 0x3ef  :   84 - 0x54
    "00010001", -- 1008 - 0x3f0  :   17 - 0x11
    "00000000", -- 1009 - 0x3f1  :    0 - 0x0
    "00000000", -- 1010 - 0x3f2  :    0 - 0x0
    "00000000", -- 1011 - 0x3f3  :    0 - 0x0
    "00000000", -- 1012 - 0x3f4  :    0 - 0x0
    "00000000", -- 1013 - 0x3f5  :    0 - 0x0
    "01000100", -- 1014 - 0x3f6  :   68 - 0x44
    "01010101", -- 1015 - 0x3f7  :   85 - 0x55
    "00000101", -- 1016 - 0x3f8  :    5 - 0x5
    "00000101", -- 1017 - 0x3f9  :    5 - 0x5
    "00000101", -- 1018 - 0x3fa  :    5 - 0x5
    "00000101", -- 1019 - 0x3fb  :    5 - 0x5
    "00000101", -- 1020 - 0x3fc  :    5 - 0x5
    "00000101", -- 1021 - 0x3fd  :    5 - 0x5
    "00000101", -- 1022 - 0x3fe  :    5 - 0x5
    "00000101"  -- 1023 - 0x3ff  :    5 - 0x5
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
