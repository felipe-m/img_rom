---   Sprites Pattern table BOTH COLOR PLANES
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
--- Autcmatically generated VHDL ROM from a NES memory file----


---  Original memory dump file name: lawnmower_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory with clock ------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_LAWN_SPR is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(12-1 downto 0);  --4096 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_LAWN_SPR;

architecture BEHAVIORAL of ROM_PTABLE_LAWN_SPR is
  signal addr_int  : natural range 0 to 2**12-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Sprite pattern Table both color planes
    "11111111", --    0 -  0x0  :  255 - 0xff -- Sprite 0x0
    "11111111", --    1 -  0x1  :  255 - 0xff
    "11111111", --    2 -  0x2  :  255 - 0xff
    "11111111", --    3 -  0x3  :  255 - 0xff
    "11111111", --    4 -  0x4  :  255 - 0xff
    "11111111", --    5 -  0x5  :  255 - 0xff
    "11111111", --    6 -  0x6  :  255 - 0xff
    "11111111", --    7 -  0x7  :  255 - 0xff
    "00000000", --    8 -  0x8  :    0 - 0x0 -- plane 1
    "00000000", --    9 -  0x9  :    0 - 0x0
    "00000000", --   10 -  0xa  :    0 - 0x0
    "00000000", --   11 -  0xb  :    0 - 0x0
    "00000000", --   12 -  0xc  :    0 - 0x0
    "00000000", --   13 -  0xd  :    0 - 0x0
    "00000000", --   14 -  0xe  :    0 - 0x0
    "00000000", --   15 -  0xf  :    0 - 0x0
    "11111111", --   16 - 0x10  :  255 - 0xff -- Sprite 0x1
    "11111111", --   17 - 0x11  :  255 - 0xff
    "11111111", --   18 - 0x12  :  255 - 0xff
    "11111111", --   19 - 0x13  :  255 - 0xff
    "11111111", --   20 - 0x14  :  255 - 0xff
    "11111111", --   21 - 0x15  :  255 - 0xff
    "11111100", --   22 - 0x16  :  252 - 0xfc
    "11111100", --   23 - 0x17  :  252 - 0xfc
    "00000000", --   24 - 0x18  :    0 - 0x0 -- plane 1
    "00000000", --   25 - 0x19  :    0 - 0x0
    "00000000", --   26 - 0x1a  :    0 - 0x0
    "00000000", --   27 - 0x1b  :    0 - 0x0
    "00000000", --   28 - 0x1c  :    0 - 0x0
    "00000111", --   29 - 0x1d  :    7 - 0x7
    "00000111", --   30 - 0x1e  :    7 - 0x7
    "00000110", --   31 - 0x1f  :    6 - 0x6
    "11111111", --   32 - 0x20  :  255 - 0xff -- Sprite 0x2
    "11111111", --   33 - 0x21  :  255 - 0xff
    "11111111", --   34 - 0x22  :  255 - 0xff
    "11111111", --   35 - 0x23  :  255 - 0xff
    "11111111", --   36 - 0x24  :  255 - 0xff
    "11111111", --   37 - 0x25  :  255 - 0xff
    "00000000", --   38 - 0x26  :    0 - 0x0
    "00000000", --   39 - 0x27  :    0 - 0x0
    "00000000", --   40 - 0x28  :    0 - 0x0 -- plane 1
    "00000000", --   41 - 0x29  :    0 - 0x0
    "00000000", --   42 - 0x2a  :    0 - 0x0
    "00000000", --   43 - 0x2b  :    0 - 0x0
    "00000000", --   44 - 0x2c  :    0 - 0x0
    "11111111", --   45 - 0x2d  :  255 - 0xff
    "11111111", --   46 - 0x2e  :  255 - 0xff
    "00000000", --   47 - 0x2f  :    0 - 0x0
    "11111111", --   48 - 0x30  :  255 - 0xff -- Sprite 0x3
    "11111111", --   49 - 0x31  :  255 - 0xff
    "11111111", --   50 - 0x32  :  255 - 0xff
    "11111111", --   51 - 0x33  :  255 - 0xff
    "11111111", --   52 - 0x34  :  255 - 0xff
    "11111111", --   53 - 0x35  :  255 - 0xff
    "00011111", --   54 - 0x36  :   31 - 0x1f
    "01000111", --   55 - 0x37  :   71 - 0x47
    "00000000", --   56 - 0x38  :    0 - 0x0 -- plane 1
    "00000000", --   57 - 0x39  :    0 - 0x0
    "00000000", --   58 - 0x3a  :    0 - 0x0
    "00000000", --   59 - 0x3b  :    0 - 0x0
    "00000000", --   60 - 0x3c  :    0 - 0x0
    "11100000", --   61 - 0x3d  :  224 - 0xe0
    "11100000", --   62 - 0x3e  :  224 - 0xe0
    "01100000", --   63 - 0x3f  :   96 - 0x60
    "11111111", --   64 - 0x40  :  255 - 0xff -- Sprite 0x4
    "11111111", --   65 - 0x41  :  255 - 0xff
    "11111111", --   66 - 0x42  :  255 - 0xff
    "11111111", --   67 - 0x43  :  255 - 0xff
    "11111111", --   68 - 0x44  :  255 - 0xff
    "11111111", --   69 - 0x45  :  255 - 0xff
    "11100000", --   70 - 0x46  :  224 - 0xe0
    "10000000", --   71 - 0x47  :  128 - 0x80
    "00000000", --   72 - 0x48  :    0 - 0x0 -- plane 1
    "00000000", --   73 - 0x49  :    0 - 0x0
    "00000000", --   74 - 0x4a  :    0 - 0x0
    "00000000", --   75 - 0x4b  :    0 - 0x0
    "00000000", --   76 - 0x4c  :    0 - 0x0
    "00011111", --   77 - 0x4d  :   31 - 0x1f
    "01111111", --   78 - 0x4e  :  127 - 0x7f
    "11110000", --   79 - 0x4f  :  240 - 0xf0
    "11111111", --   80 - 0x50  :  255 - 0xff -- Sprite 0x5
    "11111111", --   81 - 0x51  :  255 - 0xff
    "11111111", --   82 - 0x52  :  255 - 0xff
    "11111111", --   83 - 0x53  :  255 - 0xff
    "11111111", --   84 - 0x54  :  255 - 0xff
    "11110111", --   85 - 0x55  :  247 - 0xf7
    "00000001", --   86 - 0x56  :    1 - 0x1
    "00000100", --   87 - 0x57  :    4 - 0x4
    "00000000", --   88 - 0x58  :    0 - 0x0 -- plane 1
    "00000000", --   89 - 0x59  :    0 - 0x0
    "00000000", --   90 - 0x5a  :    0 - 0x0
    "00000000", --   91 - 0x5b  :    0 - 0x0
    "00000000", --   92 - 0x5c  :    0 - 0x0
    "11111000", --   93 - 0x5d  :  248 - 0xf8
    "11111110", --   94 - 0x5e  :  254 - 0xfe
    "00001111", --   95 - 0x5f  :   15 - 0xf
    "11111111", --   96 - 0x60  :  255 - 0xff -- Sprite 0x6
    "11111111", --   97 - 0x61  :  255 - 0xff
    "11111111", --   98 - 0x62  :  255 - 0xff
    "11111111", --   99 - 0x63  :  255 - 0xff
    "11111111", --  100 - 0x64  :  255 - 0xff
    "11011111", --  101 - 0x65  :  223 - 0xdf
    "00011100", --  102 - 0x66  :   28 - 0x1c
    "01000100", --  103 - 0x67  :   68 - 0x44
    "00000000", --  104 - 0x68  :    0 - 0x0 -- plane 1
    "00000000", --  105 - 0x69  :    0 - 0x0
    "00000000", --  106 - 0x6a  :    0 - 0x0
    "00000000", --  107 - 0x6b  :    0 - 0x0
    "00000000", --  108 - 0x6c  :    0 - 0x0
    "11100111", --  109 - 0x6d  :  231 - 0xe7
    "11100111", --  110 - 0x6e  :  231 - 0xe7
    "01100110", --  111 - 0x6f  :  102 - 0x66
    "11111111", --  112 - 0x70  :  255 - 0xff -- Sprite 0x7
    "11111111", --  113 - 0x71  :  255 - 0xff
    "11111111", --  114 - 0x72  :  255 - 0xff
    "11111111", --  115 - 0x73  :  255 - 0xff
    "11111111", --  116 - 0x74  :  255 - 0xff
    "10111111", --  117 - 0x75  :  191 - 0xbf
    "00111100", --  118 - 0x76  :   60 - 0x3c
    "01001100", --  119 - 0x77  :   76 - 0x4c
    "00000000", --  120 - 0x78  :    0 - 0x0 -- plane 1
    "00000000", --  121 - 0x79  :    0 - 0x0
    "00000000", --  122 - 0x7a  :    0 - 0x0
    "00000000", --  123 - 0x7b  :    0 - 0x0
    "00000000", --  124 - 0x7c  :    0 - 0x0
    "11000111", --  125 - 0x7d  :  199 - 0xc7
    "11000111", --  126 - 0x7e  :  199 - 0xc7
    "01100110", --  127 - 0x7f  :  102 - 0x66
    "11111100", --  128 - 0x80  :  252 - 0xfc -- Sprite 0x8
    "11111100", --  129 - 0x81  :  252 - 0xfc
    "11111100", --  130 - 0x82  :  252 - 0xfc
    "11111100", --  131 - 0x83  :  252 - 0xfc
    "11111100", --  132 - 0x84  :  252 - 0xfc
    "11111100", --  133 - 0x85  :  252 - 0xfc
    "11111100", --  134 - 0x86  :  252 - 0xfc
    "11111100", --  135 - 0x87  :  252 - 0xfc
    "00000110", --  136 - 0x88  :    6 - 0x6 -- plane 1
    "00000110", --  137 - 0x89  :    6 - 0x6
    "00000110", --  138 - 0x8a  :    6 - 0x6
    "00000110", --  139 - 0x8b  :    6 - 0x6
    "00000110", --  140 - 0x8c  :    6 - 0x6
    "00000110", --  141 - 0x8d  :    6 - 0x6
    "00000110", --  142 - 0x8e  :    6 - 0x6
    "00000110", --  143 - 0x8f  :    6 - 0x6
    "00010000", --  144 - 0x90  :   16 - 0x10 -- Sprite 0x9
    "00111000", --  145 - 0x91  :   56 - 0x38
    "01111100", --  146 - 0x92  :  124 - 0x7c
    "11111000", --  147 - 0x93  :  248 - 0xf8
    "01110000", --  148 - 0x94  :  112 - 0x70
    "00100010", --  149 - 0x95  :   34 - 0x22
    "00000101", --  150 - 0x96  :    5 - 0x5
    "00000010", --  151 - 0x97  :    2 - 0x2
    "11111111", --  152 - 0x98  :  255 - 0xff -- plane 1
    "11111111", --  153 - 0x99  :  255 - 0xff
    "11111111", --  154 - 0x9a  :  255 - 0xff
    "11111111", --  155 - 0x9b  :  255 - 0xff
    "11111111", --  156 - 0x9c  :  255 - 0xff
    "11111111", --  157 - 0x9d  :  255 - 0xff
    "11111111", --  158 - 0x9e  :  255 - 0xff
    "11111111", --  159 - 0x9f  :  255 - 0xff
    "01000111", --  160 - 0xa0  :   71 - 0x47 -- Sprite 0xa
    "01000111", --  161 - 0xa1  :   71 - 0x47
    "01000111", --  162 - 0xa2  :   71 - 0x47
    "01000111", --  163 - 0xa3  :   71 - 0x47
    "01000111", --  164 - 0xa4  :   71 - 0x47
    "01000111", --  165 - 0xa5  :   71 - 0x47
    "01000111", --  166 - 0xa6  :   71 - 0x47
    "01000111", --  167 - 0xa7  :   71 - 0x47
    "01100000", --  168 - 0xa8  :   96 - 0x60 -- plane 1
    "01100000", --  169 - 0xa9  :   96 - 0x60
    "01100000", --  170 - 0xaa  :   96 - 0x60
    "01100000", --  171 - 0xab  :   96 - 0x60
    "01100000", --  172 - 0xac  :   96 - 0x60
    "01100000", --  173 - 0xad  :   96 - 0x60
    "01100000", --  174 - 0xae  :   96 - 0x60
    "01100000", --  175 - 0xaf  :   96 - 0x60
    "11111111", --  176 - 0xb0  :  255 - 0xff -- Sprite 0xb
    "11111110", --  177 - 0xb1  :  254 - 0xfe
    "11111110", --  178 - 0xb2  :  254 - 0xfe
    "11111100", --  179 - 0xb3  :  252 - 0xfc
    "11111100", --  180 - 0xb4  :  252 - 0xfc
    "11111100", --  181 - 0xb5  :  252 - 0xfc
    "11111100", --  182 - 0xb6  :  252 - 0xfc
    "11111100", --  183 - 0xb7  :  252 - 0xfc
    "00000001", --  184 - 0xb8  :    1 - 0x1 -- plane 1
    "00000011", --  185 - 0xb9  :    3 - 0x3
    "00000011", --  186 - 0xba  :    3 - 0x3
    "00000111", --  187 - 0xbb  :    7 - 0x7
    "00000110", --  188 - 0xbc  :    6 - 0x6
    "00000110", --  189 - 0xbd  :    6 - 0x6
    "00000110", --  190 - 0xbe  :    6 - 0x6
    "00000110", --  191 - 0xbf  :    6 - 0x6
    "00000000", --  192 - 0xc0  :    0 - 0x0 -- Sprite 0xc
    "00001000", --  193 - 0xc1  :    8 - 0x8
    "00011100", --  194 - 0xc2  :   28 - 0x1c
    "00111000", --  195 - 0xc3  :   56 - 0x38
    "01110000", --  196 - 0xc4  :  112 - 0x70
    "00100010", --  197 - 0xc5  :   34 - 0x22
    "00000101", --  198 - 0xc6  :    5 - 0x5
    "00000010", --  199 - 0xc7  :    2 - 0x2
    "11000111", --  200 - 0xc8  :  199 - 0xc7 -- plane 1
    "10011111", --  201 - 0xc9  :  159 - 0x9f
    "00111111", --  202 - 0xca  :   63 - 0x3f
    "01111111", --  203 - 0xcb  :  127 - 0x7f
    "01111111", --  204 - 0xcc  :  127 - 0x7f
    "11111111", --  205 - 0xcd  :  255 - 0xff
    "11111111", --  206 - 0xce  :  255 - 0xff
    "11111111", --  207 - 0xcf  :  255 - 0xff
    "00000010", --  208 - 0xd0  :    2 - 0x2 -- Sprite 0xd
    "00110001", --  209 - 0xd1  :   49 - 0x31
    "01111000", --  210 - 0xd2  :  120 - 0x78
    "11111000", --  211 - 0xd3  :  248 - 0xf8
    "01110000", --  212 - 0xd4  :  112 - 0x70
    "00100010", --  213 - 0xd5  :   34 - 0x22
    "00000101", --  214 - 0xd6  :    5 - 0x5
    "00000010", --  215 - 0xd7  :    2 - 0x2
    "11100011", --  216 - 0xd8  :  227 - 0xe3 -- plane 1
    "11111001", --  217 - 0xd9  :  249 - 0xf9
    "11111100", --  218 - 0xda  :  252 - 0xfc
    "11111110", --  219 - 0xdb  :  254 - 0xfe
    "11111110", --  220 - 0xdc  :  254 - 0xfe
    "11111111", --  221 - 0xdd  :  255 - 0xff
    "11111111", --  222 - 0xde  :  255 - 0xff
    "11111111", --  223 - 0xdf  :  255 - 0xff
    "01111100", --  224 - 0xe0  :  124 - 0x7c -- Sprite 0xe
    "00111100", --  225 - 0xe1  :   60 - 0x3c
    "10011100", --  226 - 0xe2  :  156 - 0x9c
    "10001100", --  227 - 0xe3  :  140 - 0x8c
    "01001100", --  228 - 0xe4  :   76 - 0x4c
    "01000100", --  229 - 0xe5  :   68 - 0x44
    "01000100", --  230 - 0xe6  :   68 - 0x44
    "01000100", --  231 - 0xe7  :   68 - 0x44
    "10000110", --  232 - 0xe8  :  134 - 0x86 -- plane 1
    "11000110", --  233 - 0xe9  :  198 - 0xc6
    "11000110", --  234 - 0xea  :  198 - 0xc6
    "11100110", --  235 - 0xeb  :  230 - 0xe6
    "01100110", --  236 - 0xec  :  102 - 0x66
    "01100110", --  237 - 0xed  :  102 - 0x66
    "01100110", --  238 - 0xee  :  102 - 0x66
    "01100110", --  239 - 0xef  :  102 - 0x66
    "01000100", --  240 - 0xf0  :   68 - 0x44 -- Sprite 0xf
    "01000100", --  241 - 0xf1  :   68 - 0x44
    "01000100", --  242 - 0xf2  :   68 - 0x44
    "01000100", --  243 - 0xf3  :   68 - 0x44
    "01000100", --  244 - 0xf4  :   68 - 0x44
    "01000100", --  245 - 0xf5  :   68 - 0x44
    "01000100", --  246 - 0xf6  :   68 - 0x44
    "01000100", --  247 - 0xf7  :   68 - 0x44
    "01100110", --  248 - 0xf8  :  102 - 0x66 -- plane 1
    "01100110", --  249 - 0xf9  :  102 - 0x66
    "01100110", --  250 - 0xfa  :  102 - 0x66
    "01100110", --  251 - 0xfb  :  102 - 0x66
    "01100110", --  252 - 0xfc  :  102 - 0x66
    "01100110", --  253 - 0xfd  :  102 - 0x66
    "01100110", --  254 - 0xfe  :  102 - 0x66
    "01100110", --  255 - 0xff  :  102 - 0x66
    "01001100", --  256 - 0x100  :   76 - 0x4c -- Sprite 0x10
    "00100100", --  257 - 0x101  :   36 - 0x24
    "00100100", --  258 - 0x102  :   36 - 0x24
    "10010100", --  259 - 0x103  :  148 - 0x94
    "00010000", --  260 - 0x104  :   16 - 0x10
    "00001000", --  261 - 0x105  :    8 - 0x8
    "00001000", --  262 - 0x106  :    8 - 0x8
    "00000100", --  263 - 0x107  :    4 - 0x4
    "01100110", --  264 - 0x108  :  102 - 0x66 -- plane 1
    "00110110", --  265 - 0x109  :   54 - 0x36
    "10110110", --  266 - 0x10a  :  182 - 0xb6
    "10011110", --  267 - 0x10b  :  158 - 0x9e
    "11011110", --  268 - 0x10c  :  222 - 0xde
    "11001110", --  269 - 0x10d  :  206 - 0xce
    "11101110", --  270 - 0x10e  :  238 - 0xee
    "11100110", --  271 - 0x10f  :  230 - 0xe6
    "00000000", --  272 - 0x110  :    0 - 0x0 -- Sprite 0x11
    "00111100", --  273 - 0x111  :   60 - 0x3c
    "01000000", --  274 - 0x112  :   64 - 0x40
    "01000100", --  275 - 0x113  :   68 - 0x44
    "01000100", --  276 - 0x114  :   68 - 0x44
    "01000100", --  277 - 0x115  :   68 - 0x44
    "01000100", --  278 - 0x116  :   68 - 0x44
    "01000100", --  279 - 0x117  :   68 - 0x44
    "10000001", --  280 - 0x118  :  129 - 0x81 -- plane 1
    "00111100", --  281 - 0x119  :   60 - 0x3c
    "01111110", --  282 - 0x11a  :  126 - 0x7e
    "01100110", --  283 - 0x11b  :  102 - 0x66
    "01100110", --  284 - 0x11c  :  102 - 0x66
    "01100110", --  285 - 0x11d  :  102 - 0x66
    "01100110", --  286 - 0x11e  :  102 - 0x66
    "01100110", --  287 - 0x11f  :  102 - 0x66
    "00000100", --  288 - 0x120  :    4 - 0x4 -- Sprite 0x12
    "00010010", --  289 - 0x121  :   18 - 0x12
    "00110010", --  290 - 0x122  :   50 - 0x32
    "01111000", --  291 - 0x123  :  120 - 0x78
    "11111000", --  292 - 0x124  :  248 - 0xf8
    "01110000", --  293 - 0x125  :  112 - 0x70
    "00100100", --  294 - 0x126  :   36 - 0x24
    "00000000", --  295 - 0x127  :    0 - 0x0
    "11110110", --  296 - 0x128  :  246 - 0xf6 -- plane 1
    "11110010", --  297 - 0x129  :  242 - 0xf2
    "11111010", --  298 - 0x12a  :  250 - 0xfa
    "11111000", --  299 - 0x12b  :  248 - 0xf8
    "11111100", --  300 - 0x12c  :  252 - 0xfc
    "11111100", --  301 - 0x12d  :  252 - 0xfc
    "11111110", --  302 - 0x12e  :  254 - 0xfe
    "11111110", --  303 - 0x12f  :  254 - 0xfe
    "01000100", --  304 - 0x130  :   68 - 0x44 -- Sprite 0x13
    "01000100", --  305 - 0x131  :   68 - 0x44
    "01000100", --  306 - 0x132  :   68 - 0x44
    "01000100", --  307 - 0x133  :   68 - 0x44
    "01000100", --  308 - 0x134  :   68 - 0x44
    "01000100", --  309 - 0x135  :   68 - 0x44
    "01000100", --  310 - 0x136  :   68 - 0x44
    "01011100", --  311 - 0x137  :   92 - 0x5c
    "01100110", --  312 - 0x138  :  102 - 0x66 -- plane 1
    "01100110", --  313 - 0x139  :  102 - 0x66
    "01100110", --  314 - 0x13a  :  102 - 0x66
    "01100110", --  315 - 0x13b  :  102 - 0x66
    "01100110", --  316 - 0x13c  :  102 - 0x66
    "01100110", --  317 - 0x13d  :  102 - 0x66
    "01100110", --  318 - 0x13e  :  102 - 0x66
    "01111110", --  319 - 0x13f  :  126 - 0x7e
    "00010000", --  320 - 0x140  :   16 - 0x10 -- Sprite 0x14
    "00111000", --  321 - 0x141  :   56 - 0x38
    "00111100", --  322 - 0x142  :   60 - 0x3c
    "00111000", --  323 - 0x143  :   56 - 0x38
    "00010000", --  324 - 0x144  :   16 - 0x10
    "00000010", --  325 - 0x145  :    2 - 0x2
    "01000101", --  326 - 0x146  :   69 - 0x45
    "01000010", --  327 - 0x147  :   66 - 0x42
    "11111111", --  328 - 0x148  :  255 - 0xff -- plane 1
    "01111111", --  329 - 0x149  :  127 - 0x7f
    "01111111", --  330 - 0x14a  :  127 - 0x7f
    "00111111", --  331 - 0x14b  :   63 - 0x3f
    "00111111", --  332 - 0x14c  :   63 - 0x3f
    "00011111", --  333 - 0x14d  :   31 - 0x1f
    "01011111", --  334 - 0x14e  :   95 - 0x5f
    "01001111", --  335 - 0x14f  :   79 - 0x4f
    "01000100", --  336 - 0x150  :   68 - 0x44 -- Sprite 0x15
    "01000100", --  337 - 0x151  :   68 - 0x44
    "01000100", --  338 - 0x152  :   68 - 0x44
    "01000100", --  339 - 0x153  :   68 - 0x44
    "01000100", --  340 - 0x154  :   68 - 0x44
    "01011100", --  341 - 0x155  :   92 - 0x5c
    "01000000", --  342 - 0x156  :   64 - 0x40
    "00000000", --  343 - 0x157  :    0 - 0x0
    "01100110", --  344 - 0x158  :  102 - 0x66 -- plane 1
    "01100110", --  345 - 0x159  :  102 - 0x66
    "01100110", --  346 - 0x15a  :  102 - 0x66
    "01100110", --  347 - 0x15b  :  102 - 0x66
    "01100110", --  348 - 0x15c  :  102 - 0x66
    "01111110", --  349 - 0x15d  :  126 - 0x7e
    "01111110", --  350 - 0x15e  :  126 - 0x7e
    "00000000", --  351 - 0x15f  :    0 - 0x0
    "01000000", --  352 - 0x160  :   64 - 0x40 -- Sprite 0x16
    "01000000", --  353 - 0x161  :   64 - 0x40
    "00000000", --  354 - 0x162  :    0 - 0x0
    "00000000", --  355 - 0x163  :    0 - 0x0
    "00011000", --  356 - 0x164  :   24 - 0x18
    "00111000", --  357 - 0x165  :   56 - 0x38
    "00010000", --  358 - 0x166  :   16 - 0x10
    "00000000", --  359 - 0x167  :    0 - 0x0
    "01111110", --  360 - 0x168  :  126 - 0x7e -- plane 1
    "01100110", --  361 - 0x169  :  102 - 0x66
    "01000010", --  362 - 0x16a  :   66 - 0x42
    "00011000", --  363 - 0x16b  :   24 - 0x18
    "00111100", --  364 - 0x16c  :   60 - 0x3c
    "01111110", --  365 - 0x16d  :  126 - 0x7e
    "11111111", --  366 - 0x16e  :  255 - 0xff
    "11111111", --  367 - 0x16f  :  255 - 0xff
    "01000000", --  368 - 0x170  :   64 - 0x40 -- Sprite 0x17
    "01000000", --  369 - 0x171  :   64 - 0x40
    "01000000", --  370 - 0x172  :   64 - 0x40
    "01000000", --  371 - 0x173  :   64 - 0x40
    "01010000", --  372 - 0x174  :   80 - 0x50
    "01010000", --  373 - 0x175  :   80 - 0x50
    "01001000", --  374 - 0x176  :   72 - 0x48
    "01001000", --  375 - 0x177  :   72 - 0x48
    "01101111", --  376 - 0x178  :  111 - 0x6f -- plane 1
    "01100111", --  377 - 0x179  :  103 - 0x67
    "01110111", --  378 - 0x17a  :  119 - 0x77
    "01110011", --  379 - 0x17b  :  115 - 0x73
    "01111011", --  380 - 0x17c  :  123 - 0x7b
    "01111001", --  381 - 0x17d  :  121 - 0x79
    "01101101", --  382 - 0x17e  :  109 - 0x6d
    "01101100", --  383 - 0x17f  :  108 - 0x6c
    "01000111", --  384 - 0x180  :   71 - 0x47 -- Sprite 0x18
    "01000111", --  385 - 0x181  :   71 - 0x47
    "01000111", --  386 - 0x182  :   71 - 0x47
    "01000111", --  387 - 0x183  :   71 - 0x47
    "01000111", --  388 - 0x184  :   71 - 0x47
    "01011111", --  389 - 0x185  :   95 - 0x5f
    "00000000", --  390 - 0x186  :    0 - 0x0
    "00000000", --  391 - 0x187  :    0 - 0x0
    "01100000", --  392 - 0x188  :   96 - 0x60 -- plane 1
    "01100000", --  393 - 0x189  :   96 - 0x60
    "01100000", --  394 - 0x18a  :   96 - 0x60
    "01100000", --  395 - 0x18b  :   96 - 0x60
    "01100000", --  396 - 0x18c  :   96 - 0x60
    "01111111", --  397 - 0x18d  :  127 - 0x7f
    "01111111", --  398 - 0x18e  :  127 - 0x7f
    "00000000", --  399 - 0x18f  :    0 - 0x0
    "11111100", --  400 - 0x190  :  252 - 0xfc -- Sprite 0x19
    "11111100", --  401 - 0x191  :  252 - 0xfc
    "11111100", --  402 - 0x192  :  252 - 0xfc
    "11111100", --  403 - 0x193  :  252 - 0xfc
    "11111100", --  404 - 0x194  :  252 - 0xfc
    "11011100", --  405 - 0x195  :  220 - 0xdc
    "00011100", --  406 - 0x196  :   28 - 0x1c
    "01000100", --  407 - 0x197  :   68 - 0x44
    "00000110", --  408 - 0x198  :    6 - 0x6 -- plane 1
    "00000110", --  409 - 0x199  :    6 - 0x6
    "00000110", --  410 - 0x19a  :    6 - 0x6
    "00000110", --  411 - 0x19b  :    6 - 0x6
    "00000110", --  412 - 0x19c  :    6 - 0x6
    "11100110", --  413 - 0x19d  :  230 - 0xe6
    "11100110", --  414 - 0x19e  :  230 - 0xe6
    "01100110", --  415 - 0x19f  :  102 - 0x66
    "00010000", --  416 - 0x1a0  :   16 - 0x10 -- Sprite 0x1a
    "00111000", --  417 - 0x1a1  :   56 - 0x38
    "01111100", --  418 - 0x1a2  :  124 - 0x7c
    "11100000", --  419 - 0x1a3  :  224 - 0xe0
    "01000000", --  420 - 0x1a4  :   64 - 0x40
    "00000000", --  421 - 0x1a5  :    0 - 0x0
    "00010000", --  422 - 0x1a6  :   16 - 0x10
    "00100000", --  423 - 0x1a7  :   32 - 0x20
    "11111111", --  424 - 0x1a8  :  255 - 0xff -- plane 1
    "11111111", --  425 - 0x1a9  :  255 - 0xff
    "11111111", --  426 - 0x1aa  :  255 - 0xff
    "11111111", --  427 - 0x1ab  :  255 - 0xff
    "11100111", --  428 - 0x1ac  :  231 - 0xe7
    "11000011", --  429 - 0x1ad  :  195 - 0xc3
    "10011001", --  430 - 0x1ae  :  153 - 0x99
    "00111100", --  431 - 0x1af  :   60 - 0x3c
    "00000000", --  432 - 0x1b0  :    0 - 0x0 -- Sprite 0x1b
    "01111100", --  433 - 0x1b1  :  124 - 0x7c
    "01000000", --  434 - 0x1b2  :   64 - 0x40
    "01000100", --  435 - 0x1b3  :   68 - 0x44
    "01000100", --  436 - 0x1b4  :   68 - 0x44
    "01000100", --  437 - 0x1b5  :   68 - 0x44
    "01000100", --  438 - 0x1b6  :   68 - 0x44
    "01000100", --  439 - 0x1b7  :   68 - 0x44
    "00000000", --  440 - 0x1b8  :    0 - 0x0 -- plane 1
    "01111110", --  441 - 0x1b9  :  126 - 0x7e
    "01111110", --  442 - 0x1ba  :  126 - 0x7e
    "01100110", --  443 - 0x1bb  :  102 - 0x66
    "01100110", --  444 - 0x1bc  :  102 - 0x66
    "01100110", --  445 - 0x1bd  :  102 - 0x66
    "01100110", --  446 - 0x1be  :  102 - 0x66
    "01100110", --  447 - 0x1bf  :  102 - 0x66
    "00010000", --  448 - 0x1c0  :   16 - 0x10 -- Sprite 0x1c
    "00111000", --  449 - 0x1c1  :   56 - 0x38
    "01110001", --  450 - 0x1c2  :  113 - 0x71
    "11100010", --  451 - 0x1c3  :  226 - 0xe2
    "01000100", --  452 - 0x1c4  :   68 - 0x44
    "00001000", --  453 - 0x1c5  :    8 - 0x8
    "00010000", --  454 - 0x1c6  :   16 - 0x10
    "00100000", --  455 - 0x1c7  :   32 - 0x20
    "11111110", --  456 - 0x1c8  :  254 - 0xfe -- plane 1
    "11111100", --  457 - 0x1c9  :  252 - 0xfc
    "11111001", --  458 - 0x1ca  :  249 - 0xf9
    "11110011", --  459 - 0x1cb  :  243 - 0xf3
    "11100111", --  460 - 0x1cc  :  231 - 0xe7
    "11001110", --  461 - 0x1cd  :  206 - 0xce
    "10011100", --  462 - 0x1ce  :  156 - 0x9c
    "00111000", --  463 - 0x1cf  :   56 - 0x38
    "01000000", --  464 - 0x1d0  :   64 - 0x40 -- Sprite 0x1d
    "10000100", --  465 - 0x1d1  :  132 - 0x84
    "00000010", --  466 - 0x1d2  :    2 - 0x2
    "00000111", --  467 - 0x1d3  :    7 - 0x7
    "00001111", --  468 - 0x1d4  :   15 - 0xf
    "00011111", --  469 - 0x1d5  :   31 - 0x1f
    "00111111", --  470 - 0x1d6  :   63 - 0x3f
    "01111111", --  471 - 0x1d7  :  127 - 0x7f
    "01111110", --  472 - 0x1d8  :  126 - 0x7e -- plane 1
    "11100111", --  473 - 0x1d9  :  231 - 0xe7
    "11000011", --  474 - 0x1da  :  195 - 0xc3
    "10000001", --  475 - 0x1db  :  129 - 0x81
    "00000000", --  476 - 0x1dc  :    0 - 0x0
    "00000000", --  477 - 0x1dd  :    0 - 0x0
    "00000000", --  478 - 0x1de  :    0 - 0x0
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "00010000", --  480 - 0x1e0  :   16 - 0x10 -- Sprite 0x1e
    "00011000", --  481 - 0x1e1  :   24 - 0x18
    "00001100", --  482 - 0x1e2  :   12 - 0xc
    "00000110", --  483 - 0x1e3  :    6 - 0x6
    "10000000", --  484 - 0x1e4  :  128 - 0x80
    "11000000", --  485 - 0x1e5  :  192 - 0xc0
    "11100000", --  486 - 0x1e6  :  224 - 0xe0
    "11110000", --  487 - 0x1e7  :  240 - 0xf0
    "01111111", --  488 - 0x1e8  :  127 - 0x7f -- plane 1
    "00111111", --  489 - 0x1e9  :   63 - 0x3f
    "10011111", --  490 - 0x1ea  :  159 - 0x9f
    "11001111", --  491 - 0x1eb  :  207 - 0xcf
    "11100111", --  492 - 0x1ec  :  231 - 0xe7
    "01110011", --  493 - 0x1ed  :  115 - 0x73
    "00111001", --  494 - 0x1ee  :   57 - 0x39
    "00011100", --  495 - 0x1ef  :   28 - 0x1c
    "11111100", --  496 - 0x1f0  :  252 - 0xfc -- Sprite 0x1f
    "11111101", --  497 - 0x1f1  :  253 - 0xfd
    "11111100", --  498 - 0x1f2  :  252 - 0xfc
    "11111110", --  499 - 0x1f3  :  254 - 0xfe
    "11111110", --  500 - 0x1f4  :  254 - 0xfe
    "11111111", --  501 - 0x1f5  :  255 - 0xff
    "11111111", --  502 - 0x1f6  :  255 - 0xff
    "11111111", --  503 - 0x1f7  :  255 - 0xff
    "00000110", --  504 - 0x1f8  :    6 - 0x6 -- plane 1
    "00000111", --  505 - 0x1f9  :    7 - 0x7
    "00000111", --  506 - 0x1fa  :    7 - 0x7
    "00000000", --  507 - 0x1fb  :    0 - 0x0
    "00000000", --  508 - 0x1fc  :    0 - 0x0
    "00000000", --  509 - 0x1fd  :    0 - 0x0
    "00000000", --  510 - 0x1fe  :    0 - 0x0
    "00000000", --  511 - 0x1ff  :    0 - 0x0
    "00000000", --  512 - 0x200  :    0 - 0x0 -- Sprite 0x20
    "11111111", --  513 - 0x201  :  255 - 0xff
    "00000000", --  514 - 0x202  :    0 - 0x0
    "00000000", --  515 - 0x203  :    0 - 0x0
    "00000000", --  516 - 0x204  :    0 - 0x0
    "11111111", --  517 - 0x205  :  255 - 0xff
    "11111111", --  518 - 0x206  :  255 - 0xff
    "11111111", --  519 - 0x207  :  255 - 0xff
    "00000000", --  520 - 0x208  :    0 - 0x0 -- plane 1
    "11111111", --  521 - 0x209  :  255 - 0xff
    "11111111", --  522 - 0x20a  :  255 - 0xff
    "00000000", --  523 - 0x20b  :    0 - 0x0
    "00000000", --  524 - 0x20c  :    0 - 0x0
    "00000000", --  525 - 0x20d  :    0 - 0x0
    "00000000", --  526 - 0x20e  :    0 - 0x0
    "00000000", --  527 - 0x20f  :    0 - 0x0
    "01000100", --  528 - 0x210  :   68 - 0x44 -- Sprite 0x21
    "11000101", --  529 - 0x211  :  197 - 0xc5
    "00000000", --  530 - 0x212  :    0 - 0x0
    "00000110", --  531 - 0x213  :    6 - 0x6
    "00000110", --  532 - 0x214  :    6 - 0x6
    "11111111", --  533 - 0x215  :  255 - 0xff
    "11111111", --  534 - 0x216  :  255 - 0xff
    "11111111", --  535 - 0x217  :  255 - 0xff
    "01100110", --  536 - 0x218  :  102 - 0x66 -- plane 1
    "11100111", --  537 - 0x219  :  231 - 0xe7
    "11100111", --  538 - 0x21a  :  231 - 0xe7
    "00000000", --  539 - 0x21b  :    0 - 0x0
    "00000000", --  540 - 0x21c  :    0 - 0x0
    "00000000", --  541 - 0x21d  :    0 - 0x0
    "00000000", --  542 - 0x21e  :    0 - 0x0
    "00000000", --  543 - 0x21f  :    0 - 0x0
    "01000000", --  544 - 0x220  :   64 - 0x40 -- Sprite 0x22
    "10000001", --  545 - 0x221  :  129 - 0x81
    "00000011", --  546 - 0x222  :    3 - 0x3
    "00000111", --  547 - 0x223  :    7 - 0x7
    "00001111", --  548 - 0x224  :   15 - 0xf
    "11111111", --  549 - 0x225  :  255 - 0xff
    "11111111", --  550 - 0x226  :  255 - 0xff
    "11111111", --  551 - 0x227  :  255 - 0xff
    "01110000", --  552 - 0x228  :  112 - 0x70 -- plane 1
    "11100000", --  553 - 0x229  :  224 - 0xe0
    "11000000", --  554 - 0x22a  :  192 - 0xc0
    "00000000", --  555 - 0x22b  :    0 - 0x0
    "00000000", --  556 - 0x22c  :    0 - 0x0
    "00000000", --  557 - 0x22d  :    0 - 0x0
    "00000000", --  558 - 0x22e  :    0 - 0x0
    "00000000", --  559 - 0x22f  :    0 - 0x0
    "11111000", --  560 - 0x230  :  248 - 0xf8 -- Sprite 0x23
    "11111100", --  561 - 0x231  :  252 - 0xfc
    "11111110", --  562 - 0x232  :  254 - 0xfe
    "11111110", --  563 - 0x233  :  254 - 0xfe
    "11111111", --  564 - 0x234  :  255 - 0xff
    "11111111", --  565 - 0x235  :  255 - 0xff
    "11111111", --  566 - 0x236  :  255 - 0xff
    "11111111", --  567 - 0x237  :  255 - 0xff
    "00001110", --  568 - 0x238  :   14 - 0xe -- plane 1
    "00000111", --  569 - 0x239  :    7 - 0x7
    "00000011", --  570 - 0x23a  :    3 - 0x3
    "00000000", --  571 - 0x23b  :    0 - 0x0
    "00000000", --  572 - 0x23c  :    0 - 0x0
    "00000000", --  573 - 0x23d  :    0 - 0x0
    "00000000", --  574 - 0x23e  :    0 - 0x0
    "00000000", --  575 - 0x23f  :    0 - 0x0
    "01000111", --  576 - 0x240  :   71 - 0x47 -- Sprite 0x24
    "11000111", --  577 - 0x241  :  199 - 0xc7
    "00000111", --  578 - 0x242  :    7 - 0x7
    "00000111", --  579 - 0x243  :    7 - 0x7
    "00000111", --  580 - 0x244  :    7 - 0x7
    "11111111", --  581 - 0x245  :  255 - 0xff
    "11111111", --  582 - 0x246  :  255 - 0xff
    "11111111", --  583 - 0x247  :  255 - 0xff
    "01100000", --  584 - 0x248  :   96 - 0x60 -- plane 1
    "11100000", --  585 - 0x249  :  224 - 0xe0
    "11100000", --  586 - 0x24a  :  224 - 0xe0
    "00000000", --  587 - 0x24b  :    0 - 0x0
    "00000000", --  588 - 0x24c  :    0 - 0x0
    "00000000", --  589 - 0x24d  :    0 - 0x0
    "00000000", --  590 - 0x24e  :    0 - 0x0
    "00000000", --  591 - 0x24f  :    0 - 0x0
    "11111111", --  592 - 0x250  :  255 - 0xff -- Sprite 0x25
    "11111111", --  593 - 0x251  :  255 - 0xff
    "11111111", --  594 - 0x252  :  255 - 0xff
    "11111111", --  595 - 0x253  :  255 - 0xff
    "11111111", --  596 - 0x254  :  255 - 0xff
    "11111111", --  597 - 0x255  :  255 - 0xff
    "00011111", --  598 - 0x256  :   31 - 0x1f
    "00001111", --  599 - 0x257  :   15 - 0xf
    "00000000", --  600 - 0x258  :    0 - 0x0 -- plane 1
    "00000000", --  601 - 0x259  :    0 - 0x0
    "00000000", --  602 - 0x25a  :    0 - 0x0
    "00000000", --  603 - 0x25b  :    0 - 0x0
    "00000000", --  604 - 0x25c  :    0 - 0x0
    "11000000", --  605 - 0x25d  :  192 - 0xc0
    "11100000", --  606 - 0x25e  :  224 - 0xe0
    "01110000", --  607 - 0x25f  :  112 - 0x70
    "11111111", --  608 - 0x260  :  255 - 0xff -- Sprite 0x26
    "11111111", --  609 - 0x261  :  255 - 0xff
    "11111111", --  610 - 0x262  :  255 - 0xff
    "11111111", --  611 - 0x263  :  255 - 0xff
    "11111111", --  612 - 0x264  :  255 - 0xff
    "11111111", --  613 - 0x265  :  255 - 0xff
    "11111100", --  614 - 0x266  :  252 - 0xfc
    "11111000", --  615 - 0x267  :  248 - 0xf8
    "00000000", --  616 - 0x268  :    0 - 0x0 -- plane 1
    "00000000", --  617 - 0x269  :    0 - 0x0
    "00000000", --  618 - 0x26a  :    0 - 0x0
    "00000000", --  619 - 0x26b  :    0 - 0x0
    "00000000", --  620 - 0x26c  :    0 - 0x0
    "00000011", --  621 - 0x26d  :    3 - 0x3
    "00000111", --  622 - 0x26e  :    7 - 0x7
    "00001110", --  623 - 0x26f  :   14 - 0xe
    "00100111", --  624 - 0x270  :   39 - 0x27 -- Sprite 0x27
    "00010011", --  625 - 0x271  :   19 - 0x13
    "00001001", --  626 - 0x272  :    9 - 0x9
    "11000100", --  627 - 0x273  :  196 - 0xc4
    "01100010", --  628 - 0x274  :   98 - 0x62
    "00100001", --  629 - 0x275  :   33 - 0x21
    "00000000", --  630 - 0x276  :    0 - 0x0
    "00000000", --  631 - 0x277  :    0 - 0x0
    "00111000", --  632 - 0x278  :   56 - 0x38 -- plane 1
    "10011100", --  633 - 0x279  :  156 - 0x9c
    "11001110", --  634 - 0x27a  :  206 - 0xce
    "11100111", --  635 - 0x27b  :  231 - 0xe7
    "11110011", --  636 - 0x27c  :  243 - 0xf3
    "11111001", --  637 - 0x27d  :  249 - 0xf9
    "11111100", --  638 - 0x27e  :  252 - 0xfc
    "11111110", --  639 - 0x27f  :  254 - 0xfe
    "11111111", --  640 - 0x280  :  255 - 0xff -- Sprite 0x28
    "11111111", --  641 - 0x281  :  255 - 0xff
    "11111111", --  642 - 0x282  :  255 - 0xff
    "11111111", --  643 - 0x283  :  255 - 0xff
    "01111111", --  644 - 0x284  :  127 - 0x7f
    "00111110", --  645 - 0x285  :   62 - 0x3e
    "10011100", --  646 - 0x286  :  156 - 0x9c
    "01001000", --  647 - 0x287  :   72 - 0x48
    "00000000", --  648 - 0x288  :    0 - 0x0 -- plane 1
    "00000000", --  649 - 0x289  :    0 - 0x0
    "00000000", --  650 - 0x28a  :    0 - 0x0
    "00000000", --  651 - 0x28b  :    0 - 0x0
    "10000001", --  652 - 0x28c  :  129 - 0x81
    "11000011", --  653 - 0x28d  :  195 - 0xc3
    "11100111", --  654 - 0x28e  :  231 - 0xe7
    "01111110", --  655 - 0x28f  :  126 - 0x7e
    "11110000", --  656 - 0x290  :  240 - 0xf0 -- Sprite 0x29
    "11100000", --  657 - 0x291  :  224 - 0xe0
    "11000000", --  658 - 0x292  :  192 - 0xc0
    "10000000", --  659 - 0x293  :  128 - 0x80
    "00000000", --  660 - 0x294  :    0 - 0x0
    "00000010", --  661 - 0x295  :    2 - 0x2
    "00000101", --  662 - 0x296  :    5 - 0x5
    "00000010", --  663 - 0x297  :    2 - 0x2
    "00011100", --  664 - 0x298  :   28 - 0x1c -- plane 1
    "00111001", --  665 - 0x299  :   57 - 0x39
    "01110011", --  666 - 0x29a  :  115 - 0x73
    "11100111", --  667 - 0x29b  :  231 - 0xe7
    "11001111", --  668 - 0x29c  :  207 - 0xcf
    "10011111", --  669 - 0x29d  :  159 - 0x9f
    "00111111", --  670 - 0x29e  :   63 - 0x3f
    "01111111", --  671 - 0x29f  :  127 - 0x7f
    "01000111", --  672 - 0x2a0  :   71 - 0x47 -- Sprite 0x2a
    "01000110", --  673 - 0x2a1  :   70 - 0x46
    "01000110", --  674 - 0x2a2  :   70 - 0x46
    "01000100", --  675 - 0x2a3  :   68 - 0x44
    "01000100", --  676 - 0x2a4  :   68 - 0x44
    "01000100", --  677 - 0x2a5  :   68 - 0x44
    "01000100", --  678 - 0x2a6  :   68 - 0x44
    "01000100", --  679 - 0x2a7  :   68 - 0x44
    "01100001", --  680 - 0x2a8  :   97 - 0x61 -- plane 1
    "01100011", --  681 - 0x2a9  :   99 - 0x63
    "01100011", --  682 - 0x2aa  :   99 - 0x63
    "01100111", --  683 - 0x2ab  :  103 - 0x67
    "01100110", --  684 - 0x2ac  :  102 - 0x66
    "01100110", --  685 - 0x2ad  :  102 - 0x66
    "01100110", --  686 - 0x2ae  :  102 - 0x66
    "01100110", --  687 - 0x2af  :  102 - 0x66
    "01111111", --  688 - 0x2b0  :  127 - 0x7f -- Sprite 0x2b
    "00111111", --  689 - 0x2b1  :   63 - 0x3f
    "10011111", --  690 - 0x2b2  :  159 - 0x9f
    "10001111", --  691 - 0x2b3  :  143 - 0x8f
    "01001111", --  692 - 0x2b4  :   79 - 0x4f
    "01000111", --  693 - 0x2b5  :   71 - 0x47
    "01000111", --  694 - 0x2b6  :   71 - 0x47
    "01000111", --  695 - 0x2b7  :   71 - 0x47
    "10000000", --  696 - 0x2b8  :  128 - 0x80 -- plane 1
    "11000000", --  697 - 0x2b9  :  192 - 0xc0
    "11000000", --  698 - 0x2ba  :  192 - 0xc0
    "11100000", --  699 - 0x2bb  :  224 - 0xe0
    "01100000", --  700 - 0x2bc  :   96 - 0x60
    "01100000", --  701 - 0x2bd  :   96 - 0x60
    "01100000", --  702 - 0x2be  :   96 - 0x60
    "01100000", --  703 - 0x2bf  :   96 - 0x60
    "00100000", --  704 - 0x2c0  :   32 - 0x20 -- Sprite 0x2c
    "00010000", --  705 - 0x2c1  :   16 - 0x10
    "00000000", --  706 - 0x2c2  :    0 - 0x0
    "11000000", --  707 - 0x2c3  :  192 - 0xc0
    "01100000", --  708 - 0x2c4  :   96 - 0x60
    "00100010", --  709 - 0x2c5  :   34 - 0x22
    "00000101", --  710 - 0x2c6  :    5 - 0x5
    "00000010", --  711 - 0x2c7  :    2 - 0x2
    "00111100", --  712 - 0x2c8  :   60 - 0x3c -- plane 1
    "10011001", --  713 - 0x2c9  :  153 - 0x99
    "11000011", --  714 - 0x2ca  :  195 - 0xc3
    "11100111", --  715 - 0x2cb  :  231 - 0xe7
    "11111111", --  716 - 0x2cc  :  255 - 0xff
    "11111111", --  717 - 0x2cd  :  255 - 0xff
    "11111111", --  718 - 0x2ce  :  255 - 0xff
    "11111111", --  719 - 0x2cf  :  255 - 0xff
    "00000000", --  720 - 0x2d0  :    0 - 0x0 -- Sprite 0x2d
    "01111111", --  721 - 0x2d1  :  127 - 0x7f
    "01000000", --  722 - 0x2d2  :   64 - 0x40
    "01000000", --  723 - 0x2d3  :   64 - 0x40
    "01000000", --  724 - 0x2d4  :   64 - 0x40
    "01000111", --  725 - 0x2d5  :   71 - 0x47
    "01000111", --  726 - 0x2d6  :   71 - 0x47
    "01000111", --  727 - 0x2d7  :   71 - 0x47
    "00000000", --  728 - 0x2d8  :    0 - 0x0 -- plane 1
    "01111111", --  729 - 0x2d9  :  127 - 0x7f
    "01111111", --  730 - 0x2da  :  127 - 0x7f
    "01100000", --  731 - 0x2db  :   96 - 0x60
    "01100000", --  732 - 0x2dc  :   96 - 0x60
    "01100000", --  733 - 0x2dd  :   96 - 0x60
    "01100000", --  734 - 0x2de  :   96 - 0x60
    "01100000", --  735 - 0x2df  :   96 - 0x60
    "01000100", --  736 - 0x2e0  :   68 - 0x44 -- Sprite 0x2e
    "11000100", --  737 - 0x2e1  :  196 - 0xc4
    "00000100", --  738 - 0x2e2  :    4 - 0x4
    "00000100", --  739 - 0x2e3  :    4 - 0x4
    "00000100", --  740 - 0x2e4  :    4 - 0x4
    "11111100", --  741 - 0x2e5  :  252 - 0xfc
    "11111100", --  742 - 0x2e6  :  252 - 0xfc
    "11111100", --  743 - 0x2e7  :  252 - 0xfc
    "01100110", --  744 - 0x2e8  :  102 - 0x66 -- plane 1
    "11100110", --  745 - 0x2e9  :  230 - 0xe6
    "11100110", --  746 - 0x2ea  :  230 - 0xe6
    "00000110", --  747 - 0x2eb  :    6 - 0x6
    "00000110", --  748 - 0x2ec  :    6 - 0x6
    "00000110", --  749 - 0x2ed  :    6 - 0x6
    "00000110", --  750 - 0x2ee  :    6 - 0x6
    "00000110", --  751 - 0x2ef  :    6 - 0x6
    "00000001", --  752 - 0x2f0  :    1 - 0x1 -- Sprite 0x2f
    "01111100", --  753 - 0x2f1  :  124 - 0x7c
    "01000000", --  754 - 0x2f2  :   64 - 0x40
    "01000100", --  755 - 0x2f3  :   68 - 0x44
    "01000100", --  756 - 0x2f4  :   68 - 0x44
    "01000100", --  757 - 0x2f5  :   68 - 0x44
    "01000100", --  758 - 0x2f6  :   68 - 0x44
    "01000100", --  759 - 0x2f7  :   68 - 0x44
    "00000001", --  760 - 0x2f8  :    1 - 0x1 -- plane 1
    "01111100", --  761 - 0x2f9  :  124 - 0x7c
    "01111110", --  762 - 0x2fa  :  126 - 0x7e
    "01100110", --  763 - 0x2fb  :  102 - 0x66
    "01100110", --  764 - 0x2fc  :  102 - 0x66
    "01100110", --  765 - 0x2fd  :  102 - 0x66
    "01100110", --  766 - 0x2fe  :  102 - 0x66
    "01100110", --  767 - 0x2ff  :  102 - 0x66
    "00010000", --  768 - 0x300  :   16 - 0x10 -- Sprite 0x30
    "00111000", --  769 - 0x301  :   56 - 0x38
    "00111100", --  770 - 0x302  :   60 - 0x3c
    "00011000", --  771 - 0x303  :   24 - 0x18
    "00000000", --  772 - 0x304  :    0 - 0x0
    "01000010", --  773 - 0x305  :   66 - 0x42
    "01000100", --  774 - 0x306  :   68 - 0x44
    "01001000", --  775 - 0x307  :   72 - 0x48
    "11111111", --  776 - 0x308  :  255 - 0xff -- plane 1
    "11111111", --  777 - 0x309  :  255 - 0xff
    "01111110", --  778 - 0x30a  :  126 - 0x7e
    "00111100", --  779 - 0x30b  :   60 - 0x3c
    "00011000", --  780 - 0x30c  :   24 - 0x18
    "01000010", --  781 - 0x30d  :   66 - 0x42
    "01100110", --  782 - 0x30e  :  102 - 0x66
    "01111110", --  783 - 0x30f  :  126 - 0x7e
    "01000111", --  784 - 0x310  :   71 - 0x47 -- Sprite 0x31
    "01011111", --  785 - 0x311  :   95 - 0x5f
    "00000000", --  786 - 0x312  :    0 - 0x0
    "00000000", --  787 - 0x313  :    0 - 0x0
    "01110000", --  788 - 0x314  :  112 - 0x70
    "00100010", --  789 - 0x315  :   34 - 0x22
    "00000101", --  790 - 0x316  :    5 - 0x5
    "00000010", --  791 - 0x317  :    2 - 0x2
    "01100000", --  792 - 0x318  :   96 - 0x60 -- plane 1
    "01111111", --  793 - 0x319  :  127 - 0x7f
    "01111111", --  794 - 0x31a  :  127 - 0x7f
    "00000000", --  795 - 0x31b  :    0 - 0x0
    "11111111", --  796 - 0x31c  :  255 - 0xff
    "11111111", --  797 - 0x31d  :  255 - 0xff
    "11111111", --  798 - 0x31e  :  255 - 0xff
    "11111111", --  799 - 0x31f  :  255 - 0xff
    "11111111", --  800 - 0x320  :  255 - 0xff -- Sprite 0x32
    "11111111", --  801 - 0x321  :  255 - 0xff
    "00000000", --  802 - 0x322  :    0 - 0x0
    "00000000", --  803 - 0x323  :    0 - 0x0
    "01110000", --  804 - 0x324  :  112 - 0x70
    "00100010", --  805 - 0x325  :   34 - 0x22
    "00000101", --  806 - 0x326  :    5 - 0x5
    "00000010", --  807 - 0x327  :    2 - 0x2
    "00000000", --  808 - 0x328  :    0 - 0x0 -- plane 1
    "11111111", --  809 - 0x329  :  255 - 0xff
    "11111111", --  810 - 0x32a  :  255 - 0xff
    "00000000", --  811 - 0x32b  :    0 - 0x0
    "11111111", --  812 - 0x32c  :  255 - 0xff
    "11111111", --  813 - 0x32d  :  255 - 0xff
    "11111111", --  814 - 0x32e  :  255 - 0xff
    "11111111", --  815 - 0x32f  :  255 - 0xff
    "11111111", --  816 - 0x330  :  255 - 0xff -- Sprite 0x33
    "11011111", --  817 - 0x331  :  223 - 0xdf
    "00011111", --  818 - 0x332  :   31 - 0x1f
    "01000111", --  819 - 0x333  :   71 - 0x47
    "01000111", --  820 - 0x334  :   71 - 0x47
    "01000111", --  821 - 0x335  :   71 - 0x47
    "01000111", --  822 - 0x336  :   71 - 0x47
    "01000111", --  823 - 0x337  :   71 - 0x47
    "00000000", --  824 - 0x338  :    0 - 0x0 -- plane 1
    "11100000", --  825 - 0x339  :  224 - 0xe0
    "11100000", --  826 - 0x33a  :  224 - 0xe0
    "01100000", --  827 - 0x33b  :   96 - 0x60
    "01100000", --  828 - 0x33c  :   96 - 0x60
    "01100000", --  829 - 0x33d  :   96 - 0x60
    "01100000", --  830 - 0x33e  :   96 - 0x60
    "01100000", --  831 - 0x33f  :   96 - 0x60
    "01000100", --  832 - 0x340  :   68 - 0x44 -- Sprite 0x34
    "01000100", --  833 - 0x341  :   68 - 0x44
    "01000100", --  834 - 0x342  :   68 - 0x44
    "01000100", --  835 - 0x343  :   68 - 0x44
    "01000100", --  836 - 0x344  :   68 - 0x44
    "01000100", --  837 - 0x345  :   68 - 0x44
    "01000100", --  838 - 0x346  :   68 - 0x44
    "01000100", --  839 - 0x347  :   68 - 0x44
    "01111110", --  840 - 0x348  :  126 - 0x7e -- plane 1
    "01100110", --  841 - 0x349  :  102 - 0x66
    "01100110", --  842 - 0x34a  :  102 - 0x66
    "01100110", --  843 - 0x34b  :  102 - 0x66
    "01100110", --  844 - 0x34c  :  102 - 0x66
    "01100110", --  845 - 0x34d  :  102 - 0x66
    "01100110", --  846 - 0x34e  :  102 - 0x66
    "01100110", --  847 - 0x34f  :  102 - 0x66
    "00010000", --  848 - 0x350  :   16 - 0x10 -- Sprite 0x35
    "00111000", --  849 - 0x351  :   56 - 0x38
    "01111100", --  850 - 0x352  :  124 - 0x7c
    "11111000", --  851 - 0x353  :  248 - 0xf8
    "00000000", --  852 - 0x354  :    0 - 0x0
    "01111111", --  853 - 0x355  :  127 - 0x7f
    "01000000", --  854 - 0x356  :   64 - 0x40
    "01000000", --  855 - 0x357  :   64 - 0x40
    "11111111", --  856 - 0x358  :  255 - 0xff -- plane 1
    "11111111", --  857 - 0x359  :  255 - 0xff
    "11111111", --  858 - 0x35a  :  255 - 0xff
    "11111111", --  859 - 0x35b  :  255 - 0xff
    "00000000", --  860 - 0x35c  :    0 - 0x0
    "01111111", --  861 - 0x35d  :  127 - 0x7f
    "01111111", --  862 - 0x35e  :  127 - 0x7f
    "01100000", --  863 - 0x35f  :   96 - 0x60
    "00010000", --  864 - 0x360  :   16 - 0x10 -- Sprite 0x36
    "00111000", --  865 - 0x361  :   56 - 0x38
    "01111100", --  866 - 0x362  :  124 - 0x7c
    "11111000", --  867 - 0x363  :  248 - 0xf8
    "00000000", --  868 - 0x364  :    0 - 0x0
    "11111111", --  869 - 0x365  :  255 - 0xff
    "00000000", --  870 - 0x366  :    0 - 0x0
    "00000000", --  871 - 0x367  :    0 - 0x0
    "11111111", --  872 - 0x368  :  255 - 0xff -- plane 1
    "11111111", --  873 - 0x369  :  255 - 0xff
    "11111111", --  874 - 0x36a  :  255 - 0xff
    "11111111", --  875 - 0x36b  :  255 - 0xff
    "00000000", --  876 - 0x36c  :    0 - 0x0
    "11111111", --  877 - 0x36d  :  255 - 0xff
    "11111111", --  878 - 0x36e  :  255 - 0xff
    "00000000", --  879 - 0x36f  :    0 - 0x0
    "01000111", --  880 - 0x370  :   71 - 0x47 -- Sprite 0x37
    "01000111", --  881 - 0x371  :   71 - 0x47
    "01000111", --  882 - 0x372  :   71 - 0x47
    "01000111", --  883 - 0x373  :   71 - 0x47
    "01000111", --  884 - 0x374  :   71 - 0x47
    "11000111", --  885 - 0x375  :  199 - 0xc7
    "00000111", --  886 - 0x376  :    7 - 0x7
    "00000111", --  887 - 0x377  :    7 - 0x7
    "01100000", --  888 - 0x378  :   96 - 0x60 -- plane 1
    "01100000", --  889 - 0x379  :   96 - 0x60
    "01100000", --  890 - 0x37a  :   96 - 0x60
    "01100000", --  891 - 0x37b  :   96 - 0x60
    "01100000", --  892 - 0x37c  :   96 - 0x60
    "11100000", --  893 - 0x37d  :  224 - 0xe0
    "11100000", --  894 - 0x37e  :  224 - 0xe0
    "00000000", --  895 - 0x37f  :    0 - 0x0
    "01000100", --  896 - 0x380  :   68 - 0x44 -- Sprite 0x38
    "01000100", --  897 - 0x381  :   68 - 0x44
    "01000100", --  898 - 0x382  :   68 - 0x44
    "01000100", --  899 - 0x383  :   68 - 0x44
    "01000100", --  900 - 0x384  :   68 - 0x44
    "01011000", --  901 - 0x385  :   88 - 0x58
    "00000000", --  902 - 0x386  :    0 - 0x0
    "00000000", --  903 - 0x387  :    0 - 0x0
    "01100110", --  904 - 0x388  :  102 - 0x66 -- plane 1
    "01100110", --  905 - 0x389  :  102 - 0x66
    "01100110", --  906 - 0x38a  :  102 - 0x66
    "01100110", --  907 - 0x38b  :  102 - 0x66
    "01100110", --  908 - 0x38c  :  102 - 0x66
    "01111110", --  909 - 0x38d  :  126 - 0x7e
    "01111100", --  910 - 0x38e  :  124 - 0x7c
    "00000001", --  911 - 0x38f  :    1 - 0x1
    "00010000", --  912 - 0x390  :   16 - 0x10 -- Sprite 0x39
    "00111000", --  913 - 0x391  :   56 - 0x38
    "01111100", --  914 - 0x392  :  124 - 0x7c
    "11111000", --  915 - 0x393  :  248 - 0xf8
    "01110000", --  916 - 0x394  :  112 - 0x70
    "00100010", --  917 - 0x395  :   34 - 0x22
    "00000100", --  918 - 0x396  :    4 - 0x4
    "00000000", --  919 - 0x397  :    0 - 0x0
    "11111111", --  920 - 0x398  :  255 - 0xff -- plane 1
    "11111111", --  921 - 0x399  :  255 - 0xff
    "11111111", --  922 - 0x39a  :  255 - 0xff
    "11111111", --  923 - 0x39b  :  255 - 0xff
    "11111111", --  924 - 0x39c  :  255 - 0xff
    "11111111", --  925 - 0x39d  :  255 - 0xff
    "11111111", --  926 - 0x39e  :  255 - 0xff
    "11111110", --  927 - 0x39f  :  254 - 0xfe
    "01000100", --  928 - 0x3a0  :   68 - 0x44 -- Sprite 0x3a
    "01000100", --  929 - 0x3a1  :   68 - 0x44
    "01000100", --  930 - 0x3a2  :   68 - 0x44
    "01000100", --  931 - 0x3a3  :   68 - 0x44
    "01000100", --  932 - 0x3a4  :   68 - 0x44
    "01011000", --  933 - 0x3a5  :   88 - 0x58
    "00000000", --  934 - 0x3a6  :    0 - 0x0
    "00000000", --  935 - 0x3a7  :    0 - 0x0
    "01100110", --  936 - 0x3a8  :  102 - 0x66 -- plane 1
    "01100110", --  937 - 0x3a9  :  102 - 0x66
    "01100110", --  938 - 0x3aa  :  102 - 0x66
    "01100110", --  939 - 0x3ab  :  102 - 0x66
    "01100110", --  940 - 0x3ac  :  102 - 0x66
    "01111110", --  941 - 0x3ad  :  126 - 0x7e
    "00111100", --  942 - 0x3ae  :   60 - 0x3c
    "10000001", --  943 - 0x3af  :  129 - 0x81
    "01000000", --  944 - 0x3b0  :   64 - 0x40 -- Sprite 0x3b
    "01000111", --  945 - 0x3b1  :   71 - 0x47
    "01000111", --  946 - 0x3b2  :   71 - 0x47
    "01000111", --  947 - 0x3b3  :   71 - 0x47
    "01000111", --  948 - 0x3b4  :   71 - 0x47
    "01011111", --  949 - 0x3b5  :   95 - 0x5f
    "00000000", --  950 - 0x3b6  :    0 - 0x0
    "00000000", --  951 - 0x3b7  :    0 - 0x0
    "01100000", --  952 - 0x3b8  :   96 - 0x60 -- plane 1
    "01100000", --  953 - 0x3b9  :   96 - 0x60
    "01100000", --  954 - 0x3ba  :   96 - 0x60
    "01100000", --  955 - 0x3bb  :   96 - 0x60
    "01100000", --  956 - 0x3bc  :   96 - 0x60
    "01111111", --  957 - 0x3bd  :  127 - 0x7f
    "01111111", --  958 - 0x3be  :  127 - 0x7f
    "00000000", --  959 - 0x3bf  :    0 - 0x0
    "00000000", --  960 - 0x3c0  :    0 - 0x0 -- Sprite 0x3c
    "11111111", --  961 - 0x3c1  :  255 - 0xff
    "11111111", --  962 - 0x3c2  :  255 - 0xff
    "11111111", --  963 - 0x3c3  :  255 - 0xff
    "11111111", --  964 - 0x3c4  :  255 - 0xff
    "11111111", --  965 - 0x3c5  :  255 - 0xff
    "00000000", --  966 - 0x3c6  :    0 - 0x0
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "00000000", --  968 - 0x3c8  :    0 - 0x0 -- plane 1
    "00000000", --  969 - 0x3c9  :    0 - 0x0
    "00000000", --  970 - 0x3ca  :    0 - 0x0
    "00000000", --  971 - 0x3cb  :    0 - 0x0
    "00000000", --  972 - 0x3cc  :    0 - 0x0
    "11111111", --  973 - 0x3cd  :  255 - 0xff
    "11111111", --  974 - 0x3ce  :  255 - 0xff
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "00000111", --  976 - 0x3d0  :    7 - 0x7 -- Sprite 0x3d
    "11111111", --  977 - 0x3d1  :  255 - 0xff
    "11111111", --  978 - 0x3d2  :  255 - 0xff
    "11111111", --  979 - 0x3d3  :  255 - 0xff
    "11111111", --  980 - 0x3d4  :  255 - 0xff
    "11111111", --  981 - 0x3d5  :  255 - 0xff
    "00000000", --  982 - 0x3d6  :    0 - 0x0
    "00000000", --  983 - 0x3d7  :    0 - 0x0
    "00000000", --  984 - 0x3d8  :    0 - 0x0 -- plane 1
    "00000000", --  985 - 0x3d9  :    0 - 0x0
    "00000000", --  986 - 0x3da  :    0 - 0x0
    "00000000", --  987 - 0x3db  :    0 - 0x0
    "00000000", --  988 - 0x3dc  :    0 - 0x0
    "11111111", --  989 - 0x3dd  :  255 - 0xff
    "11111111", --  990 - 0x3de  :  255 - 0xff
    "00000000", --  991 - 0x3df  :    0 - 0x0
    "00010000", --  992 - 0x3e0  :   16 - 0x10 -- Sprite 0x3e
    "00111000", --  993 - 0x3e1  :   56 - 0x38
    "01110001", --  994 - 0x3e2  :  113 - 0x71
    "11100010", --  995 - 0x3e3  :  226 - 0xe2
    "01100010", --  996 - 0x3e4  :   98 - 0x62
    "00100001", --  997 - 0x3e5  :   33 - 0x21
    "00000000", --  998 - 0x3e6  :    0 - 0x0
    "00000000", --  999 - 0x3e7  :    0 - 0x0
    "11111110", -- 1000 - 0x3e8  :  254 - 0xfe -- plane 1
    "11111100", -- 1001 - 0x3e9  :  252 - 0xfc
    "11111001", -- 1002 - 0x3ea  :  249 - 0xf9
    "11110011", -- 1003 - 0x3eb  :  243 - 0xf3
    "11110011", -- 1004 - 0x3ec  :  243 - 0xf3
    "11111001", -- 1005 - 0x3ed  :  249 - 0xf9
    "11111100", -- 1006 - 0x3ee  :  252 - 0xfc
    "11111110", -- 1007 - 0x3ef  :  254 - 0xfe
    "10000111", -- 1008 - 0x3f0  :  135 - 0x87 -- Sprite 0x3f
    "10000111", -- 1009 - 0x3f1  :  135 - 0x87
    "00000111", -- 1010 - 0x3f2  :    7 - 0x7
    "00001111", -- 1011 - 0x3f3  :   15 - 0xf
    "00001111", -- 1012 - 0x3f4  :   15 - 0xf
    "00011111", -- 1013 - 0x3f5  :   31 - 0x1f
    "10011111", -- 1014 - 0x3f6  :  159 - 0x9f
    "10001111", -- 1015 - 0x3f7  :  143 - 0x8f
    "11100000", -- 1016 - 0x3f8  :  224 - 0xe0 -- plane 1
    "11000000", -- 1017 - 0x3f9  :  192 - 0xc0
    "11000000", -- 1018 - 0x3fa  :  192 - 0xc0
    "10000000", -- 1019 - 0x3fb  :  128 - 0x80
    "10000000", -- 1020 - 0x3fc  :  128 - 0x80
    "11000000", -- 1021 - 0x3fd  :  192 - 0xc0
    "11000000", -- 1022 - 0x3fe  :  192 - 0xc0
    "11100000", -- 1023 - 0x3ff  :  224 - 0xe0
    "01000100", -- 1024 - 0x400  :   68 - 0x44 -- Sprite 0x40
    "01000100", -- 1025 - 0x401  :   68 - 0x44
    "01000100", -- 1026 - 0x402  :   68 - 0x44
    "01000100", -- 1027 - 0x403  :   68 - 0x44
    "01000100", -- 1028 - 0x404  :   68 - 0x44
    "01000110", -- 1029 - 0x405  :   70 - 0x46
    "01000110", -- 1030 - 0x406  :   70 - 0x46
    "01000111", -- 1031 - 0x407  :   71 - 0x47
    "01100110", -- 1032 - 0x408  :  102 - 0x66 -- plane 1
    "01100110", -- 1033 - 0x409  :  102 - 0x66
    "01100110", -- 1034 - 0x40a  :  102 - 0x66
    "01100110", -- 1035 - 0x40b  :  102 - 0x66
    "01100111", -- 1036 - 0x40c  :  103 - 0x67
    "01100011", -- 1037 - 0x40d  :   99 - 0x63
    "01100011", -- 1038 - 0x40e  :   99 - 0x63
    "01100001", -- 1039 - 0x40f  :   97 - 0x61
    "00010000", -- 1040 - 0x410  :   16 - 0x10 -- Sprite 0x41
    "00111000", -- 1041 - 0x411  :   56 - 0x38
    "01111100", -- 1042 - 0x412  :  124 - 0x7c
    "01111000", -- 1043 - 0x413  :  120 - 0x78
    "00110000", -- 1044 - 0x414  :   48 - 0x30
    "00000010", -- 1045 - 0x415  :    2 - 0x2
    "00000101", -- 1046 - 0x416  :    5 - 0x5
    "00000010", -- 1047 - 0x417  :    2 - 0x2
    "11111111", -- 1048 - 0x418  :  255 - 0xff -- plane 1
    "11111111", -- 1049 - 0x419  :  255 - 0xff
    "11111111", -- 1050 - 0x41a  :  255 - 0xff
    "01111111", -- 1051 - 0x41b  :  127 - 0x7f
    "01111111", -- 1052 - 0x41c  :  127 - 0x7f
    "00111111", -- 1053 - 0x41d  :   63 - 0x3f
    "10011111", -- 1054 - 0x41e  :  159 - 0x9f
    "11000111", -- 1055 - 0x41f  :  199 - 0xc7
    "00010000", -- 1056 - 0x420  :   16 - 0x10 -- Sprite 0x42
    "00111000", -- 1057 - 0x421  :   56 - 0x38
    "01111100", -- 1058 - 0x422  :  124 - 0x7c
    "11111000", -- 1059 - 0x423  :  248 - 0xf8
    "01110000", -- 1060 - 0x424  :  112 - 0x70
    "00100000", -- 1061 - 0x425  :   32 - 0x20
    "00000001", -- 1062 - 0x426  :    1 - 0x1
    "00000010", -- 1063 - 0x427  :    2 - 0x2
    "11111111", -- 1064 - 0x428  :  255 - 0xff -- plane 1
    "11111111", -- 1065 - 0x429  :  255 - 0xff
    "11111111", -- 1066 - 0x42a  :  255 - 0xff
    "11111110", -- 1067 - 0x42b  :  254 - 0xfe
    "11111110", -- 1068 - 0x42c  :  254 - 0xfe
    "11111100", -- 1069 - 0x42d  :  252 - 0xfc
    "11111001", -- 1070 - 0x42e  :  249 - 0xf9
    "11100011", -- 1071 - 0x42f  :  227 - 0xe3
    "01000100", -- 1072 - 0x430  :   68 - 0x44 -- Sprite 0x43
    "01000100", -- 1073 - 0x431  :   68 - 0x44
    "01000100", -- 1074 - 0x432  :   68 - 0x44
    "01000100", -- 1075 - 0x433  :   68 - 0x44
    "10000100", -- 1076 - 0x434  :  132 - 0x84
    "10000100", -- 1077 - 0x435  :  132 - 0x84
    "00000100", -- 1078 - 0x436  :    4 - 0x4
    "00001100", -- 1079 - 0x437  :   12 - 0xc
    "01100110", -- 1080 - 0x438  :  102 - 0x66 -- plane 1
    "01100110", -- 1081 - 0x439  :  102 - 0x66
    "01100110", -- 1082 - 0x43a  :  102 - 0x66
    "01100110", -- 1083 - 0x43b  :  102 - 0x66
    "11100110", -- 1084 - 0x43c  :  230 - 0xe6
    "11000110", -- 1085 - 0x43d  :  198 - 0xc6
    "11000110", -- 1086 - 0x43e  :  198 - 0xc6
    "10000110", -- 1087 - 0x43f  :  134 - 0x86
    "00010000", -- 1088 - 0x440  :   16 - 0x10 -- Sprite 0x44
    "00111000", -- 1089 - 0x441  :   56 - 0x38
    "01111100", -- 1090 - 0x442  :  124 - 0x7c
    "11111000", -- 1091 - 0x443  :  248 - 0xf8
    "01110000", -- 1092 - 0x444  :  112 - 0x70
    "00100010", -- 1093 - 0x445  :   34 - 0x22
    "00000101", -- 1094 - 0x446  :    5 - 0x5
    "00000010", -- 1095 - 0x447  :    2 - 0x2
    "11111110", -- 1096 - 0x448  :  254 - 0xfe -- plane 1
    "11111111", -- 1097 - 0x449  :  255 - 0xff
    "11111111", -- 1098 - 0x44a  :  255 - 0xff
    "11111111", -- 1099 - 0x44b  :  255 - 0xff
    "11111111", -- 1100 - 0x44c  :  255 - 0xff
    "11111111", -- 1101 - 0x44d  :  255 - 0xff
    "11111111", -- 1102 - 0x44e  :  255 - 0xff
    "11111111", -- 1103 - 0x44f  :  255 - 0xff
    "01001111", -- 1104 - 0x450  :   79 - 0x4f -- Sprite 0x45
    "01000111", -- 1105 - 0x451  :   71 - 0x47
    "01000111", -- 1106 - 0x452  :   71 - 0x47
    "01000111", -- 1107 - 0x453  :   71 - 0x47
    "01000111", -- 1108 - 0x454  :   71 - 0x47
    "01000111", -- 1109 - 0x455  :   71 - 0x47
    "01000111", -- 1110 - 0x456  :   71 - 0x47
    "01000111", -- 1111 - 0x457  :   71 - 0x47
    "01100000", -- 1112 - 0x458  :   96 - 0x60 -- plane 1
    "01100000", -- 1113 - 0x459  :   96 - 0x60
    "01100000", -- 1114 - 0x45a  :   96 - 0x60
    "01100000", -- 1115 - 0x45b  :   96 - 0x60
    "01100000", -- 1116 - 0x45c  :   96 - 0x60
    "01100000", -- 1117 - 0x45d  :   96 - 0x60
    "01100000", -- 1118 - 0x45e  :   96 - 0x60
    "01100000", -- 1119 - 0x45f  :   96 - 0x60
    "10100000", -- 1120 - 0x460  :  160 - 0xa0 -- Sprite 0x46
    "10011111", -- 1121 - 0x461  :  159 - 0x9f
    "11000000", -- 1122 - 0x462  :  192 - 0xc0
    "11100000", -- 1123 - 0x463  :  224 - 0xe0
    "11111000", -- 1124 - 0x464  :  248 - 0xf8
    "11111111", -- 1125 - 0x465  :  255 - 0xff
    "11111111", -- 1126 - 0x466  :  255 - 0xff
    "11111111", -- 1127 - 0x467  :  255 - 0xff
    "11110000", -- 1128 - 0x468  :  240 - 0xf0 -- plane 1
    "01111111", -- 1129 - 0x469  :  127 - 0x7f
    "00011111", -- 1130 - 0x46a  :   31 - 0x1f
    "00000000", -- 1131 - 0x46b  :    0 - 0x0
    "00000000", -- 1132 - 0x46c  :    0 - 0x0
    "00000000", -- 1133 - 0x46d  :    0 - 0x0
    "00000000", -- 1134 - 0x46e  :    0 - 0x0
    "00000000", -- 1135 - 0x46f  :    0 - 0x0
    "00001100", -- 1136 - 0x470  :   12 - 0xc -- Sprite 0x47
    "11110000", -- 1137 - 0x471  :  240 - 0xf0
    "00000000", -- 1138 - 0x472  :    0 - 0x0
    "00000000", -- 1139 - 0x473  :    0 - 0x0
    "00000001", -- 1140 - 0x474  :    1 - 0x1
    "11111111", -- 1141 - 0x475  :  255 - 0xff
    "11111111", -- 1142 - 0x476  :  255 - 0xff
    "11111111", -- 1143 - 0x477  :  255 - 0xff
    "00001111", -- 1144 - 0x478  :   15 - 0xf -- plane 1
    "11111110", -- 1145 - 0x479  :  254 - 0xfe
    "11111000", -- 1146 - 0x47a  :  248 - 0xf8
    "00000000", -- 1147 - 0x47b  :    0 - 0x0
    "00000000", -- 1148 - 0x47c  :    0 - 0x0
    "00000000", -- 1149 - 0x47d  :    0 - 0x0
    "00000000", -- 1150 - 0x47e  :    0 - 0x0
    "00000000", -- 1151 - 0x47f  :    0 - 0x0
    "00001100", -- 1152 - 0x480  :   12 - 0xc -- Sprite 0x48
    "00011101", -- 1153 - 0x481  :   29 - 0x1d
    "00111000", -- 1154 - 0x482  :   56 - 0x38
    "01111110", -- 1155 - 0x483  :  126 - 0x7e
    "11111110", -- 1156 - 0x484  :  254 - 0xfe
    "11111111", -- 1157 - 0x485  :  255 - 0xff
    "11111111", -- 1158 - 0x486  :  255 - 0xff
    "11111111", -- 1159 - 0x487  :  255 - 0xff
    "00000110", -- 1160 - 0x488  :    6 - 0x6 -- plane 1
    "00000111", -- 1161 - 0x489  :    7 - 0x7
    "00000111", -- 1162 - 0x48a  :    7 - 0x7
    "00000000", -- 1163 - 0x48b  :    0 - 0x0
    "00000000", -- 1164 - 0x48c  :    0 - 0x0
    "00000000", -- 1165 - 0x48d  :    0 - 0x0
    "00000000", -- 1166 - 0x48e  :    0 - 0x0
    "00000000", -- 1167 - 0x48f  :    0 - 0x0
    "11111111", -- 1168 - 0x490  :  255 - 0xff -- Sprite 0x49
    "11111111", -- 1169 - 0x491  :  255 - 0xff
    "11111111", -- 1170 - 0x492  :  255 - 0xff
    "11111111", -- 1171 - 0x493  :  255 - 0xff
    "11111111", -- 1172 - 0x494  :  255 - 0xff
    "11111111", -- 1173 - 0x495  :  255 - 0xff
    "11111111", -- 1174 - 0x496  :  255 - 0xff
    "11111111", -- 1175 - 0x497  :  255 - 0xff
    "00000000", -- 1176 - 0x498  :    0 - 0x0 -- plane 1
    "00000000", -- 1177 - 0x499  :    0 - 0x0
    "00000000", -- 1178 - 0x49a  :    0 - 0x0
    "00000000", -- 1179 - 0x49b  :    0 - 0x0
    "00000000", -- 1180 - 0x49c  :    0 - 0x0
    "00000000", -- 1181 - 0x49d  :    0 - 0x0
    "00000000", -- 1182 - 0x49e  :    0 - 0x0
    "00000000", -- 1183 - 0x49f  :    0 - 0x0
    "11111111", -- 1184 - 0x4a0  :  255 - 0xff -- Sprite 0x4a
    "11101111", -- 1185 - 0x4a1  :  239 - 0xef
    "11111101", -- 1186 - 0x4a2  :  253 - 0xfd
    "11111111", -- 1187 - 0x4a3  :  255 - 0xff
    "11111111", -- 1188 - 0x4a4  :  255 - 0xff
    "11101111", -- 1189 - 0x4a5  :  239 - 0xef
    "11111110", -- 1190 - 0x4a6  :  254 - 0xfe
    "11111111", -- 1191 - 0x4a7  :  255 - 0xff
    "00000000", -- 1192 - 0x4a8  :    0 - 0x0 -- plane 1
    "01110110", -- 1193 - 0x4a9  :  118 - 0x76
    "01010111", -- 1194 - 0x4aa  :   87 - 0x57
    "01010101", -- 1195 - 0x4ab  :   85 - 0x55
    "01010101", -- 1196 - 0x4ac  :   85 - 0x55
    "01110101", -- 1197 - 0x4ad  :  117 - 0x75
    "01000111", -- 1198 - 0x4ae  :   71 - 0x47
    "00000000", -- 1199 - 0x4af  :    0 - 0x0
    "11111111", -- 1200 - 0x4b0  :  255 - 0xff -- Sprite 0x4b
    "11101010", -- 1201 - 0x4b1  :  234 - 0xea
    "11111111", -- 1202 - 0x4b2  :  255 - 0xff
    "10101111", -- 1203 - 0x4b3  :  175 - 0xaf
    "11111111", -- 1204 - 0x4b4  :  255 - 0xff
    "11111111", -- 1205 - 0x4b5  :  255 - 0xff
    "11111010", -- 1206 - 0x4b6  :  250 - 0xfa
    "11111111", -- 1207 - 0x4b7  :  255 - 0xff
    "00000000", -- 1208 - 0x4b8  :    0 - 0x0 -- plane 1
    "01110111", -- 1209 - 0x4b9  :  119 - 0x77
    "00010101", -- 1210 - 0x4ba  :   21 - 0x15
    "01110101", -- 1211 - 0x4bb  :  117 - 0x75
    "01000101", -- 1212 - 0x4bc  :   69 - 0x45
    "01000101", -- 1213 - 0x4bd  :   69 - 0x45
    "01110111", -- 1214 - 0x4be  :  119 - 0x77
    "00000000", -- 1215 - 0x4bf  :    0 - 0x0
    "11111111", -- 1216 - 0x4c0  :  255 - 0xff -- Sprite 0x4c
    "11111111", -- 1217 - 0x4c1  :  255 - 0xff
    "11111111", -- 1218 - 0x4c2  :  255 - 0xff
    "11111111", -- 1219 - 0x4c3  :  255 - 0xff
    "11111111", -- 1220 - 0x4c4  :  255 - 0xff
    "11111111", -- 1221 - 0x4c5  :  255 - 0xff
    "11111110", -- 1222 - 0x4c6  :  254 - 0xfe
    "11111111", -- 1223 - 0x4c7  :  255 - 0xff
    "00000000", -- 1224 - 0x4c8  :    0 - 0x0 -- plane 1
    "00100100", -- 1225 - 0x4c9  :   36 - 0x24
    "01101100", -- 1226 - 0x4ca  :  108 - 0x6c
    "00100100", -- 1227 - 0x4cb  :   36 - 0x24
    "00100100", -- 1228 - 0x4cc  :   36 - 0x24
    "00100100", -- 1229 - 0x4cd  :   36 - 0x24
    "00100101", -- 1230 - 0x4ce  :   37 - 0x25
    "00000000", -- 1231 - 0x4cf  :    0 - 0x0
    "11111111", -- 1232 - 0x4d0  :  255 - 0xff -- Sprite 0x4d
    "10111111", -- 1233 - 0x4d1  :  191 - 0xbf
    "11111110", -- 1234 - 0x4d2  :  254 - 0xfe
    "10101111", -- 1235 - 0x4d3  :  175 - 0xaf
    "11111111", -- 1236 - 0x4d4  :  255 - 0xff
    "11111111", -- 1237 - 0x4d5  :  255 - 0xff
    "11101111", -- 1238 - 0x4d6  :  239 - 0xef
    "11111111", -- 1239 - 0x4d7  :  255 - 0xff
    "00000000", -- 1240 - 0x4d8  :    0 - 0x0 -- plane 1
    "01110100", -- 1241 - 0x4d9  :  116 - 0x74
    "01000111", -- 1242 - 0x4da  :   71 - 0x47
    "01110101", -- 1243 - 0x4db  :  117 - 0x75
    "00010101", -- 1244 - 0x4dc  :   21 - 0x15
    "00010101", -- 1245 - 0x4dd  :   21 - 0x15
    "01110101", -- 1246 - 0x4de  :  117 - 0x75
    "00000000", -- 1247 - 0x4df  :    0 - 0x0
    "11111111", -- 1248 - 0x4e0  :  255 - 0xff -- Sprite 0x4e
    "11111111", -- 1249 - 0x4e1  :  255 - 0xff
    "11111011", -- 1250 - 0x4e2  :  251 - 0xfb
    "11111111", -- 1251 - 0x4e3  :  255 - 0xff
    "11111111", -- 1252 - 0x4e4  :  255 - 0xff
    "11111111", -- 1253 - 0x4e5  :  255 - 0xff
    "11111110", -- 1254 - 0x4e6  :  254 - 0xfe
    "11111111", -- 1255 - 0x4e7  :  255 - 0xff
    "00000000", -- 1256 - 0x4e8  :    0 - 0x0 -- plane 1
    "01000000", -- 1257 - 0x4e9  :   64 - 0x40
    "00011101", -- 1258 - 0x4ea  :   29 - 0x1d
    "01010101", -- 1259 - 0x4eb  :   85 - 0x55
    "01010001", -- 1260 - 0x4ec  :   81 - 0x51
    "01010001", -- 1261 - 0x4ed  :   81 - 0x51
    "01010001", -- 1262 - 0x4ee  :   81 - 0x51
    "00000000", -- 1263 - 0x4ef  :    0 - 0x0
    "11111111", -- 1264 - 0x4f0  :  255 - 0xff -- Sprite 0x4f
    "11111111", -- 1265 - 0x4f1  :  255 - 0xff
    "11110111", -- 1266 - 0x4f2  :  247 - 0xf7
    "11111110", -- 1267 - 0x4f3  :  254 - 0xfe
    "11111011", -- 1268 - 0x4f4  :  251 - 0xfb
    "11111111", -- 1269 - 0x4f5  :  255 - 0xff
    "11101111", -- 1270 - 0x4f6  :  239 - 0xef
    "11111101", -- 1271 - 0x4f7  :  253 - 0xfd
    "00000000", -- 1272 - 0x4f8  :    0 - 0x0 -- plane 1
    "00000000", -- 1273 - 0x4f9  :    0 - 0x0
    "01001000", -- 1274 - 0x4fa  :   72 - 0x48
    "01000001", -- 1275 - 0x4fb  :   65 - 0x41
    "01000100", -- 1276 - 0x4fc  :   68 - 0x44
    "01000000", -- 1277 - 0x4fd  :   64 - 0x40
    "11010000", -- 1278 - 0x4fe  :  208 - 0xd0
    "00000010", -- 1279 - 0x4ff  :    2 - 0x2
    "11111111", -- 1280 - 0x500  :  255 - 0xff -- Sprite 0x50
    "11111111", -- 1281 - 0x501  :  255 - 0xff
    "00000011", -- 1282 - 0x502  :    3 - 0x3
    "00000001", -- 1283 - 0x503  :    1 - 0x1
    "11101110", -- 1284 - 0x504  :  238 - 0xee
    "00000000", -- 1285 - 0x505  :    0 - 0x0
    "11101110", -- 1286 - 0x506  :  238 - 0xee
    "11101110", -- 1287 - 0x507  :  238 - 0xee
    "00000000", -- 1288 - 0x508  :    0 - 0x0 -- plane 1
    "00000000", -- 1289 - 0x509  :    0 - 0x0
    "11111100", -- 1290 - 0x50a  :  252 - 0xfc
    "11111110", -- 1291 - 0x50b  :  254 - 0xfe
    "11101110", -- 1292 - 0x50c  :  238 - 0xee
    "11101110", -- 1293 - 0x50d  :  238 - 0xee
    "11101110", -- 1294 - 0x50e  :  238 - 0xee
    "11101110", -- 1295 - 0x50f  :  238 - 0xee
    "11111111", -- 1296 - 0x510  :  255 - 0xff -- Sprite 0x51
    "11111111", -- 1297 - 0x511  :  255 - 0xff
    "00000011", -- 1298 - 0x512  :    3 - 0x3
    "00000001", -- 1299 - 0x513  :    1 - 0x1
    "11101110", -- 1300 - 0x514  :  238 - 0xee
    "00000000", -- 1301 - 0x515  :    0 - 0x0
    "11101110", -- 1302 - 0x516  :  238 - 0xee
    "11101110", -- 1303 - 0x517  :  238 - 0xee
    "00000000", -- 1304 - 0x518  :    0 - 0x0 -- plane 1
    "00000000", -- 1305 - 0x519  :    0 - 0x0
    "11111100", -- 1306 - 0x51a  :  252 - 0xfc
    "11111110", -- 1307 - 0x51b  :  254 - 0xfe
    "11101110", -- 1308 - 0x51c  :  238 - 0xee
    "11101110", -- 1309 - 0x51d  :  238 - 0xee
    "11101110", -- 1310 - 0x51e  :  238 - 0xee
    "11101110", -- 1311 - 0x51f  :  238 - 0xee
    "11111111", -- 1312 - 0x520  :  255 - 0xff -- Sprite 0x52
    "11111111", -- 1313 - 0x521  :  255 - 0xff
    "00000001", -- 1314 - 0x522  :    1 - 0x1
    "00000000", -- 1315 - 0x523  :    0 - 0x0
    "11100000", -- 1316 - 0x524  :  224 - 0xe0
    "00001111", -- 1317 - 0x525  :   15 - 0xf
    "11111111", -- 1318 - 0x526  :  255 - 0xff
    "11111011", -- 1319 - 0x527  :  251 - 0xfb
    "00000000", -- 1320 - 0x528  :    0 - 0x0 -- plane 1
    "00000000", -- 1321 - 0x529  :    0 - 0x0
    "11111110", -- 1322 - 0x52a  :  254 - 0xfe
    "11111110", -- 1323 - 0x52b  :  254 - 0xfe
    "11100000", -- 1324 - 0x52c  :  224 - 0xe0
    "11100000", -- 1325 - 0x52d  :  224 - 0xe0
    "11111000", -- 1326 - 0x52e  :  248 - 0xf8
    "11111000", -- 1327 - 0x52f  :  248 - 0xf8
    "11111111", -- 1328 - 0x530  :  255 - 0xff -- Sprite 0x53
    "11111111", -- 1329 - 0x531  :  255 - 0xff
    "10000011", -- 1330 - 0x532  :  131 - 0x83
    "00000001", -- 1331 - 0x533  :    1 - 0x1
    "11101110", -- 1332 - 0x534  :  238 - 0xee
    "00000000", -- 1333 - 0x535  :    0 - 0x0
    "11111111", -- 1334 - 0x536  :  255 - 0xff
    "11111111", -- 1335 - 0x537  :  255 - 0xff
    "00000000", -- 1336 - 0x538  :    0 - 0x0 -- plane 1
    "00000000", -- 1337 - 0x539  :    0 - 0x0
    "01111100", -- 1338 - 0x53a  :  124 - 0x7c
    "11111110", -- 1339 - 0x53b  :  254 - 0xfe
    "11101110", -- 1340 - 0x53c  :  238 - 0xee
    "11100000", -- 1341 - 0x53d  :  224 - 0xe0
    "11111100", -- 1342 - 0x53e  :  252 - 0xfc
    "01111110", -- 1343 - 0x53f  :  126 - 0x7e
    "11111111", -- 1344 - 0x540  :  255 - 0xff -- Sprite 0x54
    "11111111", -- 1345 - 0x541  :  255 - 0xff
    "00000001", -- 1346 - 0x542  :    1 - 0x1
    "00000000", -- 1347 - 0x543  :    0 - 0x0
    "10111000", -- 1348 - 0x544  :  184 - 0xb8
    "11000011", -- 1349 - 0x545  :  195 - 0xc3
    "11111011", -- 1350 - 0x546  :  251 - 0xfb
    "11111011", -- 1351 - 0x547  :  251 - 0xfb
    "00000000", -- 1352 - 0x548  :    0 - 0x0 -- plane 1
    "00000000", -- 1353 - 0x549  :    0 - 0x0
    "11111110", -- 1354 - 0x54a  :  254 - 0xfe
    "11111110", -- 1355 - 0x54b  :  254 - 0xfe
    "00111000", -- 1356 - 0x54c  :   56 - 0x38
    "00111000", -- 1357 - 0x54d  :   56 - 0x38
    "00111000", -- 1358 - 0x54e  :   56 - 0x38
    "00111000", -- 1359 - 0x54f  :   56 - 0x38
    "11111111", -- 1360 - 0x550  :  255 - 0xff -- Sprite 0x55
    "11111111", -- 1361 - 0x551  :  255 - 0xff
    "10000011", -- 1362 - 0x552  :  131 - 0x83
    "00000001", -- 1363 - 0x553  :    1 - 0x1
    "11101110", -- 1364 - 0x554  :  238 - 0xee
    "00000000", -- 1365 - 0x555  :    0 - 0x0
    "11101110", -- 1366 - 0x556  :  238 - 0xee
    "11101110", -- 1367 - 0x557  :  238 - 0xee
    "00000000", -- 1368 - 0x558  :    0 - 0x0 -- plane 1
    "00000000", -- 1369 - 0x559  :    0 - 0x0
    "01111100", -- 1370 - 0x55a  :  124 - 0x7c
    "11111110", -- 1371 - 0x55b  :  254 - 0xfe
    "11101110", -- 1372 - 0x55c  :  238 - 0xee
    "11101110", -- 1373 - 0x55d  :  238 - 0xee
    "11101110", -- 1374 - 0x55e  :  238 - 0xee
    "11101110", -- 1375 - 0x55f  :  238 - 0xee
    "11111111", -- 1376 - 0x560  :  255 - 0xff -- Sprite 0x56
    "11111111", -- 1377 - 0x561  :  255 - 0xff
    "00011111", -- 1378 - 0x562  :   31 - 0x1f
    "00001111", -- 1379 - 0x563  :   15 - 0xf
    "11101111", -- 1380 - 0x564  :  239 - 0xef
    "00001111", -- 1381 - 0x565  :   15 - 0xf
    "11101111", -- 1382 - 0x566  :  239 - 0xef
    "11101111", -- 1383 - 0x567  :  239 - 0xef
    "00000000", -- 1384 - 0x568  :    0 - 0x0 -- plane 1
    "00000000", -- 1385 - 0x569  :    0 - 0x0
    "11100000", -- 1386 - 0x56a  :  224 - 0xe0
    "11100000", -- 1387 - 0x56b  :  224 - 0xe0
    "11100000", -- 1388 - 0x56c  :  224 - 0xe0
    "11100000", -- 1389 - 0x56d  :  224 - 0xe0
    "11100000", -- 1390 - 0x56e  :  224 - 0xe0
    "11100000", -- 1391 - 0x56f  :  224 - 0xe0
    "11111111", -- 1392 - 0x570  :  255 - 0xff -- Sprite 0x57
    "11111111", -- 1393 - 0x571  :  255 - 0xff
    "00010001", -- 1394 - 0x572  :   17 - 0x11
    "00000000", -- 1395 - 0x573  :    0 - 0x0
    "11101110", -- 1396 - 0x574  :  238 - 0xee
    "00000000", -- 1397 - 0x575  :    0 - 0x0
    "11101110", -- 1398 - 0x576  :  238 - 0xee
    "11101110", -- 1399 - 0x577  :  238 - 0xee
    "00000000", -- 1400 - 0x578  :    0 - 0x0 -- plane 1
    "00000000", -- 1401 - 0x579  :    0 - 0x0
    "11101110", -- 1402 - 0x57a  :  238 - 0xee
    "11101110", -- 1403 - 0x57b  :  238 - 0xee
    "11101110", -- 1404 - 0x57c  :  238 - 0xee
    "11101110", -- 1405 - 0x57d  :  238 - 0xee
    "11101110", -- 1406 - 0x57e  :  238 - 0xee
    "11101110", -- 1407 - 0x57f  :  238 - 0xee
    "11111111", -- 1408 - 0x580  :  255 - 0xff -- Sprite 0x58
    "11111111", -- 1409 - 0x581  :  255 - 0xff
    "01110001", -- 1410 - 0x582  :  113 - 0x71
    "00110000", -- 1411 - 0x583  :   48 - 0x30
    "11111110", -- 1412 - 0x584  :  254 - 0xfe
    "00000000", -- 1413 - 0x585  :    0 - 0x0
    "11111110", -- 1414 - 0x586  :  254 - 0xfe
    "11101110", -- 1415 - 0x587  :  238 - 0xee
    "00000000", -- 1416 - 0x588  :    0 - 0x0 -- plane 1
    "00000000", -- 1417 - 0x589  :    0 - 0x0
    "10001110", -- 1418 - 0x58a  :  142 - 0x8e
    "11001110", -- 1419 - 0x58b  :  206 - 0xce
    "11101110", -- 1420 - 0x58c  :  238 - 0xee
    "11111110", -- 1421 - 0x58d  :  254 - 0xfe
    "11111110", -- 1422 - 0x58e  :  254 - 0xfe
    "11101110", -- 1423 - 0x58f  :  238 - 0xee
    "11111111", -- 1424 - 0x590  :  255 - 0xff -- Sprite 0x59
    "11111111", -- 1425 - 0x591  :  255 - 0xff
    "00000011", -- 1426 - 0x592  :    3 - 0x3
    "00000001", -- 1427 - 0x593  :    1 - 0x1
    "11101110", -- 1428 - 0x594  :  238 - 0xee
    "00000000", -- 1429 - 0x595  :    0 - 0x0
    "11101110", -- 1430 - 0x596  :  238 - 0xee
    "11101110", -- 1431 - 0x597  :  238 - 0xee
    "00000000", -- 1432 - 0x598  :    0 - 0x0 -- plane 1
    "00000000", -- 1433 - 0x599  :    0 - 0x0
    "11111100", -- 1434 - 0x59a  :  252 - 0xfc
    "11111110", -- 1435 - 0x59b  :  254 - 0xfe
    "11101110", -- 1436 - 0x59c  :  238 - 0xee
    "11101110", -- 1437 - 0x59d  :  238 - 0xee
    "11101110", -- 1438 - 0x59e  :  238 - 0xee
    "11101110", -- 1439 - 0x59f  :  238 - 0xee
    "11111111", -- 1440 - 0x5a0  :  255 - 0xff -- Sprite 0x5a
    "11111111", -- 1441 - 0x5a1  :  255 - 0xff
    "10000011", -- 1442 - 0x5a2  :  131 - 0x83
    "00000001", -- 1443 - 0x5a3  :    1 - 0x1
    "11101110", -- 1444 - 0x5a4  :  238 - 0xee
    "00000000", -- 1445 - 0x5a5  :    0 - 0x0
    "11101110", -- 1446 - 0x5a6  :  238 - 0xee
    "11101110", -- 1447 - 0x5a7  :  238 - 0xee
    "00000000", -- 1448 - 0x5a8  :    0 - 0x0 -- plane 1
    "00000000", -- 1449 - 0x5a9  :    0 - 0x0
    "01111100", -- 1450 - 0x5aa  :  124 - 0x7c
    "11111110", -- 1451 - 0x5ab  :  254 - 0xfe
    "11101110", -- 1452 - 0x5ac  :  238 - 0xee
    "11101110", -- 1453 - 0x5ad  :  238 - 0xee
    "11101110", -- 1454 - 0x5ae  :  238 - 0xee
    "11101110", -- 1455 - 0x5af  :  238 - 0xee
    "11111111", -- 1456 - 0x5b0  :  255 - 0xff -- Sprite 0x5b
    "11111111", -- 1457 - 0x5b1  :  255 - 0xff
    "00000001", -- 1458 - 0x5b2  :    1 - 0x1
    "00000000", -- 1459 - 0x5b3  :    0 - 0x0
    "11100000", -- 1460 - 0x5b4  :  224 - 0xe0
    "00001111", -- 1461 - 0x5b5  :   15 - 0xf
    "11111111", -- 1462 - 0x5b6  :  255 - 0xff
    "11111011", -- 1463 - 0x5b7  :  251 - 0xfb
    "00000000", -- 1464 - 0x5b8  :    0 - 0x0 -- plane 1
    "00000000", -- 1465 - 0x5b9  :    0 - 0x0
    "11111110", -- 1466 - 0x5ba  :  254 - 0xfe
    "11111110", -- 1467 - 0x5bb  :  254 - 0xfe
    "11100000", -- 1468 - 0x5bc  :  224 - 0xe0
    "11100000", -- 1469 - 0x5bd  :  224 - 0xe0
    "11111000", -- 1470 - 0x5be  :  248 - 0xf8
    "11111000", -- 1471 - 0x5bf  :  248 - 0xf8
    "11111111", -- 1472 - 0x5c0  :  255 - 0xff -- Sprite 0x5c
    "11111111", -- 1473 - 0x5c1  :  255 - 0xff
    "11111111", -- 1474 - 0x5c2  :  255 - 0xff
    "11111111", -- 1475 - 0x5c3  :  255 - 0xff
    "11111111", -- 1476 - 0x5c4  :  255 - 0xff
    "11111111", -- 1477 - 0x5c5  :  255 - 0xff
    "11111111", -- 1478 - 0x5c6  :  255 - 0xff
    "11011101", -- 1479 - 0x5c7  :  221 - 0xdd
    "00000000", -- 1480 - 0x5c8  :    0 - 0x0 -- plane 1
    "00000000", -- 1481 - 0x5c9  :    0 - 0x0
    "00000000", -- 1482 - 0x5ca  :    0 - 0x0
    "00000000", -- 1483 - 0x5cb  :    0 - 0x0
    "00000000", -- 1484 - 0x5cc  :    0 - 0x0
    "00000000", -- 1485 - 0x5cd  :    0 - 0x0
    "11001100", -- 1486 - 0x5ce  :  204 - 0xcc
    "11001100", -- 1487 - 0x5cf  :  204 - 0xcc
    "11111111", -- 1488 - 0x5d0  :  255 - 0xff -- Sprite 0x5d
    "11111111", -- 1489 - 0x5d1  :  255 - 0xff
    "00000001", -- 1490 - 0x5d2  :    1 - 0x1
    "00000000", -- 1491 - 0x5d3  :    0 - 0x0
    "11100000", -- 1492 - 0x5d4  :  224 - 0xe0
    "00001111", -- 1493 - 0x5d5  :   15 - 0xf
    "11111111", -- 1494 - 0x5d6  :  255 - 0xff
    "11111011", -- 1495 - 0x5d7  :  251 - 0xfb
    "00000000", -- 1496 - 0x5d8  :    0 - 0x0 -- plane 1
    "00000000", -- 1497 - 0x5d9  :    0 - 0x0
    "11111110", -- 1498 - 0x5da  :  254 - 0xfe
    "11111110", -- 1499 - 0x5db  :  254 - 0xfe
    "11100000", -- 1500 - 0x5dc  :  224 - 0xe0
    "11100000", -- 1501 - 0x5dd  :  224 - 0xe0
    "11111000", -- 1502 - 0x5de  :  248 - 0xf8
    "11111000", -- 1503 - 0x5df  :  248 - 0xf8
    "11111111", -- 1504 - 0x5e0  :  255 - 0xff -- Sprite 0x5e
    "11111111", -- 1505 - 0x5e1  :  255 - 0xff
    "00010001", -- 1506 - 0x5e2  :   17 - 0x11
    "00000000", -- 1507 - 0x5e3  :    0 - 0x0
    "11101110", -- 1508 - 0x5e4  :  238 - 0xee
    "00000000", -- 1509 - 0x5e5  :    0 - 0x0
    "11101110", -- 1510 - 0x5e6  :  238 - 0xee
    "11101110", -- 1511 - 0x5e7  :  238 - 0xee
    "00000000", -- 1512 - 0x5e8  :    0 - 0x0 -- plane 1
    "00000000", -- 1513 - 0x5e9  :    0 - 0x0
    "11101110", -- 1514 - 0x5ea  :  238 - 0xee
    "11101110", -- 1515 - 0x5eb  :  238 - 0xee
    "11101110", -- 1516 - 0x5ec  :  238 - 0xee
    "11101110", -- 1517 - 0x5ed  :  238 - 0xee
    "11101110", -- 1518 - 0x5ee  :  238 - 0xee
    "11101110", -- 1519 - 0x5ef  :  238 - 0xee
    "10111101", -- 1520 - 0x5f0  :  189 - 0xbd -- Sprite 0x5f
    "11111111", -- 1521 - 0x5f1  :  255 - 0xff
    "11111111", -- 1522 - 0x5f2  :  255 - 0xff
    "11111111", -- 1523 - 0x5f3  :  255 - 0xff
    "11111111", -- 1524 - 0x5f4  :  255 - 0xff
    "11111111", -- 1525 - 0x5f5  :  255 - 0xff
    "11111111", -- 1526 - 0x5f6  :  255 - 0xff
    "11111111", -- 1527 - 0x5f7  :  255 - 0xff
    "01111110", -- 1528 - 0x5f8  :  126 - 0x7e -- plane 1
    "01111110", -- 1529 - 0x5f9  :  126 - 0x7e
    "01111110", -- 1530 - 0x5fa  :  126 - 0x7e
    "01111110", -- 1531 - 0x5fb  :  126 - 0x7e
    "01111110", -- 1532 - 0x5fc  :  126 - 0x7e
    "01111110", -- 1533 - 0x5fd  :  126 - 0x7e
    "01111110", -- 1534 - 0x5fe  :  126 - 0x7e
    "01111110", -- 1535 - 0x5ff  :  126 - 0x7e
    "11101110", -- 1536 - 0x600  :  238 - 0xee -- Sprite 0x60
    "00000000", -- 1537 - 0x601  :    0 - 0x0
    "11111110", -- 1538 - 0x602  :  254 - 0xfe
    "00000000", -- 1539 - 0x603  :    0 - 0x0
    "00000001", -- 1540 - 0x604  :    1 - 0x1
    "00001111", -- 1541 - 0x605  :   15 - 0xf
    "10001111", -- 1542 - 0x606  :  143 - 0x8f
    "11111111", -- 1543 - 0x607  :  255 - 0xff
    "11101110", -- 1544 - 0x608  :  238 - 0xee -- plane 1
    "11101110", -- 1545 - 0x609  :  238 - 0xee
    "11111110", -- 1546 - 0x60a  :  254 - 0xfe
    "11111100", -- 1547 - 0x60b  :  252 - 0xfc
    "11100000", -- 1548 - 0x60c  :  224 - 0xe0
    "11100000", -- 1549 - 0x60d  :  224 - 0xe0
    "00000000", -- 1550 - 0x60e  :    0 - 0x0
    "00000000", -- 1551 - 0x60f  :    0 - 0x0
    "11101110", -- 1552 - 0x610  :  238 - 0xee -- Sprite 0x61
    "00000000", -- 1553 - 0x611  :    0 - 0x0
    "11111100", -- 1554 - 0x612  :  252 - 0xfc
    "00000001", -- 1555 - 0x613  :    1 - 0x1
    "00000001", -- 1556 - 0x614  :    1 - 0x1
    "00000000", -- 1557 - 0x615  :    0 - 0x0
    "10001000", -- 1558 - 0x616  :  136 - 0x88
    "11111111", -- 1559 - 0x617  :  255 - 0xff
    "11101110", -- 1560 - 0x618  :  238 - 0xee -- plane 1
    "11101110", -- 1561 - 0x619  :  238 - 0xee
    "11111100", -- 1562 - 0x61a  :  252 - 0xfc
    "11111100", -- 1563 - 0x61b  :  252 - 0xfc
    "11101110", -- 1564 - 0x61c  :  238 - 0xee
    "11101110", -- 1565 - 0x61d  :  238 - 0xee
    "00000000", -- 1566 - 0x61e  :    0 - 0x0
    "00000000", -- 1567 - 0x61f  :    0 - 0x0
    "11100011", -- 1568 - 0x620  :  227 - 0xe3 -- Sprite 0x62
    "00001111", -- 1569 - 0x621  :   15 - 0xf
    "11101111", -- 1570 - 0x622  :  239 - 0xef
    "00001111", -- 1571 - 0x623  :   15 - 0xf
    "00000001", -- 1572 - 0x624  :    1 - 0x1
    "00000000", -- 1573 - 0x625  :    0 - 0x0
    "10000000", -- 1574 - 0x626  :  128 - 0x80
    "11111111", -- 1575 - 0x627  :  255 - 0xff
    "11100000", -- 1576 - 0x628  :  224 - 0xe0 -- plane 1
    "11100000", -- 1577 - 0x629  :  224 - 0xe0
    "11100000", -- 1578 - 0x62a  :  224 - 0xe0
    "11100000", -- 1579 - 0x62b  :  224 - 0xe0
    "11111110", -- 1580 - 0x62c  :  254 - 0xfe
    "11111110", -- 1581 - 0x62d  :  254 - 0xfe
    "00000000", -- 1582 - 0x62e  :    0 - 0x0
    "00000000", -- 1583 - 0x62f  :    0 - 0x0
    "11001110", -- 1584 - 0x630  :  206 - 0xce -- Sprite 0x63
    "11110000", -- 1585 - 0x631  :  240 - 0xf0
    "11111110", -- 1586 - 0x632  :  254 - 0xfe
    "00010000", -- 1587 - 0x633  :   16 - 0x10
    "00000000", -- 1588 - 0x634  :    0 - 0x0
    "10000000", -- 1589 - 0x635  :  128 - 0x80
    "11000001", -- 1590 - 0x636  :  193 - 0xc1
    "11111111", -- 1591 - 0x637  :  255 - 0xff
    "00001110", -- 1592 - 0x638  :   14 - 0xe -- plane 1
    "00001110", -- 1593 - 0x639  :   14 - 0xe
    "00001110", -- 1594 - 0x63a  :   14 - 0xe
    "11101110", -- 1595 - 0x63b  :  238 - 0xee
    "11111110", -- 1596 - 0x63c  :  254 - 0xfe
    "01111100", -- 1597 - 0x63d  :  124 - 0x7c
    "00000000", -- 1598 - 0x63e  :    0 - 0x0
    "00000000", -- 1599 - 0x63f  :    0 - 0x0
    "11111011", -- 1600 - 0x640  :  251 - 0xfb -- Sprite 0x64
    "11000011", -- 1601 - 0x641  :  195 - 0xc3
    "11111011", -- 1602 - 0x642  :  251 - 0xfb
    "11000011", -- 1603 - 0x643  :  195 - 0xc3
    "11000011", -- 1604 - 0x644  :  195 - 0xc3
    "11000011", -- 1605 - 0x645  :  195 - 0xc3
    "11100011", -- 1606 - 0x646  :  227 - 0xe3
    "11111111", -- 1607 - 0x647  :  255 - 0xff
    "00111000", -- 1608 - 0x648  :   56 - 0x38 -- plane 1
    "00111000", -- 1609 - 0x649  :   56 - 0x38
    "00111000", -- 1610 - 0x64a  :   56 - 0x38
    "00111000", -- 1611 - 0x64b  :   56 - 0x38
    "00111000", -- 1612 - 0x64c  :   56 - 0x38
    "00111000", -- 1613 - 0x64d  :   56 - 0x38
    "00000000", -- 1614 - 0x64e  :    0 - 0x0
    "00000000", -- 1615 - 0x64f  :    0 - 0x0
    "11101110", -- 1616 - 0x650  :  238 - 0xee -- Sprite 0x65
    "00000000", -- 1617 - 0x651  :    0 - 0x0
    "11111110", -- 1618 - 0x652  :  254 - 0xfe
    "00000000", -- 1619 - 0x653  :    0 - 0x0
    "00000000", -- 1620 - 0x654  :    0 - 0x0
    "00000000", -- 1621 - 0x655  :    0 - 0x0
    "10001000", -- 1622 - 0x656  :  136 - 0x88
    "11111111", -- 1623 - 0x657  :  255 - 0xff
    "11101110", -- 1624 - 0x658  :  238 - 0xee -- plane 1
    "11101110", -- 1625 - 0x659  :  238 - 0xee
    "11111110", -- 1626 - 0x65a  :  254 - 0xfe
    "11111110", -- 1627 - 0x65b  :  254 - 0xfe
    "11101110", -- 1628 - 0x65c  :  238 - 0xee
    "11101110", -- 1629 - 0x65d  :  238 - 0xee
    "00000000", -- 1630 - 0x65e  :    0 - 0x0
    "00000000", -- 1631 - 0x65f  :    0 - 0x0
    "11101111", -- 1632 - 0x660  :  239 - 0xef -- Sprite 0x66
    "00001111", -- 1633 - 0x661  :   15 - 0xf
    "11101111", -- 1634 - 0x662  :  239 - 0xef
    "00000001", -- 1635 - 0x663  :    1 - 0x1
    "00000000", -- 1636 - 0x664  :    0 - 0x0
    "00000000", -- 1637 - 0x665  :    0 - 0x0
    "10000000", -- 1638 - 0x666  :  128 - 0x80
    "11111111", -- 1639 - 0x667  :  255 - 0xff
    "11100000", -- 1640 - 0x668  :  224 - 0xe0 -- plane 1
    "11100000", -- 1641 - 0x669  :  224 - 0xe0
    "11100000", -- 1642 - 0x66a  :  224 - 0xe0
    "11101110", -- 1643 - 0x66b  :  238 - 0xee
    "11111110", -- 1644 - 0x66c  :  254 - 0xfe
    "11111110", -- 1645 - 0x66d  :  254 - 0xfe
    "00000000", -- 1646 - 0x66e  :    0 - 0x0
    "00000000", -- 1647 - 0x66f  :    0 - 0x0
    "11101110", -- 1648 - 0x670  :  238 - 0xee -- Sprite 0x67
    "00000000", -- 1649 - 0x671  :    0 - 0x0
    "11111110", -- 1650 - 0x672  :  254 - 0xfe
    "00000000", -- 1651 - 0x673  :    0 - 0x0
    "00000000", -- 1652 - 0x674  :    0 - 0x0
    "00001000", -- 1653 - 0x675  :    8 - 0x8
    "10011100", -- 1654 - 0x676  :  156 - 0x9c
    "11111111", -- 1655 - 0x677  :  255 - 0xff
    "11101110", -- 1656 - 0x678  :  238 - 0xee -- plane 1
    "11101110", -- 1657 - 0x679  :  238 - 0xee
    "11111110", -- 1658 - 0x67a  :  254 - 0xfe
    "11111110", -- 1659 - 0x67b  :  254 - 0xfe
    "11101110", -- 1660 - 0x67c  :  238 - 0xee
    "11000110", -- 1661 - 0x67d  :  198 - 0xc6
    "00000000", -- 1662 - 0x67e  :    0 - 0x0
    "00000000", -- 1663 - 0x67f  :    0 - 0x0
    "11101110", -- 1664 - 0x680  :  238 - 0xee -- Sprite 0x68
    "00000000", -- 1665 - 0x681  :    0 - 0x0
    "11101110", -- 1666 - 0x682  :  238 - 0xee
    "00000000", -- 1667 - 0x683  :    0 - 0x0
    "00000000", -- 1668 - 0x684  :    0 - 0x0
    "00000000", -- 1669 - 0x685  :    0 - 0x0
    "10001000", -- 1670 - 0x686  :  136 - 0x88
    "11111111", -- 1671 - 0x687  :  255 - 0xff
    "11101110", -- 1672 - 0x688  :  238 - 0xee -- plane 1
    "11101110", -- 1673 - 0x689  :  238 - 0xee
    "11101110", -- 1674 - 0x68a  :  238 - 0xee
    "11101110", -- 1675 - 0x68b  :  238 - 0xee
    "11101110", -- 1676 - 0x68c  :  238 - 0xee
    "11101110", -- 1677 - 0x68d  :  238 - 0xee
    "00000000", -- 1678 - 0x68e  :    0 - 0x0
    "00000000", -- 1679 - 0x68f  :    0 - 0x0
    "11101110", -- 1680 - 0x690  :  238 - 0xee -- Sprite 0x69
    "00000000", -- 1681 - 0x691  :    0 - 0x0
    "11101110", -- 1682 - 0x692  :  238 - 0xee
    "00000000", -- 1683 - 0x693  :    0 - 0x0
    "00000000", -- 1684 - 0x694  :    0 - 0x0
    "00000000", -- 1685 - 0x695  :    0 - 0x0
    "10000001", -- 1686 - 0x696  :  129 - 0x81
    "11111111", -- 1687 - 0x697  :  255 - 0xff
    "11101110", -- 1688 - 0x698  :  238 - 0xee -- plane 1
    "11101110", -- 1689 - 0x699  :  238 - 0xee
    "11101110", -- 1690 - 0x69a  :  238 - 0xee
    "11101110", -- 1691 - 0x69b  :  238 - 0xee
    "11111110", -- 1692 - 0x69c  :  254 - 0xfe
    "11111100", -- 1693 - 0x69d  :  252 - 0xfc
    "00000000", -- 1694 - 0x69e  :    0 - 0x0
    "00000000", -- 1695 - 0x69f  :    0 - 0x0
    "11101110", -- 1696 - 0x6a0  :  238 - 0xee -- Sprite 0x6a
    "00000000", -- 1697 - 0x6a1  :    0 - 0x0
    "11101110", -- 1698 - 0x6a2  :  238 - 0xee
    "00000000", -- 1699 - 0x6a3  :    0 - 0x0
    "00000000", -- 1700 - 0x6a4  :    0 - 0x0
    "10000000", -- 1701 - 0x6a5  :  128 - 0x80
    "11000001", -- 1702 - 0x6a6  :  193 - 0xc1
    "11111111", -- 1703 - 0x6a7  :  255 - 0xff
    "11101110", -- 1704 - 0x6a8  :  238 - 0xee -- plane 1
    "11101110", -- 1705 - 0x6a9  :  238 - 0xee
    "11101110", -- 1706 - 0x6aa  :  238 - 0xee
    "11101110", -- 1707 - 0x6ab  :  238 - 0xee
    "11111110", -- 1708 - 0x6ac  :  254 - 0xfe
    "01111100", -- 1709 - 0x6ad  :  124 - 0x7c
    "00000000", -- 1710 - 0x6ae  :    0 - 0x0
    "00000000", -- 1711 - 0x6af  :    0 - 0x0
    "11100011", -- 1712 - 0x6b0  :  227 - 0xe3 -- Sprite 0x6b
    "00001111", -- 1713 - 0x6b1  :   15 - 0xf
    "11101111", -- 1714 - 0x6b2  :  239 - 0xef
    "00001111", -- 1715 - 0x6b3  :   15 - 0xf
    "00000001", -- 1716 - 0x6b4  :    1 - 0x1
    "00000000", -- 1717 - 0x6b5  :    0 - 0x0
    "10000000", -- 1718 - 0x6b6  :  128 - 0x80
    "11111111", -- 1719 - 0x6b7  :  255 - 0xff
    "11100000", -- 1720 - 0x6b8  :  224 - 0xe0 -- plane 1
    "11100000", -- 1721 - 0x6b9  :  224 - 0xe0
    "11100000", -- 1722 - 0x6ba  :  224 - 0xe0
    "11100000", -- 1723 - 0x6bb  :  224 - 0xe0
    "11111110", -- 1724 - 0x6bc  :  254 - 0xfe
    "11111110", -- 1725 - 0x6bd  :  254 - 0xfe
    "00000000", -- 1726 - 0x6be  :    0 - 0x0
    "00000000", -- 1727 - 0x6bf  :    0 - 0x0
    "10011001", -- 1728 - 0x6c0  :  153 - 0x99 -- Sprite 0x6c
    "11100011", -- 1729 - 0x6c1  :  227 - 0xe3
    "11110011", -- 1730 - 0x6c2  :  243 - 0xf3
    "11000111", -- 1731 - 0x6c3  :  199 - 0xc7
    "10000001", -- 1732 - 0x6c4  :  129 - 0x81
    "10001000", -- 1733 - 0x6c5  :  136 - 0x88
    "11001100", -- 1734 - 0x6c6  :  204 - 0xcc
    "11111111", -- 1735 - 0x6c7  :  255 - 0xff
    "00011000", -- 1736 - 0x6c8  :   24 - 0x18 -- plane 1
    "00011000", -- 1737 - 0x6c9  :   24 - 0x18
    "00110000", -- 1738 - 0x6ca  :   48 - 0x30
    "00110000", -- 1739 - 0x6cb  :   48 - 0x30
    "01100110", -- 1740 - 0x6cc  :  102 - 0x66
    "01100110", -- 1741 - 0x6cd  :  102 - 0x66
    "00000000", -- 1742 - 0x6ce  :    0 - 0x0
    "00000000", -- 1743 - 0x6cf  :    0 - 0x0
    "11100011", -- 1744 - 0x6d0  :  227 - 0xe3 -- Sprite 0x6d
    "00001111", -- 1745 - 0x6d1  :   15 - 0xf
    "11101111", -- 1746 - 0x6d2  :  239 - 0xef
    "00001111", -- 1747 - 0x6d3  :   15 - 0xf
    "00001111", -- 1748 - 0x6d4  :   15 - 0xf
    "00001111", -- 1749 - 0x6d5  :   15 - 0xf
    "10001111", -- 1750 - 0x6d6  :  143 - 0x8f
    "11111111", -- 1751 - 0x6d7  :  255 - 0xff
    "11100000", -- 1752 - 0x6d8  :  224 - 0xe0 -- plane 1
    "11100000", -- 1753 - 0x6d9  :  224 - 0xe0
    "11100000", -- 1754 - 0x6da  :  224 - 0xe0
    "11100000", -- 1755 - 0x6db  :  224 - 0xe0
    "11100000", -- 1756 - 0x6dc  :  224 - 0xe0
    "11100000", -- 1757 - 0x6dd  :  224 - 0xe0
    "00000000", -- 1758 - 0x6de  :    0 - 0x0
    "00000000", -- 1759 - 0x6df  :    0 - 0x0
    "11101110", -- 1760 - 0x6e0  :  238 - 0xee -- Sprite 0x6e
    "00000000", -- 1761 - 0x6e1  :    0 - 0x0
    "11101110", -- 1762 - 0x6e2  :  238 - 0xee
    "00000000", -- 1763 - 0x6e3  :    0 - 0x0
    "00000000", -- 1764 - 0x6e4  :    0 - 0x0
    "10000000", -- 1765 - 0x6e5  :  128 - 0x80
    "11000001", -- 1766 - 0x6e6  :  193 - 0xc1
    "11111111", -- 1767 - 0x6e7  :  255 - 0xff
    "11101110", -- 1768 - 0x6e8  :  238 - 0xee -- plane 1
    "11101110", -- 1769 - 0x6e9  :  238 - 0xee
    "11101110", -- 1770 - 0x6ea  :  238 - 0xee
    "11101110", -- 1771 - 0x6eb  :  238 - 0xee
    "11111110", -- 1772 - 0x6ec  :  254 - 0xfe
    "01111100", -- 1773 - 0x6ed  :  124 - 0x7c
    "00000000", -- 1774 - 0x6ee  :    0 - 0x0
    "00000000", -- 1775 - 0x6ef  :    0 - 0x0
    "11111111", -- 1776 - 0x6f0  :  255 - 0xff -- Sprite 0x6f
    "11111111", -- 1777 - 0x6f1  :  255 - 0xff
    "11111111", -- 1778 - 0x6f2  :  255 - 0xff
    "10111101", -- 1779 - 0x6f3  :  189 - 0xbd
    "11111111", -- 1780 - 0x6f4  :  255 - 0xff
    "11011011", -- 1781 - 0x6f5  :  219 - 0xdb
    "11111111", -- 1782 - 0x6f6  :  255 - 0xff
    "11111111", -- 1783 - 0x6f7  :  255 - 0xff
    "01111110", -- 1784 - 0x6f8  :  126 - 0x7e -- plane 1
    "01111110", -- 1785 - 0x6f9  :  126 - 0x7e
    "01111110", -- 1786 - 0x6fa  :  126 - 0x7e
    "01111110", -- 1787 - 0x6fb  :  126 - 0x7e
    "00111100", -- 1788 - 0x6fc  :   60 - 0x3c
    "00111100", -- 1789 - 0x6fd  :   60 - 0x3c
    "00000000", -- 1790 - 0x6fe  :    0 - 0x0
    "00000000", -- 1791 - 0x6ff  :    0 - 0x0
    "11111011", -- 1792 - 0x700  :  251 - 0xfb -- Sprite 0x70
    "11101111", -- 1793 - 0x701  :  239 - 0xef
    "11011111", -- 1794 - 0x702  :  223 - 0xdf
    "11111111", -- 1795 - 0x703  :  255 - 0xff
    "10111111", -- 1796 - 0x704  :  191 - 0xbf
    "10111111", -- 1797 - 0x705  :  191 - 0xbf
    "11111110", -- 1798 - 0x706  :  254 - 0xfe
    "11111111", -- 1799 - 0x707  :  255 - 0xff
    "00000111", -- 1800 - 0x708  :    7 - 0x7 -- plane 1
    "00011111", -- 1801 - 0x709  :   31 - 0x1f
    "00111111", -- 1802 - 0x70a  :   63 - 0x3f
    "00111111", -- 1803 - 0x70b  :   63 - 0x3f
    "01111111", -- 1804 - 0x70c  :  127 - 0x7f
    "01111111", -- 1805 - 0x70d  :  127 - 0x7f
    "01111111", -- 1806 - 0x70e  :  127 - 0x7f
    "01111110", -- 1807 - 0x70f  :  126 - 0x7e
    "11011111", -- 1808 - 0x710  :  223 - 0xdf -- Sprite 0x71
    "11110111", -- 1809 - 0x711  :  247 - 0xf7
    "11111011", -- 1810 - 0x712  :  251 - 0xfb
    "11111111", -- 1811 - 0x713  :  255 - 0xff
    "11111101", -- 1812 - 0x714  :  253 - 0xfd
    "11111101", -- 1813 - 0x715  :  253 - 0xfd
    "01111111", -- 1814 - 0x716  :  127 - 0x7f
    "11111111", -- 1815 - 0x717  :  255 - 0xff
    "11100000", -- 1816 - 0x718  :  224 - 0xe0 -- plane 1
    "11111000", -- 1817 - 0x719  :  248 - 0xf8
    "11111100", -- 1818 - 0x71a  :  252 - 0xfc
    "11111100", -- 1819 - 0x71b  :  252 - 0xfc
    "11111110", -- 1820 - 0x71c  :  254 - 0xfe
    "11111110", -- 1821 - 0x71d  :  254 - 0xfe
    "11111110", -- 1822 - 0x71e  :  254 - 0xfe
    "01111110", -- 1823 - 0x71f  :  126 - 0x7e
    "11111111", -- 1824 - 0x720  :  255 - 0xff -- Sprite 0x72
    "11111111", -- 1825 - 0x721  :  255 - 0xff
    "11111111", -- 1826 - 0x722  :  255 - 0xff
    "11111111", -- 1827 - 0x723  :  255 - 0xff
    "11111111", -- 1828 - 0x724  :  255 - 0xff
    "11111111", -- 1829 - 0x725  :  255 - 0xff
    "11111111", -- 1830 - 0x726  :  255 - 0xff
    "11111111", -- 1831 - 0x727  :  255 - 0xff
    "01111110", -- 1832 - 0x728  :  126 - 0x7e -- plane 1
    "01111110", -- 1833 - 0x729  :  126 - 0x7e
    "01111110", -- 1834 - 0x72a  :  126 - 0x7e
    "01111110", -- 1835 - 0x72b  :  126 - 0x7e
    "01111110", -- 1836 - 0x72c  :  126 - 0x7e
    "01111110", -- 1837 - 0x72d  :  126 - 0x7e
    "01111110", -- 1838 - 0x72e  :  126 - 0x7e
    "01111110", -- 1839 - 0x72f  :  126 - 0x7e
    "11111111", -- 1840 - 0x730  :  255 - 0xff -- Sprite 0x73
    "11111110", -- 1841 - 0x731  :  254 - 0xfe
    "10111111", -- 1842 - 0x732  :  191 - 0xbf
    "10111111", -- 1843 - 0x733  :  191 - 0xbf
    "11111111", -- 1844 - 0x734  :  255 - 0xff
    "11011111", -- 1845 - 0x735  :  223 - 0xdf
    "11101111", -- 1846 - 0x736  :  239 - 0xef
    "11111011", -- 1847 - 0x737  :  251 - 0xfb
    "01111110", -- 1848 - 0x738  :  126 - 0x7e -- plane 1
    "01111111", -- 1849 - 0x739  :  127 - 0x7f
    "01111111", -- 1850 - 0x73a  :  127 - 0x7f
    "01111111", -- 1851 - 0x73b  :  127 - 0x7f
    "00111111", -- 1852 - 0x73c  :   63 - 0x3f
    "00111111", -- 1853 - 0x73d  :   63 - 0x3f
    "00011111", -- 1854 - 0x73e  :   31 - 0x1f
    "00000111", -- 1855 - 0x73f  :    7 - 0x7
    "11111111", -- 1856 - 0x740  :  255 - 0xff -- Sprite 0x74
    "01111111", -- 1857 - 0x741  :  127 - 0x7f
    "11111101", -- 1858 - 0x742  :  253 - 0xfd
    "11111101", -- 1859 - 0x743  :  253 - 0xfd
    "11111111", -- 1860 - 0x744  :  255 - 0xff
    "11111011", -- 1861 - 0x745  :  251 - 0xfb
    "11110111", -- 1862 - 0x746  :  247 - 0xf7
    "11011111", -- 1863 - 0x747  :  223 - 0xdf
    "01111110", -- 1864 - 0x748  :  126 - 0x7e -- plane 1
    "11111110", -- 1865 - 0x749  :  254 - 0xfe
    "11111110", -- 1866 - 0x74a  :  254 - 0xfe
    "11111110", -- 1867 - 0x74b  :  254 - 0xfe
    "11111100", -- 1868 - 0x74c  :  252 - 0xfc
    "11111100", -- 1869 - 0x74d  :  252 - 0xfc
    "11111000", -- 1870 - 0x74e  :  248 - 0xf8
    "11100000", -- 1871 - 0x74f  :  224 - 0xe0
    "11111111", -- 1872 - 0x750  :  255 - 0xff -- Sprite 0x75
    "11111111", -- 1873 - 0x751  :  255 - 0xff
    "11111111", -- 1874 - 0x752  :  255 - 0xff
    "11111111", -- 1875 - 0x753  :  255 - 0xff
    "11111111", -- 1876 - 0x754  :  255 - 0xff
    "11111111", -- 1877 - 0x755  :  255 - 0xff
    "11111111", -- 1878 - 0x756  :  255 - 0xff
    "11111111", -- 1879 - 0x757  :  255 - 0xff
    "01111111", -- 1880 - 0x758  :  127 - 0x7f -- plane 1
    "01111111", -- 1881 - 0x759  :  127 - 0x7f
    "01111111", -- 1882 - 0x75a  :  127 - 0x7f
    "01111111", -- 1883 - 0x75b  :  127 - 0x7f
    "01111111", -- 1884 - 0x75c  :  127 - 0x7f
    "01111111", -- 1885 - 0x75d  :  127 - 0x7f
    "00000111", -- 1886 - 0x75e  :    7 - 0x7
    "00000111", -- 1887 - 0x75f  :    7 - 0x7
    "11111111", -- 1888 - 0x760  :  255 - 0xff -- Sprite 0x76
    "11111111", -- 1889 - 0x761  :  255 - 0xff
    "11111111", -- 1890 - 0x762  :  255 - 0xff
    "11111111", -- 1891 - 0x763  :  255 - 0xff
    "11111111", -- 1892 - 0x764  :  255 - 0xff
    "11111111", -- 1893 - 0x765  :  255 - 0xff
    "11111111", -- 1894 - 0x766  :  255 - 0xff
    "11111111", -- 1895 - 0x767  :  255 - 0xff
    "11111110", -- 1896 - 0x768  :  254 - 0xfe -- plane 1
    "11111110", -- 1897 - 0x769  :  254 - 0xfe
    "11111110", -- 1898 - 0x76a  :  254 - 0xfe
    "11111110", -- 1899 - 0x76b  :  254 - 0xfe
    "11111110", -- 1900 - 0x76c  :  254 - 0xfe
    "11111110", -- 1901 - 0x76d  :  254 - 0xfe
    "11100000", -- 1902 - 0x76e  :  224 - 0xe0
    "11100000", -- 1903 - 0x76f  :  224 - 0xe0
    "11111111", -- 1904 - 0x770  :  255 - 0xff -- Sprite 0x77
    "11111111", -- 1905 - 0x771  :  255 - 0xff
    "11111111", -- 1906 - 0x772  :  255 - 0xff
    "11111111", -- 1907 - 0x773  :  255 - 0xff
    "11111111", -- 1908 - 0x774  :  255 - 0xff
    "11111111", -- 1909 - 0x775  :  255 - 0xff
    "11111111", -- 1910 - 0x776  :  255 - 0xff
    "11111111", -- 1911 - 0x777  :  255 - 0xff
    "00000111", -- 1912 - 0x778  :    7 - 0x7 -- plane 1
    "00000111", -- 1913 - 0x779  :    7 - 0x7
    "00000111", -- 1914 - 0x77a  :    7 - 0x7
    "00000111", -- 1915 - 0x77b  :    7 - 0x7
    "00000111", -- 1916 - 0x77c  :    7 - 0x7
    "00000111", -- 1917 - 0x77d  :    7 - 0x7
    "00000111", -- 1918 - 0x77e  :    7 - 0x7
    "00000111", -- 1919 - 0x77f  :    7 - 0x7
    "11111111", -- 1920 - 0x780  :  255 - 0xff -- Sprite 0x78
    "11111111", -- 1921 - 0x781  :  255 - 0xff
    "11111111", -- 1922 - 0x782  :  255 - 0xff
    "11111111", -- 1923 - 0x783  :  255 - 0xff
    "11111111", -- 1924 - 0x784  :  255 - 0xff
    "11111111", -- 1925 - 0x785  :  255 - 0xff
    "11111111", -- 1926 - 0x786  :  255 - 0xff
    "11111111", -- 1927 - 0x787  :  255 - 0xff
    "11100000", -- 1928 - 0x788  :  224 - 0xe0 -- plane 1
    "11100000", -- 1929 - 0x789  :  224 - 0xe0
    "11100000", -- 1930 - 0x78a  :  224 - 0xe0
    "11100000", -- 1931 - 0x78b  :  224 - 0xe0
    "11100000", -- 1932 - 0x78c  :  224 - 0xe0
    "11100000", -- 1933 - 0x78d  :  224 - 0xe0
    "11100000", -- 1934 - 0x78e  :  224 - 0xe0
    "11100000", -- 1935 - 0x78f  :  224 - 0xe0
    "11111111", -- 1936 - 0x790  :  255 - 0xff -- Sprite 0x79
    "11111111", -- 1937 - 0x791  :  255 - 0xff
    "11111111", -- 1938 - 0x792  :  255 - 0xff
    "11111111", -- 1939 - 0x793  :  255 - 0xff
    "11111111", -- 1940 - 0x794  :  255 - 0xff
    "11111111", -- 1941 - 0x795  :  255 - 0xff
    "11111111", -- 1942 - 0x796  :  255 - 0xff
    "11111111", -- 1943 - 0x797  :  255 - 0xff
    "01111111", -- 1944 - 0x798  :  127 - 0x7f -- plane 1
    "01111111", -- 1945 - 0x799  :  127 - 0x7f
    "01111111", -- 1946 - 0x79a  :  127 - 0x7f
    "01111111", -- 1947 - 0x79b  :  127 - 0x7f
    "01111111", -- 1948 - 0x79c  :  127 - 0x7f
    "01111111", -- 1949 - 0x79d  :  127 - 0x7f
    "01111110", -- 1950 - 0x79e  :  126 - 0x7e
    "01111110", -- 1951 - 0x79f  :  126 - 0x7e
    "11111111", -- 1952 - 0x7a0  :  255 - 0xff -- Sprite 0x7a
    "11111111", -- 1953 - 0x7a1  :  255 - 0xff
    "11111111", -- 1954 - 0x7a2  :  255 - 0xff
    "11111111", -- 1955 - 0x7a3  :  255 - 0xff
    "11111111", -- 1956 - 0x7a4  :  255 - 0xff
    "11111111", -- 1957 - 0x7a5  :  255 - 0xff
    "11111111", -- 1958 - 0x7a6  :  255 - 0xff
    "11111111", -- 1959 - 0x7a7  :  255 - 0xff
    "11111110", -- 1960 - 0x7a8  :  254 - 0xfe -- plane 1
    "11111110", -- 1961 - 0x7a9  :  254 - 0xfe
    "11111110", -- 1962 - 0x7aa  :  254 - 0xfe
    "11111110", -- 1963 - 0x7ab  :  254 - 0xfe
    "11111110", -- 1964 - 0x7ac  :  254 - 0xfe
    "11111110", -- 1965 - 0x7ad  :  254 - 0xfe
    "00000000", -- 1966 - 0x7ae  :    0 - 0x0
    "00000000", -- 1967 - 0x7af  :    0 - 0x0
    "11111111", -- 1968 - 0x7b0  :  255 - 0xff -- Sprite 0x7b
    "11111111", -- 1969 - 0x7b1  :  255 - 0xff
    "11111111", -- 1970 - 0x7b2  :  255 - 0xff
    "11111111", -- 1971 - 0x7b3  :  255 - 0xff
    "11111111", -- 1972 - 0x7b4  :  255 - 0xff
    "11111111", -- 1973 - 0x7b5  :  255 - 0xff
    "11111111", -- 1974 - 0x7b6  :  255 - 0xff
    "11111111", -- 1975 - 0x7b7  :  255 - 0xff
    "01111110", -- 1976 - 0x7b8  :  126 - 0x7e -- plane 1
    "01111111", -- 1977 - 0x7b9  :  127 - 0x7f
    "01111111", -- 1978 - 0x7ba  :  127 - 0x7f
    "01111111", -- 1979 - 0x7bb  :  127 - 0x7f
    "01111111", -- 1980 - 0x7bc  :  127 - 0x7f
    "01111111", -- 1981 - 0x7bd  :  127 - 0x7f
    "01111111", -- 1982 - 0x7be  :  127 - 0x7f
    "01111110", -- 1983 - 0x7bf  :  126 - 0x7e
    "11111111", -- 1984 - 0x7c0  :  255 - 0xff -- Sprite 0x7c
    "11111111", -- 1985 - 0x7c1  :  255 - 0xff
    "11111111", -- 1986 - 0x7c2  :  255 - 0xff
    "11111111", -- 1987 - 0x7c3  :  255 - 0xff
    "11111111", -- 1988 - 0x7c4  :  255 - 0xff
    "11111111", -- 1989 - 0x7c5  :  255 - 0xff
    "11111111", -- 1990 - 0x7c6  :  255 - 0xff
    "11111111", -- 1991 - 0x7c7  :  255 - 0xff
    "00000000", -- 1992 - 0x7c8  :    0 - 0x0 -- plane 1
    "11110000", -- 1993 - 0x7c9  :  240 - 0xf0
    "11110000", -- 1994 - 0x7ca  :  240 - 0xf0
    "11110000", -- 1995 - 0x7cb  :  240 - 0xf0
    "11110000", -- 1996 - 0x7cc  :  240 - 0xf0
    "11110000", -- 1997 - 0x7cd  :  240 - 0xf0
    "11110000", -- 1998 - 0x7ce  :  240 - 0xf0
    "00000000", -- 1999 - 0x7cf  :    0 - 0x0
    "11111111", -- 2000 - 0x7d0  :  255 - 0xff -- Sprite 0x7d
    "11111111", -- 2001 - 0x7d1  :  255 - 0xff
    "11111111", -- 2002 - 0x7d2  :  255 - 0xff
    "11111111", -- 2003 - 0x7d3  :  255 - 0xff
    "11111111", -- 2004 - 0x7d4  :  255 - 0xff
    "11111111", -- 2005 - 0x7d5  :  255 - 0xff
    "11111111", -- 2006 - 0x7d6  :  255 - 0xff
    "11111111", -- 2007 - 0x7d7  :  255 - 0xff
    "01111110", -- 2008 - 0x7d8  :  126 - 0x7e -- plane 1
    "01111110", -- 2009 - 0x7d9  :  126 - 0x7e
    "01111111", -- 2010 - 0x7da  :  127 - 0x7f
    "01111111", -- 2011 - 0x7db  :  127 - 0x7f
    "01111111", -- 2012 - 0x7dc  :  127 - 0x7f
    "01111111", -- 2013 - 0x7dd  :  127 - 0x7f
    "01111111", -- 2014 - 0x7de  :  127 - 0x7f
    "01111111", -- 2015 - 0x7df  :  127 - 0x7f
    "11111111", -- 2016 - 0x7e0  :  255 - 0xff -- Sprite 0x7e
    "11111111", -- 2017 - 0x7e1  :  255 - 0xff
    "11111111", -- 2018 - 0x7e2  :  255 - 0xff
    "11111111", -- 2019 - 0x7e3  :  255 - 0xff
    "11111111", -- 2020 - 0x7e4  :  255 - 0xff
    "11111111", -- 2021 - 0x7e5  :  255 - 0xff
    "11111111", -- 2022 - 0x7e6  :  255 - 0xff
    "11111111", -- 2023 - 0x7e7  :  255 - 0xff
    "00000000", -- 2024 - 0x7e8  :    0 - 0x0 -- plane 1
    "00000000", -- 2025 - 0x7e9  :    0 - 0x0
    "11111110", -- 2026 - 0x7ea  :  254 - 0xfe
    "11111110", -- 2027 - 0x7eb  :  254 - 0xfe
    "11111110", -- 2028 - 0x7ec  :  254 - 0xfe
    "11111110", -- 2029 - 0x7ed  :  254 - 0xfe
    "11111110", -- 2030 - 0x7ee  :  254 - 0xfe
    "11111110", -- 2031 - 0x7ef  :  254 - 0xfe
    "11111111", -- 2032 - 0x7f0  :  255 - 0xff -- Sprite 0x7f
    "11111111", -- 2033 - 0x7f1  :  255 - 0xff
    "11111111", -- 2034 - 0x7f2  :  255 - 0xff
    "11111111", -- 2035 - 0x7f3  :  255 - 0xff
    "11111111", -- 2036 - 0x7f4  :  255 - 0xff
    "11111111", -- 2037 - 0x7f5  :  255 - 0xff
    "11111111", -- 2038 - 0x7f6  :  255 - 0xff
    "11111111", -- 2039 - 0x7f7  :  255 - 0xff
    "01111110", -- 2040 - 0x7f8  :  126 - 0x7e -- plane 1
    "11111110", -- 2041 - 0x7f9  :  254 - 0xfe
    "11111110", -- 2042 - 0x7fa  :  254 - 0xfe
    "11111110", -- 2043 - 0x7fb  :  254 - 0xfe
    "11111110", -- 2044 - 0x7fc  :  254 - 0xfe
    "11111110", -- 2045 - 0x7fd  :  254 - 0xfe
    "11111110", -- 2046 - 0x7fe  :  254 - 0xfe
    "01111110", -- 2047 - 0x7ff  :  126 - 0x7e
    "10111111", -- 2048 - 0x800  :  191 - 0xbf -- Sprite 0x80
    "11110111", -- 2049 - 0x801  :  247 - 0xf7
    "11111101", -- 2050 - 0x802  :  253 - 0xfd
    "11011111", -- 2051 - 0x803  :  223 - 0xdf
    "11111011", -- 2052 - 0x804  :  251 - 0xfb
    "10111111", -- 2053 - 0x805  :  191 - 0xbf
    "11111110", -- 2054 - 0x806  :  254 - 0xfe
    "11101111", -- 2055 - 0x807  :  239 - 0xef
    "01000000", -- 2056 - 0x808  :   64 - 0x40 -- plane 1
    "00001000", -- 2057 - 0x809  :    8 - 0x8
    "00000010", -- 2058 - 0x80a  :    2 - 0x2
    "00100000", -- 2059 - 0x80b  :   32 - 0x20
    "00000100", -- 2060 - 0x80c  :    4 - 0x4
    "01000000", -- 2061 - 0x80d  :   64 - 0x40
    "00000001", -- 2062 - 0x80e  :    1 - 0x1
    "00010000", -- 2063 - 0x80f  :   16 - 0x10
    "11111111", -- 2064 - 0x810  :  255 - 0xff -- Sprite 0x81
    "11101110", -- 2065 - 0x811  :  238 - 0xee
    "11111111", -- 2066 - 0x812  :  255 - 0xff
    "11011111", -- 2067 - 0x813  :  223 - 0xdf
    "01110111", -- 2068 - 0x814  :  119 - 0x77
    "11111101", -- 2069 - 0x815  :  253 - 0xfd
    "11011111", -- 2070 - 0x816  :  223 - 0xdf
    "10111111", -- 2071 - 0x817  :  191 - 0xbf
    "00000000", -- 2072 - 0x818  :    0 - 0x0 -- plane 1
    "00010001", -- 2073 - 0x819  :   17 - 0x11
    "00000000", -- 2074 - 0x81a  :    0 - 0x0
    "00100000", -- 2075 - 0x81b  :   32 - 0x20
    "10001000", -- 2076 - 0x81c  :  136 - 0x88
    "00000010", -- 2077 - 0x81d  :    2 - 0x2
    "00100000", -- 2078 - 0x81e  :   32 - 0x20
    "01000000", -- 2079 - 0x81f  :   64 - 0x40
    "11111110", -- 2080 - 0x820  :  254 - 0xfe -- Sprite 0x82
    "11101111", -- 2081 - 0x821  :  239 - 0xef
    "10111111", -- 2082 - 0x822  :  191 - 0xbf
    "11110111", -- 2083 - 0x823  :  247 - 0xf7
    "11111101", -- 2084 - 0x824  :  253 - 0xfd
    "11011111", -- 2085 - 0x825  :  223 - 0xdf
    "11111011", -- 2086 - 0x826  :  251 - 0xfb
    "10111111", -- 2087 - 0x827  :  191 - 0xbf
    "00000001", -- 2088 - 0x828  :    1 - 0x1 -- plane 1
    "00010000", -- 2089 - 0x829  :   16 - 0x10
    "01000000", -- 2090 - 0x82a  :   64 - 0x40
    "00001000", -- 2091 - 0x82b  :    8 - 0x8
    "00000010", -- 2092 - 0x82c  :    2 - 0x2
    "00100000", -- 2093 - 0x82d  :   32 - 0x20
    "00000100", -- 2094 - 0x82e  :    4 - 0x4
    "01000000", -- 2095 - 0x82f  :   64 - 0x40
    "11101111", -- 2096 - 0x830  :  239 - 0xef -- Sprite 0x83
    "11111111", -- 2097 - 0x831  :  255 - 0xff
    "10111011", -- 2098 - 0x832  :  187 - 0xbb
    "11111111", -- 2099 - 0x833  :  255 - 0xff
    "11110111", -- 2100 - 0x834  :  247 - 0xf7
    "11011101", -- 2101 - 0x835  :  221 - 0xdd
    "01111111", -- 2102 - 0x836  :  127 - 0x7f
    "11110111", -- 2103 - 0x837  :  247 - 0xf7
    "00010000", -- 2104 - 0x838  :   16 - 0x10 -- plane 1
    "00000000", -- 2105 - 0x839  :    0 - 0x0
    "01000100", -- 2106 - 0x83a  :   68 - 0x44
    "00000000", -- 2107 - 0x83b  :    0 - 0x0
    "00001000", -- 2108 - 0x83c  :    8 - 0x8
    "00100010", -- 2109 - 0x83d  :   34 - 0x22
    "10000000", -- 2110 - 0x83e  :  128 - 0x80
    "00001000", -- 2111 - 0x83f  :    8 - 0x8
    "11111111", -- 2112 - 0x840  :  255 - 0xff -- Sprite 0x84
    "11101110", -- 2113 - 0x841  :  238 - 0xee
    "11111011", -- 2114 - 0x842  :  251 - 0xfb
    "10111111", -- 2115 - 0x843  :  191 - 0xbf
    "01111111", -- 2116 - 0x844  :  127 - 0x7f
    "11101101", -- 2117 - 0x845  :  237 - 0xed
    "11111111", -- 2118 - 0x846  :  255 - 0xff
    "10111111", -- 2119 - 0x847  :  191 - 0xbf
    "00010100", -- 2120 - 0x848  :   20 - 0x14 -- plane 1
    "10110101", -- 2121 - 0x849  :  181 - 0xb5
    "01000100", -- 2122 - 0x84a  :   68 - 0x44
    "01001010", -- 2123 - 0x84b  :   74 - 0x4a
    "10010010", -- 2124 - 0x84c  :  146 - 0x92
    "10010010", -- 2125 - 0x84d  :  146 - 0x92
    "01000100", -- 2126 - 0x84e  :   68 - 0x44
    "01001001", -- 2127 - 0x84f  :   73 - 0x49
    "11111111", -- 2128 - 0x850  :  255 - 0xff -- Sprite 0x85
    "10111111", -- 2129 - 0x851  :  191 - 0xbf
    "01111101", -- 2130 - 0x852  :  125 - 0x7d
    "11110111", -- 2131 - 0x853  :  247 - 0xf7
    "11011011", -- 2132 - 0x854  :  219 - 0xdb
    "11111101", -- 2133 - 0x855  :  253 - 0xfd
    "01111110", -- 2134 - 0x856  :  126 - 0x7e
    "11111011", -- 2135 - 0x857  :  251 - 0xfb
    "01000010", -- 2136 - 0x858  :   66 - 0x42 -- plane 1
    "01001010", -- 2137 - 0x859  :   74 - 0x4a
    "11001010", -- 2138 - 0x85a  :  202 - 0xca
    "00101001", -- 2139 - 0x85b  :   41 - 0x29
    "10100110", -- 2140 - 0x85c  :  166 - 0xa6
    "10010010", -- 2141 - 0x85d  :  146 - 0x92
    "10001001", -- 2142 - 0x85e  :  137 - 0x89
    "00101101", -- 2143 - 0x85f  :   45 - 0x2d
    "11111111", -- 2144 - 0x860  :  255 - 0xff -- Sprite 0x86
    "11110111", -- 2145 - 0x861  :  247 - 0xf7
    "11111111", -- 2146 - 0x862  :  255 - 0xff
    "11011101", -- 2147 - 0x863  :  221 - 0xdd
    "01111111", -- 2148 - 0x864  :  127 - 0x7f
    "11110111", -- 2149 - 0x865  :  247 - 0xf7
    "11101111", -- 2150 - 0x866  :  239 - 0xef
    "10111101", -- 2151 - 0x867  :  189 - 0xbd
    "10001000", -- 2152 - 0x868  :  136 - 0x88 -- plane 1
    "00101001", -- 2153 - 0x869  :   41 - 0x29
    "10000010", -- 2154 - 0x86a  :  130 - 0x82
    "10110110", -- 2155 - 0x86b  :  182 - 0xb6
    "10001000", -- 2156 - 0x86c  :  136 - 0x88
    "01001001", -- 2157 - 0x86d  :   73 - 0x49
    "01010010", -- 2158 - 0x86e  :   82 - 0x52
    "01010010", -- 2159 - 0x86f  :   82 - 0x52
    "01011111", -- 2160 - 0x870  :   95 - 0x5f -- Sprite 0x87
    "11111101", -- 2161 - 0x871  :  253 - 0xfd
    "11110110", -- 2162 - 0x872  :  246 - 0xf6
    "01111111", -- 2163 - 0x873  :  127 - 0x7f
    "10011111", -- 2164 - 0x874  :  159 - 0x9f
    "11111110", -- 2165 - 0x875  :  254 - 0xfe
    "11111111", -- 2166 - 0x876  :  255 - 0xff
    "11101111", -- 2167 - 0x877  :  239 - 0xef
    "10110010", -- 2168 - 0x878  :  178 - 0xb2 -- plane 1
    "01001010", -- 2169 - 0x879  :   74 - 0x4a
    "10101001", -- 2170 - 0x87a  :  169 - 0xa9
    "10100100", -- 2171 - 0x87b  :  164 - 0xa4
    "01100010", -- 2172 - 0x87c  :   98 - 0x62
    "01001011", -- 2173 - 0x87d  :   75 - 0x4b
    "10010000", -- 2174 - 0x87e  :  144 - 0x90
    "10010010", -- 2175 - 0x87f  :  146 - 0x92
    "11111111", -- 2176 - 0x880  :  255 - 0xff -- Sprite 0x88
    "11111111", -- 2177 - 0x881  :  255 - 0xff
    "10011111", -- 2178 - 0x882  :  159 - 0x9f
    "10110011", -- 2179 - 0x883  :  179 - 0xb3
    "11110011", -- 2180 - 0x884  :  243 - 0xf3
    "11111111", -- 2181 - 0x885  :  255 - 0xff
    "11111111", -- 2182 - 0x886  :  255 - 0xff
    "11111111", -- 2183 - 0x887  :  255 - 0xff
    "00000000", -- 2184 - 0x888  :    0 - 0x0 -- plane 1
    "01100000", -- 2185 - 0x889  :   96 - 0x60
    "11111110", -- 2186 - 0x88a  :  254 - 0xfe
    "11111111", -- 2187 - 0x88b  :  255 - 0xff
    "01111111", -- 2188 - 0x88c  :  127 - 0x7f
    "00011111", -- 2189 - 0x88d  :   31 - 0x1f
    "00001110", -- 2190 - 0x88e  :   14 - 0xe
    "00000000", -- 2191 - 0x88f  :    0 - 0x0
    "11111111", -- 2192 - 0x890  :  255 - 0xff -- Sprite 0x89
    "11001111", -- 2193 - 0x891  :  207 - 0xcf
    "11011111", -- 2194 - 0x892  :  223 - 0xdf
    "11111111", -- 2195 - 0x893  :  255 - 0xff
    "11110011", -- 2196 - 0x894  :  243 - 0xf3
    "11110011", -- 2197 - 0x895  :  243 - 0xf3
    "11111111", -- 2198 - 0x896  :  255 - 0xff
    "11111111", -- 2199 - 0x897  :  255 - 0xff
    "00110000", -- 2200 - 0x898  :   48 - 0x30 -- plane 1
    "01111000", -- 2201 - 0x899  :  120 - 0x78
    "01111000", -- 2202 - 0x89a  :  120 - 0x78
    "00111110", -- 2203 - 0x89b  :   62 - 0x3e
    "00011111", -- 2204 - 0x89c  :   31 - 0x1f
    "00011111", -- 2205 - 0x89d  :   31 - 0x1f
    "00011111", -- 2206 - 0x89e  :   31 - 0x1f
    "00001110", -- 2207 - 0x89f  :   14 - 0xe
    "10111111", -- 2208 - 0x8a0  :  191 - 0xbf -- Sprite 0x8a
    "11110111", -- 2209 - 0x8a1  :  247 - 0xf7
    "11111101", -- 2210 - 0x8a2  :  253 - 0xfd
    "11111111", -- 2211 - 0x8a3  :  255 - 0xff
    "11111011", -- 2212 - 0x8a4  :  251 - 0xfb
    "10111111", -- 2213 - 0x8a5  :  191 - 0xbf
    "11111110", -- 2214 - 0x8a6  :  254 - 0xfe
    "11101111", -- 2215 - 0x8a7  :  239 - 0xef
    "01000000", -- 2216 - 0x8a8  :   64 - 0x40 -- plane 1
    "00001000", -- 2217 - 0x8a9  :    8 - 0x8
    "00000010", -- 2218 - 0x8aa  :    2 - 0x2
    "00101000", -- 2219 - 0x8ab  :   40 - 0x28
    "00010100", -- 2220 - 0x8ac  :   20 - 0x14
    "01010100", -- 2221 - 0x8ad  :   84 - 0x54
    "00000001", -- 2222 - 0x8ae  :    1 - 0x1
    "00010000", -- 2223 - 0x8af  :   16 - 0x10
    "10111111", -- 2224 - 0x8b0  :  191 - 0xbf -- Sprite 0x8b
    "11111111", -- 2225 - 0x8b1  :  255 - 0xff
    "11101110", -- 2226 - 0x8b2  :  238 - 0xee
    "11111111", -- 2227 - 0x8b3  :  255 - 0xff
    "11011111", -- 2228 - 0x8b4  :  223 - 0xdf
    "01111101", -- 2229 - 0x8b5  :  125 - 0x7d
    "11111111", -- 2230 - 0x8b6  :  255 - 0xff
    "11011111", -- 2231 - 0x8b7  :  223 - 0xdf
    "01000000", -- 2232 - 0x8b8  :   64 - 0x40 -- plane 1
    "00000000", -- 2233 - 0x8b9  :    0 - 0x0
    "10010001", -- 2234 - 0x8ba  :  145 - 0x91
    "00010100", -- 2235 - 0x8bb  :   20 - 0x14
    "00101000", -- 2236 - 0x8bc  :   40 - 0x28
    "10001010", -- 2237 - 0x8bd  :  138 - 0x8a
    "01000000", -- 2238 - 0x8be  :   64 - 0x40
    "00100000", -- 2239 - 0x8bf  :   32 - 0x20
    "11111111", -- 2240 - 0x8c0  :  255 - 0xff -- Sprite 0x8c
    "11111000", -- 2241 - 0x8c1  :  248 - 0xf8
    "11100010", -- 2242 - 0x8c2  :  226 - 0xe2
    "11010111", -- 2243 - 0x8c3  :  215 - 0xd7
    "11001111", -- 2244 - 0x8c4  :  207 - 0xcf
    "10011111", -- 2245 - 0x8c5  :  159 - 0x9f
    "10111110", -- 2246 - 0x8c6  :  190 - 0xbe
    "10011101", -- 2247 - 0x8c7  :  157 - 0x9d
    "00000000", -- 2248 - 0x8c8  :    0 - 0x0 -- plane 1
    "00000111", -- 2249 - 0x8c9  :    7 - 0x7
    "00011111", -- 2250 - 0x8ca  :   31 - 0x1f
    "00111111", -- 2251 - 0x8cb  :   63 - 0x3f
    "00111111", -- 2252 - 0x8cc  :   63 - 0x3f
    "01111111", -- 2253 - 0x8cd  :  127 - 0x7f
    "01111111", -- 2254 - 0x8ce  :  127 - 0x7f
    "01111111", -- 2255 - 0x8cf  :  127 - 0x7f
    "11111111", -- 2256 - 0x8d0  :  255 - 0xff -- Sprite 0x8d
    "00011111", -- 2257 - 0x8d1  :   31 - 0x1f
    "10100111", -- 2258 - 0x8d2  :  167 - 0xa7
    "11000011", -- 2259 - 0x8d3  :  195 - 0xc3
    "11100011", -- 2260 - 0x8d4  :  227 - 0xe3
    "01000001", -- 2261 - 0x8d5  :   65 - 0x41
    "10100001", -- 2262 - 0x8d6  :  161 - 0xa1
    "00000001", -- 2263 - 0x8d7  :    1 - 0x1
    "00000000", -- 2264 - 0x8d8  :    0 - 0x0 -- plane 1
    "11100000", -- 2265 - 0x8d9  :  224 - 0xe0
    "11111000", -- 2266 - 0x8da  :  248 - 0xf8
    "11111000", -- 2267 - 0x8db  :  248 - 0xf8
    "11110000", -- 2268 - 0x8dc  :  240 - 0xf0
    "11111000", -- 2269 - 0x8dd  :  248 - 0xf8
    "11110100", -- 2270 - 0x8de  :  244 - 0xf4
    "11111000", -- 2271 - 0x8df  :  248 - 0xf8
    "10111110", -- 2272 - 0x8e0  :  190 - 0xbe -- Sprite 0x8e
    "11111111", -- 2273 - 0x8e1  :  255 - 0xff
    "11011111", -- 2274 - 0x8e2  :  223 - 0xdf
    "11111111", -- 2275 - 0x8e3  :  255 - 0xff
    "11101111", -- 2276 - 0x8e4  :  239 - 0xef
    "11111111", -- 2277 - 0x8e5  :  255 - 0xff
    "11110111", -- 2278 - 0x8e6  :  247 - 0xf7
    "11111111", -- 2279 - 0x8e7  :  255 - 0xff
    "01111111", -- 2280 - 0x8e8  :  127 - 0x7f -- plane 1
    "00111111", -- 2281 - 0x8e9  :   63 - 0x3f
    "00111111", -- 2282 - 0x8ea  :   63 - 0x3f
    "00011111", -- 2283 - 0x8eb  :   31 - 0x1f
    "00011111", -- 2284 - 0x8ec  :   31 - 0x1f
    "00001111", -- 2285 - 0x8ed  :   15 - 0xf
    "00001111", -- 2286 - 0x8ee  :   15 - 0xf
    "00000111", -- 2287 - 0x8ef  :    7 - 0x7
    "01111101", -- 2288 - 0x8f0  :  125 - 0x7d -- Sprite 0x8f
    "11111111", -- 2289 - 0x8f1  :  255 - 0xff
    "11111011", -- 2290 - 0x8f2  :  251 - 0xfb
    "11111111", -- 2291 - 0x8f3  :  255 - 0xff
    "11110111", -- 2292 - 0x8f4  :  247 - 0xf7
    "11111111", -- 2293 - 0x8f5  :  255 - 0xff
    "11101111", -- 2294 - 0x8f6  :  239 - 0xef
    "11111111", -- 2295 - 0x8f7  :  255 - 0xff
    "11111110", -- 2296 - 0x8f8  :  254 - 0xfe -- plane 1
    "11111100", -- 2297 - 0x8f9  :  252 - 0xfc
    "11111100", -- 2298 - 0x8fa  :  252 - 0xfc
    "11111000", -- 2299 - 0x8fb  :  248 - 0xf8
    "11111000", -- 2300 - 0x8fc  :  248 - 0xf8
    "11110000", -- 2301 - 0x8fd  :  240 - 0xf0
    "11110000", -- 2302 - 0x8fe  :  240 - 0xf0
    "11100000", -- 2303 - 0x8ff  :  224 - 0xe0
    "10111110", -- 2304 - 0x900  :  190 - 0xbe -- Sprite 0x90
    "11110111", -- 2305 - 0x901  :  247 - 0xf7
    "11111111", -- 2306 - 0x902  :  255 - 0xff
    "11011111", -- 2307 - 0x903  :  223 - 0xdf
    "11111011", -- 2308 - 0x904  :  251 - 0xfb
    "11111110", -- 2309 - 0x905  :  254 - 0xfe
    "10111111", -- 2310 - 0x906  :  191 - 0xbf
    "11110111", -- 2311 - 0x907  :  247 - 0xf7
    "01000001", -- 2312 - 0x908  :   65 - 0x41 -- plane 1
    "00001000", -- 2313 - 0x909  :    8 - 0x8
    "00000000", -- 2314 - 0x90a  :    0 - 0x0
    "00100000", -- 2315 - 0x90b  :   32 - 0x20
    "00000100", -- 2316 - 0x90c  :    4 - 0x4
    "00000001", -- 2317 - 0x90d  :    1 - 0x1
    "01000000", -- 2318 - 0x90e  :   64 - 0x40
    "00001000", -- 2319 - 0x90f  :    8 - 0x8
    "11101110", -- 2320 - 0x910  :  238 - 0xee -- Sprite 0x91
    "11111111", -- 2321 - 0x911  :  255 - 0xff
    "01111011", -- 2322 - 0x912  :  123 - 0x7b
    "11111101", -- 2323 - 0x913  :  253 - 0xfd
    "11101111", -- 2324 - 0x914  :  239 - 0xef
    "11111111", -- 2325 - 0x915  :  255 - 0xff
    "10111101", -- 2326 - 0x916  :  189 - 0xbd
    "11111111", -- 2327 - 0x917  :  255 - 0xff
    "00010001", -- 2328 - 0x918  :   17 - 0x11 -- plane 1
    "00000000", -- 2329 - 0x919  :    0 - 0x0
    "10000100", -- 2330 - 0x91a  :  132 - 0x84
    "00000010", -- 2331 - 0x91b  :    2 - 0x2
    "00010000", -- 2332 - 0x91c  :   16 - 0x10
    "00000000", -- 2333 - 0x91d  :    0 - 0x0
    "01000010", -- 2334 - 0x91e  :   66 - 0x42
    "00000000", -- 2335 - 0x91f  :    0 - 0x0
    "11111011", -- 2336 - 0x920  :  251 - 0xfb -- Sprite 0x92
    "10111111", -- 2337 - 0x921  :  191 - 0xbf
    "11101111", -- 2338 - 0x922  :  239 - 0xef
    "11111101", -- 2339 - 0x923  :  253 - 0xfd
    "11111111", -- 2340 - 0x924  :  255 - 0xff
    "10111111", -- 2341 - 0x925  :  191 - 0xbf
    "11111011", -- 2342 - 0x926  :  251 - 0xfb
    "11011111", -- 2343 - 0x927  :  223 - 0xdf
    "00000100", -- 2344 - 0x928  :    4 - 0x4 -- plane 1
    "01000000", -- 2345 - 0x929  :   64 - 0x40
    "00010000", -- 2346 - 0x92a  :   16 - 0x10
    "00000010", -- 2347 - 0x92b  :    2 - 0x2
    "00000000", -- 2348 - 0x92c  :    0 - 0x0
    "01000000", -- 2349 - 0x92d  :   64 - 0x40
    "00000100", -- 2350 - 0x92e  :    4 - 0x4
    "00100000", -- 2351 - 0x92f  :   32 - 0x20
    "10111101", -- 2352 - 0x930  :  189 - 0xbd -- Sprite 0x93
    "11111111", -- 2353 - 0x931  :  255 - 0xff
    "01110111", -- 2354 - 0x932  :  119 - 0x77
    "11111110", -- 2355 - 0x933  :  254 - 0xfe
    "11011111", -- 2356 - 0x934  :  223 - 0xdf
    "11111011", -- 2357 - 0x935  :  251 - 0xfb
    "11101111", -- 2358 - 0x936  :  239 - 0xef
    "01111111", -- 2359 - 0x937  :  127 - 0x7f
    "01000010", -- 2360 - 0x938  :   66 - 0x42 -- plane 1
    "00000000", -- 2361 - 0x939  :    0 - 0x0
    "10001000", -- 2362 - 0x93a  :  136 - 0x88
    "00000001", -- 2363 - 0x93b  :    1 - 0x1
    "00100000", -- 2364 - 0x93c  :   32 - 0x20
    "00000100", -- 2365 - 0x93d  :    4 - 0x4
    "00010000", -- 2366 - 0x93e  :   16 - 0x10
    "10000000", -- 2367 - 0x93f  :  128 - 0x80
    "01111111", -- 2368 - 0x940  :  127 - 0x7f -- Sprite 0x94
    "11110111", -- 2369 - 0x941  :  247 - 0xf7
    "11011101", -- 2370 - 0x942  :  221 - 0xdd
    "01111011", -- 2371 - 0x943  :  123 - 0x7b
    "11111111", -- 2372 - 0x944  :  255 - 0xff
    "11101110", -- 2373 - 0x945  :  238 - 0xee
    "10111011", -- 2374 - 0x946  :  187 - 0xbb
    "11111101", -- 2375 - 0x947  :  253 - 0xfd
    "11001000", -- 2376 - 0x948  :  200 - 0xc8 -- plane 1
    "00101010", -- 2377 - 0x949  :   42 - 0x2a
    "10100010", -- 2378 - 0x94a  :  162 - 0xa2
    "10010100", -- 2379 - 0x94b  :  148 - 0x94
    "10010001", -- 2380 - 0x94c  :  145 - 0x91
    "01010101", -- 2381 - 0x94d  :   85 - 0x55
    "01000100", -- 2382 - 0x94e  :   68 - 0x44
    "00010010", -- 2383 - 0x94f  :   18 - 0x12
    "11010111", -- 2384 - 0x950  :  215 - 0xd7 -- Sprite 0x95
    "01111111", -- 2385 - 0x951  :  127 - 0x7f
    "11111101", -- 2386 - 0x952  :  253 - 0xfd
    "11101110", -- 2387 - 0x953  :  238 - 0xee
    "11110111", -- 2388 - 0x954  :  247 - 0xf7
    "10111011", -- 2389 - 0x955  :  187 - 0xbb
    "11101111", -- 2390 - 0x956  :  239 - 0xef
    "11110111", -- 2391 - 0x957  :  247 - 0xf7
    "10101010", -- 2392 - 0x958  :  170 - 0xaa -- plane 1
    "10100010", -- 2393 - 0x959  :  162 - 0xa2
    "00010010", -- 2394 - 0x95a  :   18 - 0x12
    "01010011", -- 2395 - 0x95b  :   83 - 0x53
    "01001100", -- 2396 - 0x95c  :   76 - 0x4c
    "01010101", -- 2397 - 0x95d  :   85 - 0x55
    "10010001", -- 2398 - 0x95e  :  145 - 0x91
    "01001000", -- 2399 - 0x95f  :   72 - 0x48
    "10111111", -- 2400 - 0x960  :  191 - 0xbf -- Sprite 0x96
    "11101110", -- 2401 - 0x961  :  238 - 0xee
    "11011011", -- 2402 - 0x962  :  219 - 0xdb
    "11111111", -- 2403 - 0x963  :  255 - 0xff
    "01110111", -- 2404 - 0x964  :  119 - 0x77
    "11011101", -- 2405 - 0x965  :  221 - 0xdd
    "11101111", -- 2406 - 0x966  :  239 - 0xef
    "11111011", -- 2407 - 0x967  :  251 - 0xfb
    "01010001", -- 2408 - 0x968  :   81 - 0x51 -- plane 1
    "00010101", -- 2409 - 0x969  :   21 - 0x15
    "10100100", -- 2410 - 0x96a  :  164 - 0xa4
    "10001100", -- 2411 - 0x96b  :  140 - 0x8c
    "10101010", -- 2412 - 0x96c  :  170 - 0xaa
    "00100010", -- 2413 - 0x96d  :   34 - 0x22
    "10010000", -- 2414 - 0x96e  :  144 - 0x90
    "01000110", -- 2415 - 0x96f  :   70 - 0x46
    "11111101", -- 2416 - 0x970  :  253 - 0xfd -- Sprite 0x97
    "11101110", -- 2417 - 0x971  :  238 - 0xee
    "11111011", -- 2418 - 0x972  :  251 - 0xfb
    "11111101", -- 2419 - 0x973  :  253 - 0xfd
    "11110101", -- 2420 - 0x974  :  245 - 0xf5
    "11011111", -- 2421 - 0x975  :  223 - 0xdf
    "01111111", -- 2422 - 0x976  :  127 - 0x7f
    "10111011", -- 2423 - 0x977  :  187 - 0xbb
    "00010011", -- 2424 - 0x978  :   19 - 0x13 -- plane 1
    "01010101", -- 2425 - 0x979  :   85 - 0x55
    "01100100", -- 2426 - 0x97a  :  100 - 0x64
    "00010010", -- 2427 - 0x97b  :   18 - 0x12
    "10101010", -- 2428 - 0x97c  :  170 - 0xaa
    "10101000", -- 2429 - 0x97d  :  168 - 0xa8
    "10000100", -- 2430 - 0x97e  :  132 - 0x84
    "11010100", -- 2431 - 0x97f  :  212 - 0xd4
    "11111111", -- 2432 - 0x980  :  255 - 0xff -- Sprite 0x98
    "11001111", -- 2433 - 0x981  :  207 - 0xcf
    "11011111", -- 2434 - 0x982  :  223 - 0xdf
    "11111111", -- 2435 - 0x983  :  255 - 0xff
    "11110011", -- 2436 - 0x984  :  243 - 0xf3
    "11110011", -- 2437 - 0x985  :  243 - 0xf3
    "11111111", -- 2438 - 0x986  :  255 - 0xff
    "11111111", -- 2439 - 0x987  :  255 - 0xff
    "00110000", -- 2440 - 0x988  :   48 - 0x30 -- plane 1
    "01111000", -- 2441 - 0x989  :  120 - 0x78
    "01111000", -- 2442 - 0x98a  :  120 - 0x78
    "00111110", -- 2443 - 0x98b  :   62 - 0x3e
    "00011111", -- 2444 - 0x98c  :   31 - 0x1f
    "00011111", -- 2445 - 0x98d  :   31 - 0x1f
    "00011111", -- 2446 - 0x98e  :   31 - 0x1f
    "00001110", -- 2447 - 0x98f  :   14 - 0xe
    "11111111", -- 2448 - 0x990  :  255 - 0xff -- Sprite 0x99
    "11111111", -- 2449 - 0x991  :  255 - 0xff
    "10011111", -- 2450 - 0x992  :  159 - 0x9f
    "10110011", -- 2451 - 0x993  :  179 - 0xb3
    "11110011", -- 2452 - 0x994  :  243 - 0xf3
    "11111111", -- 2453 - 0x995  :  255 - 0xff
    "11111111", -- 2454 - 0x996  :  255 - 0xff
    "11111111", -- 2455 - 0x997  :  255 - 0xff
    "00000000", -- 2456 - 0x998  :    0 - 0x0 -- plane 1
    "01100000", -- 2457 - 0x999  :   96 - 0x60
    "11111110", -- 2458 - 0x99a  :  254 - 0xfe
    "11111111", -- 2459 - 0x99b  :  255 - 0xff
    "01111111", -- 2460 - 0x99c  :  127 - 0x7f
    "00011111", -- 2461 - 0x99d  :   31 - 0x1f
    "00001110", -- 2462 - 0x99e  :   14 - 0xe
    "00000000", -- 2463 - 0x99f  :    0 - 0x0
    "10111111", -- 2464 - 0x9a0  :  191 - 0xbf -- Sprite 0x9a
    "11110111", -- 2465 - 0x9a1  :  247 - 0xf7
    "11111111", -- 2466 - 0x9a2  :  255 - 0xff
    "11011111", -- 2467 - 0x9a3  :  223 - 0xdf
    "11111011", -- 2468 - 0x9a4  :  251 - 0xfb
    "11111111", -- 2469 - 0x9a5  :  255 - 0xff
    "10111111", -- 2470 - 0x9a6  :  191 - 0xbf
    "11110111", -- 2471 - 0x9a7  :  247 - 0xf7
    "01000000", -- 2472 - 0x9a8  :   64 - 0x40 -- plane 1
    "00001100", -- 2473 - 0x9a9  :   12 - 0xc
    "00000000", -- 2474 - 0x9aa  :    0 - 0x0
    "00101000", -- 2475 - 0x9ab  :   40 - 0x28
    "00101100", -- 2476 - 0x9ac  :   44 - 0x2c
    "00010001", -- 2477 - 0x9ad  :   17 - 0x11
    "01000000", -- 2478 - 0x9ae  :   64 - 0x40
    "00001000", -- 2479 - 0x9af  :    8 - 0x8
    "11011111", -- 2480 - 0x9b0  :  223 - 0xdf -- Sprite 0x9b
    "11111111", -- 2481 - 0x9b1  :  255 - 0xff
    "01111011", -- 2482 - 0x9b2  :  123 - 0x7b
    "11111111", -- 2483 - 0x9b3  :  255 - 0xff
    "11101111", -- 2484 - 0x9b4  :  239 - 0xef
    "11111101", -- 2485 - 0x9b5  :  253 - 0xfd
    "10111111", -- 2486 - 0x9b6  :  191 - 0xbf
    "11111111", -- 2487 - 0x9b7  :  255 - 0xff
    "00100000", -- 2488 - 0x9b8  :   32 - 0x20 -- plane 1
    "00000000", -- 2489 - 0x9b9  :    0 - 0x0
    "10010100", -- 2490 - 0x9ba  :  148 - 0x94
    "01001000", -- 2491 - 0x9bb  :   72 - 0x48
    "00011000", -- 2492 - 0x9bc  :   24 - 0x18
    "00000110", -- 2493 - 0x9bd  :    6 - 0x6
    "01000000", -- 2494 - 0x9be  :   64 - 0x40
    "00000000", -- 2495 - 0x9bf  :    0 - 0x0
    "10111010", -- 2496 - 0x9c0  :  186 - 0xba -- Sprite 0x9c
    "10011100", -- 2497 - 0x9c1  :  156 - 0x9c
    "10101010", -- 2498 - 0x9c2  :  170 - 0xaa
    "11000000", -- 2499 - 0x9c3  :  192 - 0xc0
    "11000000", -- 2500 - 0x9c4  :  192 - 0xc0
    "11100000", -- 2501 - 0x9c5  :  224 - 0xe0
    "11111000", -- 2502 - 0x9c6  :  248 - 0xf8
    "11111111", -- 2503 - 0x9c7  :  255 - 0xff
    "01111111", -- 2504 - 0x9c8  :  127 - 0x7f -- plane 1
    "01111111", -- 2505 - 0x9c9  :  127 - 0x7f
    "01111111", -- 2506 - 0x9ca  :  127 - 0x7f
    "00111111", -- 2507 - 0x9cb  :   63 - 0x3f
    "00110101", -- 2508 - 0x9cc  :   53 - 0x35
    "00000010", -- 2509 - 0x9cd  :    2 - 0x2
    "00000000", -- 2510 - 0x9ce  :    0 - 0x0
    "00000000", -- 2511 - 0x9cf  :    0 - 0x0
    "00000001", -- 2512 - 0x9d0  :    1 - 0x1 -- Sprite 0x9d
    "00000001", -- 2513 - 0x9d1  :    1 - 0x1
    "00000001", -- 2514 - 0x9d2  :    1 - 0x1
    "00000011", -- 2515 - 0x9d3  :    3 - 0x3
    "00000011", -- 2516 - 0x9d4  :    3 - 0x3
    "00000111", -- 2517 - 0x9d5  :    7 - 0x7
    "00011111", -- 2518 - 0x9d6  :   31 - 0x1f
    "11111111", -- 2519 - 0x9d7  :  255 - 0xff
    "11110100", -- 2520 - 0x9d8  :  244 - 0xf4 -- plane 1
    "11111000", -- 2521 - 0x9d9  :  248 - 0xf8
    "11110000", -- 2522 - 0x9da  :  240 - 0xf0
    "11101000", -- 2523 - 0x9db  :  232 - 0xe8
    "01010000", -- 2524 - 0x9dc  :   80 - 0x50
    "10000000", -- 2525 - 0x9dd  :  128 - 0x80
    "00000000", -- 2526 - 0x9de  :    0 - 0x0
    "00000000", -- 2527 - 0x9df  :    0 - 0x0
    "01111101", -- 2528 - 0x9e0  :  125 - 0x7d -- Sprite 0x9e
    "11111111", -- 2529 - 0x9e1  :  255 - 0xff
    "11111011", -- 2530 - 0x9e2  :  251 - 0xfb
    "11111111", -- 2531 - 0x9e3  :  255 - 0xff
    "11111111", -- 2532 - 0x9e4  :  255 - 0xff
    "11111011", -- 2533 - 0x9e5  :  251 - 0xfb
    "11111111", -- 2534 - 0x9e6  :  255 - 0xff
    "01111101", -- 2535 - 0x9e7  :  125 - 0x7d
    "11111110", -- 2536 - 0x9e8  :  254 - 0xfe -- plane 1
    "11111100", -- 2537 - 0x9e9  :  252 - 0xfc
    "11111100", -- 2538 - 0x9ea  :  252 - 0xfc
    "11111000", -- 2539 - 0x9eb  :  248 - 0xf8
    "11111000", -- 2540 - 0x9ec  :  248 - 0xf8
    "11111100", -- 2541 - 0x9ed  :  252 - 0xfc
    "11111100", -- 2542 - 0x9ee  :  252 - 0xfc
    "11111110", -- 2543 - 0x9ef  :  254 - 0xfe
    "11111111", -- 2544 - 0x9f0  :  255 - 0xff -- Sprite 0x9f
    "11111111", -- 2545 - 0x9f1  :  255 - 0xff
    "10111101", -- 2546 - 0x9f2  :  189 - 0xbd
    "11111111", -- 2547 - 0x9f3  :  255 - 0xff
    "11111111", -- 2548 - 0x9f4  :  255 - 0xff
    "11111111", -- 2549 - 0x9f5  :  255 - 0xff
    "11111111", -- 2550 - 0x9f6  :  255 - 0xff
    "10111101", -- 2551 - 0x9f7  :  189 - 0xbd
    "00000000", -- 2552 - 0x9f8  :    0 - 0x0 -- plane 1
    "00000000", -- 2553 - 0x9f9  :    0 - 0x0
    "01111110", -- 2554 - 0x9fa  :  126 - 0x7e
    "01111110", -- 2555 - 0x9fb  :  126 - 0x7e
    "01111110", -- 2556 - 0x9fc  :  126 - 0x7e
    "01111110", -- 2557 - 0x9fd  :  126 - 0x7e
    "01111110", -- 2558 - 0x9fe  :  126 - 0x7e
    "01111110", -- 2559 - 0x9ff  :  126 - 0x7e
    "11101111", -- 2560 - 0xa00  :  239 - 0xef -- Sprite 0xa0
    "11000111", -- 2561 - 0xa01  :  199 - 0xc7
    "10000011", -- 2562 - 0xa02  :  131 - 0x83
    "00000111", -- 2563 - 0xa03  :    7 - 0x7
    "10001111", -- 2564 - 0xa04  :  143 - 0x8f
    "11011101", -- 2565 - 0xa05  :  221 - 0xdd
    "11111010", -- 2566 - 0xa06  :  250 - 0xfa
    "11111101", -- 2567 - 0xa07  :  253 - 0xfd
    "00010000", -- 2568 - 0xa08  :   16 - 0x10 -- plane 1
    "00111000", -- 2569 - 0xa09  :   56 - 0x38
    "01111100", -- 2570 - 0xa0a  :  124 - 0x7c
    "11111000", -- 2571 - 0xa0b  :  248 - 0xf8
    "01110000", -- 2572 - 0xa0c  :  112 - 0x70
    "00100010", -- 2573 - 0xa0d  :   34 - 0x22
    "00000101", -- 2574 - 0xa0e  :    5 - 0x5
    "00000010", -- 2575 - 0xa0f  :    2 - 0x2
    "11101111", -- 2576 - 0xa10  :  239 - 0xef -- Sprite 0xa1
    "11000111", -- 2577 - 0xa11  :  199 - 0xc7
    "10000011", -- 2578 - 0xa12  :  131 - 0x83
    "00011111", -- 2579 - 0xa13  :   31 - 0x1f
    "10010000", -- 2580 - 0xa14  :  144 - 0x90
    "11010100", -- 2581 - 0xa15  :  212 - 0xd4
    "11110011", -- 2582 - 0xa16  :  243 - 0xf3
    "11110010", -- 2583 - 0xa17  :  242 - 0xf2
    "00010000", -- 2584 - 0xa18  :   16 - 0x10 -- plane 1
    "00111000", -- 2585 - 0xa19  :   56 - 0x38
    "01111100", -- 2586 - 0xa1a  :  124 - 0x7c
    "11100000", -- 2587 - 0xa1b  :  224 - 0xe0
    "01100000", -- 2588 - 0xa1c  :   96 - 0x60
    "00100000", -- 2589 - 0xa1d  :   32 - 0x20
    "00000000", -- 2590 - 0xa1e  :    0 - 0x0
    "00000000", -- 2591 - 0xa1f  :    0 - 0x0
    "11101111", -- 2592 - 0xa20  :  239 - 0xef -- Sprite 0xa2
    "11000111", -- 2593 - 0xa21  :  199 - 0xc7
    "10000011", -- 2594 - 0xa22  :  131 - 0x83
    "11111111", -- 2595 - 0xa23  :  255 - 0xff
    "00000000", -- 2596 - 0xa24  :    0 - 0x0
    "00000000", -- 2597 - 0xa25  :    0 - 0x0
    "01010101", -- 2598 - 0xa26  :   85 - 0x55
    "00000000", -- 2599 - 0xa27  :    0 - 0x0
    "00010000", -- 2600 - 0xa28  :   16 - 0x10 -- plane 1
    "00111000", -- 2601 - 0xa29  :   56 - 0x38
    "01111100", -- 2602 - 0xa2a  :  124 - 0x7c
    "00000000", -- 2603 - 0xa2b  :    0 - 0x0
    "00000000", -- 2604 - 0xa2c  :    0 - 0x0
    "00000000", -- 2605 - 0xa2d  :    0 - 0x0
    "00000000", -- 2606 - 0xa2e  :    0 - 0x0
    "00000000", -- 2607 - 0xa2f  :    0 - 0x0
    "11110000", -- 2608 - 0xa30  :  240 - 0xf0 -- Sprite 0xa3
    "11010010", -- 2609 - 0xa31  :  210 - 0xd2
    "10010000", -- 2610 - 0xa32  :  144 - 0x90
    "00010010", -- 2611 - 0xa33  :   18 - 0x12
    "10010000", -- 2612 - 0xa34  :  144 - 0x90
    "11010010", -- 2613 - 0xa35  :  210 - 0xd2
    "11110000", -- 2614 - 0xa36  :  240 - 0xf0
    "11110010", -- 2615 - 0xa37  :  242 - 0xf2
    "00000000", -- 2616 - 0xa38  :    0 - 0x0 -- plane 1
    "00100000", -- 2617 - 0xa39  :   32 - 0x20
    "01100000", -- 2618 - 0xa3a  :   96 - 0x60
    "11100000", -- 2619 - 0xa3b  :  224 - 0xe0
    "01100000", -- 2620 - 0xa3c  :   96 - 0x60
    "00100000", -- 2621 - 0xa3d  :   32 - 0x20
    "00000000", -- 2622 - 0xa3e  :    0 - 0x0
    "00000000", -- 2623 - 0xa3f  :    0 - 0x0
    "11110000", -- 2624 - 0xa40  :  240 - 0xf0 -- Sprite 0xa4
    "11010011", -- 2625 - 0xa41  :  211 - 0xd3
    "10010100", -- 2626 - 0xa42  :  148 - 0x94
    "00011000", -- 2627 - 0xa43  :   24 - 0x18
    "10011111", -- 2628 - 0xa44  :  159 - 0x9f
    "11011101", -- 2629 - 0xa45  :  221 - 0xdd
    "11111010", -- 2630 - 0xa46  :  250 - 0xfa
    "11111101", -- 2631 - 0xa47  :  253 - 0xfd
    "00000000", -- 2632 - 0xa48  :    0 - 0x0 -- plane 1
    "00100000", -- 2633 - 0xa49  :   32 - 0x20
    "01100011", -- 2634 - 0xa4a  :   99 - 0x63
    "11100111", -- 2635 - 0xa4b  :  231 - 0xe7
    "01100000", -- 2636 - 0xa4c  :   96 - 0x60
    "00100010", -- 2637 - 0xa4d  :   34 - 0x22
    "00000101", -- 2638 - 0xa4e  :    5 - 0x5
    "00000010", -- 2639 - 0xa4f  :    2 - 0x2
    "00000000", -- 2640 - 0xa50  :    0 - 0x0 -- Sprite 0xa5
    "11111111", -- 2641 - 0xa51  :  255 - 0xff
    "00000000", -- 2642 - 0xa52  :    0 - 0x0
    "00000000", -- 2643 - 0xa53  :    0 - 0x0
    "11111111", -- 2644 - 0xa54  :  255 - 0xff
    "11011101", -- 2645 - 0xa55  :  221 - 0xdd
    "11111010", -- 2646 - 0xa56  :  250 - 0xfa
    "11111101", -- 2647 - 0xa57  :  253 - 0xfd
    "00000000", -- 2648 - 0xa58  :    0 - 0x0 -- plane 1
    "00000000", -- 2649 - 0xa59  :    0 - 0x0
    "11111111", -- 2650 - 0xa5a  :  255 - 0xff
    "11111111", -- 2651 - 0xa5b  :  255 - 0xff
    "00000000", -- 2652 - 0xa5c  :    0 - 0x0
    "00100010", -- 2653 - 0xa5d  :   34 - 0x22
    "00000101", -- 2654 - 0xa5e  :    5 - 0x5
    "00000010", -- 2655 - 0xa5f  :    2 - 0x2
    "11101111", -- 2656 - 0xa60  :  239 - 0xef -- Sprite 0xa6
    "11000111", -- 2657 - 0xa61  :  199 - 0xc7
    "10000011", -- 2658 - 0xa62  :  131 - 0x83
    "11111111", -- 2659 - 0xa63  :  255 - 0xff
    "00011111", -- 2660 - 0xa64  :   31 - 0x1f
    "00101101", -- 2661 - 0xa65  :   45 - 0x2d
    "01001010", -- 2662 - 0xa66  :   74 - 0x4a
    "01001101", -- 2663 - 0xa67  :   77 - 0x4d
    "00010000", -- 2664 - 0xa68  :   16 - 0x10 -- plane 1
    "00111000", -- 2665 - 0xa69  :   56 - 0x38
    "01111100", -- 2666 - 0xa6a  :  124 - 0x7c
    "00000000", -- 2667 - 0xa6b  :    0 - 0x0
    "00000000", -- 2668 - 0xa6c  :    0 - 0x0
    "00010010", -- 2669 - 0xa6d  :   18 - 0x12
    "00110101", -- 2670 - 0xa6e  :   53 - 0x35
    "00110010", -- 2671 - 0xa6f  :   50 - 0x32
    "01001111", -- 2672 - 0xa70  :   79 - 0x4f -- Sprite 0xa7
    "01001111", -- 2673 - 0xa71  :   79 - 0x4f
    "01001011", -- 2674 - 0xa72  :   75 - 0x4b
    "01001111", -- 2675 - 0xa73  :   79 - 0x4f
    "01001111", -- 2676 - 0xa74  :   79 - 0x4f
    "01001101", -- 2677 - 0xa75  :   77 - 0x4d
    "01001010", -- 2678 - 0xa76  :   74 - 0x4a
    "01001101", -- 2679 - 0xa77  :   77 - 0x4d
    "00110000", -- 2680 - 0xa78  :   48 - 0x30 -- plane 1
    "00110000", -- 2681 - 0xa79  :   48 - 0x30
    "00110100", -- 2682 - 0xa7a  :   52 - 0x34
    "00110000", -- 2683 - 0xa7b  :   48 - 0x30
    "00110000", -- 2684 - 0xa7c  :   48 - 0x30
    "00110010", -- 2685 - 0xa7d  :   50 - 0x32
    "00110101", -- 2686 - 0xa7e  :   53 - 0x35
    "00110010", -- 2687 - 0xa7f  :   50 - 0x32
    "01001111", -- 2688 - 0xa80  :   79 - 0x4f -- Sprite 0xa8
    "11001111", -- 2689 - 0xa81  :  207 - 0xcf
    "00001011", -- 2690 - 0xa82  :   11 - 0xb
    "00001111", -- 2691 - 0xa83  :   15 - 0xf
    "11111111", -- 2692 - 0xa84  :  255 - 0xff
    "11011101", -- 2693 - 0xa85  :  221 - 0xdd
    "11111010", -- 2694 - 0xa86  :  250 - 0xfa
    "11111101", -- 2695 - 0xa87  :  253 - 0xfd
    "00110000", -- 2696 - 0xa88  :   48 - 0x30 -- plane 1
    "00110000", -- 2697 - 0xa89  :   48 - 0x30
    "11110100", -- 2698 - 0xa8a  :  244 - 0xf4
    "11110000", -- 2699 - 0xa8b  :  240 - 0xf0
    "00000000", -- 2700 - 0xa8c  :    0 - 0x0
    "00100010", -- 2701 - 0xa8d  :   34 - 0x22
    "00000101", -- 2702 - 0xa8e  :    5 - 0x5
    "00000010", -- 2703 - 0xa8f  :    2 - 0x2
    "11111111", -- 2704 - 0xa90  :  255 - 0xff -- Sprite 0xa9
    "11111111", -- 2705 - 0xa91  :  255 - 0xff
    "11111111", -- 2706 - 0xa92  :  255 - 0xff
    "11111111", -- 2707 - 0xa93  :  255 - 0xff
    "11111111", -- 2708 - 0xa94  :  255 - 0xff
    "11111111", -- 2709 - 0xa95  :  255 - 0xff
    "11111111", -- 2710 - 0xa96  :  255 - 0xff
    "11111111", -- 2711 - 0xa97  :  255 - 0xff
    "00000000", -- 2712 - 0xa98  :    0 - 0x0 -- plane 1
    "00000000", -- 2713 - 0xa99  :    0 - 0x0
    "00000000", -- 2714 - 0xa9a  :    0 - 0x0
    "00000000", -- 2715 - 0xa9b  :    0 - 0x0
    "00000000", -- 2716 - 0xa9c  :    0 - 0x0
    "00000000", -- 2717 - 0xa9d  :    0 - 0x0
    "00000000", -- 2718 - 0xa9e  :    0 - 0x0
    "00000000", -- 2719 - 0xa9f  :    0 - 0x0
    "11111111", -- 2720 - 0xaa0  :  255 - 0xff -- Sprite 0xaa
    "11111111", -- 2721 - 0xaa1  :  255 - 0xff
    "10101111", -- 2722 - 0xaa2  :  175 - 0xaf
    "01010111", -- 2723 - 0xaa3  :   87 - 0x57
    "10001111", -- 2724 - 0xaa4  :  143 - 0x8f
    "11011101", -- 2725 - 0xaa5  :  221 - 0xdd
    "11111010", -- 2726 - 0xaa6  :  250 - 0xfa
    "11111101", -- 2727 - 0xaa7  :  253 - 0xfd
    "00000000", -- 2728 - 0xaa8  :    0 - 0x0 -- plane 1
    "00000000", -- 2729 - 0xaa9  :    0 - 0x0
    "01010000", -- 2730 - 0xaaa  :   80 - 0x50
    "10101000", -- 2731 - 0xaab  :  168 - 0xa8
    "01110000", -- 2732 - 0xaac  :  112 - 0x70
    "00100010", -- 2733 - 0xaad  :   34 - 0x22
    "00000101", -- 2734 - 0xaae  :    5 - 0x5
    "00000010", -- 2735 - 0xaaf  :    2 - 0x2
    "11111111", -- 2736 - 0xab0  :  255 - 0xff -- Sprite 0xab
    "00000000", -- 2737 - 0xab1  :    0 - 0x0
    "00000000", -- 2738 - 0xab2  :    0 - 0x0
    "00000000", -- 2739 - 0xab3  :    0 - 0x0
    "00000000", -- 2740 - 0xab4  :    0 - 0x0
    "00000000", -- 2741 - 0xab5  :    0 - 0x0
    "00000000", -- 2742 - 0xab6  :    0 - 0x0
    "00000000", -- 2743 - 0xab7  :    0 - 0x0
    "00000000", -- 2744 - 0xab8  :    0 - 0x0 -- plane 1
    "00000000", -- 2745 - 0xab9  :    0 - 0x0
    "00000000", -- 2746 - 0xaba  :    0 - 0x0
    "00000000", -- 2747 - 0xabb  :    0 - 0x0
    "00000000", -- 2748 - 0xabc  :    0 - 0x0
    "00000000", -- 2749 - 0xabd  :    0 - 0x0
    "00000000", -- 2750 - 0xabe  :    0 - 0x0
    "00000000", -- 2751 - 0xabf  :    0 - 0x0
    "00000000", -- 2752 - 0xac0  :    0 - 0x0 -- Sprite 0xac
    "00000000", -- 2753 - 0xac1  :    0 - 0x0
    "00000000", -- 2754 - 0xac2  :    0 - 0x0
    "00000000", -- 2755 - 0xac3  :    0 - 0x0
    "00000000", -- 2756 - 0xac4  :    0 - 0x0
    "00000000", -- 2757 - 0xac5  :    0 - 0x0
    "00000000", -- 2758 - 0xac6  :    0 - 0x0
    "00000000", -- 2759 - 0xac7  :    0 - 0x0
    "00000000", -- 2760 - 0xac8  :    0 - 0x0 -- plane 1
    "00000000", -- 2761 - 0xac9  :    0 - 0x0
    "00000000", -- 2762 - 0xaca  :    0 - 0x0
    "00000000", -- 2763 - 0xacb  :    0 - 0x0
    "00000000", -- 2764 - 0xacc  :    0 - 0x0
    "00000000", -- 2765 - 0xacd  :    0 - 0x0
    "00000000", -- 2766 - 0xace  :    0 - 0x0
    "00000000", -- 2767 - 0xacf  :    0 - 0x0
    "00000000", -- 2768 - 0xad0  :    0 - 0x0 -- Sprite 0xad
    "11111111", -- 2769 - 0xad1  :  255 - 0xff
    "00000000", -- 2770 - 0xad2  :    0 - 0x0
    "11111111", -- 2771 - 0xad3  :  255 - 0xff
    "11111111", -- 2772 - 0xad4  :  255 - 0xff
    "11111111", -- 2773 - 0xad5  :  255 - 0xff
    "11111111", -- 2774 - 0xad6  :  255 - 0xff
    "11111111", -- 2775 - 0xad7  :  255 - 0xff
    "00000000", -- 2776 - 0xad8  :    0 - 0x0 -- plane 1
    "00000000", -- 2777 - 0xad9  :    0 - 0x0
    "11111111", -- 2778 - 0xada  :  255 - 0xff
    "00000000", -- 2779 - 0xadb  :    0 - 0x0
    "00000000", -- 2780 - 0xadc  :    0 - 0x0
    "00000000", -- 2781 - 0xadd  :    0 - 0x0
    "00000000", -- 2782 - 0xade  :    0 - 0x0
    "00000000", -- 2783 - 0xadf  :    0 - 0x0
    "11111111", -- 2784 - 0xae0  :  255 - 0xff -- Sprite 0xae
    "11111111", -- 2785 - 0xae1  :  255 - 0xff
    "11111111", -- 2786 - 0xae2  :  255 - 0xff
    "11111111", -- 2787 - 0xae3  :  255 - 0xff
    "11111111", -- 2788 - 0xae4  :  255 - 0xff
    "00000000", -- 2789 - 0xae5  :    0 - 0x0
    "11111111", -- 2790 - 0xae6  :  255 - 0xff
    "00000000", -- 2791 - 0xae7  :    0 - 0x0
    "00000000", -- 2792 - 0xae8  :    0 - 0x0 -- plane 1
    "00000000", -- 2793 - 0xae9  :    0 - 0x0
    "00000000", -- 2794 - 0xaea  :    0 - 0x0
    "00000000", -- 2795 - 0xaeb  :    0 - 0x0
    "00000000", -- 2796 - 0xaec  :    0 - 0x0
    "11111111", -- 2797 - 0xaed  :  255 - 0xff
    "00000000", -- 2798 - 0xaee  :    0 - 0x0
    "00000000", -- 2799 - 0xaef  :    0 - 0x0
    "11111111", -- 2800 - 0xaf0  :  255 - 0xff -- Sprite 0xaf
    "11111111", -- 2801 - 0xaf1  :  255 - 0xff
    "11111111", -- 2802 - 0xaf2  :  255 - 0xff
    "11111111", -- 2803 - 0xaf3  :  255 - 0xff
    "11111111", -- 2804 - 0xaf4  :  255 - 0xff
    "11111111", -- 2805 - 0xaf5  :  255 - 0xff
    "11111111", -- 2806 - 0xaf6  :  255 - 0xff
    "11111111", -- 2807 - 0xaf7  :  255 - 0xff
    "00000000", -- 2808 - 0xaf8  :    0 - 0x0 -- plane 1
    "00000000", -- 2809 - 0xaf9  :    0 - 0x0
    "00000000", -- 2810 - 0xafa  :    0 - 0x0
    "00000000", -- 2811 - 0xafb  :    0 - 0x0
    "00000000", -- 2812 - 0xafc  :    0 - 0x0
    "00000000", -- 2813 - 0xafd  :    0 - 0x0
    "00000000", -- 2814 - 0xafe  :    0 - 0x0
    "00000000", -- 2815 - 0xaff  :    0 - 0x0
    "00000000", -- 2816 - 0xb00  :    0 - 0x0 -- Sprite 0xb0
    "00011111", -- 2817 - 0xb01  :   31 - 0x1f
    "00010000", -- 2818 - 0xb02  :   16 - 0x10
    "00010000", -- 2819 - 0xb03  :   16 - 0x10
    "00010000", -- 2820 - 0xb04  :   16 - 0x10
    "00010000", -- 2821 - 0xb05  :   16 - 0x10
    "00010000", -- 2822 - 0xb06  :   16 - 0x10
    "00010000", -- 2823 - 0xb07  :   16 - 0x10
    "00000000", -- 2824 - 0xb08  :    0 - 0x0 -- plane 1
    "00011111", -- 2825 - 0xb09  :   31 - 0x1f
    "00011111", -- 2826 - 0xb0a  :   31 - 0x1f
    "00011111", -- 2827 - 0xb0b  :   31 - 0x1f
    "00011111", -- 2828 - 0xb0c  :   31 - 0x1f
    "00011111", -- 2829 - 0xb0d  :   31 - 0x1f
    "00011111", -- 2830 - 0xb0e  :   31 - 0x1f
    "00011111", -- 2831 - 0xb0f  :   31 - 0x1f
    "00000000", -- 2832 - 0xb10  :    0 - 0x0 -- Sprite 0xb1
    "11111000", -- 2833 - 0xb11  :  248 - 0xf8
    "00001000", -- 2834 - 0xb12  :    8 - 0x8
    "00001000", -- 2835 - 0xb13  :    8 - 0x8
    "00001000", -- 2836 - 0xb14  :    8 - 0x8
    "00001000", -- 2837 - 0xb15  :    8 - 0x8
    "00001000", -- 2838 - 0xb16  :    8 - 0x8
    "00001000", -- 2839 - 0xb17  :    8 - 0x8
    "00000000", -- 2840 - 0xb18  :    0 - 0x0 -- plane 1
    "11110000", -- 2841 - 0xb19  :  240 - 0xf0
    "11110000", -- 2842 - 0xb1a  :  240 - 0xf0
    "11110000", -- 2843 - 0xb1b  :  240 - 0xf0
    "11110000", -- 2844 - 0xb1c  :  240 - 0xf0
    "11110000", -- 2845 - 0xb1d  :  240 - 0xf0
    "11110000", -- 2846 - 0xb1e  :  240 - 0xf0
    "11110000", -- 2847 - 0xb1f  :  240 - 0xf0
    "00010000", -- 2848 - 0xb20  :   16 - 0x10 -- Sprite 0xb2
    "00010000", -- 2849 - 0xb21  :   16 - 0x10
    "00010000", -- 2850 - 0xb22  :   16 - 0x10
    "00010000", -- 2851 - 0xb23  :   16 - 0x10
    "00011111", -- 2852 - 0xb24  :   31 - 0x1f
    "00011111", -- 2853 - 0xb25  :   31 - 0x1f
    "00001111", -- 2854 - 0xb26  :   15 - 0xf
    "00000000", -- 2855 - 0xb27  :    0 - 0x0
    "00011111", -- 2856 - 0xb28  :   31 - 0x1f -- plane 1
    "00011111", -- 2857 - 0xb29  :   31 - 0x1f
    "00011111", -- 2858 - 0xb2a  :   31 - 0x1f
    "00011111", -- 2859 - 0xb2b  :   31 - 0x1f
    "00000000", -- 2860 - 0xb2c  :    0 - 0x0
    "00000000", -- 2861 - 0xb2d  :    0 - 0x0
    "00000000", -- 2862 - 0xb2e  :    0 - 0x0
    "00000000", -- 2863 - 0xb2f  :    0 - 0x0
    "00001000", -- 2864 - 0xb30  :    8 - 0x8 -- Sprite 0xb3
    "00001000", -- 2865 - 0xb31  :    8 - 0x8
    "00001000", -- 2866 - 0xb32  :    8 - 0x8
    "00001000", -- 2867 - 0xb33  :    8 - 0x8
    "11111000", -- 2868 - 0xb34  :  248 - 0xf8
    "11111000", -- 2869 - 0xb35  :  248 - 0xf8
    "11110000", -- 2870 - 0xb36  :  240 - 0xf0
    "00000000", -- 2871 - 0xb37  :    0 - 0x0
    "11110000", -- 2872 - 0xb38  :  240 - 0xf0 -- plane 1
    "11110000", -- 2873 - 0xb39  :  240 - 0xf0
    "11110000", -- 2874 - 0xb3a  :  240 - 0xf0
    "11110000", -- 2875 - 0xb3b  :  240 - 0xf0
    "00000000", -- 2876 - 0xb3c  :    0 - 0x0
    "00000000", -- 2877 - 0xb3d  :    0 - 0x0
    "00000000", -- 2878 - 0xb3e  :    0 - 0x0
    "00000000", -- 2879 - 0xb3f  :    0 - 0x0
    "00000000", -- 2880 - 0xb40  :    0 - 0x0 -- Sprite 0xb4
    "00000000", -- 2881 - 0xb41  :    0 - 0x0
    "00111111", -- 2882 - 0xb42  :   63 - 0x3f
    "01100000", -- 2883 - 0xb43  :   96 - 0x60
    "01100000", -- 2884 - 0xb44  :   96 - 0x60
    "01100000", -- 2885 - 0xb45  :   96 - 0x60
    "01100000", -- 2886 - 0xb46  :   96 - 0x60
    "01100000", -- 2887 - 0xb47  :   96 - 0x60
    "00000000", -- 2888 - 0xb48  :    0 - 0x0 -- plane 1
    "00000000", -- 2889 - 0xb49  :    0 - 0x0
    "00111111", -- 2890 - 0xb4a  :   63 - 0x3f
    "01111111", -- 2891 - 0xb4b  :  127 - 0x7f
    "01111111", -- 2892 - 0xb4c  :  127 - 0x7f
    "01111111", -- 2893 - 0xb4d  :  127 - 0x7f
    "01111111", -- 2894 - 0xb4e  :  127 - 0x7f
    "01111111", -- 2895 - 0xb4f  :  127 - 0x7f
    "00000000", -- 2896 - 0xb50  :    0 - 0x0 -- Sprite 0xb5
    "00000000", -- 2897 - 0xb51  :    0 - 0x0
    "11111100", -- 2898 - 0xb52  :  252 - 0xfc
    "00000110", -- 2899 - 0xb53  :    6 - 0x6
    "00000110", -- 2900 - 0xb54  :    6 - 0x6
    "00000110", -- 2901 - 0xb55  :    6 - 0x6
    "00000110", -- 2902 - 0xb56  :    6 - 0x6
    "00000110", -- 2903 - 0xb57  :    6 - 0x6
    "00000000", -- 2904 - 0xb58  :    0 - 0x0 -- plane 1
    "00000000", -- 2905 - 0xb59  :    0 - 0x0
    "11111000", -- 2906 - 0xb5a  :  248 - 0xf8
    "11111000", -- 2907 - 0xb5b  :  248 - 0xf8
    "11111000", -- 2908 - 0xb5c  :  248 - 0xf8
    "11111000", -- 2909 - 0xb5d  :  248 - 0xf8
    "11111000", -- 2910 - 0xb5e  :  248 - 0xf8
    "11111000", -- 2911 - 0xb5f  :  248 - 0xf8
    "01100000", -- 2912 - 0xb60  :   96 - 0x60 -- Sprite 0xb6
    "01100000", -- 2913 - 0xb61  :   96 - 0x60
    "01100000", -- 2914 - 0xb62  :   96 - 0x60
    "01111111", -- 2915 - 0xb63  :  127 - 0x7f
    "01111111", -- 2916 - 0xb64  :  127 - 0x7f
    "00111111", -- 2917 - 0xb65  :   63 - 0x3f
    "00000000", -- 2918 - 0xb66  :    0 - 0x0
    "00000000", -- 2919 - 0xb67  :    0 - 0x0
    "01111111", -- 2920 - 0xb68  :  127 - 0x7f -- plane 1
    "01111111", -- 2921 - 0xb69  :  127 - 0x7f
    "01111111", -- 2922 - 0xb6a  :  127 - 0x7f
    "01000000", -- 2923 - 0xb6b  :   64 - 0x40
    "00000000", -- 2924 - 0xb6c  :    0 - 0x0
    "00000000", -- 2925 - 0xb6d  :    0 - 0x0
    "00000000", -- 2926 - 0xb6e  :    0 - 0x0
    "00000000", -- 2927 - 0xb6f  :    0 - 0x0
    "00000110", -- 2928 - 0xb70  :    6 - 0x6 -- Sprite 0xb7
    "00000110", -- 2929 - 0xb71  :    6 - 0x6
    "00000110", -- 2930 - 0xb72  :    6 - 0x6
    "11111110", -- 2931 - 0xb73  :  254 - 0xfe
    "11111110", -- 2932 - 0xb74  :  254 - 0xfe
    "11111100", -- 2933 - 0xb75  :  252 - 0xfc
    "00000000", -- 2934 - 0xb76  :    0 - 0x0
    "00000000", -- 2935 - 0xb77  :    0 - 0x0
    "11111000", -- 2936 - 0xb78  :  248 - 0xf8 -- plane 1
    "11111000", -- 2937 - 0xb79  :  248 - 0xf8
    "11111000", -- 2938 - 0xb7a  :  248 - 0xf8
    "00000000", -- 2939 - 0xb7b  :    0 - 0x0
    "00000000", -- 2940 - 0xb7c  :    0 - 0x0
    "00000000", -- 2941 - 0xb7d  :    0 - 0x0
    "00000000", -- 2942 - 0xb7e  :    0 - 0x0
    "00000000", -- 2943 - 0xb7f  :    0 - 0x0
    "01100000", -- 2944 - 0xb80  :   96 - 0x60 -- Sprite 0xb8
    "11110011", -- 2945 - 0xb81  :  243 - 0xf3
    "11000111", -- 2946 - 0xb82  :  199 - 0xc7
    "10000110", -- 2947 - 0xb83  :  134 - 0x86
    "00000100", -- 2948 - 0xb84  :    4 - 0x4
    "00000100", -- 2949 - 0xb85  :    4 - 0x4
    "00000111", -- 2950 - 0xb86  :    7 - 0x7
    "00000111", -- 2951 - 0xb87  :    7 - 0x7
    "00000000", -- 2952 - 0xb88  :    0 - 0x0 -- plane 1
    "00000011", -- 2953 - 0xb89  :    3 - 0x3
    "00000111", -- 2954 - 0xb8a  :    7 - 0x7
    "00000111", -- 2955 - 0xb8b  :    7 - 0x7
    "00000111", -- 2956 - 0xb8c  :    7 - 0x7
    "00000011", -- 2957 - 0xb8d  :    3 - 0x3
    "00000000", -- 2958 - 0xb8e  :    0 - 0x0
    "00000000", -- 2959 - 0xb8f  :    0 - 0x0
    "00000110", -- 2960 - 0xb90  :    6 - 0x6 -- Sprite 0xb9
    "10001111", -- 2961 - 0xb91  :  143 - 0x8f
    "11000101", -- 2962 - 0xb92  :  197 - 0xc5
    "00100011", -- 2963 - 0xb93  :   35 - 0x23
    "00101110", -- 2964 - 0xb94  :   46 - 0x2e
    "01100000", -- 2965 - 0xb95  :   96 - 0x60
    "11100001", -- 2966 - 0xb96  :  225 - 0xe1
    "11100001", -- 2967 - 0xb97  :  225 - 0xe1
    "00000000", -- 2968 - 0xb98  :    0 - 0x0 -- plane 1
    "11000001", -- 2969 - 0xb99  :  193 - 0xc1
    "11100010", -- 2970 - 0xb9a  :  226 - 0xe2
    "11001100", -- 2971 - 0xb9b  :  204 - 0xcc
    "11000000", -- 2972 - 0xb9c  :  192 - 0xc0
    "10000000", -- 2973 - 0xb9d  :  128 - 0x80
    "00000001", -- 2974 - 0xb9e  :    1 - 0x1
    "00000010", -- 2975 - 0xb9f  :    2 - 0x2
    "11001000", -- 2976 - 0xba0  :  200 - 0xc8 -- Sprite 0xba
    "11111000", -- 2977 - 0xba1  :  248 - 0xf8
    "10110000", -- 2978 - 0xba2  :  176 - 0xb0
    "00010000", -- 2979 - 0xba3  :   16 - 0x10
    "00110000", -- 2980 - 0xba4  :   48 - 0x30
    "11001000", -- 2981 - 0xba5  :  200 - 0xc8
    "11111000", -- 2982 - 0xba6  :  248 - 0xf8
    "10000000", -- 2983 - 0xba7  :  128 - 0x80
    "11110000", -- 2984 - 0xba8  :  240 - 0xf0 -- plane 1
    "00000000", -- 2985 - 0xba9  :    0 - 0x0
    "00100000", -- 2986 - 0xbaa  :   32 - 0x20
    "00100000", -- 2987 - 0xbab  :   32 - 0x20
    "00000000", -- 2988 - 0xbac  :    0 - 0x0
    "11110000", -- 2989 - 0xbad  :  240 - 0xf0
    "00000000", -- 2990 - 0xbae  :    0 - 0x0
    "00000000", -- 2991 - 0xbaf  :    0 - 0x0
    "00000011", -- 2992 - 0xbb0  :    3 - 0x3 -- Sprite 0xbb
    "00000000", -- 2993 - 0xbb1  :    0 - 0x0
    "00000000", -- 2994 - 0xbb2  :    0 - 0x0
    "01100000", -- 2995 - 0xbb3  :   96 - 0x60
    "11110000", -- 2996 - 0xbb4  :  240 - 0xf0
    "11010000", -- 2997 - 0xbb5  :  208 - 0xd0
    "10010000", -- 2998 - 0xbb6  :  144 - 0x90
    "01100000", -- 2999 - 0xbb7  :   96 - 0x60
    "00000000", -- 3000 - 0xbb8  :    0 - 0x0 -- plane 1
    "00000000", -- 3001 - 0xbb9  :    0 - 0x0
    "00000000", -- 3002 - 0xbba  :    0 - 0x0
    "00000000", -- 3003 - 0xbbb  :    0 - 0x0
    "00000000", -- 3004 - 0xbbc  :    0 - 0x0
    "01100000", -- 3005 - 0xbbd  :   96 - 0x60
    "01100000", -- 3006 - 0xbbe  :   96 - 0x60
    "00000000", -- 3007 - 0xbbf  :    0 - 0x0
    "11000011", -- 3008 - 0xbc0  :  195 - 0xc3 -- Sprite 0xbc
    "00001110", -- 3009 - 0xbc1  :   14 - 0xe
    "00000000", -- 3010 - 0xbc2  :    0 - 0x0
    "00000110", -- 3011 - 0xbc3  :    6 - 0x6
    "00001111", -- 3012 - 0xbc4  :   15 - 0xf
    "00001101", -- 3013 - 0xbc5  :   13 - 0xd
    "00001001", -- 3014 - 0xbc6  :    9 - 0x9
    "00000110", -- 3015 - 0xbc7  :    6 - 0x6
    "00001100", -- 3016 - 0xbc8  :   12 - 0xc -- plane 1
    "00000000", -- 3017 - 0xbc9  :    0 - 0x0
    "00000000", -- 3018 - 0xbca  :    0 - 0x0
    "00000000", -- 3019 - 0xbcb  :    0 - 0x0
    "00000000", -- 3020 - 0xbcc  :    0 - 0x0
    "00000110", -- 3021 - 0xbcd  :    6 - 0x6
    "00000110", -- 3022 - 0xbce  :    6 - 0x6
    "00000000", -- 3023 - 0xbcf  :    0 - 0x0
    "11100000", -- 3024 - 0xbd0  :  224 - 0xe0 -- Sprite 0xbd
    "01100011", -- 3025 - 0xbd1  :   99 - 0x63
    "11100111", -- 3026 - 0xbd2  :  231 - 0xe7
    "11100110", -- 3027 - 0xbd3  :  230 - 0xe6
    "00000100", -- 3028 - 0xbd4  :    4 - 0x4
    "00000100", -- 3029 - 0xbd5  :    4 - 0x4
    "00000111", -- 3030 - 0xbd6  :    7 - 0x7
    "00000111", -- 3031 - 0xbd7  :    7 - 0x7
    "00000000", -- 3032 - 0xbd8  :    0 - 0x0 -- plane 1
    "10000011", -- 3033 - 0xbd9  :  131 - 0x83
    "00000111", -- 3034 - 0xbda  :    7 - 0x7
    "00000111", -- 3035 - 0xbdb  :    7 - 0x7
    "00000111", -- 3036 - 0xbdc  :    7 - 0x7
    "00000011", -- 3037 - 0xbdd  :    3 - 0x3
    "00000000", -- 3038 - 0xbde  :    0 - 0x0
    "00000000", -- 3039 - 0xbdf  :    0 - 0x0
    "00000111", -- 3040 - 0xbe0  :    7 - 0x7 -- Sprite 0xbe
    "10000011", -- 3041 - 0xbe1  :  131 - 0x83
    "11000111", -- 3042 - 0xbe2  :  199 - 0xc7
    "00100111", -- 3043 - 0xbe3  :   39 - 0x27
    "00100000", -- 3044 - 0xbe4  :   32 - 0x20
    "01100000", -- 3045 - 0xbe5  :   96 - 0x60
    "11100000", -- 3046 - 0xbe6  :  224 - 0xe0
    "11100000", -- 3047 - 0xbe7  :  224 - 0xe0
    "00000000", -- 3048 - 0xbe8  :    0 - 0x0 -- plane 1
    "11000100", -- 3049 - 0xbe9  :  196 - 0xc4
    "11100000", -- 3050 - 0xbea  :  224 - 0xe0
    "11000000", -- 3051 - 0xbeb  :  192 - 0xc0
    "11000000", -- 3052 - 0xbec  :  192 - 0xc0
    "10000000", -- 3053 - 0xbed  :  128 - 0x80
    "00000000", -- 3054 - 0xbee  :    0 - 0x0
    "00000000", -- 3055 - 0xbef  :    0 - 0x0
    "00000011", -- 3056 - 0xbf0  :    3 - 0x3 -- Sprite 0xbf
    "00000000", -- 3057 - 0xbf1  :    0 - 0x0
    "00001100", -- 3058 - 0xbf2  :   12 - 0xc
    "00001100", -- 3059 - 0xbf3  :   12 - 0xc
    "11100100", -- 3060 - 0xbf4  :  228 - 0xe4
    "01101100", -- 3061 - 0xbf5  :  108 - 0x6c
    "11101101", -- 3062 - 0xbf6  :  237 - 0xed
    "11100111", -- 3063 - 0xbf7  :  231 - 0xe7
    "00000000", -- 3064 - 0xbf8  :    0 - 0x0 -- plane 1
    "00000000", -- 3065 - 0xbf9  :    0 - 0x0
    "00000000", -- 3066 - 0xbfa  :    0 - 0x0
    "00000000", -- 3067 - 0xbfb  :    0 - 0x0
    "00001000", -- 3068 - 0xbfc  :    8 - 0x8
    "10001000", -- 3069 - 0xbfd  :  136 - 0x88
    "00001011", -- 3070 - 0xbfe  :   11 - 0xb
    "00001000", -- 3071 - 0xbff  :    8 - 0x8
    "11000000", -- 3072 - 0xc00  :  192 - 0xc0 -- Sprite 0xc0
    "00000000", -- 3073 - 0xc01  :    0 - 0x0
    "00110000", -- 3074 - 0xc02  :   48 - 0x30
    "00110000", -- 3075 - 0xc03  :   48 - 0x30
    "00010111", -- 3076 - 0xc04  :   23 - 0x17
    "00110011", -- 3077 - 0xc05  :   51 - 0x33
    "01110111", -- 3078 - 0xc06  :  119 - 0x77
    "11010111", -- 3079 - 0xc07  :  215 - 0xd7
    "00000000", -- 3080 - 0xc08  :    0 - 0x0 -- plane 1
    "00000000", -- 3081 - 0xc09  :    0 - 0x0
    "00000000", -- 3082 - 0xc0a  :    0 - 0x0
    "00000000", -- 3083 - 0xc0b  :    0 - 0x0
    "00100000", -- 3084 - 0xc0c  :   32 - 0x20
    "00100100", -- 3085 - 0xc0d  :   36 - 0x24
    "10100000", -- 3086 - 0xc0e  :  160 - 0xa0
    "00100000", -- 3087 - 0xc0f  :   32 - 0x20
    "00001100", -- 3088 - 0xc10  :   12 - 0xc -- Sprite 0xc1
    "00000000", -- 3089 - 0xc11  :    0 - 0x0
    "00000000", -- 3090 - 0xc12  :    0 - 0x0
    "00000000", -- 3091 - 0xc13  :    0 - 0x0
    "00000000", -- 3092 - 0xc14  :    0 - 0x0
    "00000000", -- 3093 - 0xc15  :    0 - 0x0
    "00000000", -- 3094 - 0xc16  :    0 - 0x0
    "00000000", -- 3095 - 0xc17  :    0 - 0x0
    "00000000", -- 3096 - 0xc18  :    0 - 0x0 -- plane 1
    "00000000", -- 3097 - 0xc19  :    0 - 0x0
    "00000000", -- 3098 - 0xc1a  :    0 - 0x0
    "00000000", -- 3099 - 0xc1b  :    0 - 0x0
    "00000000", -- 3100 - 0xc1c  :    0 - 0x0
    "00000000", -- 3101 - 0xc1d  :    0 - 0x0
    "00000000", -- 3102 - 0xc1e  :    0 - 0x0
    "00000000", -- 3103 - 0xc1f  :    0 - 0x0
    "00110000", -- 3104 - 0xc20  :   48 - 0x30 -- Sprite 0xc2
    "00000000", -- 3105 - 0xc21  :    0 - 0x0
    "00000000", -- 3106 - 0xc22  :    0 - 0x0
    "00000000", -- 3107 - 0xc23  :    0 - 0x0
    "00000000", -- 3108 - 0xc24  :    0 - 0x0
    "00000000", -- 3109 - 0xc25  :    0 - 0x0
    "00000000", -- 3110 - 0xc26  :    0 - 0x0
    "00000000", -- 3111 - 0xc27  :    0 - 0x0
    "00000000", -- 3112 - 0xc28  :    0 - 0x0 -- plane 1
    "00000000", -- 3113 - 0xc29  :    0 - 0x0
    "00000000", -- 3114 - 0xc2a  :    0 - 0x0
    "00000000", -- 3115 - 0xc2b  :    0 - 0x0
    "00000000", -- 3116 - 0xc2c  :    0 - 0x0
    "00000000", -- 3117 - 0xc2d  :    0 - 0x0
    "00000000", -- 3118 - 0xc2e  :    0 - 0x0
    "00000000", -- 3119 - 0xc2f  :    0 - 0x0
    "00000000", -- 3120 - 0xc30  :    0 - 0x0 -- Sprite 0xc3
    "00000000", -- 3121 - 0xc31  :    0 - 0x0
    "00000100", -- 3122 - 0xc32  :    4 - 0x4
    "00001101", -- 3123 - 0xc33  :   13 - 0xd
    "00001111", -- 3124 - 0xc34  :   15 - 0xf
    "00001100", -- 3125 - 0xc35  :   12 - 0xc
    "00001100", -- 3126 - 0xc36  :   12 - 0xc
    "00000100", -- 3127 - 0xc37  :    4 - 0x4
    "00000000", -- 3128 - 0xc38  :    0 - 0x0 -- plane 1
    "00000000", -- 3129 - 0xc39  :    0 - 0x0
    "00001000", -- 3130 - 0xc3a  :    8 - 0x8
    "00001011", -- 3131 - 0xc3b  :   11 - 0xb
    "00001000", -- 3132 - 0xc3c  :    8 - 0x8
    "00001000", -- 3133 - 0xc3d  :    8 - 0x8
    "00001000", -- 3134 - 0xc3e  :    8 - 0x8
    "00001000", -- 3135 - 0xc3f  :    8 - 0x8
    "00000000", -- 3136 - 0xc40  :    0 - 0x0 -- Sprite 0xc4
    "00000000", -- 3137 - 0xc41  :    0 - 0x0
    "00010000", -- 3138 - 0xc42  :   16 - 0x10
    "01110000", -- 3139 - 0xc43  :  112 - 0x70
    "11110000", -- 3140 - 0xc44  :  240 - 0xf0
    "00110000", -- 3141 - 0xc45  :   48 - 0x30
    "00110000", -- 3142 - 0xc46  :   48 - 0x30
    "00010000", -- 3143 - 0xc47  :   16 - 0x10
    "00000000", -- 3144 - 0xc48  :    0 - 0x0 -- plane 1
    "00000000", -- 3145 - 0xc49  :    0 - 0x0
    "00100000", -- 3146 - 0xc4a  :   32 - 0x20
    "10100000", -- 3147 - 0xc4b  :  160 - 0xa0
    "00100000", -- 3148 - 0xc4c  :   32 - 0x20
    "00100000", -- 3149 - 0xc4d  :   32 - 0x20
    "00100000", -- 3150 - 0xc4e  :   32 - 0x20
    "00100000", -- 3151 - 0xc4f  :   32 - 0x20
    "11100100", -- 3152 - 0xc50  :  228 - 0xe4 -- Sprite 0xc5
    "00100100", -- 3153 - 0xc51  :   36 - 0x24
    "11101111", -- 3154 - 0xc52  :  239 - 0xef
    "11100111", -- 3155 - 0xc53  :  231 - 0xe7
    "00000110", -- 3156 - 0xc54  :    6 - 0x6
    "00000100", -- 3157 - 0xc55  :    4 - 0x4
    "00000100", -- 3158 - 0xc56  :    4 - 0x4
    "00000111", -- 3159 - 0xc57  :    7 - 0x7
    "00001000", -- 3160 - 0xc58  :    8 - 0x8 -- plane 1
    "11001000", -- 3161 - 0xc59  :  200 - 0xc8
    "00000011", -- 3162 - 0xc5a  :    3 - 0x3
    "00000111", -- 3163 - 0xc5b  :    7 - 0x7
    "00000111", -- 3164 - 0xc5c  :    7 - 0x7
    "00000111", -- 3165 - 0xc5d  :    7 - 0x7
    "00000011", -- 3166 - 0xc5e  :    3 - 0x3
    "00000000", -- 3167 - 0xc5f  :    0 - 0x0
    "00010111", -- 3168 - 0xc60  :   23 - 0x17 -- Sprite 0xc6
    "00010001", -- 3169 - 0xc61  :   17 - 0x11
    "10110111", -- 3170 - 0xc62  :  183 - 0xb7
    "11000111", -- 3171 - 0xc63  :  199 - 0xc7
    "00100000", -- 3172 - 0xc64  :   32 - 0x20
    "00100000", -- 3173 - 0xc65  :   32 - 0x20
    "01100000", -- 3174 - 0xc66  :   96 - 0x60
    "11100000", -- 3175 - 0xc67  :  224 - 0xe0
    "00100000", -- 3176 - 0xc68  :   32 - 0x20 -- plane 1
    "00100110", -- 3177 - 0xc69  :   38 - 0x26
    "11000000", -- 3178 - 0xc6a  :  192 - 0xc0
    "11100000", -- 3179 - 0xc6b  :  224 - 0xe0
    "11000000", -- 3180 - 0xc6c  :  192 - 0xc0
    "11000000", -- 3181 - 0xc6d  :  192 - 0xc0
    "10000000", -- 3182 - 0xc6e  :  128 - 0x80
    "00000000", -- 3183 - 0xc6f  :    0 - 0x0
    "00000111", -- 3184 - 0xc70  :    7 - 0x7 -- Sprite 0xc7
    "00000011", -- 3185 - 0xc71  :    3 - 0x3
    "00000000", -- 3186 - 0xc72  :    0 - 0x0
    "00000000", -- 3187 - 0xc73  :    0 - 0x0
    "11100000", -- 3188 - 0xc74  :  224 - 0xe0
    "00100000", -- 3189 - 0xc75  :   32 - 0x20
    "11100000", -- 3190 - 0xc76  :  224 - 0xe0
    "11100000", -- 3191 - 0xc77  :  224 - 0xe0
    "00000000", -- 3192 - 0xc78  :    0 - 0x0 -- plane 1
    "00000000", -- 3193 - 0xc79  :    0 - 0x0
    "00000000", -- 3194 - 0xc7a  :    0 - 0x0
    "00000000", -- 3195 - 0xc7b  :    0 - 0x0
    "00000000", -- 3196 - 0xc7c  :    0 - 0x0
    "11000000", -- 3197 - 0xc7d  :  192 - 0xc0
    "00000000", -- 3198 - 0xc7e  :    0 - 0x0
    "00000000", -- 3199 - 0xc7f  :    0 - 0x0
    "11100000", -- 3200 - 0xc80  :  224 - 0xe0 -- Sprite 0xc8
    "11000000", -- 3201 - 0xc81  :  192 - 0xc0
    "00000000", -- 3202 - 0xc82  :    0 - 0x0
    "00000000", -- 3203 - 0xc83  :    0 - 0x0
    "00000111", -- 3204 - 0xc84  :    7 - 0x7
    "00000001", -- 3205 - 0xc85  :    1 - 0x1
    "00000111", -- 3206 - 0xc86  :    7 - 0x7
    "00000111", -- 3207 - 0xc87  :    7 - 0x7
    "00000000", -- 3208 - 0xc88  :    0 - 0x0 -- plane 1
    "00000000", -- 3209 - 0xc89  :    0 - 0x0
    "00000000", -- 3210 - 0xc8a  :    0 - 0x0
    "00000000", -- 3211 - 0xc8b  :    0 - 0x0
    "00000000", -- 3212 - 0xc8c  :    0 - 0x0
    "00000110", -- 3213 - 0xc8d  :    6 - 0x6
    "00000000", -- 3214 - 0xc8e  :    0 - 0x0
    "00000000", -- 3215 - 0xc8f  :    0 - 0x0
    "00010011", -- 3216 - 0xc90  :   19 - 0x13 -- Sprite 0xc9
    "00011111", -- 3217 - 0xc91  :   31 - 0x1f
    "00001101", -- 3218 - 0xc92  :   13 - 0xd
    "00000100", -- 3219 - 0xc93  :    4 - 0x4
    "00001100", -- 3220 - 0xc94  :   12 - 0xc
    "00010011", -- 3221 - 0xc95  :   19 - 0x13
    "00011111", -- 3222 - 0xc96  :   31 - 0x1f
    "00000001", -- 3223 - 0xc97  :    1 - 0x1
    "00001111", -- 3224 - 0xc98  :   15 - 0xf -- plane 1
    "00000000", -- 3225 - 0xc99  :    0 - 0x0
    "00001000", -- 3226 - 0xc9a  :    8 - 0x8
    "00001000", -- 3227 - 0xc9b  :    8 - 0x8
    "00000000", -- 3228 - 0xc9c  :    0 - 0x0
    "00001111", -- 3229 - 0xc9d  :   15 - 0xf
    "00000000", -- 3230 - 0xc9e  :    0 - 0x0
    "00000000", -- 3231 - 0xc9f  :    0 - 0x0
    "01100000", -- 3232 - 0xca0  :   96 - 0x60 -- Sprite 0xca
    "11110011", -- 3233 - 0xca1  :  243 - 0xf3
    "10100111", -- 3234 - 0xca2  :  167 - 0xa7
    "11000110", -- 3235 - 0xca3  :  198 - 0xc6
    "01110100", -- 3236 - 0xca4  :  116 - 0x74
    "00000100", -- 3237 - 0xca5  :    4 - 0x4
    "10000111", -- 3238 - 0xca6  :  135 - 0x87
    "10000111", -- 3239 - 0xca7  :  135 - 0x87
    "00000000", -- 3240 - 0xca8  :    0 - 0x0 -- plane 1
    "10000011", -- 3241 - 0xca9  :  131 - 0x83
    "01000111", -- 3242 - 0xcaa  :   71 - 0x47
    "00110111", -- 3243 - 0xcab  :   55 - 0x37
    "00000111", -- 3244 - 0xcac  :    7 - 0x7
    "00000011", -- 3245 - 0xcad  :    3 - 0x3
    "10000000", -- 3246 - 0xcae  :  128 - 0x80
    "01000000", -- 3247 - 0xcaf  :   64 - 0x40
    "00000110", -- 3248 - 0xcb0  :    6 - 0x6 -- Sprite 0xcb
    "10001111", -- 3249 - 0xcb1  :  143 - 0x8f
    "11000011", -- 3250 - 0xcb2  :  195 - 0xc3
    "00100001", -- 3251 - 0xcb3  :   33 - 0x21
    "00100000", -- 3252 - 0xcb4  :   32 - 0x20
    "01100000", -- 3253 - 0xcb5  :   96 - 0x60
    "11100000", -- 3254 - 0xcb6  :  224 - 0xe0
    "11100000", -- 3255 - 0xcb7  :  224 - 0xe0
    "00000000", -- 3256 - 0xcb8  :    0 - 0x0 -- plane 1
    "11000000", -- 3257 - 0xcb9  :  192 - 0xc0
    "11100000", -- 3258 - 0xcba  :  224 - 0xe0
    "11000000", -- 3259 - 0xcbb  :  192 - 0xc0
    "11000000", -- 3260 - 0xcbc  :  192 - 0xc0
    "10000000", -- 3261 - 0xcbd  :  128 - 0x80
    "00000000", -- 3262 - 0xcbe  :    0 - 0x0
    "00000000", -- 3263 - 0xcbf  :    0 - 0x0
    "11000011", -- 3264 - 0xcc0  :  195 - 0xc3 -- Sprite 0xcc
    "01110000", -- 3265 - 0xcc1  :  112 - 0x70
    "00000000", -- 3266 - 0xcc2  :    0 - 0x0
    "01100000", -- 3267 - 0xcc3  :   96 - 0x60
    "11110000", -- 3268 - 0xcc4  :  240 - 0xf0
    "11010000", -- 3269 - 0xcc5  :  208 - 0xd0
    "10010000", -- 3270 - 0xcc6  :  144 - 0x90
    "01100000", -- 3271 - 0xcc7  :   96 - 0x60
    "00110000", -- 3272 - 0xcc8  :   48 - 0x30 -- plane 1
    "00000000", -- 3273 - 0xcc9  :    0 - 0x0
    "00000000", -- 3274 - 0xcca  :    0 - 0x0
    "00000000", -- 3275 - 0xccb  :    0 - 0x0
    "00000000", -- 3276 - 0xccc  :    0 - 0x0
    "01100000", -- 3277 - 0xccd  :   96 - 0x60
    "01100000", -- 3278 - 0xcce  :   96 - 0x60
    "00000000", -- 3279 - 0xccf  :    0 - 0x0
    "11000000", -- 3280 - 0xcd0  :  192 - 0xc0 -- Sprite 0xcd
    "00000000", -- 3281 - 0xcd1  :    0 - 0x0
    "00000000", -- 3282 - 0xcd2  :    0 - 0x0
    "00000110", -- 3283 - 0xcd3  :    6 - 0x6
    "00001111", -- 3284 - 0xcd4  :   15 - 0xf
    "00001101", -- 3285 - 0xcd5  :   13 - 0xd
    "00001001", -- 3286 - 0xcd6  :    9 - 0x9
    "00000110", -- 3287 - 0xcd7  :    6 - 0x6
    "00000000", -- 3288 - 0xcd8  :    0 - 0x0 -- plane 1
    "00000000", -- 3289 - 0xcd9  :    0 - 0x0
    "00000000", -- 3290 - 0xcda  :    0 - 0x0
    "00000000", -- 3291 - 0xcdb  :    0 - 0x0
    "00000000", -- 3292 - 0xcdc  :    0 - 0x0
    "00000110", -- 3293 - 0xcdd  :    6 - 0x6
    "00000110", -- 3294 - 0xcde  :    6 - 0x6
    "00000000", -- 3295 - 0xcdf  :    0 - 0x0
    "11111100", -- 3296 - 0xce0  :  252 - 0xfc -- Sprite 0xce
    "11000000", -- 3297 - 0xce1  :  192 - 0xc0
    "11010001", -- 3298 - 0xce2  :  209 - 0xd1
    "11000010", -- 3299 - 0xce3  :  194 - 0xc2
    "10011110", -- 3300 - 0xce4  :  158 - 0x9e
    "10111111", -- 3301 - 0xce5  :  191 - 0xbf
    "10110000", -- 3302 - 0xce6  :  176 - 0xb0
    "10110011", -- 3303 - 0xce7  :  179 - 0xb3
    "00000000", -- 3304 - 0xce8  :    0 - 0x0 -- plane 1
    "00000001", -- 3305 - 0xce9  :    1 - 0x1
    "00011011", -- 3306 - 0xcea  :   27 - 0x1b
    "00010011", -- 3307 - 0xceb  :   19 - 0x13
    "00011111", -- 3308 - 0xcec  :   31 - 0x1f
    "00111111", -- 3309 - 0xced  :   63 - 0x3f
    "00111111", -- 3310 - 0xcee  :   63 - 0x3f
    "00111111", -- 3311 - 0xcef  :   63 - 0x3f
    "00000111", -- 3312 - 0xcf0  :    7 - 0x7 -- Sprite 0xcf
    "11110011", -- 3313 - 0xcf1  :  243 - 0xf3
    "00001011", -- 3314 - 0xcf2  :   11 - 0xb
    "01111011", -- 3315 - 0xcf3  :  123 - 0x7b
    "01111011", -- 3316 - 0xcf4  :  123 - 0x7b
    "11111001", -- 3317 - 0xcf5  :  249 - 0xf9
    "00001101", -- 3318 - 0xcf6  :   13 - 0xd
    "11101101", -- 3319 - 0xcf7  :  237 - 0xed
    "00000000", -- 3320 - 0xcf8  :    0 - 0x0 -- plane 1
    "11111000", -- 3321 - 0xcf9  :  248 - 0xf8
    "00001000", -- 3322 - 0xcfa  :    8 - 0x8
    "00001000", -- 3323 - 0xcfb  :    8 - 0x8
    "00001000", -- 3324 - 0xcfc  :    8 - 0x8
    "11111000", -- 3325 - 0xcfd  :  248 - 0xf8
    "11110000", -- 3326 - 0xcfe  :  240 - 0xf0
    "11010000", -- 3327 - 0xcff  :  208 - 0xd0
    "11111111", -- 3328 - 0xd00  :  255 - 0xff -- Sprite 0xd0
    "11111111", -- 3329 - 0xd01  :  255 - 0xff
    "11111111", -- 3330 - 0xd02  :  255 - 0xff
    "11111111", -- 3331 - 0xd03  :  255 - 0xff
    "11101110", -- 3332 - 0xd04  :  238 - 0xee
    "11101110", -- 3333 - 0xd05  :  238 - 0xee
    "11101110", -- 3334 - 0xd06  :  238 - 0xee
    "11101110", -- 3335 - 0xd07  :  238 - 0xee
    "00000000", -- 3336 - 0xd08  :    0 - 0x0 -- plane 1
    "00000000", -- 3337 - 0xd09  :    0 - 0x0
    "01111100", -- 3338 - 0xd0a  :  124 - 0x7c
    "11111110", -- 3339 - 0xd0b  :  254 - 0xfe
    "11101110", -- 3340 - 0xd0c  :  238 - 0xee
    "11101110", -- 3341 - 0xd0d  :  238 - 0xee
    "11101110", -- 3342 - 0xd0e  :  238 - 0xee
    "11101110", -- 3343 - 0xd0f  :  238 - 0xee
    "11111111", -- 3344 - 0xd10  :  255 - 0xff -- Sprite 0xd1
    "11111111", -- 3345 - 0xd11  :  255 - 0xff
    "11111111", -- 3346 - 0xd12  :  255 - 0xff
    "11111011", -- 3347 - 0xd13  :  251 - 0xfb
    "11111011", -- 3348 - 0xd14  :  251 - 0xfb
    "11111011", -- 3349 - 0xd15  :  251 - 0xfb
    "11111011", -- 3350 - 0xd16  :  251 - 0xfb
    "11111011", -- 3351 - 0xd17  :  251 - 0xfb
    "00000000", -- 3352 - 0xd18  :    0 - 0x0 -- plane 1
    "00000000", -- 3353 - 0xd19  :    0 - 0x0
    "00111000", -- 3354 - 0xd1a  :   56 - 0x38
    "01111000", -- 3355 - 0xd1b  :  120 - 0x78
    "01111000", -- 3356 - 0xd1c  :  120 - 0x78
    "00111000", -- 3357 - 0xd1d  :   56 - 0x38
    "00111000", -- 3358 - 0xd1e  :   56 - 0x38
    "00111000", -- 3359 - 0xd1f  :   56 - 0x38
    "11111111", -- 3360 - 0xd20  :  255 - 0xff -- Sprite 0xd2
    "11111111", -- 3361 - 0xd21  :  255 - 0xff
    "11111111", -- 3362 - 0xd22  :  255 - 0xff
    "11111111", -- 3363 - 0xd23  :  255 - 0xff
    "11101110", -- 3364 - 0xd24  :  238 - 0xee
    "10001110", -- 3365 - 0xd25  :  142 - 0x8e
    "11111110", -- 3366 - 0xd26  :  254 - 0xfe
    "11111110", -- 3367 - 0xd27  :  254 - 0xfe
    "00000000", -- 3368 - 0xd28  :    0 - 0x0 -- plane 1
    "00000000", -- 3369 - 0xd29  :    0 - 0x0
    "01111100", -- 3370 - 0xd2a  :  124 - 0x7c
    "11111110", -- 3371 - 0xd2b  :  254 - 0xfe
    "11101110", -- 3372 - 0xd2c  :  238 - 0xee
    "00001110", -- 3373 - 0xd2d  :   14 - 0xe
    "00001110", -- 3374 - 0xd2e  :   14 - 0xe
    "01111110", -- 3375 - 0xd2f  :  126 - 0x7e
    "11111111", -- 3376 - 0xd30  :  255 - 0xff -- Sprite 0xd3
    "11111111", -- 3377 - 0xd31  :  255 - 0xff
    "11111111", -- 3378 - 0xd32  :  255 - 0xff
    "11111111", -- 3379 - 0xd33  :  255 - 0xff
    "11101110", -- 3380 - 0xd34  :  238 - 0xee
    "10001110", -- 3381 - 0xd35  :  142 - 0x8e
    "11111100", -- 3382 - 0xd36  :  252 - 0xfc
    "11111101", -- 3383 - 0xd37  :  253 - 0xfd
    "00000000", -- 3384 - 0xd38  :    0 - 0x0 -- plane 1
    "00000000", -- 3385 - 0xd39  :    0 - 0x0
    "01111100", -- 3386 - 0xd3a  :  124 - 0x7c
    "11111110", -- 3387 - 0xd3b  :  254 - 0xfe
    "11101110", -- 3388 - 0xd3c  :  238 - 0xee
    "00001110", -- 3389 - 0xd3d  :   14 - 0xe
    "00111100", -- 3390 - 0xd3e  :   60 - 0x3c
    "00111100", -- 3391 - 0xd3f  :   60 - 0x3c
    "11111111", -- 3392 - 0xd40  :  255 - 0xff -- Sprite 0xd4
    "11111111", -- 3393 - 0xd41  :  255 - 0xff
    "11111111", -- 3394 - 0xd42  :  255 - 0xff
    "11111110", -- 3395 - 0xd43  :  254 - 0xfe
    "11101110", -- 3396 - 0xd44  :  238 - 0xee
    "11101110", -- 3397 - 0xd45  :  238 - 0xee
    "11101110", -- 3398 - 0xd46  :  238 - 0xee
    "11101110", -- 3399 - 0xd47  :  238 - 0xee
    "00000000", -- 3400 - 0xd48  :    0 - 0x0 -- plane 1
    "00000000", -- 3401 - 0xd49  :    0 - 0x0
    "00111110", -- 3402 - 0xd4a  :   62 - 0x3e
    "01111110", -- 3403 - 0xd4b  :  126 - 0x7e
    "11101110", -- 3404 - 0xd4c  :  238 - 0xee
    "11101110", -- 3405 - 0xd4d  :  238 - 0xee
    "11101110", -- 3406 - 0xd4e  :  238 - 0xee
    "11101110", -- 3407 - 0xd4f  :  238 - 0xee
    "11111111", -- 3408 - 0xd50  :  255 - 0xff -- Sprite 0xd5
    "11111111", -- 3409 - 0xd51  :  255 - 0xff
    "11111111", -- 3410 - 0xd52  :  255 - 0xff
    "11111101", -- 3411 - 0xd53  :  253 - 0xfd
    "11100001", -- 3412 - 0xd54  :  225 - 0xe1
    "11101111", -- 3413 - 0xd55  :  239 - 0xef
    "11111111", -- 3414 - 0xd56  :  255 - 0xff
    "11111111", -- 3415 - 0xd57  :  255 - 0xff
    "00000000", -- 3416 - 0xd58  :    0 - 0x0 -- plane 1
    "00000000", -- 3417 - 0xd59  :    0 - 0x0
    "11111100", -- 3418 - 0xd5a  :  252 - 0xfc
    "11111100", -- 3419 - 0xd5b  :  252 - 0xfc
    "11100000", -- 3420 - 0xd5c  :  224 - 0xe0
    "11100000", -- 3421 - 0xd5d  :  224 - 0xe0
    "11111100", -- 3422 - 0xd5e  :  252 - 0xfc
    "11111110", -- 3423 - 0xd5f  :  254 - 0xfe
    "11111111", -- 3424 - 0xd60  :  255 - 0xff -- Sprite 0xd6
    "11111111", -- 3425 - 0xd61  :  255 - 0xff
    "11111111", -- 3426 - 0xd62  :  255 - 0xff
    "11111101", -- 3427 - 0xd63  :  253 - 0xfd
    "11100001", -- 3428 - 0xd64  :  225 - 0xe1
    "11101111", -- 3429 - 0xd65  :  239 - 0xef
    "11111111", -- 3430 - 0xd66  :  255 - 0xff
    "11111111", -- 3431 - 0xd67  :  255 - 0xff
    "00000000", -- 3432 - 0xd68  :    0 - 0x0 -- plane 1
    "00000000", -- 3433 - 0xd69  :    0 - 0x0
    "01111100", -- 3434 - 0xd6a  :  124 - 0x7c
    "11111100", -- 3435 - 0xd6b  :  252 - 0xfc
    "11100000", -- 3436 - 0xd6c  :  224 - 0xe0
    "11100000", -- 3437 - 0xd6d  :  224 - 0xe0
    "11111100", -- 3438 - 0xd6e  :  252 - 0xfc
    "11111110", -- 3439 - 0xd6f  :  254 - 0xfe
    "11111111", -- 3440 - 0xd70  :  255 - 0xff -- Sprite 0xd7
    "11111111", -- 3441 - 0xd71  :  255 - 0xff
    "11111111", -- 3442 - 0xd72  :  255 - 0xff
    "11111110", -- 3443 - 0xd73  :  254 - 0xfe
    "11101110", -- 3444 - 0xd74  :  238 - 0xee
    "10001110", -- 3445 - 0xd75  :  142 - 0x8e
    "11111110", -- 3446 - 0xd76  :  254 - 0xfe
    "11111100", -- 3447 - 0xd77  :  252 - 0xfc
    "00000000", -- 3448 - 0xd78  :    0 - 0x0 -- plane 1
    "00000000", -- 3449 - 0xd79  :    0 - 0x0
    "11111110", -- 3450 - 0xd7a  :  254 - 0xfe
    "11111110", -- 3451 - 0xd7b  :  254 - 0xfe
    "11101110", -- 3452 - 0xd7c  :  238 - 0xee
    "00001110", -- 3453 - 0xd7d  :   14 - 0xe
    "00001110", -- 3454 - 0xd7e  :   14 - 0xe
    "00011100", -- 3455 - 0xd7f  :   28 - 0x1c
    "11111111", -- 3456 - 0xd80  :  255 - 0xff -- Sprite 0xd8
    "11111111", -- 3457 - 0xd81  :  255 - 0xff
    "11111111", -- 3458 - 0xd82  :  255 - 0xff
    "11111111", -- 3459 - 0xd83  :  255 - 0xff
    "11101110", -- 3460 - 0xd84  :  238 - 0xee
    "11101110", -- 3461 - 0xd85  :  238 - 0xee
    "11111100", -- 3462 - 0xd86  :  252 - 0xfc
    "11111111", -- 3463 - 0xd87  :  255 - 0xff
    "00000000", -- 3464 - 0xd88  :    0 - 0x0 -- plane 1
    "00000000", -- 3465 - 0xd89  :    0 - 0x0
    "01111100", -- 3466 - 0xd8a  :  124 - 0x7c
    "11111110", -- 3467 - 0xd8b  :  254 - 0xfe
    "11101110", -- 3468 - 0xd8c  :  238 - 0xee
    "11101110", -- 3469 - 0xd8d  :  238 - 0xee
    "01111100", -- 3470 - 0xd8e  :  124 - 0x7c
    "11111110", -- 3471 - 0xd8f  :  254 - 0xfe
    "11111111", -- 3472 - 0xd90  :  255 - 0xff -- Sprite 0xd9
    "11111111", -- 3473 - 0xd91  :  255 - 0xff
    "11111111", -- 3474 - 0xd92  :  255 - 0xff
    "11111111", -- 3475 - 0xd93  :  255 - 0xff
    "11101110", -- 3476 - 0xd94  :  238 - 0xee
    "11101110", -- 3477 - 0xd95  :  238 - 0xee
    "11101110", -- 3478 - 0xd96  :  238 - 0xee
    "11101110", -- 3479 - 0xd97  :  238 - 0xee
    "00000000", -- 3480 - 0xd98  :    0 - 0x0 -- plane 1
    "00000000", -- 3481 - 0xd99  :    0 - 0x0
    "01111100", -- 3482 - 0xd9a  :  124 - 0x7c
    "11111110", -- 3483 - 0xd9b  :  254 - 0xfe
    "11101110", -- 3484 - 0xd9c  :  238 - 0xee
    "11101110", -- 3485 - 0xd9d  :  238 - 0xee
    "11101110", -- 3486 - 0xd9e  :  238 - 0xee
    "11101110", -- 3487 - 0xd9f  :  238 - 0xee
    "00000000", -- 3488 - 0xda0  :    0 - 0x0 -- Sprite 0xda
    "00000000", -- 3489 - 0xda1  :    0 - 0x0
    "00000000", -- 3490 - 0xda2  :    0 - 0x0
    "10000000", -- 3491 - 0xda3  :  128 - 0x80
    "00000000", -- 3492 - 0xda4  :    0 - 0x0
    "00000000", -- 3493 - 0xda5  :    0 - 0x0
    "00000100", -- 3494 - 0xda6  :    4 - 0x4
    "00000000", -- 3495 - 0xda7  :    0 - 0x0
    "00000000", -- 3496 - 0xda8  :    0 - 0x0 -- plane 1
    "00100000", -- 3497 - 0xda9  :   32 - 0x20
    "00000000", -- 3498 - 0xdaa  :    0 - 0x0
    "00000010", -- 3499 - 0xdab  :    2 - 0x2
    "00000000", -- 3500 - 0xdac  :    0 - 0x0
    "00100000", -- 3501 - 0xdad  :   32 - 0x20
    "00000000", -- 3502 - 0xdae  :    0 - 0x0
    "00000000", -- 3503 - 0xdaf  :    0 - 0x0
    "00000000", -- 3504 - 0xdb0  :    0 - 0x0 -- Sprite 0xdb
    "00000100", -- 3505 - 0xdb1  :    4 - 0x4
    "00000000", -- 3506 - 0xdb2  :    0 - 0x0
    "00010001", -- 3507 - 0xdb3  :   17 - 0x11
    "00000000", -- 3508 - 0xdb4  :    0 - 0x0
    "00000000", -- 3509 - 0xdb5  :    0 - 0x0
    "00000000", -- 3510 - 0xdb6  :    0 - 0x0
    "00100000", -- 3511 - 0xdb7  :   32 - 0x20
    "00100000", -- 3512 - 0xdb8  :   32 - 0x20 -- plane 1
    "00000000", -- 3513 - 0xdb9  :    0 - 0x0
    "00000000", -- 3514 - 0xdba  :    0 - 0x0
    "00000000", -- 3515 - 0xdbb  :    0 - 0x0
    "10000000", -- 3516 - 0xdbc  :  128 - 0x80
    "00000000", -- 3517 - 0xdbd  :    0 - 0x0
    "00000100", -- 3518 - 0xdbe  :    4 - 0x4
    "00000000", -- 3519 - 0xdbf  :    0 - 0x0
    "00000000", -- 3520 - 0xdc0  :    0 - 0x0 -- Sprite 0xdc
    "00000000", -- 3521 - 0xdc1  :    0 - 0x0
    "00000000", -- 3522 - 0xdc2  :    0 - 0x0
    "00100000", -- 3523 - 0xdc3  :   32 - 0x20
    "00000000", -- 3524 - 0xdc4  :    0 - 0x0
    "00000000", -- 3525 - 0xdc5  :    0 - 0x0
    "00000000", -- 3526 - 0xdc6  :    0 - 0x0
    "00000100", -- 3527 - 0xdc7  :    4 - 0x4
    "00000000", -- 3528 - 0xdc8  :    0 - 0x0 -- plane 1
    "00001000", -- 3529 - 0xdc9  :    8 - 0x8
    "00000000", -- 3530 - 0xdca  :    0 - 0x0
    "00000000", -- 3531 - 0xdcb  :    0 - 0x0
    "00000010", -- 3532 - 0xdcc  :    2 - 0x2
    "00000000", -- 3533 - 0xdcd  :    0 - 0x0
    "01000000", -- 3534 - 0xdce  :   64 - 0x40
    "00000000", -- 3535 - 0xdcf  :    0 - 0x0
    "00000000", -- 3536 - 0xdd0  :    0 - 0x0 -- Sprite 0xdd
    "00000000", -- 3537 - 0xdd1  :    0 - 0x0
    "00010001", -- 3538 - 0xdd2  :   17 - 0x11
    "00000000", -- 3539 - 0xdd3  :    0 - 0x0
    "00000000", -- 3540 - 0xdd4  :    0 - 0x0
    "10000000", -- 3541 - 0xdd5  :  128 - 0x80
    "00000000", -- 3542 - 0xdd6  :    0 - 0x0
    "00000000", -- 3543 - 0xdd7  :    0 - 0x0
    "00000000", -- 3544 - 0xdd8  :    0 - 0x0 -- plane 1
    "01000000", -- 3545 - 0xdd9  :   64 - 0x40
    "00000000", -- 3546 - 0xdda  :    0 - 0x0
    "00000000", -- 3547 - 0xddb  :    0 - 0x0
    "00000000", -- 3548 - 0xddc  :    0 - 0x0
    "00000000", -- 3549 - 0xddd  :    0 - 0x0
    "00000010", -- 3550 - 0xdde  :    2 - 0x2
    "00100000", -- 3551 - 0xddf  :   32 - 0x20
    "10110011", -- 3552 - 0xde0  :  179 - 0xb3 -- Sprite 0xde
    "10110011", -- 3553 - 0xde1  :  179 - 0xb3
    "10110011", -- 3554 - 0xde2  :  179 - 0xb3
    "10110011", -- 3555 - 0xde3  :  179 - 0xb3
    "10110000", -- 3556 - 0xde4  :  176 - 0xb0
    "10101111", -- 3557 - 0xde5  :  175 - 0xaf
    "10011111", -- 3558 - 0xde6  :  159 - 0x9f
    "11000000", -- 3559 - 0xde7  :  192 - 0xc0
    "00111110", -- 3560 - 0xde8  :   62 - 0x3e -- plane 1
    "00111111", -- 3561 - 0xde9  :   63 - 0x3f
    "00111110", -- 3562 - 0xdea  :   62 - 0x3e
    "00111100", -- 3563 - 0xdeb  :   60 - 0x3c
    "00111111", -- 3564 - 0xdec  :   63 - 0x3f
    "00110000", -- 3565 - 0xded  :   48 - 0x30
    "00000000", -- 3566 - 0xdee  :    0 - 0x0
    "00000000", -- 3567 - 0xdef  :    0 - 0x0
    "11101101", -- 3568 - 0xdf0  :  237 - 0xed -- Sprite 0xdf
    "11001101", -- 3569 - 0xdf1  :  205 - 0xcd
    "11001101", -- 3570 - 0xdf2  :  205 - 0xcd
    "00001101", -- 3571 - 0xdf3  :   13 - 0xd
    "00001101", -- 3572 - 0xdf4  :   13 - 0xd
    "11111101", -- 3573 - 0xdf5  :  253 - 0xfd
    "11111101", -- 3574 - 0xdf6  :  253 - 0xfd
    "00000011", -- 3575 - 0xdf7  :    3 - 0x3
    "00010000", -- 3576 - 0xdf8  :   16 - 0x10 -- plane 1
    "10110000", -- 3577 - 0xdf9  :  176 - 0xb0
    "00110000", -- 3578 - 0xdfa  :   48 - 0x30
    "11110000", -- 3579 - 0xdfb  :  240 - 0xf0
    "11110000", -- 3580 - 0xdfc  :  240 - 0xf0
    "00000000", -- 3581 - 0xdfd  :    0 - 0x0
    "00000000", -- 3582 - 0xdfe  :    0 - 0x0
    "00000000", -- 3583 - 0xdff  :    0 - 0x0
    "11101110", -- 3584 - 0xe00  :  238 - 0xee -- Sprite 0xe0
    "11101110", -- 3585 - 0xe01  :  238 - 0xee
    "11101110", -- 3586 - 0xe02  :  238 - 0xee
    "11101110", -- 3587 - 0xe03  :  238 - 0xee
    "11111110", -- 3588 - 0xe04  :  254 - 0xfe
    "11111100", -- 3589 - 0xe05  :  252 - 0xfc
    "11000001", -- 3590 - 0xe06  :  193 - 0xc1
    "11111111", -- 3591 - 0xe07  :  255 - 0xff
    "11101110", -- 3592 - 0xe08  :  238 - 0xee -- plane 1
    "11101110", -- 3593 - 0xe09  :  238 - 0xee
    "11101110", -- 3594 - 0xe0a  :  238 - 0xee
    "11101110", -- 3595 - 0xe0b  :  238 - 0xee
    "11111110", -- 3596 - 0xe0c  :  254 - 0xfe
    "01111100", -- 3597 - 0xe0d  :  124 - 0x7c
    "00000000", -- 3598 - 0xe0e  :    0 - 0x0
    "00000000", -- 3599 - 0xe0f  :    0 - 0x0
    "11111011", -- 3600 - 0xe10  :  251 - 0xfb -- Sprite 0xe1
    "11111011", -- 3601 - 0xe11  :  251 - 0xfb
    "11111011", -- 3602 - 0xe12  :  251 - 0xfb
    "11111011", -- 3603 - 0xe13  :  251 - 0xfb
    "11111111", -- 3604 - 0xe14  :  255 - 0xff
    "11111101", -- 3605 - 0xe15  :  253 - 0xfd
    "11000001", -- 3606 - 0xe16  :  193 - 0xc1
    "11111111", -- 3607 - 0xe17  :  255 - 0xff
    "00111000", -- 3608 - 0xe18  :   56 - 0x38 -- plane 1
    "00111000", -- 3609 - 0xe19  :   56 - 0x38
    "00111000", -- 3610 - 0xe1a  :   56 - 0x38
    "00111000", -- 3611 - 0xe1b  :   56 - 0x38
    "01111100", -- 3612 - 0xe1c  :  124 - 0x7c
    "01111100", -- 3613 - 0xe1d  :  124 - 0x7c
    "00000000", -- 3614 - 0xe1e  :    0 - 0x0
    "00000000", -- 3615 - 0xe1f  :    0 - 0x0
    "11111100", -- 3616 - 0xe20  :  252 - 0xfc -- Sprite 0xe2
    "11100001", -- 3617 - 0xe21  :  225 - 0xe1
    "11101111", -- 3618 - 0xe22  :  239 - 0xef
    "11101111", -- 3619 - 0xe23  :  239 - 0xef
    "11111111", -- 3620 - 0xe24  :  255 - 0xff
    "11111110", -- 3621 - 0xe25  :  254 - 0xfe
    "10000000", -- 3622 - 0xe26  :  128 - 0x80
    "11111111", -- 3623 - 0xe27  :  255 - 0xff
    "11111100", -- 3624 - 0xe28  :  252 - 0xfc -- plane 1
    "11100000", -- 3625 - 0xe29  :  224 - 0xe0
    "11100000", -- 3626 - 0xe2a  :  224 - 0xe0
    "11100000", -- 3627 - 0xe2b  :  224 - 0xe0
    "11111110", -- 3628 - 0xe2c  :  254 - 0xfe
    "11111110", -- 3629 - 0xe2d  :  254 - 0xfe
    "00000000", -- 3630 - 0xe2e  :    0 - 0x0
    "00000000", -- 3631 - 0xe2f  :    0 - 0x0
    "11101110", -- 3632 - 0xe30  :  238 - 0xee -- Sprite 0xe3
    "11111110", -- 3633 - 0xe31  :  254 - 0xfe
    "11111110", -- 3634 - 0xe32  :  254 - 0xfe
    "11111110", -- 3635 - 0xe33  :  254 - 0xfe
    "11111110", -- 3636 - 0xe34  :  254 - 0xfe
    "11111100", -- 3637 - 0xe35  :  252 - 0xfc
    "11000001", -- 3638 - 0xe36  :  193 - 0xc1
    "11111111", -- 3639 - 0xe37  :  255 - 0xff
    "00001110", -- 3640 - 0xe38  :   14 - 0xe -- plane 1
    "00001110", -- 3641 - 0xe39  :   14 - 0xe
    "00001110", -- 3642 - 0xe3a  :   14 - 0xe
    "11101110", -- 3643 - 0xe3b  :  238 - 0xee
    "11111110", -- 3644 - 0xe3c  :  254 - 0xfe
    "01111100", -- 3645 - 0xe3d  :  124 - 0x7c
    "00000000", -- 3646 - 0xe3e  :    0 - 0x0
    "00000000", -- 3647 - 0xe3f  :    0 - 0x0
    "11101110", -- 3648 - 0xe40  :  238 - 0xee -- Sprite 0xe4
    "11101110", -- 3649 - 0xe41  :  238 - 0xee
    "11111110", -- 3650 - 0xe42  :  254 - 0xfe
    "11111110", -- 3651 - 0xe43  :  254 - 0xfe
    "10001110", -- 3652 - 0xe44  :  142 - 0x8e
    "11111110", -- 3653 - 0xe45  :  254 - 0xfe
    "11111000", -- 3654 - 0xe46  :  248 - 0xf8
    "11111111", -- 3655 - 0xe47  :  255 - 0xff
    "11101110", -- 3656 - 0xe48  :  238 - 0xee -- plane 1
    "11101110", -- 3657 - 0xe49  :  238 - 0xee
    "11111110", -- 3658 - 0xe4a  :  254 - 0xfe
    "11111110", -- 3659 - 0xe4b  :  254 - 0xfe
    "00001110", -- 3660 - 0xe4c  :   14 - 0xe
    "00001110", -- 3661 - 0xe4d  :   14 - 0xe
    "00000000", -- 3662 - 0xe4e  :    0 - 0x0
    "00000000", -- 3663 - 0xe4f  :    0 - 0x0
    "10001110", -- 3664 - 0xe50  :  142 - 0x8e -- Sprite 0xe5
    "11111110", -- 3665 - 0xe51  :  254 - 0xfe
    "11111110", -- 3666 - 0xe52  :  254 - 0xfe
    "11111110", -- 3667 - 0xe53  :  254 - 0xfe
    "11111110", -- 3668 - 0xe54  :  254 - 0xfe
    "11111100", -- 3669 - 0xe55  :  252 - 0xfc
    "11000001", -- 3670 - 0xe56  :  193 - 0xc1
    "11111111", -- 3671 - 0xe57  :  255 - 0xff
    "00001110", -- 3672 - 0xe58  :   14 - 0xe -- plane 1
    "00001110", -- 3673 - 0xe59  :   14 - 0xe
    "00001110", -- 3674 - 0xe5a  :   14 - 0xe
    "11101110", -- 3675 - 0xe5b  :  238 - 0xee
    "11111110", -- 3676 - 0xe5c  :  254 - 0xfe
    "01111100", -- 3677 - 0xe5d  :  124 - 0x7c
    "00000000", -- 3678 - 0xe5e  :    0 - 0x0
    "00000000", -- 3679 - 0xe5f  :    0 - 0x0
    "11101110", -- 3680 - 0xe60  :  238 - 0xee -- Sprite 0xe6
    "11101110", -- 3681 - 0xe61  :  238 - 0xee
    "11101110", -- 3682 - 0xe62  :  238 - 0xee
    "11101110", -- 3683 - 0xe63  :  238 - 0xee
    "11111110", -- 3684 - 0xe64  :  254 - 0xfe
    "11111100", -- 3685 - 0xe65  :  252 - 0xfc
    "11000001", -- 3686 - 0xe66  :  193 - 0xc1
    "11111111", -- 3687 - 0xe67  :  255 - 0xff
    "11101110", -- 3688 - 0xe68  :  238 - 0xee -- plane 1
    "11101110", -- 3689 - 0xe69  :  238 - 0xee
    "11101110", -- 3690 - 0xe6a  :  238 - 0xee
    "11101110", -- 3691 - 0xe6b  :  238 - 0xee
    "11111110", -- 3692 - 0xe6c  :  254 - 0xfe
    "01111100", -- 3693 - 0xe6d  :  124 - 0x7c
    "00000000", -- 3694 - 0xe6e  :    0 - 0x0
    "00000000", -- 3695 - 0xe6f  :    0 - 0x0
    "11111101", -- 3696 - 0xe70  :  253 - 0xfd -- Sprite 0xe7
    "11111101", -- 3697 - 0xe71  :  253 - 0xfd
    "11111001", -- 3698 - 0xe72  :  249 - 0xf9
    "11111011", -- 3699 - 0xe73  :  251 - 0xfb
    "11111011", -- 3700 - 0xe74  :  251 - 0xfb
    "11111011", -- 3701 - 0xe75  :  251 - 0xfb
    "11100011", -- 3702 - 0xe76  :  227 - 0xe3
    "11111111", -- 3703 - 0xe77  :  255 - 0xff
    "00011100", -- 3704 - 0xe78  :   28 - 0x1c -- plane 1
    "00011100", -- 3705 - 0xe79  :   28 - 0x1c
    "00111000", -- 3706 - 0xe7a  :   56 - 0x38
    "00111000", -- 3707 - 0xe7b  :   56 - 0x38
    "00111000", -- 3708 - 0xe7c  :   56 - 0x38
    "00111000", -- 3709 - 0xe7d  :   56 - 0x38
    "00000000", -- 3710 - 0xe7e  :    0 - 0x0
    "00000000", -- 3711 - 0xe7f  :    0 - 0x0
    "11101110", -- 3712 - 0xe80  :  238 - 0xee -- Sprite 0xe8
    "11101110", -- 3713 - 0xe81  :  238 - 0xee
    "11101110", -- 3714 - 0xe82  :  238 - 0xee
    "11101110", -- 3715 - 0xe83  :  238 - 0xee
    "11111110", -- 3716 - 0xe84  :  254 - 0xfe
    "11111100", -- 3717 - 0xe85  :  252 - 0xfc
    "11000001", -- 3718 - 0xe86  :  193 - 0xc1
    "11111111", -- 3719 - 0xe87  :  255 - 0xff
    "11101110", -- 3720 - 0xe88  :  238 - 0xee -- plane 1
    "11101110", -- 3721 - 0xe89  :  238 - 0xee
    "11101110", -- 3722 - 0xe8a  :  238 - 0xee
    "11101110", -- 3723 - 0xe8b  :  238 - 0xee
    "11111110", -- 3724 - 0xe8c  :  254 - 0xfe
    "01111100", -- 3725 - 0xe8d  :  124 - 0x7c
    "00000000", -- 3726 - 0xe8e  :    0 - 0x0
    "00000000", -- 3727 - 0xe8f  :    0 - 0x0
    "11111110", -- 3728 - 0xe90  :  254 - 0xfe -- Sprite 0xe9
    "11111110", -- 3729 - 0xe91  :  254 - 0xfe
    "11001110", -- 3730 - 0xe92  :  206 - 0xce
    "11111110", -- 3731 - 0xe93  :  254 - 0xfe
    "11111110", -- 3732 - 0xe94  :  254 - 0xfe
    "11111100", -- 3733 - 0xe95  :  252 - 0xfc
    "11000001", -- 3734 - 0xe96  :  193 - 0xc1
    "11111111", -- 3735 - 0xe97  :  255 - 0xff
    "11111110", -- 3736 - 0xe98  :  254 - 0xfe -- plane 1
    "01111110", -- 3737 - 0xe99  :  126 - 0x7e
    "00001110", -- 3738 - 0xe9a  :   14 - 0xe
    "00001110", -- 3739 - 0xe9b  :   14 - 0xe
    "01111110", -- 3740 - 0xe9c  :  126 - 0x7e
    "01111100", -- 3741 - 0xe9d  :  124 - 0x7c
    "00000000", -- 3742 - 0xe9e  :    0 - 0x0
    "00000000", -- 3743 - 0xe9f  :    0 - 0x0
    "00000000", -- 3744 - 0xea0  :    0 - 0x0 -- Sprite 0xea
    "01110000", -- 3745 - 0xea1  :  112 - 0x70
    "00111000", -- 3746 - 0xea2  :   56 - 0x38
    "00000000", -- 3747 - 0xea3  :    0 - 0x0
    "00000010", -- 3748 - 0xea4  :    2 - 0x2
    "00000111", -- 3749 - 0xea5  :    7 - 0x7
    "00000011", -- 3750 - 0xea6  :    3 - 0x3
    "00000000", -- 3751 - 0xea7  :    0 - 0x0
    "00000000", -- 3752 - 0xea8  :    0 - 0x0 -- plane 1
    "01110000", -- 3753 - 0xea9  :  112 - 0x70
    "00111000", -- 3754 - 0xeaa  :   56 - 0x38
    "00000000", -- 3755 - 0xeab  :    0 - 0x0
    "00000010", -- 3756 - 0xeac  :    2 - 0x2
    "00000111", -- 3757 - 0xead  :    7 - 0x7
    "00000011", -- 3758 - 0xeae  :    3 - 0x3
    "00000000", -- 3759 - 0xeaf  :    0 - 0x0
    "00000000", -- 3760 - 0xeb0  :    0 - 0x0 -- Sprite 0xeb
    "00001100", -- 3761 - 0xeb1  :   12 - 0xc
    "00000110", -- 3762 - 0xeb2  :    6 - 0x6
    "00000110", -- 3763 - 0xeb3  :    6 - 0x6
    "01100000", -- 3764 - 0xeb4  :   96 - 0x60
    "01110000", -- 3765 - 0xeb5  :  112 - 0x70
    "00110000", -- 3766 - 0xeb6  :   48 - 0x30
    "00000000", -- 3767 - 0xeb7  :    0 - 0x0
    "00000000", -- 3768 - 0xeb8  :    0 - 0x0 -- plane 1
    "00001100", -- 3769 - 0xeb9  :   12 - 0xc
    "00000110", -- 3770 - 0xeba  :    6 - 0x6
    "00000110", -- 3771 - 0xebb  :    6 - 0x6
    "01100000", -- 3772 - 0xebc  :   96 - 0x60
    "01110000", -- 3773 - 0xebd  :  112 - 0x70
    "00110000", -- 3774 - 0xebe  :   48 - 0x30
    "00000000", -- 3775 - 0xebf  :    0 - 0x0
    "00000000", -- 3776 - 0xec0  :    0 - 0x0 -- Sprite 0xec
    "11000000", -- 3777 - 0xec1  :  192 - 0xc0
    "11100000", -- 3778 - 0xec2  :  224 - 0xe0
    "01100000", -- 3779 - 0xec3  :   96 - 0x60
    "00000000", -- 3780 - 0xec4  :    0 - 0x0
    "00001100", -- 3781 - 0xec5  :   12 - 0xc
    "00001110", -- 3782 - 0xec6  :   14 - 0xe
    "00000110", -- 3783 - 0xec7  :    6 - 0x6
    "00000000", -- 3784 - 0xec8  :    0 - 0x0 -- plane 1
    "11000000", -- 3785 - 0xec9  :  192 - 0xc0
    "11100000", -- 3786 - 0xeca  :  224 - 0xe0
    "01100000", -- 3787 - 0xecb  :   96 - 0x60
    "00000000", -- 3788 - 0xecc  :    0 - 0x0
    "00001100", -- 3789 - 0xecd  :   12 - 0xc
    "00001110", -- 3790 - 0xece  :   14 - 0xe
    "00000110", -- 3791 - 0xecf  :    6 - 0x6
    "01100000", -- 3792 - 0xed0  :   96 - 0x60 -- Sprite 0xed
    "01110000", -- 3793 - 0xed1  :  112 - 0x70
    "00110000", -- 3794 - 0xed2  :   48 - 0x30
    "00000000", -- 3795 - 0xed3  :    0 - 0x0
    "00000000", -- 3796 - 0xed4  :    0 - 0x0
    "00001100", -- 3797 - 0xed5  :   12 - 0xc
    "00001110", -- 3798 - 0xed6  :   14 - 0xe
    "00000110", -- 3799 - 0xed7  :    6 - 0x6
    "01100000", -- 3800 - 0xed8  :   96 - 0x60 -- plane 1
    "01110000", -- 3801 - 0xed9  :  112 - 0x70
    "00110000", -- 3802 - 0xeda  :   48 - 0x30
    "00000000", -- 3803 - 0xedb  :    0 - 0x0
    "00000000", -- 3804 - 0xedc  :    0 - 0x0
    "00001100", -- 3805 - 0xedd  :   12 - 0xc
    "00001110", -- 3806 - 0xede  :   14 - 0xe
    "00000110", -- 3807 - 0xedf  :    6 - 0x6
    "11111111", -- 3808 - 0xee0  :  255 - 0xff -- Sprite 0xee
    "11111111", -- 3809 - 0xee1  :  255 - 0xff
    "10111101", -- 3810 - 0xee2  :  189 - 0xbd
    "11111111", -- 3811 - 0xee3  :  255 - 0xff
    "11111111", -- 3812 - 0xee4  :  255 - 0xff
    "11111011", -- 3813 - 0xee5  :  251 - 0xfb
    "11111111", -- 3814 - 0xee6  :  255 - 0xff
    "11111111", -- 3815 - 0xee7  :  255 - 0xff
    "00000000", -- 3816 - 0xee8  :    0 - 0x0 -- plane 1
    "00000000", -- 3817 - 0xee9  :    0 - 0x0
    "01000010", -- 3818 - 0xeea  :   66 - 0x42
    "00000000", -- 3819 - 0xeeb  :    0 - 0x0
    "00000000", -- 3820 - 0xeec  :    0 - 0x0
    "00000100", -- 3821 - 0xeed  :    4 - 0x4
    "00000000", -- 3822 - 0xeee  :    0 - 0x0
    "00000000", -- 3823 - 0xeef  :    0 - 0x0
    "11111111", -- 3824 - 0xef0  :  255 - 0xff -- Sprite 0xef
    "11111111", -- 3825 - 0xef1  :  255 - 0xff
    "11111011", -- 3826 - 0xef2  :  251 - 0xfb
    "11111111", -- 3827 - 0xef3  :  255 - 0xff
    "11011111", -- 3828 - 0xef4  :  223 - 0xdf
    "11111111", -- 3829 - 0xef5  :  255 - 0xff
    "11111111", -- 3830 - 0xef6  :  255 - 0xff
    "11111111", -- 3831 - 0xef7  :  255 - 0xff
    "00000000", -- 3832 - 0xef8  :    0 - 0x0 -- plane 1
    "00000000", -- 3833 - 0xef9  :    0 - 0x0
    "00000100", -- 3834 - 0xefa  :    4 - 0x4
    "00000000", -- 3835 - 0xefb  :    0 - 0x0
    "00100000", -- 3836 - 0xefc  :   32 - 0x20
    "00000000", -- 3837 - 0xefd  :    0 - 0x0
    "00000000", -- 3838 - 0xefe  :    0 - 0x0
    "00000000", -- 3839 - 0xeff  :    0 - 0x0
    "00000000", -- 3840 - 0xf00  :    0 - 0x0 -- Sprite 0xf0
    "00000000", -- 3841 - 0xf01  :    0 - 0x0
    "00000000", -- 3842 - 0xf02  :    0 - 0x0
    "00000000", -- 3843 - 0xf03  :    0 - 0x0
    "00000000", -- 3844 - 0xf04  :    0 - 0x0
    "00000000", -- 3845 - 0xf05  :    0 - 0x0
    "00000000", -- 3846 - 0xf06  :    0 - 0x0
    "00000000", -- 3847 - 0xf07  :    0 - 0x0
    "00000000", -- 3848 - 0xf08  :    0 - 0x0 -- plane 1
    "00000000", -- 3849 - 0xf09  :    0 - 0x0
    "00000000", -- 3850 - 0xf0a  :    0 - 0x0
    "00000000", -- 3851 - 0xf0b  :    0 - 0x0
    "00000000", -- 3852 - 0xf0c  :    0 - 0x0
    "00000000", -- 3853 - 0xf0d  :    0 - 0x0
    "00000000", -- 3854 - 0xf0e  :    0 - 0x0
    "00000000", -- 3855 - 0xf0f  :    0 - 0x0
    "00000000", -- 3856 - 0xf10  :    0 - 0x0 -- Sprite 0xf1
    "10000000", -- 3857 - 0xf11  :  128 - 0x80
    "00000000", -- 3858 - 0xf12  :    0 - 0x0
    "00000000", -- 3859 - 0xf13  :    0 - 0x0
    "00000000", -- 3860 - 0xf14  :    0 - 0x0
    "00000000", -- 3861 - 0xf15  :    0 - 0x0
    "00000000", -- 3862 - 0xf16  :    0 - 0x0
    "00000000", -- 3863 - 0xf17  :    0 - 0x0
    "10000000", -- 3864 - 0xf18  :  128 - 0x80 -- plane 1
    "10000000", -- 3865 - 0xf19  :  128 - 0x80
    "10000000", -- 3866 - 0xf1a  :  128 - 0x80
    "10000000", -- 3867 - 0xf1b  :  128 - 0x80
    "00000000", -- 3868 - 0xf1c  :    0 - 0x0
    "00000000", -- 3869 - 0xf1d  :    0 - 0x0
    "00000000", -- 3870 - 0xf1e  :    0 - 0x0
    "00000000", -- 3871 - 0xf1f  :    0 - 0x0
    "00000000", -- 3872 - 0xf20  :    0 - 0x0 -- Sprite 0xf2
    "11000000", -- 3873 - 0xf21  :  192 - 0xc0
    "00000000", -- 3874 - 0xf22  :    0 - 0x0
    "00000000", -- 3875 - 0xf23  :    0 - 0x0
    "00000000", -- 3876 - 0xf24  :    0 - 0x0
    "00000000", -- 3877 - 0xf25  :    0 - 0x0
    "00000000", -- 3878 - 0xf26  :    0 - 0x0
    "00000000", -- 3879 - 0xf27  :    0 - 0x0
    "11000000", -- 3880 - 0xf28  :  192 - 0xc0 -- plane 1
    "11000000", -- 3881 - 0xf29  :  192 - 0xc0
    "11000000", -- 3882 - 0xf2a  :  192 - 0xc0
    "11000000", -- 3883 - 0xf2b  :  192 - 0xc0
    "00000000", -- 3884 - 0xf2c  :    0 - 0x0
    "00000000", -- 3885 - 0xf2d  :    0 - 0x0
    "00000000", -- 3886 - 0xf2e  :    0 - 0x0
    "00000000", -- 3887 - 0xf2f  :    0 - 0x0
    "00000000", -- 3888 - 0xf30  :    0 - 0x0 -- Sprite 0xf3
    "11100000", -- 3889 - 0xf31  :  224 - 0xe0
    "00000000", -- 3890 - 0xf32  :    0 - 0x0
    "00000000", -- 3891 - 0xf33  :    0 - 0x0
    "00000000", -- 3892 - 0xf34  :    0 - 0x0
    "00000000", -- 3893 - 0xf35  :    0 - 0x0
    "00000000", -- 3894 - 0xf36  :    0 - 0x0
    "00000000", -- 3895 - 0xf37  :    0 - 0x0
    "11100000", -- 3896 - 0xf38  :  224 - 0xe0 -- plane 1
    "11100000", -- 3897 - 0xf39  :  224 - 0xe0
    "11100000", -- 3898 - 0xf3a  :  224 - 0xe0
    "11100000", -- 3899 - 0xf3b  :  224 - 0xe0
    "00000000", -- 3900 - 0xf3c  :    0 - 0x0
    "00000000", -- 3901 - 0xf3d  :    0 - 0x0
    "00000000", -- 3902 - 0xf3e  :    0 - 0x0
    "00000000", -- 3903 - 0xf3f  :    0 - 0x0
    "00000000", -- 3904 - 0xf40  :    0 - 0x0 -- Sprite 0xf4
    "11110000", -- 3905 - 0xf41  :  240 - 0xf0
    "00000000", -- 3906 - 0xf42  :    0 - 0x0
    "00000000", -- 3907 - 0xf43  :    0 - 0x0
    "00000000", -- 3908 - 0xf44  :    0 - 0x0
    "00000000", -- 3909 - 0xf45  :    0 - 0x0
    "00000000", -- 3910 - 0xf46  :    0 - 0x0
    "00000000", -- 3911 - 0xf47  :    0 - 0x0
    "11110000", -- 3912 - 0xf48  :  240 - 0xf0 -- plane 1
    "11110000", -- 3913 - 0xf49  :  240 - 0xf0
    "11110000", -- 3914 - 0xf4a  :  240 - 0xf0
    "11110000", -- 3915 - 0xf4b  :  240 - 0xf0
    "00000000", -- 3916 - 0xf4c  :    0 - 0x0
    "00000000", -- 3917 - 0xf4d  :    0 - 0x0
    "00000000", -- 3918 - 0xf4e  :    0 - 0x0
    "00000000", -- 3919 - 0xf4f  :    0 - 0x0
    "00000000", -- 3920 - 0xf50  :    0 - 0x0 -- Sprite 0xf5
    "11111000", -- 3921 - 0xf51  :  248 - 0xf8
    "00000000", -- 3922 - 0xf52  :    0 - 0x0
    "00000000", -- 3923 - 0xf53  :    0 - 0x0
    "00000000", -- 3924 - 0xf54  :    0 - 0x0
    "00000000", -- 3925 - 0xf55  :    0 - 0x0
    "00000000", -- 3926 - 0xf56  :    0 - 0x0
    "00000000", -- 3927 - 0xf57  :    0 - 0x0
    "11111000", -- 3928 - 0xf58  :  248 - 0xf8 -- plane 1
    "11111000", -- 3929 - 0xf59  :  248 - 0xf8
    "11111000", -- 3930 - 0xf5a  :  248 - 0xf8
    "11111000", -- 3931 - 0xf5b  :  248 - 0xf8
    "00000000", -- 3932 - 0xf5c  :    0 - 0x0
    "00000000", -- 3933 - 0xf5d  :    0 - 0x0
    "00000000", -- 3934 - 0xf5e  :    0 - 0x0
    "00000000", -- 3935 - 0xf5f  :    0 - 0x0
    "00000000", -- 3936 - 0xf60  :    0 - 0x0 -- Sprite 0xf6
    "11111100", -- 3937 - 0xf61  :  252 - 0xfc
    "00000000", -- 3938 - 0xf62  :    0 - 0x0
    "00000000", -- 3939 - 0xf63  :    0 - 0x0
    "00000000", -- 3940 - 0xf64  :    0 - 0x0
    "00000000", -- 3941 - 0xf65  :    0 - 0x0
    "00000000", -- 3942 - 0xf66  :    0 - 0x0
    "00000000", -- 3943 - 0xf67  :    0 - 0x0
    "11111100", -- 3944 - 0xf68  :  252 - 0xfc -- plane 1
    "11111100", -- 3945 - 0xf69  :  252 - 0xfc
    "11111100", -- 3946 - 0xf6a  :  252 - 0xfc
    "11111100", -- 3947 - 0xf6b  :  252 - 0xfc
    "00000000", -- 3948 - 0xf6c  :    0 - 0x0
    "00000000", -- 3949 - 0xf6d  :    0 - 0x0
    "00000000", -- 3950 - 0xf6e  :    0 - 0x0
    "00000000", -- 3951 - 0xf6f  :    0 - 0x0
    "00000000", -- 3952 - 0xf70  :    0 - 0x0 -- Sprite 0xf7
    "11111110", -- 3953 - 0xf71  :  254 - 0xfe
    "00000000", -- 3954 - 0xf72  :    0 - 0x0
    "00000000", -- 3955 - 0xf73  :    0 - 0x0
    "00000000", -- 3956 - 0xf74  :    0 - 0x0
    "00000000", -- 3957 - 0xf75  :    0 - 0x0
    "00000000", -- 3958 - 0xf76  :    0 - 0x0
    "00000000", -- 3959 - 0xf77  :    0 - 0x0
    "11111110", -- 3960 - 0xf78  :  254 - 0xfe -- plane 1
    "11111110", -- 3961 - 0xf79  :  254 - 0xfe
    "11111110", -- 3962 - 0xf7a  :  254 - 0xfe
    "11111110", -- 3963 - 0xf7b  :  254 - 0xfe
    "00000000", -- 3964 - 0xf7c  :    0 - 0x0
    "00000000", -- 3965 - 0xf7d  :    0 - 0x0
    "00000000", -- 3966 - 0xf7e  :    0 - 0x0
    "00000000", -- 3967 - 0xf7f  :    0 - 0x0
    "00000000", -- 3968 - 0xf80  :    0 - 0x0 -- Sprite 0xf8
    "11111111", -- 3969 - 0xf81  :  255 - 0xff
    "00000000", -- 3970 - 0xf82  :    0 - 0x0
    "00000000", -- 3971 - 0xf83  :    0 - 0x0
    "00000000", -- 3972 - 0xf84  :    0 - 0x0
    "00000000", -- 3973 - 0xf85  :    0 - 0x0
    "00000000", -- 3974 - 0xf86  :    0 - 0x0
    "00000000", -- 3975 - 0xf87  :    0 - 0x0
    "11111111", -- 3976 - 0xf88  :  255 - 0xff -- plane 1
    "11111111", -- 3977 - 0xf89  :  255 - 0xff
    "11111111", -- 3978 - 0xf8a  :  255 - 0xff
    "11111111", -- 3979 - 0xf8b  :  255 - 0xff
    "00000000", -- 3980 - 0xf8c  :    0 - 0x0
    "00000000", -- 3981 - 0xf8d  :    0 - 0x0
    "00000000", -- 3982 - 0xf8e  :    0 - 0x0
    "00000000", -- 3983 - 0xf8f  :    0 - 0x0
    "11111111", -- 3984 - 0xf90  :  255 - 0xff -- Sprite 0xf9
    "11111111", -- 3985 - 0xf91  :  255 - 0xff
    "11111111", -- 3986 - 0xf92  :  255 - 0xff
    "11111111", -- 3987 - 0xf93  :  255 - 0xff
    "10000000", -- 3988 - 0xf94  :  128 - 0x80
    "10000000", -- 3989 - 0xf95  :  128 - 0x80
    "11000000", -- 3990 - 0xf96  :  192 - 0xc0
    "11000000", -- 3991 - 0xf97  :  192 - 0xc0
    "00000000", -- 3992 - 0xf98  :    0 - 0x0 -- plane 1
    "00000000", -- 3993 - 0xf99  :    0 - 0x0
    "00000000", -- 3994 - 0xf9a  :    0 - 0x0
    "00000000", -- 3995 - 0xf9b  :    0 - 0x0
    "01111111", -- 3996 - 0xf9c  :  127 - 0x7f
    "01000000", -- 3997 - 0xf9d  :   64 - 0x40
    "01000000", -- 3998 - 0xf9e  :   64 - 0x40
    "01000000", -- 3999 - 0xf9f  :   64 - 0x40
    "11111111", -- 4000 - 0xfa0  :  255 - 0xff -- Sprite 0xfa
    "11111111", -- 4001 - 0xfa1  :  255 - 0xff
    "11111111", -- 4002 - 0xfa2  :  255 - 0xff
    "11111111", -- 4003 - 0xfa3  :  255 - 0xff
    "00000000", -- 4004 - 0xfa4  :    0 - 0x0
    "00000000", -- 4005 - 0xfa5  :    0 - 0x0
    "00000000", -- 4006 - 0xfa6  :    0 - 0x0
    "00000000", -- 4007 - 0xfa7  :    0 - 0x0
    "00000000", -- 4008 - 0xfa8  :    0 - 0x0 -- plane 1
    "00000000", -- 4009 - 0xfa9  :    0 - 0x0
    "00000000", -- 4010 - 0xfaa  :    0 - 0x0
    "00000000", -- 4011 - 0xfab  :    0 - 0x0
    "11111111", -- 4012 - 0xfac  :  255 - 0xff
    "00000000", -- 4013 - 0xfad  :    0 - 0x0
    "00000000", -- 4014 - 0xfae  :    0 - 0x0
    "00000000", -- 4015 - 0xfaf  :    0 - 0x0
    "11111111", -- 4016 - 0xfb0  :  255 - 0xff -- Sprite 0xfb
    "11111111", -- 4017 - 0xfb1  :  255 - 0xff
    "11111111", -- 4018 - 0xfb2  :  255 - 0xff
    "11111111", -- 4019 - 0xfb3  :  255 - 0xff
    "00000001", -- 4020 - 0xfb4  :    1 - 0x1
    "00000000", -- 4021 - 0xfb5  :    0 - 0x0
    "00000010", -- 4022 - 0xfb6  :    2 - 0x2
    "00000010", -- 4023 - 0xfb7  :    2 - 0x2
    "00000000", -- 4024 - 0xfb8  :    0 - 0x0 -- plane 1
    "00000000", -- 4025 - 0xfb9  :    0 - 0x0
    "00000000", -- 4026 - 0xfba  :    0 - 0x0
    "00000000", -- 4027 - 0xfbb  :    0 - 0x0
    "11111110", -- 4028 - 0xfbc  :  254 - 0xfe
    "00000010", -- 4029 - 0xfbd  :    2 - 0x2
    "00000010", -- 4030 - 0xfbe  :    2 - 0x2
    "00000010", -- 4031 - 0xfbf  :    2 - 0x2
    "11000000", -- 4032 - 0xfc0  :  192 - 0xc0 -- Sprite 0xfc
    "11000000", -- 4033 - 0xfc1  :  192 - 0xc0
    "10000000", -- 4034 - 0xfc2  :  128 - 0x80
    "10000000", -- 4035 - 0xfc3  :  128 - 0x80
    "11000000", -- 4036 - 0xfc4  :  192 - 0xc0
    "11111111", -- 4037 - 0xfc5  :  255 - 0xff
    "11111111", -- 4038 - 0xfc6  :  255 - 0xff
    "11111111", -- 4039 - 0xfc7  :  255 - 0xff
    "01000000", -- 4040 - 0xfc8  :   64 - 0x40 -- plane 1
    "01000000", -- 4041 - 0xfc9  :   64 - 0x40
    "01000000", -- 4042 - 0xfca  :   64 - 0x40
    "01111111", -- 4043 - 0xfcb  :  127 - 0x7f
    "00000000", -- 4044 - 0xfcc  :    0 - 0x0
    "00000000", -- 4045 - 0xfcd  :    0 - 0x0
    "00000000", -- 4046 - 0xfce  :    0 - 0x0
    "00000000", -- 4047 - 0xfcf  :    0 - 0x0
    "00000000", -- 4048 - 0xfd0  :    0 - 0x0 -- Sprite 0xfd
    "00000000", -- 4049 - 0xfd1  :    0 - 0x0
    "00000000", -- 4050 - 0xfd2  :    0 - 0x0
    "00000000", -- 4051 - 0xfd3  :    0 - 0x0
    "00000000", -- 4052 - 0xfd4  :    0 - 0x0
    "11111111", -- 4053 - 0xfd5  :  255 - 0xff
    "11111111", -- 4054 - 0xfd6  :  255 - 0xff
    "11111111", -- 4055 - 0xfd7  :  255 - 0xff
    "00000000", -- 4056 - 0xfd8  :    0 - 0x0 -- plane 1
    "00000000", -- 4057 - 0xfd9  :    0 - 0x0
    "00000000", -- 4058 - 0xfda  :    0 - 0x0
    "11111111", -- 4059 - 0xfdb  :  255 - 0xff
    "00000000", -- 4060 - 0xfdc  :    0 - 0x0
    "00000000", -- 4061 - 0xfdd  :    0 - 0x0
    "00000000", -- 4062 - 0xfde  :    0 - 0x0
    "00000000", -- 4063 - 0xfdf  :    0 - 0x0
    "00000010", -- 4064 - 0xfe0  :    2 - 0x2 -- Sprite 0xfe
    "00000010", -- 4065 - 0xfe1  :    2 - 0x2
    "00000000", -- 4066 - 0xfe2  :    0 - 0x0
    "00000000", -- 4067 - 0xfe3  :    0 - 0x0
    "00000000", -- 4068 - 0xfe4  :    0 - 0x0
    "11111111", -- 4069 - 0xfe5  :  255 - 0xff
    "11111111", -- 4070 - 0xfe6  :  255 - 0xff
    "11111111", -- 4071 - 0xfe7  :  255 - 0xff
    "00000010", -- 4072 - 0xfe8  :    2 - 0x2 -- plane 1
    "00000010", -- 4073 - 0xfe9  :    2 - 0x2
    "00000010", -- 4074 - 0xfea  :    2 - 0x2
    "11111110", -- 4075 - 0xfeb  :  254 - 0xfe
    "00000000", -- 4076 - 0xfec  :    0 - 0x0
    "00000000", -- 4077 - 0xfed  :    0 - 0x0
    "00000000", -- 4078 - 0xfee  :    0 - 0x0
    "00000000", -- 4079 - 0xfef  :    0 - 0x0
    "11111111", -- 4080 - 0xff0  :  255 - 0xff -- Sprite 0xff
    "11111111", -- 4081 - 0xff1  :  255 - 0xff
    "11111111", -- 4082 - 0xff2  :  255 - 0xff
    "11111111", -- 4083 - 0xff3  :  255 - 0xff
    "11111111", -- 4084 - 0xff4  :  255 - 0xff
    "11111111", -- 4085 - 0xff5  :  255 - 0xff
    "11111111", -- 4086 - 0xff6  :  255 - 0xff
    "11111111", -- 4087 - 0xff7  :  255 - 0xff
    "00000000", -- 4088 - 0xff8  :    0 - 0x0 -- plane 1
    "00000000", -- 4089 - 0xff9  :    0 - 0x0
    "00000000", -- 4090 - 0xffa  :    0 - 0x0
    "00000000", -- 4091 - 0xffb  :    0 - 0x0
    "00000000", -- 4092 - 0xffc  :    0 - 0x0
    "00000000", -- 4093 - 0xffd  :    0 - 0x0
    "00000000", -- 4094 - 0xffe  :    0 - 0x0
    "00000000"  -- 4095 - 0xfff  :    0 - 0x0
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
