--------------------------------------------------------------------------------
-- Felipe Machado Sanchez
-- Departameto de Tecnologia Electronica
-- Universidad Rey Juan Carlos
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package PKG_ROM_IMGS is

  -- constant lab_20b
  -- constant monster_blue
  -- constant monster_red
  -- constant monster_green
  -- constant mario_blue
  -- constant mario_red
  -- constant mario_green
  -- constant pacman_blue
  -- constant pacman_red
  -- constant pacman_green

  type memostruct_2b is array (natural range<>) of std_logic_vector(20-1 downto 0);
  constant lab_20b : memostruct_2b := (
       "11111111100111111111",
       "10000100000000010001",
       "10110101111101010101",
       "10000000010001000101",
       "00101111010111110100",
       "10100000000000100101",
       "10110101100110101101",
       "00000101000010000000",
       "10110101111110111101",
       "10010000000000000001",
       "11010101110110111011",
       "10000100010000100001",
       "10111111011011111101",
       "10000000000000000001",
       "11111111100111111111"
        );

  --signal addr_int  : natural range 0 to 2**10-1;
  type memostruct is array (natural range<>) of std_logic_vector(4-1 downto 0);
  constant monster_blue : memostruct := (
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1100",
       "1011",
       "1011",
       "1100",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "0111",
       "0011",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0011",
       "0111",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "0100",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0100",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1001",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0111",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1000",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0110",
       "1011",
       "1111",
       "1111",
       "1101",
       "0111",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0100",
       "1011",
       "1111",
       "1111",
       "1101",
       "0111",
       "0010",
       "0010",
       "0010",
       "0010",
       "0011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1001",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0100",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1001",
       "0010",
       "0010",
       "0010",
       "0010",
       "1001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0100",
       "0010",
       "0010",
       "0010",
       "0010",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0101",
       "0010",
       "0010",
       "0010",
       "0011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1001",
       "0010",
       "0010",
       "0010",
       "0100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1001",
       "0010",
       "0010",
       "0010",
       "0010",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1100",
       "1011",
       "1011",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "0010",
       "0010",
       "0010",
       "0110",
       "1100",
       "1011",
       "1011",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "0010",
       "0010",
       "0010",
       "0010",
       "0111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1000",
       "1011",
       "1011",
       "1011",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0010",
       "0010",
       "0010",
       "0110",
       "1011",
       "1011",
       "1011",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0010",
       "0010",
       "0010",
       "0010",
       "0100",
       "1111",
       "1111",
       "1111",
       "1111",
       "0110",
       "1011",
       "1011",
       "1011",
       "1011",
       "1110",
       "1111",
       "1111",
       "1111",
       "1100",
       "0010",
       "0010",
       "0010",
       "0101",
       "1011",
       "1011",
       "1011",
       "1011",
       "1110",
       "1111",
       "1111",
       "1111",
       "1101",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1111",
       "1111",
       "1111",
       "1101",
       "0100",
       "1011",
       "1011",
       "1011",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1011",
       "0010",
       "0010",
       "0010",
       "0100",
       "1011",
       "1011",
       "1011",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1011",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1101",
       "1111",
       "1111",
       "1100",
       "0010",
       "1100",
       "1011",
       "1011",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "0111",
       "0010",
       "0010",
       "0010",
       "0010",
       "1100",
       "1011",
       "1011",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "0111",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1011",
       "1111",
       "1111",
       "1010",
       "0010",
       "1000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1010",
       "1111",
       "1111",
       "1001",
       "0010",
       "0010",
       "1001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0011",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0100",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1001",
       "1111",
       "1111",
       "0111",
       "0010",
       "0010",
       "0010",
       "0100",
       "0111",
       "1000",
       "0101",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0100",
       "0111",
       "1000",
       "0101",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0111",
       "1111",
       "1111",
       "0110",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0110",
       "1111",
       "1111",
       "0101",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0101",
       "1111",
       "1111",
       "0100",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0100",
       "1111",
       "1111",
       "0011",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0011",
       "1111",
       "1111",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1111",
       "1111",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1111",
       "1111",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1110",
       "1110",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1110",
       "1101",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "1101",
       "1101",
       "0010",
       "0010",
       "0100",
       "1100",
       "1111",
       "1101",
       "0101",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0111",
       "1110",
       "1110",
       "1000",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0101",
       "1101",
       "1111",
       "1100",
       "0100",
       "0010",
       "0010",
       "1101",
       "1100",
       "0010",
       "0101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0110",
       "0010",
       "0010",
       "0010",
       "0010",
       "1000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1001",
       "0010",
       "0010",
       "0010",
       "0010",
       "0110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0101",
       "0010",
       "1100",
       "1101",
       "0110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1000",
       "0011",
       "0100",
       "1010",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1010",
       "0100",
       "0011",
       "1000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0110",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111"
        );

  constant  monster_green : memostruct := (
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1100",
       "1011",
       "1011",
       "1100",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "0111",
       "0011",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0011",
       "0110",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "0100",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0100",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1000",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0111",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1000",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0101",
       "1011",
       "1111",
       "1111",
       "1101",
       "0111",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0011",
       "1011",
       "1111",
       "1111",
       "1101",
       "0111",
       "0001",
       "0001",
       "0001",
       "0001",
       "0011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0100",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0100",
       "0001",
       "0001",
       "0001",
       "0001",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0100",
       "0001",
       "0001",
       "0001",
       "0011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1111",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1001",
       "0001",
       "0001",
       "0001",
       "0011",
       "1111",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1001",
       "0111",
       "0111",
       "1010",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "0001",
       "0001",
       "0001",
       "0110",
       "1001",
       "0111",
       "0111",
       "1010",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "0001",
       "0001",
       "0001",
       "0001",
       "0111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0111",
       "0111",
       "0111",
       "0111",
       "0111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1101",
       "0001",
       "0001",
       "0001",
       "0101",
       "0111",
       "0111",
       "0111",
       "0111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1101",
       "0001",
       "0001",
       "0001",
       "0001",
       "0011",
       "1111",
       "1111",
       "1111",
       "1111",
       "0100",
       "0111",
       "0111",
       "0111",
       "0111",
       "1101",
       "1111",
       "1111",
       "1111",
       "1100",
       "0001",
       "0001",
       "0001",
       "0011",
       "0111",
       "0111",
       "0111",
       "0111",
       "1101",
       "1111",
       "1111",
       "1111",
       "1100",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1111",
       "1111",
       "1111",
       "1101",
       "0011",
       "0111",
       "0111",
       "0111",
       "0111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1010",
       "0001",
       "0001",
       "0001",
       "0011",
       "0111",
       "0111",
       "0111",
       "0111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1011",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1101",
       "1111",
       "1111",
       "1011",
       "0010",
       "1001",
       "0111",
       "0111",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "0111",
       "0001",
       "0001",
       "0001",
       "0010",
       "1001",
       "0111",
       "0111",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "0111",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1011",
       "1111",
       "1111",
       "1010",
       "0001",
       "1000",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0010",
       "0001",
       "0001",
       "0001",
       "0001",
       "1000",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0010",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1010",
       "1111",
       "1111",
       "1001",
       "0001",
       "0001",
       "1001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0011",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0011",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1000",
       "1111",
       "1111",
       "0111",
       "0001",
       "0001",
       "0001",
       "0011",
       "0111",
       "0111",
       "0101",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0011",
       "0111",
       "0111",
       "0101",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0111",
       "1111",
       "1111",
       "0110",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0110",
       "1111",
       "1111",
       "0101",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0101",
       "1111",
       "1111",
       "0100",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0100",
       "1111",
       "1111",
       "0011",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0011",
       "1111",
       "1111",
       "0010",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0010",
       "1111",
       "1111",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1111",
       "1111",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1110",
       "1110",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1110",
       "1101",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "1101",
       "1101",
       "0001",
       "0001",
       "0011",
       "1011",
       "1111",
       "1101",
       "0101",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0111",
       "1110",
       "1110",
       "0111",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0101",
       "1101",
       "1111",
       "1100",
       "0100",
       "0001",
       "0001",
       "1100",
       "1100",
       "0001",
       "0100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0110",
       "0001",
       "0001",
       "0001",
       "0001",
       "1000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1000",
       "0001",
       "0001",
       "0001",
       "0001",
       "0101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0101",
       "0001",
       "1100",
       "1101",
       "0101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1000",
       "0011",
       "0011",
       "1010",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1010",
       "0011",
       "0011",
       "1000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0110",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111"
        );


  constant monster_red : memostruct := (
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1100",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0100",
       "0000",
       "0000",
       "0110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "0100",
       "0000",
       "0000",
       "0110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1011",
       "0000",
       "0000",
       "0000",
       "0000",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1011",
       "0000",
       "0000",
       "0000",
       "0000",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1001",
       "0000",
       "0000",
       "0000",
       "0000",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1001",
       "0000",
       "0000",
       "0000",
       "0000",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1011",
       "0000",
       "0000",
       "0000",
       "0000",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1011",
       "0000",
       "0000",
       "0000",
       "0000",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "0110",
       "0000",
       "0000",
       "0111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "0110",
       "0000",
       "0000",
       "0111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1111",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111"
        );


  constant mario_blue : memostruct := (
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "1000",
       "0101",
       "1001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1011",
       "0010",
       "0000",
       "0001",
       "0000",
       "1000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0101",
       "0000",
       "0000",
       "0010",
       "0010",
       "0000",
       "0001",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1000",
       "0000",
       "0011",
       "0010",
       "0010",
       "0010",
       "0011",
       "0000",
       "1001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0000",
       "0011",
       "0010",
       "0010",
       "0010",
       "0010",
       "0011",
       "0000",
       "0011",
       "1010",
       "0110",
       "0100",
       "0000",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0001",
       "0000",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0001",
       "0000",
       "0000",
       "0000",
       "0011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1011",
       "0000",
       "0011",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0001",
       "0000",
       "0000",
       "0010",
       "0000",
       "0011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0011",
       "0000",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0001",
       "0010",
       "0101",
       "1001",
       "1000",
       "0111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0000",
       "0010",
       "0010",
       "0001",
       "0000",
       "0010",
       "0000",
       "0110",
       "1100",
       "1011",
       "1111",
       "1010",
       "1111",
       "1111",
       "1100",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0000",
       "0001",
       "0010",
       "0000",
       "0001",
       "0110",
       "0000",
       "0000",
       "0001",
       "1000",
       "1101",
       "1111",
       "1010",
       "1101",
       "1001",
       "1000",
       "1100",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0000",
       "0000",
       "0010",
       "0001",
       "0000",
       "1101",
       "1101",
       "1010",
       "0000",
       "0000",
       "0000",
       "1101",
       "1010",
       "0011",
       "0110",
       "0110",
       "1000",
       "1010",
       "1000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0000",
       "0000",
       "0011",
       "0000",
       "0011",
       "1111",
       "1001",
       "0111",
       "1000",
       "0000",
       "1000",
       "1110",
       "1101",
       "0000",
       "0000",
       "0000",
       "0101",
       "0110",
       "1010",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "0000",
       "0000",
       "0001",
       "0000",
       "1100",
       "1110",
       "1010",
       "1101",
       "1010",
       "1011",
       "1010",
       "1011",
       "1011",
       "0100",
       "0000",
       "0000",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0011",
       "0000",
       "0000",
       "0010",
       "1011",
       "1101",
       "1000",
       "0111",
       "1000",
       "1000",
       "1000",
       "1000",
       "1001",
       "1001",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1010",
       "0010",
       "0000",
       "0000",
       "0000",
       "0001",
       "0101",
       "0101",
       "0110",
       "0111",
       "1000",
       "0111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0010",
       "0000",
       "0001",
       "0011",
       "0100",
       "0011",
       "0001",
       "0010",
       "1010",
       "1111",
       "1111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0000",
       "0011",
       "0010",
       "0011",
       "1100",
       "1110",
       "0010",
       "0011",
       "0000",
       "1011",
       "1110",
       "1111",
       "1110",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1011",
       "1100",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "0000",
       "0010",
       "0010",
       "0001",
       "0000",
       "1111",
       "1110",
       "1111",
       "1010",
       "0111",
       "1110",
       "1111",
       "1100",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1011",
       "1011",
       "1100",
       "1101",
       "1111",
       "1100",
       "1111",
       "1001",
       "0000",
       "0010",
       "0001",
       "0000",
       "0000",
       "1011",
       "0101",
       "0001",
       "1111",
       "1000",
       "1000",
       "1111",
       "1111",
       "1011",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1011",
       "1011",
       "1101",
       "1011",
       "1111",
       "1001",
       "0000",
       "0000",
       "0000",
       "0100",
       "1101",
       "1111",
       "1010",
       "0001",
       "1110",
       "1100",
       "0110",
       "1010",
       "1101",
       "1001",
       "0111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1010",
       "1110",
       "1111",
       "1111",
       "1011",
       "1010",
       "1100",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1101",
       "1111",
       "1111",
       "1001",
       "0000",
       "0000",
       "0100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1101",
       "1111",
       "1010",
       "1010",
       "1011",
       "1100",
       "1100",
       "1100",
       "1101",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "0000",
       "0010",
       "0011",
       "0000",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0000",
       "0000",
       "1000",
       "1100",
       "1001",
       "1010",
       "1100",
       "1011",
       "1100",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1011",
       "0000",
       "0011",
       "0000",
       "0001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1010",
       "0000",
       "0011",
       "1000",
       "1100",
       "1010",
       "1001",
       "1010",
       "1100",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1111",
       "1110",
       "0000",
       "0010",
       "0000",
       "1010",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0100",
       "0000",
       "1000",
       "0110",
       "1010",
       "1100",
       "1010",
       "1010",
       "1010",
       "1010",
       "1011",
       "1100",
       "1100",
       "1101",
       "1101",
       "1110",
       "0000",
       "0000",
       "0000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0011",
       "0000",
       "1010",
       "1001",
       "0110",
       "1001",
       "1010",
       "1011",
       "1011",
       "1010",
       "1001",
       "1010",
       "1010",
       "1011",
       "1101",
       "1101",
       "0000",
       "0000",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "0000",
       "0000",
       "1010",
       "1010",
       "1010",
       "1000",
       "0111",
       "0111",
       "0111",
       "1011",
       "1100",
       "1010",
       "1001",
       "1001",
       "1100",
       "1001",
       "0000",
       "0000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0111",
       "0000",
       "0000",
       "0111",
       "1100",
       "1001",
       "1001",
       "1001",
       "1000",
       "1011",
       "1111",
       "1111",
       "1111",
       "1110",
       "1011",
       "1011",
       "0010",
       "0000",
       "1010",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0001",
       "0000",
       "0001",
       "0001",
       "1010",
       "1100",
       "1100",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1011",
       "0000",
       "0000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "0000",
       "0000",
       "0010",
       "0000",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0101",
       "0000",
       "0000",
       "0110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "0110",
       "0110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111"
        );

  constant  mario_green : memostruct := (
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "1000",
       "0101",
       "1001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1011",
       "0010",
       "0000",
       "0000",
       "0000",
       "1000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0101",
       "0000",
       "0000",
       "0001",
       "0010",
       "0000",
       "0000",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0111",
       "0000",
       "0010",
       "0001",
       "0001",
       "0010",
       "0010",
       "0000",
       "1000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0000",
       "0010",
       "0001",
       "0001",
       "0001",
       "0001",
       "0010",
       "0000",
       "0010",
       "1001",
       "0110",
       "0011",
       "0000",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0001",
       "0000",
       "0001",
       "0001",
       "0001",
       "0001",
       "0010",
       "0010",
       "0001",
       "0000",
       "0000",
       "0000",
       "0000",
       "0011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1011",
       "0000",
       "0010",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0000",
       "0000",
       "0000",
       "0010",
       "0000",
       "0011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0011",
       "0000",
       "0010",
       "0001",
       "0010",
       "0010",
       "0000",
       "0000",
       "0010",
       "0110",
       "1011",
       "1010",
       "0111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0000",
       "0001",
       "0001",
       "0000",
       "0000",
       "0000",
       "0000",
       "1000",
       "1110",
       "1111",
       "1110",
       "1000",
       "1111",
       "1111",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0000",
       "0000",
       "0010",
       "0000",
       "0000",
       "0111",
       "0001",
       "0000",
       "0011",
       "1010",
       "1111",
       "1111",
       "0111",
       "1111",
       "1011",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0000",
       "0000",
       "0010",
       "0000",
       "0000",
       "1111",
       "1111",
       "1101",
       "0000",
       "0000",
       "0001",
       "1111",
       "1110",
       "0011",
       "1000",
       "1000",
       "1010",
       "1100",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0000",
       "0000",
       "0011",
       "0000",
       "0100",
       "1111",
       "1100",
       "1001",
       "1011",
       "0000",
       "1010",
       "1111",
       "1111",
       "0000",
       "0000",
       "0000",
       "0111",
       "1000",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "0000",
       "0000",
       "0001",
       "0000",
       "1111",
       "1111",
       "1110",
       "1111",
       "1101",
       "1110",
       "1101",
       "1111",
       "1110",
       "0101",
       "0000",
       "0000",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0010",
       "0000",
       "0000",
       "0011",
       "1110",
       "1111",
       "1010",
       "1001",
       "1011",
       "1011",
       "1010",
       "1010",
       "1101",
       "1011",
       "1010",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1010",
       "0010",
       "0000",
       "0000",
       "0000",
       "0011",
       "0111",
       "1000",
       "1000",
       "1000",
       "1001",
       "1001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0001",
       "0000",
       "0010",
       "0011",
       "0011",
       "0100",
       "0101",
       "0110",
       "1100",
       "1111",
       "1111",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0000",
       "0010",
       "0000",
       "0000",
       "0100",
       "0101",
       "0000",
       "0000",
       "0000",
       "1011",
       "1101",
       "1111",
       "1110",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1010",
       "1011",
       "1101",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "0000",
       "0010",
       "0010",
       "0010",
       "0001",
       "0101",
       "1100",
       "1001",
       "0010",
       "1100",
       "1100",
       "1111",
       "1011",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1010",
       "1001",
       "1011",
       "1011",
       "1110",
       "1010",
       "1111",
       "1000",
       "0000",
       "0010",
       "0001",
       "0000",
       "0000",
       "0010",
       "1111",
       "1111",
       "1000",
       "0110",
       "1001",
       "1110",
       "1111",
       "1010",
       "1010",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1010",
       "1001",
       "1010",
       "1100",
       "1010",
       "1111",
       "0111",
       "0000",
       "0000",
       "0000",
       "0010",
       "0101",
       "0110",
       "0100",
       "1011",
       "0110",
       "0011",
       "0111",
       "1000",
       "1011",
       "1001",
       "0110",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1010",
       "1000",
       "1101",
       "1111",
       "1111",
       "0001",
       "0100",
       "0101",
       "0110",
       "0110",
       "0110",
       "0101",
       "0011",
       "0011",
       "0110",
       "1111",
       "1111",
       "1010",
       "0110",
       "0110",
       "0111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1111",
       "1110",
       "0001",
       "0100",
       "0100",
       "0101",
       "0101",
       "0101",
       "0101",
       "0110",
       "0110",
       "0101",
       "1100",
       "1101",
       "0101",
       "0111",
       "0111",
       "0000",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0000",
       "0000",
       "0001",
       "0100",
       "0011",
       "0100",
       "0101",
       "0101",
       "0101",
       "0110",
       "0110",
       "0110",
       "0110",
       "0100",
       "0001",
       "0100",
       "0110",
       "0010",
       "0100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1011",
       "0000",
       "0100",
       "0010",
       "0101",
       "0100",
       "0011",
       "0100",
       "0101",
       "0101",
       "0101",
       "0101",
       "0110",
       "0110",
       "0111",
       "0101",
       "0101",
       "0101",
       "0000",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0101",
       "0000",
       "0100",
       "0001",
       "0100",
       "0101",
       "0100",
       "0100",
       "0100",
       "0100",
       "0100",
       "0101",
       "0101",
       "0101",
       "0101",
       "0101",
       "0100",
       "0010",
       "0010",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0100",
       "0001",
       "0100",
       "0011",
       "0010",
       "0011",
       "0100",
       "0100",
       "0101",
       "0010",
       "0010",
       "0011",
       "0100",
       "0101",
       "0101",
       "0101",
       "0100",
       "0000",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "0000",
       "0011",
       "0011",
       "0100",
       "0100",
       "0011",
       "0011",
       "0010",
       "0000",
       "0110",
       "0111",
       "0001",
       "0000",
       "0010",
       "0100",
       "0101",
       "0010",
       "0001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1000",
       "0000",
       "0100",
       "0011",
       "0100",
       "0010",
       "0000",
       "0000",
       "0000",
       "1000",
       "1111",
       "1111",
       "1111",
       "1100",
       "0101",
       "0000",
       "0011",
       "0000",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0011",
       "0001",
       "0101",
       "0011",
       "0000",
       "0110",
       "1001",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1001",
       "0000",
       "0000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0000",
       "0011",
       "0101",
       "0001",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0110",
       "0001",
       "0011",
       "1000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1000",
       "1000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111"
        );


  constant mario_red : memostruct := (
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1011",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "1111",
       "1111",
       "1111",
       "1001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1011",
       "1100",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "0101",
       "1000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1010",
       "1101",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0100",
       "0110",
       "0100",
       "1001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1011",
       "1010",
       "1101",
       "1110",
       "1111",
       "1111",
       "1111",
       "1100",
       "1100",
       "1101",
       "1101",
       "1101",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1010",
       "1010",
       "1100",
       "1101",
       "1101",
       "1101",
       "1010",
       "1101",
       "1111",
       "1111",
       "1110",
       "0110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1001",
       "1010",
       "1010",
       "1001",
       "1001",
       "1011",
       "0110",
       "0101",
       "1010",
       "1101",
       "1111",
       "1111",
       "0100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1010",
       "1010",
       "1010",
       "1001",
       "1000",
       "1111",
       "1111",
       "1110",
       "0101",
       "0011",
       "0111",
       "1111",
       "1111",
       "0011",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1011",
       "1010",
       "1010",
       "1001",
       "1010",
       "1111",
       "1110",
       "1111",
       "1101",
       "0101",
       "1101",
       "1111",
       "1111",
       "0010",
       "0000",
       "0001",
       "1011",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1010",
       "1010",
       "1001",
       "0101",
       "1111",
       "1111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1000",
       "0000",
       "0000",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1011",
       "0101",
       "0100",
       "1000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1010",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1011",
       "0110",
       "0010",
       "0010",
       "0011",
       "1001",
       "1110",
       "1111",
       "1111",
       "1101",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1110",
       "1101",
       "1100",
       "1001",
       "1000",
       "0101",
       "1001",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1011",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1011",
       "0000",
       "0000",
       "1000",
       "0111",
       "1110",
       "1110",
       "1011",
       "1111",
       "1101",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1000",
       "1001",
       "1011",
       "1100",
       "1111",
       "1111",
       "1111",
       "1101",
       "1101",
       "1110",
       "1110",
       "1111",
       "1111",
       "0000",
       "0111",
       "0100",
       "0100",
       "1110",
       "1010",
       "1111",
       "1010",
       "1001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1000",
       "0111",
       "1001",
       "1001",
       "1100",
       "1001",
       "1110",
       "1010",
       "1011",
       "1001",
       "1010",
       "1111",
       "1111",
       "0010",
       "1111",
       "1111",
       "0000",
       "0100",
       "0111",
       "1100",
       "1111",
       "0111",
       "1000",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1001",
       "0111",
       "1000",
       "1011",
       "1001",
       "1110",
       "1001",
       "0101",
       "1010",
       "1111",
       "1101",
       "0100",
       "0000",
       "0001",
       "1101",
       "0010",
       "0000",
       "0111",
       "0101",
       "1000",
       "1000",
       "0110",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1001",
       "0110",
       "1011",
       "1111",
       "1111",
       "0000",
       "0001",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0011",
       "1111",
       "1111",
       "1011",
       "1110",
       "1110",
       "1010",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1111",
       "1110",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0001",
       "0000",
       "0000",
       "1011",
       "1011",
       "1011",
       "1101",
       "1011",
       "0101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0010",
       "0001",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "1010",
       "1011",
       "0110",
       "1001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "0011",
       "0110",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0001",
       "0001",
       "1010",
       "1001",
       "0011",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0111",
       "0101",
       "0011",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0001",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "1001",
       "0101",
       "0101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0110",
       "0110",
       "0001",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0001",
       "0001",
       "0000",
       "0000",
       "1001",
       "0010",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0010",
       "1000",
       "0001",
       "0000",
       "0001",
       "0001",
       "0001",
       "0000",
       "0000",
       "0100",
       "0101",
       "0000",
       "0000",
       "0000",
       "0000",
       "0011",
       "0111",
       "0101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1010",
       "0010",
       "1001",
       "0011",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0111",
       "1111",
       "1111",
       "1111",
       "1011",
       "0011",
       "0000",
       "0110",
       "0010",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0101",
       "0100",
       "1001",
       "0111",
       "0000",
       "0100",
       "1000",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1000",
       "0011",
       "0011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0001",
       "0110",
       "1001",
       "0111",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1000",
       "0110",
       "1000",
       "1010",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1010",
       "1010",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111"
        );

  constant pacman_blue : memostruct := (
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1110",
       "1011",
       "0111",
       "0100",
       "0010",
       "0010",
       "0100",
       "1000",
       "1011",
       "1110",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1011",
       "0101",
       "0010",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0000",
       "0010",
       "0110",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1000",
       "0000",
       "0000",
       "0000",
       "0001",
       "0010",
       "0010",
       "0011",
       "0010",
       "0010",
       "0001",
       "0000",
       "0000",
       "0000",
       "0000",
       "1010",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "0000",
       "0000",
       "0010",
       "0100",
       "0100",
       "0011",
       "0011",
       "0011",
       "0011",
       "0011",
       "0011",
       "0010",
       "0010",
       "0010",
       "0010",
       "0000",
       "0000",
       "0011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1011",
       "0000",
       "0000",
       "0011",
       "0011",
       "0011",
       "0011",
       "0100",
       "0100",
       "0100",
       "0100",
       "0011",
       "0011",
       "0011",
       "0011",
       "0010",
       "0010",
       "0001",
       "0001",
       "0000",
       "0000",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1011",
       "0000",
       "0010",
       "0011",
       "0011",
       "0011",
       "0100",
       "0100",
       "0100",
       "0100",
       "0100",
       "0100",
       "0100",
       "0100",
       "0011",
       "0011",
       "0011",
       "0010",
       "0001",
       "0001",
       "0001",
       "0000",
       "0000",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "0000",
       "0010",
       "0011",
       "0011",
       "0011",
       "0100",
       "0100",
       "0101",
       "0101",
       "0101",
       "0101",
       "0101",
       "0101",
       "0010",
       "0000",
       "0000",
       "0001",
       "0011",
       "0010",
       "0001",
       "0000",
       "0000",
       "0000",
       "0000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0000",
       "0000",
       "0011",
       "0011",
       "0011",
       "0100",
       "0100",
       "0101",
       "0101",
       "0101",
       "0101",
       "0101",
       "0110",
       "0110",
       "0000",
       "0000",
       "0000",
       "0000",
       "0011",
       "0010",
       "0010",
       "0001",
       "0000",
       "0001",
       "0000",
       "0001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1000",
       "0000",
       "0011",
       "0010",
       "0011",
       "0011",
       "0100",
       "0101",
       "0101",
       "0101",
       "0110",
       "0110",
       "0110",
       "0110",
       "0110",
       "0000",
       "0000",
       "0000",
       "0000",
       "0011",
       "0010",
       "0010",
       "0010",
       "0000",
       "0000",
       "0101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0000",
       "0000",
       "0010",
       "0011",
       "0011",
       "0100",
       "0100",
       "0101",
       "0101",
       "0110",
       "0110",
       "0111",
       "0111",
       "0110",
       "0110",
       "0101",
       "0001",
       "0001",
       "0011",
       "0011",
       "0011",
       "0010",
       "0000",
       "0000",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1010",
       "0000",
       "0010",
       "0010",
       "0011",
       "0011",
       "0100",
       "0100",
       "0101",
       "0101",
       "0110",
       "0111",
       "1000",
       "0111",
       "0110",
       "0110",
       "0110",
       "0110",
       "0101",
       "0100",
       "0100",
       "0000",
       "0000",
       "1000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0100",
       "0000",
       "0010",
       "0010",
       "0011",
       "0011",
       "0100",
       "0100",
       "0101",
       "0110",
       "0110",
       "0111",
       "0111",
       "0111",
       "0111",
       "0110",
       "0101",
       "0101",
       "0101",
       "0011",
       "0000",
       "0011",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1011",
       "0000",
       "0000",
       "0010",
       "0010",
       "0011",
       "0011",
       "0100",
       "0100",
       "0101",
       "0101",
       "0110",
       "0110",
       "0111",
       "0111",
       "0110",
       "0110",
       "0101",
       "0101",
       "0001",
       "0001",
       "1010",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0111",
       "0000",
       "0000",
       "0001",
       "0010",
       "0010",
       "0011",
       "0011",
       "0100",
       "0101",
       "0101",
       "0101",
       "0110",
       "0110",
       "0110",
       "0110",
       "0110",
       "0011",
       "0000",
       "0111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0011",
       "0000",
       "0000",
       "0001",
       "0010",
       "0010",
       "0011",
       "0011",
       "0011",
       "0100",
       "0101",
       "0101",
       "0101",
       "0101",
       "0101",
       "0101",
       "0001",
       "0011",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0000",
       "0000",
       "0000",
       "0001",
       "0001",
       "0010",
       "0010",
       "0011",
       "0011",
       "0100",
       "0100",
       "0101",
       "0101",
       "0101",
       "0101",
       "0011",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0000",
       "0000",
       "0000",
       "0000",
       "0001",
       "0010",
       "0010",
       "0010",
       "0011",
       "0011",
       "0100",
       "0100",
       "0100",
       "0100",
       "0100",
       "0011",
       "1010",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0100",
       "0000",
       "0000",
       "0000",
       "0001",
       "0001",
       "0010",
       "0010",
       "0011",
       "0011",
       "0011",
       "0011",
       "0011",
       "0011",
       "0011",
       "0011",
       "0000",
       "0001",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0111",
       "0000",
       "0000",
       "0000",
       "0000",
       "0001",
       "0001",
       "0010",
       "0010",
       "0010",
       "0011",
       "0011",
       "0011",
       "0011",
       "0011",
       "0011",
       "0011",
       "0010",
       "0000",
       "0101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0001",
       "0001",
       "0001",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0000",
       "0000",
       "1001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0100",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0001",
       "0001",
       "0001",
       "0001",
       "0010",
       "0010",
       "0010",
       "0010",
       "0010",
       "0001",
       "0001",
       "0010",
       "0000",
       "0000",
       "0010",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1010",
       "0000",
       "0001",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0001",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1000",
       "0000",
       "0001",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0011",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0001",
       "0000",
       "0001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "0000",
       "0000",
       "0001",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "0001",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0001",
       "0000",
       "0000",
       "0000",
       "0100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1010",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "0110",
       "0010",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0000",
       "0011",
       "0111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "0111",
       "0011",
       "0000",
       "0000",
       "0100",
       "0111",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110"
        );

  constant  pacman_green : memostruct := (
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1101",
       "1100",
       "1100",
       "1100",
       "1100",
       "1101",
       "1110",
       "1110",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1100",
       "1100",
       "1100",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1100",
       "1100",
       "1100",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1100",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1100",
       "1101",
       "1101",
       "1100",
       "1011",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1100",
       "1100",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1110",
       "1110",
       "1101",
       "1101",
       "1101",
       "1101",
       "1100",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1100",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1110",
       "1111",
       "1100",
       "1100",
       "1111",
       "1101",
       "1101",
       "1101",
       "1100",
       "1100",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1111",
       "0110",
       "0000",
       "0000",
       "0110",
       "1111",
       "1101",
       "1101",
       "1101",
       "1101",
       "1100",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1100",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1110",
       "1101",
       "1110",
       "1111",
       "0000",
       "0000",
       "0000",
       "0000",
       "1110",
       "1101",
       "1101",
       "1100",
       "1100",
       "1101",
       "1010",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "1100",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1110",
       "1101",
       "1110",
       "1110",
       "1110",
       "1111",
       "0000",
       "0000",
       "0000",
       "0000",
       "1111",
       "1101",
       "1101",
       "1101",
       "1100",
       "1011",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1110",
       "1110",
       "1110",
       "1110",
       "1101",
       "1111",
       "1101",
       "0100",
       "0100",
       "1101",
       "1111",
       "1101",
       "1101",
       "1100",
       "1100",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1100",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "1100",
       "1100",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "1100",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1100",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1100",
       "1100",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1110",
       "1110",
       "1110",
       "1110",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "1100",
       "1100",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1110",
       "1110",
       "1101",
       "1110",
       "1101",
       "1101",
       "1101",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "1100",
       "1100",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1100",
       "1100",
       "1100",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1100",
       "1100",
       "1100",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1100",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "1011",
       "1100",
       "1100",
       "1100",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1100",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1011",
       "1011",
       "1100",
       "1100",
       "1100",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1100",
       "1100",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1011",
       "1100",
       "1100",
       "1100",
       "1100",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1100",
       "1100",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "1010",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1100",
       "1101",
       "1100",
       "1100",
       "1100",
       "1100",
       "1011",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1001",
       "1011",
       "1011",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1101",
       "1100",
       "1100",
       "1100",
       "1100",
       "1011",
       "1010",
       "1010",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1001",
       "1011",
       "1011",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1011",
       "1011",
       "1011",
       "1010",
       "1000",
       "1010",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1001",
       "1010",
       "1011",
       "1011",
       "1011",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1011",
       "1011",
       "1011",
       "1010",
       "1010",
       "1010",
       "1010",
       "0110",
       "1001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1000",
       "1010",
       "1011",
       "1011",
       "1011",
       "1011",
       "1011",
       "1011",
       "1100",
       "1100",
       "1100",
       "1011",
       "1100",
       "1011",
       "1011",
       "1011",
       "1011",
       "1011",
       "1010",
       "1010",
       "1010",
       "1010",
       "1000",
       "0111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1000",
       "1010",
       "1011",
       "1011",
       "1011",
       "1011",
       "1011",
       "1011",
       "1011",
       "1011",
       "1011",
       "1011",
       "1011",
       "1011",
       "1010",
       "1010",
       "1010",
       "1010",
       "1010",
       "1010",
       "1000",
       "0111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1000",
       "1001",
       "1010",
       "1010",
       "1010",
       "1010",
       "1011",
       "1011",
       "1011",
       "1011",
       "1010",
       "1010",
       "1010",
       "1010",
       "1010",
       "1010",
       "1010",
       "1001",
       "0111",
       "0111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1001",
       "1000",
       "1001",
       "1010",
       "1010",
       "1010",
       "1010",
       "1010",
       "1010",
       "1010",
       "1010",
       "1010",
       "1010",
       "1010",
       "1001",
       "1000",
       "0110",
       "1001",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1000",
       "0111",
       "1000",
       "1001",
       "1001",
       "1010",
       "1010",
       "1010",
       "1001",
       "1001",
       "1000",
       "0111",
       "0110",
       "1000",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1011",
       "1001",
       "1001",
       "1001",
       "1001",
       "1001",
       "1001",
       "1001",
       "1001",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1010",
       "1000",
       "0111",
       "0111",
       "1000",
       "1010",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110"
        );


  constant pacman_red : memostruct := (
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0111",
       "0000",
       "0000",
       "0111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0000",
       "0000",
       "0000",
       "0000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0000",
       "0000",
       "0000",
       "0000",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "0100",
       "0101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1101",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1101",
       "1100",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1101",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1101",
       "1101",
       "1101",
       "1100",
       "1010",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1101",
       "1101",
       "1110",
       "1110",
       "1110",
       "1110",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1101",
       "1101",
       "1101",
       "1100",
       "1100",
       "1011",
       "1010",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1011",
       "1101",
       "1101",
       "1101",
       "1101",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1110",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1100",
       "1100",
       "1011",
       "1010",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1011",
       "1100",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1100",
       "1100",
       "1100",
       "1100",
       "1010",
       "1010",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1100",
       "1011",
       "1100",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1101",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1011",
       "1001",
       "1011",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "1011",
       "1010",
       "1011",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1100",
       "1011",
       "1010",
       "1001",
       "1010",
       "1101",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110",
       "1101",
       "1100",
       "1011",
       "1100",
       "1100",
       "1011",
       "1011",
       "1011",
       "1011",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1101",
       "1011",
       "1010",
       "1001",
       "1001",
       "1010",
       "1011",
       "1100",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1111",
       "1110"
        );



end PKG_ROM_IMGS;

