//-   Background Pattern table COLOR PLANE 0
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
//- Autcmatically generated verilog ROM from a NES memory file----


//-  Original memory dump file name: nova_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_PTABLE_NOVA_BG_PLN0
  (
     input     clk,   // clock
     input      [11-1:0] addr,  //2048 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Background pattern Table COLOR PLANE 0
      11'h0: dout <= 8'b00000000; //    0 :   0 - 0x0 -- Background 0x0
      11'h1: dout <= 8'b00001111; //    1 :  15 - 0xf
      11'h2: dout <= 8'b00000100; //    2 :   4 - 0x4
      11'h3: dout <= 8'b00000011; //    3 :   3 - 0x3
      11'h4: dout <= 8'b00000011; //    4 :   3 - 0x3
      11'h5: dout <= 8'b00000011; //    5 :   3 - 0x3
      11'h6: dout <= 8'b00000100; //    6 :   4 - 0x4
      11'h7: dout <= 8'b00111010; //    7 :  58 - 0x3a
      11'h8: dout <= 8'b00000000; //    8 :   0 - 0x0 -- Background 0x1
      11'h9: dout <= 8'b00111000; //    9 :  56 - 0x38
      11'hA: dout <= 8'b11000110; //   10 : 198 - 0xc6
      11'hB: dout <= 8'b11001011; //   11 : 203 - 0xcb
      11'hC: dout <= 8'b11011100; //   12 : 220 - 0xdc
      11'hD: dout <= 8'b00111010; //   13 :  58 - 0x3a
      11'hE: dout <= 8'b10011010; //   14 : 154 - 0x9a
      11'hF: dout <= 8'b10000001; //   15 : 129 - 0x81
      11'h10: dout <= 8'b01000101; //   16 :  69 - 0x45 -- Background 0x2
      11'h11: dout <= 8'b10000111; //   17 : 135 - 0x87
      11'h12: dout <= 8'b10000011; //   18 : 131 - 0x83
      11'h13: dout <= 8'b10000001; //   19 : 129 - 0x81
      11'h14: dout <= 8'b10000001; //   20 : 129 - 0x81
      11'h15: dout <= 8'b10000001; //   21 : 129 - 0x81
      11'h16: dout <= 8'b01000001; //   22 :  65 - 0x41
      11'h17: dout <= 8'b00100001; //   23 :  33 - 0x21
      11'h18: dout <= 8'b01111111; //   24 : 127 - 0x7f -- Background 0x3
      11'h19: dout <= 8'b01111110; //   25 : 126 - 0x7e
      11'h1A: dout <= 8'b11111100; //   26 : 252 - 0xfc
      11'h1B: dout <= 8'b00111000; //   27 :  56 - 0x38
      11'h1C: dout <= 8'b00011000; //   28 :  24 - 0x18
      11'h1D: dout <= 8'b10001100; //   29 : 140 - 0x8c
      11'h1E: dout <= 8'b11000100; //   30 : 196 - 0xc4
      11'h1F: dout <= 8'b11111100; //   31 : 252 - 0xfc
      11'h20: dout <= 8'b00100011; //   32 :  35 - 0x23 -- Background 0x4
      11'h21: dout <= 8'b00100011; //   33 :  35 - 0x23
      11'h22: dout <= 8'b00100001; //   34 :  33 - 0x21
      11'h23: dout <= 8'b00100000; //   35 :  32 - 0x20
      11'h24: dout <= 8'b00010011; //   36 :  19 - 0x13
      11'h25: dout <= 8'b00001100; //   37 :  12 - 0xc
      11'h26: dout <= 8'b00000000; //   38 :   0 - 0x0
      11'h27: dout <= 8'b00000000; //   39 :   0 - 0x0
      11'h28: dout <= 8'b11111100; //   40 : 252 - 0xfc -- Background 0x5
      11'h29: dout <= 8'b11111100; //   41 : 252 - 0xfc
      11'h2A: dout <= 8'b11111100; //   42 : 252 - 0xfc
      11'h2B: dout <= 8'b11111100; //   43 : 252 - 0xfc
      11'h2C: dout <= 8'b10010000; //   44 : 144 - 0x90
      11'h2D: dout <= 8'b10010000; //   45 : 144 - 0x90
      11'h2E: dout <= 8'b10001000; //   46 : 136 - 0x88
      11'h2F: dout <= 8'b11111000; //   47 : 248 - 0xf8
      11'h30: dout <= 8'b00100011; //   48 :  35 - 0x23 -- Background 0x6
      11'h31: dout <= 8'b00100011; //   49 :  35 - 0x23
      11'h32: dout <= 8'b00100001; //   50 :  33 - 0x21
      11'h33: dout <= 8'b00100000; //   51 :  32 - 0x20
      11'h34: dout <= 8'b00010011; //   52 :  19 - 0x13
      11'h35: dout <= 8'b00001101; //   53 :  13 - 0xd
      11'h36: dout <= 8'b00000010; //   54 :   2 - 0x2
      11'h37: dout <= 8'b00000001; //   55 :   1 - 0x1
      11'h38: dout <= 8'b11111100; //   56 : 252 - 0xfc -- Background 0x7
      11'h39: dout <= 8'b11111100; //   57 : 252 - 0xfc
      11'h3A: dout <= 8'b11111100; //   58 : 252 - 0xfc
      11'h3B: dout <= 8'b11111100; //   59 : 252 - 0xfc
      11'h3C: dout <= 8'b10100100; //   60 : 164 - 0xa4
      11'h3D: dout <= 8'b00100100; //   61 :  36 - 0x24
      11'h3E: dout <= 8'b01010010; //   62 :  82 - 0x52
      11'h3F: dout <= 8'b11101110; //   63 : 238 - 0xee
      11'h40: dout <= 8'b00100011; //   64 :  35 - 0x23 -- Background 0x8
      11'h41: dout <= 8'b00100011; //   65 :  35 - 0x23
      11'h42: dout <= 8'b00100001; //   66 :  33 - 0x21
      11'h43: dout <= 8'b00100000; //   67 :  32 - 0x20
      11'h44: dout <= 8'b00010011; //   68 :  19 - 0x13
      11'h45: dout <= 8'b00001101; //   69 :  13 - 0xd
      11'h46: dout <= 8'b00000001; //   70 :   1 - 0x1
      11'h47: dout <= 8'b00000001; //   71 :   1 - 0x1
      11'h48: dout <= 8'b11111110; //   72 : 254 - 0xfe -- Background 0x9
      11'h49: dout <= 8'b11111110; //   73 : 254 - 0xfe
      11'h4A: dout <= 8'b11111110; //   74 : 254 - 0xfe
      11'h4B: dout <= 8'b11111111; //   75 : 255 - 0xff
      11'h4C: dout <= 8'b10010001; //   76 : 145 - 0x91
      11'h4D: dout <= 8'b00101111; //   77 :  47 - 0x2f
      11'h4E: dout <= 8'b01000000; //   78 :  64 - 0x40
      11'h4F: dout <= 8'b11100000; //   79 : 224 - 0xe0
      11'h50: dout <= 8'b00100011; //   80 :  35 - 0x23 -- Background 0xa
      11'h51: dout <= 8'b00100011; //   81 :  35 - 0x23
      11'h52: dout <= 8'b00100001; //   82 :  33 - 0x21
      11'h53: dout <= 8'b00100000; //   83 :  32 - 0x20
      11'h54: dout <= 8'b00010011; //   84 :  19 - 0x13
      11'h55: dout <= 8'b00001110; //   85 :  14 - 0xe
      11'h56: dout <= 8'b00000001; //   86 :   1 - 0x1
      11'h57: dout <= 8'b00000000; //   87 :   0 - 0x0
      11'h58: dout <= 8'b11111110; //   88 : 254 - 0xfe -- Background 0xb
      11'h59: dout <= 8'b11111110; //   89 : 254 - 0xfe
      11'h5A: dout <= 8'b11111110; //   90 : 254 - 0xfe
      11'h5B: dout <= 8'b11111100; //   91 : 252 - 0xfc
      11'h5C: dout <= 8'b00100100; //   92 :  36 - 0x24
      11'h5D: dout <= 8'b00100010; //   93 :  34 - 0x22
      11'h5E: dout <= 8'b11010010; //   94 : 210 - 0xd2
      11'h5F: dout <= 8'b00001111; //   95 :  15 - 0xf
      11'h60: dout <= 8'b01111111; //   96 : 127 - 0x7f -- Background 0xc
      11'h61: dout <= 8'b01111110; //   97 : 126 - 0x7e
      11'h62: dout <= 8'b11111100; //   98 : 252 - 0xfc
      11'h63: dout <= 8'b00000010; //   99 :   2 - 0x2
      11'h64: dout <= 8'b00000100; //  100 :   4 - 0x4
      11'h65: dout <= 8'b11111100; //  101 : 252 - 0xfc
      11'h66: dout <= 8'b11111100; //  102 : 252 - 0xfc
      11'h67: dout <= 8'b11111110; //  103 : 254 - 0xfe
      11'h68: dout <= 8'b01000101; //  104 :  69 - 0x45 -- Background 0xd
      11'h69: dout <= 8'b10000111; //  105 : 135 - 0x87
      11'h6A: dout <= 8'b10000011; //  106 : 131 - 0x83
      11'h6B: dout <= 8'b10000010; //  107 : 130 - 0x82
      11'h6C: dout <= 8'b10000010; //  108 : 130 - 0x82
      11'h6D: dout <= 8'b10000100; //  109 : 132 - 0x84
      11'h6E: dout <= 8'b01000100; //  110 :  68 - 0x44
      11'h6F: dout <= 8'b00100100; //  111 :  36 - 0x24
      11'h70: dout <= 8'b01111111; //  112 : 127 - 0x7f -- Background 0xe
      11'h71: dout <= 8'b01111110; //  113 : 126 - 0x7e
      11'h72: dout <= 8'b11111100; //  114 : 252 - 0xfc
      11'h73: dout <= 8'b11111000; //  115 : 248 - 0xf8
      11'h74: dout <= 8'b01111000; //  116 : 120 - 0x78
      11'h75: dout <= 8'b01111100; //  117 : 124 - 0x7c
      11'h76: dout <= 8'b11111100; //  118 : 252 - 0xfc
      11'h77: dout <= 8'b11111110; //  119 : 254 - 0xfe
      11'h78: dout <= 8'b00000000; //  120 :   0 - 0x0 -- Background 0xf
      11'h79: dout <= 8'b00001111; //  121 :  15 - 0xf
      11'h7A: dout <= 8'b00000100; //  122 :   4 - 0x4
      11'h7B: dout <= 8'b00000011; //  123 :   3 - 0x3
      11'h7C: dout <= 8'b00000011; //  124 :   3 - 0x3
      11'h7D: dout <= 8'b00000011; //  125 :   3 - 0x3
      11'h7E: dout <= 8'b00000100; //  126 :   4 - 0x4
      11'h7F: dout <= 8'b00000010; //  127 :   2 - 0x2
      11'h80: dout <= 8'b00000111; //  128 :   7 - 0x7 -- Background 0x10
      11'h81: dout <= 8'b00001100; //  129 :  12 - 0xc
      11'h82: dout <= 8'b00010000; //  130 :  16 - 0x10
      11'h83: dout <= 8'b00010000; //  131 :  16 - 0x10
      11'h84: dout <= 8'b00010000; //  132 :  16 - 0x10
      11'h85: dout <= 8'b00100000; //  133 :  32 - 0x20
      11'h86: dout <= 8'b00100000; //  134 :  32 - 0x20
      11'h87: dout <= 8'b00100001; //  135 :  33 - 0x21
      11'h88: dout <= 8'b11111111; //  136 : 255 - 0xff -- Background 0x11
      11'h89: dout <= 8'b01111110; //  137 : 126 - 0x7e
      11'h8A: dout <= 8'b01111100; //  138 : 124 - 0x7c
      11'h8B: dout <= 8'b01111000; //  139 : 120 - 0x78
      11'h8C: dout <= 8'b01011000; //  140 :  88 - 0x58
      11'h8D: dout <= 8'b10001100; //  141 : 140 - 0x8c
      11'h8E: dout <= 8'b11000100; //  142 : 196 - 0xc4
      11'h8F: dout <= 8'b11111100; //  143 : 252 - 0xfc
      11'h90: dout <= 8'b00100011; //  144 :  35 - 0x23 -- Background 0x12
      11'h91: dout <= 8'b00100011; //  145 :  35 - 0x23
      11'h92: dout <= 8'b00100001; //  146 :  33 - 0x21
      11'h93: dout <= 8'b00100000; //  147 :  32 - 0x20
      11'h94: dout <= 8'b00010011; //  148 :  19 - 0x13
      11'h95: dout <= 8'b00001100; //  149 :  12 - 0xc
      11'h96: dout <= 8'b00000000; //  150 :   0 - 0x0
      11'h97: dout <= 8'b00000000; //  151 :   0 - 0x0
      11'h98: dout <= 8'b00000001; //  152 :   1 - 0x1 -- Background 0x13
      11'h99: dout <= 8'b00000001; //  153 :   1 - 0x1
      11'h9A: dout <= 8'b00000011; //  154 :   3 - 0x3
      11'h9B: dout <= 8'b00000100; //  155 :   4 - 0x4
      11'h9C: dout <= 8'b00001000; //  156 :   8 - 0x8
      11'h9D: dout <= 8'b00010000; //  157 :  16 - 0x10
      11'h9E: dout <= 8'b00010000; //  158 :  16 - 0x10
      11'h9F: dout <= 8'b00100000; //  159 :  32 - 0x20
      11'hA0: dout <= 8'b01111111; //  160 : 127 - 0x7f -- Background 0x14
      11'hA1: dout <= 8'b11111110; //  161 : 254 - 0xfe
      11'hA2: dout <= 8'b00000110; //  162 :   6 - 0x6
      11'hA3: dout <= 8'b00000001; //  163 :   1 - 0x1
      11'hA4: dout <= 8'b00000001; //  164 :   1 - 0x1
      11'hA5: dout <= 8'b00000001; //  165 :   1 - 0x1
      11'hA6: dout <= 8'b00000111; //  166 :   7 - 0x7
      11'hA7: dout <= 8'b11111110; //  167 : 254 - 0xfe
      11'hA8: dout <= 8'b00000101; //  168 :   5 - 0x5 -- Background 0x15
      11'hA9: dout <= 8'b00000101; //  169 :   5 - 0x5
      11'hAA: dout <= 8'b00000111; //  170 :   7 - 0x7
      11'hAB: dout <= 8'b00000100; //  171 :   4 - 0x4
      11'hAC: dout <= 8'b00000100; //  172 :   4 - 0x4
      11'hAD: dout <= 8'b00001111; //  173 :  15 - 0xf
      11'hAE: dout <= 8'b00110000; //  174 :  48 - 0x30
      11'hAF: dout <= 8'b01000000; //  175 :  64 - 0x40
      11'hB0: dout <= 8'b11111100; //  176 : 252 - 0xfc -- Background 0x16
      11'hB1: dout <= 8'b11111000; //  177 : 248 - 0xf8
      11'hB2: dout <= 8'b11110000; //  178 : 240 - 0xf0
      11'hB3: dout <= 8'b11100000; //  179 : 224 - 0xe0
      11'hB4: dout <= 8'b01100000; //  180 :  96 - 0x60
      11'hB5: dout <= 8'b11110000; //  181 : 240 - 0xf0
      11'hB6: dout <= 8'b00011100; //  182 :  28 - 0x1c
      11'hB7: dout <= 8'b00000010; //  183 :   2 - 0x2
      11'hB8: dout <= 8'b10000000; //  184 : 128 - 0x80 -- Background 0x17
      11'hB9: dout <= 8'b10000000; //  185 : 128 - 0x80
      11'hBA: dout <= 8'b10000000; //  186 : 128 - 0x80
      11'hBB: dout <= 8'b10000011; //  187 : 131 - 0x83
      11'hBC: dout <= 8'b01001111; //  188 :  79 - 0x4f
      11'hBD: dout <= 8'b00110010; //  189 :  50 - 0x32
      11'hBE: dout <= 8'b00000010; //  190 :   2 - 0x2
      11'hBF: dout <= 8'b00000011; //  191 :   3 - 0x3
      11'hC0: dout <= 8'b00000010; //  192 :   2 - 0x2 -- Background 0x18
      11'hC1: dout <= 8'b00000001; //  193 :   1 - 0x1
      11'hC2: dout <= 8'b00000010; //  194 :   2 - 0x2
      11'hC3: dout <= 8'b11111100; //  195 : 252 - 0xfc
      11'hC4: dout <= 8'b11000000; //  196 : 192 - 0xc0
      11'hC5: dout <= 8'b01000000; //  197 :  64 - 0x40
      11'hC6: dout <= 8'b00100000; //  198 :  32 - 0x20
      11'hC7: dout <= 8'b11100000; //  199 : 224 - 0xe0
      11'hC8: dout <= 8'b00001011; //  200 :  11 - 0xb -- Background 0x19
      11'hC9: dout <= 8'b00001011; //  201 :  11 - 0xb
      11'hCA: dout <= 8'b00001111; //  202 :  15 - 0xf
      11'hCB: dout <= 8'b00001001; //  203 :   9 - 0x9
      11'hCC: dout <= 8'b00001000; //  204 :   8 - 0x8
      11'hCD: dout <= 8'b00001001; //  205 :   9 - 0x9
      11'hCE: dout <= 8'b00001111; //  206 :  15 - 0xf
      11'hCF: dout <= 8'b00110000; //  207 :  48 - 0x30
      11'hD0: dout <= 8'b11111000; //  208 : 248 - 0xf8 -- Background 0x1a
      11'hD1: dout <= 8'b11110000; //  209 : 240 - 0xf0
      11'hD2: dout <= 8'b11100000; //  210 : 224 - 0xe0
      11'hD3: dout <= 8'b11000000; //  211 : 192 - 0xc0
      11'hD4: dout <= 8'b11000000; //  212 : 192 - 0xc0
      11'hD5: dout <= 8'b11000000; //  213 : 192 - 0xc0
      11'hD6: dout <= 8'b11111000; //  214 : 248 - 0xf8
      11'hD7: dout <= 8'b00011111; //  215 :  31 - 0x1f
      11'hD8: dout <= 8'b01000000; //  216 :  64 - 0x40 -- Background 0x1b
      11'hD9: dout <= 8'b01000000; //  217 :  64 - 0x40
      11'hDA: dout <= 8'b10000000; //  218 : 128 - 0x80
      11'hDB: dout <= 8'b10000000; //  219 : 128 - 0x80
      11'hDC: dout <= 8'b01000000; //  220 :  64 - 0x40
      11'hDD: dout <= 8'b00111111; //  221 :  63 - 0x3f
      11'hDE: dout <= 8'b00000100; //  222 :   4 - 0x4
      11'hDF: dout <= 8'b00000111; //  223 :   7 - 0x7
      11'hE0: dout <= 8'b00000000; //  224 :   0 - 0x0 -- Background 0x1c
      11'hE1: dout <= 8'b00000000; //  225 :   0 - 0x0
      11'hE2: dout <= 8'b00000000; //  226 :   0 - 0x0
      11'hE3: dout <= 8'b00000000; //  227 :   0 - 0x0
      11'hE4: dout <= 8'b00000000; //  228 :   0 - 0x0
      11'hE5: dout <= 8'b11111111; //  229 : 255 - 0xff
      11'hE6: dout <= 8'b01000000; //  230 :  64 - 0x40
      11'hE7: dout <= 8'b11000000; //  231 : 192 - 0xc0
      11'hE8: dout <= 8'b11000000; //  232 : 192 - 0xc0 -- Background 0x1d
      11'hE9: dout <= 8'b00100000; //  233 :  32 - 0x20
      11'hEA: dout <= 8'b00100000; //  234 :  32 - 0x20
      11'hEB: dout <= 8'b00100000; //  235 :  32 - 0x20
      11'hEC: dout <= 8'b01000000; //  236 :  64 - 0x40
      11'hED: dout <= 8'b10000000; //  237 : 128 - 0x80
      11'hEE: dout <= 8'b00000000; //  238 :   0 - 0x0
      11'hEF: dout <= 8'b00000000; //  239 :   0 - 0x0
      11'hF0: dout <= 8'b01111111; //  240 : 127 - 0x7f -- Background 0x1e
      11'hF1: dout <= 8'b01100010; //  241 :  98 - 0x62
      11'hF2: dout <= 8'b11000100; //  242 : 196 - 0xc4
      11'hF3: dout <= 8'b00011000; //  243 :  24 - 0x18
      11'hF4: dout <= 8'b00111100; //  244 :  60 - 0x3c
      11'hF5: dout <= 8'b11111110; //  245 : 254 - 0xfe
      11'hF6: dout <= 8'b11111110; //  246 : 254 - 0xfe
      11'hF7: dout <= 8'b11111110; //  247 : 254 - 0xfe
      11'hF8: dout <= 8'b00000000; //  248 :   0 - 0x0 -- Background 0x1f
      11'hF9: dout <= 8'b00111000; //  249 :  56 - 0x38
      11'hFA: dout <= 8'b11000110; //  250 : 198 - 0xc6
      11'hFB: dout <= 8'b11001011; //  251 : 203 - 0xcb
      11'hFC: dout <= 8'b11011100; //  252 : 220 - 0xdc
      11'hFD: dout <= 8'b00111010; //  253 :  58 - 0x3a
      11'hFE: dout <= 8'b10011010; //  254 : 154 - 0x9a
      11'hFF: dout <= 8'b11100001; //  255 : 225 - 0xe1
      11'h100: dout <= 8'b00000000; //  256 :   0 - 0x0 -- Background 0x20
      11'h101: dout <= 8'b00011100; //  257 :  28 - 0x1c
      11'h102: dout <= 8'b00010011; //  258 :  19 - 0x13
      11'h103: dout <= 8'b00001000; //  259 :   8 - 0x8
      11'h104: dout <= 8'b00010000; //  260 :  16 - 0x10
      11'h105: dout <= 8'b00001000; //  261 :   8 - 0x8
      11'h106: dout <= 8'b00010000; //  262 :  16 - 0x10
      11'h107: dout <= 8'b00010000; //  263 :  16 - 0x10
      11'h108: dout <= 8'b00000000; //  264 :   0 - 0x0 -- Background 0x21
      11'h109: dout <= 8'b00111000; //  265 :  56 - 0x38
      11'h10A: dout <= 8'b11001000; //  266 : 200 - 0xc8
      11'h10B: dout <= 8'b00010000; //  267 :  16 - 0x10
      11'h10C: dout <= 8'b00001000; //  268 :   8 - 0x8
      11'h10D: dout <= 8'b00010000; //  269 :  16 - 0x10
      11'h10E: dout <= 8'b00001000; //  270 :   8 - 0x8
      11'h10F: dout <= 8'b00001000; //  271 :   8 - 0x8
      11'h110: dout <= 8'b00001000; //  272 :   8 - 0x8 -- Background 0x22
      11'h111: dout <= 8'b00011100; //  273 :  28 - 0x1c
      11'h112: dout <= 8'b00100111; //  274 :  39 - 0x27
      11'h113: dout <= 8'b00101111; //  275 :  47 - 0x2f
      11'h114: dout <= 8'b00011111; //  276 :  31 - 0x1f
      11'h115: dout <= 8'b00001111; //  277 :  15 - 0xf
      11'h116: dout <= 8'b00001111; //  278 :  15 - 0xf
      11'h117: dout <= 8'b00001111; //  279 :  15 - 0xf
      11'h118: dout <= 8'b00010000; //  280 :  16 - 0x10 -- Background 0x23
      11'h119: dout <= 8'b00111100; //  281 :  60 - 0x3c
      11'h11A: dout <= 8'b11000010; //  282 : 194 - 0xc2
      11'h11B: dout <= 8'b10000010; //  283 : 130 - 0x82
      11'h11C: dout <= 8'b10000010; //  284 : 130 - 0x82
      11'h11D: dout <= 8'b10000010; //  285 : 130 - 0x82
      11'h11E: dout <= 8'b00010010; //  286 :  18 - 0x12
      11'h11F: dout <= 8'b00011100; //  287 :  28 - 0x1c
      11'h120: dout <= 8'b00001111; //  288 :  15 - 0xf -- Background 0x24
      11'h121: dout <= 8'b00001110; //  289 :  14 - 0xe
      11'h122: dout <= 8'b00010100; //  290 :  20 - 0x14
      11'h123: dout <= 8'b00010100; //  291 :  20 - 0x14
      11'h124: dout <= 8'b00010010; //  292 :  18 - 0x12
      11'h125: dout <= 8'b00100101; //  293 :  37 - 0x25
      11'h126: dout <= 8'b01000100; //  294 :  68 - 0x44
      11'h127: dout <= 8'b00111000; //  295 :  56 - 0x38
      11'h128: dout <= 8'b00010000; //  296 :  16 - 0x10 -- Background 0x25
      11'h129: dout <= 8'b00010000; //  297 :  16 - 0x10
      11'h12A: dout <= 8'b00010000; //  298 :  16 - 0x10
      11'h12B: dout <= 8'b00101100; //  299 :  44 - 0x2c
      11'h12C: dout <= 8'b01000100; //  300 :  68 - 0x44
      11'h12D: dout <= 8'b11000100; //  301 : 196 - 0xc4
      11'h12E: dout <= 8'b00111000; //  302 :  56 - 0x38
      11'h12F: dout <= 8'b00000000; //  303 :   0 - 0x0
      11'h130: dout <= 8'b00000000; //  304 :   0 - 0x0 -- Background 0x26
      11'h131: dout <= 8'b00000000; //  305 :   0 - 0x0
      11'h132: dout <= 8'b00000000; //  306 :   0 - 0x0
      11'h133: dout <= 8'b00000000; //  307 :   0 - 0x0
      11'h134: dout <= 8'b00000000; //  308 :   0 - 0x0
      11'h135: dout <= 8'b00000000; //  309 :   0 - 0x0
      11'h136: dout <= 8'b00000000; //  310 :   0 - 0x0
      11'h137: dout <= 8'b00000000; //  311 :   0 - 0x0
      11'h138: dout <= 8'b00000000; //  312 :   0 - 0x0 -- Background 0x27
      11'h139: dout <= 8'b00000000; //  313 :   0 - 0x0
      11'h13A: dout <= 8'b00000000; //  314 :   0 - 0x0
      11'h13B: dout <= 8'b00000000; //  315 :   0 - 0x0
      11'h13C: dout <= 8'b00000000; //  316 :   0 - 0x0
      11'h13D: dout <= 8'b00000000; //  317 :   0 - 0x0
      11'h13E: dout <= 8'b00000000; //  318 :   0 - 0x0
      11'h13F: dout <= 8'b00000000; //  319 :   0 - 0x0
      11'h140: dout <= 8'b00000000; //  320 :   0 - 0x0 -- Background 0x28
      11'h141: dout <= 8'b00000000; //  321 :   0 - 0x0
      11'h142: dout <= 8'b00000000; //  322 :   0 - 0x0
      11'h143: dout <= 8'b00000000; //  323 :   0 - 0x0
      11'h144: dout <= 8'b00000000; //  324 :   0 - 0x0
      11'h145: dout <= 8'b00000000; //  325 :   0 - 0x0
      11'h146: dout <= 8'b00000000; //  326 :   0 - 0x0
      11'h147: dout <= 8'b00000000; //  327 :   0 - 0x0
      11'h148: dout <= 8'b00100000; //  328 :  32 - 0x20 -- Background 0x29
      11'h149: dout <= 8'b00100000; //  329 :  32 - 0x20
      11'h14A: dout <= 8'b00100000; //  330 :  32 - 0x20
      11'h14B: dout <= 8'b00100000; //  331 :  32 - 0x20
      11'h14C: dout <= 8'b00010011; //  332 :  19 - 0x13
      11'h14D: dout <= 8'b00001101; //  333 :  13 - 0xd
      11'h14E: dout <= 8'b00000010; //  334 :   2 - 0x2
      11'h14F: dout <= 8'b00000001; //  335 :   1 - 0x1
      11'h150: dout <= 8'b00100000; //  336 :  32 - 0x20 -- Background 0x2a
      11'h151: dout <= 8'b00100000; //  337 :  32 - 0x20
      11'h152: dout <= 8'b00100000; //  338 :  32 - 0x20
      11'h153: dout <= 8'b00100000; //  339 :  32 - 0x20
      11'h154: dout <= 8'b00010011; //  340 :  19 - 0x13
      11'h155: dout <= 8'b00001101; //  341 :  13 - 0xd
      11'h156: dout <= 8'b00000001; //  342 :   1 - 0x1
      11'h157: dout <= 8'b00000001; //  343 :   1 - 0x1
      11'h158: dout <= 8'b00000000; //  344 :   0 - 0x0 -- Background 0x2b
      11'h159: dout <= 8'b00000000; //  345 :   0 - 0x0
      11'h15A: dout <= 8'b00000000; //  346 :   0 - 0x0
      11'h15B: dout <= 8'b00000000; //  347 :   0 - 0x0
      11'h15C: dout <= 8'b00000000; //  348 :   0 - 0x0
      11'h15D: dout <= 8'b00000000; //  349 :   0 - 0x0
      11'h15E: dout <= 8'b00000000; //  350 :   0 - 0x0
      11'h15F: dout <= 8'b00000000; //  351 :   0 - 0x0
      11'h160: dout <= 8'b00000000; //  352 :   0 - 0x0 -- Background 0x2c
      11'h161: dout <= 8'b00000000; //  353 :   0 - 0x0
      11'h162: dout <= 8'b00000000; //  354 :   0 - 0x0
      11'h163: dout <= 8'b00000000; //  355 :   0 - 0x0
      11'h164: dout <= 8'b00000000; //  356 :   0 - 0x0
      11'h165: dout <= 8'b00000000; //  357 :   0 - 0x0
      11'h166: dout <= 8'b00000000; //  358 :   0 - 0x0
      11'h167: dout <= 8'b00000000; //  359 :   0 - 0x0
      11'h168: dout <= 8'b00111100; //  360 :  60 - 0x3c -- Background 0x2d
      11'h169: dout <= 8'b00000000; //  361 :   0 - 0x0
      11'h16A: dout <= 8'b10000001; //  362 : 129 - 0x81
      11'h16B: dout <= 8'b10011001; //  363 : 153 - 0x99
      11'h16C: dout <= 8'b10011001; //  364 : 153 - 0x99
      11'h16D: dout <= 8'b10000001; //  365 : 129 - 0x81
      11'h16E: dout <= 8'b00000000; //  366 :   0 - 0x0
      11'h16F: dout <= 8'b00111100; //  367 :  60 - 0x3c
      11'h170: dout <= 8'b00000000; //  368 :   0 - 0x0 -- Background 0x2e
      11'h171: dout <= 8'b00000000; //  369 :   0 - 0x0
      11'h172: dout <= 8'b00000000; //  370 :   0 - 0x0
      11'h173: dout <= 8'b00000000; //  371 :   0 - 0x0
      11'h174: dout <= 8'b00000000; //  372 :   0 - 0x0
      11'h175: dout <= 8'b00000000; //  373 :   0 - 0x0
      11'h176: dout <= 8'b00000000; //  374 :   0 - 0x0
      11'h177: dout <= 8'b00000000; //  375 :   0 - 0x0
      11'h178: dout <= 8'b10011111; //  376 : 159 - 0x9f -- Background 0x2f
      11'h179: dout <= 8'b10011110; //  377 : 158 - 0x9e
      11'h17A: dout <= 8'b10011100; //  378 : 156 - 0x9c
      11'h17B: dout <= 8'b00011000; //  379 :  24 - 0x18
      11'h17C: dout <= 8'b00111000; //  380 :  56 - 0x38
      11'h17D: dout <= 8'b11111100; //  381 : 252 - 0xfc
      11'h17E: dout <= 8'b11111100; //  382 : 252 - 0xfc
      11'h17F: dout <= 8'b11111100; //  383 : 252 - 0xfc
      11'h180: dout <= 8'b01111111; //  384 : 127 - 0x7f -- Background 0x30
      11'h181: dout <= 8'b01111110; //  385 : 126 - 0x7e
      11'h182: dout <= 8'b11111100; //  386 : 252 - 0xfc
      11'h183: dout <= 8'b00111000; //  387 :  56 - 0x38
      11'h184: dout <= 8'b00111000; //  388 :  56 - 0x38
      11'h185: dout <= 8'b00000100; //  389 :   4 - 0x4
      11'h186: dout <= 8'b10000100; //  390 : 132 - 0x84
      11'h187: dout <= 8'b11111100; //  391 : 252 - 0xfc
      11'h188: dout <= 8'b01111111; //  392 : 127 - 0x7f -- Background 0x31
      11'h189: dout <= 8'b01111110; //  393 : 126 - 0x7e
      11'h18A: dout <= 8'b11111100; //  394 : 252 - 0xfc
      11'h18B: dout <= 8'b00111000; //  395 :  56 - 0x38
      11'h18C: dout <= 8'b00111000; //  396 :  56 - 0x38
      11'h18D: dout <= 8'b00011100; //  397 :  28 - 0x1c
      11'h18E: dout <= 8'b10000100; //  398 : 132 - 0x84
      11'h18F: dout <= 8'b11000100; //  399 : 196 - 0xc4
      11'h190: dout <= 8'b01111111; //  400 : 127 - 0x7f -- Background 0x32
      11'h191: dout <= 8'b01111110; //  401 : 126 - 0x7e
      11'h192: dout <= 8'b11111100; //  402 : 252 - 0xfc
      11'h193: dout <= 8'b00111000; //  403 :  56 - 0x38
      11'h194: dout <= 8'b00100100; //  404 :  36 - 0x24
      11'h195: dout <= 8'b00000100; //  405 :   4 - 0x4
      11'h196: dout <= 8'b10011100; //  406 : 156 - 0x9c
      11'h197: dout <= 8'b11111100; //  407 : 252 - 0xfc
      11'h198: dout <= 8'b00100011; //  408 :  35 - 0x23 -- Background 0x33
      11'h199: dout <= 8'b00100011; //  409 :  35 - 0x23
      11'h19A: dout <= 8'b00100001; //  410 :  33 - 0x21
      11'h19B: dout <= 8'b00100000; //  411 :  32 - 0x20
      11'h19C: dout <= 8'b00010011; //  412 :  19 - 0x13
      11'h19D: dout <= 8'b00001101; //  413 :  13 - 0xd
      11'h19E: dout <= 8'b00000001; //  414 :   1 - 0x1
      11'h19F: dout <= 8'b00000001; //  415 :   1 - 0x1
      11'h1A0: dout <= 8'b11111100; //  416 : 252 - 0xfc -- Background 0x34
      11'h1A1: dout <= 8'b11111100; //  417 : 252 - 0xfc
      11'h1A2: dout <= 8'b11111100; //  418 : 252 - 0xfc
      11'h1A3: dout <= 8'b11111100; //  419 : 252 - 0xfc
      11'h1A4: dout <= 8'b10100100; //  420 : 164 - 0xa4
      11'h1A5: dout <= 8'b00100100; //  421 :  36 - 0x24
      11'h1A6: dout <= 8'b00010010; //  422 :  18 - 0x12
      11'h1A7: dout <= 8'b11101110; //  423 : 238 - 0xee
      11'h1A8: dout <= 8'b00100011; //  424 :  35 - 0x23 -- Background 0x35
      11'h1A9: dout <= 8'b00100011; //  425 :  35 - 0x23
      11'h1AA: dout <= 8'b00100001; //  426 :  33 - 0x21
      11'h1AB: dout <= 8'b00100000; //  427 :  32 - 0x20
      11'h1AC: dout <= 8'b00010011; //  428 :  19 - 0x13
      11'h1AD: dout <= 8'b00001110; //  429 :  14 - 0xe
      11'h1AE: dout <= 8'b00000010; //  430 :   2 - 0x2
      11'h1AF: dout <= 8'b00000001; //  431 :   1 - 0x1
      11'h1B0: dout <= 8'b11111100; //  432 : 252 - 0xfc -- Background 0x36
      11'h1B1: dout <= 8'b11111100; //  433 : 252 - 0xfc
      11'h1B2: dout <= 8'b11111100; //  434 : 252 - 0xfc
      11'h1B3: dout <= 8'b11111100; //  435 : 252 - 0xfc
      11'h1B4: dout <= 8'b10100110; //  436 : 166 - 0xa6
      11'h1B5: dout <= 8'b00110001; //  437 :  49 - 0x31
      11'h1B6: dout <= 8'b01001001; //  438 :  73 - 0x49
      11'h1B7: dout <= 8'b11000110; //  439 : 198 - 0xc6
      11'h1B8: dout <= 8'b11111100; //  440 : 252 - 0xfc -- Background 0x37
      11'h1B9: dout <= 8'b11111100; //  441 : 252 - 0xfc
      11'h1BA: dout <= 8'b11111100; //  442 : 252 - 0xfc
      11'h1BB: dout <= 8'b11111100; //  443 : 252 - 0xfc
      11'h1BC: dout <= 8'b10100100; //  444 : 164 - 0xa4
      11'h1BD: dout <= 8'b00100100; //  445 :  36 - 0x24
      11'h1BE: dout <= 8'b00010010; //  446 :  18 - 0x12
      11'h1BF: dout <= 8'b11101110; //  447 : 238 - 0xee
      11'h1C0: dout <= 8'b00000000; //  448 :   0 - 0x0 -- Background 0x38
      11'h1C1: dout <= 8'b00000000; //  449 :   0 - 0x0
      11'h1C2: dout <= 8'b00000000; //  450 :   0 - 0x0
      11'h1C3: dout <= 8'b00000000; //  451 :   0 - 0x0
      11'h1C4: dout <= 8'b00000000; //  452 :   0 - 0x0
      11'h1C5: dout <= 8'b00000000; //  453 :   0 - 0x0
      11'h1C6: dout <= 8'b00000000; //  454 :   0 - 0x0
      11'h1C7: dout <= 8'b00000000; //  455 :   0 - 0x0
      11'h1C8: dout <= 8'b00000000; //  456 :   0 - 0x0 -- Background 0x39
      11'h1C9: dout <= 8'b00000000; //  457 :   0 - 0x0
      11'h1CA: dout <= 8'b00000000; //  458 :   0 - 0x0
      11'h1CB: dout <= 8'b00000000; //  459 :   0 - 0x0
      11'h1CC: dout <= 8'b00000000; //  460 :   0 - 0x0
      11'h1CD: dout <= 8'b00000000; //  461 :   0 - 0x0
      11'h1CE: dout <= 8'b00000000; //  462 :   0 - 0x0
      11'h1CF: dout <= 8'b00000000; //  463 :   0 - 0x0
      11'h1D0: dout <= 8'b00000000; //  464 :   0 - 0x0 -- Background 0x3a
      11'h1D1: dout <= 8'b00000000; //  465 :   0 - 0x0
      11'h1D2: dout <= 8'b00000000; //  466 :   0 - 0x0
      11'h1D3: dout <= 8'b00000000; //  467 :   0 - 0x0
      11'h1D4: dout <= 8'b00000000; //  468 :   0 - 0x0
      11'h1D5: dout <= 8'b00000000; //  469 :   0 - 0x0
      11'h1D6: dout <= 8'b00000000; //  470 :   0 - 0x0
      11'h1D7: dout <= 8'b00000000; //  471 :   0 - 0x0
      11'h1D8: dout <= 8'b00000000; //  472 :   0 - 0x0 -- Background 0x3b
      11'h1D9: dout <= 8'b00000000; //  473 :   0 - 0x0
      11'h1DA: dout <= 8'b00000000; //  474 :   0 - 0x0
      11'h1DB: dout <= 8'b00000000; //  475 :   0 - 0x0
      11'h1DC: dout <= 8'b00000000; //  476 :   0 - 0x0
      11'h1DD: dout <= 8'b00000000; //  477 :   0 - 0x0
      11'h1DE: dout <= 8'b00000000; //  478 :   0 - 0x0
      11'h1DF: dout <= 8'b00000000; //  479 :   0 - 0x0
      11'h1E0: dout <= 8'b00000000; //  480 :   0 - 0x0 -- Background 0x3c
      11'h1E1: dout <= 8'b00000000; //  481 :   0 - 0x0
      11'h1E2: dout <= 8'b00000000; //  482 :   0 - 0x0
      11'h1E3: dout <= 8'b00000000; //  483 :   0 - 0x0
      11'h1E4: dout <= 8'b00000000; //  484 :   0 - 0x0
      11'h1E5: dout <= 8'b00000000; //  485 :   0 - 0x0
      11'h1E6: dout <= 8'b00000000; //  486 :   0 - 0x0
      11'h1E7: dout <= 8'b00000000; //  487 :   0 - 0x0
      11'h1E8: dout <= 8'b00000000; //  488 :   0 - 0x0 -- Background 0x3d
      11'h1E9: dout <= 8'b00000000; //  489 :   0 - 0x0
      11'h1EA: dout <= 8'b00000000; //  490 :   0 - 0x0
      11'h1EB: dout <= 8'b00000000; //  491 :   0 - 0x0
      11'h1EC: dout <= 8'b00000000; //  492 :   0 - 0x0
      11'h1ED: dout <= 8'b00000000; //  493 :   0 - 0x0
      11'h1EE: dout <= 8'b00000000; //  494 :   0 - 0x0
      11'h1EF: dout <= 8'b00000000; //  495 :   0 - 0x0
      11'h1F0: dout <= 8'b00000000; //  496 :   0 - 0x0 -- Background 0x3e
      11'h1F1: dout <= 8'b00000000; //  497 :   0 - 0x0
      11'h1F2: dout <= 8'b00000000; //  498 :   0 - 0x0
      11'h1F3: dout <= 8'b00000000; //  499 :   0 - 0x0
      11'h1F4: dout <= 8'b00000000; //  500 :   0 - 0x0
      11'h1F5: dout <= 8'b00000000; //  501 :   0 - 0x0
      11'h1F6: dout <= 8'b00000000; //  502 :   0 - 0x0
      11'h1F7: dout <= 8'b00000000; //  503 :   0 - 0x0
      11'h1F8: dout <= 8'b00000000; //  504 :   0 - 0x0 -- Background 0x3f
      11'h1F9: dout <= 8'b00000000; //  505 :   0 - 0x0
      11'h1FA: dout <= 8'b00000000; //  506 :   0 - 0x0
      11'h1FB: dout <= 8'b00000000; //  507 :   0 - 0x0
      11'h1FC: dout <= 8'b00000000; //  508 :   0 - 0x0
      11'h1FD: dout <= 8'b00000000; //  509 :   0 - 0x0
      11'h1FE: dout <= 8'b00000000; //  510 :   0 - 0x0
      11'h1FF: dout <= 8'b00000000; //  511 :   0 - 0x0
      11'h200: dout <= 8'b00000000; //  512 :   0 - 0x0 -- Background 0x40
      11'h201: dout <= 8'b00111110; //  513 :  62 - 0x3e
      11'h202: dout <= 8'b01111111; //  514 : 127 - 0x7f
      11'h203: dout <= 8'b01111111; //  515 : 127 - 0x7f
      11'h204: dout <= 8'b01111111; //  516 : 127 - 0x7f
      11'h205: dout <= 8'b01111111; //  517 : 127 - 0x7f
      11'h206: dout <= 8'b01111111; //  518 : 127 - 0x7f
      11'h207: dout <= 8'b00111110; //  519 :  62 - 0x3e
      11'h208: dout <= 8'b00000000; //  520 :   0 - 0x0 -- Background 0x41
      11'h209: dout <= 8'b00111100; //  521 :  60 - 0x3c
      11'h20A: dout <= 8'b00011100; //  522 :  28 - 0x1c
      11'h20B: dout <= 8'b00011100; //  523 :  28 - 0x1c
      11'h20C: dout <= 8'b00011100; //  524 :  28 - 0x1c
      11'h20D: dout <= 8'b00011100; //  525 :  28 - 0x1c
      11'h20E: dout <= 8'b00011100; //  526 :  28 - 0x1c
      11'h20F: dout <= 8'b00011100; //  527 :  28 - 0x1c
      11'h210: dout <= 8'b00000000; //  528 :   0 - 0x0 -- Background 0x42
      11'h211: dout <= 8'b01111100; //  529 : 124 - 0x7c
      11'h212: dout <= 8'b01111111; //  530 : 127 - 0x7f
      11'h213: dout <= 8'b01100111; //  531 : 103 - 0x67
      11'h214: dout <= 8'b00111111; //  532 :  63 - 0x3f
      11'h215: dout <= 8'b01111110; //  533 : 126 - 0x7e
      11'h216: dout <= 8'b01111111; //  534 : 127 - 0x7f
      11'h217: dout <= 8'b01111111; //  535 : 127 - 0x7f
      11'h218: dout <= 8'b00000000; //  536 :   0 - 0x0 -- Background 0x43
      11'h219: dout <= 8'b01111110; //  537 : 126 - 0x7e
      11'h21A: dout <= 8'b01111111; //  538 : 127 - 0x7f
      11'h21B: dout <= 8'b01111111; //  539 : 127 - 0x7f
      11'h21C: dout <= 8'b00011111; //  540 :  31 - 0x1f
      11'h21D: dout <= 8'b01110111; //  541 : 119 - 0x77
      11'h21E: dout <= 8'b01111111; //  542 : 127 - 0x7f
      11'h21F: dout <= 8'b01111110; //  543 : 126 - 0x7e
      11'h220: dout <= 8'b00000000; //  544 :   0 - 0x0 -- Background 0x44
      11'h221: dout <= 8'b00001110; //  545 :  14 - 0xe
      11'h222: dout <= 8'b00011110; //  546 :  30 - 0x1e
      11'h223: dout <= 8'b00111110; //  547 :  62 - 0x3e
      11'h224: dout <= 8'b01111110; //  548 : 126 - 0x7e
      11'h225: dout <= 8'b01111111; //  549 : 127 - 0x7f
      11'h226: dout <= 8'b01111110; //  550 : 126 - 0x7e
      11'h227: dout <= 8'b00001100; //  551 :  12 - 0xc
      11'h228: dout <= 8'b00000000; //  552 :   0 - 0x0 -- Background 0x45
      11'h229: dout <= 8'b01111111; //  553 : 127 - 0x7f
      11'h22A: dout <= 8'b01111111; //  554 : 127 - 0x7f
      11'h22B: dout <= 8'b01111111; //  555 : 127 - 0x7f
      11'h22C: dout <= 8'b01111111; //  556 : 127 - 0x7f
      11'h22D: dout <= 8'b01110111; //  557 : 119 - 0x77
      11'h22E: dout <= 8'b01111111; //  558 : 127 - 0x7f
      11'h22F: dout <= 8'b01111110; //  559 : 126 - 0x7e
      11'h230: dout <= 8'b00000000; //  560 :   0 - 0x0 -- Background 0x46
      11'h231: dout <= 8'b00111110; //  561 :  62 - 0x3e
      11'h232: dout <= 8'b01111110; //  562 : 126 - 0x7e
      11'h233: dout <= 8'b01111111; //  563 : 127 - 0x7f
      11'h234: dout <= 8'b01111111; //  564 : 127 - 0x7f
      11'h235: dout <= 8'b01110111; //  565 : 119 - 0x77
      11'h236: dout <= 8'b01111111; //  566 : 127 - 0x7f
      11'h237: dout <= 8'b00111110; //  567 :  62 - 0x3e
      11'h238: dout <= 8'b00000000; //  568 :   0 - 0x0 -- Background 0x47
      11'h239: dout <= 8'b01111110; //  569 : 126 - 0x7e
      11'h23A: dout <= 8'b01111110; //  570 : 126 - 0x7e
      11'h23B: dout <= 8'b00011110; //  571 :  30 - 0x1e
      11'h23C: dout <= 8'b00011100; //  572 :  28 - 0x1c
      11'h23D: dout <= 8'b00111100; //  573 :  60 - 0x3c
      11'h23E: dout <= 8'b00111000; //  574 :  56 - 0x38
      11'h23F: dout <= 8'b00111000; //  575 :  56 - 0x38
      11'h240: dout <= 8'b00000000; //  576 :   0 - 0x0 -- Background 0x48
      11'h241: dout <= 8'b00111110; //  577 :  62 - 0x3e
      11'h242: dout <= 8'b01111111; //  578 : 127 - 0x7f
      11'h243: dout <= 8'b01111111; //  579 : 127 - 0x7f
      11'h244: dout <= 8'b01111111; //  580 : 127 - 0x7f
      11'h245: dout <= 8'b01111111; //  581 : 127 - 0x7f
      11'h246: dout <= 8'b01111111; //  582 : 127 - 0x7f
      11'h247: dout <= 8'b00111110; //  583 :  62 - 0x3e
      11'h248: dout <= 8'b00000000; //  584 :   0 - 0x0 -- Background 0x49
      11'h249: dout <= 8'b00111110; //  585 :  62 - 0x3e
      11'h24A: dout <= 8'b01111111; //  586 : 127 - 0x7f
      11'h24B: dout <= 8'b01110111; //  587 : 119 - 0x77
      11'h24C: dout <= 8'b01111111; //  588 : 127 - 0x7f
      11'h24D: dout <= 8'b01111111; //  589 : 127 - 0x7f
      11'h24E: dout <= 8'b00111111; //  590 :  63 - 0x3f
      11'h24F: dout <= 8'b00111110; //  591 :  62 - 0x3e
      11'h250: dout <= 8'b11111111; //  592 : 255 - 0xff -- Background 0x4a
      11'h251: dout <= 8'b10011001; //  593 : 153 - 0x99
      11'h252: dout <= 8'b10011001; //  594 : 153 - 0x99
      11'h253: dout <= 8'b10011001; //  595 : 153 - 0x99
      11'h254: dout <= 8'b10011001; //  596 : 153 - 0x99
      11'h255: dout <= 8'b10011001; //  597 : 153 - 0x99
      11'h256: dout <= 8'b10011001; //  598 : 153 - 0x99
      11'h257: dout <= 8'b11111111; //  599 : 255 - 0xff
      11'h258: dout <= 8'b11110000; //  600 : 240 - 0xf0 -- Background 0x4b
      11'h259: dout <= 8'b10010000; //  601 : 144 - 0x90
      11'h25A: dout <= 8'b10010000; //  602 : 144 - 0x90
      11'h25B: dout <= 8'b10010000; //  603 : 144 - 0x90
      11'h25C: dout <= 8'b10010000; //  604 : 144 - 0x90
      11'h25D: dout <= 8'b10010000; //  605 : 144 - 0x90
      11'h25E: dout <= 8'b10010000; //  606 : 144 - 0x90
      11'h25F: dout <= 8'b11110000; //  607 : 240 - 0xf0
      11'h260: dout <= 8'b11111111; //  608 : 255 - 0xff -- Background 0x4c
      11'h261: dout <= 8'b11111111; //  609 : 255 - 0xff
      11'h262: dout <= 8'b11111111; //  610 : 255 - 0xff
      11'h263: dout <= 8'b11111111; //  611 : 255 - 0xff
      11'h264: dout <= 8'b11111111; //  612 : 255 - 0xff
      11'h265: dout <= 8'b11111111; //  613 : 255 - 0xff
      11'h266: dout <= 8'b11111111; //  614 : 255 - 0xff
      11'h267: dout <= 8'b11111111; //  615 : 255 - 0xff
      11'h268: dout <= 8'b11111111; //  616 : 255 - 0xff -- Background 0x4d
      11'h269: dout <= 8'b11111111; //  617 : 255 - 0xff
      11'h26A: dout <= 8'b11111111; //  618 : 255 - 0xff
      11'h26B: dout <= 8'b11111111; //  619 : 255 - 0xff
      11'h26C: dout <= 8'b11111111; //  620 : 255 - 0xff
      11'h26D: dout <= 8'b11111111; //  621 : 255 - 0xff
      11'h26E: dout <= 8'b11111111; //  622 : 255 - 0xff
      11'h26F: dout <= 8'b11111111; //  623 : 255 - 0xff
      11'h270: dout <= 8'b11111111; //  624 : 255 - 0xff -- Background 0x4e
      11'h271: dout <= 8'b11111111; //  625 : 255 - 0xff
      11'h272: dout <= 8'b11111111; //  626 : 255 - 0xff
      11'h273: dout <= 8'b11111111; //  627 : 255 - 0xff
      11'h274: dout <= 8'b11111111; //  628 : 255 - 0xff
      11'h275: dout <= 8'b11111111; //  629 : 255 - 0xff
      11'h276: dout <= 8'b11111111; //  630 : 255 - 0xff
      11'h277: dout <= 8'b11111111; //  631 : 255 - 0xff
      11'h278: dout <= 8'b11111111; //  632 : 255 - 0xff -- Background 0x4f
      11'h279: dout <= 8'b11111111; //  633 : 255 - 0xff
      11'h27A: dout <= 8'b11111111; //  634 : 255 - 0xff
      11'h27B: dout <= 8'b11111111; //  635 : 255 - 0xff
      11'h27C: dout <= 8'b11111111; //  636 : 255 - 0xff
      11'h27D: dout <= 8'b11111111; //  637 : 255 - 0xff
      11'h27E: dout <= 8'b11111111; //  638 : 255 - 0xff
      11'h27F: dout <= 8'b11111111; //  639 : 255 - 0xff
      11'h280: dout <= 8'b00010000; //  640 :  16 - 0x10 -- Background 0x50
      11'h281: dout <= 8'b00101000; //  641 :  40 - 0x28
      11'h282: dout <= 8'b11101110; //  642 : 238 - 0xee
      11'h283: dout <= 8'b10000010; //  643 : 130 - 0x82
      11'h284: dout <= 8'b01000100; //  644 :  68 - 0x44
      11'h285: dout <= 8'b01000100; //  645 :  68 - 0x44
      11'h286: dout <= 8'b10010010; //  646 : 146 - 0x92
      11'h287: dout <= 8'b11101110; //  647 : 238 - 0xee
      11'h288: dout <= 8'b00010000; //  648 :  16 - 0x10 -- Background 0x51
      11'h289: dout <= 8'b00101000; //  649 :  40 - 0x28
      11'h28A: dout <= 8'b11101110; //  650 : 238 - 0xee
      11'h28B: dout <= 8'b10000010; //  651 : 130 - 0x82
      11'h28C: dout <= 8'b01000100; //  652 :  68 - 0x44
      11'h28D: dout <= 8'b01000100; //  653 :  68 - 0x44
      11'h28E: dout <= 8'b10010010; //  654 : 146 - 0x92
      11'h28F: dout <= 8'b11101110; //  655 : 238 - 0xee
      11'h290: dout <= 8'b00010000; //  656 :  16 - 0x10 -- Background 0x52
      11'h291: dout <= 8'b00111000; //  657 :  56 - 0x38
      11'h292: dout <= 8'b11111110; //  658 : 254 - 0xfe
      11'h293: dout <= 8'b11111110; //  659 : 254 - 0xfe
      11'h294: dout <= 8'b01111100; //  660 : 124 - 0x7c
      11'h295: dout <= 8'b01111100; //  661 : 124 - 0x7c
      11'h296: dout <= 8'b11111110; //  662 : 254 - 0xfe
      11'h297: dout <= 8'b11101110; //  663 : 238 - 0xee
      11'h298: dout <= 8'b11111111; //  664 : 255 - 0xff -- Background 0x53
      11'h299: dout <= 8'b11111111; //  665 : 255 - 0xff
      11'h29A: dout <= 8'b11111111; //  666 : 255 - 0xff
      11'h29B: dout <= 8'b11111111; //  667 : 255 - 0xff
      11'h29C: dout <= 8'b11111111; //  668 : 255 - 0xff
      11'h29D: dout <= 8'b11111111; //  669 : 255 - 0xff
      11'h29E: dout <= 8'b11111111; //  670 : 255 - 0xff
      11'h29F: dout <= 8'b11111111; //  671 : 255 - 0xff
      11'h2A0: dout <= 8'b00000000; //  672 :   0 - 0x0 -- Background 0x54
      11'h2A1: dout <= 8'b00000000; //  673 :   0 - 0x0
      11'h2A2: dout <= 8'b00000000; //  674 :   0 - 0x0
      11'h2A3: dout <= 8'b00000000; //  675 :   0 - 0x0
      11'h2A4: dout <= 8'b00000000; //  676 :   0 - 0x0
      11'h2A5: dout <= 8'b00000000; //  677 :   0 - 0x0
      11'h2A6: dout <= 8'b00000000; //  678 :   0 - 0x0
      11'h2A7: dout <= 8'b00000000; //  679 :   0 - 0x0
      11'h2A8: dout <= 8'b11111111; //  680 : 255 - 0xff -- Background 0x55
      11'h2A9: dout <= 8'b11111111; //  681 : 255 - 0xff
      11'h2AA: dout <= 8'b11111111; //  682 : 255 - 0xff
      11'h2AB: dout <= 8'b11111111; //  683 : 255 - 0xff
      11'h2AC: dout <= 8'b11111111; //  684 : 255 - 0xff
      11'h2AD: dout <= 8'b11111111; //  685 : 255 - 0xff
      11'h2AE: dout <= 8'b11111111; //  686 : 255 - 0xff
      11'h2AF: dout <= 8'b11111111; //  687 : 255 - 0xff
      11'h2B0: dout <= 8'b00101010; //  688 :  42 - 0x2a -- Background 0x56
      11'h2B1: dout <= 8'b01000101; //  689 :  69 - 0x45
      11'h2B2: dout <= 8'b00001000; //  690 :   8 - 0x8
      11'h2B3: dout <= 8'b00010101; //  691 :  21 - 0x15
      11'h2B4: dout <= 8'b00100000; //  692 :  32 - 0x20
      11'h2B5: dout <= 8'b01000101; //  693 :  69 - 0x45
      11'h2B6: dout <= 8'b10101000; //  694 : 168 - 0xa8
      11'h2B7: dout <= 8'b00000000; //  695 :   0 - 0x0
      11'h2B8: dout <= 8'b00001000; //  696 :   8 - 0x8 -- Background 0x57
      11'h2B9: dout <= 8'b01010101; //  697 :  85 - 0x55
      11'h2BA: dout <= 8'b10100000; //  698 : 160 - 0xa0
      11'h2BB: dout <= 8'b00010000; //  699 :  16 - 0x10
      11'h2BC: dout <= 8'b10000000; //  700 : 128 - 0x80
      11'h2BD: dout <= 8'b00010100; //  701 :  20 - 0x14
      11'h2BE: dout <= 8'b00100010; //  702 :  34 - 0x22
      11'h2BF: dout <= 8'b00000000; //  703 :   0 - 0x0
      11'h2C0: dout <= 8'b11111111; //  704 : 255 - 0xff -- Background 0x58
      11'h2C1: dout <= 8'b11010101; //  705 : 213 - 0xd5
      11'h2C2: dout <= 8'b10100000; //  706 : 160 - 0xa0
      11'h2C3: dout <= 8'b11010000; //  707 : 208 - 0xd0
      11'h2C4: dout <= 8'b10001111; //  708 : 143 - 0x8f
      11'h2C5: dout <= 8'b11001000; //  709 : 200 - 0xc8
      11'h2C6: dout <= 8'b10001000; //  710 : 136 - 0x88
      11'h2C7: dout <= 8'b11001000; //  711 : 200 - 0xc8
      11'h2C8: dout <= 8'b10001000; //  712 : 136 - 0x88 -- Background 0x59
      11'h2C9: dout <= 8'b11001000; //  713 : 200 - 0xc8
      11'h2CA: dout <= 8'b10001000; //  714 : 136 - 0x88
      11'h2CB: dout <= 8'b11001111; //  715 : 207 - 0xcf
      11'h2CC: dout <= 8'b10010000; //  716 : 144 - 0x90
      11'h2CD: dout <= 8'b11100000; //  717 : 224 - 0xe0
      11'h2CE: dout <= 8'b11101010; //  718 : 234 - 0xea
      11'h2CF: dout <= 8'b11111111; //  719 : 255 - 0xff
      11'h2D0: dout <= 8'b11111111; //  720 : 255 - 0xff -- Background 0x5a
      11'h2D1: dout <= 8'b01011011; //  721 :  91 - 0x5b
      11'h2D2: dout <= 8'b00000111; //  722 :   7 - 0x7
      11'h2D3: dout <= 8'b00001001; //  723 :   9 - 0x9
      11'h2D4: dout <= 8'b11110011; //  724 : 243 - 0xf3
      11'h2D5: dout <= 8'b00010001; //  725 :  17 - 0x11
      11'h2D6: dout <= 8'b00010011; //  726 :  19 - 0x13
      11'h2D7: dout <= 8'b00010001; //  727 :  17 - 0x11
      11'h2D8: dout <= 8'b00010011; //  728 :  19 - 0x13 -- Background 0x5b
      11'h2D9: dout <= 8'b00010001; //  729 :  17 - 0x11
      11'h2DA: dout <= 8'b00010011; //  730 :  19 - 0x13
      11'h2DB: dout <= 8'b11110001; //  731 : 241 - 0xf1
      11'h2DC: dout <= 8'b00001011; //  732 :  11 - 0xb
      11'h2DD: dout <= 8'b00000101; //  733 :   5 - 0x5
      11'h2DE: dout <= 8'b10101011; //  734 : 171 - 0xab
      11'h2DF: dout <= 8'b11111111; //  735 : 255 - 0xff
      11'h2E0: dout <= 8'b00011100; //  736 :  28 - 0x1c -- Background 0x5c
      11'h2E1: dout <= 8'b00100010; //  737 :  34 - 0x22
      11'h2E2: dout <= 8'b01000001; //  738 :  65 - 0x41
      11'h2E3: dout <= 8'b01000001; //  739 :  65 - 0x41
      11'h2E4: dout <= 8'b01000001; //  740 :  65 - 0x41
      11'h2E5: dout <= 8'b00100010; //  741 :  34 - 0x22
      11'h2E6: dout <= 8'b00100010; //  742 :  34 - 0x22
      11'h2E7: dout <= 8'b00011100; //  743 :  28 - 0x1c
      11'h2E8: dout <= 8'b00001000; //  744 :   8 - 0x8 -- Background 0x5d
      11'h2E9: dout <= 8'b00010000; //  745 :  16 - 0x10
      11'h2EA: dout <= 8'b00010000; //  746 :  16 - 0x10
      11'h2EB: dout <= 8'b00001000; //  747 :   8 - 0x8
      11'h2EC: dout <= 8'b00000100; //  748 :   4 - 0x4
      11'h2ED: dout <= 8'b00000100; //  749 :   4 - 0x4
      11'h2EE: dout <= 8'b00001000; //  750 :   8 - 0x8
      11'h2EF: dout <= 8'b00010000; //  751 :  16 - 0x10
      11'h2F0: dout <= 8'b00110110; //  752 :  54 - 0x36 -- Background 0x5e
      11'h2F1: dout <= 8'b01101011; //  753 : 107 - 0x6b
      11'h2F2: dout <= 8'b01001001; //  754 :  73 - 0x49
      11'h2F3: dout <= 8'b01000001; //  755 :  65 - 0x41
      11'h2F4: dout <= 8'b01000001; //  756 :  65 - 0x41
      11'h2F5: dout <= 8'b00100010; //  757 :  34 - 0x22
      11'h2F6: dout <= 8'b00010100; //  758 :  20 - 0x14
      11'h2F7: dout <= 8'b00001000; //  759 :   8 - 0x8
      11'h2F8: dout <= 8'b00111110; //  760 :  62 - 0x3e -- Background 0x5f
      11'h2F9: dout <= 8'b01101011; //  761 : 107 - 0x6b
      11'h2FA: dout <= 8'b00100010; //  762 :  34 - 0x22
      11'h2FB: dout <= 8'b01100011; //  763 :  99 - 0x63
      11'h2FC: dout <= 8'b00100010; //  764 :  34 - 0x22
      11'h2FD: dout <= 8'b01100011; //  765 :  99 - 0x63
      11'h2FE: dout <= 8'b00100010; //  766 :  34 - 0x22
      11'h2FF: dout <= 8'b01111111; //  767 : 127 - 0x7f
      11'h300: dout <= 8'b11111111; //  768 : 255 - 0xff -- Background 0x60
      11'h301: dout <= 8'b11111111; //  769 : 255 - 0xff
      11'h302: dout <= 8'b11111111; //  770 : 255 - 0xff
      11'h303: dout <= 8'b11111111; //  771 : 255 - 0xff
      11'h304: dout <= 8'b11010101; //  772 : 213 - 0xd5
      11'h305: dout <= 8'b10101010; //  773 : 170 - 0xaa
      11'h306: dout <= 8'b11010101; //  774 : 213 - 0xd5
      11'h307: dout <= 8'b11111111; //  775 : 255 - 0xff
      11'h308: dout <= 8'b11111111; //  776 : 255 - 0xff -- Background 0x61
      11'h309: dout <= 8'b11111111; //  777 : 255 - 0xff
      11'h30A: dout <= 8'b11111111; //  778 : 255 - 0xff
      11'h30B: dout <= 8'b11111111; //  779 : 255 - 0xff
      11'h30C: dout <= 8'b01010101; //  780 :  85 - 0x55
      11'h30D: dout <= 8'b10101010; //  781 : 170 - 0xaa
      11'h30E: dout <= 8'b01010101; //  782 :  85 - 0x55
      11'h30F: dout <= 8'b11111111; //  783 : 255 - 0xff
      11'h310: dout <= 8'b11111111; //  784 : 255 - 0xff -- Background 0x62
      11'h311: dout <= 8'b11111111; //  785 : 255 - 0xff
      11'h312: dout <= 8'b11111111; //  786 : 255 - 0xff
      11'h313: dout <= 8'b11111111; //  787 : 255 - 0xff
      11'h314: dout <= 8'b01010101; //  788 :  85 - 0x55
      11'h315: dout <= 8'b10101011; //  789 : 171 - 0xab
      11'h316: dout <= 8'b01010101; //  790 :  85 - 0x55
      11'h317: dout <= 8'b11111111; //  791 : 255 - 0xff
      11'h318: dout <= 8'b00000000; //  792 :   0 - 0x0 -- Background 0x63
      11'h319: dout <= 8'b00000000; //  793 :   0 - 0x0
      11'h31A: dout <= 8'b00000000; //  794 :   0 - 0x0
      11'h31B: dout <= 8'b00000000; //  795 :   0 - 0x0
      11'h31C: dout <= 8'b00000000; //  796 :   0 - 0x0
      11'h31D: dout <= 8'b00000000; //  797 :   0 - 0x0
      11'h31E: dout <= 8'b00000000; //  798 :   0 - 0x0
      11'h31F: dout <= 8'b00000000; //  799 :   0 - 0x0
      11'h320: dout <= 8'b00000001; //  800 :   1 - 0x1 -- Background 0x64
      11'h321: dout <= 8'b00000001; //  801 :   1 - 0x1
      11'h322: dout <= 8'b00000011; //  802 :   3 - 0x3
      11'h323: dout <= 8'b00000011; //  803 :   3 - 0x3
      11'h324: dout <= 8'b00000110; //  804 :   6 - 0x6
      11'h325: dout <= 8'b00000110; //  805 :   6 - 0x6
      11'h326: dout <= 8'b00001100; //  806 :  12 - 0xc
      11'h327: dout <= 8'b00001100; //  807 :  12 - 0xc
      11'h328: dout <= 8'b00011000; //  808 :  24 - 0x18 -- Background 0x65
      11'h329: dout <= 8'b00011000; //  809 :  24 - 0x18
      11'h32A: dout <= 8'b00110000; //  810 :  48 - 0x30
      11'h32B: dout <= 8'b00110000; //  811 :  48 - 0x30
      11'h32C: dout <= 8'b01100000; //  812 :  96 - 0x60
      11'h32D: dout <= 8'b01100000; //  813 :  96 - 0x60
      11'h32E: dout <= 8'b11101010; //  814 : 234 - 0xea
      11'h32F: dout <= 8'b11111111; //  815 : 255 - 0xff
      11'h330: dout <= 8'b10000000; //  816 : 128 - 0x80 -- Background 0x66
      11'h331: dout <= 8'b10000000; //  817 : 128 - 0x80
      11'h332: dout <= 8'b11000000; //  818 : 192 - 0xc0
      11'h333: dout <= 8'b01000000; //  819 :  64 - 0x40
      11'h334: dout <= 8'b10100000; //  820 : 160 - 0xa0
      11'h335: dout <= 8'b01100000; //  821 :  96 - 0x60
      11'h336: dout <= 8'b00110000; //  822 :  48 - 0x30
      11'h337: dout <= 8'b00010000; //  823 :  16 - 0x10
      11'h338: dout <= 8'b00101000; //  824 :  40 - 0x28 -- Background 0x67
      11'h339: dout <= 8'b00011000; //  825 :  24 - 0x18
      11'h33A: dout <= 8'b00001100; //  826 :  12 - 0xc
      11'h33B: dout <= 8'b00010100; //  827 :  20 - 0x14
      11'h33C: dout <= 8'b00001010; //  828 :  10 - 0xa
      11'h33D: dout <= 8'b00000110; //  829 :   6 - 0x6
      11'h33E: dout <= 8'b10101011; //  830 : 171 - 0xab
      11'h33F: dout <= 8'b11111111; //  831 : 255 - 0xff
      11'h340: dout <= 8'b00000000; //  832 :   0 - 0x0 -- Background 0x68
      11'h341: dout <= 8'b00000000; //  833 :   0 - 0x0
      11'h342: dout <= 8'b00000000; //  834 :   0 - 0x0
      11'h343: dout <= 8'b00000000; //  835 :   0 - 0x0
      11'h344: dout <= 8'b00000000; //  836 :   0 - 0x0
      11'h345: dout <= 8'b00000000; //  837 :   0 - 0x0
      11'h346: dout <= 8'b00000000; //  838 :   0 - 0x0
      11'h347: dout <= 8'b00000000; //  839 :   0 - 0x0
      11'h348: dout <= 8'b00000000; //  840 :   0 - 0x0 -- Background 0x69
      11'h349: dout <= 8'b00000000; //  841 :   0 - 0x0
      11'h34A: dout <= 8'b00000000; //  842 :   0 - 0x0
      11'h34B: dout <= 8'b00000000; //  843 :   0 - 0x0
      11'h34C: dout <= 8'b00000000; //  844 :   0 - 0x0
      11'h34D: dout <= 8'b00000000; //  845 :   0 - 0x0
      11'h34E: dout <= 8'b00000000; //  846 :   0 - 0x0
      11'h34F: dout <= 8'b00000000; //  847 :   0 - 0x0
      11'h350: dout <= 8'b00000000; //  848 :   0 - 0x0 -- Background 0x6a
      11'h351: dout <= 8'b00000000; //  849 :   0 - 0x0
      11'h352: dout <= 8'b00000000; //  850 :   0 - 0x0
      11'h353: dout <= 8'b00000000; //  851 :   0 - 0x0
      11'h354: dout <= 8'b00000000; //  852 :   0 - 0x0
      11'h355: dout <= 8'b00000000; //  853 :   0 - 0x0
      11'h356: dout <= 8'b00000000; //  854 :   0 - 0x0
      11'h357: dout <= 8'b00000000; //  855 :   0 - 0x0
      11'h358: dout <= 8'b00000000; //  856 :   0 - 0x0 -- Background 0x6b
      11'h359: dout <= 8'b00000000; //  857 :   0 - 0x0
      11'h35A: dout <= 8'b00000000; //  858 :   0 - 0x0
      11'h35B: dout <= 8'b00000000; //  859 :   0 - 0x0
      11'h35C: dout <= 8'b00000000; //  860 :   0 - 0x0
      11'h35D: dout <= 8'b00000000; //  861 :   0 - 0x0
      11'h35E: dout <= 8'b00000000; //  862 :   0 - 0x0
      11'h35F: dout <= 8'b00000000; //  863 :   0 - 0x0
      11'h360: dout <= 8'b00000000; //  864 :   0 - 0x0 -- Background 0x6c
      11'h361: dout <= 8'b00000000; //  865 :   0 - 0x0
      11'h362: dout <= 8'b00000000; //  866 :   0 - 0x0
      11'h363: dout <= 8'b00000000; //  867 :   0 - 0x0
      11'h364: dout <= 8'b00000000; //  868 :   0 - 0x0
      11'h365: dout <= 8'b00000000; //  869 :   0 - 0x0
      11'h366: dout <= 8'b00000000; //  870 :   0 - 0x0
      11'h367: dout <= 8'b00000000; //  871 :   0 - 0x0
      11'h368: dout <= 8'b00000000; //  872 :   0 - 0x0 -- Background 0x6d
      11'h369: dout <= 8'b00000000; //  873 :   0 - 0x0
      11'h36A: dout <= 8'b00000000; //  874 :   0 - 0x0
      11'h36B: dout <= 8'b00000000; //  875 :   0 - 0x0
      11'h36C: dout <= 8'b00000000; //  876 :   0 - 0x0
      11'h36D: dout <= 8'b00000000; //  877 :   0 - 0x0
      11'h36E: dout <= 8'b00000000; //  878 :   0 - 0x0
      11'h36F: dout <= 8'b00000000; //  879 :   0 - 0x0
      11'h370: dout <= 8'b00000000; //  880 :   0 - 0x0 -- Background 0x6e
      11'h371: dout <= 8'b00000000; //  881 :   0 - 0x0
      11'h372: dout <= 8'b00000000; //  882 :   0 - 0x0
      11'h373: dout <= 8'b00000000; //  883 :   0 - 0x0
      11'h374: dout <= 8'b00000000; //  884 :   0 - 0x0
      11'h375: dout <= 8'b00000000; //  885 :   0 - 0x0
      11'h376: dout <= 8'b00000000; //  886 :   0 - 0x0
      11'h377: dout <= 8'b00000000; //  887 :   0 - 0x0
      11'h378: dout <= 8'b00000000; //  888 :   0 - 0x0 -- Background 0x6f
      11'h379: dout <= 8'b00000000; //  889 :   0 - 0x0
      11'h37A: dout <= 8'b00000000; //  890 :   0 - 0x0
      11'h37B: dout <= 8'b00000000; //  891 :   0 - 0x0
      11'h37C: dout <= 8'b00000000; //  892 :   0 - 0x0
      11'h37D: dout <= 8'b00000000; //  893 :   0 - 0x0
      11'h37E: dout <= 8'b00000000; //  894 :   0 - 0x0
      11'h37F: dout <= 8'b00000000; //  895 :   0 - 0x0
      11'h380: dout <= 8'b00000000; //  896 :   0 - 0x0 -- Background 0x70
      11'h381: dout <= 8'b00000000; //  897 :   0 - 0x0
      11'h382: dout <= 8'b00000000; //  898 :   0 - 0x0
      11'h383: dout <= 8'b00000000; //  899 :   0 - 0x0
      11'h384: dout <= 8'b00000000; //  900 :   0 - 0x0
      11'h385: dout <= 8'b00000000; //  901 :   0 - 0x0
      11'h386: dout <= 8'b00000000; //  902 :   0 - 0x0
      11'h387: dout <= 8'b00000000; //  903 :   0 - 0x0
      11'h388: dout <= 8'b00000000; //  904 :   0 - 0x0 -- Background 0x71
      11'h389: dout <= 8'b00000000; //  905 :   0 - 0x0
      11'h38A: dout <= 8'b00000000; //  906 :   0 - 0x0
      11'h38B: dout <= 8'b00000000; //  907 :   0 - 0x0
      11'h38C: dout <= 8'b00000000; //  908 :   0 - 0x0
      11'h38D: dout <= 8'b00000000; //  909 :   0 - 0x0
      11'h38E: dout <= 8'b00000000; //  910 :   0 - 0x0
      11'h38F: dout <= 8'b00000000; //  911 :   0 - 0x0
      11'h390: dout <= 8'b00000000; //  912 :   0 - 0x0 -- Background 0x72
      11'h391: dout <= 8'b00000000; //  913 :   0 - 0x0
      11'h392: dout <= 8'b00000000; //  914 :   0 - 0x0
      11'h393: dout <= 8'b00000000; //  915 :   0 - 0x0
      11'h394: dout <= 8'b00000000; //  916 :   0 - 0x0
      11'h395: dout <= 8'b00000000; //  917 :   0 - 0x0
      11'h396: dout <= 8'b00000000; //  918 :   0 - 0x0
      11'h397: dout <= 8'b00000000; //  919 :   0 - 0x0
      11'h398: dout <= 8'b00000000; //  920 :   0 - 0x0 -- Background 0x73
      11'h399: dout <= 8'b00000000; //  921 :   0 - 0x0
      11'h39A: dout <= 8'b00000000; //  922 :   0 - 0x0
      11'h39B: dout <= 8'b00000000; //  923 :   0 - 0x0
      11'h39C: dout <= 8'b00000000; //  924 :   0 - 0x0
      11'h39D: dout <= 8'b00000000; //  925 :   0 - 0x0
      11'h39E: dout <= 8'b00000000; //  926 :   0 - 0x0
      11'h39F: dout <= 8'b00000000; //  927 :   0 - 0x0
      11'h3A0: dout <= 8'b00000000; //  928 :   0 - 0x0 -- Background 0x74
      11'h3A1: dout <= 8'b00000000; //  929 :   0 - 0x0
      11'h3A2: dout <= 8'b00000000; //  930 :   0 - 0x0
      11'h3A3: dout <= 8'b00000000; //  931 :   0 - 0x0
      11'h3A4: dout <= 8'b00000000; //  932 :   0 - 0x0
      11'h3A5: dout <= 8'b00000000; //  933 :   0 - 0x0
      11'h3A6: dout <= 8'b00000000; //  934 :   0 - 0x0
      11'h3A7: dout <= 8'b00000000; //  935 :   0 - 0x0
      11'h3A8: dout <= 8'b00000000; //  936 :   0 - 0x0 -- Background 0x75
      11'h3A9: dout <= 8'b00000000; //  937 :   0 - 0x0
      11'h3AA: dout <= 8'b00000000; //  938 :   0 - 0x0
      11'h3AB: dout <= 8'b00000000; //  939 :   0 - 0x0
      11'h3AC: dout <= 8'b00000000; //  940 :   0 - 0x0
      11'h3AD: dout <= 8'b00000000; //  941 :   0 - 0x0
      11'h3AE: dout <= 8'b00000000; //  942 :   0 - 0x0
      11'h3AF: dout <= 8'b00000000; //  943 :   0 - 0x0
      11'h3B0: dout <= 8'b00000000; //  944 :   0 - 0x0 -- Background 0x76
      11'h3B1: dout <= 8'b00000000; //  945 :   0 - 0x0
      11'h3B2: dout <= 8'b00000000; //  946 :   0 - 0x0
      11'h3B3: dout <= 8'b00000000; //  947 :   0 - 0x0
      11'h3B4: dout <= 8'b00000000; //  948 :   0 - 0x0
      11'h3B5: dout <= 8'b00000000; //  949 :   0 - 0x0
      11'h3B6: dout <= 8'b00000000; //  950 :   0 - 0x0
      11'h3B7: dout <= 8'b00000000; //  951 :   0 - 0x0
      11'h3B8: dout <= 8'b00000000; //  952 :   0 - 0x0 -- Background 0x77
      11'h3B9: dout <= 8'b00000000; //  953 :   0 - 0x0
      11'h3BA: dout <= 8'b00000000; //  954 :   0 - 0x0
      11'h3BB: dout <= 8'b00000000; //  955 :   0 - 0x0
      11'h3BC: dout <= 8'b00000000; //  956 :   0 - 0x0
      11'h3BD: dout <= 8'b00000000; //  957 :   0 - 0x0
      11'h3BE: dout <= 8'b00000000; //  958 :   0 - 0x0
      11'h3BF: dout <= 8'b00000000; //  959 :   0 - 0x0
      11'h3C0: dout <= 8'b00000000; //  960 :   0 - 0x0 -- Background 0x78
      11'h3C1: dout <= 8'b00000000; //  961 :   0 - 0x0
      11'h3C2: dout <= 8'b00000000; //  962 :   0 - 0x0
      11'h3C3: dout <= 8'b00000000; //  963 :   0 - 0x0
      11'h3C4: dout <= 8'b00000000; //  964 :   0 - 0x0
      11'h3C5: dout <= 8'b00000000; //  965 :   0 - 0x0
      11'h3C6: dout <= 8'b00000000; //  966 :   0 - 0x0
      11'h3C7: dout <= 8'b00000000; //  967 :   0 - 0x0
      11'h3C8: dout <= 8'b00000000; //  968 :   0 - 0x0 -- Background 0x79
      11'h3C9: dout <= 8'b00000000; //  969 :   0 - 0x0
      11'h3CA: dout <= 8'b00000000; //  970 :   0 - 0x0
      11'h3CB: dout <= 8'b00000000; //  971 :   0 - 0x0
      11'h3CC: dout <= 8'b00000000; //  972 :   0 - 0x0
      11'h3CD: dout <= 8'b00000000; //  973 :   0 - 0x0
      11'h3CE: dout <= 8'b00000000; //  974 :   0 - 0x0
      11'h3CF: dout <= 8'b00000000; //  975 :   0 - 0x0
      11'h3D0: dout <= 8'b00000000; //  976 :   0 - 0x0 -- Background 0x7a
      11'h3D1: dout <= 8'b00000000; //  977 :   0 - 0x0
      11'h3D2: dout <= 8'b00000000; //  978 :   0 - 0x0
      11'h3D3: dout <= 8'b00000000; //  979 :   0 - 0x0
      11'h3D4: dout <= 8'b00000000; //  980 :   0 - 0x0
      11'h3D5: dout <= 8'b00000000; //  981 :   0 - 0x0
      11'h3D6: dout <= 8'b00000000; //  982 :   0 - 0x0
      11'h3D7: dout <= 8'b00000000; //  983 :   0 - 0x0
      11'h3D8: dout <= 8'b00000000; //  984 :   0 - 0x0 -- Background 0x7b
      11'h3D9: dout <= 8'b00000000; //  985 :   0 - 0x0
      11'h3DA: dout <= 8'b00000000; //  986 :   0 - 0x0
      11'h3DB: dout <= 8'b00000000; //  987 :   0 - 0x0
      11'h3DC: dout <= 8'b00000000; //  988 :   0 - 0x0
      11'h3DD: dout <= 8'b00000000; //  989 :   0 - 0x0
      11'h3DE: dout <= 8'b00000000; //  990 :   0 - 0x0
      11'h3DF: dout <= 8'b00000000; //  991 :   0 - 0x0
      11'h3E0: dout <= 8'b00000000; //  992 :   0 - 0x0 -- Background 0x7c
      11'h3E1: dout <= 8'b00000000; //  993 :   0 - 0x0
      11'h3E2: dout <= 8'b00000000; //  994 :   0 - 0x0
      11'h3E3: dout <= 8'b00000000; //  995 :   0 - 0x0
      11'h3E4: dout <= 8'b00000000; //  996 :   0 - 0x0
      11'h3E5: dout <= 8'b00000000; //  997 :   0 - 0x0
      11'h3E6: dout <= 8'b00000000; //  998 :   0 - 0x0
      11'h3E7: dout <= 8'b00000000; //  999 :   0 - 0x0
      11'h3E8: dout <= 8'b00000000; // 1000 :   0 - 0x0 -- Background 0x7d
      11'h3E9: dout <= 8'b00000000; // 1001 :   0 - 0x0
      11'h3EA: dout <= 8'b00000000; // 1002 :   0 - 0x0
      11'h3EB: dout <= 8'b00000000; // 1003 :   0 - 0x0
      11'h3EC: dout <= 8'b00000000; // 1004 :   0 - 0x0
      11'h3ED: dout <= 8'b00000000; // 1005 :   0 - 0x0
      11'h3EE: dout <= 8'b00000000; // 1006 :   0 - 0x0
      11'h3EF: dout <= 8'b00000000; // 1007 :   0 - 0x0
      11'h3F0: dout <= 8'b00000000; // 1008 :   0 - 0x0 -- Background 0x7e
      11'h3F1: dout <= 8'b00000000; // 1009 :   0 - 0x0
      11'h3F2: dout <= 8'b00000000; // 1010 :   0 - 0x0
      11'h3F3: dout <= 8'b00000000; // 1011 :   0 - 0x0
      11'h3F4: dout <= 8'b00000000; // 1012 :   0 - 0x0
      11'h3F5: dout <= 8'b00000000; // 1013 :   0 - 0x0
      11'h3F6: dout <= 8'b00000000; // 1014 :   0 - 0x0
      11'h3F7: dout <= 8'b00000000; // 1015 :   0 - 0x0
      11'h3F8: dout <= 8'b00000000; // 1016 :   0 - 0x0 -- Background 0x7f
      11'h3F9: dout <= 8'b00000000; // 1017 :   0 - 0x0
      11'h3FA: dout <= 8'b00000000; // 1018 :   0 - 0x0
      11'h3FB: dout <= 8'b00000000; // 1019 :   0 - 0x0
      11'h3FC: dout <= 8'b00000000; // 1020 :   0 - 0x0
      11'h3FD: dout <= 8'b00000000; // 1021 :   0 - 0x0
      11'h3FE: dout <= 8'b00000000; // 1022 :   0 - 0x0
      11'h3FF: dout <= 8'b00000000; // 1023 :   0 - 0x0
      11'h400: dout <= 8'b00000011; // 1024 :   3 - 0x3 -- Background 0x80
      11'h401: dout <= 8'b00001111; // 1025 :  15 - 0xf
      11'h402: dout <= 8'b00011100; // 1026 :  28 - 0x1c
      11'h403: dout <= 8'b00110000; // 1027 :  48 - 0x30
      11'h404: dout <= 8'b00100000; // 1028 :  32 - 0x20
      11'h405: dout <= 8'b01000000; // 1029 :  64 - 0x40
      11'h406: dout <= 8'b01000000; // 1030 :  64 - 0x40
      11'h407: dout <= 8'b01111111; // 1031 : 127 - 0x7f
      11'h408: dout <= 8'b00000001; // 1032 :   1 - 0x1 -- Background 0x81
      11'h409: dout <= 8'b00000001; // 1033 :   1 - 0x1
      11'h40A: dout <= 8'b00000001; // 1034 :   1 - 0x1
      11'h40B: dout <= 8'b00000001; // 1035 :   1 - 0x1
      11'h40C: dout <= 8'b00000001; // 1036 :   1 - 0x1
      11'h40D: dout <= 8'b00000001; // 1037 :   1 - 0x1
      11'h40E: dout <= 8'b00000011; // 1038 :   3 - 0x3
      11'h40F: dout <= 8'b00000011; // 1039 :   3 - 0x3
      11'h410: dout <= 8'b11000000; // 1040 : 192 - 0xc0 -- Background 0x82
      11'h411: dout <= 8'b11110000; // 1041 : 240 - 0xf0
      11'h412: dout <= 8'b00111000; // 1042 :  56 - 0x38
      11'h413: dout <= 8'b00001110; // 1043 :  14 - 0xe
      11'h414: dout <= 8'b00011110; // 1044 :  30 - 0x1e
      11'h415: dout <= 8'b00011110; // 1045 :  30 - 0x1e
      11'h416: dout <= 8'b00000010; // 1046 :   2 - 0x2
      11'h417: dout <= 8'b11111110; // 1047 : 254 - 0xfe
      11'h418: dout <= 8'b10000000; // 1048 : 128 - 0x80 -- Background 0x83
      11'h419: dout <= 8'b10000000; // 1049 : 128 - 0x80
      11'h41A: dout <= 8'b10000000; // 1050 : 128 - 0x80
      11'h41B: dout <= 8'b10000000; // 1051 : 128 - 0x80
      11'h41C: dout <= 8'b10000000; // 1052 : 128 - 0x80
      11'h41D: dout <= 8'b11100000; // 1053 : 224 - 0xe0
      11'h41E: dout <= 8'b00010000; // 1054 :  16 - 0x10
      11'h41F: dout <= 8'b11110000; // 1055 : 240 - 0xf0
      11'h420: dout <= 8'b00000011; // 1056 :   3 - 0x3 -- Background 0x84
      11'h421: dout <= 8'b00001111; // 1057 :  15 - 0xf
      11'h422: dout <= 8'b00011100; // 1058 :  28 - 0x1c
      11'h423: dout <= 8'b00110000; // 1059 :  48 - 0x30
      11'h424: dout <= 8'b00100000; // 1060 :  32 - 0x20
      11'h425: dout <= 8'b01000000; // 1061 :  64 - 0x40
      11'h426: dout <= 8'b01000000; // 1062 :  64 - 0x40
      11'h427: dout <= 8'b01111111; // 1063 : 127 - 0x7f
      11'h428: dout <= 8'b00000011; // 1064 :   3 - 0x3 -- Background 0x85
      11'h429: dout <= 8'b00000110; // 1065 :   6 - 0x6
      11'h42A: dout <= 8'b00000110; // 1066 :   6 - 0x6
      11'h42B: dout <= 8'b00011100; // 1067 :  28 - 0x1c
      11'h42C: dout <= 8'b00011000; // 1068 :  24 - 0x18
      11'h42D: dout <= 8'b00110110; // 1069 :  54 - 0x36
      11'h42E: dout <= 8'b00110001; // 1070 :  49 - 0x31
      11'h42F: dout <= 8'b00001111; // 1071 :  15 - 0xf
      11'h430: dout <= 8'b11000000; // 1072 : 192 - 0xc0 -- Background 0x86
      11'h431: dout <= 8'b11110000; // 1073 : 240 - 0xf0
      11'h432: dout <= 8'b00111000; // 1074 :  56 - 0x38
      11'h433: dout <= 8'b00001110; // 1075 :  14 - 0xe
      11'h434: dout <= 8'b00011110; // 1076 :  30 - 0x1e
      11'h435: dout <= 8'b00011110; // 1077 :  30 - 0x1e
      11'h436: dout <= 8'b00000010; // 1078 :   2 - 0x2
      11'h437: dout <= 8'b11111110; // 1079 : 254 - 0xfe
      11'h438: dout <= 8'b11000000; // 1080 : 192 - 0xc0 -- Background 0x87
      11'h439: dout <= 8'b01100000; // 1081 :  96 - 0x60
      11'h43A: dout <= 8'b01100000; // 1082 :  96 - 0x60
      11'h43B: dout <= 8'b00110000; // 1083 :  48 - 0x30
      11'h43C: dout <= 8'b00111110; // 1084 :  62 - 0x3e
      11'h43D: dout <= 8'b00011001; // 1085 :  25 - 0x19
      11'h43E: dout <= 8'b00110011; // 1086 :  51 - 0x33
      11'h43F: dout <= 8'b00111100; // 1087 :  60 - 0x3c
      11'h440: dout <= 8'b00000011; // 1088 :   3 - 0x3 -- Background 0x88
      11'h441: dout <= 8'b00000111; // 1089 :   7 - 0x7
      11'h442: dout <= 8'b00000111; // 1090 :   7 - 0x7
      11'h443: dout <= 8'b00001011; // 1091 :  11 - 0xb
      11'h444: dout <= 8'b00010000; // 1092 :  16 - 0x10
      11'h445: dout <= 8'b01100000; // 1093 :  96 - 0x60
      11'h446: dout <= 8'b11110000; // 1094 : 240 - 0xf0
      11'h447: dout <= 8'b11110000; // 1095 : 240 - 0xf0
      11'h448: dout <= 8'b11110000; // 1096 : 240 - 0xf0 -- Background 0x89
      11'h449: dout <= 8'b11110000; // 1097 : 240 - 0xf0
      11'h44A: dout <= 8'b01100000; // 1098 :  96 - 0x60
      11'h44B: dout <= 8'b00010000; // 1099 :  16 - 0x10
      11'h44C: dout <= 8'b00001011; // 1100 :  11 - 0xb
      11'h44D: dout <= 8'b00000111; // 1101 :   7 - 0x7
      11'h44E: dout <= 8'b00000111; // 1102 :   7 - 0x7
      11'h44F: dout <= 8'b00000011; // 1103 :   3 - 0x3
      11'h450: dout <= 8'b00000000; // 1104 :   0 - 0x0 -- Background 0x8a
      11'h451: dout <= 8'b00011100; // 1105 :  28 - 0x1c
      11'h452: dout <= 8'b00111111; // 1106 :  63 - 0x3f
      11'h453: dout <= 8'b01111000; // 1107 : 120 - 0x78
      11'h454: dout <= 8'b01110000; // 1108 : 112 - 0x70
      11'h455: dout <= 8'b01100000; // 1109 :  96 - 0x60
      11'h456: dout <= 8'b00100000; // 1110 :  32 - 0x20
      11'h457: dout <= 8'b00100000; // 1111 :  32 - 0x20
      11'h458: dout <= 8'b00100000; // 1112 :  32 - 0x20 -- Background 0x8b
      11'h459: dout <= 8'b00100000; // 1113 :  32 - 0x20
      11'h45A: dout <= 8'b01100000; // 1114 :  96 - 0x60
      11'h45B: dout <= 8'b01110000; // 1115 : 112 - 0x70
      11'h45C: dout <= 8'b01111000; // 1116 : 120 - 0x78
      11'h45D: dout <= 8'b00111111; // 1117 :  63 - 0x3f
      11'h45E: dout <= 8'b00011100; // 1118 :  28 - 0x1c
      11'h45F: dout <= 8'b00000000; // 1119 :   0 - 0x0
      11'h460: dout <= 8'b00000011; // 1120 :   3 - 0x3 -- Background 0x8c
      11'h461: dout <= 8'b00001100; // 1121 :  12 - 0xc
      11'h462: dout <= 8'b00011110; // 1122 :  30 - 0x1e
      11'h463: dout <= 8'b00100110; // 1123 :  38 - 0x26
      11'h464: dout <= 8'b01000110; // 1124 :  70 - 0x46
      11'h465: dout <= 8'b01100100; // 1125 : 100 - 0x64
      11'h466: dout <= 8'b01110000; // 1126 : 112 - 0x70
      11'h467: dout <= 8'b11110000; // 1127 : 240 - 0xf0
      11'h468: dout <= 8'b10101010; // 1128 : 170 - 0xaa -- Background 0x8d
      11'h469: dout <= 8'b11111111; // 1129 : 255 - 0xff
      11'h46A: dout <= 8'b01111111; // 1130 : 127 - 0x7f
      11'h46B: dout <= 8'b00111001; // 1131 :  57 - 0x39
      11'h46C: dout <= 8'b00011001; // 1132 :  25 - 0x19
      11'h46D: dout <= 8'b00001011; // 1133 :  11 - 0xb
      11'h46E: dout <= 8'b00001000; // 1134 :   8 - 0x8
      11'h46F: dout <= 8'b00000111; // 1135 :   7 - 0x7
      11'h470: dout <= 8'b11000000; // 1136 : 192 - 0xc0 -- Background 0x8e
      11'h471: dout <= 8'b00110000; // 1137 :  48 - 0x30
      11'h472: dout <= 8'b00001000; // 1138 :   8 - 0x8
      11'h473: dout <= 8'b01000100; // 1139 :  68 - 0x44
      11'h474: dout <= 8'b01100010; // 1140 :  98 - 0x62
      11'h475: dout <= 8'b01100010; // 1141 :  98 - 0x62
      11'h476: dout <= 8'b00000001; // 1142 :   1 - 0x1
      11'h477: dout <= 8'b00111111; // 1143 :  63 - 0x3f
      11'h478: dout <= 8'b10001011; // 1144 : 139 - 0x8b -- Background 0x8f
      11'h479: dout <= 8'b11000001; // 1145 : 193 - 0xc1
      11'h47A: dout <= 8'b11111110; // 1146 : 254 - 0xfe
      11'h47B: dout <= 8'b11111100; // 1147 : 252 - 0xfc
      11'h47C: dout <= 8'b11110000; // 1148 : 240 - 0xf0
      11'h47D: dout <= 8'b11110000; // 1149 : 240 - 0xf0
      11'h47E: dout <= 8'b11111000; // 1150 : 248 - 0xf8
      11'h47F: dout <= 8'b11110000; // 1151 : 240 - 0xf0
      11'h480: dout <= 8'b00000011; // 1152 :   3 - 0x3 -- Background 0x90
      11'h481: dout <= 8'b00001110; // 1153 :  14 - 0xe
      11'h482: dout <= 8'b00010110; // 1154 :  22 - 0x16
      11'h483: dout <= 8'b00100110; // 1155 :  38 - 0x26
      11'h484: dout <= 8'b01100011; // 1156 :  99 - 0x63
      11'h485: dout <= 8'b01110010; // 1157 : 114 - 0x72
      11'h486: dout <= 8'b01110000; // 1158 : 112 - 0x70
      11'h487: dout <= 8'b11010000; // 1159 : 208 - 0xd0
      11'h488: dout <= 8'b10101010; // 1160 : 170 - 0xaa -- Background 0x91
      11'h489: dout <= 8'b11111111; // 1161 : 255 - 0xff
      11'h48A: dout <= 8'b01111111; // 1162 : 127 - 0x7f
      11'h48B: dout <= 8'b00111100; // 1163 :  60 - 0x3c
      11'h48C: dout <= 8'b00011100; // 1164 :  28 - 0x1c
      11'h48D: dout <= 8'b00000100; // 1165 :   4 - 0x4
      11'h48E: dout <= 8'b00000010; // 1166 :   2 - 0x2
      11'h48F: dout <= 8'b00000001; // 1167 :   1 - 0x1
      11'h490: dout <= 8'b11000000; // 1168 : 192 - 0xc0 -- Background 0x92
      11'h491: dout <= 8'b00110000; // 1169 :  48 - 0x30
      11'h492: dout <= 8'b00001000; // 1170 :   8 - 0x8
      11'h493: dout <= 8'b00100100; // 1171 :  36 - 0x24
      11'h494: dout <= 8'b00110010; // 1172 :  50 - 0x32
      11'h495: dout <= 8'b00110010; // 1173 :  50 - 0x32
      11'h496: dout <= 8'b00000001; // 1174 :   1 - 0x1
      11'h497: dout <= 8'b00011111; // 1175 :  31 - 0x1f
      11'h498: dout <= 8'b10001011; // 1176 : 139 - 0x8b -- Background 0x93
      11'h499: dout <= 8'b11000001; // 1177 : 193 - 0xc1
      11'h49A: dout <= 8'b11111110; // 1178 : 254 - 0xfe
      11'h49B: dout <= 8'b11111100; // 1179 : 252 - 0xfc
      11'h49C: dout <= 8'b11110000; // 1180 : 240 - 0xf0
      11'h49D: dout <= 8'b11000000; // 1181 : 192 - 0xc0
      11'h49E: dout <= 8'b00100000; // 1182 :  32 - 0x20
      11'h49F: dout <= 8'b11100000; // 1183 : 224 - 0xe0
      11'h4A0: dout <= 8'b00000011; // 1184 :   3 - 0x3 -- Background 0x94
      11'h4A1: dout <= 8'b00001111; // 1185 :  15 - 0xf
      11'h4A2: dout <= 8'b00010011; // 1186 :  19 - 0x13
      11'h4A3: dout <= 8'b00110001; // 1187 :  49 - 0x31
      11'h4A4: dout <= 8'b01111001; // 1188 : 121 - 0x79
      11'h4A5: dout <= 8'b01011001; // 1189 :  89 - 0x59
      11'h4A6: dout <= 8'b01001000; // 1190 :  72 - 0x48
      11'h4A7: dout <= 8'b11001100; // 1191 : 204 - 0xcc
      11'h4A8: dout <= 8'b10010101; // 1192 : 149 - 0x95 -- Background 0x95
      11'h4A9: dout <= 8'b11111111; // 1193 : 255 - 0xff
      11'h4AA: dout <= 8'b01111111; // 1194 : 127 - 0x7f
      11'h4AB: dout <= 8'b00111110; // 1195 :  62 - 0x3e
      11'h4AC: dout <= 8'b00011111; // 1196 :  31 - 0x1f
      11'h4AD: dout <= 8'b00001111; // 1197 :  15 - 0xf
      11'h4AE: dout <= 8'b00001111; // 1198 :  15 - 0xf
      11'h4AF: dout <= 8'b00000111; // 1199 :   7 - 0x7
      11'h4B0: dout <= 8'b11000000; // 1200 : 192 - 0xc0 -- Background 0x96
      11'h4B1: dout <= 8'b00110000; // 1201 :  48 - 0x30
      11'h4B2: dout <= 8'b00001000; // 1202 :   8 - 0x8
      11'h4B3: dout <= 8'b10010100; // 1203 : 148 - 0x94
      11'h4B4: dout <= 8'b10011010; // 1204 : 154 - 0x9a
      11'h4B5: dout <= 8'b00011010; // 1205 :  26 - 0x1a
      11'h4B6: dout <= 8'b00000001; // 1206 :   1 - 0x1
      11'h4B7: dout <= 8'b00001111; // 1207 :  15 - 0xf
      11'h4B8: dout <= 8'b01000101; // 1208 :  69 - 0x45 -- Background 0x97
      11'h4B9: dout <= 8'b11100001; // 1209 : 225 - 0xe1
      11'h4BA: dout <= 8'b11111110; // 1210 : 254 - 0xfe
      11'h4BB: dout <= 8'b01111100; // 1211 : 124 - 0x7c
      11'h4BC: dout <= 8'b00110000; // 1212 :  48 - 0x30
      11'h4BD: dout <= 8'b00110000; // 1213 :  48 - 0x30
      11'h4BE: dout <= 8'b10001000; // 1214 : 136 - 0x88
      11'h4BF: dout <= 8'b01111000; // 1215 : 120 - 0x78
      11'h4C0: dout <= 8'b00000001; // 1216 :   1 - 0x1 -- Background 0x98
      11'h4C1: dout <= 8'b00000000; // 1217 :   0 - 0x0
      11'h4C2: dout <= 8'b00000000; // 1218 :   0 - 0x0
      11'h4C3: dout <= 8'b00000000; // 1219 :   0 - 0x0
      11'h4C4: dout <= 8'b00000001; // 1220 :   1 - 0x1
      11'h4C5: dout <= 8'b00000001; // 1221 :   1 - 0x1
      11'h4C6: dout <= 8'b00000010; // 1222 :   2 - 0x2
      11'h4C7: dout <= 8'b00000110; // 1223 :   6 - 0x6
      11'h4C8: dout <= 8'b01111000; // 1224 : 120 - 0x78 -- Background 0x99
      11'h4C9: dout <= 8'b00101010; // 1225 :  42 - 0x2a
      11'h4CA: dout <= 8'b01010100; // 1226 :  84 - 0x54
      11'h4CB: dout <= 8'b00101001; // 1227 :  41 - 0x29
      11'h4CC: dout <= 8'b00101111; // 1228 :  47 - 0x2f
      11'h4CD: dout <= 8'b00110111; // 1229 :  55 - 0x37
      11'h4CE: dout <= 8'b00000011; // 1230 :   3 - 0x3
      11'h4CF: dout <= 8'b00000111; // 1231 :   7 - 0x7
      11'h4D0: dout <= 8'b10110000; // 1232 : 176 - 0xb0 -- Background 0x9a
      11'h4D1: dout <= 8'b11101000; // 1233 : 232 - 0xe8
      11'h4D2: dout <= 8'b10001100; // 1234 : 140 - 0x8c
      11'h4D3: dout <= 8'b10011110; // 1235 : 158 - 0x9e
      11'h4D4: dout <= 8'b00011111; // 1236 :  31 - 0x1f
      11'h4D5: dout <= 8'b00001111; // 1237 :  15 - 0xf
      11'h4D6: dout <= 8'b10010110; // 1238 : 150 - 0x96
      11'h4D7: dout <= 8'b00011100; // 1239 :  28 - 0x1c
      11'h4D8: dout <= 8'b00001100; // 1240 :  12 - 0xc -- Background 0x9b
      11'h4D9: dout <= 8'b00111000; // 1241 :  56 - 0x38
      11'h4DA: dout <= 8'b11101000; // 1242 : 232 - 0xe8
      11'h4DB: dout <= 8'b11010000; // 1243 : 208 - 0xd0
      11'h4DC: dout <= 8'b11100000; // 1244 : 224 - 0xe0
      11'h4DD: dout <= 8'b10000000; // 1245 : 128 - 0x80
      11'h4DE: dout <= 8'b00000000; // 1246 :   0 - 0x0
      11'h4DF: dout <= 8'b10000000; // 1247 : 128 - 0x80
      11'h4E0: dout <= 8'b00000001; // 1248 :   1 - 0x1 -- Background 0x9c
      11'h4E1: dout <= 8'b00000000; // 1249 :   0 - 0x0
      11'h4E2: dout <= 8'b00000000; // 1250 :   0 - 0x0
      11'h4E3: dout <= 8'b00000000; // 1251 :   0 - 0x0
      11'h4E4: dout <= 8'b00000001; // 1252 :   1 - 0x1
      11'h4E5: dout <= 8'b00000001; // 1253 :   1 - 0x1
      11'h4E6: dout <= 8'b00000010; // 1254 :   2 - 0x2
      11'h4E7: dout <= 8'b00000110; // 1255 :   6 - 0x6
      11'h4E8: dout <= 8'b01111000; // 1256 : 120 - 0x78 -- Background 0x9d
      11'h4E9: dout <= 8'b00101010; // 1257 :  42 - 0x2a
      11'h4EA: dout <= 8'b01010100; // 1258 :  84 - 0x54
      11'h4EB: dout <= 8'b00101001; // 1259 :  41 - 0x29
      11'h4EC: dout <= 8'b00101111; // 1260 :  47 - 0x2f
      11'h4ED: dout <= 8'b00111100; // 1261 :  60 - 0x3c
      11'h4EE: dout <= 8'b00011110; // 1262 :  30 - 0x1e
      11'h4EF: dout <= 8'b00000000; // 1263 :   0 - 0x0
      11'h4F0: dout <= 8'b10110000; // 1264 : 176 - 0xb0 -- Background 0x9e
      11'h4F1: dout <= 8'b11101000; // 1265 : 232 - 0xe8
      11'h4F2: dout <= 8'b10001100; // 1266 : 140 - 0x8c
      11'h4F3: dout <= 8'b10011110; // 1267 : 158 - 0x9e
      11'h4F4: dout <= 8'b00011111; // 1268 :  31 - 0x1f
      11'h4F5: dout <= 8'b00001111; // 1269 :  15 - 0xf
      11'h4F6: dout <= 8'b10010110; // 1270 : 150 - 0x96
      11'h4F7: dout <= 8'b00011100; // 1271 :  28 - 0x1c
      11'h4F8: dout <= 8'b00001100; // 1272 :  12 - 0xc -- Background 0x9f
      11'h4F9: dout <= 8'b00111000; // 1273 :  56 - 0x38
      11'h4FA: dout <= 8'b11101000; // 1274 : 232 - 0xe8
      11'h4FB: dout <= 8'b11110000; // 1275 : 240 - 0xf0
      11'h4FC: dout <= 8'b11000000; // 1276 : 192 - 0xc0
      11'h4FD: dout <= 8'b01110000; // 1277 : 112 - 0x70
      11'h4FE: dout <= 8'b11000000; // 1278 : 192 - 0xc0
      11'h4FF: dout <= 8'b00000000; // 1279 :   0 - 0x0
      11'h500: dout <= 8'b00000011; // 1280 :   3 - 0x3 -- Background 0xa0
      11'h501: dout <= 8'b00001111; // 1281 :  15 - 0xf
      11'h502: dout <= 8'b00011100; // 1282 :  28 - 0x1c
      11'h503: dout <= 8'b00110000; // 1283 :  48 - 0x30
      11'h504: dout <= 8'b01100000; // 1284 :  96 - 0x60
      11'h505: dout <= 8'b01100000; // 1285 :  96 - 0x60
      11'h506: dout <= 8'b11000000; // 1286 : 192 - 0xc0
      11'h507: dout <= 8'b11000000; // 1287 : 192 - 0xc0
      11'h508: dout <= 8'b11000000; // 1288 : 192 - 0xc0 -- Background 0xa1
      11'h509: dout <= 8'b11000000; // 1289 : 192 - 0xc0
      11'h50A: dout <= 8'b01100000; // 1290 :  96 - 0x60
      11'h50B: dout <= 8'b01100000; // 1291 :  96 - 0x60
      11'h50C: dout <= 8'b00110000; // 1292 :  48 - 0x30
      11'h50D: dout <= 8'b00011010; // 1293 :  26 - 0x1a
      11'h50E: dout <= 8'b00001101; // 1294 :  13 - 0xd
      11'h50F: dout <= 8'b00000011; // 1295 :   3 - 0x3
      11'h510: dout <= 8'b11000000; // 1296 : 192 - 0xc0 -- Background 0xa2
      11'h511: dout <= 8'b11110000; // 1297 : 240 - 0xf0
      11'h512: dout <= 8'b00111000; // 1298 :  56 - 0x38
      11'h513: dout <= 8'b00001100; // 1299 :  12 - 0xc
      11'h514: dout <= 8'b00000110; // 1300 :   6 - 0x6
      11'h515: dout <= 8'b00000010; // 1301 :   2 - 0x2
      11'h516: dout <= 8'b00000101; // 1302 :   5 - 0x5
      11'h517: dout <= 8'b00000011; // 1303 :   3 - 0x3
      11'h518: dout <= 8'b00000101; // 1304 :   5 - 0x5 -- Background 0xa3
      11'h519: dout <= 8'b00001011; // 1305 :  11 - 0xb
      11'h51A: dout <= 8'b00010110; // 1306 :  22 - 0x16
      11'h51B: dout <= 8'b00101010; // 1307 :  42 - 0x2a
      11'h51C: dout <= 8'b01010100; // 1308 :  84 - 0x54
      11'h51D: dout <= 8'b10101000; // 1309 : 168 - 0xa8
      11'h51E: dout <= 8'b01110000; // 1310 : 112 - 0x70
      11'h51F: dout <= 8'b11000000; // 1311 : 192 - 0xc0
      11'h520: dout <= 8'b00000000; // 1312 :   0 - 0x0 -- Background 0xa4
      11'h521: dout <= 8'b00001111; // 1313 :  15 - 0xf
      11'h522: dout <= 8'b00011111; // 1314 :  31 - 0x1f
      11'h523: dout <= 8'b00110001; // 1315 :  49 - 0x31
      11'h524: dout <= 8'b00111111; // 1316 :  63 - 0x3f
      11'h525: dout <= 8'b01111111; // 1317 : 127 - 0x7f
      11'h526: dout <= 8'b11111111; // 1318 : 255 - 0xff
      11'h527: dout <= 8'b11011111; // 1319 : 223 - 0xdf
      11'h528: dout <= 8'b11000000; // 1320 : 192 - 0xc0 -- Background 0xa5
      11'h529: dout <= 8'b11000111; // 1321 : 199 - 0xc7
      11'h52A: dout <= 8'b01101111; // 1322 : 111 - 0x6f
      11'h52B: dout <= 8'b01100111; // 1323 : 103 - 0x67
      11'h52C: dout <= 8'b01100011; // 1324 :  99 - 0x63
      11'h52D: dout <= 8'b00110000; // 1325 :  48 - 0x30
      11'h52E: dout <= 8'b00011000; // 1326 :  24 - 0x18
      11'h52F: dout <= 8'b00000111; // 1327 :   7 - 0x7
      11'h530: dout <= 8'b00000000; // 1328 :   0 - 0x0 -- Background 0xa6
      11'h531: dout <= 8'b11110000; // 1329 : 240 - 0xf0
      11'h532: dout <= 8'b11111000; // 1330 : 248 - 0xf8
      11'h533: dout <= 8'b10001100; // 1331 : 140 - 0x8c
      11'h534: dout <= 8'b11111100; // 1332 : 252 - 0xfc
      11'h535: dout <= 8'b11111110; // 1333 : 254 - 0xfe
      11'h536: dout <= 8'b11111101; // 1334 : 253 - 0xfd
      11'h537: dout <= 8'b11111001; // 1335 : 249 - 0xf9
      11'h538: dout <= 8'b00000011; // 1336 :   3 - 0x3 -- Background 0xa7
      11'h539: dout <= 8'b11100101; // 1337 : 229 - 0xe5
      11'h53A: dout <= 8'b11110010; // 1338 : 242 - 0xf2
      11'h53B: dout <= 8'b11100110; // 1339 : 230 - 0xe6
      11'h53C: dout <= 8'b11001010; // 1340 : 202 - 0xca
      11'h53D: dout <= 8'b00010100; // 1341 :  20 - 0x14
      11'h53E: dout <= 8'b00111000; // 1342 :  56 - 0x38
      11'h53F: dout <= 8'b11100000; // 1343 : 224 - 0xe0
      11'h540: dout <= 8'b00000000; // 1344 :   0 - 0x0 -- Background 0xa8
      11'h541: dout <= 8'b00001111; // 1345 :  15 - 0xf
      11'h542: dout <= 8'b00011111; // 1346 :  31 - 0x1f
      11'h543: dout <= 8'b00110001; // 1347 :  49 - 0x31
      11'h544: dout <= 8'b00111111; // 1348 :  63 - 0x3f
      11'h545: dout <= 8'b01111111; // 1349 : 127 - 0x7f
      11'h546: dout <= 8'b11111111; // 1350 : 255 - 0xff
      11'h547: dout <= 8'b11011111; // 1351 : 223 - 0xdf
      11'h548: dout <= 8'b11000000; // 1352 : 192 - 0xc0 -- Background 0xa9
      11'h549: dout <= 8'b11000011; // 1353 : 195 - 0xc3
      11'h54A: dout <= 8'b11000111; // 1354 : 199 - 0xc7
      11'h54B: dout <= 8'b11001111; // 1355 : 207 - 0xcf
      11'h54C: dout <= 8'b11000111; // 1356 : 199 - 0xc7
      11'h54D: dout <= 8'b11000000; // 1357 : 192 - 0xc0
      11'h54E: dout <= 8'b11100000; // 1358 : 224 - 0xe0
      11'h54F: dout <= 8'b11111111; // 1359 : 255 - 0xff
      11'h550: dout <= 8'b00000000; // 1360 :   0 - 0x0 -- Background 0xaa
      11'h551: dout <= 8'b11110000; // 1361 : 240 - 0xf0
      11'h552: dout <= 8'b11111000; // 1362 : 248 - 0xf8
      11'h553: dout <= 8'b10001100; // 1363 : 140 - 0x8c
      11'h554: dout <= 8'b11111100; // 1364 : 252 - 0xfc
      11'h555: dout <= 8'b11111110; // 1365 : 254 - 0xfe
      11'h556: dout <= 8'b11111101; // 1366 : 253 - 0xfd
      11'h557: dout <= 8'b11111001; // 1367 : 249 - 0xf9
      11'h558: dout <= 8'b00000011; // 1368 :   3 - 0x3 -- Background 0xab
      11'h559: dout <= 8'b11000101; // 1369 : 197 - 0xc5
      11'h55A: dout <= 8'b11100011; // 1370 : 227 - 0xe3
      11'h55B: dout <= 8'b11110101; // 1371 : 245 - 0xf5
      11'h55C: dout <= 8'b11100011; // 1372 : 227 - 0xe3
      11'h55D: dout <= 8'b00000101; // 1373 :   5 - 0x5
      11'h55E: dout <= 8'b00001011; // 1374 :  11 - 0xb
      11'h55F: dout <= 8'b11111111; // 1375 : 255 - 0xff
      11'h560: dout <= 8'b10000011; // 1376 : 131 - 0x83 -- Background 0xac
      11'h561: dout <= 8'b10001100; // 1377 : 140 - 0x8c
      11'h562: dout <= 8'b10010000; // 1378 : 144 - 0x90
      11'h563: dout <= 8'b10010000; // 1379 : 144 - 0x90
      11'h564: dout <= 8'b11100000; // 1380 : 224 - 0xe0
      11'h565: dout <= 8'b10100000; // 1381 : 160 - 0xa0
      11'h566: dout <= 8'b10101111; // 1382 : 175 - 0xaf
      11'h567: dout <= 8'b01101111; // 1383 : 111 - 0x6f
      11'h568: dout <= 8'b11111011; // 1384 : 251 - 0xfb -- Background 0xad
      11'h569: dout <= 8'b00000101; // 1385 :   5 - 0x5
      11'h56A: dout <= 8'b00000101; // 1386 :   5 - 0x5
      11'h56B: dout <= 8'b00000101; // 1387 :   5 - 0x5
      11'h56C: dout <= 8'b01000101; // 1388 :  69 - 0x45
      11'h56D: dout <= 8'b01100101; // 1389 : 101 - 0x65
      11'h56E: dout <= 8'b11110101; // 1390 : 245 - 0xf5
      11'h56F: dout <= 8'b11111101; // 1391 : 253 - 0xfd
      11'h570: dout <= 8'b10000011; // 1392 : 131 - 0x83 -- Background 0xae
      11'h571: dout <= 8'b10001100; // 1393 : 140 - 0x8c
      11'h572: dout <= 8'b10010000; // 1394 : 144 - 0x90
      11'h573: dout <= 8'b10010000; // 1395 : 144 - 0x90
      11'h574: dout <= 8'b11100000; // 1396 : 224 - 0xe0
      11'h575: dout <= 8'b10100000; // 1397 : 160 - 0xa0
      11'h576: dout <= 8'b10101111; // 1398 : 175 - 0xaf
      11'h577: dout <= 8'b01101111; // 1399 : 111 - 0x6f
      11'h578: dout <= 8'b11111011; // 1400 : 251 - 0xfb -- Background 0xaf
      11'h579: dout <= 8'b00000101; // 1401 :   5 - 0x5
      11'h57A: dout <= 8'b00000101; // 1402 :   5 - 0x5
      11'h57B: dout <= 8'b00000101; // 1403 :   5 - 0x5
      11'h57C: dout <= 8'b11000101; // 1404 : 197 - 0xc5
      11'h57D: dout <= 8'b11100101; // 1405 : 229 - 0xe5
      11'h57E: dout <= 8'b11110101; // 1406 : 245 - 0xf5
      11'h57F: dout <= 8'b11111101; // 1407 : 253 - 0xfd
      11'h580: dout <= 8'b00000000; // 1408 :   0 - 0x0 -- Background 0xb0
      11'h581: dout <= 8'b00000011; // 1409 :   3 - 0x3
      11'h582: dout <= 8'b00001111; // 1410 :  15 - 0xf
      11'h583: dout <= 8'b00111111; // 1411 :  63 - 0x3f
      11'h584: dout <= 8'b01111111; // 1412 : 127 - 0x7f
      11'h585: dout <= 8'b01111111; // 1413 : 127 - 0x7f
      11'h586: dout <= 8'b11111111; // 1414 : 255 - 0xff
      11'h587: dout <= 8'b11111111; // 1415 : 255 - 0xff
      11'h588: dout <= 8'b11111111; // 1416 : 255 - 0xff -- Background 0xb1
      11'h589: dout <= 8'b10001111; // 1417 : 143 - 0x8f
      11'h58A: dout <= 8'b10000000; // 1418 : 128 - 0x80
      11'h58B: dout <= 8'b11110000; // 1419 : 240 - 0xf0
      11'h58C: dout <= 8'b11111111; // 1420 : 255 - 0xff
      11'h58D: dout <= 8'b11111111; // 1421 : 255 - 0xff
      11'h58E: dout <= 8'b01111111; // 1422 : 127 - 0x7f
      11'h58F: dout <= 8'b00001111; // 1423 :  15 - 0xf
      11'h590: dout <= 8'b00000000; // 1424 :   0 - 0x0 -- Background 0xb2
      11'h591: dout <= 8'b11000000; // 1425 : 192 - 0xc0
      11'h592: dout <= 8'b11110000; // 1426 : 240 - 0xf0
      11'h593: dout <= 8'b11111100; // 1427 : 252 - 0xfc
      11'h594: dout <= 8'b11111110; // 1428 : 254 - 0xfe
      11'h595: dout <= 8'b11111110; // 1429 : 254 - 0xfe
      11'h596: dout <= 8'b11111111; // 1430 : 255 - 0xff
      11'h597: dout <= 8'b11111111; // 1431 : 255 - 0xff
      11'h598: dout <= 8'b11111111; // 1432 : 255 - 0xff -- Background 0xb3
      11'h599: dout <= 8'b11110001; // 1433 : 241 - 0xf1
      11'h59A: dout <= 8'b00000001; // 1434 :   1 - 0x1
      11'h59B: dout <= 8'b00001111; // 1435 :  15 - 0xf
      11'h59C: dout <= 8'b11111111; // 1436 : 255 - 0xff
      11'h59D: dout <= 8'b11111111; // 1437 : 255 - 0xff
      11'h59E: dout <= 8'b11111110; // 1438 : 254 - 0xfe
      11'h59F: dout <= 8'b11110000; // 1439 : 240 - 0xf0
      11'h5A0: dout <= 8'b00000000; // 1440 :   0 - 0x0 -- Background 0xb4
      11'h5A1: dout <= 8'b00000011; // 1441 :   3 - 0x3
      11'h5A2: dout <= 8'b00001110; // 1442 :  14 - 0xe
      11'h5A3: dout <= 8'b00110101; // 1443 :  53 - 0x35
      11'h5A4: dout <= 8'b01101110; // 1444 : 110 - 0x6e
      11'h5A5: dout <= 8'b01010101; // 1445 :  85 - 0x55
      11'h5A6: dout <= 8'b10111010; // 1446 : 186 - 0xba
      11'h5A7: dout <= 8'b11010111; // 1447 : 215 - 0xd7
      11'h5A8: dout <= 8'b11111010; // 1448 : 250 - 0xfa -- Background 0xb5
      11'h5A9: dout <= 8'b10001111; // 1449 : 143 - 0x8f
      11'h5AA: dout <= 8'b10000000; // 1450 : 128 - 0x80
      11'h5AB: dout <= 8'b11110000; // 1451 : 240 - 0xf0
      11'h5AC: dout <= 8'b10101111; // 1452 : 175 - 0xaf
      11'h5AD: dout <= 8'b11010101; // 1453 : 213 - 0xd5
      11'h5AE: dout <= 8'b01111010; // 1454 : 122 - 0x7a
      11'h5AF: dout <= 8'b00001111; // 1455 :  15 - 0xf
      11'h5B0: dout <= 8'b00000000; // 1456 :   0 - 0x0 -- Background 0xb6
      11'h5B1: dout <= 8'b11000000; // 1457 : 192 - 0xc0
      11'h5B2: dout <= 8'b10110000; // 1458 : 176 - 0xb0
      11'h5B3: dout <= 8'b01011100; // 1459 :  92 - 0x5c
      11'h5B4: dout <= 8'b11101010; // 1460 : 234 - 0xea
      11'h5B5: dout <= 8'b01011110; // 1461 :  94 - 0x5e
      11'h5B6: dout <= 8'b10101011; // 1462 : 171 - 0xab
      11'h5B7: dout <= 8'b01110101; // 1463 : 117 - 0x75
      11'h5B8: dout <= 8'b10101111; // 1464 : 175 - 0xaf -- Background 0xb7
      11'h5B9: dout <= 8'b11110001; // 1465 : 241 - 0xf1
      11'h5BA: dout <= 8'b00000001; // 1466 :   1 - 0x1
      11'h5BB: dout <= 8'b00001111; // 1467 :  15 - 0xf
      11'h5BC: dout <= 8'b11111011; // 1468 : 251 - 0xfb
      11'h5BD: dout <= 8'b01010101; // 1469 :  85 - 0x55
      11'h5BE: dout <= 8'b10101110; // 1470 : 174 - 0xae
      11'h5BF: dout <= 8'b11110000; // 1471 : 240 - 0xf0
      11'h5C0: dout <= 8'b00000000; // 1472 :   0 - 0x0 -- Background 0xb8
      11'h5C1: dout <= 8'b00000011; // 1473 :   3 - 0x3
      11'h5C2: dout <= 8'b00001100; // 1474 :  12 - 0xc
      11'h5C3: dout <= 8'b00110000; // 1475 :  48 - 0x30
      11'h5C4: dout <= 8'b01000100; // 1476 :  68 - 0x44
      11'h5C5: dout <= 8'b01000000; // 1477 :  64 - 0x40
      11'h5C6: dout <= 8'b10010000; // 1478 : 144 - 0x90
      11'h5C7: dout <= 8'b10000010; // 1479 : 130 - 0x82
      11'h5C8: dout <= 8'b11110000; // 1480 : 240 - 0xf0 -- Background 0xb9
      11'h5C9: dout <= 8'b11111111; // 1481 : 255 - 0xff
      11'h5CA: dout <= 8'b11111111; // 1482 : 255 - 0xff
      11'h5CB: dout <= 8'b11111111; // 1483 : 255 - 0xff
      11'h5CC: dout <= 8'b10001111; // 1484 : 143 - 0x8f
      11'h5CD: dout <= 8'b10000000; // 1485 : 128 - 0x80
      11'h5CE: dout <= 8'b01110000; // 1486 : 112 - 0x70
      11'h5CF: dout <= 8'b00001111; // 1487 :  15 - 0xf
      11'h5D0: dout <= 8'b00000000; // 1488 :   0 - 0x0 -- Background 0xba
      11'h5D1: dout <= 8'b11000000; // 1489 : 192 - 0xc0
      11'h5D2: dout <= 8'b00110000; // 1490 :  48 - 0x30
      11'h5D3: dout <= 8'b00001100; // 1491 :  12 - 0xc
      11'h5D4: dout <= 8'b01000010; // 1492 :  66 - 0x42
      11'h5D5: dout <= 8'b00001010; // 1493 :  10 - 0xa
      11'h5D6: dout <= 8'b00000001; // 1494 :   1 - 0x1
      11'h5D7: dout <= 8'b00100001; // 1495 :  33 - 0x21
      11'h5D8: dout <= 8'b00001111; // 1496 :  15 - 0xf -- Background 0xbb
      11'h5D9: dout <= 8'b11111111; // 1497 : 255 - 0xff
      11'h5DA: dout <= 8'b11111111; // 1498 : 255 - 0xff
      11'h5DB: dout <= 8'b11111111; // 1499 : 255 - 0xff
      11'h5DC: dout <= 8'b11110001; // 1500 : 241 - 0xf1
      11'h5DD: dout <= 8'b00000001; // 1501 :   1 - 0x1
      11'h5DE: dout <= 8'b00001110; // 1502 :  14 - 0xe
      11'h5DF: dout <= 8'b11110000; // 1503 : 240 - 0xf0
      11'h5E0: dout <= 8'b11110011; // 1504 : 243 - 0xf3 -- Background 0xbc
      11'h5E1: dout <= 8'b11111111; // 1505 : 255 - 0xff
      11'h5E2: dout <= 8'b11000100; // 1506 : 196 - 0xc4
      11'h5E3: dout <= 8'b11000000; // 1507 : 192 - 0xc0
      11'h5E4: dout <= 8'b01000000; // 1508 :  64 - 0x40
      11'h5E5: dout <= 8'b01100011; // 1509 :  99 - 0x63
      11'h5E6: dout <= 8'b11000111; // 1510 : 199 - 0xc7
      11'h5E7: dout <= 8'b11000110; // 1511 : 198 - 0xc6
      11'h5E8: dout <= 8'b11000110; // 1512 : 198 - 0xc6 -- Background 0xbd
      11'h5E9: dout <= 8'b11000110; // 1513 : 198 - 0xc6
      11'h5EA: dout <= 8'b01100011; // 1514 :  99 - 0x63
      11'h5EB: dout <= 8'b01000000; // 1515 :  64 - 0x40
      11'h5EC: dout <= 8'b11000000; // 1516 : 192 - 0xc0
      11'h5ED: dout <= 8'b11000100; // 1517 : 196 - 0xc4
      11'h5EE: dout <= 8'b11001100; // 1518 : 204 - 0xcc
      11'h5EF: dout <= 8'b11110011; // 1519 : 243 - 0xf3
      11'h5F0: dout <= 8'b11001111; // 1520 : 207 - 0xcf -- Background 0xbe
      11'h5F1: dout <= 8'b11111111; // 1521 : 255 - 0xff
      11'h5F2: dout <= 8'b00100001; // 1522 :  33 - 0x21
      11'h5F3: dout <= 8'b00000001; // 1523 :   1 - 0x1
      11'h5F4: dout <= 8'b00000010; // 1524 :   2 - 0x2
      11'h5F5: dout <= 8'b11000110; // 1525 : 198 - 0xc6
      11'h5F6: dout <= 8'b11100001; // 1526 : 225 - 0xe1
      11'h5F7: dout <= 8'b00100001; // 1527 :  33 - 0x21
      11'h5F8: dout <= 8'b00100001; // 1528 :  33 - 0x21 -- Background 0xbf
      11'h5F9: dout <= 8'b00100001; // 1529 :  33 - 0x21
      11'h5FA: dout <= 8'b11000110; // 1530 : 198 - 0xc6
      11'h5FB: dout <= 8'b00000010; // 1531 :   2 - 0x2
      11'h5FC: dout <= 8'b00000001; // 1532 :   1 - 0x1
      11'h5FD: dout <= 8'b00100001; // 1533 :  33 - 0x21
      11'h5FE: dout <= 8'b00110001; // 1534 :  49 - 0x31
      11'h5FF: dout <= 8'b11001111; // 1535 : 207 - 0xcf
      11'h600: dout <= 8'b00000000; // 1536 :   0 - 0x0 -- Background 0xc0
      11'h601: dout <= 8'b01010000; // 1537 :  80 - 0x50
      11'h602: dout <= 8'b10110011; // 1538 : 179 - 0xb3
      11'h603: dout <= 8'b10010111; // 1539 : 151 - 0x97
      11'h604: dout <= 8'b10011111; // 1540 : 159 - 0x9f
      11'h605: dout <= 8'b01101111; // 1541 : 111 - 0x6f
      11'h606: dout <= 8'b00011111; // 1542 :  31 - 0x1f
      11'h607: dout <= 8'b00011111; // 1543 :  31 - 0x1f
      11'h608: dout <= 8'b00011111; // 1544 :  31 - 0x1f -- Background 0xc1
      11'h609: dout <= 8'b00011111; // 1545 :  31 - 0x1f
      11'h60A: dout <= 8'b00001111; // 1546 :  15 - 0xf
      11'h60B: dout <= 8'b00000111; // 1547 :   7 - 0x7
      11'h60C: dout <= 8'b00011101; // 1548 :  29 - 0x1d
      11'h60D: dout <= 8'b00101100; // 1549 :  44 - 0x2c
      11'h60E: dout <= 8'b01010100; // 1550 :  84 - 0x54
      11'h60F: dout <= 8'b01111100; // 1551 : 124 - 0x7c
      11'h610: dout <= 8'b00000000; // 1552 :   0 - 0x0 -- Background 0xc2
      11'h611: dout <= 8'b00001010; // 1553 :  10 - 0xa
      11'h612: dout <= 8'b11001101; // 1554 : 205 - 0xcd
      11'h613: dout <= 8'b11101001; // 1555 : 233 - 0xe9
      11'h614: dout <= 8'b11111001; // 1556 : 249 - 0xf9
      11'h615: dout <= 8'b11110110; // 1557 : 246 - 0xf6
      11'h616: dout <= 8'b11110000; // 1558 : 240 - 0xf0
      11'h617: dout <= 8'b11111000; // 1559 : 248 - 0xf8
      11'h618: dout <= 8'b11111000; // 1560 : 248 - 0xf8 -- Background 0xc3
      11'h619: dout <= 8'b11111000; // 1561 : 248 - 0xf8
      11'h61A: dout <= 8'b11110000; // 1562 : 240 - 0xf0
      11'h61B: dout <= 8'b11000000; // 1563 : 192 - 0xc0
      11'h61C: dout <= 8'b10111000; // 1564 : 184 - 0xb8
      11'h61D: dout <= 8'b00110100; // 1565 :  52 - 0x34
      11'h61E: dout <= 8'b00101010; // 1566 :  42 - 0x2a
      11'h61F: dout <= 8'b00111110; // 1567 :  62 - 0x3e
      11'h620: dout <= 8'b00000101; // 1568 :   5 - 0x5 -- Background 0xc4
      11'h621: dout <= 8'b00001010; // 1569 :  10 - 0xa
      11'h622: dout <= 8'b00001000; // 1570 :   8 - 0x8
      11'h623: dout <= 8'b00001111; // 1571 :  15 - 0xf
      11'h624: dout <= 8'b00000001; // 1572 :   1 - 0x1
      11'h625: dout <= 8'b00000011; // 1573 :   3 - 0x3
      11'h626: dout <= 8'b00000111; // 1574 :   7 - 0x7
      11'h627: dout <= 8'b00001111; // 1575 :  15 - 0xf
      11'h628: dout <= 8'b00001111; // 1576 :  15 - 0xf -- Background 0xc5
      11'h629: dout <= 8'b11101111; // 1577 : 239 - 0xef
      11'h62A: dout <= 8'b11011111; // 1578 : 223 - 0xdf
      11'h62B: dout <= 8'b10101111; // 1579 : 175 - 0xaf
      11'h62C: dout <= 8'b01100111; // 1580 : 103 - 0x67
      11'h62D: dout <= 8'b00001101; // 1581 :  13 - 0xd
      11'h62E: dout <= 8'b00001010; // 1582 :  10 - 0xa
      11'h62F: dout <= 8'b00000111; // 1583 :   7 - 0x7
      11'h630: dout <= 8'b00000000; // 1584 :   0 - 0x0 -- Background 0xc6
      11'h631: dout <= 8'b10000000; // 1585 : 128 - 0x80
      11'h632: dout <= 8'b10000000; // 1586 : 128 - 0x80
      11'h633: dout <= 8'b11110000; // 1587 : 240 - 0xf0
      11'h634: dout <= 8'b11111000; // 1588 : 248 - 0xf8
      11'h635: dout <= 8'b11111100; // 1589 : 252 - 0xfc
      11'h636: dout <= 8'b11111100; // 1590 : 252 - 0xfc
      11'h637: dout <= 8'b11111100; // 1591 : 252 - 0xfc
      11'h638: dout <= 8'b11111100; // 1592 : 252 - 0xfc -- Background 0xc7
      11'h639: dout <= 8'b11111110; // 1593 : 254 - 0xfe
      11'h63A: dout <= 8'b11111001; // 1594 : 249 - 0xf9
      11'h63B: dout <= 8'b11111010; // 1595 : 250 - 0xfa
      11'h63C: dout <= 8'b11101001; // 1596 : 233 - 0xe9
      11'h63D: dout <= 8'b00001110; // 1597 :  14 - 0xe
      11'h63E: dout <= 8'b10000000; // 1598 : 128 - 0x80
      11'h63F: dout <= 8'b00000000; // 1599 :   0 - 0x0
      11'h640: dout <= 8'b00000000; // 1600 :   0 - 0x0 -- Background 0xc8
      11'h641: dout <= 8'b11000000; // 1601 : 192 - 0xc0
      11'h642: dout <= 8'b10100000; // 1602 : 160 - 0xa0
      11'h643: dout <= 8'b11010011; // 1603 : 211 - 0xd3
      11'h644: dout <= 8'b10110111; // 1604 : 183 - 0xb7
      11'h645: dout <= 8'b11111111; // 1605 : 255 - 0xff
      11'h646: dout <= 8'b00001111; // 1606 :  15 - 0xf
      11'h647: dout <= 8'b00011111; // 1607 :  31 - 0x1f
      11'h648: dout <= 8'b00011111; // 1608 :  31 - 0x1f -- Background 0xc9
      11'h649: dout <= 8'b00001111; // 1609 :  15 - 0xf
      11'h64A: dout <= 8'b11110111; // 1610 : 247 - 0xf7
      11'h64B: dout <= 8'b10110111; // 1611 : 183 - 0xb7
      11'h64C: dout <= 8'b11010011; // 1612 : 211 - 0xd3
      11'h64D: dout <= 8'b10100000; // 1613 : 160 - 0xa0
      11'h64E: dout <= 8'b11000000; // 1614 : 192 - 0xc0
      11'h64F: dout <= 8'b00000000; // 1615 :   0 - 0x0
      11'h650: dout <= 8'b00011100; // 1616 :  28 - 0x1c -- Background 0xca
      11'h651: dout <= 8'b00100010; // 1617 :  34 - 0x22
      11'h652: dout <= 8'b00100100; // 1618 :  36 - 0x24
      11'h653: dout <= 8'b11011110; // 1619 : 222 - 0xde
      11'h654: dout <= 8'b11110000; // 1620 : 240 - 0xf0
      11'h655: dout <= 8'b11111000; // 1621 : 248 - 0xf8
      11'h656: dout <= 8'b11111100; // 1622 : 252 - 0xfc
      11'h657: dout <= 8'b11111100; // 1623 : 252 - 0xfc
      11'h658: dout <= 8'b11111100; // 1624 : 252 - 0xfc -- Background 0xcb
      11'h659: dout <= 8'b11111100; // 1625 : 252 - 0xfc
      11'h65A: dout <= 8'b11111000; // 1626 : 248 - 0xf8
      11'h65B: dout <= 8'b11110000; // 1627 : 240 - 0xf0
      11'h65C: dout <= 8'b10011110; // 1628 : 158 - 0x9e
      11'h65D: dout <= 8'b00100100; // 1629 :  36 - 0x24
      11'h65E: dout <= 8'b00100010; // 1630 :  34 - 0x22
      11'h65F: dout <= 8'b00011100; // 1631 :  28 - 0x1c
      11'h660: dout <= 8'b00001110; // 1632 :  14 - 0xe -- Background 0xcc
      11'h661: dout <= 8'b00010110; // 1633 :  22 - 0x16
      11'h662: dout <= 8'b00011010; // 1634 :  26 - 0x1a
      11'h663: dout <= 8'b00000100; // 1635 :   4 - 0x4
      11'h664: dout <= 8'b01101111; // 1636 : 111 - 0x6f
      11'h665: dout <= 8'b10111111; // 1637 : 191 - 0xbf
      11'h666: dout <= 8'b11011111; // 1638 : 223 - 0xdf
      11'h667: dout <= 8'b10111111; // 1639 : 191 - 0xbf
      11'h668: dout <= 8'b01011111; // 1640 :  95 - 0x5f -- Background 0xcd
      11'h669: dout <= 8'b00011111; // 1641 :  31 - 0x1f
      11'h66A: dout <= 8'b00011111; // 1642 :  31 - 0x1f
      11'h66B: dout <= 8'b00001111; // 1643 :  15 - 0xf
      11'h66C: dout <= 8'b00111111; // 1644 :  63 - 0x3f
      11'h66D: dout <= 8'b00100011; // 1645 :  35 - 0x23
      11'h66E: dout <= 8'b00101010; // 1646 :  42 - 0x2a
      11'h66F: dout <= 8'b00010100; // 1647 :  20 - 0x14
      11'h670: dout <= 8'b00000000; // 1648 :   0 - 0x0 -- Background 0xce
      11'h671: dout <= 8'b00000000; // 1649 :   0 - 0x0
      11'h672: dout <= 8'b00000000; // 1650 :   0 - 0x0
      11'h673: dout <= 8'b00000000; // 1651 :   0 - 0x0
      11'h674: dout <= 8'b10001110; // 1652 : 142 - 0x8e
      11'h675: dout <= 8'b11001001; // 1653 : 201 - 0xc9
      11'h676: dout <= 8'b11101010; // 1654 : 234 - 0xea
      11'h677: dout <= 8'b11111001; // 1655 : 249 - 0xf9
      11'h678: dout <= 8'b11111110; // 1656 : 254 - 0xfe -- Background 0xcf
      11'h679: dout <= 8'b11111000; // 1657 : 248 - 0xf8
      11'h67A: dout <= 8'b11111000; // 1658 : 248 - 0xf8
      11'h67B: dout <= 8'b11111000; // 1659 : 248 - 0xf8
      11'h67C: dout <= 8'b11110000; // 1660 : 240 - 0xf0
      11'h67D: dout <= 8'b11100000; // 1661 : 224 - 0xe0
      11'h67E: dout <= 8'b00000000; // 1662 :   0 - 0x0
      11'h67F: dout <= 8'b00000000; // 1663 :   0 - 0x0
      11'h680: dout <= 8'b00000000; // 1664 :   0 - 0x0 -- Background 0xd0
      11'h681: dout <= 8'b00000000; // 1665 :   0 - 0x0
      11'h682: dout <= 8'b00000100; // 1666 :   4 - 0x4
      11'h683: dout <= 8'b00100110; // 1667 :  38 - 0x26
      11'h684: dout <= 8'b00101011; // 1668 :  43 - 0x2b
      11'h685: dout <= 8'b01110001; // 1669 : 113 - 0x71
      11'h686: dout <= 8'b01000000; // 1670 :  64 - 0x40
      11'h687: dout <= 8'b01000111; // 1671 :  71 - 0x47
      11'h688: dout <= 8'b10001111; // 1672 : 143 - 0x8f -- Background 0xd1
      11'h689: dout <= 8'b10001111; // 1673 : 143 - 0x8f
      11'h68A: dout <= 8'b01001111; // 1674 :  79 - 0x4f
      11'h68B: dout <= 8'b01001111; // 1675 :  79 - 0x4f
      11'h68C: dout <= 8'b00111111; // 1676 :  63 - 0x3f
      11'h68D: dout <= 8'b00010011; // 1677 :  19 - 0x13
      11'h68E: dout <= 8'b00010001; // 1678 :  17 - 0x11
      11'h68F: dout <= 8'b00011111; // 1679 :  31 - 0x1f
      11'h690: dout <= 8'b00000000; // 1680 :   0 - 0x0 -- Background 0xd2
      11'h691: dout <= 8'b10000000; // 1681 : 128 - 0x80
      11'h692: dout <= 8'b11001000; // 1682 : 200 - 0xc8
      11'h693: dout <= 8'b11010100; // 1683 : 212 - 0xd4
      11'h694: dout <= 8'b00100100; // 1684 :  36 - 0x24
      11'h695: dout <= 8'b00000010; // 1685 :   2 - 0x2
      11'h696: dout <= 8'b00000010; // 1686 :   2 - 0x2
      11'h697: dout <= 8'b11110010; // 1687 : 242 - 0xf2
      11'h698: dout <= 8'b11110010; // 1688 : 242 - 0xf2 -- Background 0xd3
      11'h699: dout <= 8'b11110010; // 1689 : 242 - 0xf2
      11'h69A: dout <= 8'b11110100; // 1690 : 244 - 0xf4
      11'h69B: dout <= 8'b11110100; // 1691 : 244 - 0xf4
      11'h69C: dout <= 8'b11110100; // 1692 : 244 - 0xf4
      11'h69D: dout <= 8'b11001000; // 1693 : 200 - 0xc8
      11'h69E: dout <= 8'b01000100; // 1694 :  68 - 0x44
      11'h69F: dout <= 8'b01111100; // 1695 : 124 - 0x7c
      11'h6A0: dout <= 8'b00000000; // 1696 :   0 - 0x0 -- Background 0xd4
      11'h6A1: dout <= 8'b00000000; // 1697 :   0 - 0x0
      11'h6A2: dout <= 8'b00000000; // 1698 :   0 - 0x0
      11'h6A3: dout <= 8'b00001001; // 1699 :   9 - 0x9
      11'h6A4: dout <= 8'b00011010; // 1700 :  26 - 0x1a
      11'h6A5: dout <= 8'b00010100; // 1701 :  20 - 0x14
      11'h6A6: dout <= 8'b00100000; // 1702 :  32 - 0x20
      11'h6A7: dout <= 8'b01000111; // 1703 :  71 - 0x47
      11'h6A8: dout <= 8'b10001111; // 1704 : 143 - 0x8f -- Background 0xd5
      11'h6A9: dout <= 8'b10001111; // 1705 : 143 - 0x8f
      11'h6AA: dout <= 8'b01001111; // 1706 :  79 - 0x4f
      11'h6AB: dout <= 8'b01001111; // 1707 :  79 - 0x4f
      11'h6AC: dout <= 8'b00111111; // 1708 :  63 - 0x3f
      11'h6AD: dout <= 8'b01000111; // 1709 :  71 - 0x47
      11'h6AE: dout <= 8'b00100010; // 1710 :  34 - 0x22
      11'h6AF: dout <= 8'b00011100; // 1711 :  28 - 0x1c
      11'h6B0: dout <= 8'b00000000; // 1712 :   0 - 0x0 -- Background 0xd6
      11'h6B1: dout <= 8'b01000000; // 1713 :  64 - 0x40
      11'h6B2: dout <= 8'b11000000; // 1714 : 192 - 0xc0
      11'h6B3: dout <= 8'b00101100; // 1715 :  44 - 0x2c
      11'h6B4: dout <= 8'b00110100; // 1716 :  52 - 0x34
      11'h6B5: dout <= 8'b00000100; // 1717 :   4 - 0x4
      11'h6B6: dout <= 8'b00000010; // 1718 :   2 - 0x2
      11'h6B7: dout <= 8'b11110010; // 1719 : 242 - 0xf2
      11'h6B8: dout <= 8'b11110010; // 1720 : 242 - 0xf2 -- Background 0xd7
      11'h6B9: dout <= 8'b11110010; // 1721 : 242 - 0xf2
      11'h6BA: dout <= 8'b11110100; // 1722 : 244 - 0xf4
      11'h6BB: dout <= 8'b11110111; // 1723 : 247 - 0xf7
      11'h6BC: dout <= 8'b11111101; // 1724 : 253 - 0xfd
      11'h6BD: dout <= 8'b11100001; // 1725 : 225 - 0xe1
      11'h6BE: dout <= 8'b00010010; // 1726 :  18 - 0x12
      11'h6BF: dout <= 8'b00001100; // 1727 :  12 - 0xc
      11'h6C0: dout <= 8'b01111000; // 1728 : 120 - 0x78 -- Background 0xd8
      11'h6C1: dout <= 8'b01001110; // 1729 :  78 - 0x4e
      11'h6C2: dout <= 8'b11000010; // 1730 : 194 - 0xc2
      11'h6C3: dout <= 8'b10011010; // 1731 : 154 - 0x9a
      11'h6C4: dout <= 8'b10011011; // 1732 : 155 - 0x9b
      11'h6C5: dout <= 8'b11011001; // 1733 : 217 - 0xd9
      11'h6C6: dout <= 8'b01100011; // 1734 :  99 - 0x63
      11'h6C7: dout <= 8'b00111110; // 1735 :  62 - 0x3e
      11'h6C8: dout <= 8'b00011110; // 1736 :  30 - 0x1e -- Background 0xd9
      11'h6C9: dout <= 8'b01110001; // 1737 : 113 - 0x71
      11'h6CA: dout <= 8'b01001001; // 1738 :  73 - 0x49
      11'h6CB: dout <= 8'b10111001; // 1739 : 185 - 0xb9
      11'h6CC: dout <= 8'b10011101; // 1740 : 157 - 0x9d
      11'h6CD: dout <= 8'b01010010; // 1741 :  82 - 0x52
      11'h6CE: dout <= 8'b01110010; // 1742 : 114 - 0x72
      11'h6CF: dout <= 8'b00011110; // 1743 :  30 - 0x1e
      11'h6D0: dout <= 8'b01100000; // 1744 :  96 - 0x60 -- Background 0xda
      11'h6D1: dout <= 8'b01011110; // 1745 :  94 - 0x5e
      11'h6D2: dout <= 8'b10001001; // 1746 : 137 - 0x89
      11'h6D3: dout <= 8'b10111101; // 1747 : 189 - 0xbd
      11'h6D4: dout <= 8'b10011101; // 1748 : 157 - 0x9d
      11'h6D5: dout <= 8'b11010011; // 1749 : 211 - 0xd3
      11'h6D6: dout <= 8'b01000110; // 1750 :  70 - 0x46
      11'h6D7: dout <= 8'b01111100; // 1751 : 124 - 0x7c
      11'h6D8: dout <= 8'b00011110; // 1752 :  30 - 0x1e -- Background 0xdb
      11'h6D9: dout <= 8'b00100011; // 1753 :  35 - 0x23
      11'h6DA: dout <= 8'b01001001; // 1754 :  73 - 0x49
      11'h6DB: dout <= 8'b10111101; // 1755 : 189 - 0xbd
      11'h6DC: dout <= 8'b10011001; // 1756 : 153 - 0x99
      11'h6DD: dout <= 8'b01000011; // 1757 :  67 - 0x43
      11'h6DE: dout <= 8'b01101110; // 1758 : 110 - 0x6e
      11'h6DF: dout <= 8'b00011000; // 1759 :  24 - 0x18
      11'h6E0: dout <= 8'b00000000; // 1760 :   0 - 0x0 -- Background 0xdc
      11'h6E1: dout <= 8'b00000000; // 1761 :   0 - 0x0
      11'h6E2: dout <= 8'b00000001; // 1762 :   1 - 0x1
      11'h6E3: dout <= 8'b00000010; // 1763 :   2 - 0x2
      11'h6E4: dout <= 8'b00000100; // 1764 :   4 - 0x4
      11'h6E5: dout <= 8'b00000010; // 1765 :   2 - 0x2
      11'h6E6: dout <= 8'b00011110; // 1766 :  30 - 0x1e
      11'h6E7: dout <= 8'b00010000; // 1767 :  16 - 0x10
      11'h6E8: dout <= 8'b00001000; // 1768 :   8 - 0x8 -- Background 0xdd
      11'h6E9: dout <= 8'b00001101; // 1769 :  13 - 0xd
      11'h6EA: dout <= 8'b00111010; // 1770 :  58 - 0x3a
      11'h6EB: dout <= 8'b00100101; // 1771 :  37 - 0x25
      11'h6EC: dout <= 8'b00011011; // 1772 :  27 - 0x1b
      11'h6ED: dout <= 8'b00001111; // 1773 :  15 - 0xf
      11'h6EE: dout <= 8'b00000111; // 1774 :   7 - 0x7
      11'h6EF: dout <= 8'b00000011; // 1775 :   3 - 0x3
      11'h6F0: dout <= 8'b00000000; // 1776 :   0 - 0x0 -- Background 0xde
      11'h6F1: dout <= 8'b00000000; // 1777 :   0 - 0x0
      11'h6F2: dout <= 8'b00000000; // 1778 :   0 - 0x0
      11'h6F3: dout <= 8'b11000000; // 1779 : 192 - 0xc0
      11'h6F4: dout <= 8'b01000000; // 1780 :  64 - 0x40
      11'h6F5: dout <= 8'b01011000; // 1781 :  88 - 0x58
      11'h6F6: dout <= 8'b01101000; // 1782 : 104 - 0x68
      11'h6F7: dout <= 8'b00001000; // 1783 :   8 - 0x8
      11'h6F8: dout <= 8'b00010000; // 1784 :  16 - 0x10 -- Background 0xdf
      11'h6F9: dout <= 8'b01011100; // 1785 :  92 - 0x5c
      11'h6FA: dout <= 8'b10101000; // 1786 : 168 - 0xa8
      11'h6FB: dout <= 8'b11011000; // 1787 : 216 - 0xd8
      11'h6FC: dout <= 8'b10111000; // 1788 : 184 - 0xb8
      11'h6FD: dout <= 8'b11110000; // 1789 : 240 - 0xf0
      11'h6FE: dout <= 8'b11100000; // 1790 : 224 - 0xe0
      11'h6FF: dout <= 8'b11000000; // 1791 : 192 - 0xc0
      11'h700: dout <= 8'b00000000; // 1792 :   0 - 0x0 -- Background 0xe0
      11'h701: dout <= 8'b00000000; // 1793 :   0 - 0x0
      11'h702: dout <= 8'b00000000; // 1794 :   0 - 0x0
      11'h703: dout <= 8'b00010011; // 1795 :  19 - 0x13
      11'h704: dout <= 8'b00010011; // 1796 :  19 - 0x13
      11'h705: dout <= 8'b00110111; // 1797 :  55 - 0x37
      11'h706: dout <= 8'b00110111; // 1798 :  55 - 0x37
      11'h707: dout <= 8'b00000111; // 1799 :   7 - 0x7
      11'h708: dout <= 8'b00000111; // 1800 :   7 - 0x7 -- Background 0xe1
      11'h709: dout <= 8'b00000100; // 1801 :   4 - 0x4
      11'h70A: dout <= 8'b00000000; // 1802 :   0 - 0x0
      11'h70B: dout <= 8'b00000000; // 1803 :   0 - 0x0
      11'h70C: dout <= 8'b00000000; // 1804 :   0 - 0x0
      11'h70D: dout <= 8'b00100000; // 1805 :  32 - 0x20
      11'h70E: dout <= 8'b01110000; // 1806 : 112 - 0x70
      11'h70F: dout <= 8'b11111000; // 1807 : 248 - 0xf8
      11'h710: dout <= 8'b00000000; // 1808 :   0 - 0x0 -- Background 0xe2
      11'h711: dout <= 8'b00000000; // 1809 :   0 - 0x0
      11'h712: dout <= 8'b00000000; // 1810 :   0 - 0x0
      11'h713: dout <= 8'b11111000; // 1811 : 248 - 0xf8
      11'h714: dout <= 8'b11111100; // 1812 : 252 - 0xfc
      11'h715: dout <= 8'b11111100; // 1813 : 252 - 0xfc
      11'h716: dout <= 8'b11111100; // 1814 : 252 - 0xfc
      11'h717: dout <= 8'b11111101; // 1815 : 253 - 0xfd
      11'h718: dout <= 8'b11111100; // 1816 : 252 - 0xfc -- Background 0xe3
      11'h719: dout <= 8'b00011100; // 1817 :  28 - 0x1c
      11'h71A: dout <= 8'b11000000; // 1818 : 192 - 0xc0
      11'h71B: dout <= 8'b11100000; // 1819 : 224 - 0xe0
      11'h71C: dout <= 8'b00000000; // 1820 :   0 - 0x0
      11'h71D: dout <= 8'b00000000; // 1821 :   0 - 0x0
      11'h71E: dout <= 8'b00000110; // 1822 :   6 - 0x6
      11'h71F: dout <= 8'b00001111; // 1823 :  15 - 0xf
      11'h720: dout <= 8'b00000000; // 1824 :   0 - 0x0 -- Background 0xe4
      11'h721: dout <= 8'b00000000; // 1825 :   0 - 0x0
      11'h722: dout <= 8'b00000000; // 1826 :   0 - 0x0
      11'h723: dout <= 8'b00010011; // 1827 :  19 - 0x13
      11'h724: dout <= 8'b00010011; // 1828 :  19 - 0x13
      11'h725: dout <= 8'b00110111; // 1829 :  55 - 0x37
      11'h726: dout <= 8'b00110111; // 1830 :  55 - 0x37
      11'h727: dout <= 8'b00000111; // 1831 :   7 - 0x7
      11'h728: dout <= 8'b00000111; // 1832 :   7 - 0x7 -- Background 0xe5
      11'h729: dout <= 8'b00000100; // 1833 :   4 - 0x4
      11'h72A: dout <= 8'b00000001; // 1834 :   1 - 0x1
      11'h72B: dout <= 8'b00000000; // 1835 :   0 - 0x0
      11'h72C: dout <= 8'b00000000; // 1836 :   0 - 0x0
      11'h72D: dout <= 8'b00100000; // 1837 :  32 - 0x20
      11'h72E: dout <= 8'b01110000; // 1838 : 112 - 0x70
      11'h72F: dout <= 8'b11111000; // 1839 : 248 - 0xf8
      11'h730: dout <= 8'b00000000; // 1840 :   0 - 0x0 -- Background 0xe6
      11'h731: dout <= 8'b00000000; // 1841 :   0 - 0x0
      11'h732: dout <= 8'b00000000; // 1842 :   0 - 0x0
      11'h733: dout <= 8'b11111100; // 1843 : 252 - 0xfc
      11'h734: dout <= 8'b11111100; // 1844 : 252 - 0xfc
      11'h735: dout <= 8'b11111100; // 1845 : 252 - 0xfc
      11'h736: dout <= 8'b11111100; // 1846 : 252 - 0xfc
      11'h737: dout <= 8'b11111101; // 1847 : 253 - 0xfd
      11'h738: dout <= 8'b11111100; // 1848 : 252 - 0xfc -- Background 0xe7
      11'h739: dout <= 8'b00001100; // 1849 :  12 - 0xc
      11'h73A: dout <= 8'b11000000; // 1850 : 192 - 0xc0
      11'h73B: dout <= 8'b11110000; // 1851 : 240 - 0xf0
      11'h73C: dout <= 8'b11110000; // 1852 : 240 - 0xf0
      11'h73D: dout <= 8'b00000000; // 1853 :   0 - 0x0
      11'h73E: dout <= 8'b00000110; // 1854 :   6 - 0x6
      11'h73F: dout <= 8'b00001111; // 1855 :  15 - 0xf
      11'h740: dout <= 8'b11111111; // 1856 : 255 - 0xff -- Background 0xe8
      11'h741: dout <= 8'b11111111; // 1857 : 255 - 0xff
      11'h742: dout <= 8'b01111111; // 1858 : 127 - 0x7f
      11'h743: dout <= 8'b01111111; // 1859 : 127 - 0x7f
      11'h744: dout <= 8'b01111111; // 1860 : 127 - 0x7f
      11'h745: dout <= 8'b00111111; // 1861 :  63 - 0x3f
      11'h746: dout <= 8'b00111111; // 1862 :  63 - 0x3f
      11'h747: dout <= 8'b00111111; // 1863 :  63 - 0x3f
      11'h748: dout <= 8'b00111100; // 1864 :  60 - 0x3c -- Background 0xe9
      11'h749: dout <= 8'b00111110; // 1865 :  62 - 0x3e
      11'h74A: dout <= 8'b00011111; // 1866 :  31 - 0x1f
      11'h74B: dout <= 8'b00001111; // 1867 :  15 - 0xf
      11'h74C: dout <= 8'b00000111; // 1868 :   7 - 0x7
      11'h74D: dout <= 8'b00000000; // 1869 :   0 - 0x0
      11'h74E: dout <= 8'b00000000; // 1870 :   0 - 0x0
      11'h74F: dout <= 8'b00000000; // 1871 :   0 - 0x0
      11'h750: dout <= 8'b11111111; // 1872 : 255 - 0xff -- Background 0xea
      11'h751: dout <= 8'b11111110; // 1873 : 254 - 0xfe
      11'h752: dout <= 8'b11111110; // 1874 : 254 - 0xfe
      11'h753: dout <= 8'b11111100; // 1875 : 252 - 0xfc
      11'h754: dout <= 8'b11111000; // 1876 : 248 - 0xf8
      11'h755: dout <= 8'b11110000; // 1877 : 240 - 0xf0
      11'h756: dout <= 8'b10110000; // 1878 : 176 - 0xb0
      11'h757: dout <= 8'b00111001; // 1879 :  57 - 0x39
      11'h758: dout <= 8'b00011111; // 1880 :  31 - 0x1f -- Background 0xeb
      11'h759: dout <= 8'b11001111; // 1881 : 207 - 0xcf
      11'h75A: dout <= 8'b11000110; // 1882 : 198 - 0xc6
      11'h75B: dout <= 8'b10000000; // 1883 : 128 - 0x80
      11'h75C: dout <= 8'b00000000; // 1884 :   0 - 0x0
      11'h75D: dout <= 8'b00000000; // 1885 :   0 - 0x0
      11'h75E: dout <= 8'b00000000; // 1886 :   0 - 0x0
      11'h75F: dout <= 8'b00000000; // 1887 :   0 - 0x0
      11'h760: dout <= 8'b00000000; // 1888 :   0 - 0x0 -- Background 0xec
      11'h761: dout <= 8'b00000000; // 1889 :   0 - 0x0
      11'h762: dout <= 8'b00000000; // 1890 :   0 - 0x0
      11'h763: dout <= 8'b00000000; // 1891 :   0 - 0x0
      11'h764: dout <= 8'b00000000; // 1892 :   0 - 0x0
      11'h765: dout <= 8'b00000000; // 1893 :   0 - 0x0
      11'h766: dout <= 8'b00001100; // 1894 :  12 - 0xc
      11'h767: dout <= 8'b00001100; // 1895 :  12 - 0xc
      11'h768: dout <= 8'b00110000; // 1896 :  48 - 0x30 -- Background 0xed
      11'h769: dout <= 8'b01000011; // 1897 :  67 - 0x43
      11'h76A: dout <= 8'b01000000; // 1898 :  64 - 0x40
      11'h76B: dout <= 8'b01100000; // 1899 :  96 - 0x60
      11'h76C: dout <= 8'b00000011; // 1900 :   3 - 0x3
      11'h76D: dout <= 8'b00000000; // 1901 :   0 - 0x0
      11'h76E: dout <= 8'b01111111; // 1902 : 127 - 0x7f
      11'h76F: dout <= 8'b00000000; // 1903 :   0 - 0x0
      11'h770: dout <= 8'b00000000; // 1904 :   0 - 0x0 -- Background 0xee
      11'h771: dout <= 8'b00000000; // 1905 :   0 - 0x0
      11'h772: dout <= 8'b00000000; // 1906 :   0 - 0x0
      11'h773: dout <= 8'b00000000; // 1907 :   0 - 0x0
      11'h774: dout <= 8'b00000000; // 1908 :   0 - 0x0
      11'h775: dout <= 8'b00000000; // 1909 :   0 - 0x0
      11'h776: dout <= 8'b00110000; // 1910 :  48 - 0x30
      11'h777: dout <= 8'b00110000; // 1911 :  48 - 0x30
      11'h778: dout <= 8'b00001110; // 1912 :  14 - 0xe -- Background 0xef
      11'h779: dout <= 8'b11001011; // 1913 : 203 - 0xcb
      11'h77A: dout <= 8'b00000000; // 1914 :   0 - 0x0
      11'h77B: dout <= 8'b00000000; // 1915 :   0 - 0x0
      11'h77C: dout <= 8'b11000000; // 1916 : 192 - 0xc0
      11'h77D: dout <= 8'b00000000; // 1917 :   0 - 0x0
      11'h77E: dout <= 8'b11111110; // 1918 : 254 - 0xfe
      11'h77F: dout <= 8'b00000000; // 1919 :   0 - 0x0
      11'h780: dout <= 8'b00000000; // 1920 :   0 - 0x0 -- Background 0xf0
      11'h781: dout <= 8'b00000000; // 1921 :   0 - 0x0
      11'h782: dout <= 8'b00000000; // 1922 :   0 - 0x0
      11'h783: dout <= 8'b00000000; // 1923 :   0 - 0x0
      11'h784: dout <= 8'b00000000; // 1924 :   0 - 0x0
      11'h785: dout <= 8'b00000000; // 1925 :   0 - 0x0
      11'h786: dout <= 8'b00001100; // 1926 :  12 - 0xc
      11'h787: dout <= 8'b00001100; // 1927 :  12 - 0xc
      11'h788: dout <= 8'b00110000; // 1928 :  48 - 0x30 -- Background 0xf1
      11'h789: dout <= 8'b00100011; // 1929 :  35 - 0x23
      11'h78A: dout <= 8'b00100000; // 1930 :  32 - 0x20
      11'h78B: dout <= 8'b01100000; // 1931 :  96 - 0x60
      11'h78C: dout <= 8'b00000011; // 1932 :   3 - 0x3
      11'h78D: dout <= 8'b00000000; // 1933 :   0 - 0x0
      11'h78E: dout <= 8'b01111111; // 1934 : 127 - 0x7f
      11'h78F: dout <= 8'b00000000; // 1935 :   0 - 0x0
      11'h790: dout <= 8'b00000000; // 1936 :   0 - 0x0 -- Background 0xf2
      11'h791: dout <= 8'b00000000; // 1937 :   0 - 0x0
      11'h792: dout <= 8'b00000000; // 1938 :   0 - 0x0
      11'h793: dout <= 8'b00000000; // 1939 :   0 - 0x0
      11'h794: dout <= 8'b00000000; // 1940 :   0 - 0x0
      11'h795: dout <= 8'b00000000; // 1941 :   0 - 0x0
      11'h796: dout <= 8'b00110000; // 1942 :  48 - 0x30
      11'h797: dout <= 8'b00110000; // 1943 :  48 - 0x30
      11'h798: dout <= 8'b00001001; // 1944 :   9 - 0x9 -- Background 0xf3
      11'h799: dout <= 8'b11001111; // 1945 : 207 - 0xcf
      11'h79A: dout <= 8'b00000000; // 1946 :   0 - 0x0
      11'h79B: dout <= 8'b00000000; // 1947 :   0 - 0x0
      11'h79C: dout <= 8'b11000000; // 1948 : 192 - 0xc0
      11'h79D: dout <= 8'b00000000; // 1949 :   0 - 0x0
      11'h79E: dout <= 8'b11111110; // 1950 : 254 - 0xfe
      11'h79F: dout <= 8'b00000000; // 1951 :   0 - 0x0
      11'h7A0: dout <= 8'b00111111; // 1952 :  63 - 0x3f -- Background 0xf4
      11'h7A1: dout <= 8'b00110101; // 1953 :  53 - 0x35
      11'h7A2: dout <= 8'b00011010; // 1954 :  26 - 0x1a
      11'h7A3: dout <= 8'b00001101; // 1955 :  13 - 0xd
      11'h7A4: dout <= 8'b00001010; // 1956 :  10 - 0xa
      11'h7A5: dout <= 8'b00001101; // 1957 :  13 - 0xd
      11'h7A6: dout <= 8'b00001000; // 1958 :   8 - 0x8
      11'h7A7: dout <= 8'b00111000; // 1959 :  56 - 0x38
      11'h7A8: dout <= 8'b01110011; // 1960 : 115 - 0x73 -- Background 0xf5
      11'h7A9: dout <= 8'b11000100; // 1961 : 196 - 0xc4
      11'h7AA: dout <= 8'b11000100; // 1962 : 196 - 0xc4
      11'h7AB: dout <= 8'b11000000; // 1963 : 192 - 0xc0
      11'h7AC: dout <= 8'b11000001; // 1964 : 193 - 0xc1
      11'h7AD: dout <= 8'b11000000; // 1965 : 192 - 0xc0
      11'h7AE: dout <= 8'b01100001; // 1966 :  97 - 0x61
      11'h7AF: dout <= 8'b00111111; // 1967 :  63 - 0x3f
      11'h7B0: dout <= 8'b11111100; // 1968 : 252 - 0xfc -- Background 0xf6
      11'h7B1: dout <= 8'b01010100; // 1969 :  84 - 0x54
      11'h7B2: dout <= 8'b10101000; // 1970 : 168 - 0xa8
      11'h7B3: dout <= 8'b01010000; // 1971 :  80 - 0x50
      11'h7B4: dout <= 8'b10110000; // 1972 : 176 - 0xb0
      11'h7B5: dout <= 8'b01010000; // 1973 :  80 - 0x50
      11'h7B6: dout <= 8'b10010000; // 1974 : 144 - 0x90
      11'h7B7: dout <= 8'b00011100; // 1975 :  28 - 0x1c
      11'h7B8: dout <= 8'b10000110; // 1976 : 134 - 0x86 -- Background 0xf7
      11'h7B9: dout <= 8'b01000010; // 1977 :  66 - 0x42
      11'h7BA: dout <= 8'b01000111; // 1978 :  71 - 0x47
      11'h7BB: dout <= 8'b01000001; // 1979 :  65 - 0x41
      11'h7BC: dout <= 8'b10000011; // 1980 : 131 - 0x83
      11'h7BD: dout <= 8'b00000001; // 1981 :   1 - 0x1
      11'h7BE: dout <= 8'b10000110; // 1982 : 134 - 0x86
      11'h7BF: dout <= 8'b11111100; // 1983 : 252 - 0xfc
      11'h7C0: dout <= 8'b11100100; // 1984 : 228 - 0xe4 -- Background 0xf8
      11'h7C1: dout <= 8'b11100100; // 1985 : 228 - 0xe4
      11'h7C2: dout <= 8'b11101111; // 1986 : 239 - 0xef
      11'h7C3: dout <= 8'b11101111; // 1987 : 239 - 0xef
      11'h7C4: dout <= 8'b11111111; // 1988 : 255 - 0xff
      11'h7C5: dout <= 8'b11111111; // 1989 : 255 - 0xff
      11'h7C6: dout <= 8'b01111111; // 1990 : 127 - 0x7f
      11'h7C7: dout <= 8'b01111111; // 1991 : 127 - 0x7f
      11'h7C8: dout <= 8'b00111111; // 1992 :  63 - 0x3f -- Background 0xf9
      11'h7C9: dout <= 8'b01111111; // 1993 : 127 - 0x7f
      11'h7CA: dout <= 8'b01111111; // 1994 : 127 - 0x7f
      11'h7CB: dout <= 8'b11111111; // 1995 : 255 - 0xff
      11'h7CC: dout <= 8'b11111111; // 1996 : 255 - 0xff
      11'h7CD: dout <= 8'b11111111; // 1997 : 255 - 0xff
      11'h7CE: dout <= 8'b11111111; // 1998 : 255 - 0xff
      11'h7CF: dout <= 8'b11111111; // 1999 : 255 - 0xff
      11'h7D0: dout <= 8'b00010011; // 2000 :  19 - 0x13 -- Background 0xfa
      11'h7D1: dout <= 8'b00010011; // 2001 :  19 - 0x13
      11'h7D2: dout <= 8'b11111011; // 2002 : 251 - 0xfb
      11'h7D3: dout <= 8'b11111011; // 2003 : 251 - 0xfb
      11'h7D4: dout <= 8'b11111111; // 2004 : 255 - 0xff
      11'h7D5: dout <= 8'b11111111; // 2005 : 255 - 0xff
      11'h7D6: dout <= 8'b11111110; // 2006 : 254 - 0xfe
      11'h7D7: dout <= 8'b11111110; // 2007 : 254 - 0xfe
      11'h7D8: dout <= 8'b11111110; // 2008 : 254 - 0xfe -- Background 0xfb
      11'h7D9: dout <= 8'b11111111; // 2009 : 255 - 0xff
      11'h7DA: dout <= 8'b11111111; // 2010 : 255 - 0xff
      11'h7DB: dout <= 8'b11111111; // 2011 : 255 - 0xff
      11'h7DC: dout <= 8'b11111111; // 2012 : 255 - 0xff
      11'h7DD: dout <= 8'b11111111; // 2013 : 255 - 0xff
      11'h7DE: dout <= 8'b11111111; // 2014 : 255 - 0xff
      11'h7DF: dout <= 8'b11111111; // 2015 : 255 - 0xff
      11'h7E0: dout <= 8'b00000000; // 2016 :   0 - 0x0 -- Background 0xfc
      11'h7E1: dout <= 8'b00000000; // 2017 :   0 - 0x0
      11'h7E2: dout <= 8'b01111100; // 2018 : 124 - 0x7c
      11'h7E3: dout <= 8'b11111110; // 2019 : 254 - 0xfe
      11'h7E4: dout <= 8'b11111110; // 2020 : 254 - 0xfe
      11'h7E5: dout <= 8'b01111100; // 2021 : 124 - 0x7c
      11'h7E6: dout <= 8'b01000100; // 2022 :  68 - 0x44
      11'h7E7: dout <= 8'b10000010; // 2023 : 130 - 0x82
      11'h7E8: dout <= 8'b10000010; // 2024 : 130 - 0x82 -- Background 0xfd
      11'h7E9: dout <= 8'b10000010; // 2025 : 130 - 0x82
      11'h7EA: dout <= 8'b10000010; // 2026 : 130 - 0x82
      11'h7EB: dout <= 8'b11000110; // 2027 : 198 - 0xc6
      11'h7EC: dout <= 8'b11111110; // 2028 : 254 - 0xfe
      11'h7ED: dout <= 8'b11111110; // 2029 : 254 - 0xfe
      11'h7EE: dout <= 8'b10111010; // 2030 : 186 - 0xba
      11'h7EF: dout <= 8'b01111100; // 2031 : 124 - 0x7c
      11'h7F0: dout <= 8'b00000000; // 2032 :   0 - 0x0 -- Background 0xfe
      11'h7F1: dout <= 8'b00011001; // 2033 :  25 - 0x19
      11'h7F2: dout <= 8'b00111110; // 2034 :  62 - 0x3e
      11'h7F3: dout <= 8'b00111100; // 2035 :  60 - 0x3c
      11'h7F4: dout <= 8'b00111100; // 2036 :  60 - 0x3c
      11'h7F5: dout <= 8'b00111100; // 2037 :  60 - 0x3c
      11'h7F6: dout <= 8'b00111110; // 2038 :  62 - 0x3e
      11'h7F7: dout <= 8'b00011001; // 2039 :  25 - 0x19
      11'h7F8: dout <= 8'b00000000; // 2040 :   0 - 0x0 -- Background 0xff
      11'h7F9: dout <= 8'b11111110; // 2041 : 254 - 0xfe
      11'h7FA: dout <= 8'b00011101; // 2042 :  29 - 0x1d
      11'h7FB: dout <= 8'b00001111; // 2043 :  15 - 0xf
      11'h7FC: dout <= 8'b00001111; // 2044 :  15 - 0xf
      11'h7FD: dout <= 8'b00001111; // 2045 :  15 - 0xf
      11'h7FE: dout <= 8'b00011101; // 2046 :  29 - 0x1d
      11'h7FF: dout <= 8'b11111110; // 2047 : 254 - 0xfe
    endcase
  end

endmodule
