--- Autcmatically generated VHDL ROM from a NES memory file----
---   NAME TABLE
-- https://wiki.nesdev.com/w/index.php/PPU_nametables
--- Only the first Name Table: 1KiB


---  Original memory dump file name: sprilo_ntable_00.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_NTABLE0_SPRILO_00 is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(10-1 downto 0);  --1024 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_NTABLE0_SPRILO_00;

architecture BEHAVIORAL of ROM_NTABLE0_SPRILO_00 is
  signal addr_int  : natural range 0 to 2**10-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
     ------- Name Table 0---------
    "11111010", --    0 -  0x0  :  250 - 0xfa -- line 0x0
    "11111010", --    1 -  0x1  :  250 - 0xfa
    "11111010", --    2 -  0x2  :  250 - 0xfa
    "11101010", --    3 -  0x3  :  234 - 0xea
    "11111010", --    4 -  0x4  :  250 - 0xfa
    "11111010", --    5 -  0x5  :  250 - 0xfa
    "11111010", --    6 -  0x6  :  250 - 0xfa
    "11111010", --    7 -  0x7  :  250 - 0xfa
    "11111010", --    8 -  0x8  :  250 - 0xfa
    "11111010", --    9 -  0x9  :  250 - 0xfa
    "11111010", --   10 -  0xa  :  250 - 0xfa
    "11111010", --   11 -  0xb  :  250 - 0xfa
    "11111010", --   12 -  0xc  :  250 - 0xfa
    "11111010", --   13 -  0xd  :  250 - 0xfa
    "11101010", --   14 -  0xe  :  234 - 0xea
    "11111010", --   15 -  0xf  :  250 - 0xfa
    "11111010", --   16 - 0x10  :  250 - 0xfa
    "11111010", --   17 - 0x11  :  250 - 0xfa
    "11111010", --   18 - 0x12  :  250 - 0xfa
    "11111010", --   19 - 0x13  :  250 - 0xfa
    "11111010", --   20 - 0x14  :  250 - 0xfa
    "11111010", --   21 - 0x15  :  250 - 0xfa
    "11111010", --   22 - 0x16  :  250 - 0xfa
    "11111010", --   23 - 0x17  :  250 - 0xfa
    "11111010", --   24 - 0x18  :  250 - 0xfa
    "11111010", --   25 - 0x19  :  250 - 0xfa
    "11111010", --   26 - 0x1a  :  250 - 0xfa
    "11111010", --   27 - 0x1b  :  250 - 0xfa
    "11111010", --   28 - 0x1c  :  250 - 0xfa
    "11111010", --   29 - 0x1d  :  250 - 0xfa
    "11111010", --   30 - 0x1e  :  250 - 0xfa
    "11111010", --   31 - 0x1f  :  250 - 0xfa
    "11111010", --   32 - 0x20  :  250 - 0xfa -- line 0x1
    "11100111", --   33 - 0x21  :  231 - 0xe7
    "11111011", --   34 - 0x22  :  251 - 0xfb
    "11111011", --   35 - 0x23  :  251 - 0xfb
    "11111011", --   36 - 0x24  :  251 - 0xfb
    "11111011", --   37 - 0x25  :  251 - 0xfb
    "11111011", --   38 - 0x26  :  251 - 0xfb
    "11111011", --   39 - 0x27  :  251 - 0xfb
    "11111011", --   40 - 0x28  :  251 - 0xfb
    "11111011", --   41 - 0x29  :  251 - 0xfb
    "11111011", --   42 - 0x2a  :  251 - 0xfb
    "11111011", --   43 - 0x2b  :  251 - 0xfb
    "11111011", --   44 - 0x2c  :  251 - 0xfb
    "11111011", --   45 - 0x2d  :  251 - 0xfb
    "11111011", --   46 - 0x2e  :  251 - 0xfb
    "11111011", --   47 - 0x2f  :  251 - 0xfb
    "11111011", --   48 - 0x30  :  251 - 0xfb
    "11111011", --   49 - 0x31  :  251 - 0xfb
    "11111011", --   50 - 0x32  :  251 - 0xfb
    "11111011", --   51 - 0x33  :  251 - 0xfb
    "11111011", --   52 - 0x34  :  251 - 0xfb
    "11111011", --   53 - 0x35  :  251 - 0xfb
    "11101000", --   54 - 0x36  :  232 - 0xe8
    "11111010", --   55 - 0x37  :  250 - 0xfa
    "11111010", --   56 - 0x38  :  250 - 0xfa
    "11101001", --   57 - 0x39  :  233 - 0xe9
    "11111001", --   58 - 0x3a  :  249 - 0xf9
    "11101001", --   59 - 0x3b  :  233 - 0xe9
    "11111010", --   60 - 0x3c  :  250 - 0xfa
    "11111010", --   61 - 0x3d  :  250 - 0xfa
    "11101001", --   62 - 0x3e  :  233 - 0xe9
    "11111010", --   63 - 0x3f  :  250 - 0xfa
    "11101010", --   64 - 0x40  :  234 - 0xea -- line 0x2
    "11111100", --   65 - 0x41  :  252 - 0xfc
    "11111111", --   66 - 0x42  :  255 - 0xff
    "11111111", --   67 - 0x43  :  255 - 0xff
    "11111111", --   68 - 0x44  :  255 - 0xff
    "11111111", --   69 - 0x45  :  255 - 0xff
    "11111111", --   70 - 0x46  :  255 - 0xff
    "11111111", --   71 - 0x47  :  255 - 0xff
    "11111111", --   72 - 0x48  :  255 - 0xff
    "11111111", --   73 - 0x49  :  255 - 0xff
    "11111111", --   74 - 0x4a  :  255 - 0xff
    "11111111", --   75 - 0x4b  :  255 - 0xff
    "11111111", --   76 - 0x4c  :  255 - 0xff
    "11111111", --   77 - 0x4d  :  255 - 0xff
    "11111111", --   78 - 0x4e  :  255 - 0xff
    "11111111", --   79 - 0x4f  :  255 - 0xff
    "11111111", --   80 - 0x50  :  255 - 0xff
    "11111111", --   81 - 0x51  :  255 - 0xff
    "11111111", --   82 - 0x52  :  255 - 0xff
    "11111111", --   83 - 0x53  :  255 - 0xff
    "11111111", --   84 - 0x54  :  255 - 0xff
    "11111111", --   85 - 0x55  :  255 - 0xff
    "11101100", --   86 - 0x56  :  236 - 0xec
    "11111010", --   87 - 0x57  :  250 - 0xfa
    "11111010", --   88 - 0x58  :  250 - 0xfa
    "11111010", --   89 - 0x59  :  250 - 0xfa
    "11111010", --   90 - 0x5a  :  250 - 0xfa
    "11111010", --   91 - 0x5b  :  250 - 0xfa
    "11111010", --   92 - 0x5c  :  250 - 0xfa
    "11101001", --   93 - 0x5d  :  233 - 0xe9
    "11111010", --   94 - 0x5e  :  250 - 0xfa
    "11111010", --   95 - 0x5f  :  250 - 0xfa
    "11111010", --   96 - 0x60  :  250 - 0xfa -- line 0x3
    "11111100", --   97 - 0x61  :  252 - 0xfc
    "11111111", --   98 - 0x62  :  255 - 0xff
    "11111111", --   99 - 0x63  :  255 - 0xff
    "11111111", --  100 - 0x64  :  255 - 0xff
    "11111111", --  101 - 0x65  :  255 - 0xff
    "11111101", --  102 - 0x66  :  253 - 0xfd
    "11111111", --  103 - 0x67  :  255 - 0xff
    "11111101", --  104 - 0x68  :  253 - 0xfd
    "11111111", --  105 - 0x69  :  255 - 0xff
    "11111101", --  106 - 0x6a  :  253 - 0xfd
    "11111111", --  107 - 0x6b  :  255 - 0xff
    "11111101", --  108 - 0x6c  :  253 - 0xfd
    "11111111", --  109 - 0x6d  :  255 - 0xff
    "11111101", --  110 - 0x6e  :  253 - 0xfd
    "11111111", --  111 - 0x6f  :  255 - 0xff
    "11111101", --  112 - 0x70  :  253 - 0xfd
    "11111111", --  113 - 0x71  :  255 - 0xff
    "11111101", --  114 - 0x72  :  253 - 0xfd
    "11111111", --  115 - 0x73  :  255 - 0xff
    "11111111", --  116 - 0x74  :  255 - 0xff
    "11111111", --  117 - 0x75  :  255 - 0xff
    "11101100", --  118 - 0x76  :  236 - 0xec
    "11111010", --  119 - 0x77  :  250 - 0xfa
    "11111010", --  120 - 0x78  :  250 - 0xfa
    "11111010", --  121 - 0x79  :  250 - 0xfa
    "11111010", --  122 - 0x7a  :  250 - 0xfa
    "11111010", --  123 - 0x7b  :  250 - 0xfa
    "11111010", --  124 - 0x7c  :  250 - 0xfa
    "11111010", --  125 - 0x7d  :  250 - 0xfa
    "11111010", --  126 - 0x7e  :  250 - 0xfa
    "11111010", --  127 - 0x7f  :  250 - 0xfa
    "11101001", --  128 - 0x80  :  233 - 0xe9 -- line 0x4
    "11111100", --  129 - 0x81  :  252 - 0xfc
    "11111111", --  130 - 0x82  :  255 - 0xff
    "11111111", --  131 - 0x83  :  255 - 0xff
    "11111111", --  132 - 0x84  :  255 - 0xff
    "11111111", --  133 - 0x85  :  255 - 0xff
    "11111101", --  134 - 0x86  :  253 - 0xfd
    "11111111", --  135 - 0x87  :  255 - 0xff
    "11111101", --  136 - 0x88  :  253 - 0xfd
    "11111111", --  137 - 0x89  :  255 - 0xff
    "11111101", --  138 - 0x8a  :  253 - 0xfd
    "11111111", --  139 - 0x8b  :  255 - 0xff
    "11111101", --  140 - 0x8c  :  253 - 0xfd
    "11111111", --  141 - 0x8d  :  255 - 0xff
    "11111101", --  142 - 0x8e  :  253 - 0xfd
    "11111111", --  143 - 0x8f  :  255 - 0xff
    "11111101", --  144 - 0x90  :  253 - 0xfd
    "11111111", --  145 - 0x91  :  255 - 0xff
    "11111101", --  146 - 0x92  :  253 - 0xfd
    "11111111", --  147 - 0x93  :  255 - 0xff
    "11111111", --  148 - 0x94  :  255 - 0xff
    "11111111", --  149 - 0x95  :  255 - 0xff
    "11101100", --  150 - 0x96  :  236 - 0xec
    "11101001", --  151 - 0x97  :  233 - 0xe9
    "11111010", --  152 - 0x98  :  250 - 0xfa
    "11111010", --  153 - 0x99  :  250 - 0xfa
    "11101010", --  154 - 0x9a  :  234 - 0xea
    "11111010", --  155 - 0x9b  :  250 - 0xfa
    "11111001", --  156 - 0x9c  :  249 - 0xf9
    "11111010", --  157 - 0x9d  :  250 - 0xfa
    "11111010", --  158 - 0x9e  :  250 - 0xfa
    "11111010", --  159 - 0x9f  :  250 - 0xfa
    "11111010", --  160 - 0xa0  :  250 - 0xfa -- line 0x5
    "11111100", --  161 - 0xa1  :  252 - 0xfc
    "11111111", --  162 - 0xa2  :  255 - 0xff
    "11111111", --  163 - 0xa3  :  255 - 0xff
    "11111111", --  164 - 0xa4  :  255 - 0xff
    "11111111", --  165 - 0xa5  :  255 - 0xff
    "11111111", --  166 - 0xa6  :  255 - 0xff
    "11111111", --  167 - 0xa7  :  255 - 0xff
    "11111111", --  168 - 0xa8  :  255 - 0xff
    "11111111", --  169 - 0xa9  :  255 - 0xff
    "11111111", --  170 - 0xaa  :  255 - 0xff
    "11111111", --  171 - 0xab  :  255 - 0xff
    "11111111", --  172 - 0xac  :  255 - 0xff
    "11111111", --  173 - 0xad  :  255 - 0xff
    "11111111", --  174 - 0xae  :  255 - 0xff
    "11111111", --  175 - 0xaf  :  255 - 0xff
    "11111111", --  176 - 0xb0  :  255 - 0xff
    "11111111", --  177 - 0xb1  :  255 - 0xff
    "11111111", --  178 - 0xb2  :  255 - 0xff
    "11111111", --  179 - 0xb3  :  255 - 0xff
    "11111111", --  180 - 0xb4  :  255 - 0xff
    "11111111", --  181 - 0xb5  :  255 - 0xff
    "11110101", --  182 - 0xb6  :  245 - 0xf5
    "11111011", --  183 - 0xb7  :  251 - 0xfb
    "11111011", --  184 - 0xb8  :  251 - 0xfb
    "11111011", --  185 - 0xb9  :  251 - 0xfb
    "11111011", --  186 - 0xba  :  251 - 0xfb
    "11111011", --  187 - 0xbb  :  251 - 0xfb
    "11111011", --  188 - 0xbc  :  251 - 0xfb
    "11111011", --  189 - 0xbd  :  251 - 0xfb
    "11101000", --  190 - 0xbe  :  232 - 0xe8
    "11111010", --  191 - 0xbf  :  250 - 0xfa
    "11111010", --  192 - 0xc0  :  250 - 0xfa -- line 0x6
    "11111100", --  193 - 0xc1  :  252 - 0xfc
    "11111111", --  194 - 0xc2  :  255 - 0xff
    "11111111", --  195 - 0xc3  :  255 - 0xff
    "11111111", --  196 - 0xc4  :  255 - 0xff
    "11111111", --  197 - 0xc5  :  255 - 0xff
    "11100101", --  198 - 0xc6  :  229 - 0xe5
    "11101011", --  199 - 0xc7  :  235 - 0xeb
    "11101011", --  200 - 0xc8  :  235 - 0xeb
    "11101011", --  201 - 0xc9  :  235 - 0xeb
    "11101011", --  202 - 0xca  :  235 - 0xeb
    "11101011", --  203 - 0xcb  :  235 - 0xeb
    "11101011", --  204 - 0xcc  :  235 - 0xeb
    "11101011", --  205 - 0xcd  :  235 - 0xeb
    "11101011", --  206 - 0xce  :  235 - 0xeb
    "11101011", --  207 - 0xcf  :  235 - 0xeb
    "11101011", --  208 - 0xd0  :  235 - 0xeb
    "11100110", --  209 - 0xd1  :  230 - 0xe6
    "11111111", --  210 - 0xd2  :  255 - 0xff
    "11111110", --  211 - 0xd3  :  254 - 0xfe
    "11111110", --  212 - 0xd4  :  254 - 0xfe
    "11111111", --  213 - 0xd5  :  255 - 0xff
    "11111111", --  214 - 0xd6  :  255 - 0xff
    "11111111", --  215 - 0xd7  :  255 - 0xff
    "11111111", --  216 - 0xd8  :  255 - 0xff
    "11111111", --  217 - 0xd9  :  255 - 0xff
    "11111111", --  218 - 0xda  :  255 - 0xff
    "11111111", --  219 - 0xdb  :  255 - 0xff
    "11111111", --  220 - 0xdc  :  255 - 0xff
    "11111111", --  221 - 0xdd  :  255 - 0xff
    "11101100", --  222 - 0xde  :  236 - 0xec
    "11111010", --  223 - 0xdf  :  250 - 0xfa
    "11111010", --  224 - 0xe0  :  250 - 0xfa -- line 0x7
    "11111100", --  225 - 0xe1  :  252 - 0xfc
    "11111111", --  226 - 0xe2  :  255 - 0xff
    "11111110", --  227 - 0xe3  :  254 - 0xfe
    "11111110", --  228 - 0xe4  :  254 - 0xfe
    "11111111", --  229 - 0xe5  :  255 - 0xff
    "11101100", --  230 - 0xe6  :  236 - 0xec
    "11111010", --  231 - 0xe7  :  250 - 0xfa
    "11111010", --  232 - 0xe8  :  250 - 0xfa
    "11111001", --  233 - 0xe9  :  249 - 0xf9
    "11111010", --  234 - 0xea  :  250 - 0xfa
    "11111010", --  235 - 0xeb  :  250 - 0xfa
    "11111010", --  236 - 0xec  :  250 - 0xfa
    "11111010", --  237 - 0xed  :  250 - 0xfa
    "11111010", --  238 - 0xee  :  250 - 0xfa
    "11111010", --  239 - 0xef  :  250 - 0xfa
    "11111010", --  240 - 0xf0  :  250 - 0xfa
    "11111100", --  241 - 0xf1  :  252 - 0xfc
    "11111111", --  242 - 0xf2  :  255 - 0xff
    "11111111", --  243 - 0xf3  :  255 - 0xff
    "11111111", --  244 - 0xf4  :  255 - 0xff
    "11111111", --  245 - 0xf5  :  255 - 0xff
    "11111101", --  246 - 0xf6  :  253 - 0xfd
    "11111111", --  247 - 0xf7  :  255 - 0xff
    "11111101", --  248 - 0xf8  :  253 - 0xfd
    "11111111", --  249 - 0xf9  :  255 - 0xff
    "11111101", --  250 - 0xfa  :  253 - 0xfd
    "11111111", --  251 - 0xfb  :  255 - 0xff
    "11111111", --  252 - 0xfc  :  255 - 0xff
    "11111111", --  253 - 0xfd  :  255 - 0xff
    "11101100", --  254 - 0xfe  :  236 - 0xec
    "11111010", --  255 - 0xff  :  250 - 0xfa
    "11111010", --  256 - 0x100  :  250 - 0xfa -- line 0x8
    "11111100", --  257 - 0x101  :  252 - 0xfc
    "11111111", --  258 - 0x102  :  255 - 0xff
    "11111111", --  259 - 0x103  :  255 - 0xff
    "11111111", --  260 - 0x104  :  255 - 0xff
    "11111111", --  261 - 0x105  :  255 - 0xff
    "11101100", --  262 - 0x106  :  236 - 0xec
    "11111010", --  263 - 0x107  :  250 - 0xfa
    "11111010", --  264 - 0x108  :  250 - 0xfa
    "11111010", --  265 - 0x109  :  250 - 0xfa
    "11111010", --  266 - 0x10a  :  250 - 0xfa
    "11111010", --  267 - 0x10b  :  250 - 0xfa
    "11111010", --  268 - 0x10c  :  250 - 0xfa
    "11111010", --  269 - 0x10d  :  250 - 0xfa
    "11111010", --  270 - 0x10e  :  250 - 0xfa
    "11111010", --  271 - 0x10f  :  250 - 0xfa
    "11111010", --  272 - 0x110  :  250 - 0xfa
    "11111100", --  273 - 0x111  :  252 - 0xfc
    "11111111", --  274 - 0x112  :  255 - 0xff
    "11111111", --  275 - 0x113  :  255 - 0xff
    "11111111", --  276 - 0x114  :  255 - 0xff
    "11111111", --  277 - 0x115  :  255 - 0xff
    "11111101", --  278 - 0x116  :  253 - 0xfd
    "11111111", --  279 - 0x117  :  255 - 0xff
    "11111101", --  280 - 0x118  :  253 - 0xfd
    "11111111", --  281 - 0x119  :  255 - 0xff
    "11111101", --  282 - 0x11a  :  253 - 0xfd
    "11111111", --  283 - 0x11b  :  255 - 0xff
    "11111111", --  284 - 0x11c  :  255 - 0xff
    "11111111", --  285 - 0x11d  :  255 - 0xff
    "11101100", --  286 - 0x11e  :  236 - 0xec
    "11111010", --  287 - 0x11f  :  250 - 0xfa
    "11111010", --  288 - 0x120  :  250 - 0xfa -- line 0x9
    "11111100", --  289 - 0x121  :  252 - 0xfc
    "11111111", --  290 - 0x122  :  255 - 0xff
    "11111110", --  291 - 0x123  :  254 - 0xfe
    "11111110", --  292 - 0x124  :  254 - 0xfe
    "11111111", --  293 - 0x125  :  255 - 0xff
    "11101100", --  294 - 0x126  :  236 - 0xec
    "11111010", --  295 - 0x127  :  250 - 0xfa
    "11111010", --  296 - 0x128  :  250 - 0xfa
    "11101001", --  297 - 0x129  :  233 - 0xe9
    "11111010", --  298 - 0x12a  :  250 - 0xfa
    "11101001", --  299 - 0x12b  :  233 - 0xe9
    "11111010", --  300 - 0x12c  :  250 - 0xfa
    "11111010", --  301 - 0x12d  :  250 - 0xfa
    "11101001", --  302 - 0x12e  :  233 - 0xe9
    "11111010", --  303 - 0x12f  :  250 - 0xfa
    "11111010", --  304 - 0x130  :  250 - 0xfa
    "11111100", --  305 - 0x131  :  252 - 0xfc
    "11111111", --  306 - 0x132  :  255 - 0xff
    "11111111", --  307 - 0x133  :  255 - 0xff
    "11111111", --  308 - 0x134  :  255 - 0xff
    "11111111", --  309 - 0x135  :  255 - 0xff
    "11111111", --  310 - 0x136  :  255 - 0xff
    "11111111", --  311 - 0x137  :  255 - 0xff
    "11111111", --  312 - 0x138  :  255 - 0xff
    "11111111", --  313 - 0x139  :  255 - 0xff
    "11111111", --  314 - 0x13a  :  255 - 0xff
    "11111111", --  315 - 0x13b  :  255 - 0xff
    "11111111", --  316 - 0x13c  :  255 - 0xff
    "11111111", --  317 - 0x13d  :  255 - 0xff
    "11101100", --  318 - 0x13e  :  236 - 0xec
    "11111010", --  319 - 0x13f  :  250 - 0xfa
    "11111010", --  320 - 0x140  :  250 - 0xfa -- line 0xa
    "11111100", --  321 - 0x141  :  252 - 0xfc
    "11111111", --  322 - 0x142  :  255 - 0xff
    "11111111", --  323 - 0x143  :  255 - 0xff
    "11111111", --  324 - 0x144  :  255 - 0xff
    "11111111", --  325 - 0x145  :  255 - 0xff
    "11101100", --  326 - 0x146  :  236 - 0xec
    "11111010", --  327 - 0x147  :  250 - 0xfa
    "11111010", --  328 - 0x148  :  250 - 0xfa
    "11111010", --  329 - 0x149  :  250 - 0xfa
    "11111010", --  330 - 0x14a  :  250 - 0xfa
    "11101001", --  331 - 0x14b  :  233 - 0xe9
    "11111010", --  332 - 0x14c  :  250 - 0xfa
    "11111010", --  333 - 0x14d  :  250 - 0xfa
    "11111010", --  334 - 0x14e  :  250 - 0xfa
    "11111010", --  335 - 0x14f  :  250 - 0xfa
    "11111010", --  336 - 0x150  :  250 - 0xfa
    "11110111", --  337 - 0x151  :  247 - 0xf7
    "11101011", --  338 - 0x152  :  235 - 0xeb
    "11101011", --  339 - 0x153  :  235 - 0xeb
    "11101011", --  340 - 0x154  :  235 - 0xeb
    "11101011", --  341 - 0x155  :  235 - 0xeb
    "11101011", --  342 - 0x156  :  235 - 0xeb
    "11101011", --  343 - 0x157  :  235 - 0xeb
    "11101011", --  344 - 0x158  :  235 - 0xeb
    "11100110", --  345 - 0x159  :  230 - 0xe6
    "11111111", --  346 - 0x15a  :  255 - 0xff
    "11111111", --  347 - 0x15b  :  255 - 0xff
    "11111111", --  348 - 0x15c  :  255 - 0xff
    "11111111", --  349 - 0x15d  :  255 - 0xff
    "11101100", --  350 - 0x15e  :  236 - 0xec
    "11111010", --  351 - 0x15f  :  250 - 0xfa
    "11111010", --  352 - 0x160  :  250 - 0xfa -- line 0xb
    "11111100", --  353 - 0x161  :  252 - 0xfc
    "11111111", --  354 - 0x162  :  255 - 0xff
    "11111110", --  355 - 0x163  :  254 - 0xfe
    "11111110", --  356 - 0x164  :  254 - 0xfe
    "11111111", --  357 - 0x165  :  255 - 0xff
    "11101100", --  358 - 0x166  :  236 - 0xec
    "11111010", --  359 - 0x167  :  250 - 0xfa
    "11111010", --  360 - 0x168  :  250 - 0xfa
    "11111010", --  361 - 0x169  :  250 - 0xfa
    "11111010", --  362 - 0x16a  :  250 - 0xfa
    "11111010", --  363 - 0x16b  :  250 - 0xfa
    "11111010", --  364 - 0x16c  :  250 - 0xfa
    "11111010", --  365 - 0x16d  :  250 - 0xfa
    "11111010", --  366 - 0x16e  :  250 - 0xfa
    "11111010", --  367 - 0x16f  :  250 - 0xfa
    "11111010", --  368 - 0x170  :  250 - 0xfa
    "11111010", --  369 - 0x171  :  250 - 0xfa
    "11111010", --  370 - 0x172  :  250 - 0xfa
    "11111010", --  371 - 0x173  :  250 - 0xfa
    "11111010", --  372 - 0x174  :  250 - 0xfa
    "11111010", --  373 - 0x175  :  250 - 0xfa
    "11111010", --  374 - 0x176  :  250 - 0xfa
    "11101001", --  375 - 0x177  :  233 - 0xe9
    "11111010", --  376 - 0x178  :  250 - 0xfa
    "11111100", --  377 - 0x179  :  252 - 0xfc
    "11111111", --  378 - 0x17a  :  255 - 0xff
    "11111110", --  379 - 0x17b  :  254 - 0xfe
    "11111110", --  380 - 0x17c  :  254 - 0xfe
    "11111111", --  381 - 0x17d  :  255 - 0xff
    "11101100", --  382 - 0x17e  :  236 - 0xec
    "11111010", --  383 - 0x17f  :  250 - 0xfa
    "11101001", --  384 - 0x180  :  233 - 0xe9 -- line 0xc
    "11111100", --  385 - 0x181  :  252 - 0xfc
    "11111111", --  386 - 0x182  :  255 - 0xff
    "11111111", --  387 - 0x183  :  255 - 0xff
    "11111111", --  388 - 0x184  :  255 - 0xff
    "11111111", --  389 - 0x185  :  255 - 0xff
    "11101100", --  390 - 0x186  :  236 - 0xec
    "11111010", --  391 - 0x187  :  250 - 0xfa
    "11111010", --  392 - 0x188  :  250 - 0xfa
    "11111010", --  393 - 0x189  :  250 - 0xfa
    "11111010", --  394 - 0x18a  :  250 - 0xfa
    "11111010", --  395 - 0x18b  :  250 - 0xfa
    "11111010", --  396 - 0x18c  :  250 - 0xfa
    "11111010", --  397 - 0x18d  :  250 - 0xfa
    "11111010", --  398 - 0x18e  :  250 - 0xfa
    "11101001", --  399 - 0x18f  :  233 - 0xe9
    "11111010", --  400 - 0x190  :  250 - 0xfa
    "11101001", --  401 - 0x191  :  233 - 0xe9
    "11111010", --  402 - 0x192  :  250 - 0xfa
    "11111010", --  403 - 0x193  :  250 - 0xfa
    "11111010", --  404 - 0x194  :  250 - 0xfa
    "11111010", --  405 - 0x195  :  250 - 0xfa
    "11111010", --  406 - 0x196  :  250 - 0xfa
    "11111010", --  407 - 0x197  :  250 - 0xfa
    "11111010", --  408 - 0x198  :  250 - 0xfa
    "11111100", --  409 - 0x199  :  252 - 0xfc
    "11111111", --  410 - 0x19a  :  255 - 0xff
    "11111111", --  411 - 0x19b  :  255 - 0xff
    "11111111", --  412 - 0x19c  :  255 - 0xff
    "11111111", --  413 - 0x19d  :  255 - 0xff
    "11101100", --  414 - 0x19e  :  236 - 0xec
    "11111010", --  415 - 0x19f  :  250 - 0xfa
    "11111010", --  416 - 0x1a0  :  250 - 0xfa -- line 0xd
    "11111100", --  417 - 0x1a1  :  252 - 0xfc
    "11111111", --  418 - 0x1a2  :  255 - 0xff
    "11111110", --  419 - 0x1a3  :  254 - 0xfe
    "11111110", --  420 - 0x1a4  :  254 - 0xfe
    "11111111", --  421 - 0x1a5  :  255 - 0xff
    "11101100", --  422 - 0x1a6  :  236 - 0xec
    "11111010", --  423 - 0x1a7  :  250 - 0xfa
    "11111001", --  424 - 0x1a8  :  249 - 0xf9
    "11111010", --  425 - 0x1a9  :  250 - 0xfa
    "11111010", --  426 - 0x1aa  :  250 - 0xfa
    "11101001", --  427 - 0x1ab  :  233 - 0xe9
    "11111010", --  428 - 0x1ac  :  250 - 0xfa
    "11111010", --  429 - 0x1ad  :  250 - 0xfa
    "11111010", --  430 - 0x1ae  :  250 - 0xfa
    "11111010", --  431 - 0x1af  :  250 - 0xfa
    "11111010", --  432 - 0x1b0  :  250 - 0xfa
    "11111010", --  433 - 0x1b1  :  250 - 0xfa
    "11111010", --  434 - 0x1b2  :  250 - 0xfa
    "11100111", --  435 - 0x1b3  :  231 - 0xe7
    "11111011", --  436 - 0x1b4  :  251 - 0xfb
    "11111011", --  437 - 0x1b5  :  251 - 0xfb
    "11111011", --  438 - 0x1b6  :  251 - 0xfb
    "11111011", --  439 - 0x1b7  :  251 - 0xfb
    "11111011", --  440 - 0x1b8  :  251 - 0xfb
    "11110110", --  441 - 0x1b9  :  246 - 0xf6
    "11111111", --  442 - 0x1ba  :  255 - 0xff
    "11111110", --  443 - 0x1bb  :  254 - 0xfe
    "11111110", --  444 - 0x1bc  :  254 - 0xfe
    "11111111", --  445 - 0x1bd  :  255 - 0xff
    "11101100", --  446 - 0x1be  :  236 - 0xec
    "11101001", --  447 - 0x1bf  :  233 - 0xe9
    "11111010", --  448 - 0x1c0  :  250 - 0xfa -- line 0xe
    "11111100", --  449 - 0x1c1  :  252 - 0xfc
    "11111111", --  450 - 0x1c2  :  255 - 0xff
    "11111111", --  451 - 0x1c3  :  255 - 0xff
    "11111111", --  452 - 0x1c4  :  255 - 0xff
    "11111111", --  453 - 0x1c5  :  255 - 0xff
    "11101100", --  454 - 0x1c6  :  236 - 0xec
    "11111010", --  455 - 0x1c7  :  250 - 0xfa
    "11111010", --  456 - 0x1c8  :  250 - 0xfa
    "11111010", --  457 - 0x1c9  :  250 - 0xfa
    "11101001", --  458 - 0x1ca  :  233 - 0xe9
    "11111010", --  459 - 0x1cb  :  250 - 0xfa
    "11111010", --  460 - 0x1cc  :  250 - 0xfa
    "11111010", --  461 - 0x1cd  :  250 - 0xfa
    "11111010", --  462 - 0x1ce  :  250 - 0xfa
    "11111010", --  463 - 0x1cf  :  250 - 0xfa
    "11111010", --  464 - 0x1d0  :  250 - 0xfa
    "11111010", --  465 - 0x1d1  :  250 - 0xfa
    "11111010", --  466 - 0x1d2  :  250 - 0xfa
    "11111100", --  467 - 0x1d3  :  252 - 0xfc
    "11111111", --  468 - 0x1d4  :  255 - 0xff
    "11111111", --  469 - 0x1d5  :  255 - 0xff
    "11111111", --  470 - 0x1d6  :  255 - 0xff
    "11111111", --  471 - 0x1d7  :  255 - 0xff
    "11111111", --  472 - 0x1d8  :  255 - 0xff
    "11111111", --  473 - 0x1d9  :  255 - 0xff
    "11111111", --  474 - 0x1da  :  255 - 0xff
    "11111111", --  475 - 0x1db  :  255 - 0xff
    "11111111", --  476 - 0x1dc  :  255 - 0xff
    "11111111", --  477 - 0x1dd  :  255 - 0xff
    "11101100", --  478 - 0x1de  :  236 - 0xec
    "11111010", --  479 - 0x1df  :  250 - 0xfa
    "11101010", --  480 - 0x1e0  :  234 - 0xea -- line 0xf
    "11111100", --  481 - 0x1e1  :  252 - 0xfc
    "11111111", --  482 - 0x1e2  :  255 - 0xff
    "11111110", --  483 - 0x1e3  :  254 - 0xfe
    "11111110", --  484 - 0x1e4  :  254 - 0xfe
    "11111111", --  485 - 0x1e5  :  255 - 0xff
    "11110101", --  486 - 0x1e6  :  245 - 0xf5
    "11111011", --  487 - 0x1e7  :  251 - 0xfb
    "11111011", --  488 - 0x1e8  :  251 - 0xfb
    "11111011", --  489 - 0x1e9  :  251 - 0xfb
    "11111011", --  490 - 0x1ea  :  251 - 0xfb
    "11111011", --  491 - 0x1eb  :  251 - 0xfb
    "11101000", --  492 - 0x1ec  :  232 - 0xe8
    "11111010", --  493 - 0x1ed  :  250 - 0xfa
    "11111010", --  494 - 0x1ee  :  250 - 0xfa
    "11111010", --  495 - 0x1ef  :  250 - 0xfa
    "11101001", --  496 - 0x1f0  :  233 - 0xe9
    "11111010", --  497 - 0x1f1  :  250 - 0xfa
    "11111010", --  498 - 0x1f2  :  250 - 0xfa
    "11111100", --  499 - 0x1f3  :  252 - 0xfc
    "11111111", --  500 - 0x1f4  :  255 - 0xff
    "11111111", --  501 - 0x1f5  :  255 - 0xff
    "11111111", --  502 - 0x1f6  :  255 - 0xff
    "11111111", --  503 - 0x1f7  :  255 - 0xff
    "11111101", --  504 - 0x1f8  :  253 - 0xfd
    "11111111", --  505 - 0x1f9  :  255 - 0xff
    "11111101", --  506 - 0x1fa  :  253 - 0xfd
    "11111111", --  507 - 0x1fb  :  255 - 0xff
    "11111111", --  508 - 0x1fc  :  255 - 0xff
    "11111111", --  509 - 0x1fd  :  255 - 0xff
    "11101100", --  510 - 0x1fe  :  236 - 0xec
    "11111010", --  511 - 0x1ff  :  250 - 0xfa
    "11111010", --  512 - 0x200  :  250 - 0xfa -- line 0x10
    "11111100", --  513 - 0x201  :  252 - 0xfc
    "11111111", --  514 - 0x202  :  255 - 0xff
    "11111111", --  515 - 0x203  :  255 - 0xff
    "11111111", --  516 - 0x204  :  255 - 0xff
    "11111111", --  517 - 0x205  :  255 - 0xff
    "11111111", --  518 - 0x206  :  255 - 0xff
    "11111111", --  519 - 0x207  :  255 - 0xff
    "11111111", --  520 - 0x208  :  255 - 0xff
    "11111111", --  521 - 0x209  :  255 - 0xff
    "11111111", --  522 - 0x20a  :  255 - 0xff
    "11111111", --  523 - 0x20b  :  255 - 0xff
    "11101100", --  524 - 0x20c  :  236 - 0xec
    "11111010", --  525 - 0x20d  :  250 - 0xfa
    "11111010", --  526 - 0x20e  :  250 - 0xfa
    "11111010", --  527 - 0x20f  :  250 - 0xfa
    "11111010", --  528 - 0x210  :  250 - 0xfa
    "11111010", --  529 - 0x211  :  250 - 0xfa
    "11111010", --  530 - 0x212  :  250 - 0xfa
    "11111100", --  531 - 0x213  :  252 - 0xfc
    "11111111", --  532 - 0x214  :  255 - 0xff
    "11111111", --  533 - 0x215  :  255 - 0xff
    "11111111", --  534 - 0x216  :  255 - 0xff
    "11111111", --  535 - 0x217  :  255 - 0xff
    "11111101", --  536 - 0x218  :  253 - 0xfd
    "11111111", --  537 - 0x219  :  255 - 0xff
    "11111101", --  538 - 0x21a  :  253 - 0xfd
    "11111111", --  539 - 0x21b  :  255 - 0xff
    "11111111", --  540 - 0x21c  :  255 - 0xff
    "11111111", --  541 - 0x21d  :  255 - 0xff
    "11101100", --  542 - 0x21e  :  236 - 0xec
    "11101010", --  543 - 0x21f  :  234 - 0xea
    "11111010", --  544 - 0x220  :  250 - 0xfa -- line 0x11
    "11111100", --  545 - 0x221  :  252 - 0xfc
    "11111111", --  546 - 0x222  :  255 - 0xff
    "11111111", --  547 - 0x223  :  255 - 0xff
    "11111111", --  548 - 0x224  :  255 - 0xff
    "11111111", --  549 - 0x225  :  255 - 0xff
    "11111101", --  550 - 0x226  :  253 - 0xfd
    "11111111", --  551 - 0x227  :  255 - 0xff
    "11111101", --  552 - 0x228  :  253 - 0xfd
    "11111111", --  553 - 0x229  :  255 - 0xff
    "11111111", --  554 - 0x22a  :  255 - 0xff
    "11111111", --  555 - 0x22b  :  255 - 0xff
    "11101100", --  556 - 0x22c  :  236 - 0xec
    "11111010", --  557 - 0x22d  :  250 - 0xfa
    "11111010", --  558 - 0x22e  :  250 - 0xfa
    "11111010", --  559 - 0x22f  :  250 - 0xfa
    "11111010", --  560 - 0x230  :  250 - 0xfa
    "11111010", --  561 - 0x231  :  250 - 0xfa
    "11111010", --  562 - 0x232  :  250 - 0xfa
    "11111100", --  563 - 0x233  :  252 - 0xfc
    "11111111", --  564 - 0x234  :  255 - 0xff
    "11111110", --  565 - 0x235  :  254 - 0xfe
    "11111110", --  566 - 0x236  :  254 - 0xfe
    "11111111", --  567 - 0x237  :  255 - 0xff
    "11111111", --  568 - 0x238  :  255 - 0xff
    "11111111", --  569 - 0x239  :  255 - 0xff
    "11111111", --  570 - 0x23a  :  255 - 0xff
    "11111111", --  571 - 0x23b  :  255 - 0xff
    "11111111", --  572 - 0x23c  :  255 - 0xff
    "11111111", --  573 - 0x23d  :  255 - 0xff
    "11101100", --  574 - 0x23e  :  236 - 0xec
    "11111010", --  575 - 0x23f  :  250 - 0xfa
    "11111010", --  576 - 0x240  :  250 - 0xfa -- line 0x12
    "11111100", --  577 - 0x241  :  252 - 0xfc
    "11111111", --  578 - 0x242  :  255 - 0xff
    "11111111", --  579 - 0x243  :  255 - 0xff
    "11111111", --  580 - 0x244  :  255 - 0xff
    "11111111", --  581 - 0x245  :  255 - 0xff
    "11111101", --  582 - 0x246  :  253 - 0xfd
    "11111111", --  583 - 0x247  :  255 - 0xff
    "11111101", --  584 - 0x248  :  253 - 0xfd
    "11111111", --  585 - 0x249  :  255 - 0xff
    "11111111", --  586 - 0x24a  :  255 - 0xff
    "11111111", --  587 - 0x24b  :  255 - 0xff
    "11101100", --  588 - 0x24c  :  236 - 0xec
    "11111010", --  589 - 0x24d  :  250 - 0xfa
    "11111010", --  590 - 0x24e  :  250 - 0xfa
    "11101001", --  591 - 0x24f  :  233 - 0xe9
    "11111010", --  592 - 0x250  :  250 - 0xfa
    "11111010", --  593 - 0x251  :  250 - 0xfa
    "11111010", --  594 - 0x252  :  250 - 0xfa
    "11111100", --  595 - 0x253  :  252 - 0xfc
    "11111111", --  596 - 0x254  :  255 - 0xff
    "11111111", --  597 - 0x255  :  255 - 0xff
    "11111111", --  598 - 0x256  :  255 - 0xff
    "11111111", --  599 - 0x257  :  255 - 0xff
    "11100101", --  600 - 0x258  :  229 - 0xe5
    "11101011", --  601 - 0x259  :  235 - 0xeb
    "11101011", --  602 - 0x25a  :  235 - 0xeb
    "11101011", --  603 - 0x25b  :  235 - 0xeb
    "11101011", --  604 - 0x25c  :  235 - 0xeb
    "11101011", --  605 - 0x25d  :  235 - 0xeb
    "11111000", --  606 - 0x25e  :  248 - 0xf8
    "11111010", --  607 - 0x25f  :  250 - 0xfa
    "11111010", --  608 - 0x260  :  250 - 0xfa -- line 0x13
    "11111100", --  609 - 0x261  :  252 - 0xfc
    "11111111", --  610 - 0x262  :  255 - 0xff
    "11111111", --  611 - 0x263  :  255 - 0xff
    "11111111", --  612 - 0x264  :  255 - 0xff
    "11111111", --  613 - 0x265  :  255 - 0xff
    "11111111", --  614 - 0x266  :  255 - 0xff
    "11111111", --  615 - 0x267  :  255 - 0xff
    "11111111", --  616 - 0x268  :  255 - 0xff
    "11111111", --  617 - 0x269  :  255 - 0xff
    "11111111", --  618 - 0x26a  :  255 - 0xff
    "11111111", --  619 - 0x26b  :  255 - 0xff
    "11101100", --  620 - 0x26c  :  236 - 0xec
    "11111010", --  621 - 0x26d  :  250 - 0xfa
    "11111010", --  622 - 0x26e  :  250 - 0xfa
    "11111010", --  623 - 0x26f  :  250 - 0xfa
    "11111010", --  624 - 0x270  :  250 - 0xfa
    "11111010", --  625 - 0x271  :  250 - 0xfa
    "11111010", --  626 - 0x272  :  250 - 0xfa
    "11111100", --  627 - 0x273  :  252 - 0xfc
    "11111111", --  628 - 0x274  :  255 - 0xff
    "11111110", --  629 - 0x275  :  254 - 0xfe
    "11111110", --  630 - 0x276  :  254 - 0xfe
    "11111111", --  631 - 0x277  :  255 - 0xff
    "11110101", --  632 - 0x278  :  245 - 0xf5
    "11111011", --  633 - 0x279  :  251 - 0xfb
    "11111011", --  634 - 0x27a  :  251 - 0xfb
    "11111011", --  635 - 0x27b  :  251 - 0xfb
    "11111011", --  636 - 0x27c  :  251 - 0xfb
    "11111011", --  637 - 0x27d  :  251 - 0xfb
    "11101000", --  638 - 0x27e  :  232 - 0xe8
    "11111010", --  639 - 0x27f  :  250 - 0xfa
    "11111010", --  640 - 0x280  :  250 - 0xfa -- line 0x14
    "11110111", --  641 - 0x281  :  247 - 0xf7
    "11101011", --  642 - 0x282  :  235 - 0xeb
    "11101011", --  643 - 0x283  :  235 - 0xeb
    "11101011", --  644 - 0x284  :  235 - 0xeb
    "11101011", --  645 - 0x285  :  235 - 0xeb
    "11101011", --  646 - 0x286  :  235 - 0xeb
    "11100110", --  647 - 0x287  :  230 - 0xe6
    "11111111", --  648 - 0x288  :  255 - 0xff
    "11111111", --  649 - 0x289  :  255 - 0xff
    "11111111", --  650 - 0x28a  :  255 - 0xff
    "11111111", --  651 - 0x28b  :  255 - 0xff
    "11101100", --  652 - 0x28c  :  236 - 0xec
    "11111010", --  653 - 0x28d  :  250 - 0xfa
    "11111010", --  654 - 0x28e  :  250 - 0xfa
    "11101001", --  655 - 0x28f  :  233 - 0xe9
    "11111010", --  656 - 0x290  :  250 - 0xfa
    "11111010", --  657 - 0x291  :  250 - 0xfa
    "11111010", --  658 - 0x292  :  250 - 0xfa
    "11111100", --  659 - 0x293  :  252 - 0xfc
    "11111111", --  660 - 0x294  :  255 - 0xff
    "11111111", --  661 - 0x295  :  255 - 0xff
    "11111111", --  662 - 0x296  :  255 - 0xff
    "11111111", --  663 - 0x297  :  255 - 0xff
    "11111111", --  664 - 0x298  :  255 - 0xff
    "11111111", --  665 - 0x299  :  255 - 0xff
    "11111111", --  666 - 0x29a  :  255 - 0xff
    "11111111", --  667 - 0x29b  :  255 - 0xff
    "11111111", --  668 - 0x29c  :  255 - 0xff
    "11111111", --  669 - 0x29d  :  255 - 0xff
    "11101100", --  670 - 0x29e  :  236 - 0xec
    "11111010", --  671 - 0x29f  :  250 - 0xfa
    "11111010", --  672 - 0x2a0  :  250 - 0xfa -- line 0x15
    "11111010", --  673 - 0x2a1  :  250 - 0xfa
    "11101010", --  674 - 0x2a2  :  234 - 0xea
    "11101001", --  675 - 0x2a3  :  233 - 0xe9
    "11111010", --  676 - 0x2a4  :  250 - 0xfa
    "11111010", --  677 - 0x2a5  :  250 - 0xfa
    "11111010", --  678 - 0x2a6  :  250 - 0xfa
    "11111100", --  679 - 0x2a7  :  252 - 0xfc
    "11111111", --  680 - 0x2a8  :  255 - 0xff
    "11111110", --  681 - 0x2a9  :  254 - 0xfe
    "11111110", --  682 - 0x2aa  :  254 - 0xfe
    "11111111", --  683 - 0x2ab  :  255 - 0xff
    "11101100", --  684 - 0x2ac  :  236 - 0xec
    "11111010", --  685 - 0x2ad  :  250 - 0xfa
    "11111010", --  686 - 0x2ae  :  250 - 0xfa
    "11111010", --  687 - 0x2af  :  250 - 0xfa
    "11111010", --  688 - 0x2b0  :  250 - 0xfa
    "11101001", --  689 - 0x2b1  :  233 - 0xe9
    "11111010", --  690 - 0x2b2  :  250 - 0xfa
    "11111100", --  691 - 0x2b3  :  252 - 0xfc
    "11111111", --  692 - 0x2b4  :  255 - 0xff
    "11111111", --  693 - 0x2b5  :  255 - 0xff
    "11111111", --  694 - 0x2b6  :  255 - 0xff
    "11111111", --  695 - 0x2b7  :  255 - 0xff
    "11111111", --  696 - 0x2b8  :  255 - 0xff
    "11111111", --  697 - 0x2b9  :  255 - 0xff
    "11111111", --  698 - 0x2ba  :  255 - 0xff
    "11111111", --  699 - 0x2bb  :  255 - 0xff
    "11111111", --  700 - 0x2bc  :  255 - 0xff
    "11111111", --  701 - 0x2bd  :  255 - 0xff
    "11101100", --  702 - 0x2be  :  236 - 0xec
    "11111010", --  703 - 0x2bf  :  250 - 0xfa
    "11111010", --  704 - 0x2c0  :  250 - 0xfa -- line 0x16
    "11111010", --  705 - 0x2c1  :  250 - 0xfa
    "11111010", --  706 - 0x2c2  :  250 - 0xfa
    "11111010", --  707 - 0x2c3  :  250 - 0xfa
    "11111010", --  708 - 0x2c4  :  250 - 0xfa
    "11111010", --  709 - 0x2c5  :  250 - 0xfa
    "11101001", --  710 - 0x2c6  :  233 - 0xe9
    "11111100", --  711 - 0x2c7  :  252 - 0xfc
    "11111111", --  712 - 0x2c8  :  255 - 0xff
    "11111111", --  713 - 0x2c9  :  255 - 0xff
    "11111111", --  714 - 0x2ca  :  255 - 0xff
    "11111111", --  715 - 0x2cb  :  255 - 0xff
    "11101100", --  716 - 0x2cc  :  236 - 0xec
    "11111010", --  717 - 0x2cd  :  250 - 0xfa
    "11111010", --  718 - 0x2ce  :  250 - 0xfa
    "11111010", --  719 - 0x2cf  :  250 - 0xfa
    "11111010", --  720 - 0x2d0  :  250 - 0xfa
    "11111010", --  721 - 0x2d1  :  250 - 0xfa
    "11111010", --  722 - 0x2d2  :  250 - 0xfa
    "11110111", --  723 - 0x2d3  :  247 - 0xf7
    "11101011", --  724 - 0x2d4  :  235 - 0xeb
    "11101011", --  725 - 0x2d5  :  235 - 0xeb
    "11101011", --  726 - 0x2d6  :  235 - 0xeb
    "11101011", --  727 - 0x2d7  :  235 - 0xeb
    "11101011", --  728 - 0x2d8  :  235 - 0xeb
    "11100110", --  729 - 0x2d9  :  230 - 0xe6
    "11111111", --  730 - 0x2da  :  255 - 0xff
    "11111111", --  731 - 0x2db  :  255 - 0xff
    "11111111", --  732 - 0x2dc  :  255 - 0xff
    "11111111", --  733 - 0x2dd  :  255 - 0xff
    "11101100", --  734 - 0x2de  :  236 - 0xec
    "11111010", --  735 - 0x2df  :  250 - 0xfa
    "11111010", --  736 - 0x2e0  :  250 - 0xfa -- line 0x17
    "11111010", --  737 - 0x2e1  :  250 - 0xfa
    "11101001", --  738 - 0x2e2  :  233 - 0xe9
    "11111010", --  739 - 0x2e3  :  250 - 0xfa
    "11111010", --  740 - 0x2e4  :  250 - 0xfa
    "11111010", --  741 - 0x2e5  :  250 - 0xfa
    "11111010", --  742 - 0x2e6  :  250 - 0xfa
    "11111100", --  743 - 0x2e7  :  252 - 0xfc
    "11111111", --  744 - 0x2e8  :  255 - 0xff
    "11111110", --  745 - 0x2e9  :  254 - 0xfe
    "11111110", --  746 - 0x2ea  :  254 - 0xfe
    "11111111", --  747 - 0x2eb  :  255 - 0xff
    "11110101", --  748 - 0x2ec  :  245 - 0xf5
    "11111011", --  749 - 0x2ed  :  251 - 0xfb
    "11111011", --  750 - 0x2ee  :  251 - 0xfb
    "11111011", --  751 - 0x2ef  :  251 - 0xfb
    "11111011", --  752 - 0x2f0  :  251 - 0xfb
    "11111011", --  753 - 0x2f1  :  251 - 0xfb
    "11111011", --  754 - 0x2f2  :  251 - 0xfb
    "11111011", --  755 - 0x2f3  :  251 - 0xfb
    "11111011", --  756 - 0x2f4  :  251 - 0xfb
    "11111011", --  757 - 0x2f5  :  251 - 0xfb
    "11111011", --  758 - 0x2f6  :  251 - 0xfb
    "11111011", --  759 - 0x2f7  :  251 - 0xfb
    "11111011", --  760 - 0x2f8  :  251 - 0xfb
    "11110110", --  761 - 0x2f9  :  246 - 0xf6
    "11111111", --  762 - 0x2fa  :  255 - 0xff
    "11111110", --  763 - 0x2fb  :  254 - 0xfe
    "11111110", --  764 - 0x2fc  :  254 - 0xfe
    "11111111", --  765 - 0x2fd  :  255 - 0xff
    "11101100", --  766 - 0x2fe  :  236 - 0xec
    "11111010", --  767 - 0x2ff  :  250 - 0xfa
    "11111010", --  768 - 0x300  :  250 - 0xfa -- line 0x18
    "11111010", --  769 - 0x301  :  250 - 0xfa
    "11111010", --  770 - 0x302  :  250 - 0xfa
    "11111010", --  771 - 0x303  :  250 - 0xfa
    "11111010", --  772 - 0x304  :  250 - 0xfa
    "11111010", --  773 - 0x305  :  250 - 0xfa
    "11111010", --  774 - 0x306  :  250 - 0xfa
    "11111100", --  775 - 0x307  :  252 - 0xfc
    "11111111", --  776 - 0x308  :  255 - 0xff
    "11111111", --  777 - 0x309  :  255 - 0xff
    "11111111", --  778 - 0x30a  :  255 - 0xff
    "11111111", --  779 - 0x30b  :  255 - 0xff
    "11111111", --  780 - 0x30c  :  255 - 0xff
    "11111111", --  781 - 0x30d  :  255 - 0xff
    "11111111", --  782 - 0x30e  :  255 - 0xff
    "11111111", --  783 - 0x30f  :  255 - 0xff
    "11111111", --  784 - 0x310  :  255 - 0xff
    "11111111", --  785 - 0x311  :  255 - 0xff
    "11101111", --  786 - 0x312  :  239 - 0xef
    "11111111", --  787 - 0x313  :  255 - 0xff
    "11111111", --  788 - 0x314  :  255 - 0xff
    "11111111", --  789 - 0x315  :  255 - 0xff
    "11111111", --  790 - 0x316  :  255 - 0xff
    "11111111", --  791 - 0x317  :  255 - 0xff
    "11111111", --  792 - 0x318  :  255 - 0xff
    "11111111", --  793 - 0x319  :  255 - 0xff
    "11111111", --  794 - 0x31a  :  255 - 0xff
    "11111111", --  795 - 0x31b  :  255 - 0xff
    "11111111", --  796 - 0x31c  :  255 - 0xff
    "11111111", --  797 - 0x31d  :  255 - 0xff
    "11101100", --  798 - 0x31e  :  236 - 0xec
    "11101001", --  799 - 0x31f  :  233 - 0xe9
    "11101010", --  800 - 0x320  :  234 - 0xea -- line 0x19
    "00001101", --  801 - 0x321  :   13 - 0xd
    "00000001", --  802 - 0x322  :    1 - 0x1
    "00000010", --  803 - 0x323  :    2 - 0x2
    "00000010", --  804 - 0x324  :    2 - 0x2
    "11111010", --  805 - 0x325  :  250 - 0xfa
    "11111010", --  806 - 0x326  :  250 - 0xfa
    "11111100", --  807 - 0x327  :  252 - 0xfc
    "11111111", --  808 - 0x328  :  255 - 0xff
    "11111111", --  809 - 0x329  :  255 - 0xff
    "11111111", --  810 - 0x32a  :  255 - 0xff
    "11111111", --  811 - 0x32b  :  255 - 0xff
    "11111101", --  812 - 0x32c  :  253 - 0xfd
    "11111111", --  813 - 0x32d  :  255 - 0xff
    "11111101", --  814 - 0x32e  :  253 - 0xfd
    "11111111", --  815 - 0x32f  :  255 - 0xff
    "11111101", --  816 - 0x330  :  253 - 0xfd
    "11111111", --  817 - 0x331  :  255 - 0xff
    "11101111", --  818 - 0x332  :  239 - 0xef
    "11111111", --  819 - 0x333  :  255 - 0xff
    "11111101", --  820 - 0x334  :  253 - 0xfd
    "11111111", --  821 - 0x335  :  255 - 0xff
    "11111101", --  822 - 0x336  :  253 - 0xfd
    "11111111", --  823 - 0x337  :  255 - 0xff
    "11111101", --  824 - 0x338  :  253 - 0xfd
    "11111111", --  825 - 0x339  :  255 - 0xff
    "11111111", --  826 - 0x33a  :  255 - 0xff
    "11111111", --  827 - 0x33b  :  255 - 0xff
    "11111111", --  828 - 0x33c  :  255 - 0xff
    "11111111", --  829 - 0x33d  :  255 - 0xff
    "11101100", --  830 - 0x33e  :  236 - 0xec
    "11111010", --  831 - 0x33f  :  250 - 0xfa
    "11111010", --  832 - 0x340  :  250 - 0xfa -- line 0x1a
    "11111010", --  833 - 0x341  :  250 - 0xfa
    "11111010", --  834 - 0x342  :  250 - 0xfa
    "11111010", --  835 - 0x343  :  250 - 0xfa
    "11111010", --  836 - 0x344  :  250 - 0xfa
    "11111010", --  837 - 0x345  :  250 - 0xfa
    "11111010", --  838 - 0x346  :  250 - 0xfa
    "11111100", --  839 - 0x347  :  252 - 0xfc
    "11111111", --  840 - 0x348  :  255 - 0xff
    "11111111", --  841 - 0x349  :  255 - 0xff
    "11111111", --  842 - 0x34a  :  255 - 0xff
    "11111111", --  843 - 0x34b  :  255 - 0xff
    "11111101", --  844 - 0x34c  :  253 - 0xfd
    "11111111", --  845 - 0x34d  :  255 - 0xff
    "11111101", --  846 - 0x34e  :  253 - 0xfd
    "11111111", --  847 - 0x34f  :  255 - 0xff
    "11111101", --  848 - 0x350  :  253 - 0xfd
    "11111111", --  849 - 0x351  :  255 - 0xff
    "11101111", --  850 - 0x352  :  239 - 0xef
    "11111111", --  851 - 0x353  :  255 - 0xff
    "11111101", --  852 - 0x354  :  253 - 0xfd
    "11111111", --  853 - 0x355  :  255 - 0xff
    "11111101", --  854 - 0x356  :  253 - 0xfd
    "11111111", --  855 - 0x357  :  255 - 0xff
    "11111101", --  856 - 0x358  :  253 - 0xfd
    "11111111", --  857 - 0x359  :  255 - 0xff
    "11111111", --  858 - 0x35a  :  255 - 0xff
    "11111111", --  859 - 0x35b  :  255 - 0xff
    "11111111", --  860 - 0x35c  :  255 - 0xff
    "11111111", --  861 - 0x35d  :  255 - 0xff
    "11101100", --  862 - 0x35e  :  236 - 0xec
    "11111010", --  863 - 0x35f  :  250 - 0xfa
    "11111010", --  864 - 0x360  :  250 - 0xfa -- line 0x1b
    "00001111", --  865 - 0x361  :   15 - 0xf
    "00000001", --  866 - 0x362  :    1 - 0x1
    "00010000", --  867 - 0x363  :   16 - 0x10
    "00000011", --  868 - 0x364  :    3 - 0x3
    "11111010", --  869 - 0x365  :  250 - 0xfa
    "11111010", --  870 - 0x366  :  250 - 0xfa
    "11111100", --  871 - 0x367  :  252 - 0xfc
    "11111111", --  872 - 0x368  :  255 - 0xff
    "11111111", --  873 - 0x369  :  255 - 0xff
    "11111111", --  874 - 0x36a  :  255 - 0xff
    "11111111", --  875 - 0x36b  :  255 - 0xff
    "11111111", --  876 - 0x36c  :  255 - 0xff
    "11111111", --  877 - 0x36d  :  255 - 0xff
    "11111111", --  878 - 0x36e  :  255 - 0xff
    "11111111", --  879 - 0x36f  :  255 - 0xff
    "11111111", --  880 - 0x370  :  255 - 0xff
    "11111111", --  881 - 0x371  :  255 - 0xff
    "11101111", --  882 - 0x372  :  239 - 0xef
    "11111111", --  883 - 0x373  :  255 - 0xff
    "11111111", --  884 - 0x374  :  255 - 0xff
    "11111111", --  885 - 0x375  :  255 - 0xff
    "11111111", --  886 - 0x376  :  255 - 0xff
    "11111111", --  887 - 0x377  :  255 - 0xff
    "11111111", --  888 - 0x378  :  255 - 0xff
    "11111111", --  889 - 0x379  :  255 - 0xff
    "11111111", --  890 - 0x37a  :  255 - 0xff
    "11111111", --  891 - 0x37b  :  255 - 0xff
    "11111111", --  892 - 0x37c  :  255 - 0xff
    "11111111", --  893 - 0x37d  :  255 - 0xff
    "11101100", --  894 - 0x37e  :  236 - 0xec
    "11111010", --  895 - 0x37f  :  250 - 0xfa
    "11111010", --  896 - 0x380  :  250 - 0xfa -- line 0x1c
    "11111010", --  897 - 0x381  :  250 - 0xfa
    "11111001", --  898 - 0x382  :  249 - 0xf9
    "11111010", --  899 - 0x383  :  250 - 0xfa
    "11111010", --  900 - 0x384  :  250 - 0xfa
    "11101010", --  901 - 0x385  :  234 - 0xea
    "11111010", --  902 - 0x386  :  250 - 0xfa
    "11110111", --  903 - 0x387  :  247 - 0xf7
    "11101011", --  904 - 0x388  :  235 - 0xeb
    "11101011", --  905 - 0x389  :  235 - 0xeb
    "11101011", --  906 - 0x38a  :  235 - 0xeb
    "11101011", --  907 - 0x38b  :  235 - 0xeb
    "11101011", --  908 - 0x38c  :  235 - 0xeb
    "11101011", --  909 - 0x38d  :  235 - 0xeb
    "11101011", --  910 - 0x38e  :  235 - 0xeb
    "11101011", --  911 - 0x38f  :  235 - 0xeb
    "11101011", --  912 - 0x390  :  235 - 0xeb
    "11101011", --  913 - 0x391  :  235 - 0xeb
    "11101011", --  914 - 0x392  :  235 - 0xeb
    "11101011", --  915 - 0x393  :  235 - 0xeb
    "11101011", --  916 - 0x394  :  235 - 0xeb
    "11101011", --  917 - 0x395  :  235 - 0xeb
    "11101011", --  918 - 0x396  :  235 - 0xeb
    "11101011", --  919 - 0x397  :  235 - 0xeb
    "11101011", --  920 - 0x398  :  235 - 0xeb
    "11101011", --  921 - 0x399  :  235 - 0xeb
    "11101011", --  922 - 0x39a  :  235 - 0xeb
    "11101011", --  923 - 0x39b  :  235 - 0xeb
    "11101011", --  924 - 0x39c  :  235 - 0xeb
    "11101011", --  925 - 0x39d  :  235 - 0xeb
    "11111000", --  926 - 0x39e  :  248 - 0xf8
    "11111010", --  927 - 0x39f  :  250 - 0xfa
    "11111010", --  928 - 0x3a0  :  250 - 0xfa -- line 0x1d
    "11111001", --  929 - 0x3a1  :  249 - 0xf9
    "11111010", --  930 - 0x3a2  :  250 - 0xfa
    "11111010", --  931 - 0x3a3  :  250 - 0xfa
    "11111010", --  932 - 0x3a4  :  250 - 0xfa
    "11111010", --  933 - 0x3a5  :  250 - 0xfa
    "11111010", --  934 - 0x3a6  :  250 - 0xfa
    "11111010", --  935 - 0x3a7  :  250 - 0xfa
    "11111010", --  936 - 0x3a8  :  250 - 0xfa
    "11111010", --  937 - 0x3a9  :  250 - 0xfa
    "11111010", --  938 - 0x3aa  :  250 - 0xfa
    "11111010", --  939 - 0x3ab  :  250 - 0xfa
    "11111010", --  940 - 0x3ac  :  250 - 0xfa
    "11111010", --  941 - 0x3ad  :  250 - 0xfa
    "11111010", --  942 - 0x3ae  :  250 - 0xfa
    "11111010", --  943 - 0x3af  :  250 - 0xfa
    "11111010", --  944 - 0x3b0  :  250 - 0xfa
    "11111010", --  945 - 0x3b1  :  250 - 0xfa
    "11111010", --  946 - 0x3b2  :  250 - 0xfa
    "11111010", --  947 - 0x3b3  :  250 - 0xfa
    "11111010", --  948 - 0x3b4  :  250 - 0xfa
    "11101001", --  949 - 0x3b5  :  233 - 0xe9
    "11111010", --  950 - 0x3b6  :  250 - 0xfa
    "11111010", --  951 - 0x3b7  :  250 - 0xfa
    "11111010", --  952 - 0x3b8  :  250 - 0xfa
    "11111010", --  953 - 0x3b9  :  250 - 0xfa
    "11111010", --  954 - 0x3ba  :  250 - 0xfa
    "11111010", --  955 - 0x3bb  :  250 - 0xfa
    "11101010", --  956 - 0x3bc  :  234 - 0xea
    "11111010", --  957 - 0x3bd  :  250 - 0xfa
    "11111010", --  958 - 0x3be  :  250 - 0xfa
    "11111010", --  959 - 0x3bf  :  250 - 0xfa
        ---- Attribute Table 0----
    "00010101", --  960 - 0x3c0  :   21 - 0x15
    "00000101", --  961 - 0x3c1  :    5 - 0x5
    "00000101", --  962 - 0x3c2  :    5 - 0x5
    "00000101", --  963 - 0x3c3  :    5 - 0x5
    "00000101", --  964 - 0x3c4  :    5 - 0x5
    "01000101", --  965 - 0x3c5  :   69 - 0x45
    "01010101", --  966 - 0x3c6  :   85 - 0x55
    "01010101", --  967 - 0x3c7  :   85 - 0x55
    "00010001", --  968 - 0x3c8  :   17 - 0x11
    "01000000", --  969 - 0x3c9  :   64 - 0x40
    "01010000", --  970 - 0x3ca  :   80 - 0x50
    "01010000", --  971 - 0x3cb  :   80 - 0x50
    "00010000", --  972 - 0x3cc  :   16 - 0x10
    "00000100", --  973 - 0x3cd  :    4 - 0x4
    "00000101", --  974 - 0x3ce  :    5 - 0x5
    "01000101", --  975 - 0x3cf  :   69 - 0x45
    "00010001", --  976 - 0x3d0  :   17 - 0x11
    "01000100", --  977 - 0x3d1  :   68 - 0x44
    "01010101", --  978 - 0x3d2  :   85 - 0x55
    "01010101", --  979 - 0x3d3  :   85 - 0x55
    "01010001", --  980 - 0x3d4  :   81 - 0x51
    "01010000", --  981 - 0x3d5  :   80 - 0x50
    "00010000", --  982 - 0x3d6  :   16 - 0x10
    "01000100", --  983 - 0x3d7  :   68 - 0x44
    "00010001", --  984 - 0x3d8  :   17 - 0x11
    "01000100", --  985 - 0x3d9  :   68 - 0x44
    "01010101", --  986 - 0x3da  :   85 - 0x55
    "01010101", --  987 - 0x3db  :   85 - 0x55
    "01010101", --  988 - 0x3dc  :   85 - 0x55
    "00000101", --  989 - 0x3dd  :    5 - 0x5
    "00000001", --  990 - 0x3de  :    1 - 0x1
    "01000100", --  991 - 0x3df  :   68 - 0x44
    "00010001", --  992 - 0x3e0  :   17 - 0x11
    "00000000", --  993 - 0x3e1  :    0 - 0x0
    "00000000", --  994 - 0x3e2  :    0 - 0x0
    "01010101", --  995 - 0x3e3  :   85 - 0x55
    "01010101", --  996 - 0x3e4  :   85 - 0x55
    "00000000", --  997 - 0x3e5  :    0 - 0x0
    "01010000", --  998 - 0x3e6  :   80 - 0x50
    "01010100", --  999 - 0x3e7  :   84 - 0x54
    "01010101", -- 1000 - 0x3e8  :   85 - 0x55
    "01010101", -- 1001 - 0x3e9  :   85 - 0x55
    "00000000", -- 1002 - 0x3ea  :    0 - 0x0
    "01010101", -- 1003 - 0x3eb  :   85 - 0x55
    "01010101", -- 1004 - 0x3ec  :   85 - 0x55
    "01010000", -- 1005 - 0x3ed  :   80 - 0x50
    "00010000", -- 1006 - 0x3ee  :   16 - 0x10
    "01000100", -- 1007 - 0x3ef  :   68 - 0x44
    "01010101", -- 1008 - 0x3f0  :   85 - 0x55
    "01010101", -- 1009 - 0x3f1  :   85 - 0x55
    "00000000", -- 1010 - 0x3f2  :    0 - 0x0
    "00000000", -- 1011 - 0x3f3  :    0 - 0x0
    "00000000", -- 1012 - 0x3f4  :    0 - 0x0
    "00000000", -- 1013 - 0x3f5  :    0 - 0x0
    "00000000", -- 1014 - 0x3f6  :    0 - 0x0
    "01000100", -- 1015 - 0x3f7  :   68 - 0x44
    "00000101", -- 1016 - 0x3f8  :    5 - 0x5
    "00000101", -- 1017 - 0x3f9  :    5 - 0x5
    "00000101", -- 1018 - 0x3fa  :    5 - 0x5
    "00000101", -- 1019 - 0x3fb  :    5 - 0x5
    "00000101", -- 1020 - 0x3fc  :    5 - 0x5
    "00000101", -- 1021 - 0x3fd  :    5 - 0x5
    "00000101", -- 1022 - 0x3fe  :    5 - 0x5
    "00000101"  -- 1023 - 0x3ff  :    5 - 0x5
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
