//- Autcmatically generated verilog ROM from a NES memory file----
//-   PATTERN TABLE
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


//-  Original memory dump file name: nova_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_PTABLE_NOVA
  (
     input     clk,   // clock
     input      [13-1:0] addr,  //8192 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Pattern Table 0---------
      13'h0: dout <= 8'b11111111; //    0 : 255 - 0xff -- Sprite 0x0
      13'h1: dout <= 8'b11111111; //    1 : 255 - 0xff
      13'h2: dout <= 8'b11000000; //    2 : 192 - 0xc0
      13'h3: dout <= 8'b11000000; //    3 : 192 - 0xc0
      13'h4: dout <= 8'b11000000; //    4 : 192 - 0xc0
      13'h5: dout <= 8'b11000000; //    5 : 192 - 0xc0
      13'h6: dout <= 8'b11010101; //    6 : 213 - 0xd5
      13'h7: dout <= 8'b11111111; //    7 : 255 - 0xff
      13'h8: dout <= 8'b00000000; //    8 :   0 - 0x0
      13'h9: dout <= 8'b01111111; //    9 : 127 - 0x7f
      13'hA: dout <= 8'b01111111; //   10 : 127 - 0x7f
      13'hB: dout <= 8'b01111111; //   11 : 127 - 0x7f
      13'hC: dout <= 8'b01111111; //   12 : 127 - 0x7f
      13'hD: dout <= 8'b01111111; //   13 : 127 - 0x7f
      13'hE: dout <= 8'b01101010; //   14 : 106 - 0x6a
      13'hF: dout <= 8'b00000000; //   15 :   0 - 0x0
      13'h10: dout <= 8'b11111111; //   16 : 255 - 0xff -- Sprite 0x1
      13'h11: dout <= 8'b11111111; //   17 : 255 - 0xff
      13'h12: dout <= 8'b11001110; //   18 : 206 - 0xce
      13'h13: dout <= 8'b11000110; //   19 : 198 - 0xc6
      13'h14: dout <= 8'b11001110; //   20 : 206 - 0xce
      13'h15: dout <= 8'b11000110; //   21 : 198 - 0xc6
      13'h16: dout <= 8'b11101110; //   22 : 238 - 0xee
      13'h17: dout <= 8'b11111111; //   23 : 255 - 0xff
      13'h18: dout <= 8'b00000000; //   24 :   0 - 0x0
      13'h19: dout <= 8'b01111011; //   25 : 123 - 0x7b
      13'h1A: dout <= 8'b01110011; //   26 : 115 - 0x73
      13'h1B: dout <= 8'b01111011; //   27 : 123 - 0x7b
      13'h1C: dout <= 8'b01110011; //   28 : 115 - 0x73
      13'h1D: dout <= 8'b01111011; //   29 : 123 - 0x7b
      13'h1E: dout <= 8'b01010011; //   30 :  83 - 0x53
      13'h1F: dout <= 8'b00000000; //   31 :   0 - 0x0
      13'h20: dout <= 8'b11111111; //   32 : 255 - 0xff -- Sprite 0x2
      13'h21: dout <= 8'b11111111; //   33 : 255 - 0xff
      13'h22: dout <= 8'b01110001; //   34 : 113 - 0x71
      13'h23: dout <= 8'b00110011; //   35 :  51 - 0x33
      13'h24: dout <= 8'b01110001; //   36 : 113 - 0x71
      13'h25: dout <= 8'b00110011; //   37 :  51 - 0x33
      13'h26: dout <= 8'b01110101; //   38 : 117 - 0x75
      13'h27: dout <= 8'b11111111; //   39 : 255 - 0xff
      13'h28: dout <= 8'b00000000; //   40 :   0 - 0x0
      13'h29: dout <= 8'b11011110; //   41 : 222 - 0xde
      13'h2A: dout <= 8'b10011110; //   42 : 158 - 0x9e
      13'h2B: dout <= 8'b11011100; //   43 : 220 - 0xdc
      13'h2C: dout <= 8'b10011110; //   44 : 158 - 0x9e
      13'h2D: dout <= 8'b11011100; //   45 : 220 - 0xdc
      13'h2E: dout <= 8'b10011010; //   46 : 154 - 0x9a
      13'h2F: dout <= 8'b00000000; //   47 :   0 - 0x0
      13'h30: dout <= 8'b11111111; //   48 : 255 - 0xff -- Sprite 0x3
      13'h31: dout <= 8'b11111111; //   49 : 255 - 0xff
      13'h32: dout <= 8'b00000011; //   50 :   3 - 0x3
      13'h33: dout <= 8'b00000001; //   51 :   1 - 0x1
      13'h34: dout <= 8'b00000011; //   52 :   3 - 0x3
      13'h35: dout <= 8'b00000001; //   53 :   1 - 0x1
      13'h36: dout <= 8'b10101011; //   54 : 171 - 0xab
      13'h37: dout <= 8'b11111111; //   55 : 255 - 0xff
      13'h38: dout <= 8'b00000000; //   56 :   0 - 0x0
      13'h39: dout <= 8'b11111110; //   57 : 254 - 0xfe
      13'h3A: dout <= 8'b11111100; //   58 : 252 - 0xfc
      13'h3B: dout <= 8'b11111110; //   59 : 254 - 0xfe
      13'h3C: dout <= 8'b11111100; //   60 : 252 - 0xfc
      13'h3D: dout <= 8'b11111110; //   61 : 254 - 0xfe
      13'h3E: dout <= 8'b01010100; //   62 :  84 - 0x54
      13'h3F: dout <= 8'b00000000; //   63 :   0 - 0x0
      13'h40: dout <= 8'b11111111; //   64 : 255 - 0xff -- Sprite 0x4
      13'h41: dout <= 8'b11111111; //   65 : 255 - 0xff
      13'h42: dout <= 8'b11100000; //   66 : 224 - 0xe0
      13'h43: dout <= 8'b11000110; //   67 : 198 - 0xc6
      13'h44: dout <= 8'b11000110; //   68 : 198 - 0xc6
      13'h45: dout <= 8'b11110110; //   69 : 246 - 0xf6
      13'h46: dout <= 8'b11110000; //   70 : 240 - 0xf0
      13'h47: dout <= 8'b11110001; //   71 : 241 - 0xf1
      13'h48: dout <= 8'b00000000; //   72 :   0 - 0x0
      13'h49: dout <= 8'b01111111; //   73 : 127 - 0x7f
      13'h4A: dout <= 8'b01011111; //   74 :  95 - 0x5f
      13'h4B: dout <= 8'b01111001; //   75 : 121 - 0x79
      13'h4C: dout <= 8'b01111001; //   76 : 121 - 0x79
      13'h4D: dout <= 8'b01001001; //   77 :  73 - 0x49
      13'h4E: dout <= 8'b01001111; //   78 :  79 - 0x4f
      13'h4F: dout <= 8'b01001110; //   79 :  78 - 0x4e
      13'h50: dout <= 8'b11000111; //   80 : 199 - 0xc7 -- Sprite 0x5
      13'h51: dout <= 8'b11001111; //   81 : 207 - 0xcf
      13'h52: dout <= 8'b11011111; //   82 : 223 - 0xdf
      13'h53: dout <= 8'b11011111; //   83 : 223 - 0xdf
      13'h54: dout <= 8'b11001110; //   84 : 206 - 0xce
      13'h55: dout <= 8'b11100000; //   85 : 224 - 0xe0
      13'h56: dout <= 8'b11111111; //   86 : 255 - 0xff
      13'h57: dout <= 8'b11111111; //   87 : 255 - 0xff
      13'h58: dout <= 8'b01111000; //   88 : 120 - 0x78
      13'h59: dout <= 8'b01110000; //   89 : 112 - 0x70
      13'h5A: dout <= 8'b01100000; //   90 :  96 - 0x60
      13'h5B: dout <= 8'b01100000; //   91 :  96 - 0x60
      13'h5C: dout <= 8'b01110001; //   92 : 113 - 0x71
      13'h5D: dout <= 8'b01011111; //   93 :  95 - 0x5f
      13'h5E: dout <= 8'b01111111; //   94 : 127 - 0x7f
      13'h5F: dout <= 8'b00000000; //   95 :   0 - 0x0
      13'h60: dout <= 8'b11111111; //   96 : 255 - 0xff -- Sprite 0x6
      13'h61: dout <= 8'b11111111; //   97 : 255 - 0xff
      13'h62: dout <= 8'b00000111; //   98 :   7 - 0x7
      13'h63: dout <= 8'b01100011; //   99 :  99 - 0x63
      13'h64: dout <= 8'b01100011; //  100 :  99 - 0x63
      13'h65: dout <= 8'b01101111; //  101 : 111 - 0x6f
      13'h66: dout <= 8'b00001111; //  102 :  15 - 0xf
      13'h67: dout <= 8'b10001111; //  103 : 143 - 0x8f
      13'h68: dout <= 8'b00000000; //  104 :   0 - 0x0
      13'h69: dout <= 8'b11111110; //  105 : 254 - 0xfe
      13'h6A: dout <= 8'b11111010; //  106 : 250 - 0xfa
      13'h6B: dout <= 8'b10011110; //  107 : 158 - 0x9e
      13'h6C: dout <= 8'b10011110; //  108 : 158 - 0x9e
      13'h6D: dout <= 8'b10010010; //  109 : 146 - 0x92
      13'h6E: dout <= 8'b11110010; //  110 : 242 - 0xf2
      13'h6F: dout <= 8'b01110010; //  111 : 114 - 0x72
      13'h70: dout <= 8'b11100011; //  112 : 227 - 0xe3 -- Sprite 0x7
      13'h71: dout <= 8'b11110011; //  113 : 243 - 0xf3
      13'h72: dout <= 8'b11111011; //  114 : 251 - 0xfb
      13'h73: dout <= 8'b11111011; //  115 : 251 - 0xfb
      13'h74: dout <= 8'b01110011; //  116 : 115 - 0x73
      13'h75: dout <= 8'b00000111; //  117 :   7 - 0x7
      13'h76: dout <= 8'b11111111; //  118 : 255 - 0xff
      13'h77: dout <= 8'b11111111; //  119 : 255 - 0xff
      13'h78: dout <= 8'b00011110; //  120 :  30 - 0x1e
      13'h79: dout <= 8'b00001110; //  121 :  14 - 0xe
      13'h7A: dout <= 8'b00000110; //  122 :   6 - 0x6
      13'h7B: dout <= 8'b00000110; //  123 :   6 - 0x6
      13'h7C: dout <= 8'b10001110; //  124 : 142 - 0x8e
      13'h7D: dout <= 8'b11111010; //  125 : 250 - 0xfa
      13'h7E: dout <= 8'b11111110; //  126 : 254 - 0xfe
      13'h7F: dout <= 8'b00000000; //  127 :   0 - 0x0
      13'h80: dout <= 8'b11111111; //  128 : 255 - 0xff -- Sprite 0x8
      13'h81: dout <= 8'b11010101; //  129 : 213 - 0xd5
      13'h82: dout <= 8'b10101010; //  130 : 170 - 0xaa
      13'h83: dout <= 8'b11010101; //  131 : 213 - 0xd5
      13'h84: dout <= 8'b10101010; //  132 : 170 - 0xaa
      13'h85: dout <= 8'b11010101; //  133 : 213 - 0xd5
      13'h86: dout <= 8'b10101010; //  134 : 170 - 0xaa
      13'h87: dout <= 8'b11010101; //  135 : 213 - 0xd5
      13'h88: dout <= 8'b00000000; //  136 :   0 - 0x0
      13'h89: dout <= 8'b01111111; //  137 : 127 - 0x7f
      13'h8A: dout <= 8'b01011111; //  138 :  95 - 0x5f
      13'h8B: dout <= 8'b01111111; //  139 : 127 - 0x7f
      13'h8C: dout <= 8'b01111111; //  140 : 127 - 0x7f
      13'h8D: dout <= 8'b01111111; //  141 : 127 - 0x7f
      13'h8E: dout <= 8'b01111111; //  142 : 127 - 0x7f
      13'h8F: dout <= 8'b01111111; //  143 : 127 - 0x7f
      13'h90: dout <= 8'b10101010; //  144 : 170 - 0xaa -- Sprite 0x9
      13'h91: dout <= 8'b11010101; //  145 : 213 - 0xd5
      13'h92: dout <= 8'b10101010; //  146 : 170 - 0xaa
      13'h93: dout <= 8'b11010101; //  147 : 213 - 0xd5
      13'h94: dout <= 8'b10101010; //  148 : 170 - 0xaa
      13'h95: dout <= 8'b11110101; //  149 : 245 - 0xf5
      13'h96: dout <= 8'b10101010; //  150 : 170 - 0xaa
      13'h97: dout <= 8'b11111111; //  151 : 255 - 0xff
      13'h98: dout <= 8'b01111111; //  152 : 127 - 0x7f
      13'h99: dout <= 8'b01111111; //  153 : 127 - 0x7f
      13'h9A: dout <= 8'b01111111; //  154 : 127 - 0x7f
      13'h9B: dout <= 8'b01111111; //  155 : 127 - 0x7f
      13'h9C: dout <= 8'b01111111; //  156 : 127 - 0x7f
      13'h9D: dout <= 8'b01011111; //  157 :  95 - 0x5f
      13'h9E: dout <= 8'b01111111; //  158 : 127 - 0x7f
      13'h9F: dout <= 8'b00000000; //  159 :   0 - 0x0
      13'hA0: dout <= 8'b11111111; //  160 : 255 - 0xff -- Sprite 0xa
      13'hA1: dout <= 8'b01010101; //  161 :  85 - 0x55
      13'hA2: dout <= 8'b10101111; //  162 : 175 - 0xaf
      13'hA3: dout <= 8'b01010101; //  163 :  85 - 0x55
      13'hA4: dout <= 8'b10101011; //  164 : 171 - 0xab
      13'hA5: dout <= 8'b01010101; //  165 :  85 - 0x55
      13'hA6: dout <= 8'b10101011; //  166 : 171 - 0xab
      13'hA7: dout <= 8'b01010101; //  167 :  85 - 0x55
      13'hA8: dout <= 8'b00000000; //  168 :   0 - 0x0
      13'hA9: dout <= 8'b11111110; //  169 : 254 - 0xfe
      13'hAA: dout <= 8'b11111010; //  170 : 250 - 0xfa
      13'hAB: dout <= 8'b11111110; //  171 : 254 - 0xfe
      13'hAC: dout <= 8'b11111110; //  172 : 254 - 0xfe
      13'hAD: dout <= 8'b11111110; //  173 : 254 - 0xfe
      13'hAE: dout <= 8'b11111110; //  174 : 254 - 0xfe
      13'hAF: dout <= 8'b11111110; //  175 : 254 - 0xfe
      13'hB0: dout <= 8'b10101011; //  176 : 171 - 0xab -- Sprite 0xb
      13'hB1: dout <= 8'b01010101; //  177 :  85 - 0x55
      13'hB2: dout <= 8'b10101011; //  178 : 171 - 0xab
      13'hB3: dout <= 8'b01010101; //  179 :  85 - 0x55
      13'hB4: dout <= 8'b10101011; //  180 : 171 - 0xab
      13'hB5: dout <= 8'b01010101; //  181 :  85 - 0x55
      13'hB6: dout <= 8'b10101011; //  182 : 171 - 0xab
      13'hB7: dout <= 8'b11111111; //  183 : 255 - 0xff
      13'hB8: dout <= 8'b11111110; //  184 : 254 - 0xfe
      13'hB9: dout <= 8'b11111110; //  185 : 254 - 0xfe
      13'hBA: dout <= 8'b11111110; //  186 : 254 - 0xfe
      13'hBB: dout <= 8'b11111110; //  187 : 254 - 0xfe
      13'hBC: dout <= 8'b11111110; //  188 : 254 - 0xfe
      13'hBD: dout <= 8'b11111010; //  189 : 250 - 0xfa
      13'hBE: dout <= 8'b11111110; //  190 : 254 - 0xfe
      13'hBF: dout <= 8'b00000000; //  191 :   0 - 0x0
      13'hC0: dout <= 8'b11111111; //  192 : 255 - 0xff -- Sprite 0xc
      13'hC1: dout <= 8'b11010101; //  193 : 213 - 0xd5
      13'hC2: dout <= 8'b10100000; //  194 : 160 - 0xa0
      13'hC3: dout <= 8'b11010000; //  195 : 208 - 0xd0
      13'hC4: dout <= 8'b10001111; //  196 : 143 - 0x8f
      13'hC5: dout <= 8'b11001000; //  197 : 200 - 0xc8
      13'hC6: dout <= 8'b10001000; //  198 : 136 - 0x88
      13'hC7: dout <= 8'b11001000; //  199 : 200 - 0xc8
      13'hC8: dout <= 8'b00000000; //  200 :   0 - 0x0
      13'hC9: dout <= 8'b00111111; //  201 :  63 - 0x3f
      13'hCA: dout <= 8'b01011111; //  202 :  95 - 0x5f
      13'hCB: dout <= 8'b01101111; //  203 : 111 - 0x6f
      13'hCC: dout <= 8'b01110000; //  204 : 112 - 0x70
      13'hCD: dout <= 8'b01110111; //  205 : 119 - 0x77
      13'hCE: dout <= 8'b01110111; //  206 : 119 - 0x77
      13'hCF: dout <= 8'b01110111; //  207 : 119 - 0x77
      13'hD0: dout <= 8'b10001000; //  208 : 136 - 0x88 -- Sprite 0xd
      13'hD1: dout <= 8'b11001000; //  209 : 200 - 0xc8
      13'hD2: dout <= 8'b10001000; //  210 : 136 - 0x88
      13'hD3: dout <= 8'b11001111; //  211 : 207 - 0xcf
      13'hD4: dout <= 8'b10010000; //  212 : 144 - 0x90
      13'hD5: dout <= 8'b11100000; //  213 : 224 - 0xe0
      13'hD6: dout <= 8'b11101010; //  214 : 234 - 0xea
      13'hD7: dout <= 8'b11111111; //  215 : 255 - 0xff
      13'hD8: dout <= 8'b01110111; //  216 : 119 - 0x77
      13'hD9: dout <= 8'b01110111; //  217 : 119 - 0x77
      13'hDA: dout <= 8'b01110111; //  218 : 119 - 0x77
      13'hDB: dout <= 8'b01110000; //  219 : 112 - 0x70
      13'hDC: dout <= 8'b01101111; //  220 : 111 - 0x6f
      13'hDD: dout <= 8'b01011111; //  221 :  95 - 0x5f
      13'hDE: dout <= 8'b00010101; //  222 :  21 - 0x15
      13'hDF: dout <= 8'b00000000; //  223 :   0 - 0x0
      13'hE0: dout <= 8'b11111111; //  224 : 255 - 0xff -- Sprite 0xe
      13'hE1: dout <= 8'b01011011; //  225 :  91 - 0x5b
      13'hE2: dout <= 8'b00000111; //  226 :   7 - 0x7
      13'hE3: dout <= 8'b00001001; //  227 :   9 - 0x9
      13'hE4: dout <= 8'b11110011; //  228 : 243 - 0xf3
      13'hE5: dout <= 8'b00010001; //  229 :  17 - 0x11
      13'hE6: dout <= 8'b00010011; //  230 :  19 - 0x13
      13'hE7: dout <= 8'b00010001; //  231 :  17 - 0x11
      13'hE8: dout <= 8'b00000000; //  232 :   0 - 0x0
      13'hE9: dout <= 8'b11111100; //  233 : 252 - 0xfc
      13'hEA: dout <= 8'b11111000; //  234 : 248 - 0xf8
      13'hEB: dout <= 8'b11110110; //  235 : 246 - 0xf6
      13'hEC: dout <= 8'b00001100; //  236 :  12 - 0xc
      13'hED: dout <= 8'b11101110; //  237 : 238 - 0xee
      13'hEE: dout <= 8'b11101100; //  238 : 236 - 0xec
      13'hEF: dout <= 8'b11101110; //  239 : 238 - 0xee
      13'hF0: dout <= 8'b00010011; //  240 :  19 - 0x13 -- Sprite 0xf
      13'hF1: dout <= 8'b00010001; //  241 :  17 - 0x11
      13'hF2: dout <= 8'b00010011; //  242 :  19 - 0x13
      13'hF3: dout <= 8'b11110001; //  243 : 241 - 0xf1
      13'hF4: dout <= 8'b00001011; //  244 :  11 - 0xb
      13'hF5: dout <= 8'b00000101; //  245 :   5 - 0x5
      13'hF6: dout <= 8'b10101011; //  246 : 171 - 0xab
      13'hF7: dout <= 8'b11111111; //  247 : 255 - 0xff
      13'hF8: dout <= 8'b11101100; //  248 : 236 - 0xec
      13'hF9: dout <= 8'b11101110; //  249 : 238 - 0xee
      13'hFA: dout <= 8'b11101100; //  250 : 236 - 0xec
      13'hFB: dout <= 8'b00001110; //  251 :  14 - 0xe
      13'hFC: dout <= 8'b11110100; //  252 : 244 - 0xf4
      13'hFD: dout <= 8'b11111010; //  253 : 250 - 0xfa
      13'hFE: dout <= 8'b01010100; //  254 :  84 - 0x54
      13'hFF: dout <= 8'b00000000; //  255 :   0 - 0x0
      13'h100: dout <= 8'b11010000; //  256 : 208 - 0xd0 -- Sprite 0x10
      13'h101: dout <= 8'b10010000; //  257 : 144 - 0x90
      13'h102: dout <= 8'b11011111; //  258 : 223 - 0xdf
      13'h103: dout <= 8'b10011010; //  259 : 154 - 0x9a
      13'h104: dout <= 8'b11010101; //  260 : 213 - 0xd5
      13'h105: dout <= 8'b10011111; //  261 : 159 - 0x9f
      13'h106: dout <= 8'b11010000; //  262 : 208 - 0xd0
      13'h107: dout <= 8'b10010000; //  263 : 144 - 0x90
      13'h108: dout <= 8'b01100000; //  264 :  96 - 0x60
      13'h109: dout <= 8'b01100000; //  265 :  96 - 0x60
      13'h10A: dout <= 8'b01100000; //  266 :  96 - 0x60
      13'h10B: dout <= 8'b01101111; //  267 : 111 - 0x6f
      13'h10C: dout <= 8'b01101010; //  268 : 106 - 0x6a
      13'h10D: dout <= 8'b01100000; //  269 :  96 - 0x60
      13'h10E: dout <= 8'b01100000; //  270 :  96 - 0x60
      13'h10F: dout <= 8'b01100000; //  271 :  96 - 0x60
      13'h110: dout <= 8'b00001001; //  272 :   9 - 0x9 -- Sprite 0x11
      13'h111: dout <= 8'b00001011; //  273 :  11 - 0xb
      13'h112: dout <= 8'b11111001; //  274 : 249 - 0xf9
      13'h113: dout <= 8'b10101011; //  275 : 171 - 0xab
      13'h114: dout <= 8'b01011001; //  276 :  89 - 0x59
      13'h115: dout <= 8'b11111011; //  277 : 251 - 0xfb
      13'h116: dout <= 8'b00001001; //  278 :   9 - 0x9
      13'h117: dout <= 8'b00001011; //  279 :  11 - 0xb
      13'h118: dout <= 8'b00000110; //  280 :   6 - 0x6
      13'h119: dout <= 8'b00000100; //  281 :   4 - 0x4
      13'h11A: dout <= 8'b00000110; //  282 :   6 - 0x6
      13'h11B: dout <= 8'b11110100; //  283 : 244 - 0xf4
      13'h11C: dout <= 8'b10100110; //  284 : 166 - 0xa6
      13'h11D: dout <= 8'b00000100; //  285 :   4 - 0x4
      13'h11E: dout <= 8'b00000110; //  286 :   6 - 0x6
      13'h11F: dout <= 8'b00000100; //  287 :   4 - 0x4
      13'h120: dout <= 8'b00011000; //  288 :  24 - 0x18 -- Sprite 0x12
      13'h121: dout <= 8'b00010100; //  289 :  20 - 0x14
      13'h122: dout <= 8'b00010100; //  290 :  20 - 0x14
      13'h123: dout <= 8'b00111010; //  291 :  58 - 0x3a
      13'h124: dout <= 8'b00111010; //  292 :  58 - 0x3a
      13'h125: dout <= 8'b01111010; //  293 : 122 - 0x7a
      13'h126: dout <= 8'b01111010; //  294 : 122 - 0x7a
      13'h127: dout <= 8'b01111010; //  295 : 122 - 0x7a
      13'h128: dout <= 8'b00000000; //  296 :   0 - 0x0
      13'h129: dout <= 8'b00001000; //  297 :   8 - 0x8
      13'h12A: dout <= 8'b00001000; //  298 :   8 - 0x8
      13'h12B: dout <= 8'b00011100; //  299 :  28 - 0x1c
      13'h12C: dout <= 8'b00011100; //  300 :  28 - 0x1c
      13'h12D: dout <= 8'b00111100; //  301 :  60 - 0x3c
      13'h12E: dout <= 8'b00111100; //  302 :  60 - 0x3c
      13'h12F: dout <= 8'b00111100; //  303 :  60 - 0x3c
      13'h130: dout <= 8'b11111011; //  304 : 251 - 0xfb -- Sprite 0x13
      13'h131: dout <= 8'b11111101; //  305 : 253 - 0xfd
      13'h132: dout <= 8'b11111101; //  306 : 253 - 0xfd
      13'h133: dout <= 8'b11111101; //  307 : 253 - 0xfd
      13'h134: dout <= 8'b11111101; //  308 : 253 - 0xfd
      13'h135: dout <= 8'b11111101; //  309 : 253 - 0xfd
      13'h136: dout <= 8'b10000001; //  310 : 129 - 0x81
      13'h137: dout <= 8'b11111111; //  311 : 255 - 0xff
      13'h138: dout <= 8'b00111100; //  312 :  60 - 0x3c
      13'h139: dout <= 8'b01111110; //  313 : 126 - 0x7e
      13'h13A: dout <= 8'b01111110; //  314 : 126 - 0x7e
      13'h13B: dout <= 8'b01111110; //  315 : 126 - 0x7e
      13'h13C: dout <= 8'b01111110; //  316 : 126 - 0x7e
      13'h13D: dout <= 8'b01111110; //  317 : 126 - 0x7e
      13'h13E: dout <= 8'b01111110; //  318 : 126 - 0x7e
      13'h13F: dout <= 8'b00000000; //  319 :   0 - 0x0
      13'h140: dout <= 8'b00000000; //  320 :   0 - 0x0 -- Sprite 0x14
      13'h141: dout <= 8'b00000111; //  321 :   7 - 0x7
      13'h142: dout <= 8'b00000010; //  322 :   2 - 0x2
      13'h143: dout <= 8'b00000100; //  323 :   4 - 0x4
      13'h144: dout <= 8'b00000011; //  324 :   3 - 0x3
      13'h145: dout <= 8'b00000011; //  325 :   3 - 0x3
      13'h146: dout <= 8'b00001101; //  326 :  13 - 0xd
      13'h147: dout <= 8'b00010111; //  327 :  23 - 0x17
      13'h148: dout <= 8'b00000000; //  328 :   0 - 0x0
      13'h149: dout <= 8'b00000000; //  329 :   0 - 0x0
      13'h14A: dout <= 8'b00000101; //  330 :   5 - 0x5
      13'h14B: dout <= 8'b00000011; //  331 :   3 - 0x3
      13'h14C: dout <= 8'b00000000; //  332 :   0 - 0x0
      13'h14D: dout <= 8'b00000000; //  333 :   0 - 0x0
      13'h14E: dout <= 8'b00000010; //  334 :   2 - 0x2
      13'h14F: dout <= 8'b00001111; //  335 :  15 - 0xf
      13'h150: dout <= 8'b00101111; //  336 :  47 - 0x2f -- Sprite 0x15
      13'h151: dout <= 8'b01001111; //  337 :  79 - 0x4f
      13'h152: dout <= 8'b01001111; //  338 :  79 - 0x4f
      13'h153: dout <= 8'b01001111; //  339 :  79 - 0x4f
      13'h154: dout <= 8'b01001111; //  340 :  79 - 0x4f
      13'h155: dout <= 8'b00100111; //  341 :  39 - 0x27
      13'h156: dout <= 8'b00010000; //  342 :  16 - 0x10
      13'h157: dout <= 8'b00001111; //  343 :  15 - 0xf
      13'h158: dout <= 8'b00011100; //  344 :  28 - 0x1c
      13'h159: dout <= 8'b00111010; //  345 :  58 - 0x3a
      13'h15A: dout <= 8'b00111100; //  346 :  60 - 0x3c
      13'h15B: dout <= 8'b00111111; //  347 :  63 - 0x3f
      13'h15C: dout <= 8'b00111000; //  348 :  56 - 0x38
      13'h15D: dout <= 8'b00011110; //  349 :  30 - 0x1e
      13'h15E: dout <= 8'b00001111; //  350 :  15 - 0xf
      13'h15F: dout <= 8'b00000000; //  351 :   0 - 0x0
      13'h160: dout <= 8'b00000000; //  352 :   0 - 0x0 -- Sprite 0x16
      13'h161: dout <= 8'b11100000; //  353 : 224 - 0xe0
      13'h162: dout <= 8'b10100000; //  354 : 160 - 0xa0
      13'h163: dout <= 8'b00100000; //  355 :  32 - 0x20
      13'h164: dout <= 8'b11000000; //  356 : 192 - 0xc0
      13'h165: dout <= 8'b01000000; //  357 :  64 - 0x40
      13'h166: dout <= 8'b00110000; //  358 :  48 - 0x30
      13'h167: dout <= 8'b11101000; //  359 : 232 - 0xe8
      13'h168: dout <= 8'b00000000; //  360 :   0 - 0x0
      13'h169: dout <= 8'b00000000; //  361 :   0 - 0x0
      13'h16A: dout <= 8'b01000000; //  362 :  64 - 0x40
      13'h16B: dout <= 8'b11000000; //  363 : 192 - 0xc0
      13'h16C: dout <= 8'b00000000; //  364 :   0 - 0x0
      13'h16D: dout <= 8'b10000000; //  365 : 128 - 0x80
      13'h16E: dout <= 8'b11000000; //  366 : 192 - 0xc0
      13'h16F: dout <= 8'b01110000; //  367 : 112 - 0x70
      13'h170: dout <= 8'b11110100; //  368 : 244 - 0xf4 -- Sprite 0x17
      13'h171: dout <= 8'b11110010; //  369 : 242 - 0xf2
      13'h172: dout <= 8'b11110010; //  370 : 242 - 0xf2
      13'h173: dout <= 8'b11110010; //  371 : 242 - 0xf2
      13'h174: dout <= 8'b11110010; //  372 : 242 - 0xf2
      13'h175: dout <= 8'b11100100; //  373 : 228 - 0xe4
      13'h176: dout <= 8'b00001000; //  374 :   8 - 0x8
      13'h177: dout <= 8'b11110000; //  375 : 240 - 0xf0
      13'h178: dout <= 8'b00011000; //  376 :  24 - 0x18
      13'h179: dout <= 8'b11111100; //  377 : 252 - 0xfc
      13'h17A: dout <= 8'b00111100; //  378 :  60 - 0x3c
      13'h17B: dout <= 8'b01011100; //  379 :  92 - 0x5c
      13'h17C: dout <= 8'b00111100; //  380 :  60 - 0x3c
      13'h17D: dout <= 8'b11111000; //  381 : 248 - 0xf8
      13'h17E: dout <= 8'b11110000; //  382 : 240 - 0xf0
      13'h17F: dout <= 8'b00000000; //  383 :   0 - 0x0
      13'h180: dout <= 8'b00111111; //  384 :  63 - 0x3f -- Sprite 0x18
      13'h181: dout <= 8'b01000000; //  385 :  64 - 0x40
      13'h182: dout <= 8'b01000000; //  386 :  64 - 0x40
      13'h183: dout <= 8'b10000000; //  387 : 128 - 0x80
      13'h184: dout <= 8'b10000000; //  388 : 128 - 0x80
      13'h185: dout <= 8'b01111111; //  389 : 127 - 0x7f
      13'h186: dout <= 8'b00000001; //  390 :   1 - 0x1
      13'h187: dout <= 8'b01111111; //  391 : 127 - 0x7f
      13'h188: dout <= 8'b00000000; //  392 :   0 - 0x0
      13'h189: dout <= 8'b00111111; //  393 :  63 - 0x3f
      13'h18A: dout <= 8'b00111111; //  394 :  63 - 0x3f
      13'h18B: dout <= 8'b01111111; //  395 : 127 - 0x7f
      13'h18C: dout <= 8'b01111111; //  396 : 127 - 0x7f
      13'h18D: dout <= 8'b00000000; //  397 :   0 - 0x0
      13'h18E: dout <= 8'b00000000; //  398 :   0 - 0x0
      13'h18F: dout <= 8'b00000000; //  399 :   0 - 0x0
      13'h190: dout <= 8'b11111100; //  400 : 252 - 0xfc -- Sprite 0x19
      13'h191: dout <= 8'b00000010; //  401 :   2 - 0x2
      13'h192: dout <= 8'b00000010; //  402 :   2 - 0x2
      13'h193: dout <= 8'b00000001; //  403 :   1 - 0x1
      13'h194: dout <= 8'b00000001; //  404 :   1 - 0x1
      13'h195: dout <= 8'b11111110; //  405 : 254 - 0xfe
      13'h196: dout <= 8'b10000000; //  406 : 128 - 0x80
      13'h197: dout <= 8'b11111110; //  407 : 254 - 0xfe
      13'h198: dout <= 8'b00000000; //  408 :   0 - 0x0
      13'h199: dout <= 8'b11111100; //  409 : 252 - 0xfc
      13'h19A: dout <= 8'b11111100; //  410 : 252 - 0xfc
      13'h19B: dout <= 8'b11111110; //  411 : 254 - 0xfe
      13'h19C: dout <= 8'b11111110; //  412 : 254 - 0xfe
      13'h19D: dout <= 8'b00000000; //  413 :   0 - 0x0
      13'h19E: dout <= 8'b00000000; //  414 :   0 - 0x0
      13'h19F: dout <= 8'b00000000; //  415 :   0 - 0x0
      13'h1A0: dout <= 8'b00000000; //  416 :   0 - 0x0 -- Sprite 0x1a
      13'h1A1: dout <= 8'b00000000; //  417 :   0 - 0x0
      13'h1A2: dout <= 8'b00111111; //  418 :  63 - 0x3f
      13'h1A3: dout <= 8'b01000000; //  419 :  64 - 0x40
      13'h1A4: dout <= 8'b01000000; //  420 :  64 - 0x40
      13'h1A5: dout <= 8'b10000000; //  421 : 128 - 0x80
      13'h1A6: dout <= 8'b10000000; //  422 : 128 - 0x80
      13'h1A7: dout <= 8'b01111111; //  423 : 127 - 0x7f
      13'h1A8: dout <= 8'b00000000; //  424 :   0 - 0x0
      13'h1A9: dout <= 8'b00000000; //  425 :   0 - 0x0
      13'h1AA: dout <= 8'b00000000; //  426 :   0 - 0x0
      13'h1AB: dout <= 8'b00111111; //  427 :  63 - 0x3f
      13'h1AC: dout <= 8'b00111111; //  428 :  63 - 0x3f
      13'h1AD: dout <= 8'b01111111; //  429 : 127 - 0x7f
      13'h1AE: dout <= 8'b01111111; //  430 : 127 - 0x7f
      13'h1AF: dout <= 8'b00000000; //  431 :   0 - 0x0
      13'h1B0: dout <= 8'b00000000; //  432 :   0 - 0x0 -- Sprite 0x1b
      13'h1B1: dout <= 8'b00000000; //  433 :   0 - 0x0
      13'h1B2: dout <= 8'b11111100; //  434 : 252 - 0xfc
      13'h1B3: dout <= 8'b00000010; //  435 :   2 - 0x2
      13'h1B4: dout <= 8'b00000010; //  436 :   2 - 0x2
      13'h1B5: dout <= 8'b00000001; //  437 :   1 - 0x1
      13'h1B6: dout <= 8'b00000001; //  438 :   1 - 0x1
      13'h1B7: dout <= 8'b11111110; //  439 : 254 - 0xfe
      13'h1B8: dout <= 8'b00000000; //  440 :   0 - 0x0
      13'h1B9: dout <= 8'b00000000; //  441 :   0 - 0x0
      13'h1BA: dout <= 8'b00000000; //  442 :   0 - 0x0
      13'h1BB: dout <= 8'b11111100; //  443 : 252 - 0xfc
      13'h1BC: dout <= 8'b11111100; //  444 : 252 - 0xfc
      13'h1BD: dout <= 8'b11111110; //  445 : 254 - 0xfe
      13'h1BE: dout <= 8'b11111110; //  446 : 254 - 0xfe
      13'h1BF: dout <= 8'b00000000; //  447 :   0 - 0x0
      13'h1C0: dout <= 8'b01111111; //  448 : 127 - 0x7f -- Sprite 0x1c
      13'h1C1: dout <= 8'b10000000; //  449 : 128 - 0x80
      13'h1C2: dout <= 8'b10000000; //  450 : 128 - 0x80
      13'h1C3: dout <= 8'b10000000; //  451 : 128 - 0x80
      13'h1C4: dout <= 8'b10011011; //  452 : 155 - 0x9b
      13'h1C5: dout <= 8'b10100100; //  453 : 164 - 0xa4
      13'h1C6: dout <= 8'b10100110; //  454 : 166 - 0xa6
      13'h1C7: dout <= 8'b10000000; //  455 : 128 - 0x80
      13'h1C8: dout <= 8'b00000000; //  456 :   0 - 0x0
      13'h1C9: dout <= 8'b01111111; //  457 : 127 - 0x7f
      13'h1CA: dout <= 8'b01111111; //  458 : 127 - 0x7f
      13'h1CB: dout <= 8'b01111111; //  459 : 127 - 0x7f
      13'h1CC: dout <= 8'b01100100; //  460 : 100 - 0x64
      13'h1CD: dout <= 8'b01011011; //  461 :  91 - 0x5b
      13'h1CE: dout <= 8'b01011001; //  462 :  89 - 0x59
      13'h1CF: dout <= 8'b01111111; //  463 : 127 - 0x7f
      13'h1D0: dout <= 8'b10000000; //  464 : 128 - 0x80 -- Sprite 0x1d
      13'h1D1: dout <= 8'b01111111; //  465 : 127 - 0x7f
      13'h1D2: dout <= 8'b00000010; //  466 :   2 - 0x2
      13'h1D3: dout <= 8'b00000010; //  467 :   2 - 0x2
      13'h1D4: dout <= 8'b00000010; //  468 :   2 - 0x2
      13'h1D5: dout <= 8'b00000010; //  469 :   2 - 0x2
      13'h1D6: dout <= 8'b00000010; //  470 :   2 - 0x2
      13'h1D7: dout <= 8'b00001111; //  471 :  15 - 0xf
      13'h1D8: dout <= 8'b01111111; //  472 : 127 - 0x7f
      13'h1D9: dout <= 8'b00000000; //  473 :   0 - 0x0
      13'h1DA: dout <= 8'b00000001; //  474 :   1 - 0x1
      13'h1DB: dout <= 8'b00000001; //  475 :   1 - 0x1
      13'h1DC: dout <= 8'b00000001; //  476 :   1 - 0x1
      13'h1DD: dout <= 8'b00000001; //  477 :   1 - 0x1
      13'h1DE: dout <= 8'b00000001; //  478 :   1 - 0x1
      13'h1DF: dout <= 8'b00000000; //  479 :   0 - 0x0
      13'h1E0: dout <= 8'b11111110; //  480 : 254 - 0xfe -- Sprite 0x1e
      13'h1E1: dout <= 8'b00000001; //  481 :   1 - 0x1
      13'h1E2: dout <= 8'b00000001; //  482 :   1 - 0x1
      13'h1E3: dout <= 8'b00000001; //  483 :   1 - 0x1
      13'h1E4: dout <= 8'b01000001; //  484 :  65 - 0x41
      13'h1E5: dout <= 8'b11110101; //  485 : 245 - 0xf5
      13'h1E6: dout <= 8'b00011101; //  486 :  29 - 0x1d
      13'h1E7: dout <= 8'b00000001; //  487 :   1 - 0x1
      13'h1E8: dout <= 8'b00000000; //  488 :   0 - 0x0
      13'h1E9: dout <= 8'b11111110; //  489 : 254 - 0xfe
      13'h1EA: dout <= 8'b11111110; //  490 : 254 - 0xfe
      13'h1EB: dout <= 8'b11111110; //  491 : 254 - 0xfe
      13'h1EC: dout <= 8'b10111110; //  492 : 190 - 0xbe
      13'h1ED: dout <= 8'b00001010; //  493 :  10 - 0xa
      13'h1EE: dout <= 8'b11100010; //  494 : 226 - 0xe2
      13'h1EF: dout <= 8'b11111110; //  495 : 254 - 0xfe
      13'h1F0: dout <= 8'b00000001; //  496 :   1 - 0x1 -- Sprite 0x1f
      13'h1F1: dout <= 8'b11111110; //  497 : 254 - 0xfe
      13'h1F2: dout <= 8'b01000000; //  498 :  64 - 0x40
      13'h1F3: dout <= 8'b01000000; //  499 :  64 - 0x40
      13'h1F4: dout <= 8'b01000000; //  500 :  64 - 0x40
      13'h1F5: dout <= 8'b01000000; //  501 :  64 - 0x40
      13'h1F6: dout <= 8'b01000000; //  502 :  64 - 0x40
      13'h1F7: dout <= 8'b11110000; //  503 : 240 - 0xf0
      13'h1F8: dout <= 8'b11111110; //  504 : 254 - 0xfe
      13'h1F9: dout <= 8'b00000000; //  505 :   0 - 0x0
      13'h1FA: dout <= 8'b10000000; //  506 : 128 - 0x80
      13'h1FB: dout <= 8'b10000000; //  507 : 128 - 0x80
      13'h1FC: dout <= 8'b10000000; //  508 : 128 - 0x80
      13'h1FD: dout <= 8'b10000000; //  509 : 128 - 0x80
      13'h1FE: dout <= 8'b10000000; //  510 : 128 - 0x80
      13'h1FF: dout <= 8'b00000000; //  511 :   0 - 0x0
      13'h200: dout <= 8'b00000111; //  512 :   7 - 0x7 -- Sprite 0x20
      13'h201: dout <= 8'b00011111; //  513 :  31 - 0x1f
      13'h202: dout <= 8'b00111111; //  514 :  63 - 0x3f
      13'h203: dout <= 8'b01111111; //  515 : 127 - 0x7f
      13'h204: dout <= 8'b01111111; //  516 : 127 - 0x7f
      13'h205: dout <= 8'b11111111; //  517 : 255 - 0xff
      13'h206: dout <= 8'b11111111; //  518 : 255 - 0xff
      13'h207: dout <= 8'b11111111; //  519 : 255 - 0xff
      13'h208: dout <= 8'b00000000; //  520 :   0 - 0x0
      13'h209: dout <= 8'b00000000; //  521 :   0 - 0x0
      13'h20A: dout <= 8'b00000000; //  522 :   0 - 0x0
      13'h20B: dout <= 8'b00000000; //  523 :   0 - 0x0
      13'h20C: dout <= 8'b00000000; //  524 :   0 - 0x0
      13'h20D: dout <= 8'b00000000; //  525 :   0 - 0x0
      13'h20E: dout <= 8'b00000000; //  526 :   0 - 0x0
      13'h20F: dout <= 8'b00000000; //  527 :   0 - 0x0
      13'h210: dout <= 8'b11100000; //  528 : 224 - 0xe0 -- Sprite 0x21
      13'h211: dout <= 8'b11111000; //  529 : 248 - 0xf8
      13'h212: dout <= 8'b11111100; //  530 : 252 - 0xfc
      13'h213: dout <= 8'b11111110; //  531 : 254 - 0xfe
      13'h214: dout <= 8'b11111110; //  532 : 254 - 0xfe
      13'h215: dout <= 8'b11111111; //  533 : 255 - 0xff
      13'h216: dout <= 8'b11111111; //  534 : 255 - 0xff
      13'h217: dout <= 8'b11111111; //  535 : 255 - 0xff
      13'h218: dout <= 8'b00000000; //  536 :   0 - 0x0
      13'h219: dout <= 8'b00000000; //  537 :   0 - 0x0
      13'h21A: dout <= 8'b00000000; //  538 :   0 - 0x0
      13'h21B: dout <= 8'b00000000; //  539 :   0 - 0x0
      13'h21C: dout <= 8'b00000000; //  540 :   0 - 0x0
      13'h21D: dout <= 8'b00000000; //  541 :   0 - 0x0
      13'h21E: dout <= 8'b00000000; //  542 :   0 - 0x0
      13'h21F: dout <= 8'b00000000; //  543 :   0 - 0x0
      13'h220: dout <= 8'b00000111; //  544 :   7 - 0x7 -- Sprite 0x22
      13'h221: dout <= 8'b00011111; //  545 :  31 - 0x1f
      13'h222: dout <= 8'b00111111; //  546 :  63 - 0x3f
      13'h223: dout <= 8'b01111111; //  547 : 127 - 0x7f
      13'h224: dout <= 8'b01111111; //  548 : 127 - 0x7f
      13'h225: dout <= 8'b11111111; //  549 : 255 - 0xff
      13'h226: dout <= 8'b11111111; //  550 : 255 - 0xff
      13'h227: dout <= 8'b11111111; //  551 : 255 - 0xff
      13'h228: dout <= 8'b00000000; //  552 :   0 - 0x0
      13'h229: dout <= 8'b00000000; //  553 :   0 - 0x0
      13'h22A: dout <= 8'b00011000; //  554 :  24 - 0x18
      13'h22B: dout <= 8'b00010000; //  555 :  16 - 0x10
      13'h22C: dout <= 8'b00011010; //  556 :  26 - 0x1a
      13'h22D: dout <= 8'b00010001; //  557 :  17 - 0x11
      13'h22E: dout <= 8'b00011010; //  558 :  26 - 0x1a
      13'h22F: dout <= 8'b00000000; //  559 :   0 - 0x0
      13'h230: dout <= 8'b11100000; //  560 : 224 - 0xe0 -- Sprite 0x23
      13'h231: dout <= 8'b11111000; //  561 : 248 - 0xf8
      13'h232: dout <= 8'b11111100; //  562 : 252 - 0xfc
      13'h233: dout <= 8'b11111110; //  563 : 254 - 0xfe
      13'h234: dout <= 8'b11111110; //  564 : 254 - 0xfe
      13'h235: dout <= 8'b11111111; //  565 : 255 - 0xff
      13'h236: dout <= 8'b11111111; //  566 : 255 - 0xff
      13'h237: dout <= 8'b11111111; //  567 : 255 - 0xff
      13'h238: dout <= 8'b00000000; //  568 :   0 - 0x0
      13'h239: dout <= 8'b00000000; //  569 :   0 - 0x0
      13'h23A: dout <= 8'b00000000; //  570 :   0 - 0x0
      13'h23B: dout <= 8'b00101000; //  571 :  40 - 0x28
      13'h23C: dout <= 8'b10001100; //  572 : 140 - 0x8c
      13'h23D: dout <= 8'b00101000; //  573 :  40 - 0x28
      13'h23E: dout <= 8'b10101100; //  574 : 172 - 0xac
      13'h23F: dout <= 8'b00000000; //  575 :   0 - 0x0
      13'h240: dout <= 8'b00000000; //  576 :   0 - 0x0 -- Sprite 0x24
      13'h241: dout <= 8'b00000000; //  577 :   0 - 0x0
      13'h242: dout <= 8'b00000000; //  578 :   0 - 0x0
      13'h243: dout <= 8'b00000000; //  579 :   0 - 0x0
      13'h244: dout <= 8'b00000000; //  580 :   0 - 0x0
      13'h245: dout <= 8'b00000000; //  581 :   0 - 0x0
      13'h246: dout <= 8'b00000000; //  582 :   0 - 0x0
      13'h247: dout <= 8'b00000000; //  583 :   0 - 0x0
      13'h248: dout <= 8'b00000000; //  584 :   0 - 0x0
      13'h249: dout <= 8'b00000000; //  585 :   0 - 0x0
      13'h24A: dout <= 8'b00000000; //  586 :   0 - 0x0
      13'h24B: dout <= 8'b00000000; //  587 :   0 - 0x0
      13'h24C: dout <= 8'b00000000; //  588 :   0 - 0x0
      13'h24D: dout <= 8'b00000000; //  589 :   0 - 0x0
      13'h24E: dout <= 8'b00000000; //  590 :   0 - 0x0
      13'h24F: dout <= 8'b00000000; //  591 :   0 - 0x0
      13'h250: dout <= 8'b00101111; //  592 :  47 - 0x2f -- Sprite 0x25
      13'h251: dout <= 8'b01001111; //  593 :  79 - 0x4f
      13'h252: dout <= 8'b01001111; //  594 :  79 - 0x4f
      13'h253: dout <= 8'b01001111; //  595 :  79 - 0x4f
      13'h254: dout <= 8'b01001111; //  596 :  79 - 0x4f
      13'h255: dout <= 8'b00100111; //  597 :  39 - 0x27
      13'h256: dout <= 8'b00010000; //  598 :  16 - 0x10
      13'h257: dout <= 8'b00001111; //  599 :  15 - 0xf
      13'h258: dout <= 8'b00011100; //  600 :  28 - 0x1c
      13'h259: dout <= 8'b00111001; //  601 :  57 - 0x39
      13'h25A: dout <= 8'b00111111; //  602 :  63 - 0x3f
      13'h25B: dout <= 8'b00111110; //  603 :  62 - 0x3e
      13'h25C: dout <= 8'b00111111; //  604 :  63 - 0x3f
      13'h25D: dout <= 8'b00011110; //  605 :  30 - 0x1e
      13'h25E: dout <= 8'b00001111; //  606 :  15 - 0xf
      13'h25F: dout <= 8'b00000000; //  607 :   0 - 0x0
      13'h260: dout <= 8'b00000000; //  608 :   0 - 0x0 -- Sprite 0x26
      13'h261: dout <= 8'b11100000; //  609 : 224 - 0xe0
      13'h262: dout <= 8'b10100000; //  610 : 160 - 0xa0
      13'h263: dout <= 8'b00100000; //  611 :  32 - 0x20
      13'h264: dout <= 8'b11000000; //  612 : 192 - 0xc0
      13'h265: dout <= 8'b01000000; //  613 :  64 - 0x40
      13'h266: dout <= 8'b00110000; //  614 :  48 - 0x30
      13'h267: dout <= 8'b11101000; //  615 : 232 - 0xe8
      13'h268: dout <= 8'b00000000; //  616 :   0 - 0x0
      13'h269: dout <= 8'b00000000; //  617 :   0 - 0x0
      13'h26A: dout <= 8'b01000000; //  618 :  64 - 0x40
      13'h26B: dout <= 8'b11000000; //  619 : 192 - 0xc0
      13'h26C: dout <= 8'b00000000; //  620 :   0 - 0x0
      13'h26D: dout <= 8'b10000000; //  621 : 128 - 0x80
      13'h26E: dout <= 8'b11000000; //  622 : 192 - 0xc0
      13'h26F: dout <= 8'b11110000; //  623 : 240 - 0xf0
      13'h270: dout <= 8'b11110100; //  624 : 244 - 0xf4 -- Sprite 0x27
      13'h271: dout <= 8'b11110010; //  625 : 242 - 0xf2
      13'h272: dout <= 8'b11110010; //  626 : 242 - 0xf2
      13'h273: dout <= 8'b11110010; //  627 : 242 - 0xf2
      13'h274: dout <= 8'b11110010; //  628 : 242 - 0xf2
      13'h275: dout <= 8'b11100100; //  629 : 228 - 0xe4
      13'h276: dout <= 8'b00001000; //  630 :   8 - 0x8
      13'h277: dout <= 8'b11110000; //  631 : 240 - 0xf0
      13'h278: dout <= 8'b00111000; //  632 :  56 - 0x38
      13'h279: dout <= 8'b10011100; //  633 : 156 - 0x9c
      13'h27A: dout <= 8'b10011100; //  634 : 156 - 0x9c
      13'h27B: dout <= 8'b00111100; //  635 :  60 - 0x3c
      13'h27C: dout <= 8'b11111100; //  636 : 252 - 0xfc
      13'h27D: dout <= 8'b01111000; //  637 : 120 - 0x78
      13'h27E: dout <= 8'b11110000; //  638 : 240 - 0xf0
      13'h27F: dout <= 8'b00000000; //  639 :   0 - 0x0
      13'h280: dout <= 8'b11111111; //  640 : 255 - 0xff -- Sprite 0x28
      13'h281: dout <= 8'b11010101; //  641 : 213 - 0xd5
      13'h282: dout <= 8'b10100011; //  642 : 163 - 0xa3
      13'h283: dout <= 8'b11010111; //  643 : 215 - 0xd7
      13'h284: dout <= 8'b10001111; //  644 : 143 - 0x8f
      13'h285: dout <= 8'b11001111; //  645 : 207 - 0xcf
      13'h286: dout <= 8'b10001011; //  646 : 139 - 0x8b
      13'h287: dout <= 8'b11001011; //  647 : 203 - 0xcb
      13'h288: dout <= 8'b00000000; //  648 :   0 - 0x0
      13'h289: dout <= 8'b00111110; //  649 :  62 - 0x3e
      13'h28A: dout <= 8'b01011101; //  650 :  93 - 0x5d
      13'h28B: dout <= 8'b01101011; //  651 : 107 - 0x6b
      13'h28C: dout <= 8'b01110101; //  652 : 117 - 0x75
      13'h28D: dout <= 8'b01110001; //  653 : 113 - 0x71
      13'h28E: dout <= 8'b01110101; //  654 : 117 - 0x75
      13'h28F: dout <= 8'b01110100; //  655 : 116 - 0x74
      13'h290: dout <= 8'b10001111; //  656 : 143 - 0x8f -- Sprite 0x29
      13'h291: dout <= 8'b11001111; //  657 : 207 - 0xcf
      13'h292: dout <= 8'b10001111; //  658 : 143 - 0x8f
      13'h293: dout <= 8'b11001111; //  659 : 207 - 0xcf
      13'h294: dout <= 8'b10010000; //  660 : 144 - 0x90
      13'h295: dout <= 8'b11100000; //  661 : 224 - 0xe0
      13'h296: dout <= 8'b11101010; //  662 : 234 - 0xea
      13'h297: dout <= 8'b11111111; //  663 : 255 - 0xff
      13'h298: dout <= 8'b01110000; //  664 : 112 - 0x70
      13'h299: dout <= 8'b01110111; //  665 : 119 - 0x77
      13'h29A: dout <= 8'b01110111; //  666 : 119 - 0x77
      13'h29B: dout <= 8'b01110000; //  667 : 112 - 0x70
      13'h29C: dout <= 8'b01101111; //  668 : 111 - 0x6f
      13'h29D: dout <= 8'b01011111; //  669 :  95 - 0x5f
      13'h29E: dout <= 8'b00010101; //  670 :  21 - 0x15
      13'h29F: dout <= 8'b00000000; //  671 :   0 - 0x0
      13'h2A0: dout <= 8'b11111111; //  672 : 255 - 0xff -- Sprite 0x2a
      13'h2A1: dout <= 8'b11011011; //  673 : 219 - 0xdb
      13'h2A2: dout <= 8'b11000111; //  674 : 199 - 0xc7
      13'h2A3: dout <= 8'b11101001; //  675 : 233 - 0xe9
      13'h2A4: dout <= 8'b11110011; //  676 : 243 - 0xf3
      13'h2A5: dout <= 8'b11110001; //  677 : 241 - 0xf1
      13'h2A6: dout <= 8'b11010011; //  678 : 211 - 0xd3
      13'h2A7: dout <= 8'b11010001; //  679 : 209 - 0xd1
      13'h2A8: dout <= 8'b00000000; //  680 :   0 - 0x0
      13'h2A9: dout <= 8'b01111100; //  681 : 124 - 0x7c
      13'h2AA: dout <= 8'b10111000; //  682 : 184 - 0xb8
      13'h2AB: dout <= 8'b11010110; //  683 : 214 - 0xd6
      13'h2AC: dout <= 8'b10101100; //  684 : 172 - 0xac
      13'h2AD: dout <= 8'b10001110; //  685 : 142 - 0x8e
      13'h2AE: dout <= 8'b10101100; //  686 : 172 - 0xac
      13'h2AF: dout <= 8'b00101110; //  687 :  46 - 0x2e
      13'h2B0: dout <= 8'b11110011; //  688 : 243 - 0xf3 -- Sprite 0x2b
      13'h2B1: dout <= 8'b11110001; //  689 : 241 - 0xf1
      13'h2B2: dout <= 8'b11110011; //  690 : 243 - 0xf3
      13'h2B3: dout <= 8'b11110001; //  691 : 241 - 0xf1
      13'h2B4: dout <= 8'b00001011; //  692 :  11 - 0xb
      13'h2B5: dout <= 8'b00000101; //  693 :   5 - 0x5
      13'h2B6: dout <= 8'b10101011; //  694 : 171 - 0xab
      13'h2B7: dout <= 8'b11111111; //  695 : 255 - 0xff
      13'h2B8: dout <= 8'b00001100; //  696 :  12 - 0xc
      13'h2B9: dout <= 8'b11101110; //  697 : 238 - 0xee
      13'h2BA: dout <= 8'b11101100; //  698 : 236 - 0xec
      13'h2BB: dout <= 8'b00001110; //  699 :  14 - 0xe
      13'h2BC: dout <= 8'b11110100; //  700 : 244 - 0xf4
      13'h2BD: dout <= 8'b11111010; //  701 : 250 - 0xfa
      13'h2BE: dout <= 8'b01010100; //  702 :  84 - 0x54
      13'h2BF: dout <= 8'b00000000; //  703 :   0 - 0x0
      13'h2C0: dout <= 8'b00000000; //  704 :   0 - 0x0 -- Sprite 0x2c
      13'h2C1: dout <= 8'b00000000; //  705 :   0 - 0x0
      13'h2C2: dout <= 8'b00000000; //  706 :   0 - 0x0
      13'h2C3: dout <= 8'b00000000; //  707 :   0 - 0x0
      13'h2C4: dout <= 8'b00000000; //  708 :   0 - 0x0
      13'h2C5: dout <= 8'b00000000; //  709 :   0 - 0x0
      13'h2C6: dout <= 8'b00000000; //  710 :   0 - 0x0
      13'h2C7: dout <= 8'b00000000; //  711 :   0 - 0x0
      13'h2C8: dout <= 8'b00000000; //  712 :   0 - 0x0
      13'h2C9: dout <= 8'b00000000; //  713 :   0 - 0x0
      13'h2CA: dout <= 8'b00000000; //  714 :   0 - 0x0
      13'h2CB: dout <= 8'b00000000; //  715 :   0 - 0x0
      13'h2CC: dout <= 8'b00000000; //  716 :   0 - 0x0
      13'h2CD: dout <= 8'b00000000; //  717 :   0 - 0x0
      13'h2CE: dout <= 8'b00000000; //  718 :   0 - 0x0
      13'h2CF: dout <= 8'b00000000; //  719 :   0 - 0x0
      13'h2D0: dout <= 8'b00101111; //  720 :  47 - 0x2f -- Sprite 0x2d
      13'h2D1: dout <= 8'b01001111; //  721 :  79 - 0x4f
      13'h2D2: dout <= 8'b01001111; //  722 :  79 - 0x4f
      13'h2D3: dout <= 8'b01001111; //  723 :  79 - 0x4f
      13'h2D4: dout <= 8'b01001111; //  724 :  79 - 0x4f
      13'h2D5: dout <= 8'b00100111; //  725 :  39 - 0x27
      13'h2D6: dout <= 8'b00010000; //  726 :  16 - 0x10
      13'h2D7: dout <= 8'b00001111; //  727 :  15 - 0xf
      13'h2D8: dout <= 8'b00011110; //  728 :  30 - 0x1e
      13'h2D9: dout <= 8'b00111110; //  729 :  62 - 0x3e
      13'h2DA: dout <= 8'b00111110; //  730 :  62 - 0x3e
      13'h2DB: dout <= 8'b00111110; //  731 :  62 - 0x3e
      13'h2DC: dout <= 8'b00111111; //  732 :  63 - 0x3f
      13'h2DD: dout <= 8'b00011110; //  733 :  30 - 0x1e
      13'h2DE: dout <= 8'b00001111; //  734 :  15 - 0xf
      13'h2DF: dout <= 8'b00000000; //  735 :   0 - 0x0
      13'h2E0: dout <= 8'b00000000; //  736 :   0 - 0x0 -- Sprite 0x2e
      13'h2E1: dout <= 8'b00000000; //  737 :   0 - 0x0
      13'h2E2: dout <= 8'b00000000; //  738 :   0 - 0x0
      13'h2E3: dout <= 8'b00000000; //  739 :   0 - 0x0
      13'h2E4: dout <= 8'b00000000; //  740 :   0 - 0x0
      13'h2E5: dout <= 8'b00000000; //  741 :   0 - 0x0
      13'h2E6: dout <= 8'b00000000; //  742 :   0 - 0x0
      13'h2E7: dout <= 8'b00000000; //  743 :   0 - 0x0
      13'h2E8: dout <= 8'b00000000; //  744 :   0 - 0x0
      13'h2E9: dout <= 8'b00000000; //  745 :   0 - 0x0
      13'h2EA: dout <= 8'b00000000; //  746 :   0 - 0x0
      13'h2EB: dout <= 8'b00000000; //  747 :   0 - 0x0
      13'h2EC: dout <= 8'b00000000; //  748 :   0 - 0x0
      13'h2ED: dout <= 8'b00000000; //  749 :   0 - 0x0
      13'h2EE: dout <= 8'b00000000; //  750 :   0 - 0x0
      13'h2EF: dout <= 8'b00000000; //  751 :   0 - 0x0
      13'h2F0: dout <= 8'b11110100; //  752 : 244 - 0xf4 -- Sprite 0x2f
      13'h2F1: dout <= 8'b11110010; //  753 : 242 - 0xf2
      13'h2F2: dout <= 8'b11110010; //  754 : 242 - 0xf2
      13'h2F3: dout <= 8'b11110010; //  755 : 242 - 0xf2
      13'h2F4: dout <= 8'b11110010; //  756 : 242 - 0xf2
      13'h2F5: dout <= 8'b11100100; //  757 : 228 - 0xe4
      13'h2F6: dout <= 8'b00001000; //  758 :   8 - 0x8
      13'h2F7: dout <= 8'b11110000; //  759 : 240 - 0xf0
      13'h2F8: dout <= 8'b01111000; //  760 : 120 - 0x78
      13'h2F9: dout <= 8'b01111100; //  761 : 124 - 0x7c
      13'h2FA: dout <= 8'b01111100; //  762 : 124 - 0x7c
      13'h2FB: dout <= 8'b01111100; //  763 : 124 - 0x7c
      13'h2FC: dout <= 8'b11111100; //  764 : 252 - 0xfc
      13'h2FD: dout <= 8'b01111000; //  765 : 120 - 0x78
      13'h2FE: dout <= 8'b11110000; //  766 : 240 - 0xf0
      13'h2FF: dout <= 8'b00000000; //  767 :   0 - 0x0
      13'h300: dout <= 8'b00011000; //  768 :  24 - 0x18 -- Sprite 0x30
      13'h301: dout <= 8'b00100100; //  769 :  36 - 0x24
      13'h302: dout <= 8'b01000010; //  770 :  66 - 0x42
      13'h303: dout <= 8'b10100101; //  771 : 165 - 0xa5
      13'h304: dout <= 8'b11100111; //  772 : 231 - 0xe7
      13'h305: dout <= 8'b00100100; //  773 :  36 - 0x24
      13'h306: dout <= 8'b00100100; //  774 :  36 - 0x24
      13'h307: dout <= 8'b00111100; //  775 :  60 - 0x3c
      13'h308: dout <= 8'b00000000; //  776 :   0 - 0x0
      13'h309: dout <= 8'b00011000; //  777 :  24 - 0x18
      13'h30A: dout <= 8'b00111100; //  778 :  60 - 0x3c
      13'h30B: dout <= 8'b01011010; //  779 :  90 - 0x5a
      13'h30C: dout <= 8'b00011000; //  780 :  24 - 0x18
      13'h30D: dout <= 8'b00011000; //  781 :  24 - 0x18
      13'h30E: dout <= 8'b00011000; //  782 :  24 - 0x18
      13'h30F: dout <= 8'b00000000; //  783 :   0 - 0x0
      13'h310: dout <= 8'b00111100; //  784 :  60 - 0x3c -- Sprite 0x31
      13'h311: dout <= 8'b00100100; //  785 :  36 - 0x24
      13'h312: dout <= 8'b00100100; //  786 :  36 - 0x24
      13'h313: dout <= 8'b01100110; //  787 : 102 - 0x66
      13'h314: dout <= 8'b10100101; //  788 : 165 - 0xa5
      13'h315: dout <= 8'b01000010; //  789 :  66 - 0x42
      13'h316: dout <= 8'b00100100; //  790 :  36 - 0x24
      13'h317: dout <= 8'b00011000; //  791 :  24 - 0x18
      13'h318: dout <= 8'b00000000; //  792 :   0 - 0x0
      13'h319: dout <= 8'b00011000; //  793 :  24 - 0x18
      13'h31A: dout <= 8'b00011000; //  794 :  24 - 0x18
      13'h31B: dout <= 8'b00011000; //  795 :  24 - 0x18
      13'h31C: dout <= 8'b01011010; //  796 :  90 - 0x5a
      13'h31D: dout <= 8'b00111100; //  797 :  60 - 0x3c
      13'h31E: dout <= 8'b00011000; //  798 :  24 - 0x18
      13'h31F: dout <= 8'b00000000; //  799 :   0 - 0x0
      13'h320: dout <= 8'b00000010; //  800 :   2 - 0x2 -- Sprite 0x32
      13'h321: dout <= 8'b00000010; //  801 :   2 - 0x2
      13'h322: dout <= 8'b00000011; //  802 :   3 - 0x3
      13'h323: dout <= 8'b00000010; //  803 :   2 - 0x2
      13'h324: dout <= 8'b00000010; //  804 :   2 - 0x2
      13'h325: dout <= 8'b00000010; //  805 :   2 - 0x2
      13'h326: dout <= 8'b00000011; //  806 :   3 - 0x3
      13'h327: dout <= 8'b00000010; //  807 :   2 - 0x2
      13'h328: dout <= 8'b00000001; //  808 :   1 - 0x1
      13'h329: dout <= 8'b00000001; //  809 :   1 - 0x1
      13'h32A: dout <= 8'b00000000; //  810 :   0 - 0x0
      13'h32B: dout <= 8'b00000001; //  811 :   1 - 0x1
      13'h32C: dout <= 8'b00000001; //  812 :   1 - 0x1
      13'h32D: dout <= 8'b00000001; //  813 :   1 - 0x1
      13'h32E: dout <= 8'b00000000; //  814 :   0 - 0x0
      13'h32F: dout <= 8'b00000001; //  815 :   1 - 0x1
      13'h330: dout <= 8'b01000000; //  816 :  64 - 0x40 -- Sprite 0x33
      13'h331: dout <= 8'b11000000; //  817 : 192 - 0xc0
      13'h332: dout <= 8'b01000000; //  818 :  64 - 0x40
      13'h333: dout <= 8'b01000000; //  819 :  64 - 0x40
      13'h334: dout <= 8'b01000000; //  820 :  64 - 0x40
      13'h335: dout <= 8'b11000000; //  821 : 192 - 0xc0
      13'h336: dout <= 8'b01000000; //  822 :  64 - 0x40
      13'h337: dout <= 8'b01000000; //  823 :  64 - 0x40
      13'h338: dout <= 8'b10000000; //  824 : 128 - 0x80
      13'h339: dout <= 8'b00000000; //  825 :   0 - 0x0
      13'h33A: dout <= 8'b10000000; //  826 : 128 - 0x80
      13'h33B: dout <= 8'b10000000; //  827 : 128 - 0x80
      13'h33C: dout <= 8'b10000000; //  828 : 128 - 0x80
      13'h33D: dout <= 8'b00000000; //  829 :   0 - 0x0
      13'h33E: dout <= 8'b10000000; //  830 : 128 - 0x80
      13'h33F: dout <= 8'b10000000; //  831 : 128 - 0x80
      13'h340: dout <= 8'b00000000; //  832 :   0 - 0x0 -- Sprite 0x34
      13'h341: dout <= 8'b00011000; //  833 :  24 - 0x18
      13'h342: dout <= 8'b00111100; //  834 :  60 - 0x3c
      13'h343: dout <= 8'b01100010; //  835 :  98 - 0x62
      13'h344: dout <= 8'b01100001; //  836 :  97 - 0x61
      13'h345: dout <= 8'b11000000; //  837 : 192 - 0xc0
      13'h346: dout <= 8'b11000000; //  838 : 192 - 0xc0
      13'h347: dout <= 8'b11000000; //  839 : 192 - 0xc0
      13'h348: dout <= 8'b00000000; //  840 :   0 - 0x0
      13'h349: dout <= 8'b00000000; //  841 :   0 - 0x0
      13'h34A: dout <= 8'b00011000; //  842 :  24 - 0x18
      13'h34B: dout <= 8'b00111100; //  843 :  60 - 0x3c
      13'h34C: dout <= 8'b00111110; //  844 :  62 - 0x3e
      13'h34D: dout <= 8'b01111111; //  845 : 127 - 0x7f
      13'h34E: dout <= 8'b01111111; //  846 : 127 - 0x7f
      13'h34F: dout <= 8'b01111111; //  847 : 127 - 0x7f
      13'h350: dout <= 8'b01100000; //  848 :  96 - 0x60 -- Sprite 0x35
      13'h351: dout <= 8'b01100000; //  849 :  96 - 0x60
      13'h352: dout <= 8'b00110000; //  850 :  48 - 0x30
      13'h353: dout <= 8'b00011000; //  851 :  24 - 0x18
      13'h354: dout <= 8'b00001100; //  852 :  12 - 0xc
      13'h355: dout <= 8'b00000110; //  853 :   6 - 0x6
      13'h356: dout <= 8'b00000010; //  854 :   2 - 0x2
      13'h357: dout <= 8'b00000001; //  855 :   1 - 0x1
      13'h358: dout <= 8'b00111111; //  856 :  63 - 0x3f
      13'h359: dout <= 8'b00111111; //  857 :  63 - 0x3f
      13'h35A: dout <= 8'b00011111; //  858 :  31 - 0x1f
      13'h35B: dout <= 8'b00001111; //  859 :  15 - 0xf
      13'h35C: dout <= 8'b00000111; //  860 :   7 - 0x7
      13'h35D: dout <= 8'b00000011; //  861 :   3 - 0x3
      13'h35E: dout <= 8'b00000001; //  862 :   1 - 0x1
      13'h35F: dout <= 8'b00000000; //  863 :   0 - 0x0
      13'h360: dout <= 8'b00000000; //  864 :   0 - 0x0 -- Sprite 0x36
      13'h361: dout <= 8'b00011000; //  865 :  24 - 0x18
      13'h362: dout <= 8'b00100100; //  866 :  36 - 0x24
      13'h363: dout <= 8'b01000010; //  867 :  66 - 0x42
      13'h364: dout <= 8'b10000010; //  868 : 130 - 0x82
      13'h365: dout <= 8'b00000001; //  869 :   1 - 0x1
      13'h366: dout <= 8'b00000001; //  870 :   1 - 0x1
      13'h367: dout <= 8'b00000001; //  871 :   1 - 0x1
      13'h368: dout <= 8'b00000000; //  872 :   0 - 0x0
      13'h369: dout <= 8'b00000000; //  873 :   0 - 0x0
      13'h36A: dout <= 8'b00011000; //  874 :  24 - 0x18
      13'h36B: dout <= 8'b00111100; //  875 :  60 - 0x3c
      13'h36C: dout <= 8'b01111100; //  876 : 124 - 0x7c
      13'h36D: dout <= 8'b11111110; //  877 : 254 - 0xfe
      13'h36E: dout <= 8'b11111110; //  878 : 254 - 0xfe
      13'h36F: dout <= 8'b11111110; //  879 : 254 - 0xfe
      13'h370: dout <= 8'b00000010; //  880 :   2 - 0x2 -- Sprite 0x37
      13'h371: dout <= 8'b00000010; //  881 :   2 - 0x2
      13'h372: dout <= 8'b00000100; //  882 :   4 - 0x4
      13'h373: dout <= 8'b00001000; //  883 :   8 - 0x8
      13'h374: dout <= 8'b00010000; //  884 :  16 - 0x10
      13'h375: dout <= 8'b00100000; //  885 :  32 - 0x20
      13'h376: dout <= 8'b01000000; //  886 :  64 - 0x40
      13'h377: dout <= 8'b10000000; //  887 : 128 - 0x80
      13'h378: dout <= 8'b11111100; //  888 : 252 - 0xfc
      13'h379: dout <= 8'b11111100; //  889 : 252 - 0xfc
      13'h37A: dout <= 8'b11111000; //  890 : 248 - 0xf8
      13'h37B: dout <= 8'b11110000; //  891 : 240 - 0xf0
      13'h37C: dout <= 8'b11100000; //  892 : 224 - 0xe0
      13'h37D: dout <= 8'b11000000; //  893 : 192 - 0xc0
      13'h37E: dout <= 8'b10000000; //  894 : 128 - 0x80
      13'h37F: dout <= 8'b00000000; //  895 :   0 - 0x0
      13'h380: dout <= 8'b00000000; //  896 :   0 - 0x0 -- Sprite 0x38
      13'h381: dout <= 8'b00000110; //  897 :   6 - 0x6
      13'h382: dout <= 8'b00001101; //  898 :  13 - 0xd
      13'h383: dout <= 8'b00001100; //  899 :  12 - 0xc
      13'h384: dout <= 8'b00001100; //  900 :  12 - 0xc
      13'h385: dout <= 8'b00000110; //  901 :   6 - 0x6
      13'h386: dout <= 8'b00000010; //  902 :   2 - 0x2
      13'h387: dout <= 8'b00000001; //  903 :   1 - 0x1
      13'h388: dout <= 8'b00000000; //  904 :   0 - 0x0
      13'h389: dout <= 8'b00000000; //  905 :   0 - 0x0
      13'h38A: dout <= 8'b00000110; //  906 :   6 - 0x6
      13'h38B: dout <= 8'b00000111; //  907 :   7 - 0x7
      13'h38C: dout <= 8'b00000111; //  908 :   7 - 0x7
      13'h38D: dout <= 8'b00000011; //  909 :   3 - 0x3
      13'h38E: dout <= 8'b00000001; //  910 :   1 - 0x1
      13'h38F: dout <= 8'b00000000; //  911 :   0 - 0x0
      13'h390: dout <= 8'b11111111; //  912 : 255 - 0xff -- Sprite 0x39
      13'h391: dout <= 8'b00000000; //  913 :   0 - 0x0
      13'h392: dout <= 8'b00000000; //  914 :   0 - 0x0
      13'h393: dout <= 8'b00000000; //  915 :   0 - 0x0
      13'h394: dout <= 8'b00000000; //  916 :   0 - 0x0
      13'h395: dout <= 8'b00000000; //  917 :   0 - 0x0
      13'h396: dout <= 8'b00000000; //  918 :   0 - 0x0
      13'h397: dout <= 8'b00000000; //  919 :   0 - 0x0
      13'h398: dout <= 8'b00000000; //  920 :   0 - 0x0
      13'h399: dout <= 8'b00000000; //  921 :   0 - 0x0
      13'h39A: dout <= 8'b00000000; //  922 :   0 - 0x0
      13'h39B: dout <= 8'b00000000; //  923 :   0 - 0x0
      13'h39C: dout <= 8'b00000000; //  924 :   0 - 0x0
      13'h39D: dout <= 8'b00000000; //  925 :   0 - 0x0
      13'h39E: dout <= 8'b00000000; //  926 :   0 - 0x0
      13'h39F: dout <= 8'b00000000; //  927 :   0 - 0x0
      13'h3A0: dout <= 8'b00000000; //  928 :   0 - 0x0 -- Sprite 0x3a
      13'h3A1: dout <= 8'b01100000; //  929 :  96 - 0x60
      13'h3A2: dout <= 8'b10010000; //  930 : 144 - 0x90
      13'h3A3: dout <= 8'b00010000; //  931 :  16 - 0x10
      13'h3A4: dout <= 8'b00010000; //  932 :  16 - 0x10
      13'h3A5: dout <= 8'b00100000; //  933 :  32 - 0x20
      13'h3A6: dout <= 8'b01000000; //  934 :  64 - 0x40
      13'h3A7: dout <= 8'b10000000; //  935 : 128 - 0x80
      13'h3A8: dout <= 8'b00000000; //  936 :   0 - 0x0
      13'h3A9: dout <= 8'b00000000; //  937 :   0 - 0x0
      13'h3AA: dout <= 8'b01100000; //  938 :  96 - 0x60
      13'h3AB: dout <= 8'b11100000; //  939 : 224 - 0xe0
      13'h3AC: dout <= 8'b11100000; //  940 : 224 - 0xe0
      13'h3AD: dout <= 8'b11000000; //  941 : 192 - 0xc0
      13'h3AE: dout <= 8'b10000000; //  942 : 128 - 0x80
      13'h3AF: dout <= 8'b00000000; //  943 :   0 - 0x0
      13'h3B0: dout <= 8'b00000000; //  944 :   0 - 0x0 -- Sprite 0x3b
      13'h3B1: dout <= 8'b01010100; //  945 :  84 - 0x54
      13'h3B2: dout <= 8'b00000010; //  946 :   2 - 0x2
      13'h3B3: dout <= 8'b01000000; //  947 :  64 - 0x40
      13'h3B4: dout <= 8'b00000010; //  948 :   2 - 0x2
      13'h3B5: dout <= 8'b01000000; //  949 :  64 - 0x40
      13'h3B6: dout <= 8'b00101010; //  950 :  42 - 0x2a
      13'h3B7: dout <= 8'b00000000; //  951 :   0 - 0x0
      13'h3B8: dout <= 8'b00000000; //  952 :   0 - 0x0
      13'h3B9: dout <= 8'b00101010; //  953 :  42 - 0x2a
      13'h3BA: dout <= 8'b01000000; //  954 :  64 - 0x40
      13'h3BB: dout <= 8'b00000010; //  955 :   2 - 0x2
      13'h3BC: dout <= 8'b01000000; //  956 :  64 - 0x40
      13'h3BD: dout <= 8'b00000010; //  957 :   2 - 0x2
      13'h3BE: dout <= 8'b01010100; //  958 :  84 - 0x54
      13'h3BF: dout <= 8'b00000000; //  959 :   0 - 0x0
      13'h3C0: dout <= 8'b11111111; //  960 : 255 - 0xff -- Sprite 0x3c
      13'h3C1: dout <= 8'b11111111; //  961 : 255 - 0xff
      13'h3C2: dout <= 8'b11111111; //  962 : 255 - 0xff
      13'h3C3: dout <= 8'b11111111; //  963 : 255 - 0xff
      13'h3C4: dout <= 8'b11111111; //  964 : 255 - 0xff
      13'h3C5: dout <= 8'b11111111; //  965 : 255 - 0xff
      13'h3C6: dout <= 8'b11111111; //  966 : 255 - 0xff
      13'h3C7: dout <= 8'b11111111; //  967 : 255 - 0xff
      13'h3C8: dout <= 8'b00000000; //  968 :   0 - 0x0
      13'h3C9: dout <= 8'b00000000; //  969 :   0 - 0x0
      13'h3CA: dout <= 8'b00000000; //  970 :   0 - 0x0
      13'h3CB: dout <= 8'b00000000; //  971 :   0 - 0x0
      13'h3CC: dout <= 8'b00000000; //  972 :   0 - 0x0
      13'h3CD: dout <= 8'b00000000; //  973 :   0 - 0x0
      13'h3CE: dout <= 8'b00000000; //  974 :   0 - 0x0
      13'h3CF: dout <= 8'b00000000; //  975 :   0 - 0x0
      13'h3D0: dout <= 8'b00000000; //  976 :   0 - 0x0 -- Sprite 0x3d
      13'h3D1: dout <= 8'b00000000; //  977 :   0 - 0x0
      13'h3D2: dout <= 8'b00000000; //  978 :   0 - 0x0
      13'h3D3: dout <= 8'b00000000; //  979 :   0 - 0x0
      13'h3D4: dout <= 8'b00000000; //  980 :   0 - 0x0
      13'h3D5: dout <= 8'b00000000; //  981 :   0 - 0x0
      13'h3D6: dout <= 8'b00000000; //  982 :   0 - 0x0
      13'h3D7: dout <= 8'b00000000; //  983 :   0 - 0x0
      13'h3D8: dout <= 8'b11111111; //  984 : 255 - 0xff
      13'h3D9: dout <= 8'b11111111; //  985 : 255 - 0xff
      13'h3DA: dout <= 8'b11111111; //  986 : 255 - 0xff
      13'h3DB: dout <= 8'b11111111; //  987 : 255 - 0xff
      13'h3DC: dout <= 8'b11111111; //  988 : 255 - 0xff
      13'h3DD: dout <= 8'b11111111; //  989 : 255 - 0xff
      13'h3DE: dout <= 8'b11111111; //  990 : 255 - 0xff
      13'h3DF: dout <= 8'b11111111; //  991 : 255 - 0xff
      13'h3E0: dout <= 8'b11111111; //  992 : 255 - 0xff -- Sprite 0x3e
      13'h3E1: dout <= 8'b11111111; //  993 : 255 - 0xff
      13'h3E2: dout <= 8'b11111111; //  994 : 255 - 0xff
      13'h3E3: dout <= 8'b11111111; //  995 : 255 - 0xff
      13'h3E4: dout <= 8'b11111111; //  996 : 255 - 0xff
      13'h3E5: dout <= 8'b11111111; //  997 : 255 - 0xff
      13'h3E6: dout <= 8'b11111111; //  998 : 255 - 0xff
      13'h3E7: dout <= 8'b11111111; //  999 : 255 - 0xff
      13'h3E8: dout <= 8'b11111111; // 1000 : 255 - 0xff
      13'h3E9: dout <= 8'b11111111; // 1001 : 255 - 0xff
      13'h3EA: dout <= 8'b11111111; // 1002 : 255 - 0xff
      13'h3EB: dout <= 8'b11111111; // 1003 : 255 - 0xff
      13'h3EC: dout <= 8'b11111111; // 1004 : 255 - 0xff
      13'h3ED: dout <= 8'b11111111; // 1005 : 255 - 0xff
      13'h3EE: dout <= 8'b11111111; // 1006 : 255 - 0xff
      13'h3EF: dout <= 8'b11111111; // 1007 : 255 - 0xff
      13'h3F0: dout <= 8'b00000000; // 1008 :   0 - 0x0 -- Sprite 0x3f
      13'h3F1: dout <= 8'b00000000; // 1009 :   0 - 0x0
      13'h3F2: dout <= 8'b00000000; // 1010 :   0 - 0x0
      13'h3F3: dout <= 8'b00000000; // 1011 :   0 - 0x0
      13'h3F4: dout <= 8'b00000000; // 1012 :   0 - 0x0
      13'h3F5: dout <= 8'b00000000; // 1013 :   0 - 0x0
      13'h3F6: dout <= 8'b00000000; // 1014 :   0 - 0x0
      13'h3F7: dout <= 8'b00000000; // 1015 :   0 - 0x0
      13'h3F8: dout <= 8'b00000000; // 1016 :   0 - 0x0
      13'h3F9: dout <= 8'b00000000; // 1017 :   0 - 0x0
      13'h3FA: dout <= 8'b00000000; // 1018 :   0 - 0x0
      13'h3FB: dout <= 8'b00000000; // 1019 :   0 - 0x0
      13'h3FC: dout <= 8'b00000000; // 1020 :   0 - 0x0
      13'h3FD: dout <= 8'b00000000; // 1021 :   0 - 0x0
      13'h3FE: dout <= 8'b00000000; // 1022 :   0 - 0x0
      13'h3FF: dout <= 8'b00000000; // 1023 :   0 - 0x0
      13'h400: dout <= 8'b00111100; // 1024 :  60 - 0x3c -- Sprite 0x40
      13'h401: dout <= 8'b01000010; // 1025 :  66 - 0x42
      13'h402: dout <= 8'b10011001; // 1026 : 153 - 0x99
      13'h403: dout <= 8'b10100101; // 1027 : 165 - 0xa5
      13'h404: dout <= 8'b10100101; // 1028 : 165 - 0xa5
      13'h405: dout <= 8'b10011010; // 1029 : 154 - 0x9a
      13'h406: dout <= 8'b01000000; // 1030 :  64 - 0x40
      13'h407: dout <= 8'b00111100; // 1031 :  60 - 0x3c
      13'h408: dout <= 8'b00000000; // 1032 :   0 - 0x0
      13'h409: dout <= 8'b00000000; // 1033 :   0 - 0x0
      13'h40A: dout <= 8'b00000000; // 1034 :   0 - 0x0
      13'h40B: dout <= 8'b00000000; // 1035 :   0 - 0x0
      13'h40C: dout <= 8'b00000000; // 1036 :   0 - 0x0
      13'h40D: dout <= 8'b00000000; // 1037 :   0 - 0x0
      13'h40E: dout <= 8'b00000000; // 1038 :   0 - 0x0
      13'h40F: dout <= 8'b00000000; // 1039 :   0 - 0x0
      13'h410: dout <= 8'b00001100; // 1040 :  12 - 0xc -- Sprite 0x41
      13'h411: dout <= 8'b00010010; // 1041 :  18 - 0x12
      13'h412: dout <= 8'b00100010; // 1042 :  34 - 0x22
      13'h413: dout <= 8'b00100010; // 1043 :  34 - 0x22
      13'h414: dout <= 8'b01111110; // 1044 : 126 - 0x7e
      13'h415: dout <= 8'b00100010; // 1045 :  34 - 0x22
      13'h416: dout <= 8'b00100100; // 1046 :  36 - 0x24
      13'h417: dout <= 8'b00000000; // 1047 :   0 - 0x0
      13'h418: dout <= 8'b00000000; // 1048 :   0 - 0x0
      13'h419: dout <= 8'b00000000; // 1049 :   0 - 0x0
      13'h41A: dout <= 8'b00000000; // 1050 :   0 - 0x0
      13'h41B: dout <= 8'b00000000; // 1051 :   0 - 0x0
      13'h41C: dout <= 8'b00000000; // 1052 :   0 - 0x0
      13'h41D: dout <= 8'b00000000; // 1053 :   0 - 0x0
      13'h41E: dout <= 8'b00000000; // 1054 :   0 - 0x0
      13'h41F: dout <= 8'b00000000; // 1055 :   0 - 0x0
      13'h420: dout <= 8'b00111100; // 1056 :  60 - 0x3c -- Sprite 0x42
      13'h421: dout <= 8'b01000010; // 1057 :  66 - 0x42
      13'h422: dout <= 8'b01010010; // 1058 :  82 - 0x52
      13'h423: dout <= 8'b00011100; // 1059 :  28 - 0x1c
      13'h424: dout <= 8'b00010010; // 1060 :  18 - 0x12
      13'h425: dout <= 8'b00110010; // 1061 :  50 - 0x32
      13'h426: dout <= 8'b00011100; // 1062 :  28 - 0x1c
      13'h427: dout <= 8'b00000000; // 1063 :   0 - 0x0
      13'h428: dout <= 8'b00000000; // 1064 :   0 - 0x0
      13'h429: dout <= 8'b00000000; // 1065 :   0 - 0x0
      13'h42A: dout <= 8'b00000000; // 1066 :   0 - 0x0
      13'h42B: dout <= 8'b00000000; // 1067 :   0 - 0x0
      13'h42C: dout <= 8'b00000000; // 1068 :   0 - 0x0
      13'h42D: dout <= 8'b00000000; // 1069 :   0 - 0x0
      13'h42E: dout <= 8'b00000000; // 1070 :   0 - 0x0
      13'h42F: dout <= 8'b00000000; // 1071 :   0 - 0x0
      13'h430: dout <= 8'b00011000; // 1072 :  24 - 0x18 -- Sprite 0x43
      13'h431: dout <= 8'b00100100; // 1073 :  36 - 0x24
      13'h432: dout <= 8'b01010100; // 1074 :  84 - 0x54
      13'h433: dout <= 8'b01001000; // 1075 :  72 - 0x48
      13'h434: dout <= 8'b01000010; // 1076 :  66 - 0x42
      13'h435: dout <= 8'b00100100; // 1077 :  36 - 0x24
      13'h436: dout <= 8'b00011000; // 1078 :  24 - 0x18
      13'h437: dout <= 8'b00000000; // 1079 :   0 - 0x0
      13'h438: dout <= 8'b00000000; // 1080 :   0 - 0x0
      13'h439: dout <= 8'b00000000; // 1081 :   0 - 0x0
      13'h43A: dout <= 8'b00000000; // 1082 :   0 - 0x0
      13'h43B: dout <= 8'b00000000; // 1083 :   0 - 0x0
      13'h43C: dout <= 8'b00000000; // 1084 :   0 - 0x0
      13'h43D: dout <= 8'b00000000; // 1085 :   0 - 0x0
      13'h43E: dout <= 8'b00000000; // 1086 :   0 - 0x0
      13'h43F: dout <= 8'b00000000; // 1087 :   0 - 0x0
      13'h440: dout <= 8'b01011000; // 1088 :  88 - 0x58 -- Sprite 0x44
      13'h441: dout <= 8'b11100100; // 1089 : 228 - 0xe4
      13'h442: dout <= 8'b01000010; // 1090 :  66 - 0x42
      13'h443: dout <= 8'b01000010; // 1091 :  66 - 0x42
      13'h444: dout <= 8'b00100010; // 1092 :  34 - 0x22
      13'h445: dout <= 8'b01100100; // 1093 : 100 - 0x64
      13'h446: dout <= 8'b00111000; // 1094 :  56 - 0x38
      13'h447: dout <= 8'b00000000; // 1095 :   0 - 0x0
      13'h448: dout <= 8'b00000000; // 1096 :   0 - 0x0
      13'h449: dout <= 8'b00000000; // 1097 :   0 - 0x0
      13'h44A: dout <= 8'b00000000; // 1098 :   0 - 0x0
      13'h44B: dout <= 8'b00000000; // 1099 :   0 - 0x0
      13'h44C: dout <= 8'b00000000; // 1100 :   0 - 0x0
      13'h44D: dout <= 8'b00000000; // 1101 :   0 - 0x0
      13'h44E: dout <= 8'b00000000; // 1102 :   0 - 0x0
      13'h44F: dout <= 8'b00000000; // 1103 :   0 - 0x0
      13'h450: dout <= 8'b00011100; // 1104 :  28 - 0x1c -- Sprite 0x45
      13'h451: dout <= 8'b00100000; // 1105 :  32 - 0x20
      13'h452: dout <= 8'b00100000; // 1106 :  32 - 0x20
      13'h453: dout <= 8'b00101100; // 1107 :  44 - 0x2c
      13'h454: dout <= 8'b01110000; // 1108 : 112 - 0x70
      13'h455: dout <= 8'b00100010; // 1109 :  34 - 0x22
      13'h456: dout <= 8'b00011100; // 1110 :  28 - 0x1c
      13'h457: dout <= 8'b00000000; // 1111 :   0 - 0x0
      13'h458: dout <= 8'b00000000; // 1112 :   0 - 0x0
      13'h459: dout <= 8'b00000000; // 1113 :   0 - 0x0
      13'h45A: dout <= 8'b00000000; // 1114 :   0 - 0x0
      13'h45B: dout <= 8'b00000000; // 1115 :   0 - 0x0
      13'h45C: dout <= 8'b00000000; // 1116 :   0 - 0x0
      13'h45D: dout <= 8'b00000000; // 1117 :   0 - 0x0
      13'h45E: dout <= 8'b00000000; // 1118 :   0 - 0x0
      13'h45F: dout <= 8'b00000000; // 1119 :   0 - 0x0
      13'h460: dout <= 8'b00011100; // 1120 :  28 - 0x1c -- Sprite 0x46
      13'h461: dout <= 8'b00100000; // 1121 :  32 - 0x20
      13'h462: dout <= 8'b00100000; // 1122 :  32 - 0x20
      13'h463: dout <= 8'b00101100; // 1123 :  44 - 0x2c
      13'h464: dout <= 8'b01110000; // 1124 : 112 - 0x70
      13'h465: dout <= 8'b00010000; // 1125 :  16 - 0x10
      13'h466: dout <= 8'b00010000; // 1126 :  16 - 0x10
      13'h467: dout <= 8'b00000000; // 1127 :   0 - 0x0
      13'h468: dout <= 8'b00000000; // 1128 :   0 - 0x0
      13'h469: dout <= 8'b00000000; // 1129 :   0 - 0x0
      13'h46A: dout <= 8'b00000000; // 1130 :   0 - 0x0
      13'h46B: dout <= 8'b00000000; // 1131 :   0 - 0x0
      13'h46C: dout <= 8'b00000000; // 1132 :   0 - 0x0
      13'h46D: dout <= 8'b00000000; // 1133 :   0 - 0x0
      13'h46E: dout <= 8'b00000000; // 1134 :   0 - 0x0
      13'h46F: dout <= 8'b00000000; // 1135 :   0 - 0x0
      13'h470: dout <= 8'b00011000; // 1136 :  24 - 0x18 -- Sprite 0x47
      13'h471: dout <= 8'b00100100; // 1137 :  36 - 0x24
      13'h472: dout <= 8'b01000000; // 1138 :  64 - 0x40
      13'h473: dout <= 8'b01001110; // 1139 :  78 - 0x4e
      13'h474: dout <= 8'b01000010; // 1140 :  66 - 0x42
      13'h475: dout <= 8'b00100100; // 1141 :  36 - 0x24
      13'h476: dout <= 8'b00011000; // 1142 :  24 - 0x18
      13'h477: dout <= 8'b00000000; // 1143 :   0 - 0x0
      13'h478: dout <= 8'b00000000; // 1144 :   0 - 0x0
      13'h479: dout <= 8'b00000000; // 1145 :   0 - 0x0
      13'h47A: dout <= 8'b00000000; // 1146 :   0 - 0x0
      13'h47B: dout <= 8'b00000000; // 1147 :   0 - 0x0
      13'h47C: dout <= 8'b00000000; // 1148 :   0 - 0x0
      13'h47D: dout <= 8'b00000000; // 1149 :   0 - 0x0
      13'h47E: dout <= 8'b00000000; // 1150 :   0 - 0x0
      13'h47F: dout <= 8'b00000000; // 1151 :   0 - 0x0
      13'h480: dout <= 8'b00100000; // 1152 :  32 - 0x20 -- Sprite 0x48
      13'h481: dout <= 8'b01000100; // 1153 :  68 - 0x44
      13'h482: dout <= 8'b01000100; // 1154 :  68 - 0x44
      13'h483: dout <= 8'b01000100; // 1155 :  68 - 0x44
      13'h484: dout <= 8'b11111100; // 1156 : 252 - 0xfc
      13'h485: dout <= 8'b01000100; // 1157 :  68 - 0x44
      13'h486: dout <= 8'b01001000; // 1158 :  72 - 0x48
      13'h487: dout <= 8'b00000000; // 1159 :   0 - 0x0
      13'h488: dout <= 8'b00000000; // 1160 :   0 - 0x0
      13'h489: dout <= 8'b00000000; // 1161 :   0 - 0x0
      13'h48A: dout <= 8'b00000000; // 1162 :   0 - 0x0
      13'h48B: dout <= 8'b00000000; // 1163 :   0 - 0x0
      13'h48C: dout <= 8'b00000000; // 1164 :   0 - 0x0
      13'h48D: dout <= 8'b00000000; // 1165 :   0 - 0x0
      13'h48E: dout <= 8'b00000000; // 1166 :   0 - 0x0
      13'h48F: dout <= 8'b00000000; // 1167 :   0 - 0x0
      13'h490: dout <= 8'b00010000; // 1168 :  16 - 0x10 -- Sprite 0x49
      13'h491: dout <= 8'b00010000; // 1169 :  16 - 0x10
      13'h492: dout <= 8'b00010000; // 1170 :  16 - 0x10
      13'h493: dout <= 8'b00010000; // 1171 :  16 - 0x10
      13'h494: dout <= 8'b00010000; // 1172 :  16 - 0x10
      13'h495: dout <= 8'b00001000; // 1173 :   8 - 0x8
      13'h496: dout <= 8'b00001000; // 1174 :   8 - 0x8
      13'h497: dout <= 8'b00000000; // 1175 :   0 - 0x0
      13'h498: dout <= 8'b00000000; // 1176 :   0 - 0x0
      13'h499: dout <= 8'b00000000; // 1177 :   0 - 0x0
      13'h49A: dout <= 8'b00000000; // 1178 :   0 - 0x0
      13'h49B: dout <= 8'b00000000; // 1179 :   0 - 0x0
      13'h49C: dout <= 8'b00000000; // 1180 :   0 - 0x0
      13'h49D: dout <= 8'b00000000; // 1181 :   0 - 0x0
      13'h49E: dout <= 8'b00000000; // 1182 :   0 - 0x0
      13'h49F: dout <= 8'b00000000; // 1183 :   0 - 0x0
      13'h4A0: dout <= 8'b00001000; // 1184 :   8 - 0x8 -- Sprite 0x4a
      13'h4A1: dout <= 8'b00001000; // 1185 :   8 - 0x8
      13'h4A2: dout <= 8'b00000100; // 1186 :   4 - 0x4
      13'h4A3: dout <= 8'b00000100; // 1187 :   4 - 0x4
      13'h4A4: dout <= 8'b01000100; // 1188 :  68 - 0x44
      13'h4A5: dout <= 8'b01001000; // 1189 :  72 - 0x48
      13'h4A6: dout <= 8'b00110000; // 1190 :  48 - 0x30
      13'h4A7: dout <= 8'b00000000; // 1191 :   0 - 0x0
      13'h4A8: dout <= 8'b00000000; // 1192 :   0 - 0x0
      13'h4A9: dout <= 8'b00000000; // 1193 :   0 - 0x0
      13'h4AA: dout <= 8'b00000000; // 1194 :   0 - 0x0
      13'h4AB: dout <= 8'b00000000; // 1195 :   0 - 0x0
      13'h4AC: dout <= 8'b00000000; // 1196 :   0 - 0x0
      13'h4AD: dout <= 8'b00000000; // 1197 :   0 - 0x0
      13'h4AE: dout <= 8'b00000000; // 1198 :   0 - 0x0
      13'h4AF: dout <= 8'b00000000; // 1199 :   0 - 0x0
      13'h4B0: dout <= 8'b01000100; // 1200 :  68 - 0x44 -- Sprite 0x4b
      13'h4B1: dout <= 8'b01000100; // 1201 :  68 - 0x44
      13'h4B2: dout <= 8'b01001000; // 1202 :  72 - 0x48
      13'h4B3: dout <= 8'b01110000; // 1203 : 112 - 0x70
      13'h4B4: dout <= 8'b01001000; // 1204 :  72 - 0x48
      13'h4B5: dout <= 8'b00100100; // 1205 :  36 - 0x24
      13'h4B6: dout <= 8'b00100010; // 1206 :  34 - 0x22
      13'h4B7: dout <= 8'b00000000; // 1207 :   0 - 0x0
      13'h4B8: dout <= 8'b00000000; // 1208 :   0 - 0x0
      13'h4B9: dout <= 8'b00000000; // 1209 :   0 - 0x0
      13'h4BA: dout <= 8'b00000000; // 1210 :   0 - 0x0
      13'h4BB: dout <= 8'b00000000; // 1211 :   0 - 0x0
      13'h4BC: dout <= 8'b00000000; // 1212 :   0 - 0x0
      13'h4BD: dout <= 8'b00000000; // 1213 :   0 - 0x0
      13'h4BE: dout <= 8'b00000000; // 1214 :   0 - 0x0
      13'h4BF: dout <= 8'b00000000; // 1215 :   0 - 0x0
      13'h4C0: dout <= 8'b00010000; // 1216 :  16 - 0x10 -- Sprite 0x4c
      13'h4C1: dout <= 8'b00100000; // 1217 :  32 - 0x20
      13'h4C2: dout <= 8'b00100000; // 1218 :  32 - 0x20
      13'h4C3: dout <= 8'b00100000; // 1219 :  32 - 0x20
      13'h4C4: dout <= 8'b01000000; // 1220 :  64 - 0x40
      13'h4C5: dout <= 8'b01000000; // 1221 :  64 - 0x40
      13'h4C6: dout <= 8'b01000110; // 1222 :  70 - 0x46
      13'h4C7: dout <= 8'b00111000; // 1223 :  56 - 0x38
      13'h4C8: dout <= 8'b00000000; // 1224 :   0 - 0x0
      13'h4C9: dout <= 8'b00000000; // 1225 :   0 - 0x0
      13'h4CA: dout <= 8'b00000000; // 1226 :   0 - 0x0
      13'h4CB: dout <= 8'b00000000; // 1227 :   0 - 0x0
      13'h4CC: dout <= 8'b00000000; // 1228 :   0 - 0x0
      13'h4CD: dout <= 8'b00000000; // 1229 :   0 - 0x0
      13'h4CE: dout <= 8'b00000000; // 1230 :   0 - 0x0
      13'h4CF: dout <= 8'b00000000; // 1231 :   0 - 0x0
      13'h4D0: dout <= 8'b00100100; // 1232 :  36 - 0x24 -- Sprite 0x4d
      13'h4D1: dout <= 8'b01011010; // 1233 :  90 - 0x5a
      13'h4D2: dout <= 8'b01011010; // 1234 :  90 - 0x5a
      13'h4D3: dout <= 8'b01011010; // 1235 :  90 - 0x5a
      13'h4D4: dout <= 8'b01000010; // 1236 :  66 - 0x42
      13'h4D5: dout <= 8'b01000010; // 1237 :  66 - 0x42
      13'h4D6: dout <= 8'b00100010; // 1238 :  34 - 0x22
      13'h4D7: dout <= 8'b00000000; // 1239 :   0 - 0x0
      13'h4D8: dout <= 8'b00000000; // 1240 :   0 - 0x0
      13'h4D9: dout <= 8'b00000000; // 1241 :   0 - 0x0
      13'h4DA: dout <= 8'b00000000; // 1242 :   0 - 0x0
      13'h4DB: dout <= 8'b00000000; // 1243 :   0 - 0x0
      13'h4DC: dout <= 8'b00000000; // 1244 :   0 - 0x0
      13'h4DD: dout <= 8'b00000000; // 1245 :   0 - 0x0
      13'h4DE: dout <= 8'b00000000; // 1246 :   0 - 0x0
      13'h4DF: dout <= 8'b00000000; // 1247 :   0 - 0x0
      13'h4E0: dout <= 8'b00100100; // 1248 :  36 - 0x24 -- Sprite 0x4e
      13'h4E1: dout <= 8'b01010010; // 1249 :  82 - 0x52
      13'h4E2: dout <= 8'b01010010; // 1250 :  82 - 0x52
      13'h4E3: dout <= 8'b01010010; // 1251 :  82 - 0x52
      13'h4E4: dout <= 8'b01010010; // 1252 :  82 - 0x52
      13'h4E5: dout <= 8'b01010010; // 1253 :  82 - 0x52
      13'h4E6: dout <= 8'b01001100; // 1254 :  76 - 0x4c
      13'h4E7: dout <= 8'b00000000; // 1255 :   0 - 0x0
      13'h4E8: dout <= 8'b00000000; // 1256 :   0 - 0x0
      13'h4E9: dout <= 8'b00000000; // 1257 :   0 - 0x0
      13'h4EA: dout <= 8'b00000000; // 1258 :   0 - 0x0
      13'h4EB: dout <= 8'b00000000; // 1259 :   0 - 0x0
      13'h4EC: dout <= 8'b00000000; // 1260 :   0 - 0x0
      13'h4ED: dout <= 8'b00000000; // 1261 :   0 - 0x0
      13'h4EE: dout <= 8'b00000000; // 1262 :   0 - 0x0
      13'h4EF: dout <= 8'b00000000; // 1263 :   0 - 0x0
      13'h4F0: dout <= 8'b00111000; // 1264 :  56 - 0x38 -- Sprite 0x4f
      13'h4F1: dout <= 8'b01000100; // 1265 :  68 - 0x44
      13'h4F2: dout <= 8'b10000010; // 1266 : 130 - 0x82
      13'h4F3: dout <= 8'b10000010; // 1267 : 130 - 0x82
      13'h4F4: dout <= 8'b10000010; // 1268 : 130 - 0x82
      13'h4F5: dout <= 8'b01000100; // 1269 :  68 - 0x44
      13'h4F6: dout <= 8'b00111000; // 1270 :  56 - 0x38
      13'h4F7: dout <= 8'b00000000; // 1271 :   0 - 0x0
      13'h4F8: dout <= 8'b00000000; // 1272 :   0 - 0x0
      13'h4F9: dout <= 8'b00000000; // 1273 :   0 - 0x0
      13'h4FA: dout <= 8'b00000000; // 1274 :   0 - 0x0
      13'h4FB: dout <= 8'b00000000; // 1275 :   0 - 0x0
      13'h4FC: dout <= 8'b00000000; // 1276 :   0 - 0x0
      13'h4FD: dout <= 8'b00000000; // 1277 :   0 - 0x0
      13'h4FE: dout <= 8'b00000000; // 1278 :   0 - 0x0
      13'h4FF: dout <= 8'b00000000; // 1279 :   0 - 0x0
      13'h500: dout <= 8'b01111111; // 1280 : 127 - 0x7f -- Sprite 0x50
      13'h501: dout <= 8'b11000000; // 1281 : 192 - 0xc0
      13'h502: dout <= 8'b10000000; // 1282 : 128 - 0x80
      13'h503: dout <= 8'b10000000; // 1283 : 128 - 0x80
      13'h504: dout <= 8'b10000000; // 1284 : 128 - 0x80
      13'h505: dout <= 8'b11000011; // 1285 : 195 - 0xc3
      13'h506: dout <= 8'b11111111; // 1286 : 255 - 0xff
      13'h507: dout <= 8'b11111111; // 1287 : 255 - 0xff
      13'h508: dout <= 8'b00000000; // 1288 :   0 - 0x0
      13'h509: dout <= 8'b00111111; // 1289 :  63 - 0x3f
      13'h50A: dout <= 8'b01111111; // 1290 : 127 - 0x7f
      13'h50B: dout <= 8'b01111111; // 1291 : 127 - 0x7f
      13'h50C: dout <= 8'b01111111; // 1292 : 127 - 0x7f
      13'h50D: dout <= 8'b00111100; // 1293 :  60 - 0x3c
      13'h50E: dout <= 8'b00000000; // 1294 :   0 - 0x0
      13'h50F: dout <= 8'b01000000; // 1295 :  64 - 0x40
      13'h510: dout <= 8'b11111110; // 1296 : 254 - 0xfe -- Sprite 0x51
      13'h511: dout <= 8'b00000011; // 1297 :   3 - 0x3
      13'h512: dout <= 8'b00000001; // 1298 :   1 - 0x1
      13'h513: dout <= 8'b00000001; // 1299 :   1 - 0x1
      13'h514: dout <= 8'b00000001; // 1300 :   1 - 0x1
      13'h515: dout <= 8'b11000011; // 1301 : 195 - 0xc3
      13'h516: dout <= 8'b11111111; // 1302 : 255 - 0xff
      13'h517: dout <= 8'b11111111; // 1303 : 255 - 0xff
      13'h518: dout <= 8'b00000000; // 1304 :   0 - 0x0
      13'h519: dout <= 8'b11111100; // 1305 : 252 - 0xfc
      13'h51A: dout <= 8'b11111110; // 1306 : 254 - 0xfe
      13'h51B: dout <= 8'b11111110; // 1307 : 254 - 0xfe
      13'h51C: dout <= 8'b11111110; // 1308 : 254 - 0xfe
      13'h51D: dout <= 8'b00111100; // 1309 :  60 - 0x3c
      13'h51E: dout <= 8'b00000000; // 1310 :   0 - 0x0
      13'h51F: dout <= 8'b00000010; // 1311 :   2 - 0x2
      13'h520: dout <= 8'b00000000; // 1312 :   0 - 0x0 -- Sprite 0x52
      13'h521: dout <= 8'b00000111; // 1313 :   7 - 0x7
      13'h522: dout <= 8'b00001100; // 1314 :  12 - 0xc
      13'h523: dout <= 8'b00011000; // 1315 :  24 - 0x18
      13'h524: dout <= 8'b00110000; // 1316 :  48 - 0x30
      13'h525: dout <= 8'b01100000; // 1317 :  96 - 0x60
      13'h526: dout <= 8'b01000000; // 1318 :  64 - 0x40
      13'h527: dout <= 8'b01001111; // 1319 :  79 - 0x4f
      13'h528: dout <= 8'b00000000; // 1320 :   0 - 0x0
      13'h529: dout <= 8'b00000000; // 1321 :   0 - 0x0
      13'h52A: dout <= 8'b00000011; // 1322 :   3 - 0x3
      13'h52B: dout <= 8'b00000111; // 1323 :   7 - 0x7
      13'h52C: dout <= 8'b00001111; // 1324 :  15 - 0xf
      13'h52D: dout <= 8'b00011111; // 1325 :  31 - 0x1f
      13'h52E: dout <= 8'b00111111; // 1326 :  63 - 0x3f
      13'h52F: dout <= 8'b00110000; // 1327 :  48 - 0x30
      13'h530: dout <= 8'b00000000; // 1328 :   0 - 0x0 -- Sprite 0x53
      13'h531: dout <= 8'b11110000; // 1329 : 240 - 0xf0
      13'h532: dout <= 8'b01010000; // 1330 :  80 - 0x50
      13'h533: dout <= 8'b01001000; // 1331 :  72 - 0x48
      13'h534: dout <= 8'b01001100; // 1332 :  76 - 0x4c
      13'h535: dout <= 8'b01000100; // 1333 :  68 - 0x44
      13'h536: dout <= 8'b10000010; // 1334 : 130 - 0x82
      13'h537: dout <= 8'b10000011; // 1335 : 131 - 0x83
      13'h538: dout <= 8'b00000000; // 1336 :   0 - 0x0
      13'h539: dout <= 8'b00000000; // 1337 :   0 - 0x0
      13'h53A: dout <= 8'b10100000; // 1338 : 160 - 0xa0
      13'h53B: dout <= 8'b10110000; // 1339 : 176 - 0xb0
      13'h53C: dout <= 8'b10110000; // 1340 : 176 - 0xb0
      13'h53D: dout <= 8'b10111000; // 1341 : 184 - 0xb8
      13'h53E: dout <= 8'b01111100; // 1342 : 124 - 0x7c
      13'h53F: dout <= 8'b01111100; // 1343 : 124 - 0x7c
      13'h540: dout <= 8'b01111111; // 1344 : 127 - 0x7f -- Sprite 0x54
      13'h541: dout <= 8'b11011110; // 1345 : 222 - 0xde
      13'h542: dout <= 8'b10001110; // 1346 : 142 - 0x8e
      13'h543: dout <= 8'b11000101; // 1347 : 197 - 0xc5
      13'h544: dout <= 8'b10010010; // 1348 : 146 - 0x92
      13'h545: dout <= 8'b11000111; // 1349 : 199 - 0xc7
      13'h546: dout <= 8'b11100010; // 1350 : 226 - 0xe2
      13'h547: dout <= 8'b11010000; // 1351 : 208 - 0xd0
      13'h548: dout <= 8'b00000000; // 1352 :   0 - 0x0
      13'h549: dout <= 8'b00100001; // 1353 :  33 - 0x21
      13'h54A: dout <= 8'b01110001; // 1354 : 113 - 0x71
      13'h54B: dout <= 8'b00111010; // 1355 :  58 - 0x3a
      13'h54C: dout <= 8'b01101101; // 1356 : 109 - 0x6d
      13'h54D: dout <= 8'b00111000; // 1357 :  56 - 0x38
      13'h54E: dout <= 8'b00011101; // 1358 :  29 - 0x1d
      13'h54F: dout <= 8'b00101111; // 1359 :  47 - 0x2f
      13'h550: dout <= 8'b11111111; // 1360 : 255 - 0xff -- Sprite 0x55
      13'h551: dout <= 8'b11011110; // 1361 : 222 - 0xde
      13'h552: dout <= 8'b10001110; // 1362 : 142 - 0x8e
      13'h553: dout <= 8'b11000101; // 1363 : 197 - 0xc5
      13'h554: dout <= 8'b10010010; // 1364 : 146 - 0x92
      13'h555: dout <= 8'b01000111; // 1365 :  71 - 0x47
      13'h556: dout <= 8'b11100010; // 1366 : 226 - 0xe2
      13'h557: dout <= 8'b01010000; // 1367 :  80 - 0x50
      13'h558: dout <= 8'b00000000; // 1368 :   0 - 0x0
      13'h559: dout <= 8'b00100001; // 1369 :  33 - 0x21
      13'h55A: dout <= 8'b01110001; // 1370 : 113 - 0x71
      13'h55B: dout <= 8'b00111010; // 1371 :  58 - 0x3a
      13'h55C: dout <= 8'b01101101; // 1372 : 109 - 0x6d
      13'h55D: dout <= 8'b10111000; // 1373 : 184 - 0xb8
      13'h55E: dout <= 8'b00011101; // 1374 :  29 - 0x1d
      13'h55F: dout <= 8'b10101111; // 1375 : 175 - 0xaf
      13'h560: dout <= 8'b11111110; // 1376 : 254 - 0xfe -- Sprite 0x56
      13'h561: dout <= 8'b11011111; // 1377 : 223 - 0xdf
      13'h562: dout <= 8'b10001111; // 1378 : 143 - 0x8f
      13'h563: dout <= 8'b11000101; // 1379 : 197 - 0xc5
      13'h564: dout <= 8'b10010011; // 1380 : 147 - 0x93
      13'h565: dout <= 8'b01000111; // 1381 :  71 - 0x47
      13'h566: dout <= 8'b11100011; // 1382 : 227 - 0xe3
      13'h567: dout <= 8'b01010001; // 1383 :  81 - 0x51
      13'h568: dout <= 8'b00000000; // 1384 :   0 - 0x0
      13'h569: dout <= 8'b00100000; // 1385 :  32 - 0x20
      13'h56A: dout <= 8'b01110000; // 1386 : 112 - 0x70
      13'h56B: dout <= 8'b00111010; // 1387 :  58 - 0x3a
      13'h56C: dout <= 8'b01101100; // 1388 : 108 - 0x6c
      13'h56D: dout <= 8'b10111000; // 1389 : 184 - 0xb8
      13'h56E: dout <= 8'b00011100; // 1390 :  28 - 0x1c
      13'h56F: dout <= 8'b10101110; // 1391 : 174 - 0xae
      13'h570: dout <= 8'b01111111; // 1392 : 127 - 0x7f -- Sprite 0x57
      13'h571: dout <= 8'b10000000; // 1393 : 128 - 0x80
      13'h572: dout <= 8'b10110011; // 1394 : 179 - 0xb3
      13'h573: dout <= 8'b01001100; // 1395 :  76 - 0x4c
      13'h574: dout <= 8'b00111111; // 1396 :  63 - 0x3f
      13'h575: dout <= 8'b00000011; // 1397 :   3 - 0x3
      13'h576: dout <= 8'b00000000; // 1398 :   0 - 0x0
      13'h577: dout <= 8'b00000000; // 1399 :   0 - 0x0
      13'h578: dout <= 8'b00000000; // 1400 :   0 - 0x0
      13'h579: dout <= 8'b01111111; // 1401 : 127 - 0x7f
      13'h57A: dout <= 8'b01001100; // 1402 :  76 - 0x4c
      13'h57B: dout <= 8'b00110011; // 1403 :  51 - 0x33
      13'h57C: dout <= 8'b00000000; // 1404 :   0 - 0x0
      13'h57D: dout <= 8'b00000000; // 1405 :   0 - 0x0
      13'h57E: dout <= 8'b00000000; // 1406 :   0 - 0x0
      13'h57F: dout <= 8'b00000000; // 1407 :   0 - 0x0
      13'h580: dout <= 8'b11111111; // 1408 : 255 - 0xff -- Sprite 0x58
      13'h581: dout <= 8'b00000000; // 1409 :   0 - 0x0
      13'h582: dout <= 8'b00110011; // 1410 :  51 - 0x33
      13'h583: dout <= 8'b11001100; // 1411 : 204 - 0xcc
      13'h584: dout <= 8'b00110011; // 1412 :  51 - 0x33
      13'h585: dout <= 8'b11111111; // 1413 : 255 - 0xff
      13'h586: dout <= 8'b00000000; // 1414 :   0 - 0x0
      13'h587: dout <= 8'b00000000; // 1415 :   0 - 0x0
      13'h588: dout <= 8'b00000000; // 1416 :   0 - 0x0
      13'h589: dout <= 8'b11111111; // 1417 : 255 - 0xff
      13'h58A: dout <= 8'b11001100; // 1418 : 204 - 0xcc
      13'h58B: dout <= 8'b00110011; // 1419 :  51 - 0x33
      13'h58C: dout <= 8'b11001100; // 1420 : 204 - 0xcc
      13'h58D: dout <= 8'b00000000; // 1421 :   0 - 0x0
      13'h58E: dout <= 8'b00000000; // 1422 :   0 - 0x0
      13'h58F: dout <= 8'b00000000; // 1423 :   0 - 0x0
      13'h590: dout <= 8'b11111110; // 1424 : 254 - 0xfe -- Sprite 0x59
      13'h591: dout <= 8'b00000001; // 1425 :   1 - 0x1
      13'h592: dout <= 8'b00110011; // 1426 :  51 - 0x33
      13'h593: dout <= 8'b11001110; // 1427 : 206 - 0xce
      13'h594: dout <= 8'b00111100; // 1428 :  60 - 0x3c
      13'h595: dout <= 8'b11000000; // 1429 : 192 - 0xc0
      13'h596: dout <= 8'b00000000; // 1430 :   0 - 0x0
      13'h597: dout <= 8'b00000000; // 1431 :   0 - 0x0
      13'h598: dout <= 8'b00000000; // 1432 :   0 - 0x0
      13'h599: dout <= 8'b11111110; // 1433 : 254 - 0xfe
      13'h59A: dout <= 8'b11001100; // 1434 : 204 - 0xcc
      13'h59B: dout <= 8'b00110000; // 1435 :  48 - 0x30
      13'h59C: dout <= 8'b11000000; // 1436 : 192 - 0xc0
      13'h59D: dout <= 8'b00000000; // 1437 :   0 - 0x0
      13'h59E: dout <= 8'b00000000; // 1438 :   0 - 0x0
      13'h59F: dout <= 8'b00000000; // 1439 :   0 - 0x0
      13'h5A0: dout <= 8'b00000000; // 1440 :   0 - 0x0 -- Sprite 0x5a
      13'h5A1: dout <= 8'b00000000; // 1441 :   0 - 0x0
      13'h5A2: dout <= 8'b00000000; // 1442 :   0 - 0x0
      13'h5A3: dout <= 8'b00000000; // 1443 :   0 - 0x0
      13'h5A4: dout <= 8'b00000000; // 1444 :   0 - 0x0
      13'h5A5: dout <= 8'b00000000; // 1445 :   0 - 0x0
      13'h5A6: dout <= 8'b00000000; // 1446 :   0 - 0x0
      13'h5A7: dout <= 8'b00000000; // 1447 :   0 - 0x0
      13'h5A8: dout <= 8'b00000000; // 1448 :   0 - 0x0
      13'h5A9: dout <= 8'b00000000; // 1449 :   0 - 0x0
      13'h5AA: dout <= 8'b00000000; // 1450 :   0 - 0x0
      13'h5AB: dout <= 8'b00000000; // 1451 :   0 - 0x0
      13'h5AC: dout <= 8'b00000000; // 1452 :   0 - 0x0
      13'h5AD: dout <= 8'b00000000; // 1453 :   0 - 0x0
      13'h5AE: dout <= 8'b00000000; // 1454 :   0 - 0x0
      13'h5AF: dout <= 8'b00000000; // 1455 :   0 - 0x0
      13'h5B0: dout <= 8'b00000000; // 1456 :   0 - 0x0 -- Sprite 0x5b
      13'h5B1: dout <= 8'b00000000; // 1457 :   0 - 0x0
      13'h5B2: dout <= 8'b00000000; // 1458 :   0 - 0x0
      13'h5B3: dout <= 8'b00000001; // 1459 :   1 - 0x1
      13'h5B4: dout <= 8'b00000011; // 1460 :   3 - 0x3
      13'h5B5: dout <= 8'b00000011; // 1461 :   3 - 0x3
      13'h5B6: dout <= 8'b00000111; // 1462 :   7 - 0x7
      13'h5B7: dout <= 8'b00111111; // 1463 :  63 - 0x3f
      13'h5B8: dout <= 8'b00000000; // 1464 :   0 - 0x0
      13'h5B9: dout <= 8'b00000000; // 1465 :   0 - 0x0
      13'h5BA: dout <= 8'b00000000; // 1466 :   0 - 0x0
      13'h5BB: dout <= 8'b00000000; // 1467 :   0 - 0x0
      13'h5BC: dout <= 8'b00000001; // 1468 :   1 - 0x1
      13'h5BD: dout <= 8'b00000001; // 1469 :   1 - 0x1
      13'h5BE: dout <= 8'b00000011; // 1470 :   3 - 0x3
      13'h5BF: dout <= 8'b00000011; // 1471 :   3 - 0x3
      13'h5C0: dout <= 8'b00000000; // 1472 :   0 - 0x0 -- Sprite 0x5c
      13'h5C1: dout <= 8'b00000001; // 1473 :   1 - 0x1
      13'h5C2: dout <= 8'b01111111; // 1474 : 127 - 0x7f
      13'h5C3: dout <= 8'b11111111; // 1475 : 255 - 0xff
      13'h5C4: dout <= 8'b11111111; // 1476 : 255 - 0xff
      13'h5C5: dout <= 8'b11111111; // 1477 : 255 - 0xff
      13'h5C6: dout <= 8'b11111111; // 1478 : 255 - 0xff
      13'h5C7: dout <= 8'b11111111; // 1479 : 255 - 0xff
      13'h5C8: dout <= 8'b00000000; // 1480 :   0 - 0x0
      13'h5C9: dout <= 8'b00000000; // 1481 :   0 - 0x0
      13'h5CA: dout <= 8'b00000001; // 1482 :   1 - 0x1
      13'h5CB: dout <= 8'b01111110; // 1483 : 126 - 0x7e
      13'h5CC: dout <= 8'b11111111; // 1484 : 255 - 0xff
      13'h5CD: dout <= 8'b11111111; // 1485 : 255 - 0xff
      13'h5CE: dout <= 8'b11111111; // 1486 : 255 - 0xff
      13'h5CF: dout <= 8'b11111111; // 1487 : 255 - 0xff
      13'h5D0: dout <= 8'b11111111; // 1488 : 255 - 0xff -- Sprite 0x5d
      13'h5D1: dout <= 8'b11111111; // 1489 : 255 - 0xff
      13'h5D2: dout <= 8'b11111111; // 1490 : 255 - 0xff
      13'h5D3: dout <= 8'b11111111; // 1491 : 255 - 0xff
      13'h5D4: dout <= 8'b11111111; // 1492 : 255 - 0xff
      13'h5D5: dout <= 8'b11111111; // 1493 : 255 - 0xff
      13'h5D6: dout <= 8'b11111111; // 1494 : 255 - 0xff
      13'h5D7: dout <= 8'b11111111; // 1495 : 255 - 0xff
      13'h5D8: dout <= 8'b00000000; // 1496 :   0 - 0x0
      13'h5D9: dout <= 8'b11111111; // 1497 : 255 - 0xff
      13'h5DA: dout <= 8'b11111111; // 1498 : 255 - 0xff
      13'h5DB: dout <= 8'b11111111; // 1499 : 255 - 0xff
      13'h5DC: dout <= 8'b01111111; // 1500 : 127 - 0x7f
      13'h5DD: dout <= 8'b11111111; // 1501 : 255 - 0xff
      13'h5DE: dout <= 8'b11111111; // 1502 : 255 - 0xff
      13'h5DF: dout <= 8'b11111111; // 1503 : 255 - 0xff
      13'h5E0: dout <= 8'b00000000; // 1504 :   0 - 0x0 -- Sprite 0x5e
      13'h5E1: dout <= 8'b10000000; // 1505 : 128 - 0x80
      13'h5E2: dout <= 8'b11111110; // 1506 : 254 - 0xfe
      13'h5E3: dout <= 8'b11111111; // 1507 : 255 - 0xff
      13'h5E4: dout <= 8'b11111111; // 1508 : 255 - 0xff
      13'h5E5: dout <= 8'b11111111; // 1509 : 255 - 0xff
      13'h5E6: dout <= 8'b11111111; // 1510 : 255 - 0xff
      13'h5E7: dout <= 8'b11111111; // 1511 : 255 - 0xff
      13'h5E8: dout <= 8'b00000000; // 1512 :   0 - 0x0
      13'h5E9: dout <= 8'b00000000; // 1513 :   0 - 0x0
      13'h5EA: dout <= 8'b10000000; // 1514 : 128 - 0x80
      13'h5EB: dout <= 8'b01111110; // 1515 : 126 - 0x7e
      13'h5EC: dout <= 8'b10111111; // 1516 : 191 - 0xbf
      13'h5ED: dout <= 8'b11111111; // 1517 : 255 - 0xff
      13'h5EE: dout <= 8'b11111111; // 1518 : 255 - 0xff
      13'h5EF: dout <= 8'b11111111; // 1519 : 255 - 0xff
      13'h5F0: dout <= 8'b00000000; // 1520 :   0 - 0x0 -- Sprite 0x5f
      13'h5F1: dout <= 8'b00000000; // 1521 :   0 - 0x0
      13'h5F2: dout <= 8'b00000000; // 1522 :   0 - 0x0
      13'h5F3: dout <= 8'b10000000; // 1523 : 128 - 0x80
      13'h5F4: dout <= 8'b11000000; // 1524 : 192 - 0xc0
      13'h5F5: dout <= 8'b11000000; // 1525 : 192 - 0xc0
      13'h5F6: dout <= 8'b11100000; // 1526 : 224 - 0xe0
      13'h5F7: dout <= 8'b11111000; // 1527 : 248 - 0xf8
      13'h5F8: dout <= 8'b00000000; // 1528 :   0 - 0x0
      13'h5F9: dout <= 8'b00000000; // 1529 :   0 - 0x0
      13'h5FA: dout <= 8'b00000000; // 1530 :   0 - 0x0
      13'h5FB: dout <= 8'b00000000; // 1531 :   0 - 0x0
      13'h5FC: dout <= 8'b10000000; // 1532 : 128 - 0x80
      13'h5FD: dout <= 8'b10000000; // 1533 : 128 - 0x80
      13'h5FE: dout <= 8'b11000000; // 1534 : 192 - 0xc0
      13'h5FF: dout <= 8'b11000000; // 1535 : 192 - 0xc0
      13'h600: dout <= 8'b11111111; // 1536 : 255 - 0xff -- Sprite 0x60
      13'h601: dout <= 8'b11111111; // 1537 : 255 - 0xff
      13'h602: dout <= 8'b11111111; // 1538 : 255 - 0xff
      13'h603: dout <= 8'b11111111; // 1539 : 255 - 0xff
      13'h604: dout <= 8'b11111111; // 1540 : 255 - 0xff
      13'h605: dout <= 8'b11111111; // 1541 : 255 - 0xff
      13'h606: dout <= 8'b11111111; // 1542 : 255 - 0xff
      13'h607: dout <= 8'b11111111; // 1543 : 255 - 0xff
      13'h608: dout <= 8'b01111111; // 1544 : 127 - 0x7f
      13'h609: dout <= 8'b01111111; // 1545 : 127 - 0x7f
      13'h60A: dout <= 8'b01111101; // 1546 : 125 - 0x7d
      13'h60B: dout <= 8'b01111111; // 1547 : 127 - 0x7f
      13'h60C: dout <= 8'b00111111; // 1548 :  63 - 0x3f
      13'h60D: dout <= 8'b01111111; // 1549 : 127 - 0x7f
      13'h60E: dout <= 8'b01111111; // 1550 : 127 - 0x7f
      13'h60F: dout <= 8'b01110111; // 1551 : 119 - 0x77
      13'h610: dout <= 8'b11111111; // 1552 : 255 - 0xff -- Sprite 0x61
      13'h611: dout <= 8'b11111111; // 1553 : 255 - 0xff
      13'h612: dout <= 8'b11111111; // 1554 : 255 - 0xff
      13'h613: dout <= 8'b11111111; // 1555 : 255 - 0xff
      13'h614: dout <= 8'b11111111; // 1556 : 255 - 0xff
      13'h615: dout <= 8'b11111111; // 1557 : 255 - 0xff
      13'h616: dout <= 8'b11111111; // 1558 : 255 - 0xff
      13'h617: dout <= 8'b11111111; // 1559 : 255 - 0xff
      13'h618: dout <= 8'b11111110; // 1560 : 254 - 0xfe
      13'h619: dout <= 8'b11111110; // 1561 : 254 - 0xfe
      13'h61A: dout <= 8'b11111100; // 1562 : 252 - 0xfc
      13'h61B: dout <= 8'b11111110; // 1563 : 254 - 0xfe
      13'h61C: dout <= 8'b10111110; // 1564 : 190 - 0xbe
      13'h61D: dout <= 8'b11111110; // 1565 : 254 - 0xfe
      13'h61E: dout <= 8'b11111110; // 1566 : 254 - 0xfe
      13'h61F: dout <= 8'b11110110; // 1567 : 246 - 0xf6
      13'h620: dout <= 8'b01111000; // 1568 : 120 - 0x78 -- Sprite 0x62
      13'h621: dout <= 8'b01100000; // 1569 :  96 - 0x60
      13'h622: dout <= 8'b01000000; // 1570 :  64 - 0x40
      13'h623: dout <= 8'b01000000; // 1571 :  64 - 0x40
      13'h624: dout <= 8'b01000000; // 1572 :  64 - 0x40
      13'h625: dout <= 8'b01100000; // 1573 :  96 - 0x60
      13'h626: dout <= 8'b00110000; // 1574 :  48 - 0x30
      13'h627: dout <= 8'b00011111; // 1575 :  31 - 0x1f
      13'h628: dout <= 8'b00000111; // 1576 :   7 - 0x7
      13'h629: dout <= 8'b00011111; // 1577 :  31 - 0x1f
      13'h62A: dout <= 8'b00111111; // 1578 :  63 - 0x3f
      13'h62B: dout <= 8'b00111111; // 1579 :  63 - 0x3f
      13'h62C: dout <= 8'b00111111; // 1580 :  63 - 0x3f
      13'h62D: dout <= 8'b00011111; // 1581 :  31 - 0x1f
      13'h62E: dout <= 8'b00001111; // 1582 :  15 - 0xf
      13'h62F: dout <= 8'b00000000; // 1583 :   0 - 0x0
      13'h630: dout <= 8'b10000001; // 1584 : 129 - 0x81 -- Sprite 0x63
      13'h631: dout <= 8'b10000011; // 1585 : 131 - 0x83
      13'h632: dout <= 8'b11000001; // 1586 : 193 - 0xc1
      13'h633: dout <= 8'b01000011; // 1587 :  67 - 0x43
      13'h634: dout <= 8'b01000001; // 1588 :  65 - 0x41
      13'h635: dout <= 8'b01100011; // 1589 :  99 - 0x63
      13'h636: dout <= 8'b00100110; // 1590 :  38 - 0x26
      13'h637: dout <= 8'b11111000; // 1591 : 248 - 0xf8
      13'h638: dout <= 8'b01111110; // 1592 : 126 - 0x7e
      13'h639: dout <= 8'b01111100; // 1593 : 124 - 0x7c
      13'h63A: dout <= 8'b00111110; // 1594 :  62 - 0x3e
      13'h63B: dout <= 8'b10111100; // 1595 : 188 - 0xbc
      13'h63C: dout <= 8'b10111110; // 1596 : 190 - 0xbe
      13'h63D: dout <= 8'b10011100; // 1597 : 156 - 0x9c
      13'h63E: dout <= 8'b11011000; // 1598 : 216 - 0xd8
      13'h63F: dout <= 8'b00000000; // 1599 :   0 - 0x0
      13'h640: dout <= 8'b10111001; // 1600 : 185 - 0xb9 -- Sprite 0x64
      13'h641: dout <= 8'b10010100; // 1601 : 148 - 0x94
      13'h642: dout <= 8'b10001110; // 1602 : 142 - 0x8e
      13'h643: dout <= 8'b11000101; // 1603 : 197 - 0xc5
      13'h644: dout <= 8'b10010010; // 1604 : 146 - 0x92
      13'h645: dout <= 8'b11000111; // 1605 : 199 - 0xc7
      13'h646: dout <= 8'b11100010; // 1606 : 226 - 0xe2
      13'h647: dout <= 8'b11010000; // 1607 : 208 - 0xd0
      13'h648: dout <= 8'b01000110; // 1608 :  70 - 0x46
      13'h649: dout <= 8'b01101011; // 1609 : 107 - 0x6b
      13'h64A: dout <= 8'b01110001; // 1610 : 113 - 0x71
      13'h64B: dout <= 8'b00111010; // 1611 :  58 - 0x3a
      13'h64C: dout <= 8'b01101101; // 1612 : 109 - 0x6d
      13'h64D: dout <= 8'b00111000; // 1613 :  56 - 0x38
      13'h64E: dout <= 8'b00011101; // 1614 :  29 - 0x1d
      13'h64F: dout <= 8'b00101111; // 1615 :  47 - 0x2f
      13'h650: dout <= 8'b10111001; // 1616 : 185 - 0xb9 -- Sprite 0x65
      13'h651: dout <= 8'b00010100; // 1617 :  20 - 0x14
      13'h652: dout <= 8'b10001110; // 1618 : 142 - 0x8e
      13'h653: dout <= 8'b11000101; // 1619 : 197 - 0xc5
      13'h654: dout <= 8'b10010010; // 1620 : 146 - 0x92
      13'h655: dout <= 8'b01000111; // 1621 :  71 - 0x47
      13'h656: dout <= 8'b11100010; // 1622 : 226 - 0xe2
      13'h657: dout <= 8'b01010000; // 1623 :  80 - 0x50
      13'h658: dout <= 8'b01000110; // 1624 :  70 - 0x46
      13'h659: dout <= 8'b11101011; // 1625 : 235 - 0xeb
      13'h65A: dout <= 8'b01110001; // 1626 : 113 - 0x71
      13'h65B: dout <= 8'b00111010; // 1627 :  58 - 0x3a
      13'h65C: dout <= 8'b01101101; // 1628 : 109 - 0x6d
      13'h65D: dout <= 8'b10111000; // 1629 : 184 - 0xb8
      13'h65E: dout <= 8'b00011101; // 1630 :  29 - 0x1d
      13'h65F: dout <= 8'b10101111; // 1631 : 175 - 0xaf
      13'h660: dout <= 8'b10111001; // 1632 : 185 - 0xb9 -- Sprite 0x66
      13'h661: dout <= 8'b00010101; // 1633 :  21 - 0x15
      13'h662: dout <= 8'b10001111; // 1634 : 143 - 0x8f
      13'h663: dout <= 8'b11000101; // 1635 : 197 - 0xc5
      13'h664: dout <= 8'b10010011; // 1636 : 147 - 0x93
      13'h665: dout <= 8'b01000111; // 1637 :  71 - 0x47
      13'h666: dout <= 8'b11100011; // 1638 : 227 - 0xe3
      13'h667: dout <= 8'b01010001; // 1639 :  81 - 0x51
      13'h668: dout <= 8'b01000110; // 1640 :  70 - 0x46
      13'h669: dout <= 8'b11101010; // 1641 : 234 - 0xea
      13'h66A: dout <= 8'b01110000; // 1642 : 112 - 0x70
      13'h66B: dout <= 8'b00111010; // 1643 :  58 - 0x3a
      13'h66C: dout <= 8'b01101100; // 1644 : 108 - 0x6c
      13'h66D: dout <= 8'b10111000; // 1645 : 184 - 0xb8
      13'h66E: dout <= 8'b00011100; // 1646 :  28 - 0x1c
      13'h66F: dout <= 8'b10101110; // 1647 : 174 - 0xae
      13'h670: dout <= 8'b01111111; // 1648 : 127 - 0x7f -- Sprite 0x67
      13'h671: dout <= 8'b10000000; // 1649 : 128 - 0x80
      13'h672: dout <= 8'b11001100; // 1650 : 204 - 0xcc
      13'h673: dout <= 8'b01111111; // 1651 : 127 - 0x7f
      13'h674: dout <= 8'b00111111; // 1652 :  63 - 0x3f
      13'h675: dout <= 8'b00000011; // 1653 :   3 - 0x3
      13'h676: dout <= 8'b00000000; // 1654 :   0 - 0x0
      13'h677: dout <= 8'b00000000; // 1655 :   0 - 0x0
      13'h678: dout <= 8'b00000000; // 1656 :   0 - 0x0
      13'h679: dout <= 8'b01111111; // 1657 : 127 - 0x7f
      13'h67A: dout <= 8'b01111111; // 1658 : 127 - 0x7f
      13'h67B: dout <= 8'b00110011; // 1659 :  51 - 0x33
      13'h67C: dout <= 8'b00000000; // 1660 :   0 - 0x0
      13'h67D: dout <= 8'b00000000; // 1661 :   0 - 0x0
      13'h67E: dout <= 8'b00000000; // 1662 :   0 - 0x0
      13'h67F: dout <= 8'b00000000; // 1663 :   0 - 0x0
      13'h680: dout <= 8'b11111111; // 1664 : 255 - 0xff -- Sprite 0x68
      13'h681: dout <= 8'b00000000; // 1665 :   0 - 0x0
      13'h682: dout <= 8'b11001100; // 1666 : 204 - 0xcc
      13'h683: dout <= 8'b00110011; // 1667 :  51 - 0x33
      13'h684: dout <= 8'b11111111; // 1668 : 255 - 0xff
      13'h685: dout <= 8'b11111111; // 1669 : 255 - 0xff
      13'h686: dout <= 8'b00000000; // 1670 :   0 - 0x0
      13'h687: dout <= 8'b00000000; // 1671 :   0 - 0x0
      13'h688: dout <= 8'b00000000; // 1672 :   0 - 0x0
      13'h689: dout <= 8'b11111111; // 1673 : 255 - 0xff
      13'h68A: dout <= 8'b11111111; // 1674 : 255 - 0xff
      13'h68B: dout <= 8'b11111111; // 1675 : 255 - 0xff
      13'h68C: dout <= 8'b11001100; // 1676 : 204 - 0xcc
      13'h68D: dout <= 8'b00000000; // 1677 :   0 - 0x0
      13'h68E: dout <= 8'b00000000; // 1678 :   0 - 0x0
      13'h68F: dout <= 8'b00000000; // 1679 :   0 - 0x0
      13'h690: dout <= 8'b11111110; // 1680 : 254 - 0xfe -- Sprite 0x69
      13'h691: dout <= 8'b00000001; // 1681 :   1 - 0x1
      13'h692: dout <= 8'b11001101; // 1682 : 205 - 0xcd
      13'h693: dout <= 8'b00111110; // 1683 :  62 - 0x3e
      13'h694: dout <= 8'b11111100; // 1684 : 252 - 0xfc
      13'h695: dout <= 8'b11000000; // 1685 : 192 - 0xc0
      13'h696: dout <= 8'b00000000; // 1686 :   0 - 0x0
      13'h697: dout <= 8'b00000000; // 1687 :   0 - 0x0
      13'h698: dout <= 8'b00000000; // 1688 :   0 - 0x0
      13'h699: dout <= 8'b11111110; // 1689 : 254 - 0xfe
      13'h69A: dout <= 8'b11111110; // 1690 : 254 - 0xfe
      13'h69B: dout <= 8'b11110000; // 1691 : 240 - 0xf0
      13'h69C: dout <= 8'b11000000; // 1692 : 192 - 0xc0
      13'h69D: dout <= 8'b00000000; // 1693 :   0 - 0x0
      13'h69E: dout <= 8'b00000000; // 1694 :   0 - 0x0
      13'h69F: dout <= 8'b00000000; // 1695 :   0 - 0x0
      13'h6A0: dout <= 8'b00000000; // 1696 :   0 - 0x0 -- Sprite 0x6a
      13'h6A1: dout <= 8'b00000000; // 1697 :   0 - 0x0
      13'h6A2: dout <= 8'b00000000; // 1698 :   0 - 0x0
      13'h6A3: dout <= 8'b00000000; // 1699 :   0 - 0x0
      13'h6A4: dout <= 8'b00000000; // 1700 :   0 - 0x0
      13'h6A5: dout <= 8'b00000000; // 1701 :   0 - 0x0
      13'h6A6: dout <= 8'b00000000; // 1702 :   0 - 0x0
      13'h6A7: dout <= 8'b00000000; // 1703 :   0 - 0x0
      13'h6A8: dout <= 8'b00000000; // 1704 :   0 - 0x0
      13'h6A9: dout <= 8'b00000000; // 1705 :   0 - 0x0
      13'h6AA: dout <= 8'b00000000; // 1706 :   0 - 0x0
      13'h6AB: dout <= 8'b00000000; // 1707 :   0 - 0x0
      13'h6AC: dout <= 8'b00000000; // 1708 :   0 - 0x0
      13'h6AD: dout <= 8'b00000000; // 1709 :   0 - 0x0
      13'h6AE: dout <= 8'b00000000; // 1710 :   0 - 0x0
      13'h6AF: dout <= 8'b00000000; // 1711 :   0 - 0x0
      13'h6B0: dout <= 8'b01111111; // 1712 : 127 - 0x7f -- Sprite 0x6b
      13'h6B1: dout <= 8'b11111111; // 1713 : 255 - 0xff
      13'h6B2: dout <= 8'b11111111; // 1714 : 255 - 0xff
      13'h6B3: dout <= 8'b11111111; // 1715 : 255 - 0xff
      13'h6B4: dout <= 8'b01111111; // 1716 : 127 - 0x7f
      13'h6B5: dout <= 8'b00110000; // 1717 :  48 - 0x30
      13'h6B6: dout <= 8'b00001111; // 1718 :  15 - 0xf
      13'h6B7: dout <= 8'b00000000; // 1719 :   0 - 0x0
      13'h6B8: dout <= 8'b00111101; // 1720 :  61 - 0x3d
      13'h6B9: dout <= 8'b01111111; // 1721 : 127 - 0x7f
      13'h6BA: dout <= 8'b01111111; // 1722 : 127 - 0x7f
      13'h6BB: dout <= 8'b01111111; // 1723 : 127 - 0x7f
      13'h6BC: dout <= 8'b00111111; // 1724 :  63 - 0x3f
      13'h6BD: dout <= 8'b00001111; // 1725 :  15 - 0xf
      13'h6BE: dout <= 8'b00000000; // 1726 :   0 - 0x0
      13'h6BF: dout <= 8'b00000000; // 1727 :   0 - 0x0
      13'h6C0: dout <= 8'b11111111; // 1728 : 255 - 0xff -- Sprite 0x6c
      13'h6C1: dout <= 8'b11111111; // 1729 : 255 - 0xff
      13'h6C2: dout <= 8'b11111111; // 1730 : 255 - 0xff
      13'h6C3: dout <= 8'b11111111; // 1731 : 255 - 0xff
      13'h6C4: dout <= 8'b11111111; // 1732 : 255 - 0xff
      13'h6C5: dout <= 8'b11111110; // 1733 : 254 - 0xfe
      13'h6C6: dout <= 8'b00000001; // 1734 :   1 - 0x1
      13'h6C7: dout <= 8'b11111110; // 1735 : 254 - 0xfe
      13'h6C8: dout <= 8'b11111111; // 1736 : 255 - 0xff
      13'h6C9: dout <= 8'b11111111; // 1737 : 255 - 0xff
      13'h6CA: dout <= 8'b11111111; // 1738 : 255 - 0xff
      13'h6CB: dout <= 8'b11111111; // 1739 : 255 - 0xff
      13'h6CC: dout <= 8'b11111111; // 1740 : 255 - 0xff
      13'h6CD: dout <= 8'b11111111; // 1741 : 255 - 0xff
      13'h6CE: dout <= 8'b11111110; // 1742 : 254 - 0xfe
      13'h6CF: dout <= 8'b00000000; // 1743 :   0 - 0x0
      13'h6D0: dout <= 8'b00000000; // 1744 :   0 - 0x0 -- Sprite 0x6d
      13'h6D1: dout <= 8'b00000000; // 1745 :   0 - 0x0
      13'h6D2: dout <= 8'b00000000; // 1746 :   0 - 0x0
      13'h6D3: dout <= 8'b00000000; // 1747 :   0 - 0x0
      13'h6D4: dout <= 8'b00000000; // 1748 :   0 - 0x0
      13'h6D5: dout <= 8'b00000000; // 1749 :   0 - 0x0
      13'h6D6: dout <= 8'b00000000; // 1750 :   0 - 0x0
      13'h6D7: dout <= 8'b00000000; // 1751 :   0 - 0x0
      13'h6D8: dout <= 8'b00000000; // 1752 :   0 - 0x0
      13'h6D9: dout <= 8'b00000000; // 1753 :   0 - 0x0
      13'h6DA: dout <= 8'b00000000; // 1754 :   0 - 0x0
      13'h6DB: dout <= 8'b00000000; // 1755 :   0 - 0x0
      13'h6DC: dout <= 8'b00000000; // 1756 :   0 - 0x0
      13'h6DD: dout <= 8'b00000000; // 1757 :   0 - 0x0
      13'h6DE: dout <= 8'b00000000; // 1758 :   0 - 0x0
      13'h6DF: dout <= 8'b00000000; // 1759 :   0 - 0x0
      13'h6E0: dout <= 8'b00000000; // 1760 :   0 - 0x0 -- Sprite 0x6e
      13'h6E1: dout <= 8'b00000000; // 1761 :   0 - 0x0
      13'h6E2: dout <= 8'b00000000; // 1762 :   0 - 0x0
      13'h6E3: dout <= 8'b00000000; // 1763 :   0 - 0x0
      13'h6E4: dout <= 8'b00000000; // 1764 :   0 - 0x0
      13'h6E5: dout <= 8'b00000000; // 1765 :   0 - 0x0
      13'h6E6: dout <= 8'b00000000; // 1766 :   0 - 0x0
      13'h6E7: dout <= 8'b00000000; // 1767 :   0 - 0x0
      13'h6E8: dout <= 8'b00000000; // 1768 :   0 - 0x0
      13'h6E9: dout <= 8'b00000000; // 1769 :   0 - 0x0
      13'h6EA: dout <= 8'b00000000; // 1770 :   0 - 0x0
      13'h6EB: dout <= 8'b00000000; // 1771 :   0 - 0x0
      13'h6EC: dout <= 8'b00000000; // 1772 :   0 - 0x0
      13'h6ED: dout <= 8'b00000000; // 1773 :   0 - 0x0
      13'h6EE: dout <= 8'b00000000; // 1774 :   0 - 0x0
      13'h6EF: dout <= 8'b00000000; // 1775 :   0 - 0x0
      13'h6F0: dout <= 8'b11111100; // 1776 : 252 - 0xfc -- Sprite 0x6f
      13'h6F1: dout <= 8'b11111110; // 1777 : 254 - 0xfe
      13'h6F2: dout <= 8'b11111111; // 1778 : 255 - 0xff
      13'h6F3: dout <= 8'b11111111; // 1779 : 255 - 0xff
      13'h6F4: dout <= 8'b11110010; // 1780 : 242 - 0xf2
      13'h6F5: dout <= 8'b00001100; // 1781 :  12 - 0xc
      13'h6F6: dout <= 8'b11110000; // 1782 : 240 - 0xf0
      13'h6F7: dout <= 8'b00000000; // 1783 :   0 - 0x0
      13'h6F8: dout <= 8'b10111000; // 1784 : 184 - 0xb8
      13'h6F9: dout <= 8'b11111100; // 1785 : 252 - 0xfc
      13'h6FA: dout <= 8'b11111110; // 1786 : 254 - 0xfe
      13'h6FB: dout <= 8'b11111110; // 1787 : 254 - 0xfe
      13'h6FC: dout <= 8'b11111100; // 1788 : 252 - 0xfc
      13'h6FD: dout <= 8'b11110000; // 1789 : 240 - 0xf0
      13'h6FE: dout <= 8'b00000000; // 1790 :   0 - 0x0
      13'h6FF: dout <= 8'b00000000; // 1791 :   0 - 0x0
      13'h700: dout <= 8'b01111111; // 1792 : 127 - 0x7f -- Sprite 0x70
      13'h701: dout <= 8'b11000000; // 1793 : 192 - 0xc0
      13'h702: dout <= 8'b10000000; // 1794 : 128 - 0x80
      13'h703: dout <= 8'b10000000; // 1795 : 128 - 0x80
      13'h704: dout <= 8'b11100011; // 1796 : 227 - 0xe3
      13'h705: dout <= 8'b11111111; // 1797 : 255 - 0xff
      13'h706: dout <= 8'b11111111; // 1798 : 255 - 0xff
      13'h707: dout <= 8'b11111111; // 1799 : 255 - 0xff
      13'h708: dout <= 8'b00000000; // 1800 :   0 - 0x0
      13'h709: dout <= 8'b00111111; // 1801 :  63 - 0x3f
      13'h70A: dout <= 8'b01111111; // 1802 : 127 - 0x7f
      13'h70B: dout <= 8'b01111111; // 1803 : 127 - 0x7f
      13'h70C: dout <= 8'b00011100; // 1804 :  28 - 0x1c
      13'h70D: dout <= 8'b00000000; // 1805 :   0 - 0x0
      13'h70E: dout <= 8'b00000000; // 1806 :   0 - 0x0
      13'h70F: dout <= 8'b00000000; // 1807 :   0 - 0x0
      13'h710: dout <= 8'b11111111; // 1808 : 255 - 0xff -- Sprite 0x71
      13'h711: dout <= 8'b00000000; // 1809 :   0 - 0x0
      13'h712: dout <= 8'b00000000; // 1810 :   0 - 0x0
      13'h713: dout <= 8'b00000000; // 1811 :   0 - 0x0
      13'h714: dout <= 8'b00000000; // 1812 :   0 - 0x0
      13'h715: dout <= 8'b11000011; // 1813 : 195 - 0xc3
      13'h716: dout <= 8'b11111111; // 1814 : 255 - 0xff
      13'h717: dout <= 8'b11111111; // 1815 : 255 - 0xff
      13'h718: dout <= 8'b00000000; // 1816 :   0 - 0x0
      13'h719: dout <= 8'b11111111; // 1817 : 255 - 0xff
      13'h71A: dout <= 8'b11111111; // 1818 : 255 - 0xff
      13'h71B: dout <= 8'b11111111; // 1819 : 255 - 0xff
      13'h71C: dout <= 8'b11111111; // 1820 : 255 - 0xff
      13'h71D: dout <= 8'b00111100; // 1821 :  60 - 0x3c
      13'h71E: dout <= 8'b00000000; // 1822 :   0 - 0x0
      13'h71F: dout <= 8'b00000000; // 1823 :   0 - 0x0
      13'h720: dout <= 8'b11111110; // 1824 : 254 - 0xfe -- Sprite 0x72
      13'h721: dout <= 8'b00000011; // 1825 :   3 - 0x3
      13'h722: dout <= 8'b00000001; // 1826 :   1 - 0x1
      13'h723: dout <= 8'b00000001; // 1827 :   1 - 0x1
      13'h724: dout <= 8'b11000111; // 1828 : 199 - 0xc7
      13'h725: dout <= 8'b11111111; // 1829 : 255 - 0xff
      13'h726: dout <= 8'b11111111; // 1830 : 255 - 0xff
      13'h727: dout <= 8'b11111111; // 1831 : 255 - 0xff
      13'h728: dout <= 8'b00000000; // 1832 :   0 - 0x0
      13'h729: dout <= 8'b11111100; // 1833 : 252 - 0xfc
      13'h72A: dout <= 8'b11111110; // 1834 : 254 - 0xfe
      13'h72B: dout <= 8'b11111110; // 1835 : 254 - 0xfe
      13'h72C: dout <= 8'b00111000; // 1836 :  56 - 0x38
      13'h72D: dout <= 8'b00000000; // 1837 :   0 - 0x0
      13'h72E: dout <= 8'b00000000; // 1838 :   0 - 0x0
      13'h72F: dout <= 8'b00000000; // 1839 :   0 - 0x0
      13'h730: dout <= 8'b11111111; // 1840 : 255 - 0xff -- Sprite 0x73
      13'h731: dout <= 8'b11111111; // 1841 : 255 - 0xff
      13'h732: dout <= 8'b11111111; // 1842 : 255 - 0xff
      13'h733: dout <= 8'b11111111; // 1843 : 255 - 0xff
      13'h734: dout <= 8'b11111111; // 1844 : 255 - 0xff
      13'h735: dout <= 8'b11111111; // 1845 : 255 - 0xff
      13'h736: dout <= 8'b11111111; // 1846 : 255 - 0xff
      13'h737: dout <= 8'b11111111; // 1847 : 255 - 0xff
      13'h738: dout <= 8'b11111111; // 1848 : 255 - 0xff
      13'h739: dout <= 8'b11111111; // 1849 : 255 - 0xff
      13'h73A: dout <= 8'b11111101; // 1850 : 253 - 0xfd
      13'h73B: dout <= 8'b11111111; // 1851 : 255 - 0xff
      13'h73C: dout <= 8'b10111111; // 1852 : 191 - 0xbf
      13'h73D: dout <= 8'b11111111; // 1853 : 255 - 0xff
      13'h73E: dout <= 8'b11111111; // 1854 : 255 - 0xff
      13'h73F: dout <= 8'b11110111; // 1855 : 247 - 0xf7
      13'h740: dout <= 8'b10111001; // 1856 : 185 - 0xb9 -- Sprite 0x74
      13'h741: dout <= 8'b10010100; // 1857 : 148 - 0x94
      13'h742: dout <= 8'b10001110; // 1858 : 142 - 0x8e
      13'h743: dout <= 8'b11000101; // 1859 : 197 - 0xc5
      13'h744: dout <= 8'b10010010; // 1860 : 146 - 0x92
      13'h745: dout <= 8'b11000111; // 1861 : 199 - 0xc7
      13'h746: dout <= 8'b11100010; // 1862 : 226 - 0xe2
      13'h747: dout <= 8'b01111111; // 1863 : 127 - 0x7f
      13'h748: dout <= 8'b01000110; // 1864 :  70 - 0x46
      13'h749: dout <= 8'b01101011; // 1865 : 107 - 0x6b
      13'h74A: dout <= 8'b01110001; // 1866 : 113 - 0x71
      13'h74B: dout <= 8'b00111010; // 1867 :  58 - 0x3a
      13'h74C: dout <= 8'b01101101; // 1868 : 109 - 0x6d
      13'h74D: dout <= 8'b00111000; // 1869 :  56 - 0x38
      13'h74E: dout <= 8'b00011101; // 1870 :  29 - 0x1d
      13'h74F: dout <= 8'b00000000; // 1871 :   0 - 0x0
      13'h750: dout <= 8'b10111001; // 1872 : 185 - 0xb9 -- Sprite 0x75
      13'h751: dout <= 8'b00010100; // 1873 :  20 - 0x14
      13'h752: dout <= 8'b10001110; // 1874 : 142 - 0x8e
      13'h753: dout <= 8'b11000101; // 1875 : 197 - 0xc5
      13'h754: dout <= 8'b10010010; // 1876 : 146 - 0x92
      13'h755: dout <= 8'b01000111; // 1877 :  71 - 0x47
      13'h756: dout <= 8'b11100010; // 1878 : 226 - 0xe2
      13'h757: dout <= 8'b11111111; // 1879 : 255 - 0xff
      13'h758: dout <= 8'b01000110; // 1880 :  70 - 0x46
      13'h759: dout <= 8'b11101011; // 1881 : 235 - 0xeb
      13'h75A: dout <= 8'b01110001; // 1882 : 113 - 0x71
      13'h75B: dout <= 8'b00111010; // 1883 :  58 - 0x3a
      13'h75C: dout <= 8'b01101101; // 1884 : 109 - 0x6d
      13'h75D: dout <= 8'b10111000; // 1885 : 184 - 0xb8
      13'h75E: dout <= 8'b00011101; // 1886 :  29 - 0x1d
      13'h75F: dout <= 8'b00000000; // 1887 :   0 - 0x0
      13'h760: dout <= 8'b10111001; // 1888 : 185 - 0xb9 -- Sprite 0x76
      13'h761: dout <= 8'b00010101; // 1889 :  21 - 0x15
      13'h762: dout <= 8'b10001111; // 1890 : 143 - 0x8f
      13'h763: dout <= 8'b11000101; // 1891 : 197 - 0xc5
      13'h764: dout <= 8'b10010011; // 1892 : 147 - 0x93
      13'h765: dout <= 8'b01000111; // 1893 :  71 - 0x47
      13'h766: dout <= 8'b11100011; // 1894 : 227 - 0xe3
      13'h767: dout <= 8'b11111110; // 1895 : 254 - 0xfe
      13'h768: dout <= 8'b01000110; // 1896 :  70 - 0x46
      13'h769: dout <= 8'b11101010; // 1897 : 234 - 0xea
      13'h76A: dout <= 8'b01110000; // 1898 : 112 - 0x70
      13'h76B: dout <= 8'b00111010; // 1899 :  58 - 0x3a
      13'h76C: dout <= 8'b01101100; // 1900 : 108 - 0x6c
      13'h76D: dout <= 8'b10111000; // 1901 : 184 - 0xb8
      13'h76E: dout <= 8'b00011100; // 1902 :  28 - 0x1c
      13'h76F: dout <= 8'b00000000; // 1903 :   0 - 0x0
      13'h770: dout <= 8'b11111111; // 1904 : 255 - 0xff -- Sprite 0x77
      13'h771: dout <= 8'b11111111; // 1905 : 255 - 0xff
      13'h772: dout <= 8'b11111111; // 1906 : 255 - 0xff
      13'h773: dout <= 8'b11111111; // 1907 : 255 - 0xff
      13'h774: dout <= 8'b11111111; // 1908 : 255 - 0xff
      13'h775: dout <= 8'b11111111; // 1909 : 255 - 0xff
      13'h776: dout <= 8'b11111111; // 1910 : 255 - 0xff
      13'h777: dout <= 8'b11111111; // 1911 : 255 - 0xff
      13'h778: dout <= 8'b10000001; // 1912 : 129 - 0x81
      13'h779: dout <= 8'b11111111; // 1913 : 255 - 0xff
      13'h77A: dout <= 8'b11111101; // 1914 : 253 - 0xfd
      13'h77B: dout <= 8'b11111111; // 1915 : 255 - 0xff
      13'h77C: dout <= 8'b10111111; // 1916 : 191 - 0xbf
      13'h77D: dout <= 8'b11111111; // 1917 : 255 - 0xff
      13'h77E: dout <= 8'b11111111; // 1918 : 255 - 0xff
      13'h77F: dout <= 8'b11110111; // 1919 : 247 - 0xf7
      13'h780: dout <= 8'b00000000; // 1920 :   0 - 0x0 -- Sprite 0x78
      13'h781: dout <= 8'b00000000; // 1921 :   0 - 0x0
      13'h782: dout <= 8'b00000000; // 1922 :   0 - 0x0
      13'h783: dout <= 8'b00000000; // 1923 :   0 - 0x0
      13'h784: dout <= 8'b00000000; // 1924 :   0 - 0x0
      13'h785: dout <= 8'b00000000; // 1925 :   0 - 0x0
      13'h786: dout <= 8'b00000000; // 1926 :   0 - 0x0
      13'h787: dout <= 8'b00000000; // 1927 :   0 - 0x0
      13'h788: dout <= 8'b00000000; // 1928 :   0 - 0x0
      13'h789: dout <= 8'b00000000; // 1929 :   0 - 0x0
      13'h78A: dout <= 8'b00000000; // 1930 :   0 - 0x0
      13'h78B: dout <= 8'b00000000; // 1931 :   0 - 0x0
      13'h78C: dout <= 8'b00000000; // 1932 :   0 - 0x0
      13'h78D: dout <= 8'b00000000; // 1933 :   0 - 0x0
      13'h78E: dout <= 8'b00000000; // 1934 :   0 - 0x0
      13'h78F: dout <= 8'b00000000; // 1935 :   0 - 0x0
      13'h790: dout <= 8'b00000000; // 1936 :   0 - 0x0 -- Sprite 0x79
      13'h791: dout <= 8'b00000000; // 1937 :   0 - 0x0
      13'h792: dout <= 8'b00000000; // 1938 :   0 - 0x0
      13'h793: dout <= 8'b00000000; // 1939 :   0 - 0x0
      13'h794: dout <= 8'b00000000; // 1940 :   0 - 0x0
      13'h795: dout <= 8'b00000000; // 1941 :   0 - 0x0
      13'h796: dout <= 8'b00000000; // 1942 :   0 - 0x0
      13'h797: dout <= 8'b00000000; // 1943 :   0 - 0x0
      13'h798: dout <= 8'b00000000; // 1944 :   0 - 0x0
      13'h799: dout <= 8'b00000000; // 1945 :   0 - 0x0
      13'h79A: dout <= 8'b00000000; // 1946 :   0 - 0x0
      13'h79B: dout <= 8'b00000000; // 1947 :   0 - 0x0
      13'h79C: dout <= 8'b00000000; // 1948 :   0 - 0x0
      13'h79D: dout <= 8'b00000000; // 1949 :   0 - 0x0
      13'h79E: dout <= 8'b00000000; // 1950 :   0 - 0x0
      13'h79F: dout <= 8'b00000000; // 1951 :   0 - 0x0
      13'h7A0: dout <= 8'b00000000; // 1952 :   0 - 0x0 -- Sprite 0x7a
      13'h7A1: dout <= 8'b00000000; // 1953 :   0 - 0x0
      13'h7A2: dout <= 8'b00000000; // 1954 :   0 - 0x0
      13'h7A3: dout <= 8'b00000000; // 1955 :   0 - 0x0
      13'h7A4: dout <= 8'b00000000; // 1956 :   0 - 0x0
      13'h7A5: dout <= 8'b00000000; // 1957 :   0 - 0x0
      13'h7A6: dout <= 8'b00000000; // 1958 :   0 - 0x0
      13'h7A7: dout <= 8'b00000000; // 1959 :   0 - 0x0
      13'h7A8: dout <= 8'b00000000; // 1960 :   0 - 0x0
      13'h7A9: dout <= 8'b00000000; // 1961 :   0 - 0x0
      13'h7AA: dout <= 8'b00000000; // 1962 :   0 - 0x0
      13'h7AB: dout <= 8'b00000000; // 1963 :   0 - 0x0
      13'h7AC: dout <= 8'b00000000; // 1964 :   0 - 0x0
      13'h7AD: dout <= 8'b00000000; // 1965 :   0 - 0x0
      13'h7AE: dout <= 8'b00000000; // 1966 :   0 - 0x0
      13'h7AF: dout <= 8'b00000000; // 1967 :   0 - 0x0
      13'h7B0: dout <= 8'b00000000; // 1968 :   0 - 0x0 -- Sprite 0x7b
      13'h7B1: dout <= 8'b00000000; // 1969 :   0 - 0x0
      13'h7B2: dout <= 8'b00000000; // 1970 :   0 - 0x0
      13'h7B3: dout <= 8'b00000000; // 1971 :   0 - 0x0
      13'h7B4: dout <= 8'b00000000; // 1972 :   0 - 0x0
      13'h7B5: dout <= 8'b00000000; // 1973 :   0 - 0x0
      13'h7B6: dout <= 8'b00000000; // 1974 :   0 - 0x0
      13'h7B7: dout <= 8'b00000000; // 1975 :   0 - 0x0
      13'h7B8: dout <= 8'b00000000; // 1976 :   0 - 0x0
      13'h7B9: dout <= 8'b00000000; // 1977 :   0 - 0x0
      13'h7BA: dout <= 8'b00000000; // 1978 :   0 - 0x0
      13'h7BB: dout <= 8'b00000000; // 1979 :   0 - 0x0
      13'h7BC: dout <= 8'b00000000; // 1980 :   0 - 0x0
      13'h7BD: dout <= 8'b00000000; // 1981 :   0 - 0x0
      13'h7BE: dout <= 8'b00000000; // 1982 :   0 - 0x0
      13'h7BF: dout <= 8'b00000000; // 1983 :   0 - 0x0
      13'h7C0: dout <= 8'b00100010; // 1984 :  34 - 0x22 -- Sprite 0x7c
      13'h7C1: dout <= 8'b01010101; // 1985 :  85 - 0x55
      13'h7C2: dout <= 8'b10101010; // 1986 : 170 - 0xaa
      13'h7C3: dout <= 8'b00000101; // 1987 :   5 - 0x5
      13'h7C4: dout <= 8'b00000100; // 1988 :   4 - 0x4
      13'h7C5: dout <= 8'b00001010; // 1989 :  10 - 0xa
      13'h7C6: dout <= 8'b01010000; // 1990 :  80 - 0x50
      13'h7C7: dout <= 8'b00000010; // 1991 :   2 - 0x2
      13'h7C8: dout <= 8'b00000000; // 1992 :   0 - 0x0
      13'h7C9: dout <= 8'b00100010; // 1993 :  34 - 0x22
      13'h7CA: dout <= 8'b01110111; // 1994 : 119 - 0x77
      13'h7CB: dout <= 8'b11111111; // 1995 : 255 - 0xff
      13'h7CC: dout <= 8'b11111011; // 1996 : 251 - 0xfb
      13'h7CD: dout <= 8'b11110101; // 1997 : 245 - 0xf5
      13'h7CE: dout <= 8'b11101111; // 1998 : 239 - 0xef
      13'h7CF: dout <= 8'b11111111; // 1999 : 255 - 0xff
      13'h7D0: dout <= 8'b01110011; // 2000 : 115 - 0x73 -- Sprite 0x7d
      13'h7D1: dout <= 8'b11111111; // 2001 : 255 - 0xff
      13'h7D2: dout <= 8'b11111111; // 2002 : 255 - 0xff
      13'h7D3: dout <= 8'b10111101; // 2003 : 189 - 0xbd
      13'h7D4: dout <= 8'b01101110; // 2004 : 110 - 0x6e
      13'h7D5: dout <= 8'b00001010; // 2005 :  10 - 0xa
      13'h7D6: dout <= 8'b01010000; // 2006 :  80 - 0x50
      13'h7D7: dout <= 8'b00000010; // 2007 :   2 - 0x2
      13'h7D8: dout <= 8'b00000000; // 2008 :   0 - 0x0
      13'h7D9: dout <= 8'b01110011; // 2009 : 115 - 0x73
      13'h7DA: dout <= 8'b11111111; // 2010 : 255 - 0xff
      13'h7DB: dout <= 8'b11111111; // 2011 : 255 - 0xff
      13'h7DC: dout <= 8'b11111011; // 2012 : 251 - 0xfb
      13'h7DD: dout <= 8'b11111101; // 2013 : 253 - 0xfd
      13'h7DE: dout <= 8'b11101111; // 2014 : 239 - 0xef
      13'h7DF: dout <= 8'b11111111; // 2015 : 255 - 0xff
      13'h7E0: dout <= 8'b00100000; // 2016 :  32 - 0x20 -- Sprite 0x7e
      13'h7E1: dout <= 8'b01010000; // 2017 :  80 - 0x50
      13'h7E2: dout <= 8'b10000100; // 2018 : 132 - 0x84
      13'h7E3: dout <= 8'b00000000; // 2019 :   0 - 0x0
      13'h7E4: dout <= 8'b00100100; // 2020 :  36 - 0x24
      13'h7E5: dout <= 8'b01011010; // 2021 :  90 - 0x5a
      13'h7E6: dout <= 8'b00010000; // 2022 :  16 - 0x10
      13'h7E7: dout <= 8'b00000000; // 2023 :   0 - 0x0
      13'h7E8: dout <= 8'b11011111; // 2024 : 223 - 0xdf
      13'h7E9: dout <= 8'b10101111; // 2025 : 175 - 0xaf
      13'h7EA: dout <= 8'b01111111; // 2026 : 127 - 0x7f
      13'h7EB: dout <= 8'b11111111; // 2027 : 255 - 0xff
      13'h7EC: dout <= 8'b11111011; // 2028 : 251 - 0xfb
      13'h7ED: dout <= 8'b11110101; // 2029 : 245 - 0xf5
      13'h7EE: dout <= 8'b11101111; // 2030 : 239 - 0xef
      13'h7EF: dout <= 8'b11111111; // 2031 : 255 - 0xff
      13'h7F0: dout <= 8'b11111111; // 2032 : 255 - 0xff -- Sprite 0x7f
      13'h7F1: dout <= 8'b01010000; // 2033 :  80 - 0x50
      13'h7F2: dout <= 8'b10000100; // 2034 : 132 - 0x84
      13'h7F3: dout <= 8'b00000000; // 2035 :   0 - 0x0
      13'h7F4: dout <= 8'b00100100; // 2036 :  36 - 0x24
      13'h7F5: dout <= 8'b01011010; // 2037 :  90 - 0x5a
      13'h7F6: dout <= 8'b00010000; // 2038 :  16 - 0x10
      13'h7F7: dout <= 8'b00000000; // 2039 :   0 - 0x0
      13'h7F8: dout <= 8'b00000000; // 2040 :   0 - 0x0
      13'h7F9: dout <= 8'b10101111; // 2041 : 175 - 0xaf
      13'h7FA: dout <= 8'b01111111; // 2042 : 127 - 0x7f
      13'h7FB: dout <= 8'b11111111; // 2043 : 255 - 0xff
      13'h7FC: dout <= 8'b11111011; // 2044 : 251 - 0xfb
      13'h7FD: dout <= 8'b11110101; // 2045 : 245 - 0xf5
      13'h7FE: dout <= 8'b11101111; // 2046 : 239 - 0xef
      13'h7FF: dout <= 8'b11111111; // 2047 : 255 - 0xff
      13'h800: dout <= 8'b11111111; // 2048 : 255 - 0xff -- Sprite 0x80
      13'h801: dout <= 8'b10000000; // 2049 : 128 - 0x80
      13'h802: dout <= 8'b11001111; // 2050 : 207 - 0xcf
      13'h803: dout <= 8'b01001000; // 2051 :  72 - 0x48
      13'h804: dout <= 8'b11001111; // 2052 : 207 - 0xcf
      13'h805: dout <= 8'b10000000; // 2053 : 128 - 0x80
      13'h806: dout <= 8'b11001111; // 2054 : 207 - 0xcf
      13'h807: dout <= 8'b01001000; // 2055 :  72 - 0x48
      13'h808: dout <= 8'b00000000; // 2056 :   0 - 0x0
      13'h809: dout <= 8'b01111111; // 2057 : 127 - 0x7f
      13'h80A: dout <= 8'b00110000; // 2058 :  48 - 0x30
      13'h80B: dout <= 8'b00110000; // 2059 :  48 - 0x30
      13'h80C: dout <= 8'b00110000; // 2060 :  48 - 0x30
      13'h80D: dout <= 8'b01111111; // 2061 : 127 - 0x7f
      13'h80E: dout <= 8'b00110000; // 2062 :  48 - 0x30
      13'h80F: dout <= 8'b00110000; // 2063 :  48 - 0x30
      13'h810: dout <= 8'b11111111; // 2064 : 255 - 0xff -- Sprite 0x81
      13'h811: dout <= 8'b10000000; // 2065 : 128 - 0x80
      13'h812: dout <= 8'b11111111; // 2066 : 255 - 0xff
      13'h813: dout <= 8'b10000000; // 2067 : 128 - 0x80
      13'h814: dout <= 8'b10000000; // 2068 : 128 - 0x80
      13'h815: dout <= 8'b11011111; // 2069 : 223 - 0xdf
      13'h816: dout <= 8'b10110000; // 2070 : 176 - 0xb0
      13'h817: dout <= 8'b11000000; // 2071 : 192 - 0xc0
      13'h818: dout <= 8'b00000000; // 2072 :   0 - 0x0
      13'h819: dout <= 8'b01111111; // 2073 : 127 - 0x7f
      13'h81A: dout <= 8'b00000000; // 2074 :   0 - 0x0
      13'h81B: dout <= 8'b01111111; // 2075 : 127 - 0x7f
      13'h81C: dout <= 8'b01111111; // 2076 : 127 - 0x7f
      13'h81D: dout <= 8'b00100000; // 2077 :  32 - 0x20
      13'h81E: dout <= 8'b01000000; // 2078 :  64 - 0x40
      13'h81F: dout <= 8'b00000000; // 2079 :   0 - 0x0
      13'h820: dout <= 8'b11111111; // 2080 : 255 - 0xff -- Sprite 0x82
      13'h821: dout <= 8'b00000001; // 2081 :   1 - 0x1
      13'h822: dout <= 8'b11110011; // 2082 : 243 - 0xf3
      13'h823: dout <= 8'b00010010; // 2083 :  18 - 0x12
      13'h824: dout <= 8'b11110011; // 2084 : 243 - 0xf3
      13'h825: dout <= 8'b00000001; // 2085 :   1 - 0x1
      13'h826: dout <= 8'b11110011; // 2086 : 243 - 0xf3
      13'h827: dout <= 8'b00010010; // 2087 :  18 - 0x12
      13'h828: dout <= 8'b00000000; // 2088 :   0 - 0x0
      13'h829: dout <= 8'b11111110; // 2089 : 254 - 0xfe
      13'h82A: dout <= 8'b00001100; // 2090 :  12 - 0xc
      13'h82B: dout <= 8'b00001100; // 2091 :  12 - 0xc
      13'h82C: dout <= 8'b00001100; // 2092 :  12 - 0xc
      13'h82D: dout <= 8'b11111110; // 2093 : 254 - 0xfe
      13'h82E: dout <= 8'b00001100; // 2094 :  12 - 0xc
      13'h82F: dout <= 8'b00001100; // 2095 :  12 - 0xc
      13'h830: dout <= 8'b11111111; // 2096 : 255 - 0xff -- Sprite 0x83
      13'h831: dout <= 8'b00000000; // 2097 :   0 - 0x0
      13'h832: dout <= 8'b11111111; // 2098 : 255 - 0xff
      13'h833: dout <= 8'b00000000; // 2099 :   0 - 0x0
      13'h834: dout <= 8'b00000000; // 2100 :   0 - 0x0
      13'h835: dout <= 8'b11111111; // 2101 : 255 - 0xff
      13'h836: dout <= 8'b00000000; // 2102 :   0 - 0x0
      13'h837: dout <= 8'b00000000; // 2103 :   0 - 0x0
      13'h838: dout <= 8'b00000000; // 2104 :   0 - 0x0
      13'h839: dout <= 8'b11111111; // 2105 : 255 - 0xff
      13'h83A: dout <= 8'b00000000; // 2106 :   0 - 0x0
      13'h83B: dout <= 8'b11111111; // 2107 : 255 - 0xff
      13'h83C: dout <= 8'b11111111; // 2108 : 255 - 0xff
      13'h83D: dout <= 8'b00000000; // 2109 :   0 - 0x0
      13'h83E: dout <= 8'b00000000; // 2110 :   0 - 0x0
      13'h83F: dout <= 8'b00000000; // 2111 :   0 - 0x0
      13'h840: dout <= 8'b11111111; // 2112 : 255 - 0xff -- Sprite 0x84
      13'h841: dout <= 8'b10000010; // 2113 : 130 - 0x82
      13'h842: dout <= 8'b00010000; // 2114 :  16 - 0x10
      13'h843: dout <= 8'b00000000; // 2115 :   0 - 0x0
      13'h844: dout <= 8'b00000000; // 2116 :   0 - 0x0
      13'h845: dout <= 8'b00010000; // 2117 :  16 - 0x10
      13'h846: dout <= 8'b01000100; // 2118 :  68 - 0x44
      13'h847: dout <= 8'b11111111; // 2119 : 255 - 0xff
      13'h848: dout <= 8'b00000000; // 2120 :   0 - 0x0
      13'h849: dout <= 8'b11111111; // 2121 : 255 - 0xff
      13'h84A: dout <= 8'b11111111; // 2122 : 255 - 0xff
      13'h84B: dout <= 8'b11111111; // 2123 : 255 - 0xff
      13'h84C: dout <= 8'b11111111; // 2124 : 255 - 0xff
      13'h84D: dout <= 8'b11101111; // 2125 : 239 - 0xef
      13'h84E: dout <= 8'b10111011; // 2126 : 187 - 0xbb
      13'h84F: dout <= 8'b00000000; // 2127 :   0 - 0x0
      13'h850: dout <= 8'b11111111; // 2128 : 255 - 0xff -- Sprite 0x85
      13'h851: dout <= 8'b00000001; // 2129 :   1 - 0x1
      13'h852: dout <= 8'b11111111; // 2130 : 255 - 0xff
      13'h853: dout <= 8'b00000001; // 2131 :   1 - 0x1
      13'h854: dout <= 8'b00000001; // 2132 :   1 - 0x1
      13'h855: dout <= 8'b11110011; // 2133 : 243 - 0xf3
      13'h856: dout <= 8'b00001101; // 2134 :  13 - 0xd
      13'h857: dout <= 8'b00000011; // 2135 :   3 - 0x3
      13'h858: dout <= 8'b00000000; // 2136 :   0 - 0x0
      13'h859: dout <= 8'b11111110; // 2137 : 254 - 0xfe
      13'h85A: dout <= 8'b00000000; // 2138 :   0 - 0x0
      13'h85B: dout <= 8'b11111110; // 2139 : 254 - 0xfe
      13'h85C: dout <= 8'b11111110; // 2140 : 254 - 0xfe
      13'h85D: dout <= 8'b00001100; // 2141 :  12 - 0xc
      13'h85E: dout <= 8'b00000010; // 2142 :   2 - 0x2
      13'h85F: dout <= 8'b00000000; // 2143 :   0 - 0x0
      13'h860: dout <= 8'b00000000; // 2144 :   0 - 0x0 -- Sprite 0x86
      13'h861: dout <= 8'b00000000; // 2145 :   0 - 0x0
      13'h862: dout <= 8'b00000000; // 2146 :   0 - 0x0
      13'h863: dout <= 8'b00000000; // 2147 :   0 - 0x0
      13'h864: dout <= 8'b00000000; // 2148 :   0 - 0x0
      13'h865: dout <= 8'b00000000; // 2149 :   0 - 0x0
      13'h866: dout <= 8'b00000000; // 2150 :   0 - 0x0
      13'h867: dout <= 8'b00000000; // 2151 :   0 - 0x0
      13'h868: dout <= 8'b00000000; // 2152 :   0 - 0x0
      13'h869: dout <= 8'b00000000; // 2153 :   0 - 0x0
      13'h86A: dout <= 8'b00000000; // 2154 :   0 - 0x0
      13'h86B: dout <= 8'b00000000; // 2155 :   0 - 0x0
      13'h86C: dout <= 8'b00000000; // 2156 :   0 - 0x0
      13'h86D: dout <= 8'b00000000; // 2157 :   0 - 0x0
      13'h86E: dout <= 8'b00000000; // 2158 :   0 - 0x0
      13'h86F: dout <= 8'b00000000; // 2159 :   0 - 0x0
      13'h870: dout <= 8'b00000000; // 2160 :   0 - 0x0 -- Sprite 0x87
      13'h871: dout <= 8'b00000000; // 2161 :   0 - 0x0
      13'h872: dout <= 8'b00000000; // 2162 :   0 - 0x0
      13'h873: dout <= 8'b00000000; // 2163 :   0 - 0x0
      13'h874: dout <= 8'b00000000; // 2164 :   0 - 0x0
      13'h875: dout <= 8'b00000000; // 2165 :   0 - 0x0
      13'h876: dout <= 8'b00000000; // 2166 :   0 - 0x0
      13'h877: dout <= 8'b00000000; // 2167 :   0 - 0x0
      13'h878: dout <= 8'b00000000; // 2168 :   0 - 0x0
      13'h879: dout <= 8'b00000000; // 2169 :   0 - 0x0
      13'h87A: dout <= 8'b00000000; // 2170 :   0 - 0x0
      13'h87B: dout <= 8'b00000000; // 2171 :   0 - 0x0
      13'h87C: dout <= 8'b00000000; // 2172 :   0 - 0x0
      13'h87D: dout <= 8'b00000000; // 2173 :   0 - 0x0
      13'h87E: dout <= 8'b00000000; // 2174 :   0 - 0x0
      13'h87F: dout <= 8'b00000000; // 2175 :   0 - 0x0
      13'h880: dout <= 8'b00000111; // 2176 :   7 - 0x7 -- Sprite 0x88
      13'h881: dout <= 8'b00011110; // 2177 :  30 - 0x1e
      13'h882: dout <= 8'b00101111; // 2178 :  47 - 0x2f
      13'h883: dout <= 8'b01010011; // 2179 :  83 - 0x53
      13'h884: dout <= 8'b01101110; // 2180 : 110 - 0x6e
      13'h885: dout <= 8'b11011011; // 2181 : 219 - 0xdb
      13'h886: dout <= 8'b11111010; // 2182 : 250 - 0xfa
      13'h887: dout <= 8'b11010101; // 2183 : 213 - 0xd5
      13'h888: dout <= 8'b00000000; // 2184 :   0 - 0x0
      13'h889: dout <= 8'b00000111; // 2185 :   7 - 0x7
      13'h88A: dout <= 8'b00011111; // 2186 :  31 - 0x1f
      13'h88B: dout <= 8'b00111100; // 2187 :  60 - 0x3c
      13'h88C: dout <= 8'b00110001; // 2188 :  49 - 0x31
      13'h88D: dout <= 8'b01110100; // 2189 : 116 - 0x74
      13'h88E: dout <= 8'b01100101; // 2190 : 101 - 0x65
      13'h88F: dout <= 8'b01101010; // 2191 : 106 - 0x6a
      13'h890: dout <= 8'b10111011; // 2192 : 187 - 0xbb -- Sprite 0x89
      13'h891: dout <= 8'b11110010; // 2193 : 242 - 0xf2
      13'h892: dout <= 8'b11011101; // 2194 : 221 - 0xdd
      13'h893: dout <= 8'b01001111; // 2195 :  79 - 0x4f
      13'h894: dout <= 8'b01111011; // 2196 : 123 - 0x7b
      13'h895: dout <= 8'b00110010; // 2197 :  50 - 0x32
      13'h896: dout <= 8'b00011111; // 2198 :  31 - 0x1f
      13'h897: dout <= 8'b00000111; // 2199 :   7 - 0x7
      13'h898: dout <= 8'b01100100; // 2200 : 100 - 0x64
      13'h899: dout <= 8'b01101101; // 2201 : 109 - 0x6d
      13'h89A: dout <= 8'b01110010; // 2202 : 114 - 0x72
      13'h89B: dout <= 8'b00110000; // 2203 :  48 - 0x30
      13'h89C: dout <= 8'b00111100; // 2204 :  60 - 0x3c
      13'h89D: dout <= 8'b00011111; // 2205 :  31 - 0x1f
      13'h89E: dout <= 8'b00000111; // 2206 :   7 - 0x7
      13'h89F: dout <= 8'b00000000; // 2207 :   0 - 0x0
      13'h8A0: dout <= 8'b11100000; // 2208 : 224 - 0xe0 -- Sprite 0x8a
      13'h8A1: dout <= 8'b11011000; // 2209 : 216 - 0xd8
      13'h8A2: dout <= 8'b01010100; // 2210 :  84 - 0x54
      13'h8A3: dout <= 8'b11101010; // 2211 : 234 - 0xea
      13'h8A4: dout <= 8'b10111010; // 2212 : 186 - 0xba
      13'h8A5: dout <= 8'b10010011; // 2213 : 147 - 0x93
      13'h8A6: dout <= 8'b11011111; // 2214 : 223 - 0xdf
      13'h8A7: dout <= 8'b10111101; // 2215 : 189 - 0xbd
      13'h8A8: dout <= 8'b00000000; // 2216 :   0 - 0x0
      13'h8A9: dout <= 8'b11100000; // 2217 : 224 - 0xe0
      13'h8AA: dout <= 8'b11111000; // 2218 : 248 - 0xf8
      13'h8AB: dout <= 8'b00111100; // 2219 :  60 - 0x3c
      13'h8AC: dout <= 8'b01001100; // 2220 :  76 - 0x4c
      13'h8AD: dout <= 8'b01101110; // 2221 : 110 - 0x6e
      13'h8AE: dout <= 8'b00100110; // 2222 :  38 - 0x26
      13'h8AF: dout <= 8'b01000110; // 2223 :  70 - 0x46
      13'h8B0: dout <= 8'b01101011; // 2224 : 107 - 0x6b -- Sprite 0x8b
      13'h8B1: dout <= 8'b10011111; // 2225 : 159 - 0x9f
      13'h8B2: dout <= 8'b01011101; // 2226 :  93 - 0x5d
      13'h8B3: dout <= 8'b10110110; // 2227 : 182 - 0xb6
      13'h8B4: dout <= 8'b11101010; // 2228 : 234 - 0xea
      13'h8B5: dout <= 8'b11001100; // 2229 : 204 - 0xcc
      13'h8B6: dout <= 8'b01111000; // 2230 : 120 - 0x78
      13'h8B7: dout <= 8'b11100000; // 2231 : 224 - 0xe0
      13'h8B8: dout <= 8'b10010110; // 2232 : 150 - 0x96
      13'h8B9: dout <= 8'b01100110; // 2233 : 102 - 0x66
      13'h8BA: dout <= 8'b10101110; // 2234 : 174 - 0xae
      13'h8BB: dout <= 8'b01001100; // 2235 :  76 - 0x4c
      13'h8BC: dout <= 8'b00111100; // 2236 :  60 - 0x3c
      13'h8BD: dout <= 8'b11111000; // 2237 : 248 - 0xf8
      13'h8BE: dout <= 8'b11100000; // 2238 : 224 - 0xe0
      13'h8BF: dout <= 8'b00000000; // 2239 :   0 - 0x0
      13'h8C0: dout <= 8'b00000111; // 2240 :   7 - 0x7 -- Sprite 0x8c
      13'h8C1: dout <= 8'b00011000; // 2241 :  24 - 0x18
      13'h8C2: dout <= 8'b00100011; // 2242 :  35 - 0x23
      13'h8C3: dout <= 8'b01001100; // 2243 :  76 - 0x4c
      13'h8C4: dout <= 8'b01110000; // 2244 : 112 - 0x70
      13'h8C5: dout <= 8'b10100001; // 2245 : 161 - 0xa1
      13'h8C6: dout <= 8'b10100110; // 2246 : 166 - 0xa6
      13'h8C7: dout <= 8'b10101000; // 2247 : 168 - 0xa8
      13'h8C8: dout <= 8'b00000000; // 2248 :   0 - 0x0
      13'h8C9: dout <= 8'b00000111; // 2249 :   7 - 0x7
      13'h8CA: dout <= 8'b00011111; // 2250 :  31 - 0x1f
      13'h8CB: dout <= 8'b00111111; // 2251 :  63 - 0x3f
      13'h8CC: dout <= 8'b00111111; // 2252 :  63 - 0x3f
      13'h8CD: dout <= 8'b01111111; // 2253 : 127 - 0x7f
      13'h8CE: dout <= 8'b01111111; // 2254 : 127 - 0x7f
      13'h8CF: dout <= 8'b01111111; // 2255 : 127 - 0x7f
      13'h8D0: dout <= 8'b10100101; // 2256 : 165 - 0xa5 -- Sprite 0x8d
      13'h8D1: dout <= 8'b10100010; // 2257 : 162 - 0xa2
      13'h8D2: dout <= 8'b10010000; // 2258 : 144 - 0x90
      13'h8D3: dout <= 8'b01001000; // 2259 :  72 - 0x48
      13'h8D4: dout <= 8'b01000111; // 2260 :  71 - 0x47
      13'h8D5: dout <= 8'b00100000; // 2261 :  32 - 0x20
      13'h8D6: dout <= 8'b00011001; // 2262 :  25 - 0x19
      13'h8D7: dout <= 8'b00000111; // 2263 :   7 - 0x7
      13'h8D8: dout <= 8'b01111111; // 2264 : 127 - 0x7f
      13'h8D9: dout <= 8'b01111111; // 2265 : 127 - 0x7f
      13'h8DA: dout <= 8'b01111111; // 2266 : 127 - 0x7f
      13'h8DB: dout <= 8'b00111111; // 2267 :  63 - 0x3f
      13'h8DC: dout <= 8'b00111111; // 2268 :  63 - 0x3f
      13'h8DD: dout <= 8'b00011111; // 2269 :  31 - 0x1f
      13'h8DE: dout <= 8'b00000111; // 2270 :   7 - 0x7
      13'h8DF: dout <= 8'b00000000; // 2271 :   0 - 0x0
      13'h8E0: dout <= 8'b11100000; // 2272 : 224 - 0xe0 -- Sprite 0x8e
      13'h8E1: dout <= 8'b00011000; // 2273 :  24 - 0x18
      13'h8E2: dout <= 8'b00000100; // 2274 :   4 - 0x4
      13'h8E3: dout <= 8'b11000010; // 2275 : 194 - 0xc2
      13'h8E4: dout <= 8'b00110010; // 2276 :  50 - 0x32
      13'h8E5: dout <= 8'b00001001; // 2277 :   9 - 0x9
      13'h8E6: dout <= 8'b11000101; // 2278 : 197 - 0xc5
      13'h8E7: dout <= 8'b00100101; // 2279 :  37 - 0x25
      13'h8E8: dout <= 8'b00000000; // 2280 :   0 - 0x0
      13'h8E9: dout <= 8'b11100000; // 2281 : 224 - 0xe0
      13'h8EA: dout <= 8'b11111000; // 2282 : 248 - 0xf8
      13'h8EB: dout <= 8'b11111100; // 2283 : 252 - 0xfc
      13'h8EC: dout <= 8'b11111100; // 2284 : 252 - 0xfc
      13'h8ED: dout <= 8'b11111110; // 2285 : 254 - 0xfe
      13'h8EE: dout <= 8'b11111110; // 2286 : 254 - 0xfe
      13'h8EF: dout <= 8'b11111110; // 2287 : 254 - 0xfe
      13'h8F0: dout <= 8'b10100101; // 2288 : 165 - 0xa5 -- Sprite 0x8f
      13'h8F1: dout <= 8'b01100101; // 2289 : 101 - 0x65
      13'h8F2: dout <= 8'b01000101; // 2290 :  69 - 0x45
      13'h8F3: dout <= 8'b10001010; // 2291 : 138 - 0x8a
      13'h8F4: dout <= 8'b10010010; // 2292 : 146 - 0x92
      13'h8F5: dout <= 8'b00100100; // 2293 :  36 - 0x24
      13'h8F6: dout <= 8'b11011000; // 2294 : 216 - 0xd8
      13'h8F7: dout <= 8'b11100000; // 2295 : 224 - 0xe0
      13'h8F8: dout <= 8'b11111110; // 2296 : 254 - 0xfe
      13'h8F9: dout <= 8'b11111110; // 2297 : 254 - 0xfe
      13'h8FA: dout <= 8'b11111110; // 2298 : 254 - 0xfe
      13'h8FB: dout <= 8'b11111100; // 2299 : 252 - 0xfc
      13'h8FC: dout <= 8'b11111100; // 2300 : 252 - 0xfc
      13'h8FD: dout <= 8'b11111000; // 2301 : 248 - 0xf8
      13'h8FE: dout <= 8'b11100000; // 2302 : 224 - 0xe0
      13'h8FF: dout <= 8'b00000000; // 2303 :   0 - 0x0
      13'h900: dout <= 8'b00000000; // 2304 :   0 - 0x0 -- Sprite 0x90
      13'h901: dout <= 8'b00000000; // 2305 :   0 - 0x0
      13'h902: dout <= 8'b00100000; // 2306 :  32 - 0x20
      13'h903: dout <= 8'b00110000; // 2307 :  48 - 0x30
      13'h904: dout <= 8'b00101100; // 2308 :  44 - 0x2c
      13'h905: dout <= 8'b00100010; // 2309 :  34 - 0x22
      13'h906: dout <= 8'b00010001; // 2310 :  17 - 0x11
      13'h907: dout <= 8'b00001000; // 2311 :   8 - 0x8
      13'h908: dout <= 8'b00000000; // 2312 :   0 - 0x0
      13'h909: dout <= 8'b00000000; // 2313 :   0 - 0x0
      13'h90A: dout <= 8'b00000000; // 2314 :   0 - 0x0
      13'h90B: dout <= 8'b00000000; // 2315 :   0 - 0x0
      13'h90C: dout <= 8'b00010000; // 2316 :  16 - 0x10
      13'h90D: dout <= 8'b00011100; // 2317 :  28 - 0x1c
      13'h90E: dout <= 8'b00001110; // 2318 :  14 - 0xe
      13'h90F: dout <= 8'b00000111; // 2319 :   7 - 0x7
      13'h910: dout <= 8'b00000100; // 2320 :   4 - 0x4 -- Sprite 0x91
      13'h911: dout <= 8'b11110010; // 2321 : 242 - 0xf2
      13'h912: dout <= 8'b11001111; // 2322 : 207 - 0xcf
      13'h913: dout <= 8'b00110000; // 2323 :  48 - 0x30
      13'h914: dout <= 8'b00001100; // 2324 :  12 - 0xc
      13'h915: dout <= 8'b11111111; // 2325 : 255 - 0xff
      13'h916: dout <= 8'b10000000; // 2326 : 128 - 0x80
      13'h917: dout <= 8'b11111111; // 2327 : 255 - 0xff
      13'h918: dout <= 8'b00000011; // 2328 :   3 - 0x3
      13'h919: dout <= 8'b00000001; // 2329 :   1 - 0x1
      13'h91A: dout <= 8'b00110000; // 2330 :  48 - 0x30
      13'h91B: dout <= 8'b00001111; // 2331 :  15 - 0xf
      13'h91C: dout <= 8'b00000011; // 2332 :   3 - 0x3
      13'h91D: dout <= 8'b00000000; // 2333 :   0 - 0x0
      13'h91E: dout <= 8'b01111111; // 2334 : 127 - 0x7f
      13'h91F: dout <= 8'b00000000; // 2335 :   0 - 0x0
      13'h920: dout <= 8'b01000010; // 2336 :  66 - 0x42 -- Sprite 0x92
      13'h921: dout <= 8'b10100101; // 2337 : 165 - 0xa5
      13'h922: dout <= 8'b10100101; // 2338 : 165 - 0xa5
      13'h923: dout <= 8'b10011001; // 2339 : 153 - 0x99
      13'h924: dout <= 8'b10011001; // 2340 : 153 - 0x99
      13'h925: dout <= 8'b10011001; // 2341 : 153 - 0x99
      13'h926: dout <= 8'b00000001; // 2342 :   1 - 0x1
      13'h927: dout <= 8'b00000000; // 2343 :   0 - 0x0
      13'h928: dout <= 8'b00000000; // 2344 :   0 - 0x0
      13'h929: dout <= 8'b01000010; // 2345 :  66 - 0x42
      13'h92A: dout <= 8'b01000010; // 2346 :  66 - 0x42
      13'h92B: dout <= 8'b01100110; // 2347 : 102 - 0x66
      13'h92C: dout <= 8'b01100110; // 2348 : 102 - 0x66
      13'h92D: dout <= 8'b01100110; // 2349 : 102 - 0x66
      13'h92E: dout <= 8'b11111110; // 2350 : 254 - 0xfe
      13'h92F: dout <= 8'b11111111; // 2351 : 255 - 0xff
      13'h930: dout <= 8'b11111111; // 2352 : 255 - 0xff -- Sprite 0x93
      13'h931: dout <= 8'b11111111; // 2353 : 255 - 0xff
      13'h932: dout <= 8'b11111111; // 2354 : 255 - 0xff
      13'h933: dout <= 8'b10000001; // 2355 : 129 - 0x81
      13'h934: dout <= 8'b11111111; // 2356 : 255 - 0xff
      13'h935: dout <= 8'b11111111; // 2357 : 255 - 0xff
      13'h936: dout <= 8'b11111111; // 2358 : 255 - 0xff
      13'h937: dout <= 8'b10000001; // 2359 : 129 - 0x81
      13'h938: dout <= 8'b01111110; // 2360 : 126 - 0x7e
      13'h939: dout <= 8'b01111110; // 2361 : 126 - 0x7e
      13'h93A: dout <= 8'b01111110; // 2362 : 126 - 0x7e
      13'h93B: dout <= 8'b01111110; // 2363 : 126 - 0x7e
      13'h93C: dout <= 8'b01111110; // 2364 : 126 - 0x7e
      13'h93D: dout <= 8'b01111110; // 2365 : 126 - 0x7e
      13'h93E: dout <= 8'b01111110; // 2366 : 126 - 0x7e
      13'h93F: dout <= 8'b01111110; // 2367 : 126 - 0x7e
      13'h940: dout <= 8'b00000000; // 2368 :   0 - 0x0 -- Sprite 0x94
      13'h941: dout <= 8'b00000000; // 2369 :   0 - 0x0
      13'h942: dout <= 8'b00000100; // 2370 :   4 - 0x4
      13'h943: dout <= 8'b00001100; // 2371 :  12 - 0xc
      13'h944: dout <= 8'b00110100; // 2372 :  52 - 0x34
      13'h945: dout <= 8'b01000100; // 2373 :  68 - 0x44
      13'h946: dout <= 8'b10001000; // 2374 : 136 - 0x88
      13'h947: dout <= 8'b00010000; // 2375 :  16 - 0x10
      13'h948: dout <= 8'b00000000; // 2376 :   0 - 0x0
      13'h949: dout <= 8'b00000000; // 2377 :   0 - 0x0
      13'h94A: dout <= 8'b00000000; // 2378 :   0 - 0x0
      13'h94B: dout <= 8'b00000000; // 2379 :   0 - 0x0
      13'h94C: dout <= 8'b00001000; // 2380 :   8 - 0x8
      13'h94D: dout <= 8'b00111000; // 2381 :  56 - 0x38
      13'h94E: dout <= 8'b01110000; // 2382 : 112 - 0x70
      13'h94F: dout <= 8'b11100000; // 2383 : 224 - 0xe0
      13'h950: dout <= 8'b00100000; // 2384 :  32 - 0x20 -- Sprite 0x95
      13'h951: dout <= 8'b01001111; // 2385 :  79 - 0x4f
      13'h952: dout <= 8'b11110011; // 2386 : 243 - 0xf3
      13'h953: dout <= 8'b00001100; // 2387 :  12 - 0xc
      13'h954: dout <= 8'b00110000; // 2388 :  48 - 0x30
      13'h955: dout <= 8'b11111111; // 2389 : 255 - 0xff
      13'h956: dout <= 8'b00000001; // 2390 :   1 - 0x1
      13'h957: dout <= 8'b11111111; // 2391 : 255 - 0xff
      13'h958: dout <= 8'b11000000; // 2392 : 192 - 0xc0
      13'h959: dout <= 8'b10000000; // 2393 : 128 - 0x80
      13'h95A: dout <= 8'b00001100; // 2394 :  12 - 0xc
      13'h95B: dout <= 8'b11110000; // 2395 : 240 - 0xf0
      13'h95C: dout <= 8'b11000000; // 2396 : 192 - 0xc0
      13'h95D: dout <= 8'b00000000; // 2397 :   0 - 0x0
      13'h95E: dout <= 8'b11111110; // 2398 : 254 - 0xfe
      13'h95F: dout <= 8'b00000000; // 2399 :   0 - 0x0
      13'h960: dout <= 8'b01111111; // 2400 : 127 - 0x7f -- Sprite 0x96
      13'h961: dout <= 8'b11111111; // 2401 : 255 - 0xff
      13'h962: dout <= 8'b11111111; // 2402 : 255 - 0xff
      13'h963: dout <= 8'b11111111; // 2403 : 255 - 0xff
      13'h964: dout <= 8'b11111011; // 2404 : 251 - 0xfb
      13'h965: dout <= 8'b11111111; // 2405 : 255 - 0xff
      13'h966: dout <= 8'b11111111; // 2406 : 255 - 0xff
      13'h967: dout <= 8'b11111111; // 2407 : 255 - 0xff
      13'h968: dout <= 8'b00000000; // 2408 :   0 - 0x0
      13'h969: dout <= 8'b00111111; // 2409 :  63 - 0x3f
      13'h96A: dout <= 8'b01111111; // 2410 : 127 - 0x7f
      13'h96B: dout <= 8'b01111111; // 2411 : 127 - 0x7f
      13'h96C: dout <= 8'b01111111; // 2412 : 127 - 0x7f
      13'h96D: dout <= 8'b01111111; // 2413 : 127 - 0x7f
      13'h96E: dout <= 8'b01111111; // 2414 : 127 - 0x7f
      13'h96F: dout <= 8'b01111111; // 2415 : 127 - 0x7f
      13'h970: dout <= 8'b11111111; // 2416 : 255 - 0xff -- Sprite 0x97
      13'h971: dout <= 8'b11111111; // 2417 : 255 - 0xff
      13'h972: dout <= 8'b11111111; // 2418 : 255 - 0xff
      13'h973: dout <= 8'b11111111; // 2419 : 255 - 0xff
      13'h974: dout <= 8'b11111111; // 2420 : 255 - 0xff
      13'h975: dout <= 8'b11111111; // 2421 : 255 - 0xff
      13'h976: dout <= 8'b11111110; // 2422 : 254 - 0xfe
      13'h977: dout <= 8'b11111111; // 2423 : 255 - 0xff
      13'h978: dout <= 8'b01111111; // 2424 : 127 - 0x7f
      13'h979: dout <= 8'b01111111; // 2425 : 127 - 0x7f
      13'h97A: dout <= 8'b00111111; // 2426 :  63 - 0x3f
      13'h97B: dout <= 8'b01111111; // 2427 : 127 - 0x7f
      13'h97C: dout <= 8'b01111111; // 2428 : 127 - 0x7f
      13'h97D: dout <= 8'b01111111; // 2429 : 127 - 0x7f
      13'h97E: dout <= 8'b01111111; // 2430 : 127 - 0x7f
      13'h97F: dout <= 8'b01111111; // 2431 : 127 - 0x7f
      13'h980: dout <= 8'b11111111; // 2432 : 255 - 0xff -- Sprite 0x98
      13'h981: dout <= 8'b10111111; // 2433 : 191 - 0xbf
      13'h982: dout <= 8'b11111111; // 2434 : 255 - 0xff
      13'h983: dout <= 8'b11111111; // 2435 : 255 - 0xff
      13'h984: dout <= 8'b11111011; // 2436 : 251 - 0xfb
      13'h985: dout <= 8'b11111111; // 2437 : 255 - 0xff
      13'h986: dout <= 8'b11111111; // 2438 : 255 - 0xff
      13'h987: dout <= 8'b11111111; // 2439 : 255 - 0xff
      13'h988: dout <= 8'b00000000; // 2440 :   0 - 0x0
      13'h989: dout <= 8'b11011111; // 2441 : 223 - 0xdf
      13'h98A: dout <= 8'b11111111; // 2442 : 255 - 0xff
      13'h98B: dout <= 8'b11111111; // 2443 : 255 - 0xff
      13'h98C: dout <= 8'b11111111; // 2444 : 255 - 0xff
      13'h98D: dout <= 8'b11111111; // 2445 : 255 - 0xff
      13'h98E: dout <= 8'b11111111; // 2446 : 255 - 0xff
      13'h98F: dout <= 8'b11111111; // 2447 : 255 - 0xff
      13'h990: dout <= 8'b11111111; // 2448 : 255 - 0xff -- Sprite 0x99
      13'h991: dout <= 8'b11111111; // 2449 : 255 - 0xff
      13'h992: dout <= 8'b11111111; // 2450 : 255 - 0xff
      13'h993: dout <= 8'b11111111; // 2451 : 255 - 0xff
      13'h994: dout <= 8'b11111111; // 2452 : 255 - 0xff
      13'h995: dout <= 8'b11111111; // 2453 : 255 - 0xff
      13'h996: dout <= 8'b11111110; // 2454 : 254 - 0xfe
      13'h997: dout <= 8'b11111111; // 2455 : 255 - 0xff
      13'h998: dout <= 8'b11111111; // 2456 : 255 - 0xff
      13'h999: dout <= 8'b11111111; // 2457 : 255 - 0xff
      13'h99A: dout <= 8'b10111111; // 2458 : 191 - 0xbf
      13'h99B: dout <= 8'b11111111; // 2459 : 255 - 0xff
      13'h99C: dout <= 8'b11111111; // 2460 : 255 - 0xff
      13'h99D: dout <= 8'b11111111; // 2461 : 255 - 0xff
      13'h99E: dout <= 8'b11111111; // 2462 : 255 - 0xff
      13'h99F: dout <= 8'b11111111; // 2463 : 255 - 0xff
      13'h9A0: dout <= 8'b11111110; // 2464 : 254 - 0xfe -- Sprite 0x9a
      13'h9A1: dout <= 8'b11111111; // 2465 : 255 - 0xff
      13'h9A2: dout <= 8'b11111111; // 2466 : 255 - 0xff
      13'h9A3: dout <= 8'b11111111; // 2467 : 255 - 0xff
      13'h9A4: dout <= 8'b11111011; // 2468 : 251 - 0xfb
      13'h9A5: dout <= 8'b11111111; // 2469 : 255 - 0xff
      13'h9A6: dout <= 8'b11111111; // 2470 : 255 - 0xff
      13'h9A7: dout <= 8'b11111111; // 2471 : 255 - 0xff
      13'h9A8: dout <= 8'b00000000; // 2472 :   0 - 0x0
      13'h9A9: dout <= 8'b10111100; // 2473 : 188 - 0xbc
      13'h9AA: dout <= 8'b11111110; // 2474 : 254 - 0xfe
      13'h9AB: dout <= 8'b11111110; // 2475 : 254 - 0xfe
      13'h9AC: dout <= 8'b11111110; // 2476 : 254 - 0xfe
      13'h9AD: dout <= 8'b11111110; // 2477 : 254 - 0xfe
      13'h9AE: dout <= 8'b11111110; // 2478 : 254 - 0xfe
      13'h9AF: dout <= 8'b11111110; // 2479 : 254 - 0xfe
      13'h9B0: dout <= 8'b11111111; // 2480 : 255 - 0xff -- Sprite 0x9b
      13'h9B1: dout <= 8'b11111111; // 2481 : 255 - 0xff
      13'h9B2: dout <= 8'b11111111; // 2482 : 255 - 0xff
      13'h9B3: dout <= 8'b11111111; // 2483 : 255 - 0xff
      13'h9B4: dout <= 8'b11111111; // 2484 : 255 - 0xff
      13'h9B5: dout <= 8'b11111111; // 2485 : 255 - 0xff
      13'h9B6: dout <= 8'b11111111; // 2486 : 255 - 0xff
      13'h9B7: dout <= 8'b11111111; // 2487 : 255 - 0xff
      13'h9B8: dout <= 8'b11111110; // 2488 : 254 - 0xfe
      13'h9B9: dout <= 8'b11111110; // 2489 : 254 - 0xfe
      13'h9BA: dout <= 8'b10111110; // 2490 : 190 - 0xbe
      13'h9BB: dout <= 8'b11111110; // 2491 : 254 - 0xfe
      13'h9BC: dout <= 8'b11111110; // 2492 : 254 - 0xfe
      13'h9BD: dout <= 8'b11111110; // 2493 : 254 - 0xfe
      13'h9BE: dout <= 8'b11111110; // 2494 : 254 - 0xfe
      13'h9BF: dout <= 8'b11111110; // 2495 : 254 - 0xfe
      13'h9C0: dout <= 8'b11111111; // 2496 : 255 - 0xff -- Sprite 0x9c
      13'h9C1: dout <= 8'b11111111; // 2497 : 255 - 0xff
      13'h9C2: dout <= 8'b10100000; // 2498 : 160 - 0xa0
      13'h9C3: dout <= 8'b10010000; // 2499 : 144 - 0x90
      13'h9C4: dout <= 8'b10001000; // 2500 : 136 - 0x88
      13'h9C5: dout <= 8'b10000100; // 2501 : 132 - 0x84
      13'h9C6: dout <= 8'b01101010; // 2502 : 106 - 0x6a
      13'h9C7: dout <= 8'b00111111; // 2503 :  63 - 0x3f
      13'h9C8: dout <= 8'b00000000; // 2504 :   0 - 0x0
      13'h9C9: dout <= 8'b00111111; // 2505 :  63 - 0x3f
      13'h9CA: dout <= 8'b01011111; // 2506 :  95 - 0x5f
      13'h9CB: dout <= 8'b01101111; // 2507 : 111 - 0x6f
      13'h9CC: dout <= 8'b01110111; // 2508 : 119 - 0x77
      13'h9CD: dout <= 8'b01111011; // 2509 : 123 - 0x7b
      13'h9CE: dout <= 8'b00010101; // 2510 :  21 - 0x15
      13'h9CF: dout <= 8'b00000000; // 2511 :   0 - 0x0
      13'h9D0: dout <= 8'b11111111; // 2512 : 255 - 0xff -- Sprite 0x9d
      13'h9D1: dout <= 8'b11111111; // 2513 : 255 - 0xff
      13'h9D2: dout <= 8'b00100001; // 2514 :  33 - 0x21
      13'h9D3: dout <= 8'b00010001; // 2515 :  17 - 0x11
      13'h9D4: dout <= 8'b00001001; // 2516 :   9 - 0x9
      13'h9D5: dout <= 8'b00000101; // 2517 :   5 - 0x5
      13'h9D6: dout <= 8'b10101010; // 2518 : 170 - 0xaa
      13'h9D7: dout <= 8'b11111100; // 2519 : 252 - 0xfc
      13'h9D8: dout <= 8'b00000000; // 2520 :   0 - 0x0
      13'h9D9: dout <= 8'b10111110; // 2521 : 190 - 0xbe
      13'h9DA: dout <= 8'b11011110; // 2522 : 222 - 0xde
      13'h9DB: dout <= 8'b11101110; // 2523 : 238 - 0xee
      13'h9DC: dout <= 8'b11110110; // 2524 : 246 - 0xf6
      13'h9DD: dout <= 8'b11111010; // 2525 : 250 - 0xfa
      13'h9DE: dout <= 8'b01010100; // 2526 :  84 - 0x54
      13'h9DF: dout <= 8'b00000000; // 2527 :   0 - 0x0
      13'h9E0: dout <= 8'b11111111; // 2528 : 255 - 0xff -- Sprite 0x9e
      13'h9E1: dout <= 8'b11111111; // 2529 : 255 - 0xff
      13'h9E2: dout <= 8'b00100000; // 2530 :  32 - 0x20
      13'h9E3: dout <= 8'b00010000; // 2531 :  16 - 0x10
      13'h9E4: dout <= 8'b00001000; // 2532 :   8 - 0x8
      13'h9E5: dout <= 8'b00000100; // 2533 :   4 - 0x4
      13'h9E6: dout <= 8'b10101010; // 2534 : 170 - 0xaa
      13'h9E7: dout <= 8'b11111111; // 2535 : 255 - 0xff
      13'h9E8: dout <= 8'b00000000; // 2536 :   0 - 0x0
      13'h9E9: dout <= 8'b10111111; // 2537 : 191 - 0xbf
      13'h9EA: dout <= 8'b11011111; // 2538 : 223 - 0xdf
      13'h9EB: dout <= 8'b11101111; // 2539 : 239 - 0xef
      13'h9EC: dout <= 8'b11110111; // 2540 : 247 - 0xf7
      13'h9ED: dout <= 8'b11111011; // 2541 : 251 - 0xfb
      13'h9EE: dout <= 8'b01010101; // 2542 :  85 - 0x55
      13'h9EF: dout <= 8'b00000000; // 2543 :   0 - 0x0
      13'h9F0: dout <= 8'b00000000; // 2544 :   0 - 0x0 -- Sprite 0x9f
      13'h9F1: dout <= 8'b00000000; // 2545 :   0 - 0x0
      13'h9F2: dout <= 8'b00000000; // 2546 :   0 - 0x0
      13'h9F3: dout <= 8'b00000000; // 2547 :   0 - 0x0
      13'h9F4: dout <= 8'b00000000; // 2548 :   0 - 0x0
      13'h9F5: dout <= 8'b00000000; // 2549 :   0 - 0x0
      13'h9F6: dout <= 8'b00000000; // 2550 :   0 - 0x0
      13'h9F7: dout <= 8'b00000000; // 2551 :   0 - 0x0
      13'h9F8: dout <= 8'b00000000; // 2552 :   0 - 0x0
      13'h9F9: dout <= 8'b00000000; // 2553 :   0 - 0x0
      13'h9FA: dout <= 8'b00000000; // 2554 :   0 - 0x0
      13'h9FB: dout <= 8'b00000000; // 2555 :   0 - 0x0
      13'h9FC: dout <= 8'b00000000; // 2556 :   0 - 0x0
      13'h9FD: dout <= 8'b00000000; // 2557 :   0 - 0x0
      13'h9FE: dout <= 8'b00000000; // 2558 :   0 - 0x0
      13'h9FF: dout <= 8'b00000000; // 2559 :   0 - 0x0
      13'hA00: dout <= 8'b11111111; // 2560 : 255 - 0xff -- Sprite 0xa0
      13'hA01: dout <= 8'b11010101; // 2561 : 213 - 0xd5
      13'hA02: dout <= 8'b11111111; // 2562 : 255 - 0xff
      13'hA03: dout <= 8'b00000010; // 2563 :   2 - 0x2
      13'hA04: dout <= 8'b00000010; // 2564 :   2 - 0x2
      13'hA05: dout <= 8'b00000010; // 2565 :   2 - 0x2
      13'hA06: dout <= 8'b00000010; // 2566 :   2 - 0x2
      13'hA07: dout <= 8'b00000010; // 2567 :   2 - 0x2
      13'hA08: dout <= 8'b00000000; // 2568 :   0 - 0x0
      13'hA09: dout <= 8'b01111111; // 2569 : 127 - 0x7f
      13'hA0A: dout <= 8'b00000000; // 2570 :   0 - 0x0
      13'hA0B: dout <= 8'b00000001; // 2571 :   1 - 0x1
      13'hA0C: dout <= 8'b00000001; // 2572 :   1 - 0x1
      13'hA0D: dout <= 8'b00000001; // 2573 :   1 - 0x1
      13'hA0E: dout <= 8'b00000001; // 2574 :   1 - 0x1
      13'hA0F: dout <= 8'b00000001; // 2575 :   1 - 0x1
      13'hA10: dout <= 8'b00000010; // 2576 :   2 - 0x2 -- Sprite 0xa1
      13'hA11: dout <= 8'b00000010; // 2577 :   2 - 0x2
      13'hA12: dout <= 8'b00000010; // 2578 :   2 - 0x2
      13'hA13: dout <= 8'b00000010; // 2579 :   2 - 0x2
      13'hA14: dout <= 8'b00000010; // 2580 :   2 - 0x2
      13'hA15: dout <= 8'b00000010; // 2581 :   2 - 0x2
      13'hA16: dout <= 8'b00000010; // 2582 :   2 - 0x2
      13'hA17: dout <= 8'b00000010; // 2583 :   2 - 0x2
      13'hA18: dout <= 8'b00000001; // 2584 :   1 - 0x1
      13'hA19: dout <= 8'b00000001; // 2585 :   1 - 0x1
      13'hA1A: dout <= 8'b00000001; // 2586 :   1 - 0x1
      13'hA1B: dout <= 8'b00000001; // 2587 :   1 - 0x1
      13'hA1C: dout <= 8'b00000001; // 2588 :   1 - 0x1
      13'hA1D: dout <= 8'b00000001; // 2589 :   1 - 0x1
      13'hA1E: dout <= 8'b00000001; // 2590 :   1 - 0x1
      13'hA1F: dout <= 8'b00000001; // 2591 :   1 - 0x1
      13'hA20: dout <= 8'b11111111; // 2592 : 255 - 0xff -- Sprite 0xa2
      13'hA21: dout <= 8'b01010101; // 2593 :  85 - 0x55
      13'hA22: dout <= 8'b11111111; // 2594 : 255 - 0xff
      13'hA23: dout <= 8'b01000000; // 2595 :  64 - 0x40
      13'hA24: dout <= 8'b01000000; // 2596 :  64 - 0x40
      13'hA25: dout <= 8'b01000000; // 2597 :  64 - 0x40
      13'hA26: dout <= 8'b01000000; // 2598 :  64 - 0x40
      13'hA27: dout <= 8'b01000000; // 2599 :  64 - 0x40
      13'hA28: dout <= 8'b00000000; // 2600 :   0 - 0x0
      13'hA29: dout <= 8'b11111110; // 2601 : 254 - 0xfe
      13'hA2A: dout <= 8'b00000000; // 2602 :   0 - 0x0
      13'hA2B: dout <= 8'b10000000; // 2603 : 128 - 0x80
      13'hA2C: dout <= 8'b10000000; // 2604 : 128 - 0x80
      13'hA2D: dout <= 8'b10000000; // 2605 : 128 - 0x80
      13'hA2E: dout <= 8'b10000000; // 2606 : 128 - 0x80
      13'hA2F: dout <= 8'b10000000; // 2607 : 128 - 0x80
      13'hA30: dout <= 8'b01000000; // 2608 :  64 - 0x40 -- Sprite 0xa3
      13'hA31: dout <= 8'b01000000; // 2609 :  64 - 0x40
      13'hA32: dout <= 8'b01000000; // 2610 :  64 - 0x40
      13'hA33: dout <= 8'b01000000; // 2611 :  64 - 0x40
      13'hA34: dout <= 8'b01000000; // 2612 :  64 - 0x40
      13'hA35: dout <= 8'b01000000; // 2613 :  64 - 0x40
      13'hA36: dout <= 8'b01000000; // 2614 :  64 - 0x40
      13'hA37: dout <= 8'b01000000; // 2615 :  64 - 0x40
      13'hA38: dout <= 8'b10000000; // 2616 : 128 - 0x80
      13'hA39: dout <= 8'b10000000; // 2617 : 128 - 0x80
      13'hA3A: dout <= 8'b10000000; // 2618 : 128 - 0x80
      13'hA3B: dout <= 8'b10000000; // 2619 : 128 - 0x80
      13'hA3C: dout <= 8'b10000000; // 2620 : 128 - 0x80
      13'hA3D: dout <= 8'b10000000; // 2621 : 128 - 0x80
      13'hA3E: dout <= 8'b10000000; // 2622 : 128 - 0x80
      13'hA3F: dout <= 8'b10000000; // 2623 : 128 - 0x80
      13'hA40: dout <= 8'b00110001; // 2624 :  49 - 0x31 -- Sprite 0xa4
      13'hA41: dout <= 8'b01001000; // 2625 :  72 - 0x48
      13'hA42: dout <= 8'b01000101; // 2626 :  69 - 0x45
      13'hA43: dout <= 8'b10000101; // 2627 : 133 - 0x85
      13'hA44: dout <= 8'b10000011; // 2628 : 131 - 0x83
      13'hA45: dout <= 8'b10000010; // 2629 : 130 - 0x82
      13'hA46: dout <= 8'b01100010; // 2630 :  98 - 0x62
      13'hA47: dout <= 8'b00010010; // 2631 :  18 - 0x12
      13'hA48: dout <= 8'b00000000; // 2632 :   0 - 0x0
      13'hA49: dout <= 8'b00110000; // 2633 :  48 - 0x30
      13'hA4A: dout <= 8'b00111000; // 2634 :  56 - 0x38
      13'hA4B: dout <= 8'b01111000; // 2635 : 120 - 0x78
      13'hA4C: dout <= 8'b01111100; // 2636 : 124 - 0x7c
      13'hA4D: dout <= 8'b01111101; // 2637 : 125 - 0x7d
      13'hA4E: dout <= 8'b00011101; // 2638 :  29 - 0x1d
      13'hA4F: dout <= 8'b00001101; // 2639 :  13 - 0xd
      13'hA50: dout <= 8'b00110010; // 2640 :  50 - 0x32 -- Sprite 0xa5
      13'hA51: dout <= 8'b00100010; // 2641 :  34 - 0x22
      13'hA52: dout <= 8'b01000010; // 2642 :  66 - 0x42
      13'hA53: dout <= 8'b01000000; // 2643 :  64 - 0x40
      13'hA54: dout <= 8'b01000000; // 2644 :  64 - 0x40
      13'hA55: dout <= 8'b00100000; // 2645 :  32 - 0x20
      13'hA56: dout <= 8'b00011110; // 2646 :  30 - 0x1e
      13'hA57: dout <= 8'b00000111; // 2647 :   7 - 0x7
      13'hA58: dout <= 8'b00001101; // 2648 :  13 - 0xd
      13'hA59: dout <= 8'b00011101; // 2649 :  29 - 0x1d
      13'hA5A: dout <= 8'b00111101; // 2650 :  61 - 0x3d
      13'hA5B: dout <= 8'b00111111; // 2651 :  63 - 0x3f
      13'hA5C: dout <= 8'b00111111; // 2652 :  63 - 0x3f
      13'hA5D: dout <= 8'b00011111; // 2653 :  31 - 0x1f
      13'hA5E: dout <= 8'b00000001; // 2654 :   1 - 0x1
      13'hA5F: dout <= 8'b00000000; // 2655 :   0 - 0x0
      13'hA60: dout <= 8'b10000000; // 2656 : 128 - 0x80 -- Sprite 0xa6
      13'hA61: dout <= 8'b11100000; // 2657 : 224 - 0xe0
      13'hA62: dout <= 8'b00111000; // 2658 :  56 - 0x38
      13'hA63: dout <= 8'b00100100; // 2659 :  36 - 0x24
      13'hA64: dout <= 8'b00000100; // 2660 :   4 - 0x4
      13'hA65: dout <= 8'b00001000; // 2661 :   8 - 0x8
      13'hA66: dout <= 8'b00110000; // 2662 :  48 - 0x30
      13'hA67: dout <= 8'b00100000; // 2663 :  32 - 0x20
      13'hA68: dout <= 8'b00000000; // 2664 :   0 - 0x0
      13'hA69: dout <= 8'b00000000; // 2665 :   0 - 0x0
      13'hA6A: dout <= 8'b11100000; // 2666 : 224 - 0xe0
      13'hA6B: dout <= 8'b11111000; // 2667 : 248 - 0xf8
      13'hA6C: dout <= 8'b11111000; // 2668 : 248 - 0xf8
      13'hA6D: dout <= 8'b11110000; // 2669 : 240 - 0xf0
      13'hA6E: dout <= 8'b11000000; // 2670 : 192 - 0xc0
      13'hA6F: dout <= 8'b11000000; // 2671 : 192 - 0xc0
      13'hA70: dout <= 8'b00110000; // 2672 :  48 - 0x30 -- Sprite 0xa7
      13'hA71: dout <= 8'b00001000; // 2673 :   8 - 0x8
      13'hA72: dout <= 8'b00001000; // 2674 :   8 - 0x8
      13'hA73: dout <= 8'b00110000; // 2675 :  48 - 0x30
      13'hA74: dout <= 8'b00100000; // 2676 :  32 - 0x20
      13'hA75: dout <= 8'b00100000; // 2677 :  32 - 0x20
      13'hA76: dout <= 8'b00110000; // 2678 :  48 - 0x30
      13'hA77: dout <= 8'b11110000; // 2679 : 240 - 0xf0
      13'hA78: dout <= 8'b11000000; // 2680 : 192 - 0xc0
      13'hA79: dout <= 8'b11110000; // 2681 : 240 - 0xf0
      13'hA7A: dout <= 8'b11110000; // 2682 : 240 - 0xf0
      13'hA7B: dout <= 8'b11000000; // 2683 : 192 - 0xc0
      13'hA7C: dout <= 8'b11000000; // 2684 : 192 - 0xc0
      13'hA7D: dout <= 8'b11000000; // 2685 : 192 - 0xc0
      13'hA7E: dout <= 8'b11000000; // 2686 : 192 - 0xc0
      13'hA7F: dout <= 8'b00000000; // 2687 :   0 - 0x0
      13'hA80: dout <= 8'b11111111; // 2688 : 255 - 0xff -- Sprite 0xa8
      13'hA81: dout <= 8'b11010010; // 2689 : 210 - 0xd2
      13'hA82: dout <= 8'b11110100; // 2690 : 244 - 0xf4
      13'hA83: dout <= 8'b11011000; // 2691 : 216 - 0xd8
      13'hA84: dout <= 8'b11111000; // 2692 : 248 - 0xf8
      13'hA85: dout <= 8'b11010100; // 2693 : 212 - 0xd4
      13'hA86: dout <= 8'b11110010; // 2694 : 242 - 0xf2
      13'hA87: dout <= 8'b11010001; // 2695 : 209 - 0xd1
      13'hA88: dout <= 8'b00000000; // 2696 :   0 - 0x0
      13'hA89: dout <= 8'b01100000; // 2697 :  96 - 0x60
      13'hA8A: dout <= 8'b01100000; // 2698 :  96 - 0x60
      13'hA8B: dout <= 8'b01100000; // 2699 :  96 - 0x60
      13'hA8C: dout <= 8'b01100000; // 2700 :  96 - 0x60
      13'hA8D: dout <= 8'b01100000; // 2701 :  96 - 0x60
      13'hA8E: dout <= 8'b01100000; // 2702 :  96 - 0x60
      13'hA8F: dout <= 8'b01100000; // 2703 :  96 - 0x60
      13'hA90: dout <= 8'b11110001; // 2704 : 241 - 0xf1 -- Sprite 0xa9
      13'hA91: dout <= 8'b11010010; // 2705 : 210 - 0xd2
      13'hA92: dout <= 8'b11110100; // 2706 : 244 - 0xf4
      13'hA93: dout <= 8'b11011000; // 2707 : 216 - 0xd8
      13'hA94: dout <= 8'b11111000; // 2708 : 248 - 0xf8
      13'hA95: dout <= 8'b11010100; // 2709 : 212 - 0xd4
      13'hA96: dout <= 8'b11110010; // 2710 : 242 - 0xf2
      13'hA97: dout <= 8'b11111111; // 2711 : 255 - 0xff
      13'hA98: dout <= 8'b01100000; // 2712 :  96 - 0x60
      13'hA99: dout <= 8'b01100000; // 2713 :  96 - 0x60
      13'hA9A: dout <= 8'b01100000; // 2714 :  96 - 0x60
      13'hA9B: dout <= 8'b01100000; // 2715 :  96 - 0x60
      13'hA9C: dout <= 8'b01100000; // 2716 :  96 - 0x60
      13'hA9D: dout <= 8'b01100000; // 2717 :  96 - 0x60
      13'hA9E: dout <= 8'b01100000; // 2718 :  96 - 0x60
      13'hA9F: dout <= 8'b00000000; // 2719 :   0 - 0x0
      13'hAA0: dout <= 8'b11111111; // 2720 : 255 - 0xff -- Sprite 0xaa
      13'hAA1: dout <= 8'b01000010; // 2721 :  66 - 0x42
      13'hAA2: dout <= 8'b00100100; // 2722 :  36 - 0x24
      13'hAA3: dout <= 8'b00011000; // 2723 :  24 - 0x18
      13'hAA4: dout <= 8'b00011000; // 2724 :  24 - 0x18
      13'hAA5: dout <= 8'b00100100; // 2725 :  36 - 0x24
      13'hAA6: dout <= 8'b01000010; // 2726 :  66 - 0x42
      13'hAA7: dout <= 8'b10000001; // 2727 : 129 - 0x81
      13'hAA8: dout <= 8'b00000000; // 2728 :   0 - 0x0
      13'hAA9: dout <= 8'b00000000; // 2729 :   0 - 0x0
      13'hAAA: dout <= 8'b00000000; // 2730 :   0 - 0x0
      13'hAAB: dout <= 8'b00000000; // 2731 :   0 - 0x0
      13'hAAC: dout <= 8'b00000000; // 2732 :   0 - 0x0
      13'hAAD: dout <= 8'b00000000; // 2733 :   0 - 0x0
      13'hAAE: dout <= 8'b00000000; // 2734 :   0 - 0x0
      13'hAAF: dout <= 8'b00000000; // 2735 :   0 - 0x0
      13'hAB0: dout <= 8'b10000001; // 2736 : 129 - 0x81 -- Sprite 0xab
      13'hAB1: dout <= 8'b01000010; // 2737 :  66 - 0x42
      13'hAB2: dout <= 8'b00100100; // 2738 :  36 - 0x24
      13'hAB3: dout <= 8'b00011000; // 2739 :  24 - 0x18
      13'hAB4: dout <= 8'b00011000; // 2740 :  24 - 0x18
      13'hAB5: dout <= 8'b00100100; // 2741 :  36 - 0x24
      13'hAB6: dout <= 8'b01000010; // 2742 :  66 - 0x42
      13'hAB7: dout <= 8'b11111111; // 2743 : 255 - 0xff
      13'hAB8: dout <= 8'b00000000; // 2744 :   0 - 0x0
      13'hAB9: dout <= 8'b00000000; // 2745 :   0 - 0x0
      13'hABA: dout <= 8'b00000000; // 2746 :   0 - 0x0
      13'hABB: dout <= 8'b00000000; // 2747 :   0 - 0x0
      13'hABC: dout <= 8'b00000000; // 2748 :   0 - 0x0
      13'hABD: dout <= 8'b00000000; // 2749 :   0 - 0x0
      13'hABE: dout <= 8'b00000000; // 2750 :   0 - 0x0
      13'hABF: dout <= 8'b00000000; // 2751 :   0 - 0x0
      13'hAC0: dout <= 8'b11111111; // 2752 : 255 - 0xff -- Sprite 0xac
      13'hAC1: dout <= 8'b01001101; // 2753 :  77 - 0x4d
      13'hAC2: dout <= 8'b00101111; // 2754 :  47 - 0x2f
      13'hAC3: dout <= 8'b00011101; // 2755 :  29 - 0x1d
      13'hAC4: dout <= 8'b00011111; // 2756 :  31 - 0x1f
      13'hAC5: dout <= 8'b00101101; // 2757 :  45 - 0x2d
      13'hAC6: dout <= 8'b01001111; // 2758 :  79 - 0x4f
      13'hAC7: dout <= 8'b10001101; // 2759 : 141 - 0x8d
      13'hAC8: dout <= 8'b00000000; // 2760 :   0 - 0x0
      13'hAC9: dout <= 8'b00000110; // 2761 :   6 - 0x6
      13'hACA: dout <= 8'b00000110; // 2762 :   6 - 0x6
      13'hACB: dout <= 8'b00000110; // 2763 :   6 - 0x6
      13'hACC: dout <= 8'b00000110; // 2764 :   6 - 0x6
      13'hACD: dout <= 8'b00000110; // 2765 :   6 - 0x6
      13'hACE: dout <= 8'b00000110; // 2766 :   6 - 0x6
      13'hACF: dout <= 8'b00000110; // 2767 :   6 - 0x6
      13'hAD0: dout <= 8'b10001111; // 2768 : 143 - 0x8f -- Sprite 0xad
      13'hAD1: dout <= 8'b01001101; // 2769 :  77 - 0x4d
      13'hAD2: dout <= 8'b00101111; // 2770 :  47 - 0x2f
      13'hAD3: dout <= 8'b00011101; // 2771 :  29 - 0x1d
      13'hAD4: dout <= 8'b00011111; // 2772 :  31 - 0x1f
      13'hAD5: dout <= 8'b00101101; // 2773 :  45 - 0x2d
      13'hAD6: dout <= 8'b01001111; // 2774 :  79 - 0x4f
      13'hAD7: dout <= 8'b11111111; // 2775 : 255 - 0xff
      13'hAD8: dout <= 8'b00000110; // 2776 :   6 - 0x6
      13'hAD9: dout <= 8'b00000110; // 2777 :   6 - 0x6
      13'hADA: dout <= 8'b00000110; // 2778 :   6 - 0x6
      13'hADB: dout <= 8'b00000110; // 2779 :   6 - 0x6
      13'hADC: dout <= 8'b00000110; // 2780 :   6 - 0x6
      13'hADD: dout <= 8'b00000110; // 2781 :   6 - 0x6
      13'hADE: dout <= 8'b00000110; // 2782 :   6 - 0x6
      13'hADF: dout <= 8'b00000000; // 2783 :   0 - 0x0
      13'hAE0: dout <= 8'b00000001; // 2784 :   1 - 0x1 -- Sprite 0xae
      13'hAE1: dout <= 8'b00000011; // 2785 :   3 - 0x3
      13'hAE2: dout <= 8'b00000110; // 2786 :   6 - 0x6
      13'hAE3: dout <= 8'b00000111; // 2787 :   7 - 0x7
      13'hAE4: dout <= 8'b00000111; // 2788 :   7 - 0x7
      13'hAE5: dout <= 8'b00000111; // 2789 :   7 - 0x7
      13'hAE6: dout <= 8'b00000110; // 2790 :   6 - 0x6
      13'hAE7: dout <= 8'b00000111; // 2791 :   7 - 0x7
      13'hAE8: dout <= 8'b00000000; // 2792 :   0 - 0x0
      13'hAE9: dout <= 8'b00000001; // 2793 :   1 - 0x1
      13'hAEA: dout <= 8'b00000011; // 2794 :   3 - 0x3
      13'hAEB: dout <= 8'b00000010; // 2795 :   2 - 0x2
      13'hAEC: dout <= 8'b00000010; // 2796 :   2 - 0x2
      13'hAED: dout <= 8'b00000000; // 2797 :   0 - 0x0
      13'hAEE: dout <= 8'b00000011; // 2798 :   3 - 0x3
      13'hAEF: dout <= 8'b00000010; // 2799 :   2 - 0x2
      13'hAF0: dout <= 8'b00000110; // 2800 :   6 - 0x6 -- Sprite 0xaf
      13'hAF1: dout <= 8'b00000110; // 2801 :   6 - 0x6
      13'hAF2: dout <= 8'b00001110; // 2802 :  14 - 0xe
      13'hAF3: dout <= 8'b00001111; // 2803 :  15 - 0xf
      13'hAF4: dout <= 8'b00001110; // 2804 :  14 - 0xe
      13'hAF5: dout <= 8'b00011010; // 2805 :  26 - 0x1a
      13'hAF6: dout <= 8'b00011011; // 2806 :  27 - 0x1b
      13'hAF7: dout <= 8'b00001111; // 2807 :  15 - 0xf
      13'hAF8: dout <= 8'b00000001; // 2808 :   1 - 0x1
      13'hAF9: dout <= 8'b00000011; // 2809 :   3 - 0x3
      13'hAFA: dout <= 8'b00000101; // 2810 :   5 - 0x5
      13'hAFB: dout <= 8'b00000100; // 2811 :   4 - 0x4
      13'hAFC: dout <= 8'b00000101; // 2812 :   5 - 0x5
      13'hAFD: dout <= 8'b00001101; // 2813 :  13 - 0xd
      13'hAFE: dout <= 8'b00001100; // 2814 :  12 - 0xc
      13'hAFF: dout <= 8'b00000001; // 2815 :   1 - 0x1
      13'hB00: dout <= 8'b00000000; // 2816 :   0 - 0x0 -- Sprite 0xb0
      13'hB01: dout <= 8'b11000000; // 2817 : 192 - 0xc0
      13'hB02: dout <= 8'b11110000; // 2818 : 240 - 0xf0
      13'hB03: dout <= 8'b10001000; // 2819 : 136 - 0x88
      13'hB04: dout <= 8'b00010100; // 2820 :  20 - 0x14
      13'hB05: dout <= 8'b01101000; // 2821 : 104 - 0x68
      13'hB06: dout <= 8'b10101000; // 2822 : 168 - 0xa8
      13'hB07: dout <= 8'b00101100; // 2823 :  44 - 0x2c
      13'hB08: dout <= 8'b00000000; // 2824 :   0 - 0x0
      13'hB09: dout <= 8'b00000000; // 2825 :   0 - 0x0
      13'hB0A: dout <= 8'b01000000; // 2826 :  64 - 0x40
      13'hB0B: dout <= 8'b11110000; // 2827 : 240 - 0xf0
      13'hB0C: dout <= 8'b11101000; // 2828 : 232 - 0xe8
      13'hB0D: dout <= 8'b10010000; // 2829 : 144 - 0x90
      13'hB0E: dout <= 8'b01010000; // 2830 :  80 - 0x50
      13'hB0F: dout <= 8'b11010000; // 2831 : 208 - 0xd0
      13'hB10: dout <= 8'b00000100; // 2832 :   4 - 0x4 -- Sprite 0xb1
      13'hB11: dout <= 8'b00111000; // 2833 :  56 - 0x38
      13'hB12: dout <= 8'b00010000; // 2834 :  16 - 0x10
      13'hB13: dout <= 8'b10100000; // 2835 : 160 - 0xa0
      13'hB14: dout <= 8'b01100000; // 2836 :  96 - 0x60
      13'hB15: dout <= 8'b00100000; // 2837 :  32 - 0x20
      13'hB16: dout <= 8'b00010000; // 2838 :  16 - 0x10
      13'hB17: dout <= 8'b10001000; // 2839 : 136 - 0x88
      13'hB18: dout <= 8'b11111000; // 2840 : 248 - 0xf8
      13'hB19: dout <= 8'b11000000; // 2841 : 192 - 0xc0
      13'hB1A: dout <= 8'b11100000; // 2842 : 224 - 0xe0
      13'hB1B: dout <= 8'b01000000; // 2843 :  64 - 0x40
      13'hB1C: dout <= 8'b10000000; // 2844 : 128 - 0x80
      13'hB1D: dout <= 8'b11000000; // 2845 : 192 - 0xc0
      13'hB1E: dout <= 8'b11100000; // 2846 : 224 - 0xe0
      13'hB1F: dout <= 8'b01110000; // 2847 : 112 - 0x70
      13'hB20: dout <= 8'b00001111; // 2848 :  15 - 0xf -- Sprite 0xb2
      13'hB21: dout <= 8'b00011011; // 2849 :  27 - 0x1b
      13'hB22: dout <= 8'b00011011; // 2850 :  27 - 0x1b
      13'hB23: dout <= 8'b00001110; // 2851 :  14 - 0xe
      13'hB24: dout <= 8'b00000110; // 2852 :   6 - 0x6
      13'hB25: dout <= 8'b00001100; // 2853 :  12 - 0xc
      13'hB26: dout <= 8'b00001100; // 2854 :  12 - 0xc
      13'hB27: dout <= 8'b00111111; // 2855 :  63 - 0x3f
      13'hB28: dout <= 8'b00000001; // 2856 :   1 - 0x1
      13'hB29: dout <= 8'b00001101; // 2857 :  13 - 0xd
      13'hB2A: dout <= 8'b00001101; // 2858 :  13 - 0xd
      13'hB2B: dout <= 8'b00000011; // 2859 :   3 - 0x3
      13'hB2C: dout <= 8'b00000011; // 2860 :   3 - 0x3
      13'hB2D: dout <= 8'b00000111; // 2861 :   7 - 0x7
      13'hB2E: dout <= 8'b00000111; // 2862 :   7 - 0x7
      13'hB2F: dout <= 8'b00000000; // 2863 :   0 - 0x0
      13'hB30: dout <= 8'b01111111; // 2864 : 127 - 0x7f -- Sprite 0xb3
      13'hB31: dout <= 8'b01100000; // 2865 :  96 - 0x60
      13'hB32: dout <= 8'b01100000; // 2866 :  96 - 0x60
      13'hB33: dout <= 8'b01100000; // 2867 :  96 - 0x60
      13'hB34: dout <= 8'b01100000; // 2868 :  96 - 0x60
      13'hB35: dout <= 8'b01100000; // 2869 :  96 - 0x60
      13'hB36: dout <= 8'b01101010; // 2870 : 106 - 0x6a
      13'hB37: dout <= 8'b01111111; // 2871 : 127 - 0x7f
      13'hB38: dout <= 8'b00111111; // 2872 :  63 - 0x3f
      13'hB39: dout <= 8'b00111111; // 2873 :  63 - 0x3f
      13'hB3A: dout <= 8'b00111111; // 2874 :  63 - 0x3f
      13'hB3B: dout <= 8'b00111111; // 2875 :  63 - 0x3f
      13'hB3C: dout <= 8'b00111111; // 2876 :  63 - 0x3f
      13'hB3D: dout <= 8'b00111111; // 2877 :  63 - 0x3f
      13'hB3E: dout <= 8'b00110101; // 2878 :  53 - 0x35
      13'hB3F: dout <= 8'b00000000; // 2879 :   0 - 0x0
      13'hB40: dout <= 8'b01001000; // 2880 :  72 - 0x48 -- Sprite 0xb4
      13'hB41: dout <= 8'b00110000; // 2881 :  48 - 0x30
      13'hB42: dout <= 8'b00010000; // 2882 :  16 - 0x10
      13'hB43: dout <= 8'b00010000; // 2883 :  16 - 0x10
      13'hB44: dout <= 8'b00001000; // 2884 :   8 - 0x8
      13'hB45: dout <= 8'b00001000; // 2885 :   8 - 0x8
      13'hB46: dout <= 8'b00001000; // 2886 :   8 - 0x8
      13'hB47: dout <= 8'b11111100; // 2887 : 252 - 0xfc
      13'hB48: dout <= 8'b10110000; // 2888 : 176 - 0xb0
      13'hB49: dout <= 8'b11000000; // 2889 : 192 - 0xc0
      13'hB4A: dout <= 8'b11100000; // 2890 : 224 - 0xe0
      13'hB4B: dout <= 8'b11100000; // 2891 : 224 - 0xe0
      13'hB4C: dout <= 8'b11110000; // 2892 : 240 - 0xf0
      13'hB4D: dout <= 8'b11110000; // 2893 : 240 - 0xf0
      13'hB4E: dout <= 8'b11110000; // 2894 : 240 - 0xf0
      13'hB4F: dout <= 8'b00000000; // 2895 :   0 - 0x0
      13'hB50: dout <= 8'b11111110; // 2896 : 254 - 0xfe -- Sprite 0xb5
      13'hB51: dout <= 8'b00000110; // 2897 :   6 - 0x6
      13'hB52: dout <= 8'b00000010; // 2898 :   2 - 0x2
      13'hB53: dout <= 8'b00000110; // 2899 :   6 - 0x6
      13'hB54: dout <= 8'b00000010; // 2900 :   2 - 0x2
      13'hB55: dout <= 8'b00000110; // 2901 :   6 - 0x6
      13'hB56: dout <= 8'b10101010; // 2902 : 170 - 0xaa
      13'hB57: dout <= 8'b11111110; // 2903 : 254 - 0xfe
      13'hB58: dout <= 8'b11111100; // 2904 : 252 - 0xfc
      13'hB59: dout <= 8'b11111000; // 2905 : 248 - 0xf8
      13'hB5A: dout <= 8'b11111100; // 2906 : 252 - 0xfc
      13'hB5B: dout <= 8'b11111000; // 2907 : 248 - 0xf8
      13'hB5C: dout <= 8'b11111100; // 2908 : 252 - 0xfc
      13'hB5D: dout <= 8'b11111000; // 2909 : 248 - 0xf8
      13'hB5E: dout <= 8'b01010100; // 2910 :  84 - 0x54
      13'hB5F: dout <= 8'b00000000; // 2911 :   0 - 0x0
      13'hB60: dout <= 8'b11111111; // 2912 : 255 - 0xff -- Sprite 0xb6
      13'hB61: dout <= 8'b10000000; // 2913 : 128 - 0x80
      13'hB62: dout <= 8'b10000000; // 2914 : 128 - 0x80
      13'hB63: dout <= 8'b10000000; // 2915 : 128 - 0x80
      13'hB64: dout <= 8'b10000000; // 2916 : 128 - 0x80
      13'hB65: dout <= 8'b10000000; // 2917 : 128 - 0x80
      13'hB66: dout <= 8'b10010101; // 2918 : 149 - 0x95
      13'hB67: dout <= 8'b11111111; // 2919 : 255 - 0xff
      13'hB68: dout <= 8'b00000000; // 2920 :   0 - 0x0
      13'hB69: dout <= 8'b01111111; // 2921 : 127 - 0x7f
      13'hB6A: dout <= 8'b01111111; // 2922 : 127 - 0x7f
      13'hB6B: dout <= 8'b01111111; // 2923 : 127 - 0x7f
      13'hB6C: dout <= 8'b01111111; // 2924 : 127 - 0x7f
      13'hB6D: dout <= 8'b01111111; // 2925 : 127 - 0x7f
      13'hB6E: dout <= 8'b01101010; // 2926 : 106 - 0x6a
      13'hB6F: dout <= 8'b00000000; // 2927 :   0 - 0x0
      13'hB70: dout <= 8'b11111111; // 2928 : 255 - 0xff -- Sprite 0xb7
      13'hB71: dout <= 8'b10000100; // 2929 : 132 - 0x84
      13'hB72: dout <= 8'b10001100; // 2930 : 140 - 0x8c
      13'hB73: dout <= 8'b10000100; // 2931 : 132 - 0x84
      13'hB74: dout <= 8'b10001100; // 2932 : 140 - 0x8c
      13'hB75: dout <= 8'b10000100; // 2933 : 132 - 0x84
      13'hB76: dout <= 8'b10101100; // 2934 : 172 - 0xac
      13'hB77: dout <= 8'b11111111; // 2935 : 255 - 0xff
      13'hB78: dout <= 8'b00000000; // 2936 :   0 - 0x0
      13'hB79: dout <= 8'b01111011; // 2937 : 123 - 0x7b
      13'hB7A: dout <= 8'b01110011; // 2938 : 115 - 0x73
      13'hB7B: dout <= 8'b01111011; // 2939 : 123 - 0x7b
      13'hB7C: dout <= 8'b01110011; // 2940 : 115 - 0x73
      13'hB7D: dout <= 8'b01111011; // 2941 : 123 - 0x7b
      13'hB7E: dout <= 8'b01010011; // 2942 :  83 - 0x53
      13'hB7F: dout <= 8'b00000000; // 2943 :   0 - 0x0
      13'hB80: dout <= 8'b11111111; // 2944 : 255 - 0xff -- Sprite 0xb8
      13'hB81: dout <= 8'b00100001; // 2945 :  33 - 0x21
      13'hB82: dout <= 8'b01100001; // 2946 :  97 - 0x61
      13'hB83: dout <= 8'b00100011; // 2947 :  35 - 0x23
      13'hB84: dout <= 8'b01100001; // 2948 :  97 - 0x61
      13'hB85: dout <= 8'b00100011; // 2949 :  35 - 0x23
      13'hB86: dout <= 8'b01100101; // 2950 : 101 - 0x65
      13'hB87: dout <= 8'b11111111; // 2951 : 255 - 0xff
      13'hB88: dout <= 8'b00000000; // 2952 :   0 - 0x0
      13'hB89: dout <= 8'b11011110; // 2953 : 222 - 0xde
      13'hB8A: dout <= 8'b10011110; // 2954 : 158 - 0x9e
      13'hB8B: dout <= 8'b11011100; // 2955 : 220 - 0xdc
      13'hB8C: dout <= 8'b10011110; // 2956 : 158 - 0x9e
      13'hB8D: dout <= 8'b11011100; // 2957 : 220 - 0xdc
      13'hB8E: dout <= 8'b10011010; // 2958 : 154 - 0x9a
      13'hB8F: dout <= 8'b00000000; // 2959 :   0 - 0x0
      13'hB90: dout <= 8'b11111111; // 2960 : 255 - 0xff -- Sprite 0xb9
      13'hB91: dout <= 8'b00000001; // 2961 :   1 - 0x1
      13'hB92: dout <= 8'b00000011; // 2962 :   3 - 0x3
      13'hB93: dout <= 8'b00000001; // 2963 :   1 - 0x1
      13'hB94: dout <= 8'b00000011; // 2964 :   3 - 0x3
      13'hB95: dout <= 8'b00000001; // 2965 :   1 - 0x1
      13'hB96: dout <= 8'b10101011; // 2966 : 171 - 0xab
      13'hB97: dout <= 8'b11111111; // 2967 : 255 - 0xff
      13'hB98: dout <= 8'b00000000; // 2968 :   0 - 0x0
      13'hB99: dout <= 8'b11111110; // 2969 : 254 - 0xfe
      13'hB9A: dout <= 8'b11111100; // 2970 : 252 - 0xfc
      13'hB9B: dout <= 8'b11111110; // 2971 : 254 - 0xfe
      13'hB9C: dout <= 8'b11111100; // 2972 : 252 - 0xfc
      13'hB9D: dout <= 8'b11111110; // 2973 : 254 - 0xfe
      13'hB9E: dout <= 8'b01010100; // 2974 :  84 - 0x54
      13'hB9F: dout <= 8'b00000000; // 2975 :   0 - 0x0
      13'hBA0: dout <= 8'b11111111; // 2976 : 255 - 0xff -- Sprite 0xba
      13'hBA1: dout <= 8'b11010101; // 2977 : 213 - 0xd5
      13'hBA2: dout <= 8'b10101010; // 2978 : 170 - 0xaa
      13'hBA3: dout <= 8'b11111111; // 2979 : 255 - 0xff
      13'hBA4: dout <= 8'b10000000; // 2980 : 128 - 0x80
      13'hBA5: dout <= 8'b10000000; // 2981 : 128 - 0x80
      13'hBA6: dout <= 8'b10010101; // 2982 : 149 - 0x95
      13'hBA7: dout <= 8'b11111111; // 2983 : 255 - 0xff
      13'hBA8: dout <= 8'b00000000; // 2984 :   0 - 0x0
      13'hBA9: dout <= 8'b01111111; // 2985 : 127 - 0x7f
      13'hBAA: dout <= 8'b01111111; // 2986 : 127 - 0x7f
      13'hBAB: dout <= 8'b00000000; // 2987 :   0 - 0x0
      13'hBAC: dout <= 8'b01111111; // 2988 : 127 - 0x7f
      13'hBAD: dout <= 8'b01111111; // 2989 : 127 - 0x7f
      13'hBAE: dout <= 8'b01101010; // 2990 : 106 - 0x6a
      13'hBAF: dout <= 8'b00000000; // 2991 :   0 - 0x0
      13'hBB0: dout <= 8'b00000000; // 2992 :   0 - 0x0 -- Sprite 0xbb
      13'hBB1: dout <= 8'b00000000; // 2993 :   0 - 0x0
      13'hBB2: dout <= 8'b00000000; // 2994 :   0 - 0x0
      13'hBB3: dout <= 8'b00000000; // 2995 :   0 - 0x0
      13'hBB4: dout <= 8'b00000000; // 2996 :   0 - 0x0
      13'hBB5: dout <= 8'b00000000; // 2997 :   0 - 0x0
      13'hBB6: dout <= 8'b00000000; // 2998 :   0 - 0x0
      13'hBB7: dout <= 8'b00000000; // 2999 :   0 - 0x0
      13'hBB8: dout <= 8'b00000000; // 3000 :   0 - 0x0
      13'hBB9: dout <= 8'b00000000; // 3001 :   0 - 0x0
      13'hBBA: dout <= 8'b00000000; // 3002 :   0 - 0x0
      13'hBBB: dout <= 8'b00000000; // 3003 :   0 - 0x0
      13'hBBC: dout <= 8'b00000000; // 3004 :   0 - 0x0
      13'hBBD: dout <= 8'b00000000; // 3005 :   0 - 0x0
      13'hBBE: dout <= 8'b00000000; // 3006 :   0 - 0x0
      13'hBBF: dout <= 8'b00000000; // 3007 :   0 - 0x0
      13'hBC0: dout <= 8'b11111111; // 3008 : 255 - 0xff -- Sprite 0xbc
      13'hBC1: dout <= 8'b01010101; // 3009 :  85 - 0x55
      13'hBC2: dout <= 8'b10101011; // 3010 : 171 - 0xab
      13'hBC3: dout <= 8'b11111111; // 3011 : 255 - 0xff
      13'hBC4: dout <= 8'b01100001; // 3012 :  97 - 0x61
      13'hBC5: dout <= 8'b00100011; // 3013 :  35 - 0x23
      13'hBC6: dout <= 8'b01100101; // 3014 : 101 - 0x65
      13'hBC7: dout <= 8'b11111111; // 3015 : 255 - 0xff
      13'hBC8: dout <= 8'b00000000; // 3016 :   0 - 0x0
      13'hBC9: dout <= 8'b11111110; // 3017 : 254 - 0xfe
      13'hBCA: dout <= 8'b11111110; // 3018 : 254 - 0xfe
      13'hBCB: dout <= 8'b00000000; // 3019 :   0 - 0x0
      13'hBCC: dout <= 8'b10011110; // 3020 : 158 - 0x9e
      13'hBCD: dout <= 8'b11011100; // 3021 : 220 - 0xdc
      13'hBCE: dout <= 8'b10011010; // 3022 : 154 - 0x9a
      13'hBCF: dout <= 8'b00000000; // 3023 :   0 - 0x0
      13'hBD0: dout <= 8'b00000000; // 3024 :   0 - 0x0 -- Sprite 0xbd
      13'hBD1: dout <= 8'b00000000; // 3025 :   0 - 0x0
      13'hBD2: dout <= 8'b00000000; // 3026 :   0 - 0x0
      13'hBD3: dout <= 8'b00000000; // 3027 :   0 - 0x0
      13'hBD4: dout <= 8'b00000000; // 3028 :   0 - 0x0
      13'hBD5: dout <= 8'b00000000; // 3029 :   0 - 0x0
      13'hBD6: dout <= 8'b00000000; // 3030 :   0 - 0x0
      13'hBD7: dout <= 8'b00000000; // 3031 :   0 - 0x0
      13'hBD8: dout <= 8'b00000000; // 3032 :   0 - 0x0
      13'hBD9: dout <= 8'b00000000; // 3033 :   0 - 0x0
      13'hBDA: dout <= 8'b00000000; // 3034 :   0 - 0x0
      13'hBDB: dout <= 8'b00000000; // 3035 :   0 - 0x0
      13'hBDC: dout <= 8'b00000000; // 3036 :   0 - 0x0
      13'hBDD: dout <= 8'b00000000; // 3037 :   0 - 0x0
      13'hBDE: dout <= 8'b00000000; // 3038 :   0 - 0x0
      13'hBDF: dout <= 8'b00000000; // 3039 :   0 - 0x0
      13'hBE0: dout <= 8'b00000000; // 3040 :   0 - 0x0 -- Sprite 0xbe
      13'hBE1: dout <= 8'b00000000; // 3041 :   0 - 0x0
      13'hBE2: dout <= 8'b00000000; // 3042 :   0 - 0x0
      13'hBE3: dout <= 8'b00000000; // 3043 :   0 - 0x0
      13'hBE4: dout <= 8'b00000000; // 3044 :   0 - 0x0
      13'hBE5: dout <= 8'b00000000; // 3045 :   0 - 0x0
      13'hBE6: dout <= 8'b00000000; // 3046 :   0 - 0x0
      13'hBE7: dout <= 8'b00000000; // 3047 :   0 - 0x0
      13'hBE8: dout <= 8'b00000000; // 3048 :   0 - 0x0
      13'hBE9: dout <= 8'b00000000; // 3049 :   0 - 0x0
      13'hBEA: dout <= 8'b00000000; // 3050 :   0 - 0x0
      13'hBEB: dout <= 8'b00000000; // 3051 :   0 - 0x0
      13'hBEC: dout <= 8'b00000000; // 3052 :   0 - 0x0
      13'hBED: dout <= 8'b00000000; // 3053 :   0 - 0x0
      13'hBEE: dout <= 8'b00000000; // 3054 :   0 - 0x0
      13'hBEF: dout <= 8'b00000000; // 3055 :   0 - 0x0
      13'hBF0: dout <= 8'b00000000; // 3056 :   0 - 0x0 -- Sprite 0xbf
      13'hBF1: dout <= 8'b00000000; // 3057 :   0 - 0x0
      13'hBF2: dout <= 8'b00000000; // 3058 :   0 - 0x0
      13'hBF3: dout <= 8'b00000000; // 3059 :   0 - 0x0
      13'hBF4: dout <= 8'b00000000; // 3060 :   0 - 0x0
      13'hBF5: dout <= 8'b00000000; // 3061 :   0 - 0x0
      13'hBF6: dout <= 8'b00000000; // 3062 :   0 - 0x0
      13'hBF7: dout <= 8'b00000000; // 3063 :   0 - 0x0
      13'hBF8: dout <= 8'b00000000; // 3064 :   0 - 0x0
      13'hBF9: dout <= 8'b00000000; // 3065 :   0 - 0x0
      13'hBFA: dout <= 8'b00000000; // 3066 :   0 - 0x0
      13'hBFB: dout <= 8'b00000000; // 3067 :   0 - 0x0
      13'hBFC: dout <= 8'b00000000; // 3068 :   0 - 0x0
      13'hBFD: dout <= 8'b00000000; // 3069 :   0 - 0x0
      13'hBFE: dout <= 8'b00000000; // 3070 :   0 - 0x0
      13'hBFF: dout <= 8'b00000000; // 3071 :   0 - 0x0
      13'hC00: dout <= 8'b00000000; // 3072 :   0 - 0x0 -- Sprite 0xc0
      13'hC01: dout <= 8'b00000000; // 3073 :   0 - 0x0
      13'hC02: dout <= 8'b00000000; // 3074 :   0 - 0x0
      13'hC03: dout <= 8'b00000000; // 3075 :   0 - 0x0
      13'hC04: dout <= 8'b00000000; // 3076 :   0 - 0x0
      13'hC05: dout <= 8'b00000000; // 3077 :   0 - 0x0
      13'hC06: dout <= 8'b00000000; // 3078 :   0 - 0x0
      13'hC07: dout <= 8'b00000000; // 3079 :   0 - 0x0
      13'hC08: dout <= 8'b00000000; // 3080 :   0 - 0x0
      13'hC09: dout <= 8'b00000000; // 3081 :   0 - 0x0
      13'hC0A: dout <= 8'b00000000; // 3082 :   0 - 0x0
      13'hC0B: dout <= 8'b00000000; // 3083 :   0 - 0x0
      13'hC0C: dout <= 8'b00000000; // 3084 :   0 - 0x0
      13'hC0D: dout <= 8'b00000000; // 3085 :   0 - 0x0
      13'hC0E: dout <= 8'b00000000; // 3086 :   0 - 0x0
      13'hC0F: dout <= 8'b00000000; // 3087 :   0 - 0x0
      13'hC10: dout <= 8'b00000000; // 3088 :   0 - 0x0 -- Sprite 0xc1
      13'hC11: dout <= 8'b00000000; // 3089 :   0 - 0x0
      13'hC12: dout <= 8'b00000000; // 3090 :   0 - 0x0
      13'hC13: dout <= 8'b00000000; // 3091 :   0 - 0x0
      13'hC14: dout <= 8'b00000000; // 3092 :   0 - 0x0
      13'hC15: dout <= 8'b00000000; // 3093 :   0 - 0x0
      13'hC16: dout <= 8'b00000000; // 3094 :   0 - 0x0
      13'hC17: dout <= 8'b00000000; // 3095 :   0 - 0x0
      13'hC18: dout <= 8'b00000000; // 3096 :   0 - 0x0
      13'hC19: dout <= 8'b00000000; // 3097 :   0 - 0x0
      13'hC1A: dout <= 8'b00000000; // 3098 :   0 - 0x0
      13'hC1B: dout <= 8'b00000000; // 3099 :   0 - 0x0
      13'hC1C: dout <= 8'b00000000; // 3100 :   0 - 0x0
      13'hC1D: dout <= 8'b00000000; // 3101 :   0 - 0x0
      13'hC1E: dout <= 8'b00000000; // 3102 :   0 - 0x0
      13'hC1F: dout <= 8'b00000000; // 3103 :   0 - 0x0
      13'hC20: dout <= 8'b00000000; // 3104 :   0 - 0x0 -- Sprite 0xc2
      13'hC21: dout <= 8'b00000000; // 3105 :   0 - 0x0
      13'hC22: dout <= 8'b00000000; // 3106 :   0 - 0x0
      13'hC23: dout <= 8'b00000000; // 3107 :   0 - 0x0
      13'hC24: dout <= 8'b00000000; // 3108 :   0 - 0x0
      13'hC25: dout <= 8'b00000000; // 3109 :   0 - 0x0
      13'hC26: dout <= 8'b00000000; // 3110 :   0 - 0x0
      13'hC27: dout <= 8'b00000000; // 3111 :   0 - 0x0
      13'hC28: dout <= 8'b00000000; // 3112 :   0 - 0x0
      13'hC29: dout <= 8'b00000000; // 3113 :   0 - 0x0
      13'hC2A: dout <= 8'b00000000; // 3114 :   0 - 0x0
      13'hC2B: dout <= 8'b00000000; // 3115 :   0 - 0x0
      13'hC2C: dout <= 8'b00000000; // 3116 :   0 - 0x0
      13'hC2D: dout <= 8'b00000000; // 3117 :   0 - 0x0
      13'hC2E: dout <= 8'b00000000; // 3118 :   0 - 0x0
      13'hC2F: dout <= 8'b00000000; // 3119 :   0 - 0x0
      13'hC30: dout <= 8'b00000000; // 3120 :   0 - 0x0 -- Sprite 0xc3
      13'hC31: dout <= 8'b00000000; // 3121 :   0 - 0x0
      13'hC32: dout <= 8'b00000000; // 3122 :   0 - 0x0
      13'hC33: dout <= 8'b00000000; // 3123 :   0 - 0x0
      13'hC34: dout <= 8'b00000000; // 3124 :   0 - 0x0
      13'hC35: dout <= 8'b00000000; // 3125 :   0 - 0x0
      13'hC36: dout <= 8'b00000000; // 3126 :   0 - 0x0
      13'hC37: dout <= 8'b00000000; // 3127 :   0 - 0x0
      13'hC38: dout <= 8'b00000000; // 3128 :   0 - 0x0
      13'hC39: dout <= 8'b00000000; // 3129 :   0 - 0x0
      13'hC3A: dout <= 8'b00000000; // 3130 :   0 - 0x0
      13'hC3B: dout <= 8'b00000000; // 3131 :   0 - 0x0
      13'hC3C: dout <= 8'b00000000; // 3132 :   0 - 0x0
      13'hC3D: dout <= 8'b00000000; // 3133 :   0 - 0x0
      13'hC3E: dout <= 8'b00000000; // 3134 :   0 - 0x0
      13'hC3F: dout <= 8'b00000000; // 3135 :   0 - 0x0
      13'hC40: dout <= 8'b00000000; // 3136 :   0 - 0x0 -- Sprite 0xc4
      13'hC41: dout <= 8'b00000000; // 3137 :   0 - 0x0
      13'hC42: dout <= 8'b00000000; // 3138 :   0 - 0x0
      13'hC43: dout <= 8'b00000000; // 3139 :   0 - 0x0
      13'hC44: dout <= 8'b00000000; // 3140 :   0 - 0x0
      13'hC45: dout <= 8'b00000000; // 3141 :   0 - 0x0
      13'hC46: dout <= 8'b00000000; // 3142 :   0 - 0x0
      13'hC47: dout <= 8'b00000000; // 3143 :   0 - 0x0
      13'hC48: dout <= 8'b00000000; // 3144 :   0 - 0x0
      13'hC49: dout <= 8'b00000000; // 3145 :   0 - 0x0
      13'hC4A: dout <= 8'b00000000; // 3146 :   0 - 0x0
      13'hC4B: dout <= 8'b00000000; // 3147 :   0 - 0x0
      13'hC4C: dout <= 8'b00000000; // 3148 :   0 - 0x0
      13'hC4D: dout <= 8'b00000000; // 3149 :   0 - 0x0
      13'hC4E: dout <= 8'b00000000; // 3150 :   0 - 0x0
      13'hC4F: dout <= 8'b00000000; // 3151 :   0 - 0x0
      13'hC50: dout <= 8'b00000000; // 3152 :   0 - 0x0 -- Sprite 0xc5
      13'hC51: dout <= 8'b00000000; // 3153 :   0 - 0x0
      13'hC52: dout <= 8'b00000001; // 3154 :   1 - 0x1
      13'hC53: dout <= 8'b00000110; // 3155 :   6 - 0x6
      13'hC54: dout <= 8'b00001010; // 3156 :  10 - 0xa
      13'hC55: dout <= 8'b00010100; // 3157 :  20 - 0x14
      13'hC56: dout <= 8'b00010000; // 3158 :  16 - 0x10
      13'hC57: dout <= 8'b00101000; // 3159 :  40 - 0x28
      13'hC58: dout <= 8'b00000000; // 3160 :   0 - 0x0
      13'hC59: dout <= 8'b00000000; // 3161 :   0 - 0x0
      13'hC5A: dout <= 8'b00000000; // 3162 :   0 - 0x0
      13'hC5B: dout <= 8'b00000001; // 3163 :   1 - 0x1
      13'hC5C: dout <= 8'b00000111; // 3164 :   7 - 0x7
      13'hC5D: dout <= 8'b00001111; // 3165 :  15 - 0xf
      13'hC5E: dout <= 8'b00001111; // 3166 :  15 - 0xf
      13'hC5F: dout <= 8'b00011111; // 3167 :  31 - 0x1f
      13'hC60: dout <= 8'b00011111; // 3168 :  31 - 0x1f -- Sprite 0xc6
      13'hC61: dout <= 8'b01100000; // 3169 :  96 - 0x60
      13'hC62: dout <= 8'b10100000; // 3170 : 160 - 0xa0
      13'hC63: dout <= 8'b01000000; // 3171 :  64 - 0x40
      13'hC64: dout <= 8'b00000000; // 3172 :   0 - 0x0
      13'hC65: dout <= 8'b00000000; // 3173 :   0 - 0x0
      13'hC66: dout <= 8'b00000000; // 3174 :   0 - 0x0
      13'hC67: dout <= 8'b00000000; // 3175 :   0 - 0x0
      13'hC68: dout <= 8'b00000000; // 3176 :   0 - 0x0
      13'hC69: dout <= 8'b00011111; // 3177 :  31 - 0x1f
      13'hC6A: dout <= 8'b01111111; // 3178 : 127 - 0x7f
      13'hC6B: dout <= 8'b11111111; // 3179 : 255 - 0xff
      13'hC6C: dout <= 8'b11111111; // 3180 : 255 - 0xff
      13'hC6D: dout <= 8'b11111111; // 3181 : 255 - 0xff
      13'hC6E: dout <= 8'b11111111; // 3182 : 255 - 0xff
      13'hC6F: dout <= 8'b11111111; // 3183 : 255 - 0xff
      13'hC70: dout <= 8'b00110000; // 3184 :  48 - 0x30 -- Sprite 0xc7
      13'hC71: dout <= 8'b01000000; // 3185 :  64 - 0x40
      13'hC72: dout <= 8'b01100000; // 3186 :  96 - 0x60
      13'hC73: dout <= 8'b11000000; // 3187 : 192 - 0xc0
      13'hC74: dout <= 8'b10000000; // 3188 : 128 - 0x80
      13'hC75: dout <= 8'b10100000; // 3189 : 160 - 0xa0
      13'hC76: dout <= 8'b11000000; // 3190 : 192 - 0xc0
      13'hC77: dout <= 8'b10000000; // 3191 : 128 - 0x80
      13'hC78: dout <= 8'b00011111; // 3192 :  31 - 0x1f
      13'hC79: dout <= 8'b00111111; // 3193 :  63 - 0x3f
      13'hC7A: dout <= 8'b00111111; // 3194 :  63 - 0x3f
      13'hC7B: dout <= 8'b01111111; // 3195 : 127 - 0x7f
      13'hC7C: dout <= 8'b01111111; // 3196 : 127 - 0x7f
      13'hC7D: dout <= 8'b01111111; // 3197 : 127 - 0x7f
      13'hC7E: dout <= 8'b01111111; // 3198 : 127 - 0x7f
      13'hC7F: dout <= 8'b01111111; // 3199 : 127 - 0x7f
      13'hC80: dout <= 8'b11111111; // 3200 : 255 - 0xff -- Sprite 0xc8
      13'hC81: dout <= 8'b00000000; // 3201 :   0 - 0x0
      13'hC82: dout <= 8'b00000000; // 3202 :   0 - 0x0
      13'hC83: dout <= 8'b00000000; // 3203 :   0 - 0x0
      13'hC84: dout <= 8'b00000000; // 3204 :   0 - 0x0
      13'hC85: dout <= 8'b00000000; // 3205 :   0 - 0x0
      13'hC86: dout <= 8'b00000000; // 3206 :   0 - 0x0
      13'hC87: dout <= 8'b00000000; // 3207 :   0 - 0x0
      13'hC88: dout <= 8'b00000000; // 3208 :   0 - 0x0
      13'hC89: dout <= 8'b11111111; // 3209 : 255 - 0xff
      13'hC8A: dout <= 8'b11111111; // 3210 : 255 - 0xff
      13'hC8B: dout <= 8'b11111111; // 3211 : 255 - 0xff
      13'hC8C: dout <= 8'b11111111; // 3212 : 255 - 0xff
      13'hC8D: dout <= 8'b11111111; // 3213 : 255 - 0xff
      13'hC8E: dout <= 8'b11111111; // 3214 : 255 - 0xff
      13'hC8F: dout <= 8'b11111111; // 3215 : 255 - 0xff
      13'hC90: dout <= 8'b00010100; // 3216 :  20 - 0x14 -- Sprite 0xc9
      13'hC91: dout <= 8'b00101010; // 3217 :  42 - 0x2a
      13'hC92: dout <= 8'b00010110; // 3218 :  22 - 0x16
      13'hC93: dout <= 8'b00101011; // 3219 :  43 - 0x2b
      13'hC94: dout <= 8'b00010101; // 3220 :  21 - 0x15
      13'hC95: dout <= 8'b00101011; // 3221 :  43 - 0x2b
      13'hC96: dout <= 8'b00010101; // 3222 :  21 - 0x15
      13'hC97: dout <= 8'b00101011; // 3223 :  43 - 0x2b
      13'hC98: dout <= 8'b11101000; // 3224 : 232 - 0xe8
      13'hC99: dout <= 8'b11010100; // 3225 : 212 - 0xd4
      13'hC9A: dout <= 8'b11101000; // 3226 : 232 - 0xe8
      13'hC9B: dout <= 8'b11010100; // 3227 : 212 - 0xd4
      13'hC9C: dout <= 8'b11101010; // 3228 : 234 - 0xea
      13'hC9D: dout <= 8'b11010100; // 3229 : 212 - 0xd4
      13'hC9E: dout <= 8'b11101010; // 3230 : 234 - 0xea
      13'hC9F: dout <= 8'b11010100; // 3231 : 212 - 0xd4
      13'hCA0: dout <= 8'b00000000; // 3232 :   0 - 0x0 -- Sprite 0xca
      13'hCA1: dout <= 8'b00000100; // 3233 :   4 - 0x4
      13'hCA2: dout <= 8'b00000100; // 3234 :   4 - 0x4
      13'hCA3: dout <= 8'b00000101; // 3235 :   5 - 0x5
      13'hCA4: dout <= 8'b00010101; // 3236 :  21 - 0x15
      13'hCA5: dout <= 8'b00010101; // 3237 :  21 - 0x15
      13'hCA6: dout <= 8'b01010101; // 3238 :  85 - 0x55
      13'hCA7: dout <= 8'b01010101; // 3239 :  85 - 0x55
      13'hCA8: dout <= 8'b00000000; // 3240 :   0 - 0x0
      13'hCA9: dout <= 8'b00000000; // 3241 :   0 - 0x0
      13'hCAA: dout <= 8'b00000000; // 3242 :   0 - 0x0
      13'hCAB: dout <= 8'b00000000; // 3243 :   0 - 0x0
      13'hCAC: dout <= 8'b00000000; // 3244 :   0 - 0x0
      13'hCAD: dout <= 8'b00000000; // 3245 :   0 - 0x0
      13'hCAE: dout <= 8'b00000000; // 3246 :   0 - 0x0
      13'hCAF: dout <= 8'b00000000; // 3247 :   0 - 0x0
      13'hCB0: dout <= 8'b00000000; // 3248 :   0 - 0x0 -- Sprite 0xcb
      13'hCB1: dout <= 8'b00000000; // 3249 :   0 - 0x0
      13'hCB2: dout <= 8'b00010000; // 3250 :  16 - 0x10
      13'hCB3: dout <= 8'b00010000; // 3251 :  16 - 0x10
      13'hCB4: dout <= 8'b01010001; // 3252 :  81 - 0x51
      13'hCB5: dout <= 8'b01010101; // 3253 :  85 - 0x55
      13'hCB6: dout <= 8'b01010101; // 3254 :  85 - 0x55
      13'hCB7: dout <= 8'b01010101; // 3255 :  85 - 0x55
      13'hCB8: dout <= 8'b00000000; // 3256 :   0 - 0x0
      13'hCB9: dout <= 8'b00000000; // 3257 :   0 - 0x0
      13'hCBA: dout <= 8'b00000000; // 3258 :   0 - 0x0
      13'hCBB: dout <= 8'b00000000; // 3259 :   0 - 0x0
      13'hCBC: dout <= 8'b00000000; // 3260 :   0 - 0x0
      13'hCBD: dout <= 8'b00000000; // 3261 :   0 - 0x0
      13'hCBE: dout <= 8'b00000000; // 3262 :   0 - 0x0
      13'hCBF: dout <= 8'b00000000; // 3263 :   0 - 0x0
      13'hCC0: dout <= 8'b00000000; // 3264 :   0 - 0x0 -- Sprite 0xcc
      13'hCC1: dout <= 8'b00000000; // 3265 :   0 - 0x0
      13'hCC2: dout <= 8'b00000000; // 3266 :   0 - 0x0
      13'hCC3: dout <= 8'b00000101; // 3267 :   5 - 0x5
      13'hCC4: dout <= 8'b00001111; // 3268 :  15 - 0xf
      13'hCC5: dout <= 8'b00000111; // 3269 :   7 - 0x7
      13'hCC6: dout <= 8'b00000011; // 3270 :   3 - 0x3
      13'hCC7: dout <= 8'b00000001; // 3271 :   1 - 0x1
      13'hCC8: dout <= 8'b00000000; // 3272 :   0 - 0x0
      13'hCC9: dout <= 8'b00000000; // 3273 :   0 - 0x0
      13'hCCA: dout <= 8'b00000000; // 3274 :   0 - 0x0
      13'hCCB: dout <= 8'b00000000; // 3275 :   0 - 0x0
      13'hCCC: dout <= 8'b00000101; // 3276 :   5 - 0x5
      13'hCCD: dout <= 8'b00000010; // 3277 :   2 - 0x2
      13'hCCE: dout <= 8'b00000001; // 3278 :   1 - 0x1
      13'hCCF: dout <= 8'b00000000; // 3279 :   0 - 0x0
      13'hCD0: dout <= 8'b00000000; // 3280 :   0 - 0x0 -- Sprite 0xcd
      13'hCD1: dout <= 8'b00000000; // 3281 :   0 - 0x0
      13'hCD2: dout <= 8'b10000000; // 3282 : 128 - 0x80
      13'hCD3: dout <= 8'b11010000; // 3283 : 208 - 0xd0
      13'hCD4: dout <= 8'b11111000; // 3284 : 248 - 0xf8
      13'hCD5: dout <= 8'b11110000; // 3285 : 240 - 0xf0
      13'hCD6: dout <= 8'b11100000; // 3286 : 224 - 0xe0
      13'hCD7: dout <= 8'b11000000; // 3287 : 192 - 0xc0
      13'hCD8: dout <= 8'b00000000; // 3288 :   0 - 0x0
      13'hCD9: dout <= 8'b00000000; // 3289 :   0 - 0x0
      13'hCDA: dout <= 8'b00000000; // 3290 :   0 - 0x0
      13'hCDB: dout <= 8'b10000000; // 3291 : 128 - 0x80
      13'hCDC: dout <= 8'b01010000; // 3292 :  80 - 0x50
      13'hCDD: dout <= 8'b10100000; // 3293 : 160 - 0xa0
      13'hCDE: dout <= 8'b01000000; // 3294 :  64 - 0x40
      13'hCDF: dout <= 8'b10000000; // 3295 : 128 - 0x80
      13'hCE0: dout <= 8'b00000000; // 3296 :   0 - 0x0 -- Sprite 0xce
      13'hCE1: dout <= 8'b00000000; // 3297 :   0 - 0x0
      13'hCE2: dout <= 8'b00000000; // 3298 :   0 - 0x0
      13'hCE3: dout <= 8'b01111000; // 3299 : 120 - 0x78
      13'hCE4: dout <= 8'b11001111; // 3300 : 207 - 0xcf
      13'hCE5: dout <= 8'b10000000; // 3301 : 128 - 0x80
      13'hCE6: dout <= 8'b11001111; // 3302 : 207 - 0xcf
      13'hCE7: dout <= 8'b01001000; // 3303 :  72 - 0x48
      13'hCE8: dout <= 8'b00000000; // 3304 :   0 - 0x0
      13'hCE9: dout <= 8'b00000000; // 3305 :   0 - 0x0
      13'hCEA: dout <= 8'b00000000; // 3306 :   0 - 0x0
      13'hCEB: dout <= 8'b00000000; // 3307 :   0 - 0x0
      13'hCEC: dout <= 8'b00110000; // 3308 :  48 - 0x30
      13'hCED: dout <= 8'b01111111; // 3309 : 127 - 0x7f
      13'hCEE: dout <= 8'b00110000; // 3310 :  48 - 0x30
      13'hCEF: dout <= 8'b00110000; // 3311 :  48 - 0x30
      13'hCF0: dout <= 8'b00000000; // 3312 :   0 - 0x0 -- Sprite 0xcf
      13'hCF1: dout <= 8'b00000000; // 3313 :   0 - 0x0
      13'hCF2: dout <= 8'b00000000; // 3314 :   0 - 0x0
      13'hCF3: dout <= 8'b00011110; // 3315 :  30 - 0x1e
      13'hCF4: dout <= 8'b11110011; // 3316 : 243 - 0xf3
      13'hCF5: dout <= 8'b00000001; // 3317 :   1 - 0x1
      13'hCF6: dout <= 8'b11110011; // 3318 : 243 - 0xf3
      13'hCF7: dout <= 8'b00010010; // 3319 :  18 - 0x12
      13'hCF8: dout <= 8'b00000000; // 3320 :   0 - 0x0
      13'hCF9: dout <= 8'b00000000; // 3321 :   0 - 0x0
      13'hCFA: dout <= 8'b00000000; // 3322 :   0 - 0x0
      13'hCFB: dout <= 8'b00000000; // 3323 :   0 - 0x0
      13'hCFC: dout <= 8'b00001100; // 3324 :  12 - 0xc
      13'hCFD: dout <= 8'b11111110; // 3325 : 254 - 0xfe
      13'hCFE: dout <= 8'b00001100; // 3326 :  12 - 0xc
      13'hCFF: dout <= 8'b00001100; // 3327 :  12 - 0xc
      13'hD00: dout <= 8'b00000000; // 3328 :   0 - 0x0 -- Sprite 0xd0
      13'hD01: dout <= 8'b00000000; // 3329 :   0 - 0x0
      13'hD02: dout <= 8'b00000000; // 3330 :   0 - 0x0
      13'hD03: dout <= 8'b00000000; // 3331 :   0 - 0x0
      13'hD04: dout <= 8'b00000000; // 3332 :   0 - 0x0
      13'hD05: dout <= 8'b00000000; // 3333 :   0 - 0x0
      13'hD06: dout <= 8'b00000000; // 3334 :   0 - 0x0
      13'hD07: dout <= 8'b00000000; // 3335 :   0 - 0x0
      13'hD08: dout <= 8'b00000000; // 3336 :   0 - 0x0
      13'hD09: dout <= 8'b00000000; // 3337 :   0 - 0x0
      13'hD0A: dout <= 8'b00000000; // 3338 :   0 - 0x0
      13'hD0B: dout <= 8'b00000000; // 3339 :   0 - 0x0
      13'hD0C: dout <= 8'b00000000; // 3340 :   0 - 0x0
      13'hD0D: dout <= 8'b00000000; // 3341 :   0 - 0x0
      13'hD0E: dout <= 8'b00000000; // 3342 :   0 - 0x0
      13'hD0F: dout <= 8'b00000000; // 3343 :   0 - 0x0
      13'hD10: dout <= 8'b00000000; // 3344 :   0 - 0x0 -- Sprite 0xd1
      13'hD11: dout <= 8'b00000000; // 3345 :   0 - 0x0
      13'hD12: dout <= 8'b00000000; // 3346 :   0 - 0x0
      13'hD13: dout <= 8'b00000000; // 3347 :   0 - 0x0
      13'hD14: dout <= 8'b00000000; // 3348 :   0 - 0x0
      13'hD15: dout <= 8'b00000000; // 3349 :   0 - 0x0
      13'hD16: dout <= 8'b00000000; // 3350 :   0 - 0x0
      13'hD17: dout <= 8'b00000000; // 3351 :   0 - 0x0
      13'hD18: dout <= 8'b00000000; // 3352 :   0 - 0x0
      13'hD19: dout <= 8'b00000000; // 3353 :   0 - 0x0
      13'hD1A: dout <= 8'b00000000; // 3354 :   0 - 0x0
      13'hD1B: dout <= 8'b00000000; // 3355 :   0 - 0x0
      13'hD1C: dout <= 8'b00000000; // 3356 :   0 - 0x0
      13'hD1D: dout <= 8'b00000000; // 3357 :   0 - 0x0
      13'hD1E: dout <= 8'b00000000; // 3358 :   0 - 0x0
      13'hD1F: dout <= 8'b00000000; // 3359 :   0 - 0x0
      13'hD20: dout <= 8'b00001000; // 3360 :   8 - 0x8 -- Sprite 0xd2
      13'hD21: dout <= 8'b00001100; // 3361 :  12 - 0xc
      13'hD22: dout <= 8'b00001000; // 3362 :   8 - 0x8
      13'hD23: dout <= 8'b00001000; // 3363 :   8 - 0x8
      13'hD24: dout <= 8'b00001010; // 3364 :  10 - 0xa
      13'hD25: dout <= 8'b00001000; // 3365 :   8 - 0x8
      13'hD26: dout <= 8'b00001000; // 3366 :   8 - 0x8
      13'hD27: dout <= 8'b00001100; // 3367 :  12 - 0xc
      13'hD28: dout <= 8'b00000111; // 3368 :   7 - 0x7
      13'hD29: dout <= 8'b00000111; // 3369 :   7 - 0x7
      13'hD2A: dout <= 8'b00000111; // 3370 :   7 - 0x7
      13'hD2B: dout <= 8'b00000111; // 3371 :   7 - 0x7
      13'hD2C: dout <= 8'b00000111; // 3372 :   7 - 0x7
      13'hD2D: dout <= 8'b00000111; // 3373 :   7 - 0x7
      13'hD2E: dout <= 8'b00000111; // 3374 :   7 - 0x7
      13'hD2F: dout <= 8'b00000111; // 3375 :   7 - 0x7
      13'hD30: dout <= 8'b00010000; // 3376 :  16 - 0x10 -- Sprite 0xd3
      13'hD31: dout <= 8'b00010000; // 3377 :  16 - 0x10
      13'hD32: dout <= 8'b00110000; // 3378 :  48 - 0x30
      13'hD33: dout <= 8'b00010000; // 3379 :  16 - 0x10
      13'hD34: dout <= 8'b01010000; // 3380 :  80 - 0x50
      13'hD35: dout <= 8'b00010000; // 3381 :  16 - 0x10
      13'hD36: dout <= 8'b00110000; // 3382 :  48 - 0x30
      13'hD37: dout <= 8'b00010000; // 3383 :  16 - 0x10
      13'hD38: dout <= 8'b11100000; // 3384 : 224 - 0xe0
      13'hD39: dout <= 8'b11100000; // 3385 : 224 - 0xe0
      13'hD3A: dout <= 8'b11000000; // 3386 : 192 - 0xc0
      13'hD3B: dout <= 8'b11100000; // 3387 : 224 - 0xe0
      13'hD3C: dout <= 8'b10100000; // 3388 : 160 - 0xa0
      13'hD3D: dout <= 8'b11100000; // 3389 : 224 - 0xe0
      13'hD3E: dout <= 8'b11000000; // 3390 : 192 - 0xc0
      13'hD3F: dout <= 8'b11100000; // 3391 : 224 - 0xe0
      13'hD40: dout <= 8'b00000000; // 3392 :   0 - 0x0 -- Sprite 0xd4
      13'hD41: dout <= 8'b00000000; // 3393 :   0 - 0x0
      13'hD42: dout <= 8'b00000000; // 3394 :   0 - 0x0
      13'hD43: dout <= 8'b00000000; // 3395 :   0 - 0x0
      13'hD44: dout <= 8'b00000000; // 3396 :   0 - 0x0
      13'hD45: dout <= 8'b00000000; // 3397 :   0 - 0x0
      13'hD46: dout <= 8'b00000000; // 3398 :   0 - 0x0
      13'hD47: dout <= 8'b00000000; // 3399 :   0 - 0x0
      13'hD48: dout <= 8'b00000000; // 3400 :   0 - 0x0
      13'hD49: dout <= 8'b00000000; // 3401 :   0 - 0x0
      13'hD4A: dout <= 8'b00000000; // 3402 :   0 - 0x0
      13'hD4B: dout <= 8'b00000000; // 3403 :   0 - 0x0
      13'hD4C: dout <= 8'b00000000; // 3404 :   0 - 0x0
      13'hD4D: dout <= 8'b00000000; // 3405 :   0 - 0x0
      13'hD4E: dout <= 8'b00000000; // 3406 :   0 - 0x0
      13'hD4F: dout <= 8'b00000000; // 3407 :   0 - 0x0
      13'hD50: dout <= 8'b11111000; // 3408 : 248 - 0xf8 -- Sprite 0xd5
      13'hD51: dout <= 8'b00000110; // 3409 :   6 - 0x6
      13'hD52: dout <= 8'b00000001; // 3410 :   1 - 0x1
      13'hD53: dout <= 8'b00000000; // 3411 :   0 - 0x0
      13'hD54: dout <= 8'b00000000; // 3412 :   0 - 0x0
      13'hD55: dout <= 8'b00000000; // 3413 :   0 - 0x0
      13'hD56: dout <= 8'b00000000; // 3414 :   0 - 0x0
      13'hD57: dout <= 8'b00000000; // 3415 :   0 - 0x0
      13'hD58: dout <= 8'b00000000; // 3416 :   0 - 0x0
      13'hD59: dout <= 8'b11111000; // 3417 : 248 - 0xf8
      13'hD5A: dout <= 8'b11111110; // 3418 : 254 - 0xfe
      13'hD5B: dout <= 8'b11111111; // 3419 : 255 - 0xff
      13'hD5C: dout <= 8'b11111111; // 3420 : 255 - 0xff
      13'hD5D: dout <= 8'b11111111; // 3421 : 255 - 0xff
      13'hD5E: dout <= 8'b11111111; // 3422 : 255 - 0xff
      13'hD5F: dout <= 8'b11111111; // 3423 : 255 - 0xff
      13'hD60: dout <= 8'b00000000; // 3424 :   0 - 0x0 -- Sprite 0xd6
      13'hD61: dout <= 8'b00000000; // 3425 :   0 - 0x0
      13'hD62: dout <= 8'b10000000; // 3426 : 128 - 0x80
      13'hD63: dout <= 8'b01100000; // 3427 :  96 - 0x60
      13'hD64: dout <= 8'b01010000; // 3428 :  80 - 0x50
      13'hD65: dout <= 8'b10101000; // 3429 : 168 - 0xa8
      13'hD66: dout <= 8'b01011000; // 3430 :  88 - 0x58
      13'hD67: dout <= 8'b00101100; // 3431 :  44 - 0x2c
      13'hD68: dout <= 8'b00000000; // 3432 :   0 - 0x0
      13'hD69: dout <= 8'b00000000; // 3433 :   0 - 0x0
      13'hD6A: dout <= 8'b00000000; // 3434 :   0 - 0x0
      13'hD6B: dout <= 8'b10000000; // 3435 : 128 - 0x80
      13'hD6C: dout <= 8'b10100000; // 3436 : 160 - 0xa0
      13'hD6D: dout <= 8'b01010000; // 3437 :  80 - 0x50
      13'hD6E: dout <= 8'b10100000; // 3438 : 160 - 0xa0
      13'hD6F: dout <= 8'b11010000; // 3439 : 208 - 0xd0
      13'hD70: dout <= 8'b10100000; // 3440 : 160 - 0xa0 -- Sprite 0xd7
      13'hD71: dout <= 8'b11000000; // 3441 : 192 - 0xc0
      13'hD72: dout <= 8'b10000000; // 3442 : 128 - 0x80
      13'hD73: dout <= 8'b01010000; // 3443 :  80 - 0x50
      13'hD74: dout <= 8'b01100000; // 3444 :  96 - 0x60
      13'hD75: dout <= 8'b00111000; // 3445 :  56 - 0x38
      13'hD76: dout <= 8'b00001000; // 3446 :   8 - 0x8
      13'hD77: dout <= 8'b00000111; // 3447 :   7 - 0x7
      13'hD78: dout <= 8'b01111111; // 3448 : 127 - 0x7f
      13'hD79: dout <= 8'b01111111; // 3449 : 127 - 0x7f
      13'hD7A: dout <= 8'b01111111; // 3450 : 127 - 0x7f
      13'hD7B: dout <= 8'b00111111; // 3451 :  63 - 0x3f
      13'hD7C: dout <= 8'b00111111; // 3452 :  63 - 0x3f
      13'hD7D: dout <= 8'b00001111; // 3453 :  15 - 0xf
      13'hD7E: dout <= 8'b00000111; // 3454 :   7 - 0x7
      13'hD7F: dout <= 8'b00000000; // 3455 :   0 - 0x0
      13'hD80: dout <= 8'b00000000; // 3456 :   0 - 0x0 -- Sprite 0xd8
      13'hD81: dout <= 8'b00000000; // 3457 :   0 - 0x0
      13'hD82: dout <= 8'b00000000; // 3458 :   0 - 0x0
      13'hD83: dout <= 8'b00000000; // 3459 :   0 - 0x0
      13'hD84: dout <= 8'b00000000; // 3460 :   0 - 0x0
      13'hD85: dout <= 8'b00000000; // 3461 :   0 - 0x0
      13'hD86: dout <= 8'b00000000; // 3462 :   0 - 0x0
      13'hD87: dout <= 8'b11111111; // 3463 : 255 - 0xff
      13'hD88: dout <= 8'b11111111; // 3464 : 255 - 0xff
      13'hD89: dout <= 8'b11111111; // 3465 : 255 - 0xff
      13'hD8A: dout <= 8'b11111111; // 3466 : 255 - 0xff
      13'hD8B: dout <= 8'b11111111; // 3467 : 255 - 0xff
      13'hD8C: dout <= 8'b11111111; // 3468 : 255 - 0xff
      13'hD8D: dout <= 8'b11111111; // 3469 : 255 - 0xff
      13'hD8E: dout <= 8'b11111111; // 3470 : 255 - 0xff
      13'hD8F: dout <= 8'b00000000; // 3471 :   0 - 0x0
      13'hD90: dout <= 8'b00010101; // 3472 :  21 - 0x15 -- Sprite 0xd9
      13'hD91: dout <= 8'b00101011; // 3473 :  43 - 0x2b
      13'hD92: dout <= 8'b00010101; // 3474 :  21 - 0x15
      13'hD93: dout <= 8'b00101010; // 3475 :  42 - 0x2a
      13'hD94: dout <= 8'b01010110; // 3476 :  86 - 0x56
      13'hD95: dout <= 8'b10101100; // 3477 : 172 - 0xac
      13'hD96: dout <= 8'b01010000; // 3478 :  80 - 0x50
      13'hD97: dout <= 8'b11100000; // 3479 : 224 - 0xe0
      13'hD98: dout <= 8'b11101010; // 3480 : 234 - 0xea
      13'hD99: dout <= 8'b11010100; // 3481 : 212 - 0xd4
      13'hD9A: dout <= 8'b11101010; // 3482 : 234 - 0xea
      13'hD9B: dout <= 8'b11010100; // 3483 : 212 - 0xd4
      13'hD9C: dout <= 8'b10101000; // 3484 : 168 - 0xa8
      13'hD9D: dout <= 8'b01010000; // 3485 :  80 - 0x50
      13'hD9E: dout <= 8'b10100000; // 3486 : 160 - 0xa0
      13'hD9F: dout <= 8'b00000000; // 3487 :   0 - 0x0
      13'hDA0: dout <= 8'b00000001; // 3488 :   1 - 0x1 -- Sprite 0xda
      13'hDA1: dout <= 8'b00001101; // 3489 :  13 - 0xd
      13'hDA2: dout <= 8'b00010011; // 3490 :  19 - 0x13
      13'hDA3: dout <= 8'b00001101; // 3491 :  13 - 0xd
      13'hDA4: dout <= 8'b00000001; // 3492 :   1 - 0x1
      13'hDA5: dout <= 8'b00000001; // 3493 :   1 - 0x1
      13'hDA6: dout <= 8'b00000001; // 3494 :   1 - 0x1
      13'hDA7: dout <= 8'b00000001; // 3495 :   1 - 0x1
      13'hDA8: dout <= 8'b00000000; // 3496 :   0 - 0x0
      13'hDA9: dout <= 8'b00000000; // 3497 :   0 - 0x0
      13'hDAA: dout <= 8'b00001100; // 3498 :  12 - 0xc
      13'hDAB: dout <= 8'b00000000; // 3499 :   0 - 0x0
      13'hDAC: dout <= 8'b00000000; // 3500 :   0 - 0x0
      13'hDAD: dout <= 8'b00000000; // 3501 :   0 - 0x0
      13'hDAE: dout <= 8'b00000000; // 3502 :   0 - 0x0
      13'hDAF: dout <= 8'b00000000; // 3503 :   0 - 0x0
      13'hDB0: dout <= 8'b11000000; // 3504 : 192 - 0xc0 -- Sprite 0xdb
      13'hDB1: dout <= 8'b01000000; // 3505 :  64 - 0x40
      13'hDB2: dout <= 8'b01000000; // 3506 :  64 - 0x40
      13'hDB3: dout <= 8'b01011000; // 3507 :  88 - 0x58
      13'hDB4: dout <= 8'b01100100; // 3508 : 100 - 0x64
      13'hDB5: dout <= 8'b01011000; // 3509 :  88 - 0x58
      13'hDB6: dout <= 8'b01000000; // 3510 :  64 - 0x40
      13'hDB7: dout <= 8'b01000000; // 3511 :  64 - 0x40
      13'hDB8: dout <= 8'b00000000; // 3512 :   0 - 0x0
      13'hDB9: dout <= 8'b10000000; // 3513 : 128 - 0x80
      13'hDBA: dout <= 8'b10000000; // 3514 : 128 - 0x80
      13'hDBB: dout <= 8'b10000000; // 3515 : 128 - 0x80
      13'hDBC: dout <= 8'b10011000; // 3516 : 152 - 0x98
      13'hDBD: dout <= 8'b10000000; // 3517 : 128 - 0x80
      13'hDBE: dout <= 8'b10000000; // 3518 : 128 - 0x80
      13'hDBF: dout <= 8'b10000000; // 3519 : 128 - 0x80
      13'hDC0: dout <= 8'b00000000; // 3520 :   0 - 0x0 -- Sprite 0xdc
      13'hDC1: dout <= 8'b00000000; // 3521 :   0 - 0x0
      13'hDC2: dout <= 8'b00000000; // 3522 :   0 - 0x0
      13'hDC3: dout <= 8'b00000110; // 3523 :   6 - 0x6
      13'hDC4: dout <= 8'b00000111; // 3524 :   7 - 0x7
      13'hDC5: dout <= 8'b00000111; // 3525 :   7 - 0x7
      13'hDC6: dout <= 8'b00000111; // 3526 :   7 - 0x7
      13'hDC7: dout <= 8'b00000011; // 3527 :   3 - 0x3
      13'hDC8: dout <= 8'b00000000; // 3528 :   0 - 0x0
      13'hDC9: dout <= 8'b00000000; // 3529 :   0 - 0x0
      13'hDCA: dout <= 8'b00000000; // 3530 :   0 - 0x0
      13'hDCB: dout <= 8'b00000000; // 3531 :   0 - 0x0
      13'hDCC: dout <= 8'b00000010; // 3532 :   2 - 0x2
      13'hDCD: dout <= 8'b00000011; // 3533 :   3 - 0x3
      13'hDCE: dout <= 8'b00000011; // 3534 :   3 - 0x3
      13'hDCF: dout <= 8'b00000001; // 3535 :   1 - 0x1
      13'hDD0: dout <= 8'b00000000; // 3536 :   0 - 0x0 -- Sprite 0xdd
      13'hDD1: dout <= 8'b00000000; // 3537 :   0 - 0x0
      13'hDD2: dout <= 8'b00000000; // 3538 :   0 - 0x0
      13'hDD3: dout <= 8'b10110000; // 3539 : 176 - 0xb0
      13'hDD4: dout <= 8'b11110000; // 3540 : 240 - 0xf0
      13'hDD5: dout <= 8'b11110000; // 3541 : 240 - 0xf0
      13'hDD6: dout <= 8'b11110000; // 3542 : 240 - 0xf0
      13'hDD7: dout <= 8'b11100000; // 3543 : 224 - 0xe0
      13'hDD8: dout <= 8'b00000000; // 3544 :   0 - 0x0
      13'hDD9: dout <= 8'b00000000; // 3545 :   0 - 0x0
      13'hDDA: dout <= 8'b00000000; // 3546 :   0 - 0x0
      13'hDDB: dout <= 8'b00000000; // 3547 :   0 - 0x0
      13'hDDC: dout <= 8'b10100000; // 3548 : 160 - 0xa0
      13'hDDD: dout <= 8'b11100000; // 3549 : 224 - 0xe0
      13'hDDE: dout <= 8'b11100000; // 3550 : 224 - 0xe0
      13'hDDF: dout <= 8'b11000000; // 3551 : 192 - 0xc0
      13'hDE0: dout <= 8'b11001111; // 3552 : 207 - 0xcf -- Sprite 0xde
      13'hDE1: dout <= 8'b10000000; // 3553 : 128 - 0x80
      13'hDE2: dout <= 8'b11001111; // 3554 : 207 - 0xcf
      13'hDE3: dout <= 8'b01001000; // 3555 :  72 - 0x48
      13'hDE4: dout <= 8'b01001000; // 3556 :  72 - 0x48
      13'hDE5: dout <= 8'b01001000; // 3557 :  72 - 0x48
      13'hDE6: dout <= 8'b01001000; // 3558 :  72 - 0x48
      13'hDE7: dout <= 8'b01001000; // 3559 :  72 - 0x48
      13'hDE8: dout <= 8'b00110000; // 3560 :  48 - 0x30
      13'hDE9: dout <= 8'b01111111; // 3561 : 127 - 0x7f
      13'hDEA: dout <= 8'b00110000; // 3562 :  48 - 0x30
      13'hDEB: dout <= 8'b00110000; // 3563 :  48 - 0x30
      13'hDEC: dout <= 8'b00110000; // 3564 :  48 - 0x30
      13'hDED: dout <= 8'b00110000; // 3565 :  48 - 0x30
      13'hDEE: dout <= 8'b00110000; // 3566 :  48 - 0x30
      13'hDEF: dout <= 8'b00110000; // 3567 :  48 - 0x30
      13'hDF0: dout <= 8'b11110011; // 3568 : 243 - 0xf3 -- Sprite 0xdf
      13'hDF1: dout <= 8'b00000001; // 3569 :   1 - 0x1
      13'hDF2: dout <= 8'b11110011; // 3570 : 243 - 0xf3
      13'hDF3: dout <= 8'b00010010; // 3571 :  18 - 0x12
      13'hDF4: dout <= 8'b00010010; // 3572 :  18 - 0x12
      13'hDF5: dout <= 8'b00010010; // 3573 :  18 - 0x12
      13'hDF6: dout <= 8'b00010010; // 3574 :  18 - 0x12
      13'hDF7: dout <= 8'b00010010; // 3575 :  18 - 0x12
      13'hDF8: dout <= 8'b00001100; // 3576 :  12 - 0xc
      13'hDF9: dout <= 8'b11111110; // 3577 : 254 - 0xfe
      13'hDFA: dout <= 8'b00001100; // 3578 :  12 - 0xc
      13'hDFB: dout <= 8'b00001100; // 3579 :  12 - 0xc
      13'hDFC: dout <= 8'b00001100; // 3580 :  12 - 0xc
      13'hDFD: dout <= 8'b00001100; // 3581 :  12 - 0xc
      13'hDFE: dout <= 8'b00001100; // 3582 :  12 - 0xc
      13'hDFF: dout <= 8'b00001100; // 3583 :  12 - 0xc
      13'hE00: dout <= 8'b00000000; // 3584 :   0 - 0x0 -- Sprite 0xe0
      13'hE01: dout <= 8'b00000000; // 3585 :   0 - 0x0
      13'hE02: dout <= 8'b00000000; // 3586 :   0 - 0x0
      13'hE03: dout <= 8'b00000000; // 3587 :   0 - 0x0
      13'hE04: dout <= 8'b00000000; // 3588 :   0 - 0x0
      13'hE05: dout <= 8'b00000000; // 3589 :   0 - 0x0
      13'hE06: dout <= 8'b00000000; // 3590 :   0 - 0x0
      13'hE07: dout <= 8'b00000000; // 3591 :   0 - 0x0
      13'hE08: dout <= 8'b00000000; // 3592 :   0 - 0x0
      13'hE09: dout <= 8'b00000000; // 3593 :   0 - 0x0
      13'hE0A: dout <= 8'b00000000; // 3594 :   0 - 0x0
      13'hE0B: dout <= 8'b00000000; // 3595 :   0 - 0x0
      13'hE0C: dout <= 8'b00000000; // 3596 :   0 - 0x0
      13'hE0D: dout <= 8'b00000000; // 3597 :   0 - 0x0
      13'hE0E: dout <= 8'b00000000; // 3598 :   0 - 0x0
      13'hE0F: dout <= 8'b00000000; // 3599 :   0 - 0x0
      13'hE10: dout <= 8'b00000000; // 3600 :   0 - 0x0 -- Sprite 0xe1
      13'hE11: dout <= 8'b00000000; // 3601 :   0 - 0x0
      13'hE12: dout <= 8'b00000000; // 3602 :   0 - 0x0
      13'hE13: dout <= 8'b00000000; // 3603 :   0 - 0x0
      13'hE14: dout <= 8'b00000000; // 3604 :   0 - 0x0
      13'hE15: dout <= 8'b00000000; // 3605 :   0 - 0x0
      13'hE16: dout <= 8'b00000000; // 3606 :   0 - 0x0
      13'hE17: dout <= 8'b00000000; // 3607 :   0 - 0x0
      13'hE18: dout <= 8'b00000000; // 3608 :   0 - 0x0
      13'hE19: dout <= 8'b00000000; // 3609 :   0 - 0x0
      13'hE1A: dout <= 8'b00000000; // 3610 :   0 - 0x0
      13'hE1B: dout <= 8'b00000000; // 3611 :   0 - 0x0
      13'hE1C: dout <= 8'b00000000; // 3612 :   0 - 0x0
      13'hE1D: dout <= 8'b00000000; // 3613 :   0 - 0x0
      13'hE1E: dout <= 8'b00000000; // 3614 :   0 - 0x0
      13'hE1F: dout <= 8'b00000000; // 3615 :   0 - 0x0
      13'hE20: dout <= 8'b00000000; // 3616 :   0 - 0x0 -- Sprite 0xe2
      13'hE21: dout <= 8'b00000000; // 3617 :   0 - 0x0
      13'hE22: dout <= 8'b00000000; // 3618 :   0 - 0x0
      13'hE23: dout <= 8'b00000000; // 3619 :   0 - 0x0
      13'hE24: dout <= 8'b00000000; // 3620 :   0 - 0x0
      13'hE25: dout <= 8'b00000000; // 3621 :   0 - 0x0
      13'hE26: dout <= 8'b00000000; // 3622 :   0 - 0x0
      13'hE27: dout <= 8'b00000000; // 3623 :   0 - 0x0
      13'hE28: dout <= 8'b00000000; // 3624 :   0 - 0x0
      13'hE29: dout <= 8'b00000000; // 3625 :   0 - 0x0
      13'hE2A: dout <= 8'b00000000; // 3626 :   0 - 0x0
      13'hE2B: dout <= 8'b00000000; // 3627 :   0 - 0x0
      13'hE2C: dout <= 8'b00000000; // 3628 :   0 - 0x0
      13'hE2D: dout <= 8'b00000000; // 3629 :   0 - 0x0
      13'hE2E: dout <= 8'b00000000; // 3630 :   0 - 0x0
      13'hE2F: dout <= 8'b00000000; // 3631 :   0 - 0x0
      13'hE30: dout <= 8'b00000000; // 3632 :   0 - 0x0 -- Sprite 0xe3
      13'hE31: dout <= 8'b00000000; // 3633 :   0 - 0x0
      13'hE32: dout <= 8'b00000000; // 3634 :   0 - 0x0
      13'hE33: dout <= 8'b00000000; // 3635 :   0 - 0x0
      13'hE34: dout <= 8'b00000000; // 3636 :   0 - 0x0
      13'hE35: dout <= 8'b00000000; // 3637 :   0 - 0x0
      13'hE36: dout <= 8'b00000000; // 3638 :   0 - 0x0
      13'hE37: dout <= 8'b00000000; // 3639 :   0 - 0x0
      13'hE38: dout <= 8'b00000000; // 3640 :   0 - 0x0
      13'hE39: dout <= 8'b00000000; // 3641 :   0 - 0x0
      13'hE3A: dout <= 8'b00000000; // 3642 :   0 - 0x0
      13'hE3B: dout <= 8'b00000000; // 3643 :   0 - 0x0
      13'hE3C: dout <= 8'b00000000; // 3644 :   0 - 0x0
      13'hE3D: dout <= 8'b00000000; // 3645 :   0 - 0x0
      13'hE3E: dout <= 8'b00000000; // 3646 :   0 - 0x0
      13'hE3F: dout <= 8'b00000000; // 3647 :   0 - 0x0
      13'hE40: dout <= 8'b00000000; // 3648 :   0 - 0x0 -- Sprite 0xe4
      13'hE41: dout <= 8'b00000000; // 3649 :   0 - 0x0
      13'hE42: dout <= 8'b00000000; // 3650 :   0 - 0x0
      13'hE43: dout <= 8'b00000000; // 3651 :   0 - 0x0
      13'hE44: dout <= 8'b00000000; // 3652 :   0 - 0x0
      13'hE45: dout <= 8'b00000000; // 3653 :   0 - 0x0
      13'hE46: dout <= 8'b00000000; // 3654 :   0 - 0x0
      13'hE47: dout <= 8'b00000000; // 3655 :   0 - 0x0
      13'hE48: dout <= 8'b00000000; // 3656 :   0 - 0x0
      13'hE49: dout <= 8'b00000000; // 3657 :   0 - 0x0
      13'hE4A: dout <= 8'b00000000; // 3658 :   0 - 0x0
      13'hE4B: dout <= 8'b00000000; // 3659 :   0 - 0x0
      13'hE4C: dout <= 8'b00000000; // 3660 :   0 - 0x0
      13'hE4D: dout <= 8'b00000000; // 3661 :   0 - 0x0
      13'hE4E: dout <= 8'b00000000; // 3662 :   0 - 0x0
      13'hE4F: dout <= 8'b00000000; // 3663 :   0 - 0x0
      13'hE50: dout <= 8'b00000000; // 3664 :   0 - 0x0 -- Sprite 0xe5
      13'hE51: dout <= 8'b00000000; // 3665 :   0 - 0x0
      13'hE52: dout <= 8'b00000000; // 3666 :   0 - 0x0
      13'hE53: dout <= 8'b00000000; // 3667 :   0 - 0x0
      13'hE54: dout <= 8'b00000000; // 3668 :   0 - 0x0
      13'hE55: dout <= 8'b00000000; // 3669 :   0 - 0x0
      13'hE56: dout <= 8'b00000000; // 3670 :   0 - 0x0
      13'hE57: dout <= 8'b00000000; // 3671 :   0 - 0x0
      13'hE58: dout <= 8'b00000000; // 3672 :   0 - 0x0
      13'hE59: dout <= 8'b00000000; // 3673 :   0 - 0x0
      13'hE5A: dout <= 8'b00000000; // 3674 :   0 - 0x0
      13'hE5B: dout <= 8'b00000000; // 3675 :   0 - 0x0
      13'hE5C: dout <= 8'b00000000; // 3676 :   0 - 0x0
      13'hE5D: dout <= 8'b00000000; // 3677 :   0 - 0x0
      13'hE5E: dout <= 8'b00000000; // 3678 :   0 - 0x0
      13'hE5F: dout <= 8'b00000000; // 3679 :   0 - 0x0
      13'hE60: dout <= 8'b00000000; // 3680 :   0 - 0x0 -- Sprite 0xe6
      13'hE61: dout <= 8'b00000000; // 3681 :   0 - 0x0
      13'hE62: dout <= 8'b00000000; // 3682 :   0 - 0x0
      13'hE63: dout <= 8'b00000000; // 3683 :   0 - 0x0
      13'hE64: dout <= 8'b00000000; // 3684 :   0 - 0x0
      13'hE65: dout <= 8'b00000000; // 3685 :   0 - 0x0
      13'hE66: dout <= 8'b00000000; // 3686 :   0 - 0x0
      13'hE67: dout <= 8'b00000000; // 3687 :   0 - 0x0
      13'hE68: dout <= 8'b00000000; // 3688 :   0 - 0x0
      13'hE69: dout <= 8'b00000000; // 3689 :   0 - 0x0
      13'hE6A: dout <= 8'b00000000; // 3690 :   0 - 0x0
      13'hE6B: dout <= 8'b00000000; // 3691 :   0 - 0x0
      13'hE6C: dout <= 8'b00000000; // 3692 :   0 - 0x0
      13'hE6D: dout <= 8'b00000000; // 3693 :   0 - 0x0
      13'hE6E: dout <= 8'b00000000; // 3694 :   0 - 0x0
      13'hE6F: dout <= 8'b00000000; // 3695 :   0 - 0x0
      13'hE70: dout <= 8'b00000000; // 3696 :   0 - 0x0 -- Sprite 0xe7
      13'hE71: dout <= 8'b00000000; // 3697 :   0 - 0x0
      13'hE72: dout <= 8'b00000000; // 3698 :   0 - 0x0
      13'hE73: dout <= 8'b00000000; // 3699 :   0 - 0x0
      13'hE74: dout <= 8'b00000000; // 3700 :   0 - 0x0
      13'hE75: dout <= 8'b00000000; // 3701 :   0 - 0x0
      13'hE76: dout <= 8'b00000000; // 3702 :   0 - 0x0
      13'hE77: dout <= 8'b00000000; // 3703 :   0 - 0x0
      13'hE78: dout <= 8'b00000000; // 3704 :   0 - 0x0
      13'hE79: dout <= 8'b00000000; // 3705 :   0 - 0x0
      13'hE7A: dout <= 8'b00000000; // 3706 :   0 - 0x0
      13'hE7B: dout <= 8'b00000000; // 3707 :   0 - 0x0
      13'hE7C: dout <= 8'b00000000; // 3708 :   0 - 0x0
      13'hE7D: dout <= 8'b00000000; // 3709 :   0 - 0x0
      13'hE7E: dout <= 8'b00000000; // 3710 :   0 - 0x0
      13'hE7F: dout <= 8'b00000000; // 3711 :   0 - 0x0
      13'hE80: dout <= 8'b00000000; // 3712 :   0 - 0x0 -- Sprite 0xe8
      13'hE81: dout <= 8'b00000000; // 3713 :   0 - 0x0
      13'hE82: dout <= 8'b00000000; // 3714 :   0 - 0x0
      13'hE83: dout <= 8'b00000000; // 3715 :   0 - 0x0
      13'hE84: dout <= 8'b00000000; // 3716 :   0 - 0x0
      13'hE85: dout <= 8'b00000000; // 3717 :   0 - 0x0
      13'hE86: dout <= 8'b00000000; // 3718 :   0 - 0x0
      13'hE87: dout <= 8'b00000000; // 3719 :   0 - 0x0
      13'hE88: dout <= 8'b00000000; // 3720 :   0 - 0x0
      13'hE89: dout <= 8'b00000000; // 3721 :   0 - 0x0
      13'hE8A: dout <= 8'b00000000; // 3722 :   0 - 0x0
      13'hE8B: dout <= 8'b00000000; // 3723 :   0 - 0x0
      13'hE8C: dout <= 8'b00000000; // 3724 :   0 - 0x0
      13'hE8D: dout <= 8'b00000000; // 3725 :   0 - 0x0
      13'hE8E: dout <= 8'b00000000; // 3726 :   0 - 0x0
      13'hE8F: dout <= 8'b00000000; // 3727 :   0 - 0x0
      13'hE90: dout <= 8'b00000000; // 3728 :   0 - 0x0 -- Sprite 0xe9
      13'hE91: dout <= 8'b00000000; // 3729 :   0 - 0x0
      13'hE92: dout <= 8'b00000000; // 3730 :   0 - 0x0
      13'hE93: dout <= 8'b00000000; // 3731 :   0 - 0x0
      13'hE94: dout <= 8'b00000000; // 3732 :   0 - 0x0
      13'hE95: dout <= 8'b00000000; // 3733 :   0 - 0x0
      13'hE96: dout <= 8'b00000000; // 3734 :   0 - 0x0
      13'hE97: dout <= 8'b00000000; // 3735 :   0 - 0x0
      13'hE98: dout <= 8'b00000000; // 3736 :   0 - 0x0
      13'hE99: dout <= 8'b00000000; // 3737 :   0 - 0x0
      13'hE9A: dout <= 8'b00000000; // 3738 :   0 - 0x0
      13'hE9B: dout <= 8'b00000000; // 3739 :   0 - 0x0
      13'hE9C: dout <= 8'b00000000; // 3740 :   0 - 0x0
      13'hE9D: dout <= 8'b00000000; // 3741 :   0 - 0x0
      13'hE9E: dout <= 8'b00000000; // 3742 :   0 - 0x0
      13'hE9F: dout <= 8'b00000000; // 3743 :   0 - 0x0
      13'hEA0: dout <= 8'b00000000; // 3744 :   0 - 0x0 -- Sprite 0xea
      13'hEA1: dout <= 8'b00000000; // 3745 :   0 - 0x0
      13'hEA2: dout <= 8'b00000000; // 3746 :   0 - 0x0
      13'hEA3: dout <= 8'b00000000; // 3747 :   0 - 0x0
      13'hEA4: dout <= 8'b00000000; // 3748 :   0 - 0x0
      13'hEA5: dout <= 8'b00000000; // 3749 :   0 - 0x0
      13'hEA6: dout <= 8'b00000000; // 3750 :   0 - 0x0
      13'hEA7: dout <= 8'b00000000; // 3751 :   0 - 0x0
      13'hEA8: dout <= 8'b00000000; // 3752 :   0 - 0x0
      13'hEA9: dout <= 8'b00000000; // 3753 :   0 - 0x0
      13'hEAA: dout <= 8'b00000000; // 3754 :   0 - 0x0
      13'hEAB: dout <= 8'b00000000; // 3755 :   0 - 0x0
      13'hEAC: dout <= 8'b00000000; // 3756 :   0 - 0x0
      13'hEAD: dout <= 8'b00000000; // 3757 :   0 - 0x0
      13'hEAE: dout <= 8'b00000000; // 3758 :   0 - 0x0
      13'hEAF: dout <= 8'b00000000; // 3759 :   0 - 0x0
      13'hEB0: dout <= 8'b00000000; // 3760 :   0 - 0x0 -- Sprite 0xeb
      13'hEB1: dout <= 8'b00000000; // 3761 :   0 - 0x0
      13'hEB2: dout <= 8'b00000000; // 3762 :   0 - 0x0
      13'hEB3: dout <= 8'b00000000; // 3763 :   0 - 0x0
      13'hEB4: dout <= 8'b00000000; // 3764 :   0 - 0x0
      13'hEB5: dout <= 8'b00000000; // 3765 :   0 - 0x0
      13'hEB6: dout <= 8'b00000000; // 3766 :   0 - 0x0
      13'hEB7: dout <= 8'b00000000; // 3767 :   0 - 0x0
      13'hEB8: dout <= 8'b00000000; // 3768 :   0 - 0x0
      13'hEB9: dout <= 8'b00000000; // 3769 :   0 - 0x0
      13'hEBA: dout <= 8'b00000000; // 3770 :   0 - 0x0
      13'hEBB: dout <= 8'b00000000; // 3771 :   0 - 0x0
      13'hEBC: dout <= 8'b00000000; // 3772 :   0 - 0x0
      13'hEBD: dout <= 8'b00000000; // 3773 :   0 - 0x0
      13'hEBE: dout <= 8'b00000000; // 3774 :   0 - 0x0
      13'hEBF: dout <= 8'b00000000; // 3775 :   0 - 0x0
      13'hEC0: dout <= 8'b00000000; // 3776 :   0 - 0x0 -- Sprite 0xec
      13'hEC1: dout <= 8'b00000000; // 3777 :   0 - 0x0
      13'hEC2: dout <= 8'b00000000; // 3778 :   0 - 0x0
      13'hEC3: dout <= 8'b00000000; // 3779 :   0 - 0x0
      13'hEC4: dout <= 8'b00000000; // 3780 :   0 - 0x0
      13'hEC5: dout <= 8'b00000000; // 3781 :   0 - 0x0
      13'hEC6: dout <= 8'b00000000; // 3782 :   0 - 0x0
      13'hEC7: dout <= 8'b00000000; // 3783 :   0 - 0x0
      13'hEC8: dout <= 8'b00000000; // 3784 :   0 - 0x0
      13'hEC9: dout <= 8'b00000000; // 3785 :   0 - 0x0
      13'hECA: dout <= 8'b00000000; // 3786 :   0 - 0x0
      13'hECB: dout <= 8'b00000000; // 3787 :   0 - 0x0
      13'hECC: dout <= 8'b00000000; // 3788 :   0 - 0x0
      13'hECD: dout <= 8'b00000000; // 3789 :   0 - 0x0
      13'hECE: dout <= 8'b00000000; // 3790 :   0 - 0x0
      13'hECF: dout <= 8'b00000000; // 3791 :   0 - 0x0
      13'hED0: dout <= 8'b00000000; // 3792 :   0 - 0x0 -- Sprite 0xed
      13'hED1: dout <= 8'b00000000; // 3793 :   0 - 0x0
      13'hED2: dout <= 8'b00000000; // 3794 :   0 - 0x0
      13'hED3: dout <= 8'b00000000; // 3795 :   0 - 0x0
      13'hED4: dout <= 8'b00000000; // 3796 :   0 - 0x0
      13'hED5: dout <= 8'b00000000; // 3797 :   0 - 0x0
      13'hED6: dout <= 8'b00000000; // 3798 :   0 - 0x0
      13'hED7: dout <= 8'b00000000; // 3799 :   0 - 0x0
      13'hED8: dout <= 8'b00000000; // 3800 :   0 - 0x0
      13'hED9: dout <= 8'b00000000; // 3801 :   0 - 0x0
      13'hEDA: dout <= 8'b00000000; // 3802 :   0 - 0x0
      13'hEDB: dout <= 8'b00000000; // 3803 :   0 - 0x0
      13'hEDC: dout <= 8'b00000000; // 3804 :   0 - 0x0
      13'hEDD: dout <= 8'b00000000; // 3805 :   0 - 0x0
      13'hEDE: dout <= 8'b00000000; // 3806 :   0 - 0x0
      13'hEDF: dout <= 8'b00000000; // 3807 :   0 - 0x0
      13'hEE0: dout <= 8'b00000000; // 3808 :   0 - 0x0 -- Sprite 0xee
      13'hEE1: dout <= 8'b00000000; // 3809 :   0 - 0x0
      13'hEE2: dout <= 8'b00000000; // 3810 :   0 - 0x0
      13'hEE3: dout <= 8'b00000000; // 3811 :   0 - 0x0
      13'hEE4: dout <= 8'b00000000; // 3812 :   0 - 0x0
      13'hEE5: dout <= 8'b00000000; // 3813 :   0 - 0x0
      13'hEE6: dout <= 8'b00000000; // 3814 :   0 - 0x0
      13'hEE7: dout <= 8'b00000000; // 3815 :   0 - 0x0
      13'hEE8: dout <= 8'b00000000; // 3816 :   0 - 0x0
      13'hEE9: dout <= 8'b00000000; // 3817 :   0 - 0x0
      13'hEEA: dout <= 8'b00000000; // 3818 :   0 - 0x0
      13'hEEB: dout <= 8'b00000000; // 3819 :   0 - 0x0
      13'hEEC: dout <= 8'b00000000; // 3820 :   0 - 0x0
      13'hEED: dout <= 8'b00000000; // 3821 :   0 - 0x0
      13'hEEE: dout <= 8'b00000000; // 3822 :   0 - 0x0
      13'hEEF: dout <= 8'b00000000; // 3823 :   0 - 0x0
      13'hEF0: dout <= 8'b00000000; // 3824 :   0 - 0x0 -- Sprite 0xef
      13'hEF1: dout <= 8'b00000000; // 3825 :   0 - 0x0
      13'hEF2: dout <= 8'b00000000; // 3826 :   0 - 0x0
      13'hEF3: dout <= 8'b00000000; // 3827 :   0 - 0x0
      13'hEF4: dout <= 8'b00000000; // 3828 :   0 - 0x0
      13'hEF5: dout <= 8'b00000000; // 3829 :   0 - 0x0
      13'hEF6: dout <= 8'b00000000; // 3830 :   0 - 0x0
      13'hEF7: dout <= 8'b00000000; // 3831 :   0 - 0x0
      13'hEF8: dout <= 8'b00000000; // 3832 :   0 - 0x0
      13'hEF9: dout <= 8'b00000000; // 3833 :   0 - 0x0
      13'hEFA: dout <= 8'b00000000; // 3834 :   0 - 0x0
      13'hEFB: dout <= 8'b00000000; // 3835 :   0 - 0x0
      13'hEFC: dout <= 8'b00000000; // 3836 :   0 - 0x0
      13'hEFD: dout <= 8'b00000000; // 3837 :   0 - 0x0
      13'hEFE: dout <= 8'b00000000; // 3838 :   0 - 0x0
      13'hEFF: dout <= 8'b00000000; // 3839 :   0 - 0x0
      13'hF00: dout <= 8'b00000000; // 3840 :   0 - 0x0 -- Sprite 0xf0
      13'hF01: dout <= 8'b00000000; // 3841 :   0 - 0x0
      13'hF02: dout <= 8'b00000000; // 3842 :   0 - 0x0
      13'hF03: dout <= 8'b00000000; // 3843 :   0 - 0x0
      13'hF04: dout <= 8'b00000000; // 3844 :   0 - 0x0
      13'hF05: dout <= 8'b00000000; // 3845 :   0 - 0x0
      13'hF06: dout <= 8'b00000000; // 3846 :   0 - 0x0
      13'hF07: dout <= 8'b00000000; // 3847 :   0 - 0x0
      13'hF08: dout <= 8'b00000000; // 3848 :   0 - 0x0
      13'hF09: dout <= 8'b00000000; // 3849 :   0 - 0x0
      13'hF0A: dout <= 8'b00000000; // 3850 :   0 - 0x0
      13'hF0B: dout <= 8'b00000000; // 3851 :   0 - 0x0
      13'hF0C: dout <= 8'b00000000; // 3852 :   0 - 0x0
      13'hF0D: dout <= 8'b00000000; // 3853 :   0 - 0x0
      13'hF0E: dout <= 8'b00000000; // 3854 :   0 - 0x0
      13'hF0F: dout <= 8'b00000000; // 3855 :   0 - 0x0
      13'hF10: dout <= 8'b00000000; // 3856 :   0 - 0x0 -- Sprite 0xf1
      13'hF11: dout <= 8'b00000000; // 3857 :   0 - 0x0
      13'hF12: dout <= 8'b00000000; // 3858 :   0 - 0x0
      13'hF13: dout <= 8'b00000000; // 3859 :   0 - 0x0
      13'hF14: dout <= 8'b00000000; // 3860 :   0 - 0x0
      13'hF15: dout <= 8'b00000000; // 3861 :   0 - 0x0
      13'hF16: dout <= 8'b00000000; // 3862 :   0 - 0x0
      13'hF17: dout <= 8'b00000000; // 3863 :   0 - 0x0
      13'hF18: dout <= 8'b00000000; // 3864 :   0 - 0x0
      13'hF19: dout <= 8'b00000000; // 3865 :   0 - 0x0
      13'hF1A: dout <= 8'b00000000; // 3866 :   0 - 0x0
      13'hF1B: dout <= 8'b00000000; // 3867 :   0 - 0x0
      13'hF1C: dout <= 8'b00000000; // 3868 :   0 - 0x0
      13'hF1D: dout <= 8'b00000000; // 3869 :   0 - 0x0
      13'hF1E: dout <= 8'b00000000; // 3870 :   0 - 0x0
      13'hF1F: dout <= 8'b00000000; // 3871 :   0 - 0x0
      13'hF20: dout <= 8'b00000000; // 3872 :   0 - 0x0 -- Sprite 0xf2
      13'hF21: dout <= 8'b00000000; // 3873 :   0 - 0x0
      13'hF22: dout <= 8'b00000000; // 3874 :   0 - 0x0
      13'hF23: dout <= 8'b00000000; // 3875 :   0 - 0x0
      13'hF24: dout <= 8'b00000000; // 3876 :   0 - 0x0
      13'hF25: dout <= 8'b00000000; // 3877 :   0 - 0x0
      13'hF26: dout <= 8'b00000000; // 3878 :   0 - 0x0
      13'hF27: dout <= 8'b00000000; // 3879 :   0 - 0x0
      13'hF28: dout <= 8'b00000000; // 3880 :   0 - 0x0
      13'hF29: dout <= 8'b00000000; // 3881 :   0 - 0x0
      13'hF2A: dout <= 8'b00000000; // 3882 :   0 - 0x0
      13'hF2B: dout <= 8'b00000000; // 3883 :   0 - 0x0
      13'hF2C: dout <= 8'b00000000; // 3884 :   0 - 0x0
      13'hF2D: dout <= 8'b00000000; // 3885 :   0 - 0x0
      13'hF2E: dout <= 8'b00000000; // 3886 :   0 - 0x0
      13'hF2F: dout <= 8'b00000000; // 3887 :   0 - 0x0
      13'hF30: dout <= 8'b00000000; // 3888 :   0 - 0x0 -- Sprite 0xf3
      13'hF31: dout <= 8'b00000000; // 3889 :   0 - 0x0
      13'hF32: dout <= 8'b00000000; // 3890 :   0 - 0x0
      13'hF33: dout <= 8'b00000000; // 3891 :   0 - 0x0
      13'hF34: dout <= 8'b00000000; // 3892 :   0 - 0x0
      13'hF35: dout <= 8'b00000000; // 3893 :   0 - 0x0
      13'hF36: dout <= 8'b00000000; // 3894 :   0 - 0x0
      13'hF37: dout <= 8'b00000000; // 3895 :   0 - 0x0
      13'hF38: dout <= 8'b00000000; // 3896 :   0 - 0x0
      13'hF39: dout <= 8'b00000000; // 3897 :   0 - 0x0
      13'hF3A: dout <= 8'b00000000; // 3898 :   0 - 0x0
      13'hF3B: dout <= 8'b00000000; // 3899 :   0 - 0x0
      13'hF3C: dout <= 8'b00000000; // 3900 :   0 - 0x0
      13'hF3D: dout <= 8'b00000000; // 3901 :   0 - 0x0
      13'hF3E: dout <= 8'b00000000; // 3902 :   0 - 0x0
      13'hF3F: dout <= 8'b00000000; // 3903 :   0 - 0x0
      13'hF40: dout <= 8'b00000000; // 3904 :   0 - 0x0 -- Sprite 0xf4
      13'hF41: dout <= 8'b00000000; // 3905 :   0 - 0x0
      13'hF42: dout <= 8'b00000000; // 3906 :   0 - 0x0
      13'hF43: dout <= 8'b00000000; // 3907 :   0 - 0x0
      13'hF44: dout <= 8'b00000000; // 3908 :   0 - 0x0
      13'hF45: dout <= 8'b00000000; // 3909 :   0 - 0x0
      13'hF46: dout <= 8'b00000000; // 3910 :   0 - 0x0
      13'hF47: dout <= 8'b00000000; // 3911 :   0 - 0x0
      13'hF48: dout <= 8'b00000000; // 3912 :   0 - 0x0
      13'hF49: dout <= 8'b00000000; // 3913 :   0 - 0x0
      13'hF4A: dout <= 8'b00000000; // 3914 :   0 - 0x0
      13'hF4B: dout <= 8'b00000000; // 3915 :   0 - 0x0
      13'hF4C: dout <= 8'b00000000; // 3916 :   0 - 0x0
      13'hF4D: dout <= 8'b00000000; // 3917 :   0 - 0x0
      13'hF4E: dout <= 8'b00000000; // 3918 :   0 - 0x0
      13'hF4F: dout <= 8'b00000000; // 3919 :   0 - 0x0
      13'hF50: dout <= 8'b00000000; // 3920 :   0 - 0x0 -- Sprite 0xf5
      13'hF51: dout <= 8'b00000000; // 3921 :   0 - 0x0
      13'hF52: dout <= 8'b00000000; // 3922 :   0 - 0x0
      13'hF53: dout <= 8'b00000000; // 3923 :   0 - 0x0
      13'hF54: dout <= 8'b00000000; // 3924 :   0 - 0x0
      13'hF55: dout <= 8'b00000000; // 3925 :   0 - 0x0
      13'hF56: dout <= 8'b00000000; // 3926 :   0 - 0x0
      13'hF57: dout <= 8'b00000000; // 3927 :   0 - 0x0
      13'hF58: dout <= 8'b00000000; // 3928 :   0 - 0x0
      13'hF59: dout <= 8'b00000000; // 3929 :   0 - 0x0
      13'hF5A: dout <= 8'b00000000; // 3930 :   0 - 0x0
      13'hF5B: dout <= 8'b00000000; // 3931 :   0 - 0x0
      13'hF5C: dout <= 8'b00000000; // 3932 :   0 - 0x0
      13'hF5D: dout <= 8'b00000000; // 3933 :   0 - 0x0
      13'hF5E: dout <= 8'b00000000; // 3934 :   0 - 0x0
      13'hF5F: dout <= 8'b00000000; // 3935 :   0 - 0x0
      13'hF60: dout <= 8'b00000000; // 3936 :   0 - 0x0 -- Sprite 0xf6
      13'hF61: dout <= 8'b00000000; // 3937 :   0 - 0x0
      13'hF62: dout <= 8'b00000000; // 3938 :   0 - 0x0
      13'hF63: dout <= 8'b00000000; // 3939 :   0 - 0x0
      13'hF64: dout <= 8'b00000000; // 3940 :   0 - 0x0
      13'hF65: dout <= 8'b00000000; // 3941 :   0 - 0x0
      13'hF66: dout <= 8'b00000000; // 3942 :   0 - 0x0
      13'hF67: dout <= 8'b00000000; // 3943 :   0 - 0x0
      13'hF68: dout <= 8'b00000000; // 3944 :   0 - 0x0
      13'hF69: dout <= 8'b00000000; // 3945 :   0 - 0x0
      13'hF6A: dout <= 8'b00000000; // 3946 :   0 - 0x0
      13'hF6B: dout <= 8'b00000000; // 3947 :   0 - 0x0
      13'hF6C: dout <= 8'b00000000; // 3948 :   0 - 0x0
      13'hF6D: dout <= 8'b00000000; // 3949 :   0 - 0x0
      13'hF6E: dout <= 8'b00000000; // 3950 :   0 - 0x0
      13'hF6F: dout <= 8'b00000000; // 3951 :   0 - 0x0
      13'hF70: dout <= 8'b00000000; // 3952 :   0 - 0x0 -- Sprite 0xf7
      13'hF71: dout <= 8'b00000000; // 3953 :   0 - 0x0
      13'hF72: dout <= 8'b00000000; // 3954 :   0 - 0x0
      13'hF73: dout <= 8'b00000000; // 3955 :   0 - 0x0
      13'hF74: dout <= 8'b00000000; // 3956 :   0 - 0x0
      13'hF75: dout <= 8'b00000000; // 3957 :   0 - 0x0
      13'hF76: dout <= 8'b00000000; // 3958 :   0 - 0x0
      13'hF77: dout <= 8'b00000000; // 3959 :   0 - 0x0
      13'hF78: dout <= 8'b00000000; // 3960 :   0 - 0x0
      13'hF79: dout <= 8'b00000000; // 3961 :   0 - 0x0
      13'hF7A: dout <= 8'b00000000; // 3962 :   0 - 0x0
      13'hF7B: dout <= 8'b00000000; // 3963 :   0 - 0x0
      13'hF7C: dout <= 8'b00000000; // 3964 :   0 - 0x0
      13'hF7D: dout <= 8'b00000000; // 3965 :   0 - 0x0
      13'hF7E: dout <= 8'b00000000; // 3966 :   0 - 0x0
      13'hF7F: dout <= 8'b00000000; // 3967 :   0 - 0x0
      13'hF80: dout <= 8'b00000000; // 3968 :   0 - 0x0 -- Sprite 0xf8
      13'hF81: dout <= 8'b00000000; // 3969 :   0 - 0x0
      13'hF82: dout <= 8'b00000000; // 3970 :   0 - 0x0
      13'hF83: dout <= 8'b00000000; // 3971 :   0 - 0x0
      13'hF84: dout <= 8'b00000000; // 3972 :   0 - 0x0
      13'hF85: dout <= 8'b00000000; // 3973 :   0 - 0x0
      13'hF86: dout <= 8'b00000000; // 3974 :   0 - 0x0
      13'hF87: dout <= 8'b00000000; // 3975 :   0 - 0x0
      13'hF88: dout <= 8'b00000000; // 3976 :   0 - 0x0
      13'hF89: dout <= 8'b00000000; // 3977 :   0 - 0x0
      13'hF8A: dout <= 8'b00000000; // 3978 :   0 - 0x0
      13'hF8B: dout <= 8'b00000000; // 3979 :   0 - 0x0
      13'hF8C: dout <= 8'b00000000; // 3980 :   0 - 0x0
      13'hF8D: dout <= 8'b00000000; // 3981 :   0 - 0x0
      13'hF8E: dout <= 8'b00000000; // 3982 :   0 - 0x0
      13'hF8F: dout <= 8'b00000000; // 3983 :   0 - 0x0
      13'hF90: dout <= 8'b00000000; // 3984 :   0 - 0x0 -- Sprite 0xf9
      13'hF91: dout <= 8'b00000000; // 3985 :   0 - 0x0
      13'hF92: dout <= 8'b00000000; // 3986 :   0 - 0x0
      13'hF93: dout <= 8'b00000000; // 3987 :   0 - 0x0
      13'hF94: dout <= 8'b00000000; // 3988 :   0 - 0x0
      13'hF95: dout <= 8'b00000000; // 3989 :   0 - 0x0
      13'hF96: dout <= 8'b00000000; // 3990 :   0 - 0x0
      13'hF97: dout <= 8'b00000000; // 3991 :   0 - 0x0
      13'hF98: dout <= 8'b00000000; // 3992 :   0 - 0x0
      13'hF99: dout <= 8'b00000000; // 3993 :   0 - 0x0
      13'hF9A: dout <= 8'b00000000; // 3994 :   0 - 0x0
      13'hF9B: dout <= 8'b00000000; // 3995 :   0 - 0x0
      13'hF9C: dout <= 8'b00000000; // 3996 :   0 - 0x0
      13'hF9D: dout <= 8'b00000000; // 3997 :   0 - 0x0
      13'hF9E: dout <= 8'b00000000; // 3998 :   0 - 0x0
      13'hF9F: dout <= 8'b00000000; // 3999 :   0 - 0x0
      13'hFA0: dout <= 8'b00000000; // 4000 :   0 - 0x0 -- Sprite 0xfa
      13'hFA1: dout <= 8'b00000000; // 4001 :   0 - 0x0
      13'hFA2: dout <= 8'b00000000; // 4002 :   0 - 0x0
      13'hFA3: dout <= 8'b00000000; // 4003 :   0 - 0x0
      13'hFA4: dout <= 8'b00000000; // 4004 :   0 - 0x0
      13'hFA5: dout <= 8'b00000000; // 4005 :   0 - 0x0
      13'hFA6: dout <= 8'b00000000; // 4006 :   0 - 0x0
      13'hFA7: dout <= 8'b00000000; // 4007 :   0 - 0x0
      13'hFA8: dout <= 8'b00000000; // 4008 :   0 - 0x0
      13'hFA9: dout <= 8'b00000000; // 4009 :   0 - 0x0
      13'hFAA: dout <= 8'b00000000; // 4010 :   0 - 0x0
      13'hFAB: dout <= 8'b00000000; // 4011 :   0 - 0x0
      13'hFAC: dout <= 8'b00000000; // 4012 :   0 - 0x0
      13'hFAD: dout <= 8'b00000000; // 4013 :   0 - 0x0
      13'hFAE: dout <= 8'b00000000; // 4014 :   0 - 0x0
      13'hFAF: dout <= 8'b00000000; // 4015 :   0 - 0x0
      13'hFB0: dout <= 8'b00000000; // 4016 :   0 - 0x0 -- Sprite 0xfb
      13'hFB1: dout <= 8'b00000000; // 4017 :   0 - 0x0
      13'hFB2: dout <= 8'b00000000; // 4018 :   0 - 0x0
      13'hFB3: dout <= 8'b00000000; // 4019 :   0 - 0x0
      13'hFB4: dout <= 8'b00000000; // 4020 :   0 - 0x0
      13'hFB5: dout <= 8'b00000000; // 4021 :   0 - 0x0
      13'hFB6: dout <= 8'b00000000; // 4022 :   0 - 0x0
      13'hFB7: dout <= 8'b00000000; // 4023 :   0 - 0x0
      13'hFB8: dout <= 8'b00000000; // 4024 :   0 - 0x0
      13'hFB9: dout <= 8'b00000000; // 4025 :   0 - 0x0
      13'hFBA: dout <= 8'b00000000; // 4026 :   0 - 0x0
      13'hFBB: dout <= 8'b00000000; // 4027 :   0 - 0x0
      13'hFBC: dout <= 8'b00000000; // 4028 :   0 - 0x0
      13'hFBD: dout <= 8'b00000000; // 4029 :   0 - 0x0
      13'hFBE: dout <= 8'b00000000; // 4030 :   0 - 0x0
      13'hFBF: dout <= 8'b00000000; // 4031 :   0 - 0x0
      13'hFC0: dout <= 8'b00000000; // 4032 :   0 - 0x0 -- Sprite 0xfc
      13'hFC1: dout <= 8'b00000000; // 4033 :   0 - 0x0
      13'hFC2: dout <= 8'b10001110; // 4034 : 142 - 0x8e
      13'hFC3: dout <= 8'b10001010; // 4035 : 138 - 0x8a
      13'hFC4: dout <= 8'b10001010; // 4036 : 138 - 0x8a
      13'hFC5: dout <= 8'b10001010; // 4037 : 138 - 0x8a
      13'hFC6: dout <= 8'b10001010; // 4038 : 138 - 0x8a
      13'hFC7: dout <= 8'b11101110; // 4039 : 238 - 0xee
      13'hFC8: dout <= 8'b00000000; // 4040 :   0 - 0x0
      13'hFC9: dout <= 8'b00000000; // 4041 :   0 - 0x0
      13'hFCA: dout <= 8'b00000000; // 4042 :   0 - 0x0
      13'hFCB: dout <= 8'b00000000; // 4043 :   0 - 0x0
      13'hFCC: dout <= 8'b00000000; // 4044 :   0 - 0x0
      13'hFCD: dout <= 8'b00000000; // 4045 :   0 - 0x0
      13'hFCE: dout <= 8'b00000000; // 4046 :   0 - 0x0
      13'hFCF: dout <= 8'b00000000; // 4047 :   0 - 0x0
      13'hFD0: dout <= 8'b00000000; // 4048 :   0 - 0x0 -- Sprite 0xfd
      13'hFD1: dout <= 8'b00000000; // 4049 :   0 - 0x0
      13'hFD2: dout <= 8'b01001100; // 4050 :  76 - 0x4c
      13'hFD3: dout <= 8'b10101010; // 4051 : 170 - 0xaa
      13'hFD4: dout <= 8'b10101010; // 4052 : 170 - 0xaa
      13'hFD5: dout <= 8'b11101010; // 4053 : 234 - 0xea
      13'hFD6: dout <= 8'b10101010; // 4054 : 170 - 0xaa
      13'hFD7: dout <= 8'b10101100; // 4055 : 172 - 0xac
      13'hFD8: dout <= 8'b00000000; // 4056 :   0 - 0x0
      13'hFD9: dout <= 8'b00000000; // 4057 :   0 - 0x0
      13'hFDA: dout <= 8'b00000000; // 4058 :   0 - 0x0
      13'hFDB: dout <= 8'b00000000; // 4059 :   0 - 0x0
      13'hFDC: dout <= 8'b00000000; // 4060 :   0 - 0x0
      13'hFDD: dout <= 8'b00000000; // 4061 :   0 - 0x0
      13'hFDE: dout <= 8'b00000000; // 4062 :   0 - 0x0
      13'hFDF: dout <= 8'b00000000; // 4063 :   0 - 0x0
      13'hFE0: dout <= 8'b00000000; // 4064 :   0 - 0x0 -- Sprite 0xfe
      13'hFE1: dout <= 8'b00000000; // 4065 :   0 - 0x0
      13'hFE2: dout <= 8'b11101100; // 4066 : 236 - 0xec
      13'hFE3: dout <= 8'b01001010; // 4067 :  74 - 0x4a
      13'hFE4: dout <= 8'b01001010; // 4068 :  74 - 0x4a
      13'hFE5: dout <= 8'b01001010; // 4069 :  74 - 0x4a
      13'hFE6: dout <= 8'b01001010; // 4070 :  74 - 0x4a
      13'hFE7: dout <= 8'b11101010; // 4071 : 234 - 0xea
      13'hFE8: dout <= 8'b00000000; // 4072 :   0 - 0x0
      13'hFE9: dout <= 8'b00000000; // 4073 :   0 - 0x0
      13'hFEA: dout <= 8'b00000000; // 4074 :   0 - 0x0
      13'hFEB: dout <= 8'b00000000; // 4075 :   0 - 0x0
      13'hFEC: dout <= 8'b00000000; // 4076 :   0 - 0x0
      13'hFED: dout <= 8'b00000000; // 4077 :   0 - 0x0
      13'hFEE: dout <= 8'b00000000; // 4078 :   0 - 0x0
      13'hFEF: dout <= 8'b00000000; // 4079 :   0 - 0x0
      13'hFF0: dout <= 8'b00000000; // 4080 :   0 - 0x0 -- Sprite 0xff
      13'hFF1: dout <= 8'b00000000; // 4081 :   0 - 0x0
      13'hFF2: dout <= 8'b01100000; // 4082 :  96 - 0x60
      13'hFF3: dout <= 8'b10001000; // 4083 : 136 - 0x88
      13'hFF4: dout <= 8'b10100000; // 4084 : 160 - 0xa0
      13'hFF5: dout <= 8'b10100000; // 4085 : 160 - 0xa0
      13'hFF6: dout <= 8'b10101000; // 4086 : 168 - 0xa8
      13'hFF7: dout <= 8'b01000000; // 4087 :  64 - 0x40
      13'hFF8: dout <= 8'b00000000; // 4088 :   0 - 0x0
      13'hFF9: dout <= 8'b00000000; // 4089 :   0 - 0x0
      13'hFFA: dout <= 8'b00000000; // 4090 :   0 - 0x0
      13'hFFB: dout <= 8'b00000000; // 4091 :   0 - 0x0
      13'hFFC: dout <= 8'b00000000; // 4092 :   0 - 0x0
      13'hFFD: dout <= 8'b00000000; // 4093 :   0 - 0x0
      13'hFFE: dout <= 8'b00000000; // 4094 :   0 - 0x0
      13'hFFF: dout <= 8'b00000000; // 4095 :   0 - 0x0
          // Pattern Table 1---------
      13'h1000: dout <= 8'b00000000; // 4096 :   0 - 0x0 -- Background 0x0
      13'h1001: dout <= 8'b00001111; // 4097 :  15 - 0xf
      13'h1002: dout <= 8'b00000100; // 4098 :   4 - 0x4
      13'h1003: dout <= 8'b00000011; // 4099 :   3 - 0x3
      13'h1004: dout <= 8'b00000011; // 4100 :   3 - 0x3
      13'h1005: dout <= 8'b00000011; // 4101 :   3 - 0x3
      13'h1006: dout <= 8'b00000100; // 4102 :   4 - 0x4
      13'h1007: dout <= 8'b00111010; // 4103 :  58 - 0x3a
      13'h1008: dout <= 8'b00000000; // 4104 :   0 - 0x0
      13'h1009: dout <= 8'b00000000; // 4105 :   0 - 0x0
      13'h100A: dout <= 8'b00000011; // 4106 :   3 - 0x3
      13'h100B: dout <= 8'b00000001; // 4107 :   1 - 0x1
      13'h100C: dout <= 8'b00000001; // 4108 :   1 - 0x1
      13'h100D: dout <= 8'b00000000; // 4109 :   0 - 0x0
      13'h100E: dout <= 8'b00000011; // 4110 :   3 - 0x3
      13'h100F: dout <= 8'b00000001; // 4111 :   1 - 0x1
      13'h1010: dout <= 8'b00000000; // 4112 :   0 - 0x0 -- Background 0x1
      13'h1011: dout <= 8'b00111000; // 4113 :  56 - 0x38
      13'h1012: dout <= 8'b11000110; // 4114 : 198 - 0xc6
      13'h1013: dout <= 8'b11001011; // 4115 : 203 - 0xcb
      13'h1014: dout <= 8'b11011100; // 4116 : 220 - 0xdc
      13'h1015: dout <= 8'b00111010; // 4117 :  58 - 0x3a
      13'h1016: dout <= 8'b10011010; // 4118 : 154 - 0x9a
      13'h1017: dout <= 8'b10000001; // 4119 : 129 - 0x81
      13'h1018: dout <= 8'b00000000; // 4120 :   0 - 0x0
      13'h1019: dout <= 8'b00000000; // 4121 :   0 - 0x0
      13'h101A: dout <= 8'b00111000; // 4122 :  56 - 0x38
      13'h101B: dout <= 8'b10110100; // 4123 : 180 - 0xb4
      13'h101C: dout <= 8'b10101000; // 4124 : 168 - 0xa8
      13'h101D: dout <= 8'b11010100; // 4125 : 212 - 0xd4
      13'h101E: dout <= 8'b01110100; // 4126 : 116 - 0x74
      13'h101F: dout <= 8'b01111110; // 4127 : 126 - 0x7e
      13'h1020: dout <= 8'b01000101; // 4128 :  69 - 0x45 -- Background 0x2
      13'h1021: dout <= 8'b10000111; // 4129 : 135 - 0x87
      13'h1022: dout <= 8'b10000011; // 4130 : 131 - 0x83
      13'h1023: dout <= 8'b10000001; // 4131 : 129 - 0x81
      13'h1024: dout <= 8'b10000001; // 4132 : 129 - 0x81
      13'h1025: dout <= 8'b10000001; // 4133 : 129 - 0x81
      13'h1026: dout <= 8'b01000001; // 4134 :  65 - 0x41
      13'h1027: dout <= 8'b00100001; // 4135 :  33 - 0x21
      13'h1028: dout <= 8'b00111000; // 4136 :  56 - 0x38
      13'h1029: dout <= 8'b01111000; // 4137 : 120 - 0x78
      13'h102A: dout <= 8'b01111100; // 4138 : 124 - 0x7c
      13'h102B: dout <= 8'b01111110; // 4139 : 126 - 0x7e
      13'h102C: dout <= 8'b01111110; // 4140 : 126 - 0x7e
      13'h102D: dout <= 8'b01111110; // 4141 : 126 - 0x7e
      13'h102E: dout <= 8'b00111110; // 4142 :  62 - 0x3e
      13'h102F: dout <= 8'b00011110; // 4143 :  30 - 0x1e
      13'h1030: dout <= 8'b01111111; // 4144 : 127 - 0x7f -- Background 0x3
      13'h1031: dout <= 8'b01111110; // 4145 : 126 - 0x7e
      13'h1032: dout <= 8'b11111100; // 4146 : 252 - 0xfc
      13'h1033: dout <= 8'b00111000; // 4147 :  56 - 0x38
      13'h1034: dout <= 8'b00011000; // 4148 :  24 - 0x18
      13'h1035: dout <= 8'b10001100; // 4149 : 140 - 0x8c
      13'h1036: dout <= 8'b11000100; // 4150 : 196 - 0xc4
      13'h1037: dout <= 8'b11111100; // 4151 : 252 - 0xfc
      13'h1038: dout <= 8'b11110110; // 4152 : 246 - 0xf6
      13'h1039: dout <= 8'b11110000; // 4153 : 240 - 0xf0
      13'h103A: dout <= 8'b00111000; // 4154 :  56 - 0x38
      13'h103B: dout <= 8'b11010000; // 4155 : 208 - 0xd0
      13'h103C: dout <= 8'b11100000; // 4156 : 224 - 0xe0
      13'h103D: dout <= 8'b01110000; // 4157 : 112 - 0x70
      13'h103E: dout <= 8'b10111000; // 4158 : 184 - 0xb8
      13'h103F: dout <= 8'b01000000; // 4159 :  64 - 0x40
      13'h1040: dout <= 8'b00100011; // 4160 :  35 - 0x23 -- Background 0x4
      13'h1041: dout <= 8'b00100011; // 4161 :  35 - 0x23
      13'h1042: dout <= 8'b00100001; // 4162 :  33 - 0x21
      13'h1043: dout <= 8'b00100000; // 4163 :  32 - 0x20
      13'h1044: dout <= 8'b00010011; // 4164 :  19 - 0x13
      13'h1045: dout <= 8'b00001100; // 4165 :  12 - 0xc
      13'h1046: dout <= 8'b00000000; // 4166 :   0 - 0x0
      13'h1047: dout <= 8'b00000000; // 4167 :   0 - 0x0
      13'h1048: dout <= 8'b00011100; // 4168 :  28 - 0x1c
      13'h1049: dout <= 8'b00011100; // 4169 :  28 - 0x1c
      13'h104A: dout <= 8'b00011110; // 4170 :  30 - 0x1e
      13'h104B: dout <= 8'b00011111; // 4171 :  31 - 0x1f
      13'h104C: dout <= 8'b00001100; // 4172 :  12 - 0xc
      13'h104D: dout <= 8'b00000000; // 4173 :   0 - 0x0
      13'h104E: dout <= 8'b00000000; // 4174 :   0 - 0x0
      13'h104F: dout <= 8'b00000000; // 4175 :   0 - 0x0
      13'h1050: dout <= 8'b11111100; // 4176 : 252 - 0xfc -- Background 0x5
      13'h1051: dout <= 8'b11111100; // 4177 : 252 - 0xfc
      13'h1052: dout <= 8'b11111100; // 4178 : 252 - 0xfc
      13'h1053: dout <= 8'b11111100; // 4179 : 252 - 0xfc
      13'h1054: dout <= 8'b10010000; // 4180 : 144 - 0x90
      13'h1055: dout <= 8'b10010000; // 4181 : 144 - 0x90
      13'h1056: dout <= 8'b10001000; // 4182 : 136 - 0x88
      13'h1057: dout <= 8'b11111000; // 4183 : 248 - 0xf8
      13'h1058: dout <= 8'b10101000; // 4184 : 168 - 0xa8
      13'h1059: dout <= 8'b01010000; // 4185 :  80 - 0x50
      13'h105A: dout <= 8'b10101000; // 4186 : 168 - 0xa8
      13'h105B: dout <= 8'b00000000; // 4187 :   0 - 0x0
      13'h105C: dout <= 8'b01100000; // 4188 :  96 - 0x60
      13'h105D: dout <= 8'b01100000; // 4189 :  96 - 0x60
      13'h105E: dout <= 8'b01110000; // 4190 : 112 - 0x70
      13'h105F: dout <= 8'b00000000; // 4191 :   0 - 0x0
      13'h1060: dout <= 8'b00100011; // 4192 :  35 - 0x23 -- Background 0x6
      13'h1061: dout <= 8'b00100011; // 4193 :  35 - 0x23
      13'h1062: dout <= 8'b00100001; // 4194 :  33 - 0x21
      13'h1063: dout <= 8'b00100000; // 4195 :  32 - 0x20
      13'h1064: dout <= 8'b00010011; // 4196 :  19 - 0x13
      13'h1065: dout <= 8'b00001101; // 4197 :  13 - 0xd
      13'h1066: dout <= 8'b00000010; // 4198 :   2 - 0x2
      13'h1067: dout <= 8'b00000001; // 4199 :   1 - 0x1
      13'h1068: dout <= 8'b00011100; // 4200 :  28 - 0x1c
      13'h1069: dout <= 8'b00011100; // 4201 :  28 - 0x1c
      13'h106A: dout <= 8'b00011110; // 4202 :  30 - 0x1e
      13'h106B: dout <= 8'b00011111; // 4203 :  31 - 0x1f
      13'h106C: dout <= 8'b00001100; // 4204 :  12 - 0xc
      13'h106D: dout <= 8'b00000000; // 4205 :   0 - 0x0
      13'h106E: dout <= 8'b00000001; // 4206 :   1 - 0x1
      13'h106F: dout <= 8'b00000000; // 4207 :   0 - 0x0
      13'h1070: dout <= 8'b11111100; // 4208 : 252 - 0xfc -- Background 0x7
      13'h1071: dout <= 8'b11111100; // 4209 : 252 - 0xfc
      13'h1072: dout <= 8'b11111100; // 4210 : 252 - 0xfc
      13'h1073: dout <= 8'b11111100; // 4211 : 252 - 0xfc
      13'h1074: dout <= 8'b10100100; // 4212 : 164 - 0xa4
      13'h1075: dout <= 8'b00100100; // 4213 :  36 - 0x24
      13'h1076: dout <= 8'b01010010; // 4214 :  82 - 0x52
      13'h1077: dout <= 8'b11101110; // 4215 : 238 - 0xee
      13'h1078: dout <= 8'b10101000; // 4216 : 168 - 0xa8
      13'h1079: dout <= 8'b01010000; // 4217 :  80 - 0x50
      13'h107A: dout <= 8'b10101000; // 4218 : 168 - 0xa8
      13'h107B: dout <= 8'b00000000; // 4219 :   0 - 0x0
      13'h107C: dout <= 8'b01011000; // 4220 :  88 - 0x58
      13'h107D: dout <= 8'b11011000; // 4221 : 216 - 0xd8
      13'h107E: dout <= 8'b10001100; // 4222 : 140 - 0x8c
      13'h107F: dout <= 8'b00000000; // 4223 :   0 - 0x0
      13'h1080: dout <= 8'b00100011; // 4224 :  35 - 0x23 -- Background 0x8
      13'h1081: dout <= 8'b00100011; // 4225 :  35 - 0x23
      13'h1082: dout <= 8'b00100001; // 4226 :  33 - 0x21
      13'h1083: dout <= 8'b00100000; // 4227 :  32 - 0x20
      13'h1084: dout <= 8'b00010011; // 4228 :  19 - 0x13
      13'h1085: dout <= 8'b00001101; // 4229 :  13 - 0xd
      13'h1086: dout <= 8'b00000001; // 4230 :   1 - 0x1
      13'h1087: dout <= 8'b00000001; // 4231 :   1 - 0x1
      13'h1088: dout <= 8'b00011100; // 4232 :  28 - 0x1c
      13'h1089: dout <= 8'b00011100; // 4233 :  28 - 0x1c
      13'h108A: dout <= 8'b00011110; // 4234 :  30 - 0x1e
      13'h108B: dout <= 8'b00011111; // 4235 :  31 - 0x1f
      13'h108C: dout <= 8'b00001100; // 4236 :  12 - 0xc
      13'h108D: dout <= 8'b00000000; // 4237 :   0 - 0x0
      13'h108E: dout <= 8'b00000000; // 4238 :   0 - 0x0
      13'h108F: dout <= 8'b00000000; // 4239 :   0 - 0x0
      13'h1090: dout <= 8'b11111110; // 4240 : 254 - 0xfe -- Background 0x9
      13'h1091: dout <= 8'b11111110; // 4241 : 254 - 0xfe
      13'h1092: dout <= 8'b11111110; // 4242 : 254 - 0xfe
      13'h1093: dout <= 8'b11111111; // 4243 : 255 - 0xff
      13'h1094: dout <= 8'b10010001; // 4244 : 145 - 0x91
      13'h1095: dout <= 8'b00101111; // 4245 :  47 - 0x2f
      13'h1096: dout <= 8'b01000000; // 4246 :  64 - 0x40
      13'h1097: dout <= 8'b11100000; // 4247 : 224 - 0xe0
      13'h1098: dout <= 8'b10101000; // 4248 : 168 - 0xa8
      13'h1099: dout <= 8'b01010100; // 4249 :  84 - 0x54
      13'h109A: dout <= 8'b10101000; // 4250 : 168 - 0xa8
      13'h109B: dout <= 8'b00000000; // 4251 :   0 - 0x0
      13'h109C: dout <= 8'b01101110; // 4252 : 110 - 0x6e
      13'h109D: dout <= 8'b11000000; // 4253 : 192 - 0xc0
      13'h109E: dout <= 8'b10000000; // 4254 : 128 - 0x80
      13'h109F: dout <= 8'b00000000; // 4255 :   0 - 0x0
      13'h10A0: dout <= 8'b00100011; // 4256 :  35 - 0x23 -- Background 0xa
      13'h10A1: dout <= 8'b00100011; // 4257 :  35 - 0x23
      13'h10A2: dout <= 8'b00100001; // 4258 :  33 - 0x21
      13'h10A3: dout <= 8'b00100000; // 4259 :  32 - 0x20
      13'h10A4: dout <= 8'b00010011; // 4260 :  19 - 0x13
      13'h10A5: dout <= 8'b00001110; // 4261 :  14 - 0xe
      13'h10A6: dout <= 8'b00000001; // 4262 :   1 - 0x1
      13'h10A7: dout <= 8'b00000000; // 4263 :   0 - 0x0
      13'h10A8: dout <= 8'b00011100; // 4264 :  28 - 0x1c
      13'h10A9: dout <= 8'b00011100; // 4265 :  28 - 0x1c
      13'h10AA: dout <= 8'b00011110; // 4266 :  30 - 0x1e
      13'h10AB: dout <= 8'b00011111; // 4267 :  31 - 0x1f
      13'h10AC: dout <= 8'b00001100; // 4268 :  12 - 0xc
      13'h10AD: dout <= 8'b00000001; // 4269 :   1 - 0x1
      13'h10AE: dout <= 8'b00000000; // 4270 :   0 - 0x0
      13'h10AF: dout <= 8'b00000000; // 4271 :   0 - 0x0
      13'h10B0: dout <= 8'b11111110; // 4272 : 254 - 0xfe -- Background 0xb
      13'h10B1: dout <= 8'b11111110; // 4273 : 254 - 0xfe
      13'h10B2: dout <= 8'b11111110; // 4274 : 254 - 0xfe
      13'h10B3: dout <= 8'b11111100; // 4275 : 252 - 0xfc
      13'h10B4: dout <= 8'b00100100; // 4276 :  36 - 0x24
      13'h10B5: dout <= 8'b00100010; // 4277 :  34 - 0x22
      13'h10B6: dout <= 8'b11010010; // 4278 : 210 - 0xd2
      13'h10B7: dout <= 8'b00001111; // 4279 :  15 - 0xf
      13'h10B8: dout <= 8'b10101000; // 4280 : 168 - 0xa8
      13'h10B9: dout <= 8'b01010100; // 4281 :  84 - 0x54
      13'h10BA: dout <= 8'b10101000; // 4282 : 168 - 0xa8
      13'h10BB: dout <= 8'b00000000; // 4283 :   0 - 0x0
      13'h10BC: dout <= 8'b11011000; // 4284 : 216 - 0xd8
      13'h10BD: dout <= 8'b11011100; // 4285 : 220 - 0xdc
      13'h10BE: dout <= 8'b00001100; // 4286 :  12 - 0xc
      13'h10BF: dout <= 8'b00000000; // 4287 :   0 - 0x0
      13'h10C0: dout <= 8'b01111111; // 4288 : 127 - 0x7f -- Background 0xc
      13'h10C1: dout <= 8'b01111110; // 4289 : 126 - 0x7e
      13'h10C2: dout <= 8'b11111100; // 4290 : 252 - 0xfc
      13'h10C3: dout <= 8'b00000010; // 4291 :   2 - 0x2
      13'h10C4: dout <= 8'b00000100; // 4292 :   4 - 0x4
      13'h10C5: dout <= 8'b11111100; // 4293 : 252 - 0xfc
      13'h10C6: dout <= 8'b11111100; // 4294 : 252 - 0xfc
      13'h10C7: dout <= 8'b11111110; // 4295 : 254 - 0xfe
      13'h10C8: dout <= 8'b11110110; // 4296 : 246 - 0xf6
      13'h10C9: dout <= 8'b11110000; // 4297 : 240 - 0xf0
      13'h10CA: dout <= 8'b00000000; // 4298 :   0 - 0x0
      13'h10CB: dout <= 8'b11111100; // 4299 : 252 - 0xfc
      13'h10CC: dout <= 8'b11111000; // 4300 : 248 - 0xf8
      13'h10CD: dout <= 8'b00000000; // 4301 :   0 - 0x0
      13'h10CE: dout <= 8'b10101000; // 4302 : 168 - 0xa8
      13'h10CF: dout <= 8'b01010100; // 4303 :  84 - 0x54
      13'h10D0: dout <= 8'b01000101; // 4304 :  69 - 0x45 -- Background 0xd
      13'h10D1: dout <= 8'b10000111; // 4305 : 135 - 0x87
      13'h10D2: dout <= 8'b10000011; // 4306 : 131 - 0x83
      13'h10D3: dout <= 8'b10000010; // 4307 : 130 - 0x82
      13'h10D4: dout <= 8'b10000010; // 4308 : 130 - 0x82
      13'h10D5: dout <= 8'b10000100; // 4309 : 132 - 0x84
      13'h10D6: dout <= 8'b01000100; // 4310 :  68 - 0x44
      13'h10D7: dout <= 8'b00100100; // 4311 :  36 - 0x24
      13'h10D8: dout <= 8'b00111000; // 4312 :  56 - 0x38
      13'h10D9: dout <= 8'b01111000; // 4313 : 120 - 0x78
      13'h10DA: dout <= 8'b01111100; // 4314 : 124 - 0x7c
      13'h10DB: dout <= 8'b01111101; // 4315 : 125 - 0x7d
      13'h10DC: dout <= 8'b01111101; // 4316 : 125 - 0x7d
      13'h10DD: dout <= 8'b01111011; // 4317 : 123 - 0x7b
      13'h10DE: dout <= 8'b00111011; // 4318 :  59 - 0x3b
      13'h10DF: dout <= 8'b00011011; // 4319 :  27 - 0x1b
      13'h10E0: dout <= 8'b01111111; // 4320 : 127 - 0x7f -- Background 0xe
      13'h10E1: dout <= 8'b01111110; // 4321 : 126 - 0x7e
      13'h10E2: dout <= 8'b11111100; // 4322 : 252 - 0xfc
      13'h10E3: dout <= 8'b11111000; // 4323 : 248 - 0xf8
      13'h10E4: dout <= 8'b01111000; // 4324 : 120 - 0x78
      13'h10E5: dout <= 8'b01111100; // 4325 : 124 - 0x7c
      13'h10E6: dout <= 8'b11111100; // 4326 : 252 - 0xfc
      13'h10E7: dout <= 8'b11111110; // 4327 : 254 - 0xfe
      13'h10E8: dout <= 8'b11110110; // 4328 : 246 - 0xf6
      13'h10E9: dout <= 8'b11110000; // 4329 : 240 - 0xf0
      13'h10EA: dout <= 8'b01111000; // 4330 : 120 - 0x78
      13'h10EB: dout <= 8'b01110000; // 4331 : 112 - 0x70
      13'h10EC: dout <= 8'b10100000; // 4332 : 160 - 0xa0
      13'h10ED: dout <= 8'b10010000; // 4333 : 144 - 0x90
      13'h10EE: dout <= 8'b00101000; // 4334 :  40 - 0x28
      13'h10EF: dout <= 8'b01010100; // 4335 :  84 - 0x54
      13'h10F0: dout <= 8'b00000000; // 4336 :   0 - 0x0 -- Background 0xf
      13'h10F1: dout <= 8'b00001111; // 4337 :  15 - 0xf
      13'h10F2: dout <= 8'b00000100; // 4338 :   4 - 0x4
      13'h10F3: dout <= 8'b00000011; // 4339 :   3 - 0x3
      13'h10F4: dout <= 8'b00000011; // 4340 :   3 - 0x3
      13'h10F5: dout <= 8'b00000011; // 4341 :   3 - 0x3
      13'h10F6: dout <= 8'b00000100; // 4342 :   4 - 0x4
      13'h10F7: dout <= 8'b00000010; // 4343 :   2 - 0x2
      13'h10F8: dout <= 8'b00000000; // 4344 :   0 - 0x0
      13'h10F9: dout <= 8'b00000000; // 4345 :   0 - 0x0
      13'h10FA: dout <= 8'b00000011; // 4346 :   3 - 0x3
      13'h10FB: dout <= 8'b00000001; // 4347 :   1 - 0x1
      13'h10FC: dout <= 8'b00000001; // 4348 :   1 - 0x1
      13'h10FD: dout <= 8'b00000000; // 4349 :   0 - 0x0
      13'h10FE: dout <= 8'b00000011; // 4350 :   3 - 0x3
      13'h10FF: dout <= 8'b00000001; // 4351 :   1 - 0x1
      13'h1100: dout <= 8'b00000111; // 4352 :   7 - 0x7 -- Background 0x10
      13'h1101: dout <= 8'b00001100; // 4353 :  12 - 0xc
      13'h1102: dout <= 8'b00010000; // 4354 :  16 - 0x10
      13'h1103: dout <= 8'b00010000; // 4355 :  16 - 0x10
      13'h1104: dout <= 8'b00010000; // 4356 :  16 - 0x10
      13'h1105: dout <= 8'b00100000; // 4357 :  32 - 0x20
      13'h1106: dout <= 8'b00100000; // 4358 :  32 - 0x20
      13'h1107: dout <= 8'b00100001; // 4359 :  33 - 0x21
      13'h1108: dout <= 8'b00000000; // 4360 :   0 - 0x0
      13'h1109: dout <= 8'b00000011; // 4361 :   3 - 0x3
      13'h110A: dout <= 8'b00001111; // 4362 :  15 - 0xf
      13'h110B: dout <= 8'b00001111; // 4363 :  15 - 0xf
      13'h110C: dout <= 8'b00001111; // 4364 :  15 - 0xf
      13'h110D: dout <= 8'b00011111; // 4365 :  31 - 0x1f
      13'h110E: dout <= 8'b00011111; // 4366 :  31 - 0x1f
      13'h110F: dout <= 8'b00011110; // 4367 :  30 - 0x1e
      13'h1110: dout <= 8'b11111111; // 4368 : 255 - 0xff -- Background 0x11
      13'h1111: dout <= 8'b01111110; // 4369 : 126 - 0x7e
      13'h1112: dout <= 8'b01111100; // 4370 : 124 - 0x7c
      13'h1113: dout <= 8'b01111000; // 4371 : 120 - 0x78
      13'h1114: dout <= 8'b01011000; // 4372 :  88 - 0x58
      13'h1115: dout <= 8'b10001100; // 4373 : 140 - 0x8c
      13'h1116: dout <= 8'b11000100; // 4374 : 196 - 0xc4
      13'h1117: dout <= 8'b11111100; // 4375 : 252 - 0xfc
      13'h1118: dout <= 8'b00110110; // 4376 :  54 - 0x36
      13'h1119: dout <= 8'b10110000; // 4377 : 176 - 0xb0
      13'h111A: dout <= 8'b10111000; // 4378 : 184 - 0xb8
      13'h111B: dout <= 8'b10010000; // 4379 : 144 - 0x90
      13'h111C: dout <= 8'b10100000; // 4380 : 160 - 0xa0
      13'h111D: dout <= 8'b01110000; // 4381 : 112 - 0x70
      13'h111E: dout <= 8'b00111000; // 4382 :  56 - 0x38
      13'h111F: dout <= 8'b01000000; // 4383 :  64 - 0x40
      13'h1120: dout <= 8'b00100011; // 4384 :  35 - 0x23 -- Background 0x12
      13'h1121: dout <= 8'b00100011; // 4385 :  35 - 0x23
      13'h1122: dout <= 8'b00100001; // 4386 :  33 - 0x21
      13'h1123: dout <= 8'b00100000; // 4387 :  32 - 0x20
      13'h1124: dout <= 8'b00010011; // 4388 :  19 - 0x13
      13'h1125: dout <= 8'b00001100; // 4389 :  12 - 0xc
      13'h1126: dout <= 8'b00000000; // 4390 :   0 - 0x0
      13'h1127: dout <= 8'b00000000; // 4391 :   0 - 0x0
      13'h1128: dout <= 8'b00011100; // 4392 :  28 - 0x1c
      13'h1129: dout <= 8'b00011100; // 4393 :  28 - 0x1c
      13'h112A: dout <= 8'b00011110; // 4394 :  30 - 0x1e
      13'h112B: dout <= 8'b00011111; // 4395 :  31 - 0x1f
      13'h112C: dout <= 8'b00001100; // 4396 :  12 - 0xc
      13'h112D: dout <= 8'b00000000; // 4397 :   0 - 0x0
      13'h112E: dout <= 8'b00000000; // 4398 :   0 - 0x0
      13'h112F: dout <= 8'b00000000; // 4399 :   0 - 0x0
      13'h1130: dout <= 8'b00000001; // 4400 :   1 - 0x1 -- Background 0x13
      13'h1131: dout <= 8'b00000001; // 4401 :   1 - 0x1
      13'h1132: dout <= 8'b00000011; // 4402 :   3 - 0x3
      13'h1133: dout <= 8'b00000100; // 4403 :   4 - 0x4
      13'h1134: dout <= 8'b00001000; // 4404 :   8 - 0x8
      13'h1135: dout <= 8'b00010000; // 4405 :  16 - 0x10
      13'h1136: dout <= 8'b00010000; // 4406 :  16 - 0x10
      13'h1137: dout <= 8'b00100000; // 4407 :  32 - 0x20
      13'h1138: dout <= 8'b00000000; // 4408 :   0 - 0x0
      13'h1139: dout <= 8'b00000000; // 4409 :   0 - 0x0
      13'h113A: dout <= 8'b00000000; // 4410 :   0 - 0x0
      13'h113B: dout <= 8'b00000011; // 4411 :   3 - 0x3
      13'h113C: dout <= 8'b00000111; // 4412 :   7 - 0x7
      13'h113D: dout <= 8'b00001111; // 4413 :  15 - 0xf
      13'h113E: dout <= 8'b00001111; // 4414 :  15 - 0xf
      13'h113F: dout <= 8'b00011111; // 4415 :  31 - 0x1f
      13'h1140: dout <= 8'b01111111; // 4416 : 127 - 0x7f -- Background 0x14
      13'h1141: dout <= 8'b11111110; // 4417 : 254 - 0xfe
      13'h1142: dout <= 8'b00000110; // 4418 :   6 - 0x6
      13'h1143: dout <= 8'b00000001; // 4419 :   1 - 0x1
      13'h1144: dout <= 8'b00000001; // 4420 :   1 - 0x1
      13'h1145: dout <= 8'b00000001; // 4421 :   1 - 0x1
      13'h1146: dout <= 8'b00000111; // 4422 :   7 - 0x7
      13'h1147: dout <= 8'b11111110; // 4423 : 254 - 0xfe
      13'h1148: dout <= 8'b11110110; // 4424 : 246 - 0xf6
      13'h1149: dout <= 8'b00000000; // 4425 :   0 - 0x0
      13'h114A: dout <= 8'b11111000; // 4426 : 248 - 0xf8
      13'h114B: dout <= 8'b11111110; // 4427 : 254 - 0xfe
      13'h114C: dout <= 8'b11111110; // 4428 : 254 - 0xfe
      13'h114D: dout <= 8'b11111110; // 4429 : 254 - 0xfe
      13'h114E: dout <= 8'b11111000; // 4430 : 248 - 0xf8
      13'h114F: dout <= 8'b00000000; // 4431 :   0 - 0x0
      13'h1150: dout <= 8'b00000101; // 4432 :   5 - 0x5 -- Background 0x15
      13'h1151: dout <= 8'b00000101; // 4433 :   5 - 0x5
      13'h1152: dout <= 8'b00000111; // 4434 :   7 - 0x7
      13'h1153: dout <= 8'b00000100; // 4435 :   4 - 0x4
      13'h1154: dout <= 8'b00000100; // 4436 :   4 - 0x4
      13'h1155: dout <= 8'b00001111; // 4437 :  15 - 0xf
      13'h1156: dout <= 8'b00110000; // 4438 :  48 - 0x30
      13'h1157: dout <= 8'b01000000; // 4439 :  64 - 0x40
      13'h1158: dout <= 8'b00000011; // 4440 :   3 - 0x3
      13'h1159: dout <= 8'b00000011; // 4441 :   3 - 0x3
      13'h115A: dout <= 8'b00000000; // 4442 :   0 - 0x0
      13'h115B: dout <= 8'b00000011; // 4443 :   3 - 0x3
      13'h115C: dout <= 8'b00000011; // 4444 :   3 - 0x3
      13'h115D: dout <= 8'b00000000; // 4445 :   0 - 0x0
      13'h115E: dout <= 8'b00001111; // 4446 :  15 - 0xf
      13'h115F: dout <= 8'b00111111; // 4447 :  63 - 0x3f
      13'h1160: dout <= 8'b11111100; // 4448 : 252 - 0xfc -- Background 0x16
      13'h1161: dout <= 8'b11111000; // 4449 : 248 - 0xf8
      13'h1162: dout <= 8'b11110000; // 4450 : 240 - 0xf0
      13'h1163: dout <= 8'b11100000; // 4451 : 224 - 0xe0
      13'h1164: dout <= 8'b01100000; // 4452 :  96 - 0x60
      13'h1165: dout <= 8'b11110000; // 4453 : 240 - 0xf0
      13'h1166: dout <= 8'b00011100; // 4454 :  28 - 0x1c
      13'h1167: dout <= 8'b00000010; // 4455 :   2 - 0x2
      13'h1168: dout <= 8'b11011000; // 4456 : 216 - 0xd8
      13'h1169: dout <= 8'b11000000; // 4457 : 192 - 0xc0
      13'h116A: dout <= 8'b11100000; // 4458 : 224 - 0xe0
      13'h116B: dout <= 8'b01000000; // 4459 :  64 - 0x40
      13'h116C: dout <= 8'b10000000; // 4460 : 128 - 0x80
      13'h116D: dout <= 8'b00000000; // 4461 :   0 - 0x0
      13'h116E: dout <= 8'b11100000; // 4462 : 224 - 0xe0
      13'h116F: dout <= 8'b11111100; // 4463 : 252 - 0xfc
      13'h1170: dout <= 8'b10000000; // 4464 : 128 - 0x80 -- Background 0x17
      13'h1171: dout <= 8'b10000000; // 4465 : 128 - 0x80
      13'h1172: dout <= 8'b10000000; // 4466 : 128 - 0x80
      13'h1173: dout <= 8'b10000011; // 4467 : 131 - 0x83
      13'h1174: dout <= 8'b01001111; // 4468 :  79 - 0x4f
      13'h1175: dout <= 8'b00110010; // 4469 :  50 - 0x32
      13'h1176: dout <= 8'b00000010; // 4470 :   2 - 0x2
      13'h1177: dout <= 8'b00000011; // 4471 :   3 - 0x3
      13'h1178: dout <= 8'b01111111; // 4472 : 127 - 0x7f
      13'h1179: dout <= 8'b01111111; // 4473 : 127 - 0x7f
      13'h117A: dout <= 8'b01111111; // 4474 : 127 - 0x7f
      13'h117B: dout <= 8'b01111100; // 4475 : 124 - 0x7c
      13'h117C: dout <= 8'b00110000; // 4476 :  48 - 0x30
      13'h117D: dout <= 8'b00000001; // 4477 :   1 - 0x1
      13'h117E: dout <= 8'b00000001; // 4478 :   1 - 0x1
      13'h117F: dout <= 8'b00000000; // 4479 :   0 - 0x0
      13'h1180: dout <= 8'b00000010; // 4480 :   2 - 0x2 -- Background 0x18
      13'h1181: dout <= 8'b00000001; // 4481 :   1 - 0x1
      13'h1182: dout <= 8'b00000010; // 4482 :   2 - 0x2
      13'h1183: dout <= 8'b11111100; // 4483 : 252 - 0xfc
      13'h1184: dout <= 8'b11000000; // 4484 : 192 - 0xc0
      13'h1185: dout <= 8'b01000000; // 4485 :  64 - 0x40
      13'h1186: dout <= 8'b00100000; // 4486 :  32 - 0x20
      13'h1187: dout <= 8'b11100000; // 4487 : 224 - 0xe0
      13'h1188: dout <= 8'b11111100; // 4488 : 252 - 0xfc
      13'h1189: dout <= 8'b11111110; // 4489 : 254 - 0xfe
      13'h118A: dout <= 8'b11111100; // 4490 : 252 - 0xfc
      13'h118B: dout <= 8'b00000000; // 4491 :   0 - 0x0
      13'h118C: dout <= 8'b00000000; // 4492 :   0 - 0x0
      13'h118D: dout <= 8'b10000000; // 4493 : 128 - 0x80
      13'h118E: dout <= 8'b11000000; // 4494 : 192 - 0xc0
      13'h118F: dout <= 8'b00000000; // 4495 :   0 - 0x0
      13'h1190: dout <= 8'b00001011; // 4496 :  11 - 0xb -- Background 0x19
      13'h1191: dout <= 8'b00001011; // 4497 :  11 - 0xb
      13'h1192: dout <= 8'b00001111; // 4498 :  15 - 0xf
      13'h1193: dout <= 8'b00001001; // 4499 :   9 - 0x9
      13'h1194: dout <= 8'b00001000; // 4500 :   8 - 0x8
      13'h1195: dout <= 8'b00001001; // 4501 :   9 - 0x9
      13'h1196: dout <= 8'b00001111; // 4502 :  15 - 0xf
      13'h1197: dout <= 8'b00110000; // 4503 :  48 - 0x30
      13'h1198: dout <= 8'b00000111; // 4504 :   7 - 0x7
      13'h1199: dout <= 8'b00000111; // 4505 :   7 - 0x7
      13'h119A: dout <= 8'b00000001; // 4506 :   1 - 0x1
      13'h119B: dout <= 8'b00000110; // 4507 :   6 - 0x6
      13'h119C: dout <= 8'b00000111; // 4508 :   7 - 0x7
      13'h119D: dout <= 8'b00000110; // 4509 :   6 - 0x6
      13'h119E: dout <= 8'b00000000; // 4510 :   0 - 0x0
      13'h119F: dout <= 8'b00001111; // 4511 :  15 - 0xf
      13'h11A0: dout <= 8'b11111000; // 4512 : 248 - 0xf8 -- Background 0x1a
      13'h11A1: dout <= 8'b11110000; // 4513 : 240 - 0xf0
      13'h11A2: dout <= 8'b11100000; // 4514 : 224 - 0xe0
      13'h11A3: dout <= 8'b11000000; // 4515 : 192 - 0xc0
      13'h11A4: dout <= 8'b11000000; // 4516 : 192 - 0xc0
      13'h11A5: dout <= 8'b11000000; // 4517 : 192 - 0xc0
      13'h11A6: dout <= 8'b11111000; // 4518 : 248 - 0xf8
      13'h11A7: dout <= 8'b00011111; // 4519 :  31 - 0x1f
      13'h11A8: dout <= 8'b10110000; // 4520 : 176 - 0xb0
      13'h11A9: dout <= 8'b10000000; // 4521 : 128 - 0x80
      13'h11AA: dout <= 8'b11000000; // 4522 : 192 - 0xc0
      13'h11AB: dout <= 8'b10000000; // 4523 : 128 - 0x80
      13'h11AC: dout <= 8'b00000000; // 4524 :   0 - 0x0
      13'h11AD: dout <= 8'b00000000; // 4525 :   0 - 0x0
      13'h11AE: dout <= 8'b00000000; // 4526 :   0 - 0x0
      13'h11AF: dout <= 8'b11100000; // 4527 : 224 - 0xe0
      13'h11B0: dout <= 8'b01000000; // 4528 :  64 - 0x40 -- Background 0x1b
      13'h11B1: dout <= 8'b01000000; // 4529 :  64 - 0x40
      13'h11B2: dout <= 8'b10000000; // 4530 : 128 - 0x80
      13'h11B3: dout <= 8'b10000000; // 4531 : 128 - 0x80
      13'h11B4: dout <= 8'b01000000; // 4532 :  64 - 0x40
      13'h11B5: dout <= 8'b00111111; // 4533 :  63 - 0x3f
      13'h11B6: dout <= 8'b00000100; // 4534 :   4 - 0x4
      13'h11B7: dout <= 8'b00000111; // 4535 :   7 - 0x7
      13'h11B8: dout <= 8'b00111111; // 4536 :  63 - 0x3f
      13'h11B9: dout <= 8'b00111111; // 4537 :  63 - 0x3f
      13'h11BA: dout <= 8'b01111111; // 4538 : 127 - 0x7f
      13'h11BB: dout <= 8'b01111111; // 4539 : 127 - 0x7f
      13'h11BC: dout <= 8'b00111111; // 4540 :  63 - 0x3f
      13'h11BD: dout <= 8'b00000000; // 4541 :   0 - 0x0
      13'h11BE: dout <= 8'b00000011; // 4542 :   3 - 0x3
      13'h11BF: dout <= 8'b00000000; // 4543 :   0 - 0x0
      13'h11C0: dout <= 8'b00000000; // 4544 :   0 - 0x0 -- Background 0x1c
      13'h11C1: dout <= 8'b00000000; // 4545 :   0 - 0x0
      13'h11C2: dout <= 8'b00000000; // 4546 :   0 - 0x0
      13'h11C3: dout <= 8'b00000000; // 4547 :   0 - 0x0
      13'h11C4: dout <= 8'b00000000; // 4548 :   0 - 0x0
      13'h11C5: dout <= 8'b11111111; // 4549 : 255 - 0xff
      13'h11C6: dout <= 8'b01000000; // 4550 :  64 - 0x40
      13'h11C7: dout <= 8'b11000000; // 4551 : 192 - 0xc0
      13'h11C8: dout <= 8'b11111111; // 4552 : 255 - 0xff
      13'h11C9: dout <= 8'b11111111; // 4553 : 255 - 0xff
      13'h11CA: dout <= 8'b11111111; // 4554 : 255 - 0xff
      13'h11CB: dout <= 8'b11111111; // 4555 : 255 - 0xff
      13'h11CC: dout <= 8'b11111111; // 4556 : 255 - 0xff
      13'h11CD: dout <= 8'b00000000; // 4557 :   0 - 0x0
      13'h11CE: dout <= 8'b10000000; // 4558 : 128 - 0x80
      13'h11CF: dout <= 8'b00000000; // 4559 :   0 - 0x0
      13'h11D0: dout <= 8'b11000000; // 4560 : 192 - 0xc0 -- Background 0x1d
      13'h11D1: dout <= 8'b00100000; // 4561 :  32 - 0x20
      13'h11D2: dout <= 8'b00100000; // 4562 :  32 - 0x20
      13'h11D3: dout <= 8'b00100000; // 4563 :  32 - 0x20
      13'h11D4: dout <= 8'b01000000; // 4564 :  64 - 0x40
      13'h11D5: dout <= 8'b10000000; // 4565 : 128 - 0x80
      13'h11D6: dout <= 8'b00000000; // 4566 :   0 - 0x0
      13'h11D7: dout <= 8'b00000000; // 4567 :   0 - 0x0
      13'h11D8: dout <= 8'b00000000; // 4568 :   0 - 0x0
      13'h11D9: dout <= 8'b11000000; // 4569 : 192 - 0xc0
      13'h11DA: dout <= 8'b11000000; // 4570 : 192 - 0xc0
      13'h11DB: dout <= 8'b11000000; // 4571 : 192 - 0xc0
      13'h11DC: dout <= 8'b10000000; // 4572 : 128 - 0x80
      13'h11DD: dout <= 8'b00000000; // 4573 :   0 - 0x0
      13'h11DE: dout <= 8'b00000000; // 4574 :   0 - 0x0
      13'h11DF: dout <= 8'b00000000; // 4575 :   0 - 0x0
      13'h11E0: dout <= 8'b01111111; // 4576 : 127 - 0x7f -- Background 0x1e
      13'h11E1: dout <= 8'b01100010; // 4577 :  98 - 0x62
      13'h11E2: dout <= 8'b11000100; // 4578 : 196 - 0xc4
      13'h11E3: dout <= 8'b00011000; // 4579 :  24 - 0x18
      13'h11E4: dout <= 8'b00111100; // 4580 :  60 - 0x3c
      13'h11E5: dout <= 8'b11111110; // 4581 : 254 - 0xfe
      13'h11E6: dout <= 8'b11111110; // 4582 : 254 - 0xfe
      13'h11E7: dout <= 8'b11111110; // 4583 : 254 - 0xfe
      13'h11E8: dout <= 8'b11100000; // 4584 : 224 - 0xe0
      13'h11E9: dout <= 8'b10011100; // 4585 : 156 - 0x9c
      13'h11EA: dout <= 8'b00111000; // 4586 :  56 - 0x38
      13'h11EB: dout <= 8'b11100000; // 4587 : 224 - 0xe0
      13'h11EC: dout <= 8'b11001000; // 4588 : 200 - 0xc8
      13'h11ED: dout <= 8'b00010100; // 4589 :  20 - 0x14
      13'h11EE: dout <= 8'b10101000; // 4590 : 168 - 0xa8
      13'h11EF: dout <= 8'b01010100; // 4591 :  84 - 0x54
      13'h11F0: dout <= 8'b00000000; // 4592 :   0 - 0x0 -- Background 0x1f
      13'h11F1: dout <= 8'b00111000; // 4593 :  56 - 0x38
      13'h11F2: dout <= 8'b11000110; // 4594 : 198 - 0xc6
      13'h11F3: dout <= 8'b11001011; // 4595 : 203 - 0xcb
      13'h11F4: dout <= 8'b11011100; // 4596 : 220 - 0xdc
      13'h11F5: dout <= 8'b00111010; // 4597 :  58 - 0x3a
      13'h11F6: dout <= 8'b10011010; // 4598 : 154 - 0x9a
      13'h11F7: dout <= 8'b11100001; // 4599 : 225 - 0xe1
      13'h11F8: dout <= 8'b00000000; // 4600 :   0 - 0x0
      13'h11F9: dout <= 8'b00000000; // 4601 :   0 - 0x0
      13'h11FA: dout <= 8'b00111000; // 4602 :  56 - 0x38
      13'h11FB: dout <= 8'b10110100; // 4603 : 180 - 0xb4
      13'h11FC: dout <= 8'b10101000; // 4604 : 168 - 0xa8
      13'h11FD: dout <= 8'b11010100; // 4605 : 212 - 0xd4
      13'h11FE: dout <= 8'b01110100; // 4606 : 116 - 0x74
      13'h11FF: dout <= 8'b00011110; // 4607 :  30 - 0x1e
      13'h1200: dout <= 8'b00000000; // 4608 :   0 - 0x0 -- Background 0x20
      13'h1201: dout <= 8'b00011100; // 4609 :  28 - 0x1c
      13'h1202: dout <= 8'b00010011; // 4610 :  19 - 0x13
      13'h1203: dout <= 8'b00001000; // 4611 :   8 - 0x8
      13'h1204: dout <= 8'b00010000; // 4612 :  16 - 0x10
      13'h1205: dout <= 8'b00001000; // 4613 :   8 - 0x8
      13'h1206: dout <= 8'b00010000; // 4614 :  16 - 0x10
      13'h1207: dout <= 8'b00010000; // 4615 :  16 - 0x10
      13'h1208: dout <= 8'b00000000; // 4616 :   0 - 0x0
      13'h1209: dout <= 8'b00000000; // 4617 :   0 - 0x0
      13'h120A: dout <= 8'b00001100; // 4618 :  12 - 0xc
      13'h120B: dout <= 8'b00000111; // 4619 :   7 - 0x7
      13'h120C: dout <= 8'b00001111; // 4620 :  15 - 0xf
      13'h120D: dout <= 8'b00000111; // 4621 :   7 - 0x7
      13'h120E: dout <= 8'b00001111; // 4622 :  15 - 0xf
      13'h120F: dout <= 8'b00001111; // 4623 :  15 - 0xf
      13'h1210: dout <= 8'b00000000; // 4624 :   0 - 0x0 -- Background 0x21
      13'h1211: dout <= 8'b00111000; // 4625 :  56 - 0x38
      13'h1212: dout <= 8'b11001000; // 4626 : 200 - 0xc8
      13'h1213: dout <= 8'b00010000; // 4627 :  16 - 0x10
      13'h1214: dout <= 8'b00001000; // 4628 :   8 - 0x8
      13'h1215: dout <= 8'b00010000; // 4629 :  16 - 0x10
      13'h1216: dout <= 8'b00001000; // 4630 :   8 - 0x8
      13'h1217: dout <= 8'b00001000; // 4631 :   8 - 0x8
      13'h1218: dout <= 8'b00000000; // 4632 :   0 - 0x0
      13'h1219: dout <= 8'b00000000; // 4633 :   0 - 0x0
      13'h121A: dout <= 8'b00110000; // 4634 :  48 - 0x30
      13'h121B: dout <= 8'b11100000; // 4635 : 224 - 0xe0
      13'h121C: dout <= 8'b11110000; // 4636 : 240 - 0xf0
      13'h121D: dout <= 8'b11100000; // 4637 : 224 - 0xe0
      13'h121E: dout <= 8'b11110000; // 4638 : 240 - 0xf0
      13'h121F: dout <= 8'b11110000; // 4639 : 240 - 0xf0
      13'h1220: dout <= 8'b00001000; // 4640 :   8 - 0x8 -- Background 0x22
      13'h1221: dout <= 8'b00011100; // 4641 :  28 - 0x1c
      13'h1222: dout <= 8'b00100111; // 4642 :  39 - 0x27
      13'h1223: dout <= 8'b00101111; // 4643 :  47 - 0x2f
      13'h1224: dout <= 8'b00011111; // 4644 :  31 - 0x1f
      13'h1225: dout <= 8'b00001111; // 4645 :  15 - 0xf
      13'h1226: dout <= 8'b00001111; // 4646 :  15 - 0xf
      13'h1227: dout <= 8'b00001111; // 4647 :  15 - 0xf
      13'h1228: dout <= 8'b00000111; // 4648 :   7 - 0x7
      13'h1229: dout <= 8'b00000011; // 4649 :   3 - 0x3
      13'h122A: dout <= 8'b00011000; // 4650 :  24 - 0x18
      13'h122B: dout <= 8'b00010101; // 4651 :  21 - 0x15
      13'h122C: dout <= 8'b00000010; // 4652 :   2 - 0x2
      13'h122D: dout <= 8'b00000101; // 4653 :   5 - 0x5
      13'h122E: dout <= 8'b00000010; // 4654 :   2 - 0x2
      13'h122F: dout <= 8'b00000100; // 4655 :   4 - 0x4
      13'h1230: dout <= 8'b00010000; // 4656 :  16 - 0x10 -- Background 0x23
      13'h1231: dout <= 8'b00111100; // 4657 :  60 - 0x3c
      13'h1232: dout <= 8'b11000010; // 4658 : 194 - 0xc2
      13'h1233: dout <= 8'b10000010; // 4659 : 130 - 0x82
      13'h1234: dout <= 8'b10000010; // 4660 : 130 - 0x82
      13'h1235: dout <= 8'b10000010; // 4661 : 130 - 0x82
      13'h1236: dout <= 8'b00010010; // 4662 :  18 - 0x12
      13'h1237: dout <= 8'b00011100; // 4663 :  28 - 0x1c
      13'h1238: dout <= 8'b11100000; // 4664 : 224 - 0xe0
      13'h1239: dout <= 8'b11000000; // 4665 : 192 - 0xc0
      13'h123A: dout <= 8'b00111100; // 4666 :  60 - 0x3c
      13'h123B: dout <= 8'b01111100; // 4667 : 124 - 0x7c
      13'h123C: dout <= 8'b01111100; // 4668 : 124 - 0x7c
      13'h123D: dout <= 8'b01111100; // 4669 : 124 - 0x7c
      13'h123E: dout <= 8'b11101100; // 4670 : 236 - 0xec
      13'h123F: dout <= 8'b11100000; // 4671 : 224 - 0xe0
      13'h1240: dout <= 8'b00001111; // 4672 :  15 - 0xf -- Background 0x24
      13'h1241: dout <= 8'b00001110; // 4673 :  14 - 0xe
      13'h1242: dout <= 8'b00010100; // 4674 :  20 - 0x14
      13'h1243: dout <= 8'b00010100; // 4675 :  20 - 0x14
      13'h1244: dout <= 8'b00010010; // 4676 :  18 - 0x12
      13'h1245: dout <= 8'b00100101; // 4677 :  37 - 0x25
      13'h1246: dout <= 8'b01000100; // 4678 :  68 - 0x44
      13'h1247: dout <= 8'b00111000; // 4679 :  56 - 0x38
      13'h1248: dout <= 8'b00000010; // 4680 :   2 - 0x2
      13'h1249: dout <= 8'b00000101; // 4681 :   5 - 0x5
      13'h124A: dout <= 8'b00001011; // 4682 :  11 - 0xb
      13'h124B: dout <= 8'b00001011; // 4683 :  11 - 0xb
      13'h124C: dout <= 8'b00001101; // 4684 :  13 - 0xd
      13'h124D: dout <= 8'b00011000; // 4685 :  24 - 0x18
      13'h124E: dout <= 8'b00111000; // 4686 :  56 - 0x38
      13'h124F: dout <= 8'b00000000; // 4687 :   0 - 0x0
      13'h1250: dout <= 8'b00010000; // 4688 :  16 - 0x10 -- Background 0x25
      13'h1251: dout <= 8'b00010000; // 4689 :  16 - 0x10
      13'h1252: dout <= 8'b00010000; // 4690 :  16 - 0x10
      13'h1253: dout <= 8'b00101100; // 4691 :  44 - 0x2c
      13'h1254: dout <= 8'b01000100; // 4692 :  68 - 0x44
      13'h1255: dout <= 8'b11000100; // 4693 : 196 - 0xc4
      13'h1256: dout <= 8'b00111000; // 4694 :  56 - 0x38
      13'h1257: dout <= 8'b00000000; // 4695 :   0 - 0x0
      13'h1258: dout <= 8'b11100000; // 4696 : 224 - 0xe0
      13'h1259: dout <= 8'b11100000; // 4697 : 224 - 0xe0
      13'h125A: dout <= 8'b11100000; // 4698 : 224 - 0xe0
      13'h125B: dout <= 8'b11010000; // 4699 : 208 - 0xd0
      13'h125C: dout <= 8'b10111000; // 4700 : 184 - 0xb8
      13'h125D: dout <= 8'b00111000; // 4701 :  56 - 0x38
      13'h125E: dout <= 8'b00000000; // 4702 :   0 - 0x0
      13'h125F: dout <= 8'b00000000; // 4703 :   0 - 0x0
      13'h1260: dout <= 8'b00000000; // 4704 :   0 - 0x0 -- Background 0x26
      13'h1261: dout <= 8'b00000000; // 4705 :   0 - 0x0
      13'h1262: dout <= 8'b00000000; // 4706 :   0 - 0x0
      13'h1263: dout <= 8'b00000000; // 4707 :   0 - 0x0
      13'h1264: dout <= 8'b00000000; // 4708 :   0 - 0x0
      13'h1265: dout <= 8'b00000000; // 4709 :   0 - 0x0
      13'h1266: dout <= 8'b00000000; // 4710 :   0 - 0x0
      13'h1267: dout <= 8'b00000000; // 4711 :   0 - 0x0
      13'h1268: dout <= 8'b00000000; // 4712 :   0 - 0x0
      13'h1269: dout <= 8'b00000000; // 4713 :   0 - 0x0
      13'h126A: dout <= 8'b00000000; // 4714 :   0 - 0x0
      13'h126B: dout <= 8'b00000000; // 4715 :   0 - 0x0
      13'h126C: dout <= 8'b00000000; // 4716 :   0 - 0x0
      13'h126D: dout <= 8'b00000000; // 4717 :   0 - 0x0
      13'h126E: dout <= 8'b00000000; // 4718 :   0 - 0x0
      13'h126F: dout <= 8'b00000000; // 4719 :   0 - 0x0
      13'h1270: dout <= 8'b00000000; // 4720 :   0 - 0x0 -- Background 0x27
      13'h1271: dout <= 8'b00000000; // 4721 :   0 - 0x0
      13'h1272: dout <= 8'b00000000; // 4722 :   0 - 0x0
      13'h1273: dout <= 8'b00000000; // 4723 :   0 - 0x0
      13'h1274: dout <= 8'b00000000; // 4724 :   0 - 0x0
      13'h1275: dout <= 8'b00000000; // 4725 :   0 - 0x0
      13'h1276: dout <= 8'b00000000; // 4726 :   0 - 0x0
      13'h1277: dout <= 8'b00000000; // 4727 :   0 - 0x0
      13'h1278: dout <= 8'b00000000; // 4728 :   0 - 0x0
      13'h1279: dout <= 8'b00000000; // 4729 :   0 - 0x0
      13'h127A: dout <= 8'b00000000; // 4730 :   0 - 0x0
      13'h127B: dout <= 8'b00000000; // 4731 :   0 - 0x0
      13'h127C: dout <= 8'b00000000; // 4732 :   0 - 0x0
      13'h127D: dout <= 8'b00000000; // 4733 :   0 - 0x0
      13'h127E: dout <= 8'b00000000; // 4734 :   0 - 0x0
      13'h127F: dout <= 8'b00000000; // 4735 :   0 - 0x0
      13'h1280: dout <= 8'b00000000; // 4736 :   0 - 0x0 -- Background 0x28
      13'h1281: dout <= 8'b00000000; // 4737 :   0 - 0x0
      13'h1282: dout <= 8'b00000000; // 4738 :   0 - 0x0
      13'h1283: dout <= 8'b00000000; // 4739 :   0 - 0x0
      13'h1284: dout <= 8'b00000000; // 4740 :   0 - 0x0
      13'h1285: dout <= 8'b00000000; // 4741 :   0 - 0x0
      13'h1286: dout <= 8'b00000000; // 4742 :   0 - 0x0
      13'h1287: dout <= 8'b00000000; // 4743 :   0 - 0x0
      13'h1288: dout <= 8'b00000000; // 4744 :   0 - 0x0
      13'h1289: dout <= 8'b00000000; // 4745 :   0 - 0x0
      13'h128A: dout <= 8'b00000000; // 4746 :   0 - 0x0
      13'h128B: dout <= 8'b00000000; // 4747 :   0 - 0x0
      13'h128C: dout <= 8'b00000000; // 4748 :   0 - 0x0
      13'h128D: dout <= 8'b00000000; // 4749 :   0 - 0x0
      13'h128E: dout <= 8'b00000000; // 4750 :   0 - 0x0
      13'h128F: dout <= 8'b00000000; // 4751 :   0 - 0x0
      13'h1290: dout <= 8'b00100000; // 4752 :  32 - 0x20 -- Background 0x29
      13'h1291: dout <= 8'b00100000; // 4753 :  32 - 0x20
      13'h1292: dout <= 8'b00100000; // 4754 :  32 - 0x20
      13'h1293: dout <= 8'b00100000; // 4755 :  32 - 0x20
      13'h1294: dout <= 8'b00010011; // 4756 :  19 - 0x13
      13'h1295: dout <= 8'b00001101; // 4757 :  13 - 0xd
      13'h1296: dout <= 8'b00000010; // 4758 :   2 - 0x2
      13'h1297: dout <= 8'b00000001; // 4759 :   1 - 0x1
      13'h1298: dout <= 8'b00011111; // 4760 :  31 - 0x1f
      13'h1299: dout <= 8'b00011111; // 4761 :  31 - 0x1f
      13'h129A: dout <= 8'b00011111; // 4762 :  31 - 0x1f
      13'h129B: dout <= 8'b00011111; // 4763 :  31 - 0x1f
      13'h129C: dout <= 8'b00001100; // 4764 :  12 - 0xc
      13'h129D: dout <= 8'b00000000; // 4765 :   0 - 0x0
      13'h129E: dout <= 8'b00000001; // 4766 :   1 - 0x1
      13'h129F: dout <= 8'b00000000; // 4767 :   0 - 0x0
      13'h12A0: dout <= 8'b00100000; // 4768 :  32 - 0x20 -- Background 0x2a
      13'h12A1: dout <= 8'b00100000; // 4769 :  32 - 0x20
      13'h12A2: dout <= 8'b00100000; // 4770 :  32 - 0x20
      13'h12A3: dout <= 8'b00100000; // 4771 :  32 - 0x20
      13'h12A4: dout <= 8'b00010011; // 4772 :  19 - 0x13
      13'h12A5: dout <= 8'b00001101; // 4773 :  13 - 0xd
      13'h12A6: dout <= 8'b00000001; // 4774 :   1 - 0x1
      13'h12A7: dout <= 8'b00000001; // 4775 :   1 - 0x1
      13'h12A8: dout <= 8'b00011111; // 4776 :  31 - 0x1f
      13'h12A9: dout <= 8'b00011111; // 4777 :  31 - 0x1f
      13'h12AA: dout <= 8'b00011111; // 4778 :  31 - 0x1f
      13'h12AB: dout <= 8'b00011111; // 4779 :  31 - 0x1f
      13'h12AC: dout <= 8'b00001100; // 4780 :  12 - 0xc
      13'h12AD: dout <= 8'b00000000; // 4781 :   0 - 0x0
      13'h12AE: dout <= 8'b00000000; // 4782 :   0 - 0x0
      13'h12AF: dout <= 8'b00000000; // 4783 :   0 - 0x0
      13'h12B0: dout <= 8'b00000000; // 4784 :   0 - 0x0 -- Background 0x2b
      13'h12B1: dout <= 8'b00000000; // 4785 :   0 - 0x0
      13'h12B2: dout <= 8'b00000000; // 4786 :   0 - 0x0
      13'h12B3: dout <= 8'b00000000; // 4787 :   0 - 0x0
      13'h12B4: dout <= 8'b00000000; // 4788 :   0 - 0x0
      13'h12B5: dout <= 8'b00000000; // 4789 :   0 - 0x0
      13'h12B6: dout <= 8'b00000000; // 4790 :   0 - 0x0
      13'h12B7: dout <= 8'b00000000; // 4791 :   0 - 0x0
      13'h12B8: dout <= 8'b00000000; // 4792 :   0 - 0x0
      13'h12B9: dout <= 8'b00000000; // 4793 :   0 - 0x0
      13'h12BA: dout <= 8'b00000000; // 4794 :   0 - 0x0
      13'h12BB: dout <= 8'b00000000; // 4795 :   0 - 0x0
      13'h12BC: dout <= 8'b00000000; // 4796 :   0 - 0x0
      13'h12BD: dout <= 8'b00000000; // 4797 :   0 - 0x0
      13'h12BE: dout <= 8'b00000000; // 4798 :   0 - 0x0
      13'h12BF: dout <= 8'b00000000; // 4799 :   0 - 0x0
      13'h12C0: dout <= 8'b00000000; // 4800 :   0 - 0x0 -- Background 0x2c
      13'h12C1: dout <= 8'b00000000; // 4801 :   0 - 0x0
      13'h12C2: dout <= 8'b00000000; // 4802 :   0 - 0x0
      13'h12C3: dout <= 8'b00000000; // 4803 :   0 - 0x0
      13'h12C4: dout <= 8'b00000000; // 4804 :   0 - 0x0
      13'h12C5: dout <= 8'b00000000; // 4805 :   0 - 0x0
      13'h12C6: dout <= 8'b00000000; // 4806 :   0 - 0x0
      13'h12C7: dout <= 8'b00000000; // 4807 :   0 - 0x0
      13'h12C8: dout <= 8'b00000000; // 4808 :   0 - 0x0
      13'h12C9: dout <= 8'b00000000; // 4809 :   0 - 0x0
      13'h12CA: dout <= 8'b00000000; // 4810 :   0 - 0x0
      13'h12CB: dout <= 8'b00000000; // 4811 :   0 - 0x0
      13'h12CC: dout <= 8'b00000000; // 4812 :   0 - 0x0
      13'h12CD: dout <= 8'b00000000; // 4813 :   0 - 0x0
      13'h12CE: dout <= 8'b00000000; // 4814 :   0 - 0x0
      13'h12CF: dout <= 8'b00000000; // 4815 :   0 - 0x0
      13'h12D0: dout <= 8'b00111100; // 4816 :  60 - 0x3c -- Background 0x2d
      13'h12D1: dout <= 8'b00000000; // 4817 :   0 - 0x0
      13'h12D2: dout <= 8'b10000001; // 4818 : 129 - 0x81
      13'h12D3: dout <= 8'b10011001; // 4819 : 153 - 0x99
      13'h12D4: dout <= 8'b10011001; // 4820 : 153 - 0x99
      13'h12D5: dout <= 8'b10000001; // 4821 : 129 - 0x81
      13'h12D6: dout <= 8'b00000000; // 4822 :   0 - 0x0
      13'h12D7: dout <= 8'b00111100; // 4823 :  60 - 0x3c
      13'h12D8: dout <= 8'b00000000; // 4824 :   0 - 0x0
      13'h12D9: dout <= 8'b01111110; // 4825 : 126 - 0x7e
      13'h12DA: dout <= 8'b01000010; // 4826 :  66 - 0x42
      13'h12DB: dout <= 8'b01000010; // 4827 :  66 - 0x42
      13'h12DC: dout <= 8'b01000010; // 4828 :  66 - 0x42
      13'h12DD: dout <= 8'b01000010; // 4829 :  66 - 0x42
      13'h12DE: dout <= 8'b01111110; // 4830 : 126 - 0x7e
      13'h12DF: dout <= 8'b00000000; // 4831 :   0 - 0x0
      13'h12E0: dout <= 8'b00000000; // 4832 :   0 - 0x0 -- Background 0x2e
      13'h12E1: dout <= 8'b00000000; // 4833 :   0 - 0x0
      13'h12E2: dout <= 8'b00000000; // 4834 :   0 - 0x0
      13'h12E3: dout <= 8'b00000000; // 4835 :   0 - 0x0
      13'h12E4: dout <= 8'b00000000; // 4836 :   0 - 0x0
      13'h12E5: dout <= 8'b00000000; // 4837 :   0 - 0x0
      13'h12E6: dout <= 8'b00000000; // 4838 :   0 - 0x0
      13'h12E7: dout <= 8'b00000000; // 4839 :   0 - 0x0
      13'h12E8: dout <= 8'b00000000; // 4840 :   0 - 0x0
      13'h12E9: dout <= 8'b00000000; // 4841 :   0 - 0x0
      13'h12EA: dout <= 8'b00000000; // 4842 :   0 - 0x0
      13'h12EB: dout <= 8'b00000000; // 4843 :   0 - 0x0
      13'h12EC: dout <= 8'b00000000; // 4844 :   0 - 0x0
      13'h12ED: dout <= 8'b00000000; // 4845 :   0 - 0x0
      13'h12EE: dout <= 8'b00000000; // 4846 :   0 - 0x0
      13'h12EF: dout <= 8'b00000000; // 4847 :   0 - 0x0
      13'h12F0: dout <= 8'b10011111; // 4848 : 159 - 0x9f -- Background 0x2f
      13'h12F1: dout <= 8'b10011110; // 4849 : 158 - 0x9e
      13'h12F2: dout <= 8'b10011100; // 4850 : 156 - 0x9c
      13'h12F3: dout <= 8'b00011000; // 4851 :  24 - 0x18
      13'h12F4: dout <= 8'b00111000; // 4852 :  56 - 0x38
      13'h12F5: dout <= 8'b11111100; // 4853 : 252 - 0xfc
      13'h12F6: dout <= 8'b11111100; // 4854 : 252 - 0xfc
      13'h12F7: dout <= 8'b11111100; // 4855 : 252 - 0xfc
      13'h12F8: dout <= 8'b01100110; // 4856 : 102 - 0x66
      13'h12F9: dout <= 8'b01100000; // 4857 :  96 - 0x60
      13'h12FA: dout <= 8'b01101000; // 4858 : 104 - 0x68
      13'h12FB: dout <= 8'b11100000; // 4859 : 224 - 0xe0
      13'h12FC: dout <= 8'b11000000; // 4860 : 192 - 0xc0
      13'h12FD: dout <= 8'b00010000; // 4861 :  16 - 0x10
      13'h12FE: dout <= 8'b00101000; // 4862 :  40 - 0x28
      13'h12FF: dout <= 8'b01010000; // 4863 :  80 - 0x50
      13'h1300: dout <= 8'b01111111; // 4864 : 127 - 0x7f -- Background 0x30
      13'h1301: dout <= 8'b01111110; // 4865 : 126 - 0x7e
      13'h1302: dout <= 8'b11111100; // 4866 : 252 - 0xfc
      13'h1303: dout <= 8'b00111000; // 4867 :  56 - 0x38
      13'h1304: dout <= 8'b00111000; // 4868 :  56 - 0x38
      13'h1305: dout <= 8'b00000100; // 4869 :   4 - 0x4
      13'h1306: dout <= 8'b10000100; // 4870 : 132 - 0x84
      13'h1307: dout <= 8'b11111100; // 4871 : 252 - 0xfc
      13'h1308: dout <= 8'b11110110; // 4872 : 246 - 0xf6
      13'h1309: dout <= 8'b11110000; // 4873 : 240 - 0xf0
      13'h130A: dout <= 8'b00111000; // 4874 :  56 - 0x38
      13'h130B: dout <= 8'b11010000; // 4875 : 208 - 0xd0
      13'h130C: dout <= 8'b11000000; // 4876 : 192 - 0xc0
      13'h130D: dout <= 8'b11111000; // 4877 : 248 - 0xf8
      13'h130E: dout <= 8'b01111000; // 4878 : 120 - 0x78
      13'h130F: dout <= 8'b00000000; // 4879 :   0 - 0x0
      13'h1310: dout <= 8'b01111111; // 4880 : 127 - 0x7f -- Background 0x31
      13'h1311: dout <= 8'b01111110; // 4881 : 126 - 0x7e
      13'h1312: dout <= 8'b11111100; // 4882 : 252 - 0xfc
      13'h1313: dout <= 8'b00111000; // 4883 :  56 - 0x38
      13'h1314: dout <= 8'b00111000; // 4884 :  56 - 0x38
      13'h1315: dout <= 8'b00011100; // 4885 :  28 - 0x1c
      13'h1316: dout <= 8'b10000100; // 4886 : 132 - 0x84
      13'h1317: dout <= 8'b11000100; // 4887 : 196 - 0xc4
      13'h1318: dout <= 8'b11110110; // 4888 : 246 - 0xf6
      13'h1319: dout <= 8'b11110000; // 4889 : 240 - 0xf0
      13'h131A: dout <= 8'b00111000; // 4890 :  56 - 0x38
      13'h131B: dout <= 8'b11010000; // 4891 : 208 - 0xd0
      13'h131C: dout <= 8'b11000000; // 4892 : 192 - 0xc0
      13'h131D: dout <= 8'b11100000; // 4893 : 224 - 0xe0
      13'h131E: dout <= 8'b01111000; // 4894 : 120 - 0x78
      13'h131F: dout <= 8'b00111000; // 4895 :  56 - 0x38
      13'h1320: dout <= 8'b01111111; // 4896 : 127 - 0x7f -- Background 0x32
      13'h1321: dout <= 8'b01111110; // 4897 : 126 - 0x7e
      13'h1322: dout <= 8'b11111100; // 4898 : 252 - 0xfc
      13'h1323: dout <= 8'b00111000; // 4899 :  56 - 0x38
      13'h1324: dout <= 8'b00100100; // 4900 :  36 - 0x24
      13'h1325: dout <= 8'b00000100; // 4901 :   4 - 0x4
      13'h1326: dout <= 8'b10011100; // 4902 : 156 - 0x9c
      13'h1327: dout <= 8'b11111100; // 4903 : 252 - 0xfc
      13'h1328: dout <= 8'b11110110; // 4904 : 246 - 0xf6
      13'h1329: dout <= 8'b11110000; // 4905 : 240 - 0xf0
      13'h132A: dout <= 8'b00111000; // 4906 :  56 - 0x38
      13'h132B: dout <= 8'b11000000; // 4907 : 192 - 0xc0
      13'h132C: dout <= 8'b11011000; // 4908 : 216 - 0xd8
      13'h132D: dout <= 8'b11111000; // 4909 : 248 - 0xf8
      13'h132E: dout <= 8'b01100000; // 4910 :  96 - 0x60
      13'h132F: dout <= 8'b00010000; // 4911 :  16 - 0x10
      13'h1330: dout <= 8'b00100011; // 4912 :  35 - 0x23 -- Background 0x33
      13'h1331: dout <= 8'b00100011; // 4913 :  35 - 0x23
      13'h1332: dout <= 8'b00100001; // 4914 :  33 - 0x21
      13'h1333: dout <= 8'b00100000; // 4915 :  32 - 0x20
      13'h1334: dout <= 8'b00010011; // 4916 :  19 - 0x13
      13'h1335: dout <= 8'b00001101; // 4917 :  13 - 0xd
      13'h1336: dout <= 8'b00000001; // 4918 :   1 - 0x1
      13'h1337: dout <= 8'b00000001; // 4919 :   1 - 0x1
      13'h1338: dout <= 8'b00011100; // 4920 :  28 - 0x1c
      13'h1339: dout <= 8'b00011100; // 4921 :  28 - 0x1c
      13'h133A: dout <= 8'b00011110; // 4922 :  30 - 0x1e
      13'h133B: dout <= 8'b00011111; // 4923 :  31 - 0x1f
      13'h133C: dout <= 8'b00001100; // 4924 :  12 - 0xc
      13'h133D: dout <= 8'b00000000; // 4925 :   0 - 0x0
      13'h133E: dout <= 8'b00000000; // 4926 :   0 - 0x0
      13'h133F: dout <= 8'b00000000; // 4927 :   0 - 0x0
      13'h1340: dout <= 8'b11111100; // 4928 : 252 - 0xfc -- Background 0x34
      13'h1341: dout <= 8'b11111100; // 4929 : 252 - 0xfc
      13'h1342: dout <= 8'b11111100; // 4930 : 252 - 0xfc
      13'h1343: dout <= 8'b11111100; // 4931 : 252 - 0xfc
      13'h1344: dout <= 8'b10100100; // 4932 : 164 - 0xa4
      13'h1345: dout <= 8'b00100100; // 4933 :  36 - 0x24
      13'h1346: dout <= 8'b00010010; // 4934 :  18 - 0x12
      13'h1347: dout <= 8'b11101110; // 4935 : 238 - 0xee
      13'h1348: dout <= 8'b10000000; // 4936 : 128 - 0x80
      13'h1349: dout <= 8'b01010000; // 4937 :  80 - 0x50
      13'h134A: dout <= 8'b10101000; // 4938 : 168 - 0xa8
      13'h134B: dout <= 8'b00000000; // 4939 :   0 - 0x0
      13'h134C: dout <= 8'b01011000; // 4940 :  88 - 0x58
      13'h134D: dout <= 8'b11011000; // 4941 : 216 - 0xd8
      13'h134E: dout <= 8'b11101100; // 4942 : 236 - 0xec
      13'h134F: dout <= 8'b00000000; // 4943 :   0 - 0x0
      13'h1350: dout <= 8'b00100011; // 4944 :  35 - 0x23 -- Background 0x35
      13'h1351: dout <= 8'b00100011; // 4945 :  35 - 0x23
      13'h1352: dout <= 8'b00100001; // 4946 :  33 - 0x21
      13'h1353: dout <= 8'b00100000; // 4947 :  32 - 0x20
      13'h1354: dout <= 8'b00010011; // 4948 :  19 - 0x13
      13'h1355: dout <= 8'b00001110; // 4949 :  14 - 0xe
      13'h1356: dout <= 8'b00000010; // 4950 :   2 - 0x2
      13'h1357: dout <= 8'b00000001; // 4951 :   1 - 0x1
      13'h1358: dout <= 8'b00011100; // 4952 :  28 - 0x1c
      13'h1359: dout <= 8'b00011100; // 4953 :  28 - 0x1c
      13'h135A: dout <= 8'b00011110; // 4954 :  30 - 0x1e
      13'h135B: dout <= 8'b00011111; // 4955 :  31 - 0x1f
      13'h135C: dout <= 8'b00001100; // 4956 :  12 - 0xc
      13'h135D: dout <= 8'b00000001; // 4957 :   1 - 0x1
      13'h135E: dout <= 8'b00000001; // 4958 :   1 - 0x1
      13'h135F: dout <= 8'b00000000; // 4959 :   0 - 0x0
      13'h1360: dout <= 8'b11111100; // 4960 : 252 - 0xfc -- Background 0x36
      13'h1361: dout <= 8'b11111100; // 4961 : 252 - 0xfc
      13'h1362: dout <= 8'b11111100; // 4962 : 252 - 0xfc
      13'h1363: dout <= 8'b11111100; // 4963 : 252 - 0xfc
      13'h1364: dout <= 8'b10100110; // 4964 : 166 - 0xa6
      13'h1365: dout <= 8'b00110001; // 4965 :  49 - 0x31
      13'h1366: dout <= 8'b01001001; // 4966 :  73 - 0x49
      13'h1367: dout <= 8'b11000110; // 4967 : 198 - 0xc6
      13'h1368: dout <= 8'b10101000; // 4968 : 168 - 0xa8
      13'h1369: dout <= 8'b01010000; // 4969 :  80 - 0x50
      13'h136A: dout <= 8'b10101000; // 4970 : 168 - 0xa8
      13'h136B: dout <= 8'b00000000; // 4971 :   0 - 0x0
      13'h136C: dout <= 8'b01011000; // 4972 :  88 - 0x58
      13'h136D: dout <= 8'b11001110; // 4973 : 206 - 0xce
      13'h136E: dout <= 8'b10000110; // 4974 : 134 - 0x86
      13'h136F: dout <= 8'b00000000; // 4975 :   0 - 0x0
      13'h1370: dout <= 8'b11111100; // 4976 : 252 - 0xfc -- Background 0x37
      13'h1371: dout <= 8'b11111100; // 4977 : 252 - 0xfc
      13'h1372: dout <= 8'b11111100; // 4978 : 252 - 0xfc
      13'h1373: dout <= 8'b11111100; // 4979 : 252 - 0xfc
      13'h1374: dout <= 8'b10100100; // 4980 : 164 - 0xa4
      13'h1375: dout <= 8'b00100100; // 4981 :  36 - 0x24
      13'h1376: dout <= 8'b00010010; // 4982 :  18 - 0x12
      13'h1377: dout <= 8'b11101110; // 4983 : 238 - 0xee
      13'h1378: dout <= 8'b10101000; // 4984 : 168 - 0xa8
      13'h1379: dout <= 8'b01010000; // 4985 :  80 - 0x50
      13'h137A: dout <= 8'b10101000; // 4986 : 168 - 0xa8
      13'h137B: dout <= 8'b00000000; // 4987 :   0 - 0x0
      13'h137C: dout <= 8'b01011000; // 4988 :  88 - 0x58
      13'h137D: dout <= 8'b11011000; // 4989 : 216 - 0xd8
      13'h137E: dout <= 8'b11101100; // 4990 : 236 - 0xec
      13'h137F: dout <= 8'b00000000; // 4991 :   0 - 0x0
      13'h1380: dout <= 8'b00000000; // 4992 :   0 - 0x0 -- Background 0x38
      13'h1381: dout <= 8'b00000000; // 4993 :   0 - 0x0
      13'h1382: dout <= 8'b00000000; // 4994 :   0 - 0x0
      13'h1383: dout <= 8'b00000000; // 4995 :   0 - 0x0
      13'h1384: dout <= 8'b00000000; // 4996 :   0 - 0x0
      13'h1385: dout <= 8'b00000000; // 4997 :   0 - 0x0
      13'h1386: dout <= 8'b00000000; // 4998 :   0 - 0x0
      13'h1387: dout <= 8'b00000000; // 4999 :   0 - 0x0
      13'h1388: dout <= 8'b00000000; // 5000 :   0 - 0x0
      13'h1389: dout <= 8'b00000000; // 5001 :   0 - 0x0
      13'h138A: dout <= 8'b00000000; // 5002 :   0 - 0x0
      13'h138B: dout <= 8'b00000000; // 5003 :   0 - 0x0
      13'h138C: dout <= 8'b00000000; // 5004 :   0 - 0x0
      13'h138D: dout <= 8'b00000000; // 5005 :   0 - 0x0
      13'h138E: dout <= 8'b00000000; // 5006 :   0 - 0x0
      13'h138F: dout <= 8'b00000000; // 5007 :   0 - 0x0
      13'h1390: dout <= 8'b00000000; // 5008 :   0 - 0x0 -- Background 0x39
      13'h1391: dout <= 8'b00000000; // 5009 :   0 - 0x0
      13'h1392: dout <= 8'b00000000; // 5010 :   0 - 0x0
      13'h1393: dout <= 8'b00000000; // 5011 :   0 - 0x0
      13'h1394: dout <= 8'b00000000; // 5012 :   0 - 0x0
      13'h1395: dout <= 8'b00000000; // 5013 :   0 - 0x0
      13'h1396: dout <= 8'b00000000; // 5014 :   0 - 0x0
      13'h1397: dout <= 8'b00000000; // 5015 :   0 - 0x0
      13'h1398: dout <= 8'b00000000; // 5016 :   0 - 0x0
      13'h1399: dout <= 8'b00000000; // 5017 :   0 - 0x0
      13'h139A: dout <= 8'b00000000; // 5018 :   0 - 0x0
      13'h139B: dout <= 8'b00000000; // 5019 :   0 - 0x0
      13'h139C: dout <= 8'b00000000; // 5020 :   0 - 0x0
      13'h139D: dout <= 8'b00000000; // 5021 :   0 - 0x0
      13'h139E: dout <= 8'b00000000; // 5022 :   0 - 0x0
      13'h139F: dout <= 8'b00000000; // 5023 :   0 - 0x0
      13'h13A0: dout <= 8'b00000000; // 5024 :   0 - 0x0 -- Background 0x3a
      13'h13A1: dout <= 8'b00000000; // 5025 :   0 - 0x0
      13'h13A2: dout <= 8'b00000000; // 5026 :   0 - 0x0
      13'h13A3: dout <= 8'b00000000; // 5027 :   0 - 0x0
      13'h13A4: dout <= 8'b00000000; // 5028 :   0 - 0x0
      13'h13A5: dout <= 8'b00000000; // 5029 :   0 - 0x0
      13'h13A6: dout <= 8'b00000000; // 5030 :   0 - 0x0
      13'h13A7: dout <= 8'b00000000; // 5031 :   0 - 0x0
      13'h13A8: dout <= 8'b00000000; // 5032 :   0 - 0x0
      13'h13A9: dout <= 8'b00000000; // 5033 :   0 - 0x0
      13'h13AA: dout <= 8'b00000000; // 5034 :   0 - 0x0
      13'h13AB: dout <= 8'b00000000; // 5035 :   0 - 0x0
      13'h13AC: dout <= 8'b00000000; // 5036 :   0 - 0x0
      13'h13AD: dout <= 8'b00000000; // 5037 :   0 - 0x0
      13'h13AE: dout <= 8'b00000000; // 5038 :   0 - 0x0
      13'h13AF: dout <= 8'b00000000; // 5039 :   0 - 0x0
      13'h13B0: dout <= 8'b00000000; // 5040 :   0 - 0x0 -- Background 0x3b
      13'h13B1: dout <= 8'b00000000; // 5041 :   0 - 0x0
      13'h13B2: dout <= 8'b00000000; // 5042 :   0 - 0x0
      13'h13B3: dout <= 8'b00000000; // 5043 :   0 - 0x0
      13'h13B4: dout <= 8'b00000000; // 5044 :   0 - 0x0
      13'h13B5: dout <= 8'b00000000; // 5045 :   0 - 0x0
      13'h13B6: dout <= 8'b00000000; // 5046 :   0 - 0x0
      13'h13B7: dout <= 8'b00000000; // 5047 :   0 - 0x0
      13'h13B8: dout <= 8'b00000000; // 5048 :   0 - 0x0
      13'h13B9: dout <= 8'b00000000; // 5049 :   0 - 0x0
      13'h13BA: dout <= 8'b00000000; // 5050 :   0 - 0x0
      13'h13BB: dout <= 8'b00000000; // 5051 :   0 - 0x0
      13'h13BC: dout <= 8'b00000000; // 5052 :   0 - 0x0
      13'h13BD: dout <= 8'b00000000; // 5053 :   0 - 0x0
      13'h13BE: dout <= 8'b00000000; // 5054 :   0 - 0x0
      13'h13BF: dout <= 8'b00000000; // 5055 :   0 - 0x0
      13'h13C0: dout <= 8'b00000000; // 5056 :   0 - 0x0 -- Background 0x3c
      13'h13C1: dout <= 8'b00000000; // 5057 :   0 - 0x0
      13'h13C2: dout <= 8'b00000000; // 5058 :   0 - 0x0
      13'h13C3: dout <= 8'b00000000; // 5059 :   0 - 0x0
      13'h13C4: dout <= 8'b00000000; // 5060 :   0 - 0x0
      13'h13C5: dout <= 8'b00000000; // 5061 :   0 - 0x0
      13'h13C6: dout <= 8'b00000000; // 5062 :   0 - 0x0
      13'h13C7: dout <= 8'b00000000; // 5063 :   0 - 0x0
      13'h13C8: dout <= 8'b00000000; // 5064 :   0 - 0x0
      13'h13C9: dout <= 8'b00000000; // 5065 :   0 - 0x0
      13'h13CA: dout <= 8'b00000000; // 5066 :   0 - 0x0
      13'h13CB: dout <= 8'b00000000; // 5067 :   0 - 0x0
      13'h13CC: dout <= 8'b00000000; // 5068 :   0 - 0x0
      13'h13CD: dout <= 8'b00000000; // 5069 :   0 - 0x0
      13'h13CE: dout <= 8'b00000000; // 5070 :   0 - 0x0
      13'h13CF: dout <= 8'b00000000; // 5071 :   0 - 0x0
      13'h13D0: dout <= 8'b00000000; // 5072 :   0 - 0x0 -- Background 0x3d
      13'h13D1: dout <= 8'b00000000; // 5073 :   0 - 0x0
      13'h13D2: dout <= 8'b00000000; // 5074 :   0 - 0x0
      13'h13D3: dout <= 8'b00000000; // 5075 :   0 - 0x0
      13'h13D4: dout <= 8'b00000000; // 5076 :   0 - 0x0
      13'h13D5: dout <= 8'b00000000; // 5077 :   0 - 0x0
      13'h13D6: dout <= 8'b00000000; // 5078 :   0 - 0x0
      13'h13D7: dout <= 8'b00000000; // 5079 :   0 - 0x0
      13'h13D8: dout <= 8'b00000000; // 5080 :   0 - 0x0
      13'h13D9: dout <= 8'b00000000; // 5081 :   0 - 0x0
      13'h13DA: dout <= 8'b00000000; // 5082 :   0 - 0x0
      13'h13DB: dout <= 8'b00000000; // 5083 :   0 - 0x0
      13'h13DC: dout <= 8'b00000000; // 5084 :   0 - 0x0
      13'h13DD: dout <= 8'b00000000; // 5085 :   0 - 0x0
      13'h13DE: dout <= 8'b00000000; // 5086 :   0 - 0x0
      13'h13DF: dout <= 8'b00000000; // 5087 :   0 - 0x0
      13'h13E0: dout <= 8'b00000000; // 5088 :   0 - 0x0 -- Background 0x3e
      13'h13E1: dout <= 8'b00000000; // 5089 :   0 - 0x0
      13'h13E2: dout <= 8'b00000000; // 5090 :   0 - 0x0
      13'h13E3: dout <= 8'b00000000; // 5091 :   0 - 0x0
      13'h13E4: dout <= 8'b00000000; // 5092 :   0 - 0x0
      13'h13E5: dout <= 8'b00000000; // 5093 :   0 - 0x0
      13'h13E6: dout <= 8'b00000000; // 5094 :   0 - 0x0
      13'h13E7: dout <= 8'b00000000; // 5095 :   0 - 0x0
      13'h13E8: dout <= 8'b00000000; // 5096 :   0 - 0x0
      13'h13E9: dout <= 8'b00000000; // 5097 :   0 - 0x0
      13'h13EA: dout <= 8'b00000000; // 5098 :   0 - 0x0
      13'h13EB: dout <= 8'b00000000; // 5099 :   0 - 0x0
      13'h13EC: dout <= 8'b00000000; // 5100 :   0 - 0x0
      13'h13ED: dout <= 8'b00000000; // 5101 :   0 - 0x0
      13'h13EE: dout <= 8'b00000000; // 5102 :   0 - 0x0
      13'h13EF: dout <= 8'b00000000; // 5103 :   0 - 0x0
      13'h13F0: dout <= 8'b00000000; // 5104 :   0 - 0x0 -- Background 0x3f
      13'h13F1: dout <= 8'b00000000; // 5105 :   0 - 0x0
      13'h13F2: dout <= 8'b00000000; // 5106 :   0 - 0x0
      13'h13F3: dout <= 8'b00000000; // 5107 :   0 - 0x0
      13'h13F4: dout <= 8'b00000000; // 5108 :   0 - 0x0
      13'h13F5: dout <= 8'b00000000; // 5109 :   0 - 0x0
      13'h13F6: dout <= 8'b00000000; // 5110 :   0 - 0x0
      13'h13F7: dout <= 8'b00000000; // 5111 :   0 - 0x0
      13'h13F8: dout <= 8'b00000000; // 5112 :   0 - 0x0
      13'h13F9: dout <= 8'b00000000; // 5113 :   0 - 0x0
      13'h13FA: dout <= 8'b00000000; // 5114 :   0 - 0x0
      13'h13FB: dout <= 8'b00000000; // 5115 :   0 - 0x0
      13'h13FC: dout <= 8'b00000000; // 5116 :   0 - 0x0
      13'h13FD: dout <= 8'b00000000; // 5117 :   0 - 0x0
      13'h13FE: dout <= 8'b00000000; // 5118 :   0 - 0x0
      13'h13FF: dout <= 8'b00000000; // 5119 :   0 - 0x0
      13'h1400: dout <= 8'b00000000; // 5120 :   0 - 0x0 -- Background 0x40
      13'h1401: dout <= 8'b00111110; // 5121 :  62 - 0x3e
      13'h1402: dout <= 8'b01111111; // 5122 : 127 - 0x7f
      13'h1403: dout <= 8'b01111111; // 5123 : 127 - 0x7f
      13'h1404: dout <= 8'b01111111; // 5124 : 127 - 0x7f
      13'h1405: dout <= 8'b01111111; // 5125 : 127 - 0x7f
      13'h1406: dout <= 8'b01111111; // 5126 : 127 - 0x7f
      13'h1407: dout <= 8'b00111110; // 5127 :  62 - 0x3e
      13'h1408: dout <= 8'b00111100; // 5128 :  60 - 0x3c
      13'h1409: dout <= 8'b01111100; // 5129 : 124 - 0x7c
      13'h140A: dout <= 8'b11100110; // 5130 : 230 - 0xe6
      13'h140B: dout <= 8'b11101110; // 5131 : 238 - 0xee
      13'h140C: dout <= 8'b11110110; // 5132 : 246 - 0xf6
      13'h140D: dout <= 8'b11100110; // 5133 : 230 - 0xe6
      13'h140E: dout <= 8'b00111100; // 5134 :  60 - 0x3c
      13'h140F: dout <= 8'b00000000; // 5135 :   0 - 0x0
      13'h1410: dout <= 8'b00000000; // 5136 :   0 - 0x0 -- Background 0x41
      13'h1411: dout <= 8'b00111100; // 5137 :  60 - 0x3c
      13'h1412: dout <= 8'b00011100; // 5138 :  28 - 0x1c
      13'h1413: dout <= 8'b00011100; // 5139 :  28 - 0x1c
      13'h1414: dout <= 8'b00011100; // 5140 :  28 - 0x1c
      13'h1415: dout <= 8'b00011100; // 5141 :  28 - 0x1c
      13'h1416: dout <= 8'b00011100; // 5142 :  28 - 0x1c
      13'h1417: dout <= 8'b00011100; // 5143 :  28 - 0x1c
      13'h1418: dout <= 8'b00111000; // 5144 :  56 - 0x38
      13'h1419: dout <= 8'b01111000; // 5145 : 120 - 0x78
      13'h141A: dout <= 8'b00111000; // 5146 :  56 - 0x38
      13'h141B: dout <= 8'b00111000; // 5147 :  56 - 0x38
      13'h141C: dout <= 8'b00111000; // 5148 :  56 - 0x38
      13'h141D: dout <= 8'b00111000; // 5149 :  56 - 0x38
      13'h141E: dout <= 8'b00111000; // 5150 :  56 - 0x38
      13'h141F: dout <= 8'b00000000; // 5151 :   0 - 0x0
      13'h1420: dout <= 8'b00000000; // 5152 :   0 - 0x0 -- Background 0x42
      13'h1421: dout <= 8'b01111100; // 5153 : 124 - 0x7c
      13'h1422: dout <= 8'b01111111; // 5154 : 127 - 0x7f
      13'h1423: dout <= 8'b01100111; // 5155 : 103 - 0x67
      13'h1424: dout <= 8'b00111111; // 5156 :  63 - 0x3f
      13'h1425: dout <= 8'b01111110; // 5157 : 126 - 0x7e
      13'h1426: dout <= 8'b01111111; // 5158 : 127 - 0x7f
      13'h1427: dout <= 8'b01111111; // 5159 : 127 - 0x7f
      13'h1428: dout <= 8'b01111100; // 5160 : 124 - 0x7c
      13'h1429: dout <= 8'b11111110; // 5161 : 254 - 0xfe
      13'h142A: dout <= 8'b11100110; // 5162 : 230 - 0xe6
      13'h142B: dout <= 8'b00011110; // 5163 :  30 - 0x1e
      13'h142C: dout <= 8'b01111100; // 5164 : 124 - 0x7c
      13'h142D: dout <= 8'b11100000; // 5165 : 224 - 0xe0
      13'h142E: dout <= 8'b11111110; // 5166 : 254 - 0xfe
      13'h142F: dout <= 8'b00000000; // 5167 :   0 - 0x0
      13'h1430: dout <= 8'b00000000; // 5168 :   0 - 0x0 -- Background 0x43
      13'h1431: dout <= 8'b01111110; // 5169 : 126 - 0x7e
      13'h1432: dout <= 8'b01111111; // 5170 : 127 - 0x7f
      13'h1433: dout <= 8'b01111111; // 5171 : 127 - 0x7f
      13'h1434: dout <= 8'b00011111; // 5172 :  31 - 0x1f
      13'h1435: dout <= 8'b01110111; // 5173 : 119 - 0x77
      13'h1436: dout <= 8'b01111111; // 5174 : 127 - 0x7f
      13'h1437: dout <= 8'b01111110; // 5175 : 126 - 0x7e
      13'h1438: dout <= 8'b01111100; // 5176 : 124 - 0x7c
      13'h1439: dout <= 8'b11111100; // 5177 : 252 - 0xfc
      13'h143A: dout <= 8'b11100110; // 5178 : 230 - 0xe6
      13'h143B: dout <= 8'b00011100; // 5179 :  28 - 0x1c
      13'h143C: dout <= 8'b01100110; // 5180 : 102 - 0x66
      13'h143D: dout <= 8'b11101110; // 5181 : 238 - 0xee
      13'h143E: dout <= 8'b11111100; // 5182 : 252 - 0xfc
      13'h143F: dout <= 8'b00000000; // 5183 :   0 - 0x0
      13'h1440: dout <= 8'b00000000; // 5184 :   0 - 0x0 -- Background 0x44
      13'h1441: dout <= 8'b00001110; // 5185 :  14 - 0xe
      13'h1442: dout <= 8'b00011110; // 5186 :  30 - 0x1e
      13'h1443: dout <= 8'b00111110; // 5187 :  62 - 0x3e
      13'h1444: dout <= 8'b01111110; // 5188 : 126 - 0x7e
      13'h1445: dout <= 8'b01111111; // 5189 : 127 - 0x7f
      13'h1446: dout <= 8'b01111110; // 5190 : 126 - 0x7e
      13'h1447: dout <= 8'b00001100; // 5191 :  12 - 0xc
      13'h1448: dout <= 8'b00001100; // 5192 :  12 - 0xc
      13'h1449: dout <= 8'b00011100; // 5193 :  28 - 0x1c
      13'h144A: dout <= 8'b00111100; // 5194 :  60 - 0x3c
      13'h144B: dout <= 8'b01111100; // 5195 : 124 - 0x7c
      13'h144C: dout <= 8'b11101100; // 5196 : 236 - 0xec
      13'h144D: dout <= 8'b11111110; // 5197 : 254 - 0xfe
      13'h144E: dout <= 8'b00001100; // 5198 :  12 - 0xc
      13'h144F: dout <= 8'b00000000; // 5199 :   0 - 0x0
      13'h1450: dout <= 8'b00000000; // 5200 :   0 - 0x0 -- Background 0x45
      13'h1451: dout <= 8'b01111111; // 5201 : 127 - 0x7f
      13'h1452: dout <= 8'b01111111; // 5202 : 127 - 0x7f
      13'h1453: dout <= 8'b01111111; // 5203 : 127 - 0x7f
      13'h1454: dout <= 8'b01111111; // 5204 : 127 - 0x7f
      13'h1455: dout <= 8'b01110111; // 5205 : 119 - 0x77
      13'h1456: dout <= 8'b01111111; // 5206 : 127 - 0x7f
      13'h1457: dout <= 8'b01111110; // 5207 : 126 - 0x7e
      13'h1458: dout <= 8'b11111110; // 5208 : 254 - 0xfe
      13'h1459: dout <= 8'b11111110; // 5209 : 254 - 0xfe
      13'h145A: dout <= 8'b11100000; // 5210 : 224 - 0xe0
      13'h145B: dout <= 8'b11111110; // 5211 : 254 - 0xfe
      13'h145C: dout <= 8'b00000110; // 5212 :   6 - 0x6
      13'h145D: dout <= 8'b11101110; // 5213 : 238 - 0xee
      13'h145E: dout <= 8'b11111100; // 5214 : 252 - 0xfc
      13'h145F: dout <= 8'b00000000; // 5215 :   0 - 0x0
      13'h1460: dout <= 8'b00000000; // 5216 :   0 - 0x0 -- Background 0x46
      13'h1461: dout <= 8'b00111110; // 5217 :  62 - 0x3e
      13'h1462: dout <= 8'b01111110; // 5218 : 126 - 0x7e
      13'h1463: dout <= 8'b01111111; // 5219 : 127 - 0x7f
      13'h1464: dout <= 8'b01111111; // 5220 : 127 - 0x7f
      13'h1465: dout <= 8'b01110111; // 5221 : 119 - 0x77
      13'h1466: dout <= 8'b01111111; // 5222 : 127 - 0x7f
      13'h1467: dout <= 8'b00111110; // 5223 :  62 - 0x3e
      13'h1468: dout <= 8'b00111100; // 5224 :  60 - 0x3c
      13'h1469: dout <= 8'b01111100; // 5225 : 124 - 0x7c
      13'h146A: dout <= 8'b11100000; // 5226 : 224 - 0xe0
      13'h146B: dout <= 8'b11111110; // 5227 : 254 - 0xfe
      13'h146C: dout <= 8'b11100110; // 5228 : 230 - 0xe6
      13'h146D: dout <= 8'b11101110; // 5229 : 238 - 0xee
      13'h146E: dout <= 8'b00111100; // 5230 :  60 - 0x3c
      13'h146F: dout <= 8'b00000000; // 5231 :   0 - 0x0
      13'h1470: dout <= 8'b00000000; // 5232 :   0 - 0x0 -- Background 0x47
      13'h1471: dout <= 8'b01111110; // 5233 : 126 - 0x7e
      13'h1472: dout <= 8'b01111110; // 5234 : 126 - 0x7e
      13'h1473: dout <= 8'b00011110; // 5235 :  30 - 0x1e
      13'h1474: dout <= 8'b00011100; // 5236 :  28 - 0x1c
      13'h1475: dout <= 8'b00111100; // 5237 :  60 - 0x3c
      13'h1476: dout <= 8'b00111000; // 5238 :  56 - 0x38
      13'h1477: dout <= 8'b00111000; // 5239 :  56 - 0x38
      13'h1478: dout <= 8'b11111110; // 5240 : 254 - 0xfe
      13'h1479: dout <= 8'b11111100; // 5241 : 252 - 0xfc
      13'h147A: dout <= 8'b00001100; // 5242 :  12 - 0xc
      13'h147B: dout <= 8'b00111000; // 5243 :  56 - 0x38
      13'h147C: dout <= 8'b00111000; // 5244 :  56 - 0x38
      13'h147D: dout <= 8'b01110000; // 5245 : 112 - 0x70
      13'h147E: dout <= 8'b01110000; // 5246 : 112 - 0x70
      13'h147F: dout <= 8'b00000000; // 5247 :   0 - 0x0
      13'h1480: dout <= 8'b00000000; // 5248 :   0 - 0x0 -- Background 0x48
      13'h1481: dout <= 8'b00111110; // 5249 :  62 - 0x3e
      13'h1482: dout <= 8'b01111111; // 5250 : 127 - 0x7f
      13'h1483: dout <= 8'b01111111; // 5251 : 127 - 0x7f
      13'h1484: dout <= 8'b01111111; // 5252 : 127 - 0x7f
      13'h1485: dout <= 8'b01111111; // 5253 : 127 - 0x7f
      13'h1486: dout <= 8'b01111111; // 5254 : 127 - 0x7f
      13'h1487: dout <= 8'b00111110; // 5255 :  62 - 0x3e
      13'h1488: dout <= 8'b00111110; // 5256 :  62 - 0x3e
      13'h1489: dout <= 8'b01111100; // 5257 : 124 - 0x7c
      13'h148A: dout <= 8'b11100110; // 5258 : 230 - 0xe6
      13'h148B: dout <= 8'b10111100; // 5259 : 188 - 0xbc
      13'h148C: dout <= 8'b11100110; // 5260 : 230 - 0xe6
      13'h148D: dout <= 8'b11101110; // 5261 : 238 - 0xee
      13'h148E: dout <= 8'b00111100; // 5262 :  60 - 0x3c
      13'h148F: dout <= 8'b00000000; // 5263 :   0 - 0x0
      13'h1490: dout <= 8'b00000000; // 5264 :   0 - 0x0 -- Background 0x49
      13'h1491: dout <= 8'b00111110; // 5265 :  62 - 0x3e
      13'h1492: dout <= 8'b01111111; // 5266 : 127 - 0x7f
      13'h1493: dout <= 8'b01110111; // 5267 : 119 - 0x77
      13'h1494: dout <= 8'b01111111; // 5268 : 127 - 0x7f
      13'h1495: dout <= 8'b01111111; // 5269 : 127 - 0x7f
      13'h1496: dout <= 8'b00111111; // 5270 :  63 - 0x3f
      13'h1497: dout <= 8'b00111110; // 5271 :  62 - 0x3e
      13'h1498: dout <= 8'b00111100; // 5272 :  60 - 0x3c
      13'h1499: dout <= 8'b01111100; // 5273 : 124 - 0x7c
      13'h149A: dout <= 8'b11100110; // 5274 : 230 - 0xe6
      13'h149B: dout <= 8'b11101110; // 5275 : 238 - 0xee
      13'h149C: dout <= 8'b11111110; // 5276 : 254 - 0xfe
      13'h149D: dout <= 8'b10000110; // 5277 : 134 - 0x86
      13'h149E: dout <= 8'b01111100; // 5278 : 124 - 0x7c
      13'h149F: dout <= 8'b01000000; // 5279 :  64 - 0x40
      13'h14A0: dout <= 8'b11111111; // 5280 : 255 - 0xff -- Background 0x4a
      13'h14A1: dout <= 8'b10011001; // 5281 : 153 - 0x99
      13'h14A2: dout <= 8'b10011001; // 5282 : 153 - 0x99
      13'h14A3: dout <= 8'b10011001; // 5283 : 153 - 0x99
      13'h14A4: dout <= 8'b10011001; // 5284 : 153 - 0x99
      13'h14A5: dout <= 8'b10011001; // 5285 : 153 - 0x99
      13'h14A6: dout <= 8'b10011001; // 5286 : 153 - 0x99
      13'h14A7: dout <= 8'b11111111; // 5287 : 255 - 0xff
      13'h14A8: dout <= 8'b11101110; // 5288 : 238 - 0xee
      13'h14A9: dout <= 8'b11101110; // 5289 : 238 - 0xee
      13'h14AA: dout <= 8'b11101110; // 5290 : 238 - 0xee
      13'h14AB: dout <= 8'b11101110; // 5291 : 238 - 0xee
      13'h14AC: dout <= 8'b11101110; // 5292 : 238 - 0xee
      13'h14AD: dout <= 8'b11101110; // 5293 : 238 - 0xee
      13'h14AE: dout <= 8'b11101110; // 5294 : 238 - 0xee
      13'h14AF: dout <= 8'b10001000; // 5295 : 136 - 0x88
      13'h14B0: dout <= 8'b11110000; // 5296 : 240 - 0xf0 -- Background 0x4b
      13'h14B1: dout <= 8'b10010000; // 5297 : 144 - 0x90
      13'h14B2: dout <= 8'b10010000; // 5298 : 144 - 0x90
      13'h14B3: dout <= 8'b10010000; // 5299 : 144 - 0x90
      13'h14B4: dout <= 8'b10010000; // 5300 : 144 - 0x90
      13'h14B5: dout <= 8'b10010000; // 5301 : 144 - 0x90
      13'h14B6: dout <= 8'b10010000; // 5302 : 144 - 0x90
      13'h14B7: dout <= 8'b11110000; // 5303 : 240 - 0xf0
      13'h14B8: dout <= 8'b11100000; // 5304 : 224 - 0xe0
      13'h14B9: dout <= 8'b11100000; // 5305 : 224 - 0xe0
      13'h14BA: dout <= 8'b11100000; // 5306 : 224 - 0xe0
      13'h14BB: dout <= 8'b11100000; // 5307 : 224 - 0xe0
      13'h14BC: dout <= 8'b11100000; // 5308 : 224 - 0xe0
      13'h14BD: dout <= 8'b11100000; // 5309 : 224 - 0xe0
      13'h14BE: dout <= 8'b11100000; // 5310 : 224 - 0xe0
      13'h14BF: dout <= 8'b10000000; // 5311 : 128 - 0x80
      13'h14C0: dout <= 8'b11111111; // 5312 : 255 - 0xff -- Background 0x4c
      13'h14C1: dout <= 8'b11111111; // 5313 : 255 - 0xff
      13'h14C2: dout <= 8'b11111111; // 5314 : 255 - 0xff
      13'h14C3: dout <= 8'b11111111; // 5315 : 255 - 0xff
      13'h14C4: dout <= 8'b11111111; // 5316 : 255 - 0xff
      13'h14C5: dout <= 8'b11111111; // 5317 : 255 - 0xff
      13'h14C6: dout <= 8'b11111111; // 5318 : 255 - 0xff
      13'h14C7: dout <= 8'b11111111; // 5319 : 255 - 0xff
      13'h14C8: dout <= 8'b00000000; // 5320 :   0 - 0x0
      13'h14C9: dout <= 8'b01111111; // 5321 : 127 - 0x7f
      13'h14CA: dout <= 8'b01111111; // 5322 : 127 - 0x7f
      13'h14CB: dout <= 8'b01111111; // 5323 : 127 - 0x7f
      13'h14CC: dout <= 8'b01111111; // 5324 : 127 - 0x7f
      13'h14CD: dout <= 8'b01111111; // 5325 : 127 - 0x7f
      13'h14CE: dout <= 8'b01111111; // 5326 : 127 - 0x7f
      13'h14CF: dout <= 8'b01111111; // 5327 : 127 - 0x7f
      13'h14D0: dout <= 8'b11111111; // 5328 : 255 - 0xff -- Background 0x4d
      13'h14D1: dout <= 8'b11111111; // 5329 : 255 - 0xff
      13'h14D2: dout <= 8'b11111111; // 5330 : 255 - 0xff
      13'h14D3: dout <= 8'b11111111; // 5331 : 255 - 0xff
      13'h14D4: dout <= 8'b11111111; // 5332 : 255 - 0xff
      13'h14D5: dout <= 8'b11111111; // 5333 : 255 - 0xff
      13'h14D6: dout <= 8'b11111111; // 5334 : 255 - 0xff
      13'h14D7: dout <= 8'b11111111; // 5335 : 255 - 0xff
      13'h14D8: dout <= 8'b01111111; // 5336 : 127 - 0x7f
      13'h14D9: dout <= 8'b01111111; // 5337 : 127 - 0x7f
      13'h14DA: dout <= 8'b01111111; // 5338 : 127 - 0x7f
      13'h14DB: dout <= 8'b01111111; // 5339 : 127 - 0x7f
      13'h14DC: dout <= 8'b01111111; // 5340 : 127 - 0x7f
      13'h14DD: dout <= 8'b01111111; // 5341 : 127 - 0x7f
      13'h14DE: dout <= 8'b01111111; // 5342 : 127 - 0x7f
      13'h14DF: dout <= 8'b00000000; // 5343 :   0 - 0x0
      13'h14E0: dout <= 8'b11111111; // 5344 : 255 - 0xff -- Background 0x4e
      13'h14E1: dout <= 8'b11111111; // 5345 : 255 - 0xff
      13'h14E2: dout <= 8'b11111111; // 5346 : 255 - 0xff
      13'h14E3: dout <= 8'b11111111; // 5347 : 255 - 0xff
      13'h14E4: dout <= 8'b11111111; // 5348 : 255 - 0xff
      13'h14E5: dout <= 8'b11111111; // 5349 : 255 - 0xff
      13'h14E6: dout <= 8'b11111111; // 5350 : 255 - 0xff
      13'h14E7: dout <= 8'b11111111; // 5351 : 255 - 0xff
      13'h14E8: dout <= 8'b00000000; // 5352 :   0 - 0x0
      13'h14E9: dout <= 8'b11111110; // 5353 : 254 - 0xfe
      13'h14EA: dout <= 8'b11111110; // 5354 : 254 - 0xfe
      13'h14EB: dout <= 8'b11111110; // 5355 : 254 - 0xfe
      13'h14EC: dout <= 8'b11111110; // 5356 : 254 - 0xfe
      13'h14ED: dout <= 8'b11111110; // 5357 : 254 - 0xfe
      13'h14EE: dout <= 8'b11111110; // 5358 : 254 - 0xfe
      13'h14EF: dout <= 8'b11111110; // 5359 : 254 - 0xfe
      13'h14F0: dout <= 8'b11111111; // 5360 : 255 - 0xff -- Background 0x4f
      13'h14F1: dout <= 8'b11111111; // 5361 : 255 - 0xff
      13'h14F2: dout <= 8'b11111111; // 5362 : 255 - 0xff
      13'h14F3: dout <= 8'b11111111; // 5363 : 255 - 0xff
      13'h14F4: dout <= 8'b11111111; // 5364 : 255 - 0xff
      13'h14F5: dout <= 8'b11111111; // 5365 : 255 - 0xff
      13'h14F6: dout <= 8'b11111111; // 5366 : 255 - 0xff
      13'h14F7: dout <= 8'b11111111; // 5367 : 255 - 0xff
      13'h14F8: dout <= 8'b11111110; // 5368 : 254 - 0xfe
      13'h14F9: dout <= 8'b11111110; // 5369 : 254 - 0xfe
      13'h14FA: dout <= 8'b11111110; // 5370 : 254 - 0xfe
      13'h14FB: dout <= 8'b11111110; // 5371 : 254 - 0xfe
      13'h14FC: dout <= 8'b11111110; // 5372 : 254 - 0xfe
      13'h14FD: dout <= 8'b11111110; // 5373 : 254 - 0xfe
      13'h14FE: dout <= 8'b11111110; // 5374 : 254 - 0xfe
      13'h14FF: dout <= 8'b00000000; // 5375 :   0 - 0x0
      13'h1500: dout <= 8'b00010000; // 5376 :  16 - 0x10 -- Background 0x50
      13'h1501: dout <= 8'b00101000; // 5377 :  40 - 0x28
      13'h1502: dout <= 8'b11101110; // 5378 : 238 - 0xee
      13'h1503: dout <= 8'b10000010; // 5379 : 130 - 0x82
      13'h1504: dout <= 8'b01000100; // 5380 :  68 - 0x44
      13'h1505: dout <= 8'b01000100; // 5381 :  68 - 0x44
      13'h1506: dout <= 8'b10010010; // 5382 : 146 - 0x92
      13'h1507: dout <= 8'b11101110; // 5383 : 238 - 0xee
      13'h1508: dout <= 8'b00000000; // 5384 :   0 - 0x0
      13'h1509: dout <= 8'b00000000; // 5385 :   0 - 0x0
      13'h150A: dout <= 8'b00000000; // 5386 :   0 - 0x0
      13'h150B: dout <= 8'b00000000; // 5387 :   0 - 0x0
      13'h150C: dout <= 8'b00000000; // 5388 :   0 - 0x0
      13'h150D: dout <= 8'b00000000; // 5389 :   0 - 0x0
      13'h150E: dout <= 8'b00000000; // 5390 :   0 - 0x0
      13'h150F: dout <= 8'b00000000; // 5391 :   0 - 0x0
      13'h1510: dout <= 8'b00010000; // 5392 :  16 - 0x10 -- Background 0x51
      13'h1511: dout <= 8'b00101000; // 5393 :  40 - 0x28
      13'h1512: dout <= 8'b11101110; // 5394 : 238 - 0xee
      13'h1513: dout <= 8'b10000010; // 5395 : 130 - 0x82
      13'h1514: dout <= 8'b01000100; // 5396 :  68 - 0x44
      13'h1515: dout <= 8'b01000100; // 5397 :  68 - 0x44
      13'h1516: dout <= 8'b10010010; // 5398 : 146 - 0x92
      13'h1517: dout <= 8'b11101110; // 5399 : 238 - 0xee
      13'h1518: dout <= 8'b00000000; // 5400 :   0 - 0x0
      13'h1519: dout <= 8'b00010000; // 5401 :  16 - 0x10
      13'h151A: dout <= 8'b00010000; // 5402 :  16 - 0x10
      13'h151B: dout <= 8'b01111100; // 5403 : 124 - 0x7c
      13'h151C: dout <= 8'b00111000; // 5404 :  56 - 0x38
      13'h151D: dout <= 8'b00111000; // 5405 :  56 - 0x38
      13'h151E: dout <= 8'b01101100; // 5406 : 108 - 0x6c
      13'h151F: dout <= 8'b00000000; // 5407 :   0 - 0x0
      13'h1520: dout <= 8'b00010000; // 5408 :  16 - 0x10 -- Background 0x52
      13'h1521: dout <= 8'b00111000; // 5409 :  56 - 0x38
      13'h1522: dout <= 8'b11111110; // 5410 : 254 - 0xfe
      13'h1523: dout <= 8'b11111110; // 5411 : 254 - 0xfe
      13'h1524: dout <= 8'b01111100; // 5412 : 124 - 0x7c
      13'h1525: dout <= 8'b01111100; // 5413 : 124 - 0x7c
      13'h1526: dout <= 8'b11111110; // 5414 : 254 - 0xfe
      13'h1527: dout <= 8'b11101110; // 5415 : 238 - 0xee
      13'h1528: dout <= 8'b00000000; // 5416 :   0 - 0x0
      13'h1529: dout <= 8'b00010000; // 5417 :  16 - 0x10
      13'h152A: dout <= 8'b00010000; // 5418 :  16 - 0x10
      13'h152B: dout <= 8'b01111100; // 5419 : 124 - 0x7c
      13'h152C: dout <= 8'b00111000; // 5420 :  56 - 0x38
      13'h152D: dout <= 8'b00111000; // 5421 :  56 - 0x38
      13'h152E: dout <= 8'b01101100; // 5422 : 108 - 0x6c
      13'h152F: dout <= 8'b00000000; // 5423 :   0 - 0x0
      13'h1530: dout <= 8'b11111111; // 5424 : 255 - 0xff -- Background 0x53
      13'h1531: dout <= 8'b11111111; // 5425 : 255 - 0xff
      13'h1532: dout <= 8'b11111111; // 5426 : 255 - 0xff
      13'h1533: dout <= 8'b11111111; // 5427 : 255 - 0xff
      13'h1534: dout <= 8'b11111111; // 5428 : 255 - 0xff
      13'h1535: dout <= 8'b11111111; // 5429 : 255 - 0xff
      13'h1536: dout <= 8'b11111111; // 5430 : 255 - 0xff
      13'h1537: dout <= 8'b11111111; // 5431 : 255 - 0xff
      13'h1538: dout <= 8'b00000000; // 5432 :   0 - 0x0
      13'h1539: dout <= 8'b00000000; // 5433 :   0 - 0x0
      13'h153A: dout <= 8'b00000000; // 5434 :   0 - 0x0
      13'h153B: dout <= 8'b00000000; // 5435 :   0 - 0x0
      13'h153C: dout <= 8'b00000000; // 5436 :   0 - 0x0
      13'h153D: dout <= 8'b00000000; // 5437 :   0 - 0x0
      13'h153E: dout <= 8'b00000000; // 5438 :   0 - 0x0
      13'h153F: dout <= 8'b00000000; // 5439 :   0 - 0x0
      13'h1540: dout <= 8'b00000000; // 5440 :   0 - 0x0 -- Background 0x54
      13'h1541: dout <= 8'b00000000; // 5441 :   0 - 0x0
      13'h1542: dout <= 8'b00000000; // 5442 :   0 - 0x0
      13'h1543: dout <= 8'b00000000; // 5443 :   0 - 0x0
      13'h1544: dout <= 8'b00000000; // 5444 :   0 - 0x0
      13'h1545: dout <= 8'b00000000; // 5445 :   0 - 0x0
      13'h1546: dout <= 8'b00000000; // 5446 :   0 - 0x0
      13'h1547: dout <= 8'b00000000; // 5447 :   0 - 0x0
      13'h1548: dout <= 8'b11111111; // 5448 : 255 - 0xff
      13'h1549: dout <= 8'b11111111; // 5449 : 255 - 0xff
      13'h154A: dout <= 8'b11111111; // 5450 : 255 - 0xff
      13'h154B: dout <= 8'b11111111; // 5451 : 255 - 0xff
      13'h154C: dout <= 8'b11111111; // 5452 : 255 - 0xff
      13'h154D: dout <= 8'b11111111; // 5453 : 255 - 0xff
      13'h154E: dout <= 8'b11111111; // 5454 : 255 - 0xff
      13'h154F: dout <= 8'b11111111; // 5455 : 255 - 0xff
      13'h1550: dout <= 8'b11111111; // 5456 : 255 - 0xff -- Background 0x55
      13'h1551: dout <= 8'b11111111; // 5457 : 255 - 0xff
      13'h1552: dout <= 8'b11111111; // 5458 : 255 - 0xff
      13'h1553: dout <= 8'b11111111; // 5459 : 255 - 0xff
      13'h1554: dout <= 8'b11111111; // 5460 : 255 - 0xff
      13'h1555: dout <= 8'b11111111; // 5461 : 255 - 0xff
      13'h1556: dout <= 8'b11111111; // 5462 : 255 - 0xff
      13'h1557: dout <= 8'b11111111; // 5463 : 255 - 0xff
      13'h1558: dout <= 8'b11111111; // 5464 : 255 - 0xff
      13'h1559: dout <= 8'b11111111; // 5465 : 255 - 0xff
      13'h155A: dout <= 8'b11111111; // 5466 : 255 - 0xff
      13'h155B: dout <= 8'b11111111; // 5467 : 255 - 0xff
      13'h155C: dout <= 8'b11111111; // 5468 : 255 - 0xff
      13'h155D: dout <= 8'b11111111; // 5469 : 255 - 0xff
      13'h155E: dout <= 8'b11111111; // 5470 : 255 - 0xff
      13'h155F: dout <= 8'b11111111; // 5471 : 255 - 0xff
      13'h1560: dout <= 8'b00101010; // 5472 :  42 - 0x2a -- Background 0x56
      13'h1561: dout <= 8'b01000101; // 5473 :  69 - 0x45
      13'h1562: dout <= 8'b00001000; // 5474 :   8 - 0x8
      13'h1563: dout <= 8'b00010101; // 5475 :  21 - 0x15
      13'h1564: dout <= 8'b00100000; // 5476 :  32 - 0x20
      13'h1565: dout <= 8'b01000101; // 5477 :  69 - 0x45
      13'h1566: dout <= 8'b10101000; // 5478 : 168 - 0xa8
      13'h1567: dout <= 8'b00000000; // 5479 :   0 - 0x0
      13'h1568: dout <= 8'b00000010; // 5480 :   2 - 0x2
      13'h1569: dout <= 8'b00000101; // 5481 :   5 - 0x5
      13'h156A: dout <= 8'b10101010; // 5482 : 170 - 0xaa
      13'h156B: dout <= 8'b01010001; // 5483 :  81 - 0x51
      13'h156C: dout <= 8'b10101010; // 5484 : 170 - 0xaa
      13'h156D: dout <= 8'b01010001; // 5485 :  81 - 0x51
      13'h156E: dout <= 8'b10100010; // 5486 : 162 - 0xa2
      13'h156F: dout <= 8'b00000100; // 5487 :   4 - 0x4
      13'h1570: dout <= 8'b00001000; // 5488 :   8 - 0x8 -- Background 0x57
      13'h1571: dout <= 8'b01010101; // 5489 :  85 - 0x55
      13'h1572: dout <= 8'b10100000; // 5490 : 160 - 0xa0
      13'h1573: dout <= 8'b00010000; // 5491 :  16 - 0x10
      13'h1574: dout <= 8'b10000000; // 5492 : 128 - 0x80
      13'h1575: dout <= 8'b00010100; // 5493 :  20 - 0x14
      13'h1576: dout <= 8'b00100010; // 5494 :  34 - 0x22
      13'h1577: dout <= 8'b00000000; // 5495 :   0 - 0x0
      13'h1578: dout <= 8'b00001000; // 5496 :   8 - 0x8
      13'h1579: dout <= 8'b01010101; // 5497 :  85 - 0x55
      13'h157A: dout <= 8'b00101010; // 5498 :  42 - 0x2a
      13'h157B: dout <= 8'b01010101; // 5499 :  85 - 0x55
      13'h157C: dout <= 8'b00101010; // 5500 :  42 - 0x2a
      13'h157D: dout <= 8'b01000101; // 5501 :  69 - 0x45
      13'h157E: dout <= 8'b00001010; // 5502 :  10 - 0xa
      13'h157F: dout <= 8'b00010000; // 5503 :  16 - 0x10
      13'h1580: dout <= 8'b11111111; // 5504 : 255 - 0xff -- Background 0x58
      13'h1581: dout <= 8'b11010101; // 5505 : 213 - 0xd5
      13'h1582: dout <= 8'b10100000; // 5506 : 160 - 0xa0
      13'h1583: dout <= 8'b11010000; // 5507 : 208 - 0xd0
      13'h1584: dout <= 8'b10001111; // 5508 : 143 - 0x8f
      13'h1585: dout <= 8'b11001000; // 5509 : 200 - 0xc8
      13'h1586: dout <= 8'b10001000; // 5510 : 136 - 0x88
      13'h1587: dout <= 8'b11001000; // 5511 : 200 - 0xc8
      13'h1588: dout <= 8'b00000000; // 5512 :   0 - 0x0
      13'h1589: dout <= 8'b00111111; // 5513 :  63 - 0x3f
      13'h158A: dout <= 8'b01011111; // 5514 :  95 - 0x5f
      13'h158B: dout <= 8'b01101111; // 5515 : 111 - 0x6f
      13'h158C: dout <= 8'b01110000; // 5516 : 112 - 0x70
      13'h158D: dout <= 8'b01110111; // 5517 : 119 - 0x77
      13'h158E: dout <= 8'b01110111; // 5518 : 119 - 0x77
      13'h158F: dout <= 8'b01110111; // 5519 : 119 - 0x77
      13'h1590: dout <= 8'b10001000; // 5520 : 136 - 0x88 -- Background 0x59
      13'h1591: dout <= 8'b11001000; // 5521 : 200 - 0xc8
      13'h1592: dout <= 8'b10001000; // 5522 : 136 - 0x88
      13'h1593: dout <= 8'b11001111; // 5523 : 207 - 0xcf
      13'h1594: dout <= 8'b10010000; // 5524 : 144 - 0x90
      13'h1595: dout <= 8'b11100000; // 5525 : 224 - 0xe0
      13'h1596: dout <= 8'b11101010; // 5526 : 234 - 0xea
      13'h1597: dout <= 8'b11111111; // 5527 : 255 - 0xff
      13'h1598: dout <= 8'b01110111; // 5528 : 119 - 0x77
      13'h1599: dout <= 8'b01110111; // 5529 : 119 - 0x77
      13'h159A: dout <= 8'b01110111; // 5530 : 119 - 0x77
      13'h159B: dout <= 8'b01110000; // 5531 : 112 - 0x70
      13'h159C: dout <= 8'b01101111; // 5532 : 111 - 0x6f
      13'h159D: dout <= 8'b01011111; // 5533 :  95 - 0x5f
      13'h159E: dout <= 8'b00010101; // 5534 :  21 - 0x15
      13'h159F: dout <= 8'b00000000; // 5535 :   0 - 0x0
      13'h15A0: dout <= 8'b11111111; // 5536 : 255 - 0xff -- Background 0x5a
      13'h15A1: dout <= 8'b01011011; // 5537 :  91 - 0x5b
      13'h15A2: dout <= 8'b00000111; // 5538 :   7 - 0x7
      13'h15A3: dout <= 8'b00001001; // 5539 :   9 - 0x9
      13'h15A4: dout <= 8'b11110011; // 5540 : 243 - 0xf3
      13'h15A5: dout <= 8'b00010001; // 5541 :  17 - 0x11
      13'h15A6: dout <= 8'b00010011; // 5542 :  19 - 0x13
      13'h15A7: dout <= 8'b00010001; // 5543 :  17 - 0x11
      13'h15A8: dout <= 8'b00000000; // 5544 :   0 - 0x0
      13'h15A9: dout <= 8'b11111100; // 5545 : 252 - 0xfc
      13'h15AA: dout <= 8'b11111000; // 5546 : 248 - 0xf8
      13'h15AB: dout <= 8'b11110110; // 5547 : 246 - 0xf6
      13'h15AC: dout <= 8'b00001100; // 5548 :  12 - 0xc
      13'h15AD: dout <= 8'b11101110; // 5549 : 238 - 0xee
      13'h15AE: dout <= 8'b11101100; // 5550 : 236 - 0xec
      13'h15AF: dout <= 8'b11101110; // 5551 : 238 - 0xee
      13'h15B0: dout <= 8'b00010011; // 5552 :  19 - 0x13 -- Background 0x5b
      13'h15B1: dout <= 8'b00010001; // 5553 :  17 - 0x11
      13'h15B2: dout <= 8'b00010011; // 5554 :  19 - 0x13
      13'h15B3: dout <= 8'b11110001; // 5555 : 241 - 0xf1
      13'h15B4: dout <= 8'b00001011; // 5556 :  11 - 0xb
      13'h15B5: dout <= 8'b00000101; // 5557 :   5 - 0x5
      13'h15B6: dout <= 8'b10101011; // 5558 : 171 - 0xab
      13'h15B7: dout <= 8'b11111111; // 5559 : 255 - 0xff
      13'h15B8: dout <= 8'b11101100; // 5560 : 236 - 0xec
      13'h15B9: dout <= 8'b11101110; // 5561 : 238 - 0xee
      13'h15BA: dout <= 8'b11101100; // 5562 : 236 - 0xec
      13'h15BB: dout <= 8'b00001110; // 5563 :  14 - 0xe
      13'h15BC: dout <= 8'b11110100; // 5564 : 244 - 0xf4
      13'h15BD: dout <= 8'b11111010; // 5565 : 250 - 0xfa
      13'h15BE: dout <= 8'b01010100; // 5566 :  84 - 0x54
      13'h15BF: dout <= 8'b00000000; // 5567 :   0 - 0x0
      13'h15C0: dout <= 8'b00011100; // 5568 :  28 - 0x1c -- Background 0x5c
      13'h15C1: dout <= 8'b00100010; // 5569 :  34 - 0x22
      13'h15C2: dout <= 8'b01000001; // 5570 :  65 - 0x41
      13'h15C3: dout <= 8'b01000001; // 5571 :  65 - 0x41
      13'h15C4: dout <= 8'b01000001; // 5572 :  65 - 0x41
      13'h15C5: dout <= 8'b00100010; // 5573 :  34 - 0x22
      13'h15C6: dout <= 8'b00100010; // 5574 :  34 - 0x22
      13'h15C7: dout <= 8'b00011100; // 5575 :  28 - 0x1c
      13'h15C8: dout <= 8'b00000000; // 5576 :   0 - 0x0
      13'h15C9: dout <= 8'b00011100; // 5577 :  28 - 0x1c
      13'h15CA: dout <= 8'b00111110; // 5578 :  62 - 0x3e
      13'h15CB: dout <= 8'b00111110; // 5579 :  62 - 0x3e
      13'h15CC: dout <= 8'b00111110; // 5580 :  62 - 0x3e
      13'h15CD: dout <= 8'b00011100; // 5581 :  28 - 0x1c
      13'h15CE: dout <= 8'b00011100; // 5582 :  28 - 0x1c
      13'h15CF: dout <= 8'b00000000; // 5583 :   0 - 0x0
      13'h15D0: dout <= 8'b00001000; // 5584 :   8 - 0x8 -- Background 0x5d
      13'h15D1: dout <= 8'b00010000; // 5585 :  16 - 0x10
      13'h15D2: dout <= 8'b00010000; // 5586 :  16 - 0x10
      13'h15D3: dout <= 8'b00001000; // 5587 :   8 - 0x8
      13'h15D4: dout <= 8'b00000100; // 5588 :   4 - 0x4
      13'h15D5: dout <= 8'b00000100; // 5589 :   4 - 0x4
      13'h15D6: dout <= 8'b00001000; // 5590 :   8 - 0x8
      13'h15D7: dout <= 8'b00010000; // 5591 :  16 - 0x10
      13'h15D8: dout <= 8'b00000000; // 5592 :   0 - 0x0
      13'h15D9: dout <= 8'b00000000; // 5593 :   0 - 0x0
      13'h15DA: dout <= 8'b00000000; // 5594 :   0 - 0x0
      13'h15DB: dout <= 8'b00000000; // 5595 :   0 - 0x0
      13'h15DC: dout <= 8'b00000000; // 5596 :   0 - 0x0
      13'h15DD: dout <= 8'b00000000; // 5597 :   0 - 0x0
      13'h15DE: dout <= 8'b00000000; // 5598 :   0 - 0x0
      13'h15DF: dout <= 8'b00000000; // 5599 :   0 - 0x0
      13'h15E0: dout <= 8'b00110110; // 5600 :  54 - 0x36 -- Background 0x5e
      13'h15E1: dout <= 8'b01101011; // 5601 : 107 - 0x6b
      13'h15E2: dout <= 8'b01001001; // 5602 :  73 - 0x49
      13'h15E3: dout <= 8'b01000001; // 5603 :  65 - 0x41
      13'h15E4: dout <= 8'b01000001; // 5604 :  65 - 0x41
      13'h15E5: dout <= 8'b00100010; // 5605 :  34 - 0x22
      13'h15E6: dout <= 8'b00010100; // 5606 :  20 - 0x14
      13'h15E7: dout <= 8'b00001000; // 5607 :   8 - 0x8
      13'h15E8: dout <= 8'b00000000; // 5608 :   0 - 0x0
      13'h15E9: dout <= 8'b00010100; // 5609 :  20 - 0x14
      13'h15EA: dout <= 8'b00110110; // 5610 :  54 - 0x36
      13'h15EB: dout <= 8'b00111110; // 5611 :  62 - 0x3e
      13'h15EC: dout <= 8'b00111110; // 5612 :  62 - 0x3e
      13'h15ED: dout <= 8'b00011100; // 5613 :  28 - 0x1c
      13'h15EE: dout <= 8'b00001000; // 5614 :   8 - 0x8
      13'h15EF: dout <= 8'b00000000; // 5615 :   0 - 0x0
      13'h15F0: dout <= 8'b00111110; // 5616 :  62 - 0x3e -- Background 0x5f
      13'h15F1: dout <= 8'b01101011; // 5617 : 107 - 0x6b
      13'h15F2: dout <= 8'b00100010; // 5618 :  34 - 0x22
      13'h15F3: dout <= 8'b01100011; // 5619 :  99 - 0x63
      13'h15F4: dout <= 8'b00100010; // 5620 :  34 - 0x22
      13'h15F5: dout <= 8'b01100011; // 5621 :  99 - 0x63
      13'h15F6: dout <= 8'b00100010; // 5622 :  34 - 0x22
      13'h15F7: dout <= 8'b01111111; // 5623 : 127 - 0x7f
      13'h15F8: dout <= 8'b00000000; // 5624 :   0 - 0x0
      13'h15F9: dout <= 8'b00010100; // 5625 :  20 - 0x14
      13'h15FA: dout <= 8'b00011100; // 5626 :  28 - 0x1c
      13'h15FB: dout <= 8'b00011100; // 5627 :  28 - 0x1c
      13'h15FC: dout <= 8'b00011100; // 5628 :  28 - 0x1c
      13'h15FD: dout <= 8'b00011100; // 5629 :  28 - 0x1c
      13'h15FE: dout <= 8'b00011100; // 5630 :  28 - 0x1c
      13'h15FF: dout <= 8'b00000000; // 5631 :   0 - 0x0
      13'h1600: dout <= 8'b11111111; // 5632 : 255 - 0xff -- Background 0x60
      13'h1601: dout <= 8'b11111111; // 5633 : 255 - 0xff
      13'h1602: dout <= 8'b11111111; // 5634 : 255 - 0xff
      13'h1603: dout <= 8'b11111111; // 5635 : 255 - 0xff
      13'h1604: dout <= 8'b11010101; // 5636 : 213 - 0xd5
      13'h1605: dout <= 8'b10101010; // 5637 : 170 - 0xaa
      13'h1606: dout <= 8'b11010101; // 5638 : 213 - 0xd5
      13'h1607: dout <= 8'b11111111; // 5639 : 255 - 0xff
      13'h1608: dout <= 8'b00000000; // 5640 :   0 - 0x0
      13'h1609: dout <= 8'b01111111; // 5641 : 127 - 0x7f
      13'h160A: dout <= 8'b01111111; // 5642 : 127 - 0x7f
      13'h160B: dout <= 8'b01111111; // 5643 : 127 - 0x7f
      13'h160C: dout <= 8'b01111111; // 5644 : 127 - 0x7f
      13'h160D: dout <= 8'b01111111; // 5645 : 127 - 0x7f
      13'h160E: dout <= 8'b00101010; // 5646 :  42 - 0x2a
      13'h160F: dout <= 8'b00000000; // 5647 :   0 - 0x0
      13'h1610: dout <= 8'b11111111; // 5648 : 255 - 0xff -- Background 0x61
      13'h1611: dout <= 8'b11111111; // 5649 : 255 - 0xff
      13'h1612: dout <= 8'b11111111; // 5650 : 255 - 0xff
      13'h1613: dout <= 8'b11111111; // 5651 : 255 - 0xff
      13'h1614: dout <= 8'b01010101; // 5652 :  85 - 0x55
      13'h1615: dout <= 8'b10101010; // 5653 : 170 - 0xaa
      13'h1616: dout <= 8'b01010101; // 5654 :  85 - 0x55
      13'h1617: dout <= 8'b11111111; // 5655 : 255 - 0xff
      13'h1618: dout <= 8'b00000000; // 5656 :   0 - 0x0
      13'h1619: dout <= 8'b11111111; // 5657 : 255 - 0xff
      13'h161A: dout <= 8'b11111111; // 5658 : 255 - 0xff
      13'h161B: dout <= 8'b11111111; // 5659 : 255 - 0xff
      13'h161C: dout <= 8'b11111111; // 5660 : 255 - 0xff
      13'h161D: dout <= 8'b11111111; // 5661 : 255 - 0xff
      13'h161E: dout <= 8'b10101010; // 5662 : 170 - 0xaa
      13'h161F: dout <= 8'b00000000; // 5663 :   0 - 0x0
      13'h1620: dout <= 8'b11111111; // 5664 : 255 - 0xff -- Background 0x62
      13'h1621: dout <= 8'b11111111; // 5665 : 255 - 0xff
      13'h1622: dout <= 8'b11111111; // 5666 : 255 - 0xff
      13'h1623: dout <= 8'b11111111; // 5667 : 255 - 0xff
      13'h1624: dout <= 8'b01010101; // 5668 :  85 - 0x55
      13'h1625: dout <= 8'b10101011; // 5669 : 171 - 0xab
      13'h1626: dout <= 8'b01010101; // 5670 :  85 - 0x55
      13'h1627: dout <= 8'b11111111; // 5671 : 255 - 0xff
      13'h1628: dout <= 8'b00000000; // 5672 :   0 - 0x0
      13'h1629: dout <= 8'b11111110; // 5673 : 254 - 0xfe
      13'h162A: dout <= 8'b11111110; // 5674 : 254 - 0xfe
      13'h162B: dout <= 8'b11111110; // 5675 : 254 - 0xfe
      13'h162C: dout <= 8'b11111110; // 5676 : 254 - 0xfe
      13'h162D: dout <= 8'b11111110; // 5677 : 254 - 0xfe
      13'h162E: dout <= 8'b10101010; // 5678 : 170 - 0xaa
      13'h162F: dout <= 8'b00000000; // 5679 :   0 - 0x0
      13'h1630: dout <= 8'b00000000; // 5680 :   0 - 0x0 -- Background 0x63
      13'h1631: dout <= 8'b00000000; // 5681 :   0 - 0x0
      13'h1632: dout <= 8'b00000000; // 5682 :   0 - 0x0
      13'h1633: dout <= 8'b00000000; // 5683 :   0 - 0x0
      13'h1634: dout <= 8'b00000000; // 5684 :   0 - 0x0
      13'h1635: dout <= 8'b00000000; // 5685 :   0 - 0x0
      13'h1636: dout <= 8'b00000000; // 5686 :   0 - 0x0
      13'h1637: dout <= 8'b00000000; // 5687 :   0 - 0x0
      13'h1638: dout <= 8'b00000000; // 5688 :   0 - 0x0
      13'h1639: dout <= 8'b00000000; // 5689 :   0 - 0x0
      13'h163A: dout <= 8'b00000000; // 5690 :   0 - 0x0
      13'h163B: dout <= 8'b00000000; // 5691 :   0 - 0x0
      13'h163C: dout <= 8'b00000000; // 5692 :   0 - 0x0
      13'h163D: dout <= 8'b00000000; // 5693 :   0 - 0x0
      13'h163E: dout <= 8'b00000000; // 5694 :   0 - 0x0
      13'h163F: dout <= 8'b00000000; // 5695 :   0 - 0x0
      13'h1640: dout <= 8'b00000001; // 5696 :   1 - 0x1 -- Background 0x64
      13'h1641: dout <= 8'b00000001; // 5697 :   1 - 0x1
      13'h1642: dout <= 8'b00000011; // 5698 :   3 - 0x3
      13'h1643: dout <= 8'b00000011; // 5699 :   3 - 0x3
      13'h1644: dout <= 8'b00000110; // 5700 :   6 - 0x6
      13'h1645: dout <= 8'b00000110; // 5701 :   6 - 0x6
      13'h1646: dout <= 8'b00001100; // 5702 :  12 - 0xc
      13'h1647: dout <= 8'b00001100; // 5703 :  12 - 0xc
      13'h1648: dout <= 8'b00000000; // 5704 :   0 - 0x0
      13'h1649: dout <= 8'b00000000; // 5705 :   0 - 0x0
      13'h164A: dout <= 8'b00000001; // 5706 :   1 - 0x1
      13'h164B: dout <= 8'b00000001; // 5707 :   1 - 0x1
      13'h164C: dout <= 8'b00000011; // 5708 :   3 - 0x3
      13'h164D: dout <= 8'b00000011; // 5709 :   3 - 0x3
      13'h164E: dout <= 8'b00000111; // 5710 :   7 - 0x7
      13'h164F: dout <= 8'b00000111; // 5711 :   7 - 0x7
      13'h1650: dout <= 8'b00011000; // 5712 :  24 - 0x18 -- Background 0x65
      13'h1651: dout <= 8'b00011000; // 5713 :  24 - 0x18
      13'h1652: dout <= 8'b00110000; // 5714 :  48 - 0x30
      13'h1653: dout <= 8'b00110000; // 5715 :  48 - 0x30
      13'h1654: dout <= 8'b01100000; // 5716 :  96 - 0x60
      13'h1655: dout <= 8'b01100000; // 5717 :  96 - 0x60
      13'h1656: dout <= 8'b11101010; // 5718 : 234 - 0xea
      13'h1657: dout <= 8'b11111111; // 5719 : 255 - 0xff
      13'h1658: dout <= 8'b00001111; // 5720 :  15 - 0xf
      13'h1659: dout <= 8'b00001111; // 5721 :  15 - 0xf
      13'h165A: dout <= 8'b00011111; // 5722 :  31 - 0x1f
      13'h165B: dout <= 8'b00011111; // 5723 :  31 - 0x1f
      13'h165C: dout <= 8'b00111111; // 5724 :  63 - 0x3f
      13'h165D: dout <= 8'b00111111; // 5725 :  63 - 0x3f
      13'h165E: dout <= 8'b01010101; // 5726 :  85 - 0x55
      13'h165F: dout <= 8'b00000000; // 5727 :   0 - 0x0
      13'h1660: dout <= 8'b10000000; // 5728 : 128 - 0x80 -- Background 0x66
      13'h1661: dout <= 8'b10000000; // 5729 : 128 - 0x80
      13'h1662: dout <= 8'b11000000; // 5730 : 192 - 0xc0
      13'h1663: dout <= 8'b01000000; // 5731 :  64 - 0x40
      13'h1664: dout <= 8'b10100000; // 5732 : 160 - 0xa0
      13'h1665: dout <= 8'b01100000; // 5733 :  96 - 0x60
      13'h1666: dout <= 8'b00110000; // 5734 :  48 - 0x30
      13'h1667: dout <= 8'b00010000; // 5735 :  16 - 0x10
      13'h1668: dout <= 8'b00000000; // 5736 :   0 - 0x0
      13'h1669: dout <= 8'b00000000; // 5737 :   0 - 0x0
      13'h166A: dout <= 8'b00000000; // 5738 :   0 - 0x0
      13'h166B: dout <= 8'b10000000; // 5739 : 128 - 0x80
      13'h166C: dout <= 8'b01000000; // 5740 :  64 - 0x40
      13'h166D: dout <= 8'b10000000; // 5741 : 128 - 0x80
      13'h166E: dout <= 8'b11000000; // 5742 : 192 - 0xc0
      13'h166F: dout <= 8'b11100000; // 5743 : 224 - 0xe0
      13'h1670: dout <= 8'b00101000; // 5744 :  40 - 0x28 -- Background 0x67
      13'h1671: dout <= 8'b00011000; // 5745 :  24 - 0x18
      13'h1672: dout <= 8'b00001100; // 5746 :  12 - 0xc
      13'h1673: dout <= 8'b00010100; // 5747 :  20 - 0x14
      13'h1674: dout <= 8'b00001010; // 5748 :  10 - 0xa
      13'h1675: dout <= 8'b00000110; // 5749 :   6 - 0x6
      13'h1676: dout <= 8'b10101011; // 5750 : 171 - 0xab
      13'h1677: dout <= 8'b11111111; // 5751 : 255 - 0xff
      13'h1678: dout <= 8'b11010000; // 5752 : 208 - 0xd0
      13'h1679: dout <= 8'b11100000; // 5753 : 224 - 0xe0
      13'h167A: dout <= 8'b11110000; // 5754 : 240 - 0xf0
      13'h167B: dout <= 8'b11101000; // 5755 : 232 - 0xe8
      13'h167C: dout <= 8'b11110100; // 5756 : 244 - 0xf4
      13'h167D: dout <= 8'b11111000; // 5757 : 248 - 0xf8
      13'h167E: dout <= 8'b01010100; // 5758 :  84 - 0x54
      13'h167F: dout <= 8'b00000000; // 5759 :   0 - 0x0
      13'h1680: dout <= 8'b00000000; // 5760 :   0 - 0x0 -- Background 0x68
      13'h1681: dout <= 8'b00000000; // 5761 :   0 - 0x0
      13'h1682: dout <= 8'b00000000; // 5762 :   0 - 0x0
      13'h1683: dout <= 8'b00000000; // 5763 :   0 - 0x0
      13'h1684: dout <= 8'b00000000; // 5764 :   0 - 0x0
      13'h1685: dout <= 8'b00000000; // 5765 :   0 - 0x0
      13'h1686: dout <= 8'b00000000; // 5766 :   0 - 0x0
      13'h1687: dout <= 8'b00000000; // 5767 :   0 - 0x0
      13'h1688: dout <= 8'b00000000; // 5768 :   0 - 0x0
      13'h1689: dout <= 8'b00000000; // 5769 :   0 - 0x0
      13'h168A: dout <= 8'b00000000; // 5770 :   0 - 0x0
      13'h168B: dout <= 8'b00000000; // 5771 :   0 - 0x0
      13'h168C: dout <= 8'b00000000; // 5772 :   0 - 0x0
      13'h168D: dout <= 8'b00000000; // 5773 :   0 - 0x0
      13'h168E: dout <= 8'b00000000; // 5774 :   0 - 0x0
      13'h168F: dout <= 8'b00000000; // 5775 :   0 - 0x0
      13'h1690: dout <= 8'b00000000; // 5776 :   0 - 0x0 -- Background 0x69
      13'h1691: dout <= 8'b00000000; // 5777 :   0 - 0x0
      13'h1692: dout <= 8'b00000000; // 5778 :   0 - 0x0
      13'h1693: dout <= 8'b00000000; // 5779 :   0 - 0x0
      13'h1694: dout <= 8'b00000000; // 5780 :   0 - 0x0
      13'h1695: dout <= 8'b00000000; // 5781 :   0 - 0x0
      13'h1696: dout <= 8'b00000000; // 5782 :   0 - 0x0
      13'h1697: dout <= 8'b00000000; // 5783 :   0 - 0x0
      13'h1698: dout <= 8'b00000000; // 5784 :   0 - 0x0
      13'h1699: dout <= 8'b00000000; // 5785 :   0 - 0x0
      13'h169A: dout <= 8'b00000000; // 5786 :   0 - 0x0
      13'h169B: dout <= 8'b00000000; // 5787 :   0 - 0x0
      13'h169C: dout <= 8'b00000000; // 5788 :   0 - 0x0
      13'h169D: dout <= 8'b00000000; // 5789 :   0 - 0x0
      13'h169E: dout <= 8'b00000000; // 5790 :   0 - 0x0
      13'h169F: dout <= 8'b00000000; // 5791 :   0 - 0x0
      13'h16A0: dout <= 8'b00000000; // 5792 :   0 - 0x0 -- Background 0x6a
      13'h16A1: dout <= 8'b00000000; // 5793 :   0 - 0x0
      13'h16A2: dout <= 8'b00000000; // 5794 :   0 - 0x0
      13'h16A3: dout <= 8'b00000000; // 5795 :   0 - 0x0
      13'h16A4: dout <= 8'b00000000; // 5796 :   0 - 0x0
      13'h16A5: dout <= 8'b00000000; // 5797 :   0 - 0x0
      13'h16A6: dout <= 8'b00000000; // 5798 :   0 - 0x0
      13'h16A7: dout <= 8'b00000000; // 5799 :   0 - 0x0
      13'h16A8: dout <= 8'b00000000; // 5800 :   0 - 0x0
      13'h16A9: dout <= 8'b00000000; // 5801 :   0 - 0x0
      13'h16AA: dout <= 8'b00000000; // 5802 :   0 - 0x0
      13'h16AB: dout <= 8'b00000000; // 5803 :   0 - 0x0
      13'h16AC: dout <= 8'b00000000; // 5804 :   0 - 0x0
      13'h16AD: dout <= 8'b00000000; // 5805 :   0 - 0x0
      13'h16AE: dout <= 8'b00000000; // 5806 :   0 - 0x0
      13'h16AF: dout <= 8'b00000000; // 5807 :   0 - 0x0
      13'h16B0: dout <= 8'b00000000; // 5808 :   0 - 0x0 -- Background 0x6b
      13'h16B1: dout <= 8'b00000000; // 5809 :   0 - 0x0
      13'h16B2: dout <= 8'b00000000; // 5810 :   0 - 0x0
      13'h16B3: dout <= 8'b00000000; // 5811 :   0 - 0x0
      13'h16B4: dout <= 8'b00000000; // 5812 :   0 - 0x0
      13'h16B5: dout <= 8'b00000000; // 5813 :   0 - 0x0
      13'h16B6: dout <= 8'b00000000; // 5814 :   0 - 0x0
      13'h16B7: dout <= 8'b00000000; // 5815 :   0 - 0x0
      13'h16B8: dout <= 8'b00000000; // 5816 :   0 - 0x0
      13'h16B9: dout <= 8'b00000000; // 5817 :   0 - 0x0
      13'h16BA: dout <= 8'b00000000; // 5818 :   0 - 0x0
      13'h16BB: dout <= 8'b00000000; // 5819 :   0 - 0x0
      13'h16BC: dout <= 8'b00000000; // 5820 :   0 - 0x0
      13'h16BD: dout <= 8'b00000000; // 5821 :   0 - 0x0
      13'h16BE: dout <= 8'b00000000; // 5822 :   0 - 0x0
      13'h16BF: dout <= 8'b00000000; // 5823 :   0 - 0x0
      13'h16C0: dout <= 8'b00000000; // 5824 :   0 - 0x0 -- Background 0x6c
      13'h16C1: dout <= 8'b00000000; // 5825 :   0 - 0x0
      13'h16C2: dout <= 8'b00000000; // 5826 :   0 - 0x0
      13'h16C3: dout <= 8'b00000000; // 5827 :   0 - 0x0
      13'h16C4: dout <= 8'b00000000; // 5828 :   0 - 0x0
      13'h16C5: dout <= 8'b00000000; // 5829 :   0 - 0x0
      13'h16C6: dout <= 8'b00000000; // 5830 :   0 - 0x0
      13'h16C7: dout <= 8'b00000000; // 5831 :   0 - 0x0
      13'h16C8: dout <= 8'b00000000; // 5832 :   0 - 0x0
      13'h16C9: dout <= 8'b00000000; // 5833 :   0 - 0x0
      13'h16CA: dout <= 8'b00000000; // 5834 :   0 - 0x0
      13'h16CB: dout <= 8'b00000000; // 5835 :   0 - 0x0
      13'h16CC: dout <= 8'b00000000; // 5836 :   0 - 0x0
      13'h16CD: dout <= 8'b00000000; // 5837 :   0 - 0x0
      13'h16CE: dout <= 8'b00000000; // 5838 :   0 - 0x0
      13'h16CF: dout <= 8'b00000000; // 5839 :   0 - 0x0
      13'h16D0: dout <= 8'b00000000; // 5840 :   0 - 0x0 -- Background 0x6d
      13'h16D1: dout <= 8'b00000000; // 5841 :   0 - 0x0
      13'h16D2: dout <= 8'b00000000; // 5842 :   0 - 0x0
      13'h16D3: dout <= 8'b00000000; // 5843 :   0 - 0x0
      13'h16D4: dout <= 8'b00000000; // 5844 :   0 - 0x0
      13'h16D5: dout <= 8'b00000000; // 5845 :   0 - 0x0
      13'h16D6: dout <= 8'b00000000; // 5846 :   0 - 0x0
      13'h16D7: dout <= 8'b00000000; // 5847 :   0 - 0x0
      13'h16D8: dout <= 8'b00000000; // 5848 :   0 - 0x0
      13'h16D9: dout <= 8'b00000000; // 5849 :   0 - 0x0
      13'h16DA: dout <= 8'b00000000; // 5850 :   0 - 0x0
      13'h16DB: dout <= 8'b00000000; // 5851 :   0 - 0x0
      13'h16DC: dout <= 8'b00000000; // 5852 :   0 - 0x0
      13'h16DD: dout <= 8'b00000000; // 5853 :   0 - 0x0
      13'h16DE: dout <= 8'b00000000; // 5854 :   0 - 0x0
      13'h16DF: dout <= 8'b00000000; // 5855 :   0 - 0x0
      13'h16E0: dout <= 8'b00000000; // 5856 :   0 - 0x0 -- Background 0x6e
      13'h16E1: dout <= 8'b00000000; // 5857 :   0 - 0x0
      13'h16E2: dout <= 8'b00000000; // 5858 :   0 - 0x0
      13'h16E3: dout <= 8'b00000000; // 5859 :   0 - 0x0
      13'h16E4: dout <= 8'b00000000; // 5860 :   0 - 0x0
      13'h16E5: dout <= 8'b00000000; // 5861 :   0 - 0x0
      13'h16E6: dout <= 8'b00000000; // 5862 :   0 - 0x0
      13'h16E7: dout <= 8'b00000000; // 5863 :   0 - 0x0
      13'h16E8: dout <= 8'b00000000; // 5864 :   0 - 0x0
      13'h16E9: dout <= 8'b00000000; // 5865 :   0 - 0x0
      13'h16EA: dout <= 8'b00000000; // 5866 :   0 - 0x0
      13'h16EB: dout <= 8'b00000000; // 5867 :   0 - 0x0
      13'h16EC: dout <= 8'b00000000; // 5868 :   0 - 0x0
      13'h16ED: dout <= 8'b00000000; // 5869 :   0 - 0x0
      13'h16EE: dout <= 8'b00000000; // 5870 :   0 - 0x0
      13'h16EF: dout <= 8'b00000000; // 5871 :   0 - 0x0
      13'h16F0: dout <= 8'b00000000; // 5872 :   0 - 0x0 -- Background 0x6f
      13'h16F1: dout <= 8'b00000000; // 5873 :   0 - 0x0
      13'h16F2: dout <= 8'b00000000; // 5874 :   0 - 0x0
      13'h16F3: dout <= 8'b00000000; // 5875 :   0 - 0x0
      13'h16F4: dout <= 8'b00000000; // 5876 :   0 - 0x0
      13'h16F5: dout <= 8'b00000000; // 5877 :   0 - 0x0
      13'h16F6: dout <= 8'b00000000; // 5878 :   0 - 0x0
      13'h16F7: dout <= 8'b00000000; // 5879 :   0 - 0x0
      13'h16F8: dout <= 8'b00000000; // 5880 :   0 - 0x0
      13'h16F9: dout <= 8'b00000000; // 5881 :   0 - 0x0
      13'h16FA: dout <= 8'b00000000; // 5882 :   0 - 0x0
      13'h16FB: dout <= 8'b00000000; // 5883 :   0 - 0x0
      13'h16FC: dout <= 8'b00000000; // 5884 :   0 - 0x0
      13'h16FD: dout <= 8'b00000000; // 5885 :   0 - 0x0
      13'h16FE: dout <= 8'b00000000; // 5886 :   0 - 0x0
      13'h16FF: dout <= 8'b00000000; // 5887 :   0 - 0x0
      13'h1700: dout <= 8'b00000000; // 5888 :   0 - 0x0 -- Background 0x70
      13'h1701: dout <= 8'b00000000; // 5889 :   0 - 0x0
      13'h1702: dout <= 8'b00000000; // 5890 :   0 - 0x0
      13'h1703: dout <= 8'b00000000; // 5891 :   0 - 0x0
      13'h1704: dout <= 8'b00000000; // 5892 :   0 - 0x0
      13'h1705: dout <= 8'b00000000; // 5893 :   0 - 0x0
      13'h1706: dout <= 8'b00000000; // 5894 :   0 - 0x0
      13'h1707: dout <= 8'b00000000; // 5895 :   0 - 0x0
      13'h1708: dout <= 8'b00000000; // 5896 :   0 - 0x0
      13'h1709: dout <= 8'b00000000; // 5897 :   0 - 0x0
      13'h170A: dout <= 8'b00000000; // 5898 :   0 - 0x0
      13'h170B: dout <= 8'b00000000; // 5899 :   0 - 0x0
      13'h170C: dout <= 8'b00000000; // 5900 :   0 - 0x0
      13'h170D: dout <= 8'b00000000; // 5901 :   0 - 0x0
      13'h170E: dout <= 8'b00000000; // 5902 :   0 - 0x0
      13'h170F: dout <= 8'b00000000; // 5903 :   0 - 0x0
      13'h1710: dout <= 8'b00000000; // 5904 :   0 - 0x0 -- Background 0x71
      13'h1711: dout <= 8'b00000000; // 5905 :   0 - 0x0
      13'h1712: dout <= 8'b00000000; // 5906 :   0 - 0x0
      13'h1713: dout <= 8'b00000000; // 5907 :   0 - 0x0
      13'h1714: dout <= 8'b00000000; // 5908 :   0 - 0x0
      13'h1715: dout <= 8'b00000000; // 5909 :   0 - 0x0
      13'h1716: dout <= 8'b00000000; // 5910 :   0 - 0x0
      13'h1717: dout <= 8'b00000000; // 5911 :   0 - 0x0
      13'h1718: dout <= 8'b00000000; // 5912 :   0 - 0x0
      13'h1719: dout <= 8'b00000000; // 5913 :   0 - 0x0
      13'h171A: dout <= 8'b00000000; // 5914 :   0 - 0x0
      13'h171B: dout <= 8'b00000000; // 5915 :   0 - 0x0
      13'h171C: dout <= 8'b00000000; // 5916 :   0 - 0x0
      13'h171D: dout <= 8'b00000000; // 5917 :   0 - 0x0
      13'h171E: dout <= 8'b00000000; // 5918 :   0 - 0x0
      13'h171F: dout <= 8'b00000000; // 5919 :   0 - 0x0
      13'h1720: dout <= 8'b00000000; // 5920 :   0 - 0x0 -- Background 0x72
      13'h1721: dout <= 8'b00000000; // 5921 :   0 - 0x0
      13'h1722: dout <= 8'b00000000; // 5922 :   0 - 0x0
      13'h1723: dout <= 8'b00000000; // 5923 :   0 - 0x0
      13'h1724: dout <= 8'b00000000; // 5924 :   0 - 0x0
      13'h1725: dout <= 8'b00000000; // 5925 :   0 - 0x0
      13'h1726: dout <= 8'b00000000; // 5926 :   0 - 0x0
      13'h1727: dout <= 8'b00000000; // 5927 :   0 - 0x0
      13'h1728: dout <= 8'b00000000; // 5928 :   0 - 0x0
      13'h1729: dout <= 8'b00000000; // 5929 :   0 - 0x0
      13'h172A: dout <= 8'b00000000; // 5930 :   0 - 0x0
      13'h172B: dout <= 8'b00000000; // 5931 :   0 - 0x0
      13'h172C: dout <= 8'b00000000; // 5932 :   0 - 0x0
      13'h172D: dout <= 8'b00000000; // 5933 :   0 - 0x0
      13'h172E: dout <= 8'b00000000; // 5934 :   0 - 0x0
      13'h172F: dout <= 8'b00000000; // 5935 :   0 - 0x0
      13'h1730: dout <= 8'b00000000; // 5936 :   0 - 0x0 -- Background 0x73
      13'h1731: dout <= 8'b00000000; // 5937 :   0 - 0x0
      13'h1732: dout <= 8'b00000000; // 5938 :   0 - 0x0
      13'h1733: dout <= 8'b00000000; // 5939 :   0 - 0x0
      13'h1734: dout <= 8'b00000000; // 5940 :   0 - 0x0
      13'h1735: dout <= 8'b00000000; // 5941 :   0 - 0x0
      13'h1736: dout <= 8'b00000000; // 5942 :   0 - 0x0
      13'h1737: dout <= 8'b00000000; // 5943 :   0 - 0x0
      13'h1738: dout <= 8'b00000000; // 5944 :   0 - 0x0
      13'h1739: dout <= 8'b00000000; // 5945 :   0 - 0x0
      13'h173A: dout <= 8'b00000000; // 5946 :   0 - 0x0
      13'h173B: dout <= 8'b00000000; // 5947 :   0 - 0x0
      13'h173C: dout <= 8'b00000000; // 5948 :   0 - 0x0
      13'h173D: dout <= 8'b00000000; // 5949 :   0 - 0x0
      13'h173E: dout <= 8'b00000000; // 5950 :   0 - 0x0
      13'h173F: dout <= 8'b00000000; // 5951 :   0 - 0x0
      13'h1740: dout <= 8'b00000000; // 5952 :   0 - 0x0 -- Background 0x74
      13'h1741: dout <= 8'b00000000; // 5953 :   0 - 0x0
      13'h1742: dout <= 8'b00000000; // 5954 :   0 - 0x0
      13'h1743: dout <= 8'b00000000; // 5955 :   0 - 0x0
      13'h1744: dout <= 8'b00000000; // 5956 :   0 - 0x0
      13'h1745: dout <= 8'b00000000; // 5957 :   0 - 0x0
      13'h1746: dout <= 8'b00000000; // 5958 :   0 - 0x0
      13'h1747: dout <= 8'b00000000; // 5959 :   0 - 0x0
      13'h1748: dout <= 8'b00000000; // 5960 :   0 - 0x0
      13'h1749: dout <= 8'b00000000; // 5961 :   0 - 0x0
      13'h174A: dout <= 8'b00000000; // 5962 :   0 - 0x0
      13'h174B: dout <= 8'b00000000; // 5963 :   0 - 0x0
      13'h174C: dout <= 8'b00000000; // 5964 :   0 - 0x0
      13'h174D: dout <= 8'b00000000; // 5965 :   0 - 0x0
      13'h174E: dout <= 8'b00000000; // 5966 :   0 - 0x0
      13'h174F: dout <= 8'b00000000; // 5967 :   0 - 0x0
      13'h1750: dout <= 8'b00000000; // 5968 :   0 - 0x0 -- Background 0x75
      13'h1751: dout <= 8'b00000000; // 5969 :   0 - 0x0
      13'h1752: dout <= 8'b00000000; // 5970 :   0 - 0x0
      13'h1753: dout <= 8'b00000000; // 5971 :   0 - 0x0
      13'h1754: dout <= 8'b00000000; // 5972 :   0 - 0x0
      13'h1755: dout <= 8'b00000000; // 5973 :   0 - 0x0
      13'h1756: dout <= 8'b00000000; // 5974 :   0 - 0x0
      13'h1757: dout <= 8'b00000000; // 5975 :   0 - 0x0
      13'h1758: dout <= 8'b00000000; // 5976 :   0 - 0x0
      13'h1759: dout <= 8'b00000000; // 5977 :   0 - 0x0
      13'h175A: dout <= 8'b00000000; // 5978 :   0 - 0x0
      13'h175B: dout <= 8'b00000000; // 5979 :   0 - 0x0
      13'h175C: dout <= 8'b00000000; // 5980 :   0 - 0x0
      13'h175D: dout <= 8'b00000000; // 5981 :   0 - 0x0
      13'h175E: dout <= 8'b00000000; // 5982 :   0 - 0x0
      13'h175F: dout <= 8'b00000000; // 5983 :   0 - 0x0
      13'h1760: dout <= 8'b00000000; // 5984 :   0 - 0x0 -- Background 0x76
      13'h1761: dout <= 8'b00000000; // 5985 :   0 - 0x0
      13'h1762: dout <= 8'b00000000; // 5986 :   0 - 0x0
      13'h1763: dout <= 8'b00000000; // 5987 :   0 - 0x0
      13'h1764: dout <= 8'b00000000; // 5988 :   0 - 0x0
      13'h1765: dout <= 8'b00000000; // 5989 :   0 - 0x0
      13'h1766: dout <= 8'b00000000; // 5990 :   0 - 0x0
      13'h1767: dout <= 8'b00000000; // 5991 :   0 - 0x0
      13'h1768: dout <= 8'b00000000; // 5992 :   0 - 0x0
      13'h1769: dout <= 8'b00000000; // 5993 :   0 - 0x0
      13'h176A: dout <= 8'b00000000; // 5994 :   0 - 0x0
      13'h176B: dout <= 8'b00000000; // 5995 :   0 - 0x0
      13'h176C: dout <= 8'b00000000; // 5996 :   0 - 0x0
      13'h176D: dout <= 8'b00000000; // 5997 :   0 - 0x0
      13'h176E: dout <= 8'b00000000; // 5998 :   0 - 0x0
      13'h176F: dout <= 8'b00000000; // 5999 :   0 - 0x0
      13'h1770: dout <= 8'b00000000; // 6000 :   0 - 0x0 -- Background 0x77
      13'h1771: dout <= 8'b00000000; // 6001 :   0 - 0x0
      13'h1772: dout <= 8'b00000000; // 6002 :   0 - 0x0
      13'h1773: dout <= 8'b00000000; // 6003 :   0 - 0x0
      13'h1774: dout <= 8'b00000000; // 6004 :   0 - 0x0
      13'h1775: dout <= 8'b00000000; // 6005 :   0 - 0x0
      13'h1776: dout <= 8'b00000000; // 6006 :   0 - 0x0
      13'h1777: dout <= 8'b00000000; // 6007 :   0 - 0x0
      13'h1778: dout <= 8'b00000000; // 6008 :   0 - 0x0
      13'h1779: dout <= 8'b00000000; // 6009 :   0 - 0x0
      13'h177A: dout <= 8'b00000000; // 6010 :   0 - 0x0
      13'h177B: dout <= 8'b00000000; // 6011 :   0 - 0x0
      13'h177C: dout <= 8'b00000000; // 6012 :   0 - 0x0
      13'h177D: dout <= 8'b00000000; // 6013 :   0 - 0x0
      13'h177E: dout <= 8'b00000000; // 6014 :   0 - 0x0
      13'h177F: dout <= 8'b00000000; // 6015 :   0 - 0x0
      13'h1780: dout <= 8'b00000000; // 6016 :   0 - 0x0 -- Background 0x78
      13'h1781: dout <= 8'b00000000; // 6017 :   0 - 0x0
      13'h1782: dout <= 8'b00000000; // 6018 :   0 - 0x0
      13'h1783: dout <= 8'b00000000; // 6019 :   0 - 0x0
      13'h1784: dout <= 8'b00000000; // 6020 :   0 - 0x0
      13'h1785: dout <= 8'b00000000; // 6021 :   0 - 0x0
      13'h1786: dout <= 8'b00000000; // 6022 :   0 - 0x0
      13'h1787: dout <= 8'b00000000; // 6023 :   0 - 0x0
      13'h1788: dout <= 8'b00000000; // 6024 :   0 - 0x0
      13'h1789: dout <= 8'b00000000; // 6025 :   0 - 0x0
      13'h178A: dout <= 8'b00000000; // 6026 :   0 - 0x0
      13'h178B: dout <= 8'b00000000; // 6027 :   0 - 0x0
      13'h178C: dout <= 8'b00000000; // 6028 :   0 - 0x0
      13'h178D: dout <= 8'b00000000; // 6029 :   0 - 0x0
      13'h178E: dout <= 8'b00000000; // 6030 :   0 - 0x0
      13'h178F: dout <= 8'b00000000; // 6031 :   0 - 0x0
      13'h1790: dout <= 8'b00000000; // 6032 :   0 - 0x0 -- Background 0x79
      13'h1791: dout <= 8'b00000000; // 6033 :   0 - 0x0
      13'h1792: dout <= 8'b00000000; // 6034 :   0 - 0x0
      13'h1793: dout <= 8'b00000000; // 6035 :   0 - 0x0
      13'h1794: dout <= 8'b00000000; // 6036 :   0 - 0x0
      13'h1795: dout <= 8'b00000000; // 6037 :   0 - 0x0
      13'h1796: dout <= 8'b00000000; // 6038 :   0 - 0x0
      13'h1797: dout <= 8'b00000000; // 6039 :   0 - 0x0
      13'h1798: dout <= 8'b00000000; // 6040 :   0 - 0x0
      13'h1799: dout <= 8'b00000000; // 6041 :   0 - 0x0
      13'h179A: dout <= 8'b00000000; // 6042 :   0 - 0x0
      13'h179B: dout <= 8'b00000000; // 6043 :   0 - 0x0
      13'h179C: dout <= 8'b00000000; // 6044 :   0 - 0x0
      13'h179D: dout <= 8'b00000000; // 6045 :   0 - 0x0
      13'h179E: dout <= 8'b00000000; // 6046 :   0 - 0x0
      13'h179F: dout <= 8'b00000000; // 6047 :   0 - 0x0
      13'h17A0: dout <= 8'b00000000; // 6048 :   0 - 0x0 -- Background 0x7a
      13'h17A1: dout <= 8'b00000000; // 6049 :   0 - 0x0
      13'h17A2: dout <= 8'b00000000; // 6050 :   0 - 0x0
      13'h17A3: dout <= 8'b00000000; // 6051 :   0 - 0x0
      13'h17A4: dout <= 8'b00000000; // 6052 :   0 - 0x0
      13'h17A5: dout <= 8'b00000000; // 6053 :   0 - 0x0
      13'h17A6: dout <= 8'b00000000; // 6054 :   0 - 0x0
      13'h17A7: dout <= 8'b00000000; // 6055 :   0 - 0x0
      13'h17A8: dout <= 8'b00000000; // 6056 :   0 - 0x0
      13'h17A9: dout <= 8'b00000000; // 6057 :   0 - 0x0
      13'h17AA: dout <= 8'b00000000; // 6058 :   0 - 0x0
      13'h17AB: dout <= 8'b00000000; // 6059 :   0 - 0x0
      13'h17AC: dout <= 8'b00000000; // 6060 :   0 - 0x0
      13'h17AD: dout <= 8'b00000000; // 6061 :   0 - 0x0
      13'h17AE: dout <= 8'b00000000; // 6062 :   0 - 0x0
      13'h17AF: dout <= 8'b00000000; // 6063 :   0 - 0x0
      13'h17B0: dout <= 8'b00000000; // 6064 :   0 - 0x0 -- Background 0x7b
      13'h17B1: dout <= 8'b00000000; // 6065 :   0 - 0x0
      13'h17B2: dout <= 8'b00000000; // 6066 :   0 - 0x0
      13'h17B3: dout <= 8'b00000000; // 6067 :   0 - 0x0
      13'h17B4: dout <= 8'b00000000; // 6068 :   0 - 0x0
      13'h17B5: dout <= 8'b00000000; // 6069 :   0 - 0x0
      13'h17B6: dout <= 8'b00000000; // 6070 :   0 - 0x0
      13'h17B7: dout <= 8'b00000000; // 6071 :   0 - 0x0
      13'h17B8: dout <= 8'b00000000; // 6072 :   0 - 0x0
      13'h17B9: dout <= 8'b00000000; // 6073 :   0 - 0x0
      13'h17BA: dout <= 8'b00000000; // 6074 :   0 - 0x0
      13'h17BB: dout <= 8'b00000000; // 6075 :   0 - 0x0
      13'h17BC: dout <= 8'b00000000; // 6076 :   0 - 0x0
      13'h17BD: dout <= 8'b00000000; // 6077 :   0 - 0x0
      13'h17BE: dout <= 8'b00000000; // 6078 :   0 - 0x0
      13'h17BF: dout <= 8'b00000000; // 6079 :   0 - 0x0
      13'h17C0: dout <= 8'b00000000; // 6080 :   0 - 0x0 -- Background 0x7c
      13'h17C1: dout <= 8'b00000000; // 6081 :   0 - 0x0
      13'h17C2: dout <= 8'b00000000; // 6082 :   0 - 0x0
      13'h17C3: dout <= 8'b00000000; // 6083 :   0 - 0x0
      13'h17C4: dout <= 8'b00000000; // 6084 :   0 - 0x0
      13'h17C5: dout <= 8'b00000000; // 6085 :   0 - 0x0
      13'h17C6: dout <= 8'b00000000; // 6086 :   0 - 0x0
      13'h17C7: dout <= 8'b00000000; // 6087 :   0 - 0x0
      13'h17C8: dout <= 8'b00000000; // 6088 :   0 - 0x0
      13'h17C9: dout <= 8'b00000000; // 6089 :   0 - 0x0
      13'h17CA: dout <= 8'b00000000; // 6090 :   0 - 0x0
      13'h17CB: dout <= 8'b00000000; // 6091 :   0 - 0x0
      13'h17CC: dout <= 8'b00000000; // 6092 :   0 - 0x0
      13'h17CD: dout <= 8'b00000000; // 6093 :   0 - 0x0
      13'h17CE: dout <= 8'b00000000; // 6094 :   0 - 0x0
      13'h17CF: dout <= 8'b00000000; // 6095 :   0 - 0x0
      13'h17D0: dout <= 8'b00000000; // 6096 :   0 - 0x0 -- Background 0x7d
      13'h17D1: dout <= 8'b00000000; // 6097 :   0 - 0x0
      13'h17D2: dout <= 8'b00000000; // 6098 :   0 - 0x0
      13'h17D3: dout <= 8'b00000000; // 6099 :   0 - 0x0
      13'h17D4: dout <= 8'b00000000; // 6100 :   0 - 0x0
      13'h17D5: dout <= 8'b00000000; // 6101 :   0 - 0x0
      13'h17D6: dout <= 8'b00000000; // 6102 :   0 - 0x0
      13'h17D7: dout <= 8'b00000000; // 6103 :   0 - 0x0
      13'h17D8: dout <= 8'b00000000; // 6104 :   0 - 0x0
      13'h17D9: dout <= 8'b00000000; // 6105 :   0 - 0x0
      13'h17DA: dout <= 8'b00000000; // 6106 :   0 - 0x0
      13'h17DB: dout <= 8'b00000000; // 6107 :   0 - 0x0
      13'h17DC: dout <= 8'b00000000; // 6108 :   0 - 0x0
      13'h17DD: dout <= 8'b00000000; // 6109 :   0 - 0x0
      13'h17DE: dout <= 8'b00000000; // 6110 :   0 - 0x0
      13'h17DF: dout <= 8'b00000000; // 6111 :   0 - 0x0
      13'h17E0: dout <= 8'b00000000; // 6112 :   0 - 0x0 -- Background 0x7e
      13'h17E1: dout <= 8'b00000000; // 6113 :   0 - 0x0
      13'h17E2: dout <= 8'b00000000; // 6114 :   0 - 0x0
      13'h17E3: dout <= 8'b00000000; // 6115 :   0 - 0x0
      13'h17E4: dout <= 8'b00000000; // 6116 :   0 - 0x0
      13'h17E5: dout <= 8'b00000000; // 6117 :   0 - 0x0
      13'h17E6: dout <= 8'b00000000; // 6118 :   0 - 0x0
      13'h17E7: dout <= 8'b00000000; // 6119 :   0 - 0x0
      13'h17E8: dout <= 8'b00000000; // 6120 :   0 - 0x0
      13'h17E9: dout <= 8'b00000000; // 6121 :   0 - 0x0
      13'h17EA: dout <= 8'b00000000; // 6122 :   0 - 0x0
      13'h17EB: dout <= 8'b00000000; // 6123 :   0 - 0x0
      13'h17EC: dout <= 8'b00000000; // 6124 :   0 - 0x0
      13'h17ED: dout <= 8'b00000000; // 6125 :   0 - 0x0
      13'h17EE: dout <= 8'b00000000; // 6126 :   0 - 0x0
      13'h17EF: dout <= 8'b00000000; // 6127 :   0 - 0x0
      13'h17F0: dout <= 8'b00000000; // 6128 :   0 - 0x0 -- Background 0x7f
      13'h17F1: dout <= 8'b00000000; // 6129 :   0 - 0x0
      13'h17F2: dout <= 8'b00000000; // 6130 :   0 - 0x0
      13'h17F3: dout <= 8'b00000000; // 6131 :   0 - 0x0
      13'h17F4: dout <= 8'b00000000; // 6132 :   0 - 0x0
      13'h17F5: dout <= 8'b00000000; // 6133 :   0 - 0x0
      13'h17F6: dout <= 8'b00000000; // 6134 :   0 - 0x0
      13'h17F7: dout <= 8'b00000000; // 6135 :   0 - 0x0
      13'h17F8: dout <= 8'b00000000; // 6136 :   0 - 0x0
      13'h17F9: dout <= 8'b00000000; // 6137 :   0 - 0x0
      13'h17FA: dout <= 8'b00000000; // 6138 :   0 - 0x0
      13'h17FB: dout <= 8'b00000000; // 6139 :   0 - 0x0
      13'h17FC: dout <= 8'b00000000; // 6140 :   0 - 0x0
      13'h17FD: dout <= 8'b00000000; // 6141 :   0 - 0x0
      13'h17FE: dout <= 8'b00000000; // 6142 :   0 - 0x0
      13'h17FF: dout <= 8'b00000000; // 6143 :   0 - 0x0
      13'h1800: dout <= 8'b00000011; // 6144 :   3 - 0x3 -- Background 0x80
      13'h1801: dout <= 8'b00001111; // 6145 :  15 - 0xf
      13'h1802: dout <= 8'b00011100; // 6146 :  28 - 0x1c
      13'h1803: dout <= 8'b00110000; // 6147 :  48 - 0x30
      13'h1804: dout <= 8'b00100000; // 6148 :  32 - 0x20
      13'h1805: dout <= 8'b01000000; // 6149 :  64 - 0x40
      13'h1806: dout <= 8'b01000000; // 6150 :  64 - 0x40
      13'h1807: dout <= 8'b01111111; // 6151 : 127 - 0x7f
      13'h1808: dout <= 8'b00000000; // 6152 :   0 - 0x0
      13'h1809: dout <= 8'b00000011; // 6153 :   3 - 0x3
      13'h180A: dout <= 8'b00001111; // 6154 :  15 - 0xf
      13'h180B: dout <= 8'b00011111; // 6155 :  31 - 0x1f
      13'h180C: dout <= 8'b00011111; // 6156 :  31 - 0x1f
      13'h180D: dout <= 8'b00111111; // 6157 :  63 - 0x3f
      13'h180E: dout <= 8'b00111111; // 6158 :  63 - 0x3f
      13'h180F: dout <= 8'b00000000; // 6159 :   0 - 0x0
      13'h1810: dout <= 8'b00000001; // 6160 :   1 - 0x1 -- Background 0x81
      13'h1811: dout <= 8'b00000001; // 6161 :   1 - 0x1
      13'h1812: dout <= 8'b00000001; // 6162 :   1 - 0x1
      13'h1813: dout <= 8'b00000001; // 6163 :   1 - 0x1
      13'h1814: dout <= 8'b00000001; // 6164 :   1 - 0x1
      13'h1815: dout <= 8'b00000001; // 6165 :   1 - 0x1
      13'h1816: dout <= 8'b00000011; // 6166 :   3 - 0x3
      13'h1817: dout <= 8'b00000011; // 6167 :   3 - 0x3
      13'h1818: dout <= 8'b00000000; // 6168 :   0 - 0x0
      13'h1819: dout <= 8'b00000000; // 6169 :   0 - 0x0
      13'h181A: dout <= 8'b00000000; // 6170 :   0 - 0x0
      13'h181B: dout <= 8'b00000000; // 6171 :   0 - 0x0
      13'h181C: dout <= 8'b00000000; // 6172 :   0 - 0x0
      13'h181D: dout <= 8'b00000000; // 6173 :   0 - 0x0
      13'h181E: dout <= 8'b00000000; // 6174 :   0 - 0x0
      13'h181F: dout <= 8'b00000000; // 6175 :   0 - 0x0
      13'h1820: dout <= 8'b11000000; // 6176 : 192 - 0xc0 -- Background 0x82
      13'h1821: dout <= 8'b11110000; // 6177 : 240 - 0xf0
      13'h1822: dout <= 8'b00111000; // 6178 :  56 - 0x38
      13'h1823: dout <= 8'b00001110; // 6179 :  14 - 0xe
      13'h1824: dout <= 8'b00011110; // 6180 :  30 - 0x1e
      13'h1825: dout <= 8'b00011110; // 6181 :  30 - 0x1e
      13'h1826: dout <= 8'b00000010; // 6182 :   2 - 0x2
      13'h1827: dout <= 8'b11111110; // 6183 : 254 - 0xfe
      13'h1828: dout <= 8'b00000000; // 6184 :   0 - 0x0
      13'h1829: dout <= 8'b11000000; // 6185 : 192 - 0xc0
      13'h182A: dout <= 8'b11110000; // 6186 : 240 - 0xf0
      13'h182B: dout <= 8'b11110000; // 6187 : 240 - 0xf0
      13'h182C: dout <= 8'b11101100; // 6188 : 236 - 0xec
      13'h182D: dout <= 8'b11100000; // 6189 : 224 - 0xe0
      13'h182E: dout <= 8'b11111100; // 6190 : 252 - 0xfc
      13'h182F: dout <= 8'b00000000; // 6191 :   0 - 0x0
      13'h1830: dout <= 8'b10000000; // 6192 : 128 - 0x80 -- Background 0x83
      13'h1831: dout <= 8'b10000000; // 6193 : 128 - 0x80
      13'h1832: dout <= 8'b10000000; // 6194 : 128 - 0x80
      13'h1833: dout <= 8'b10000000; // 6195 : 128 - 0x80
      13'h1834: dout <= 8'b10000000; // 6196 : 128 - 0x80
      13'h1835: dout <= 8'b11100000; // 6197 : 224 - 0xe0
      13'h1836: dout <= 8'b00010000; // 6198 :  16 - 0x10
      13'h1837: dout <= 8'b11110000; // 6199 : 240 - 0xf0
      13'h1838: dout <= 8'b00000000; // 6200 :   0 - 0x0
      13'h1839: dout <= 8'b00000000; // 6201 :   0 - 0x0
      13'h183A: dout <= 8'b00000000; // 6202 :   0 - 0x0
      13'h183B: dout <= 8'b00000000; // 6203 :   0 - 0x0
      13'h183C: dout <= 8'b00000000; // 6204 :   0 - 0x0
      13'h183D: dout <= 8'b00000000; // 6205 :   0 - 0x0
      13'h183E: dout <= 8'b11100000; // 6206 : 224 - 0xe0
      13'h183F: dout <= 8'b00000000; // 6207 :   0 - 0x0
      13'h1840: dout <= 8'b00000011; // 6208 :   3 - 0x3 -- Background 0x84
      13'h1841: dout <= 8'b00001111; // 6209 :  15 - 0xf
      13'h1842: dout <= 8'b00011100; // 6210 :  28 - 0x1c
      13'h1843: dout <= 8'b00110000; // 6211 :  48 - 0x30
      13'h1844: dout <= 8'b00100000; // 6212 :  32 - 0x20
      13'h1845: dout <= 8'b01000000; // 6213 :  64 - 0x40
      13'h1846: dout <= 8'b01000000; // 6214 :  64 - 0x40
      13'h1847: dout <= 8'b01111111; // 6215 : 127 - 0x7f
      13'h1848: dout <= 8'b00000000; // 6216 :   0 - 0x0
      13'h1849: dout <= 8'b00000011; // 6217 :   3 - 0x3
      13'h184A: dout <= 8'b00001111; // 6218 :  15 - 0xf
      13'h184B: dout <= 8'b00011111; // 6219 :  31 - 0x1f
      13'h184C: dout <= 8'b00011111; // 6220 :  31 - 0x1f
      13'h184D: dout <= 8'b00111111; // 6221 :  63 - 0x3f
      13'h184E: dout <= 8'b00111111; // 6222 :  63 - 0x3f
      13'h184F: dout <= 8'b00000000; // 6223 :   0 - 0x0
      13'h1850: dout <= 8'b00000011; // 6224 :   3 - 0x3 -- Background 0x85
      13'h1851: dout <= 8'b00000110; // 6225 :   6 - 0x6
      13'h1852: dout <= 8'b00000110; // 6226 :   6 - 0x6
      13'h1853: dout <= 8'b00011100; // 6227 :  28 - 0x1c
      13'h1854: dout <= 8'b00011000; // 6228 :  24 - 0x18
      13'h1855: dout <= 8'b00110110; // 6229 :  54 - 0x36
      13'h1856: dout <= 8'b00110001; // 6230 :  49 - 0x31
      13'h1857: dout <= 8'b00001111; // 6231 :  15 - 0xf
      13'h1858: dout <= 8'b00000000; // 6232 :   0 - 0x0
      13'h1859: dout <= 8'b00000000; // 6233 :   0 - 0x0
      13'h185A: dout <= 8'b00000000; // 6234 :   0 - 0x0
      13'h185B: dout <= 8'b00000000; // 6235 :   0 - 0x0
      13'h185C: dout <= 8'b00000000; // 6236 :   0 - 0x0
      13'h185D: dout <= 8'b00001000; // 6237 :   8 - 0x8
      13'h185E: dout <= 8'b00001110; // 6238 :  14 - 0xe
      13'h185F: dout <= 8'b00000000; // 6239 :   0 - 0x0
      13'h1860: dout <= 8'b11000000; // 6240 : 192 - 0xc0 -- Background 0x86
      13'h1861: dout <= 8'b11110000; // 6241 : 240 - 0xf0
      13'h1862: dout <= 8'b00111000; // 6242 :  56 - 0x38
      13'h1863: dout <= 8'b00001110; // 6243 :  14 - 0xe
      13'h1864: dout <= 8'b00011110; // 6244 :  30 - 0x1e
      13'h1865: dout <= 8'b00011110; // 6245 :  30 - 0x1e
      13'h1866: dout <= 8'b00000010; // 6246 :   2 - 0x2
      13'h1867: dout <= 8'b11111110; // 6247 : 254 - 0xfe
      13'h1868: dout <= 8'b00000000; // 6248 :   0 - 0x0
      13'h1869: dout <= 8'b11000000; // 6249 : 192 - 0xc0
      13'h186A: dout <= 8'b11110000; // 6250 : 240 - 0xf0
      13'h186B: dout <= 8'b11110000; // 6251 : 240 - 0xf0
      13'h186C: dout <= 8'b11101100; // 6252 : 236 - 0xec
      13'h186D: dout <= 8'b11100000; // 6253 : 224 - 0xe0
      13'h186E: dout <= 8'b11111100; // 6254 : 252 - 0xfc
      13'h186F: dout <= 8'b00000000; // 6255 :   0 - 0x0
      13'h1870: dout <= 8'b11000000; // 6256 : 192 - 0xc0 -- Background 0x87
      13'h1871: dout <= 8'b01100000; // 6257 :  96 - 0x60
      13'h1872: dout <= 8'b01100000; // 6258 :  96 - 0x60
      13'h1873: dout <= 8'b00110000; // 6259 :  48 - 0x30
      13'h1874: dout <= 8'b00111110; // 6260 :  62 - 0x3e
      13'h1875: dout <= 8'b00011001; // 6261 :  25 - 0x19
      13'h1876: dout <= 8'b00110011; // 6262 :  51 - 0x33
      13'h1877: dout <= 8'b00111100; // 6263 :  60 - 0x3c
      13'h1878: dout <= 8'b00000000; // 6264 :   0 - 0x0
      13'h1879: dout <= 8'b00000000; // 6265 :   0 - 0x0
      13'h187A: dout <= 8'b00000000; // 6266 :   0 - 0x0
      13'h187B: dout <= 8'b00000000; // 6267 :   0 - 0x0
      13'h187C: dout <= 8'b00000000; // 6268 :   0 - 0x0
      13'h187D: dout <= 8'b00000110; // 6269 :   6 - 0x6
      13'h187E: dout <= 8'b00001100; // 6270 :  12 - 0xc
      13'h187F: dout <= 8'b00000000; // 6271 :   0 - 0x0
      13'h1880: dout <= 8'b00000011; // 6272 :   3 - 0x3 -- Background 0x88
      13'h1881: dout <= 8'b00000111; // 6273 :   7 - 0x7
      13'h1882: dout <= 8'b00000111; // 6274 :   7 - 0x7
      13'h1883: dout <= 8'b00001011; // 6275 :  11 - 0xb
      13'h1884: dout <= 8'b00010000; // 6276 :  16 - 0x10
      13'h1885: dout <= 8'b01100000; // 6277 :  96 - 0x60
      13'h1886: dout <= 8'b11110000; // 6278 : 240 - 0xf0
      13'h1887: dout <= 8'b11110000; // 6279 : 240 - 0xf0
      13'h1888: dout <= 8'b00000000; // 6280 :   0 - 0x0
      13'h1889: dout <= 8'b00000011; // 6281 :   3 - 0x3
      13'h188A: dout <= 8'b00000011; // 6282 :   3 - 0x3
      13'h188B: dout <= 8'b00000100; // 6283 :   4 - 0x4
      13'h188C: dout <= 8'b00001111; // 6284 :  15 - 0xf
      13'h188D: dout <= 8'b00011111; // 6285 :  31 - 0x1f
      13'h188E: dout <= 8'b01101111; // 6286 : 111 - 0x6f
      13'h188F: dout <= 8'b01101111; // 6287 : 111 - 0x6f
      13'h1890: dout <= 8'b11110000; // 6288 : 240 - 0xf0 -- Background 0x89
      13'h1891: dout <= 8'b11110000; // 6289 : 240 - 0xf0
      13'h1892: dout <= 8'b01100000; // 6290 :  96 - 0x60
      13'h1893: dout <= 8'b00010000; // 6291 :  16 - 0x10
      13'h1894: dout <= 8'b00001011; // 6292 :  11 - 0xb
      13'h1895: dout <= 8'b00000111; // 6293 :   7 - 0x7
      13'h1896: dout <= 8'b00000111; // 6294 :   7 - 0x7
      13'h1897: dout <= 8'b00000011; // 6295 :   3 - 0x3
      13'h1898: dout <= 8'b01101111; // 6296 : 111 - 0x6f
      13'h1899: dout <= 8'b01101111; // 6297 : 111 - 0x6f
      13'h189A: dout <= 8'b00011111; // 6298 :  31 - 0x1f
      13'h189B: dout <= 8'b00001111; // 6299 :  15 - 0xf
      13'h189C: dout <= 8'b00000100; // 6300 :   4 - 0x4
      13'h189D: dout <= 8'b00000011; // 6301 :   3 - 0x3
      13'h189E: dout <= 8'b00000011; // 6302 :   3 - 0x3
      13'h189F: dout <= 8'b00000000; // 6303 :   0 - 0x0
      13'h18A0: dout <= 8'b00000000; // 6304 :   0 - 0x0 -- Background 0x8a
      13'h18A1: dout <= 8'b00011100; // 6305 :  28 - 0x1c
      13'h18A2: dout <= 8'b00111111; // 6306 :  63 - 0x3f
      13'h18A3: dout <= 8'b01111000; // 6307 : 120 - 0x78
      13'h18A4: dout <= 8'b01110000; // 6308 : 112 - 0x70
      13'h18A5: dout <= 8'b01100000; // 6309 :  96 - 0x60
      13'h18A6: dout <= 8'b00100000; // 6310 :  32 - 0x20
      13'h18A7: dout <= 8'b00100000; // 6311 :  32 - 0x20
      13'h18A8: dout <= 8'b00000000; // 6312 :   0 - 0x0
      13'h18A9: dout <= 8'b00000000; // 6313 :   0 - 0x0
      13'h18AA: dout <= 8'b00011000; // 6314 :  24 - 0x18
      13'h18AB: dout <= 8'b00110111; // 6315 :  55 - 0x37
      13'h18AC: dout <= 8'b00101111; // 6316 :  47 - 0x2f
      13'h18AD: dout <= 8'b00011111; // 6317 :  31 - 0x1f
      13'h18AE: dout <= 8'b00011111; // 6318 :  31 - 0x1f
      13'h18AF: dout <= 8'b00011111; // 6319 :  31 - 0x1f
      13'h18B0: dout <= 8'b00100000; // 6320 :  32 - 0x20 -- Background 0x8b
      13'h18B1: dout <= 8'b00100000; // 6321 :  32 - 0x20
      13'h18B2: dout <= 8'b01100000; // 6322 :  96 - 0x60
      13'h18B3: dout <= 8'b01110000; // 6323 : 112 - 0x70
      13'h18B4: dout <= 8'b01111000; // 6324 : 120 - 0x78
      13'h18B5: dout <= 8'b00111111; // 6325 :  63 - 0x3f
      13'h18B6: dout <= 8'b00011100; // 6326 :  28 - 0x1c
      13'h18B7: dout <= 8'b00000000; // 6327 :   0 - 0x0
      13'h18B8: dout <= 8'b00011111; // 6328 :  31 - 0x1f
      13'h18B9: dout <= 8'b00011111; // 6329 :  31 - 0x1f
      13'h18BA: dout <= 8'b00011111; // 6330 :  31 - 0x1f
      13'h18BB: dout <= 8'b00101111; // 6331 :  47 - 0x2f
      13'h18BC: dout <= 8'b00110111; // 6332 :  55 - 0x37
      13'h18BD: dout <= 8'b00011000; // 6333 :  24 - 0x18
      13'h18BE: dout <= 8'b00000000; // 6334 :   0 - 0x0
      13'h18BF: dout <= 8'b00000000; // 6335 :   0 - 0x0
      13'h18C0: dout <= 8'b00000011; // 6336 :   3 - 0x3 -- Background 0x8c
      13'h18C1: dout <= 8'b00001100; // 6337 :  12 - 0xc
      13'h18C2: dout <= 8'b00011110; // 6338 :  30 - 0x1e
      13'h18C3: dout <= 8'b00100110; // 6339 :  38 - 0x26
      13'h18C4: dout <= 8'b01000110; // 6340 :  70 - 0x46
      13'h18C5: dout <= 8'b01100100; // 6341 : 100 - 0x64
      13'h18C6: dout <= 8'b01110000; // 6342 : 112 - 0x70
      13'h18C7: dout <= 8'b11110000; // 6343 : 240 - 0xf0
      13'h18C8: dout <= 8'b00000000; // 6344 :   0 - 0x0
      13'h18C9: dout <= 8'b00000011; // 6345 :   3 - 0x3
      13'h18CA: dout <= 8'b00000001; // 6346 :   1 - 0x1
      13'h18CB: dout <= 8'b00011001; // 6347 :  25 - 0x19
      13'h18CC: dout <= 8'b00111001; // 6348 :  57 - 0x39
      13'h18CD: dout <= 8'b00011011; // 6349 :  27 - 0x1b
      13'h18CE: dout <= 8'b00001111; // 6350 :  15 - 0xf
      13'h18CF: dout <= 8'b00001111; // 6351 :  15 - 0xf
      13'h18D0: dout <= 8'b10101010; // 6352 : 170 - 0xaa -- Background 0x8d
      13'h18D1: dout <= 8'b11111111; // 6353 : 255 - 0xff
      13'h18D2: dout <= 8'b01111111; // 6354 : 127 - 0x7f
      13'h18D3: dout <= 8'b00111001; // 6355 :  57 - 0x39
      13'h18D4: dout <= 8'b00011001; // 6356 :  25 - 0x19
      13'h18D5: dout <= 8'b00001011; // 6357 :  11 - 0xb
      13'h18D6: dout <= 8'b00001000; // 6358 :   8 - 0x8
      13'h18D7: dout <= 8'b00000111; // 6359 :   7 - 0x7
      13'h18D8: dout <= 8'b01111111; // 6360 : 127 - 0x7f
      13'h18D9: dout <= 8'b01111111; // 6361 : 127 - 0x7f
      13'h18DA: dout <= 8'b00111111; // 6362 :  63 - 0x3f
      13'h18DB: dout <= 8'b00010111; // 6363 :  23 - 0x17
      13'h18DC: dout <= 8'b00000110; // 6364 :   6 - 0x6
      13'h18DD: dout <= 8'b00000100; // 6365 :   4 - 0x4
      13'h18DE: dout <= 8'b00000111; // 6366 :   7 - 0x7
      13'h18DF: dout <= 8'b00000000; // 6367 :   0 - 0x0
      13'h18E0: dout <= 8'b11000000; // 6368 : 192 - 0xc0 -- Background 0x8e
      13'h18E1: dout <= 8'b00110000; // 6369 :  48 - 0x30
      13'h18E2: dout <= 8'b00001000; // 6370 :   8 - 0x8
      13'h18E3: dout <= 8'b01000100; // 6371 :  68 - 0x44
      13'h18E4: dout <= 8'b01100010; // 6372 :  98 - 0x62
      13'h18E5: dout <= 8'b01100010; // 6373 :  98 - 0x62
      13'h18E6: dout <= 8'b00000001; // 6374 :   1 - 0x1
      13'h18E7: dout <= 8'b00111111; // 6375 :  63 - 0x3f
      13'h18E8: dout <= 8'b00000000; // 6376 :   0 - 0x0
      13'h18E9: dout <= 8'b11000000; // 6377 : 192 - 0xc0
      13'h18EA: dout <= 8'b11110000; // 6378 : 240 - 0xf0
      13'h18EB: dout <= 8'b10111000; // 6379 : 184 - 0xb8
      13'h18EC: dout <= 8'b10011100; // 6380 : 156 - 0x9c
      13'h18ED: dout <= 8'b11111100; // 6381 : 252 - 0xfc
      13'h18EE: dout <= 8'b11111110; // 6382 : 254 - 0xfe
      13'h18EF: dout <= 8'b11000000; // 6383 : 192 - 0xc0
      13'h18F0: dout <= 8'b10001011; // 6384 : 139 - 0x8b -- Background 0x8f
      13'h18F1: dout <= 8'b11000001; // 6385 : 193 - 0xc1
      13'h18F2: dout <= 8'b11111110; // 6386 : 254 - 0xfe
      13'h18F3: dout <= 8'b11111100; // 6387 : 252 - 0xfc
      13'h18F4: dout <= 8'b11110000; // 6388 : 240 - 0xf0
      13'h18F5: dout <= 8'b11110000; // 6389 : 240 - 0xf0
      13'h18F6: dout <= 8'b11111000; // 6390 : 248 - 0xf8
      13'h18F7: dout <= 8'b11110000; // 6391 : 240 - 0xf0
      13'h18F8: dout <= 8'b11111110; // 6392 : 254 - 0xfe
      13'h18F9: dout <= 8'b11111110; // 6393 : 254 - 0xfe
      13'h18FA: dout <= 8'b11111000; // 6394 : 248 - 0xf8
      13'h18FB: dout <= 8'b11110000; // 6395 : 240 - 0xf0
      13'h18FC: dout <= 8'b11000000; // 6396 : 192 - 0xc0
      13'h18FD: dout <= 8'b00000000; // 6397 :   0 - 0x0
      13'h18FE: dout <= 8'b00000000; // 6398 :   0 - 0x0
      13'h18FF: dout <= 8'b10000000; // 6399 : 128 - 0x80
      13'h1900: dout <= 8'b00000011; // 6400 :   3 - 0x3 -- Background 0x90
      13'h1901: dout <= 8'b00001110; // 6401 :  14 - 0xe
      13'h1902: dout <= 8'b00010110; // 6402 :  22 - 0x16
      13'h1903: dout <= 8'b00100110; // 6403 :  38 - 0x26
      13'h1904: dout <= 8'b01100011; // 6404 :  99 - 0x63
      13'h1905: dout <= 8'b01110010; // 6405 : 114 - 0x72
      13'h1906: dout <= 8'b01110000; // 6406 : 112 - 0x70
      13'h1907: dout <= 8'b11010000; // 6407 : 208 - 0xd0
      13'h1908: dout <= 8'b00000000; // 6408 :   0 - 0x0
      13'h1909: dout <= 8'b00000001; // 6409 :   1 - 0x1
      13'h190A: dout <= 8'b00001001; // 6410 :   9 - 0x9
      13'h190B: dout <= 8'b00011001; // 6411 :  25 - 0x19
      13'h190C: dout <= 8'b00011100; // 6412 :  28 - 0x1c
      13'h190D: dout <= 8'b00001101; // 6413 :  13 - 0xd
      13'h190E: dout <= 8'b00001111; // 6414 :  15 - 0xf
      13'h190F: dout <= 8'b00101111; // 6415 :  47 - 0x2f
      13'h1910: dout <= 8'b10101010; // 6416 : 170 - 0xaa -- Background 0x91
      13'h1911: dout <= 8'b11111111; // 6417 : 255 - 0xff
      13'h1912: dout <= 8'b01111111; // 6418 : 127 - 0x7f
      13'h1913: dout <= 8'b00111100; // 6419 :  60 - 0x3c
      13'h1914: dout <= 8'b00011100; // 6420 :  28 - 0x1c
      13'h1915: dout <= 8'b00000100; // 6421 :   4 - 0x4
      13'h1916: dout <= 8'b00000010; // 6422 :   2 - 0x2
      13'h1917: dout <= 8'b00000001; // 6423 :   1 - 0x1
      13'h1918: dout <= 8'b01111111; // 6424 : 127 - 0x7f
      13'h1919: dout <= 8'b01111111; // 6425 : 127 - 0x7f
      13'h191A: dout <= 8'b00111111; // 6426 :  63 - 0x3f
      13'h191B: dout <= 8'b00011011; // 6427 :  27 - 0x1b
      13'h191C: dout <= 8'b00000011; // 6428 :   3 - 0x3
      13'h191D: dout <= 8'b00000011; // 6429 :   3 - 0x3
      13'h191E: dout <= 8'b00000001; // 6430 :   1 - 0x1
      13'h191F: dout <= 8'b00000000; // 6431 :   0 - 0x0
      13'h1920: dout <= 8'b11000000; // 6432 : 192 - 0xc0 -- Background 0x92
      13'h1921: dout <= 8'b00110000; // 6433 :  48 - 0x30
      13'h1922: dout <= 8'b00001000; // 6434 :   8 - 0x8
      13'h1923: dout <= 8'b00100100; // 6435 :  36 - 0x24
      13'h1924: dout <= 8'b00110010; // 6436 :  50 - 0x32
      13'h1925: dout <= 8'b00110010; // 6437 :  50 - 0x32
      13'h1926: dout <= 8'b00000001; // 6438 :   1 - 0x1
      13'h1927: dout <= 8'b00011111; // 6439 :  31 - 0x1f
      13'h1928: dout <= 8'b00000000; // 6440 :   0 - 0x0
      13'h1929: dout <= 8'b11000000; // 6441 : 192 - 0xc0
      13'h192A: dout <= 8'b11110000; // 6442 : 240 - 0xf0
      13'h192B: dout <= 8'b11011000; // 6443 : 216 - 0xd8
      13'h192C: dout <= 8'b11001100; // 6444 : 204 - 0xcc
      13'h192D: dout <= 8'b11111100; // 6445 : 252 - 0xfc
      13'h192E: dout <= 8'b11111110; // 6446 : 254 - 0xfe
      13'h192F: dout <= 8'b11100000; // 6447 : 224 - 0xe0
      13'h1930: dout <= 8'b10001011; // 6448 : 139 - 0x8b -- Background 0x93
      13'h1931: dout <= 8'b11000001; // 6449 : 193 - 0xc1
      13'h1932: dout <= 8'b11111110; // 6450 : 254 - 0xfe
      13'h1933: dout <= 8'b11111100; // 6451 : 252 - 0xfc
      13'h1934: dout <= 8'b11110000; // 6452 : 240 - 0xf0
      13'h1935: dout <= 8'b11000000; // 6453 : 192 - 0xc0
      13'h1936: dout <= 8'b00100000; // 6454 :  32 - 0x20
      13'h1937: dout <= 8'b11100000; // 6455 : 224 - 0xe0
      13'h1938: dout <= 8'b11111110; // 6456 : 254 - 0xfe
      13'h1939: dout <= 8'b11111110; // 6457 : 254 - 0xfe
      13'h193A: dout <= 8'b11111000; // 6458 : 248 - 0xf8
      13'h193B: dout <= 8'b01110000; // 6459 : 112 - 0x70
      13'h193C: dout <= 8'b01000000; // 6460 :  64 - 0x40
      13'h193D: dout <= 8'b00000000; // 6461 :   0 - 0x0
      13'h193E: dout <= 8'b11000000; // 6462 : 192 - 0xc0
      13'h193F: dout <= 8'b00100000; // 6463 :  32 - 0x20
      13'h1940: dout <= 8'b00000011; // 6464 :   3 - 0x3 -- Background 0x94
      13'h1941: dout <= 8'b00001111; // 6465 :  15 - 0xf
      13'h1942: dout <= 8'b00010011; // 6466 :  19 - 0x13
      13'h1943: dout <= 8'b00110001; // 6467 :  49 - 0x31
      13'h1944: dout <= 8'b01111001; // 6468 : 121 - 0x79
      13'h1945: dout <= 8'b01011001; // 6469 :  89 - 0x59
      13'h1946: dout <= 8'b01001000; // 6470 :  72 - 0x48
      13'h1947: dout <= 8'b11001100; // 6471 : 204 - 0xcc
      13'h1948: dout <= 8'b00000000; // 6472 :   0 - 0x0
      13'h1949: dout <= 8'b00000000; // 6473 :   0 - 0x0
      13'h194A: dout <= 8'b00001100; // 6474 :  12 - 0xc
      13'h194B: dout <= 8'b00001110; // 6475 :  14 - 0xe
      13'h194C: dout <= 8'b00000110; // 6476 :   6 - 0x6
      13'h194D: dout <= 8'b00100110; // 6477 :  38 - 0x26
      13'h194E: dout <= 8'b00110111; // 6478 :  55 - 0x37
      13'h194F: dout <= 8'b00110011; // 6479 :  51 - 0x33
      13'h1950: dout <= 8'b10010101; // 6480 : 149 - 0x95 -- Background 0x95
      13'h1951: dout <= 8'b11111111; // 6481 : 255 - 0xff
      13'h1952: dout <= 8'b01111111; // 6482 : 127 - 0x7f
      13'h1953: dout <= 8'b00111110; // 6483 :  62 - 0x3e
      13'h1954: dout <= 8'b00011111; // 6484 :  31 - 0x1f
      13'h1955: dout <= 8'b00001111; // 6485 :  15 - 0xf
      13'h1956: dout <= 8'b00001111; // 6486 :  15 - 0xf
      13'h1957: dout <= 8'b00000111; // 6487 :   7 - 0x7
      13'h1958: dout <= 8'b01111111; // 6488 : 127 - 0x7f
      13'h1959: dout <= 8'b01111111; // 6489 : 127 - 0x7f
      13'h195A: dout <= 8'b00111111; // 6490 :  63 - 0x3f
      13'h195B: dout <= 8'b00011111; // 6491 :  31 - 0x1f
      13'h195C: dout <= 8'b00001110; // 6492 :  14 - 0xe
      13'h195D: dout <= 8'b00000000; // 6493 :   0 - 0x0
      13'h195E: dout <= 8'b00000000; // 6494 :   0 - 0x0
      13'h195F: dout <= 8'b00000000; // 6495 :   0 - 0x0
      13'h1960: dout <= 8'b11000000; // 6496 : 192 - 0xc0 -- Background 0x96
      13'h1961: dout <= 8'b00110000; // 6497 :  48 - 0x30
      13'h1962: dout <= 8'b00001000; // 6498 :   8 - 0x8
      13'h1963: dout <= 8'b10010100; // 6499 : 148 - 0x94
      13'h1964: dout <= 8'b10011010; // 6500 : 154 - 0x9a
      13'h1965: dout <= 8'b00011010; // 6501 :  26 - 0x1a
      13'h1966: dout <= 8'b00000001; // 6502 :   1 - 0x1
      13'h1967: dout <= 8'b00001111; // 6503 :  15 - 0xf
      13'h1968: dout <= 8'b00000000; // 6504 :   0 - 0x0
      13'h1969: dout <= 8'b11000000; // 6505 : 192 - 0xc0
      13'h196A: dout <= 8'b11110000; // 6506 : 240 - 0xf0
      13'h196B: dout <= 8'b01101000; // 6507 : 104 - 0x68
      13'h196C: dout <= 8'b01100100; // 6508 : 100 - 0x64
      13'h196D: dout <= 8'b11111100; // 6509 : 252 - 0xfc
      13'h196E: dout <= 8'b11111110; // 6510 : 254 - 0xfe
      13'h196F: dout <= 8'b11110000; // 6511 : 240 - 0xf0
      13'h1970: dout <= 8'b01000101; // 6512 :  69 - 0x45 -- Background 0x97
      13'h1971: dout <= 8'b11100001; // 6513 : 225 - 0xe1
      13'h1972: dout <= 8'b11111110; // 6514 : 254 - 0xfe
      13'h1973: dout <= 8'b01111100; // 6515 : 124 - 0x7c
      13'h1974: dout <= 8'b00110000; // 6516 :  48 - 0x30
      13'h1975: dout <= 8'b00110000; // 6517 :  48 - 0x30
      13'h1976: dout <= 8'b10001000; // 6518 : 136 - 0x88
      13'h1977: dout <= 8'b01111000; // 6519 : 120 - 0x78
      13'h1978: dout <= 8'b11111111; // 6520 : 255 - 0xff
      13'h1979: dout <= 8'b11111110; // 6521 : 254 - 0xfe
      13'h197A: dout <= 8'b11111100; // 6522 : 252 - 0xfc
      13'h197B: dout <= 8'b10110000; // 6523 : 176 - 0xb0
      13'h197C: dout <= 8'b11000000; // 6524 : 192 - 0xc0
      13'h197D: dout <= 8'b11000000; // 6525 : 192 - 0xc0
      13'h197E: dout <= 8'b01110000; // 6526 : 112 - 0x70
      13'h197F: dout <= 8'b00001000; // 6527 :   8 - 0x8
      13'h1980: dout <= 8'b00000001; // 6528 :   1 - 0x1 -- Background 0x98
      13'h1981: dout <= 8'b00000000; // 6529 :   0 - 0x0
      13'h1982: dout <= 8'b00000000; // 6530 :   0 - 0x0
      13'h1983: dout <= 8'b00000000; // 6531 :   0 - 0x0
      13'h1984: dout <= 8'b00000001; // 6532 :   1 - 0x1
      13'h1985: dout <= 8'b00000001; // 6533 :   1 - 0x1
      13'h1986: dout <= 8'b00000010; // 6534 :   2 - 0x2
      13'h1987: dout <= 8'b00000110; // 6535 :   6 - 0x6
      13'h1988: dout <= 8'b00000000; // 6536 :   0 - 0x0
      13'h1989: dout <= 8'b00000001; // 6537 :   1 - 0x1
      13'h198A: dout <= 8'b00000000; // 6538 :   0 - 0x0
      13'h198B: dout <= 8'b00000000; // 6539 :   0 - 0x0
      13'h198C: dout <= 8'b00000000; // 6540 :   0 - 0x0
      13'h198D: dout <= 8'b00000000; // 6541 :   0 - 0x0
      13'h198E: dout <= 8'b00000001; // 6542 :   1 - 0x1
      13'h198F: dout <= 8'b00000011; // 6543 :   3 - 0x3
      13'h1990: dout <= 8'b01111000; // 6544 : 120 - 0x78 -- Background 0x99
      13'h1991: dout <= 8'b00101010; // 6545 :  42 - 0x2a
      13'h1992: dout <= 8'b01010100; // 6546 :  84 - 0x54
      13'h1993: dout <= 8'b00101001; // 6547 :  41 - 0x29
      13'h1994: dout <= 8'b00101111; // 6548 :  47 - 0x2f
      13'h1995: dout <= 8'b00110111; // 6549 :  55 - 0x37
      13'h1996: dout <= 8'b00000011; // 6550 :   3 - 0x3
      13'h1997: dout <= 8'b00000111; // 6551 :   7 - 0x7
      13'h1998: dout <= 8'b00000111; // 6552 :   7 - 0x7
      13'h1999: dout <= 8'b00010111; // 6553 :  23 - 0x17
      13'h199A: dout <= 8'b00101111; // 6554 :  47 - 0x2f
      13'h199B: dout <= 8'b00011110; // 6555 :  30 - 0x1e
      13'h199C: dout <= 8'b00010001; // 6556 :  17 - 0x11
      13'h199D: dout <= 8'b00000000; // 6557 :   0 - 0x0
      13'h199E: dout <= 8'b00000001; // 6558 :   1 - 0x1
      13'h199F: dout <= 8'b00000000; // 6559 :   0 - 0x0
      13'h19A0: dout <= 8'b10110000; // 6560 : 176 - 0xb0 -- Background 0x9a
      13'h19A1: dout <= 8'b11101000; // 6561 : 232 - 0xe8
      13'h19A2: dout <= 8'b10001100; // 6562 : 140 - 0x8c
      13'h19A3: dout <= 8'b10011110; // 6563 : 158 - 0x9e
      13'h19A4: dout <= 8'b00011111; // 6564 :  31 - 0x1f
      13'h19A5: dout <= 8'b00001111; // 6565 :  15 - 0xf
      13'h19A6: dout <= 8'b10010110; // 6566 : 150 - 0x96
      13'h19A7: dout <= 8'b00011100; // 6567 :  28 - 0x1c
      13'h19A8: dout <= 8'b00000000; // 6568 :   0 - 0x0
      13'h19A9: dout <= 8'b00010000; // 6569 :  16 - 0x10
      13'h19AA: dout <= 8'b01111000; // 6570 : 120 - 0x78
      13'h19AB: dout <= 8'b01110100; // 6571 : 116 - 0x74
      13'h19AC: dout <= 8'b11111110; // 6572 : 254 - 0xfe
      13'h19AD: dout <= 8'b11111000; // 6573 : 248 - 0xf8
      13'h19AE: dout <= 8'b11111100; // 6574 : 252 - 0xfc
      13'h19AF: dout <= 8'b11111000; // 6575 : 248 - 0xf8
      13'h19B0: dout <= 8'b00001100; // 6576 :  12 - 0xc -- Background 0x9b
      13'h19B1: dout <= 8'b00111000; // 6577 :  56 - 0x38
      13'h19B2: dout <= 8'b11101000; // 6578 : 232 - 0xe8
      13'h19B3: dout <= 8'b11010000; // 6579 : 208 - 0xd0
      13'h19B4: dout <= 8'b11100000; // 6580 : 224 - 0xe0
      13'h19B5: dout <= 8'b10000000; // 6581 : 128 - 0x80
      13'h19B6: dout <= 8'b00000000; // 6582 :   0 - 0x0
      13'h19B7: dout <= 8'b10000000; // 6583 : 128 - 0x80
      13'h19B8: dout <= 8'b11111000; // 6584 : 248 - 0xf8
      13'h19B9: dout <= 8'b11010000; // 6585 : 208 - 0xd0
      13'h19BA: dout <= 8'b00110000; // 6586 :  48 - 0x30
      13'h19BB: dout <= 8'b01100000; // 6587 :  96 - 0x60
      13'h19BC: dout <= 8'b10000000; // 6588 : 128 - 0x80
      13'h19BD: dout <= 8'b00000000; // 6589 :   0 - 0x0
      13'h19BE: dout <= 8'b00000000; // 6590 :   0 - 0x0
      13'h19BF: dout <= 8'b00000000; // 6591 :   0 - 0x0
      13'h19C0: dout <= 8'b00000001; // 6592 :   1 - 0x1 -- Background 0x9c
      13'h19C1: dout <= 8'b00000000; // 6593 :   0 - 0x0
      13'h19C2: dout <= 8'b00000000; // 6594 :   0 - 0x0
      13'h19C3: dout <= 8'b00000000; // 6595 :   0 - 0x0
      13'h19C4: dout <= 8'b00000001; // 6596 :   1 - 0x1
      13'h19C5: dout <= 8'b00000001; // 6597 :   1 - 0x1
      13'h19C6: dout <= 8'b00000010; // 6598 :   2 - 0x2
      13'h19C7: dout <= 8'b00000110; // 6599 :   6 - 0x6
      13'h19C8: dout <= 8'b00000000; // 6600 :   0 - 0x0
      13'h19C9: dout <= 8'b00000001; // 6601 :   1 - 0x1
      13'h19CA: dout <= 8'b00000000; // 6602 :   0 - 0x0
      13'h19CB: dout <= 8'b00000000; // 6603 :   0 - 0x0
      13'h19CC: dout <= 8'b00000000; // 6604 :   0 - 0x0
      13'h19CD: dout <= 8'b00000000; // 6605 :   0 - 0x0
      13'h19CE: dout <= 8'b00000001; // 6606 :   1 - 0x1
      13'h19CF: dout <= 8'b00000011; // 6607 :   3 - 0x3
      13'h19D0: dout <= 8'b01111000; // 6608 : 120 - 0x78 -- Background 0x9d
      13'h19D1: dout <= 8'b00101010; // 6609 :  42 - 0x2a
      13'h19D2: dout <= 8'b01010100; // 6610 :  84 - 0x54
      13'h19D3: dout <= 8'b00101001; // 6611 :  41 - 0x29
      13'h19D4: dout <= 8'b00101111; // 6612 :  47 - 0x2f
      13'h19D5: dout <= 8'b00111100; // 6613 :  60 - 0x3c
      13'h19D6: dout <= 8'b00011110; // 6614 :  30 - 0x1e
      13'h19D7: dout <= 8'b00000000; // 6615 :   0 - 0x0
      13'h19D8: dout <= 8'b00000111; // 6616 :   7 - 0x7
      13'h19D9: dout <= 8'b00010111; // 6617 :  23 - 0x17
      13'h19DA: dout <= 8'b00101111; // 6618 :  47 - 0x2f
      13'h19DB: dout <= 8'b00011110; // 6619 :  30 - 0x1e
      13'h19DC: dout <= 8'b00010000; // 6620 :  16 - 0x10
      13'h19DD: dout <= 8'b00000100; // 6621 :   4 - 0x4
      13'h19DE: dout <= 8'b00000000; // 6622 :   0 - 0x0
      13'h19DF: dout <= 8'b00000000; // 6623 :   0 - 0x0
      13'h19E0: dout <= 8'b10110000; // 6624 : 176 - 0xb0 -- Background 0x9e
      13'h19E1: dout <= 8'b11101000; // 6625 : 232 - 0xe8
      13'h19E2: dout <= 8'b10001100; // 6626 : 140 - 0x8c
      13'h19E3: dout <= 8'b10011110; // 6627 : 158 - 0x9e
      13'h19E4: dout <= 8'b00011111; // 6628 :  31 - 0x1f
      13'h19E5: dout <= 8'b00001111; // 6629 :  15 - 0xf
      13'h19E6: dout <= 8'b10010110; // 6630 : 150 - 0x96
      13'h19E7: dout <= 8'b00011100; // 6631 :  28 - 0x1c
      13'h19E8: dout <= 8'b00000000; // 6632 :   0 - 0x0
      13'h19E9: dout <= 8'b00010000; // 6633 :  16 - 0x10
      13'h19EA: dout <= 8'b01111000; // 6634 : 120 - 0x78
      13'h19EB: dout <= 8'b01110100; // 6635 : 116 - 0x74
      13'h19EC: dout <= 8'b11111110; // 6636 : 254 - 0xfe
      13'h19ED: dout <= 8'b11111000; // 6637 : 248 - 0xf8
      13'h19EE: dout <= 8'b11111100; // 6638 : 252 - 0xfc
      13'h19EF: dout <= 8'b11111000; // 6639 : 248 - 0xf8
      13'h19F0: dout <= 8'b00001100; // 6640 :  12 - 0xc -- Background 0x9f
      13'h19F1: dout <= 8'b00111000; // 6641 :  56 - 0x38
      13'h19F2: dout <= 8'b11101000; // 6642 : 232 - 0xe8
      13'h19F3: dout <= 8'b11110000; // 6643 : 240 - 0xf0
      13'h19F4: dout <= 8'b11000000; // 6644 : 192 - 0xc0
      13'h19F5: dout <= 8'b01110000; // 6645 : 112 - 0x70
      13'h19F6: dout <= 8'b11000000; // 6646 : 192 - 0xc0
      13'h19F7: dout <= 8'b00000000; // 6647 :   0 - 0x0
      13'h19F8: dout <= 8'b11111000; // 6648 : 248 - 0xf8
      13'h19F9: dout <= 8'b11010000; // 6649 : 208 - 0xd0
      13'h19FA: dout <= 8'b00110000; // 6650 :  48 - 0x30
      13'h19FB: dout <= 8'b11000000; // 6651 : 192 - 0xc0
      13'h19FC: dout <= 8'b00000000; // 6652 :   0 - 0x0
      13'h19FD: dout <= 8'b00000000; // 6653 :   0 - 0x0
      13'h19FE: dout <= 8'b00000000; // 6654 :   0 - 0x0
      13'h19FF: dout <= 8'b00000000; // 6655 :   0 - 0x0
      13'h1A00: dout <= 8'b00000011; // 6656 :   3 - 0x3 -- Background 0xa0
      13'h1A01: dout <= 8'b00001111; // 6657 :  15 - 0xf
      13'h1A02: dout <= 8'b00011100; // 6658 :  28 - 0x1c
      13'h1A03: dout <= 8'b00110000; // 6659 :  48 - 0x30
      13'h1A04: dout <= 8'b01100000; // 6660 :  96 - 0x60
      13'h1A05: dout <= 8'b01100000; // 6661 :  96 - 0x60
      13'h1A06: dout <= 8'b11000000; // 6662 : 192 - 0xc0
      13'h1A07: dout <= 8'b11000000; // 6663 : 192 - 0xc0
      13'h1A08: dout <= 8'b00000000; // 6664 :   0 - 0x0
      13'h1A09: dout <= 8'b00000011; // 6665 :   3 - 0x3
      13'h1A0A: dout <= 8'b00001111; // 6666 :  15 - 0xf
      13'h1A0B: dout <= 8'b00011111; // 6667 :  31 - 0x1f
      13'h1A0C: dout <= 8'b00111111; // 6668 :  63 - 0x3f
      13'h1A0D: dout <= 8'b00111111; // 6669 :  63 - 0x3f
      13'h1A0E: dout <= 8'b01111111; // 6670 : 127 - 0x7f
      13'h1A0F: dout <= 8'b01111111; // 6671 : 127 - 0x7f
      13'h1A10: dout <= 8'b11000000; // 6672 : 192 - 0xc0 -- Background 0xa1
      13'h1A11: dout <= 8'b11000000; // 6673 : 192 - 0xc0
      13'h1A12: dout <= 8'b01100000; // 6674 :  96 - 0x60
      13'h1A13: dout <= 8'b01100000; // 6675 :  96 - 0x60
      13'h1A14: dout <= 8'b00110000; // 6676 :  48 - 0x30
      13'h1A15: dout <= 8'b00011010; // 6677 :  26 - 0x1a
      13'h1A16: dout <= 8'b00001101; // 6678 :  13 - 0xd
      13'h1A17: dout <= 8'b00000011; // 6679 :   3 - 0x3
      13'h1A18: dout <= 8'b01111111; // 6680 : 127 - 0x7f
      13'h1A19: dout <= 8'b01111111; // 6681 : 127 - 0x7f
      13'h1A1A: dout <= 8'b00111111; // 6682 :  63 - 0x3f
      13'h1A1B: dout <= 8'b00111111; // 6683 :  63 - 0x3f
      13'h1A1C: dout <= 8'b00011111; // 6684 :  31 - 0x1f
      13'h1A1D: dout <= 8'b00000101; // 6685 :   5 - 0x5
      13'h1A1E: dout <= 8'b00000010; // 6686 :   2 - 0x2
      13'h1A1F: dout <= 8'b00000000; // 6687 :   0 - 0x0
      13'h1A20: dout <= 8'b11000000; // 6688 : 192 - 0xc0 -- Background 0xa2
      13'h1A21: dout <= 8'b11110000; // 6689 : 240 - 0xf0
      13'h1A22: dout <= 8'b00111000; // 6690 :  56 - 0x38
      13'h1A23: dout <= 8'b00001100; // 6691 :  12 - 0xc
      13'h1A24: dout <= 8'b00000110; // 6692 :   6 - 0x6
      13'h1A25: dout <= 8'b00000010; // 6693 :   2 - 0x2
      13'h1A26: dout <= 8'b00000101; // 6694 :   5 - 0x5
      13'h1A27: dout <= 8'b00000011; // 6695 :   3 - 0x3
      13'h1A28: dout <= 8'b00000000; // 6696 :   0 - 0x0
      13'h1A29: dout <= 8'b11000000; // 6697 : 192 - 0xc0
      13'h1A2A: dout <= 8'b11110000; // 6698 : 240 - 0xf0
      13'h1A2B: dout <= 8'b11111000; // 6699 : 248 - 0xf8
      13'h1A2C: dout <= 8'b11111000; // 6700 : 248 - 0xf8
      13'h1A2D: dout <= 8'b11111100; // 6701 : 252 - 0xfc
      13'h1A2E: dout <= 8'b11111010; // 6702 : 250 - 0xfa
      13'h1A2F: dout <= 8'b11111100; // 6703 : 252 - 0xfc
      13'h1A30: dout <= 8'b00000101; // 6704 :   5 - 0x5 -- Background 0xa3
      13'h1A31: dout <= 8'b00001011; // 6705 :  11 - 0xb
      13'h1A32: dout <= 8'b00010110; // 6706 :  22 - 0x16
      13'h1A33: dout <= 8'b00101010; // 6707 :  42 - 0x2a
      13'h1A34: dout <= 8'b01010100; // 6708 :  84 - 0x54
      13'h1A35: dout <= 8'b10101000; // 6709 : 168 - 0xa8
      13'h1A36: dout <= 8'b01110000; // 6710 : 112 - 0x70
      13'h1A37: dout <= 8'b11000000; // 6711 : 192 - 0xc0
      13'h1A38: dout <= 8'b11111010; // 6712 : 250 - 0xfa
      13'h1A39: dout <= 8'b11110100; // 6713 : 244 - 0xf4
      13'h1A3A: dout <= 8'b11101000; // 6714 : 232 - 0xe8
      13'h1A3B: dout <= 8'b11010100; // 6715 : 212 - 0xd4
      13'h1A3C: dout <= 8'b10101000; // 6716 : 168 - 0xa8
      13'h1A3D: dout <= 8'b01010000; // 6717 :  80 - 0x50
      13'h1A3E: dout <= 8'b10000000; // 6718 : 128 - 0x80
      13'h1A3F: dout <= 8'b00000000; // 6719 :   0 - 0x0
      13'h1A40: dout <= 8'b00000000; // 6720 :   0 - 0x0 -- Background 0xa4
      13'h1A41: dout <= 8'b00001111; // 6721 :  15 - 0xf
      13'h1A42: dout <= 8'b00011111; // 6722 :  31 - 0x1f
      13'h1A43: dout <= 8'b00110001; // 6723 :  49 - 0x31
      13'h1A44: dout <= 8'b00111111; // 6724 :  63 - 0x3f
      13'h1A45: dout <= 8'b01111111; // 6725 : 127 - 0x7f
      13'h1A46: dout <= 8'b11111111; // 6726 : 255 - 0xff
      13'h1A47: dout <= 8'b11011111; // 6727 : 223 - 0xdf
      13'h1A48: dout <= 8'b00000000; // 6728 :   0 - 0x0
      13'h1A49: dout <= 8'b00000000; // 6729 :   0 - 0x0
      13'h1A4A: dout <= 8'b00000000; // 6730 :   0 - 0x0
      13'h1A4B: dout <= 8'b00001110; // 6731 :  14 - 0xe
      13'h1A4C: dout <= 8'b00000000; // 6732 :   0 - 0x0
      13'h1A4D: dout <= 8'b00001010; // 6733 :  10 - 0xa
      13'h1A4E: dout <= 8'b01001010; // 6734 :  74 - 0x4a
      13'h1A4F: dout <= 8'b01100000; // 6735 :  96 - 0x60
      13'h1A50: dout <= 8'b11000000; // 6736 : 192 - 0xc0 -- Background 0xa5
      13'h1A51: dout <= 8'b11000111; // 6737 : 199 - 0xc7
      13'h1A52: dout <= 8'b01101111; // 6738 : 111 - 0x6f
      13'h1A53: dout <= 8'b01100111; // 6739 : 103 - 0x67
      13'h1A54: dout <= 8'b01100011; // 6740 :  99 - 0x63
      13'h1A55: dout <= 8'b00110000; // 6741 :  48 - 0x30
      13'h1A56: dout <= 8'b00011000; // 6742 :  24 - 0x18
      13'h1A57: dout <= 8'b00000111; // 6743 :   7 - 0x7
      13'h1A58: dout <= 8'b01111111; // 6744 : 127 - 0x7f
      13'h1A59: dout <= 8'b01111000; // 6745 : 120 - 0x78
      13'h1A5A: dout <= 8'b00110111; // 6746 :  55 - 0x37
      13'h1A5B: dout <= 8'b00111011; // 6747 :  59 - 0x3b
      13'h1A5C: dout <= 8'b00111100; // 6748 :  60 - 0x3c
      13'h1A5D: dout <= 8'b00011111; // 6749 :  31 - 0x1f
      13'h1A5E: dout <= 8'b00000111; // 6750 :   7 - 0x7
      13'h1A5F: dout <= 8'b00000000; // 6751 :   0 - 0x0
      13'h1A60: dout <= 8'b00000000; // 6752 :   0 - 0x0 -- Background 0xa6
      13'h1A61: dout <= 8'b11110000; // 6753 : 240 - 0xf0
      13'h1A62: dout <= 8'b11111000; // 6754 : 248 - 0xf8
      13'h1A63: dout <= 8'b10001100; // 6755 : 140 - 0x8c
      13'h1A64: dout <= 8'b11111100; // 6756 : 252 - 0xfc
      13'h1A65: dout <= 8'b11111110; // 6757 : 254 - 0xfe
      13'h1A66: dout <= 8'b11111101; // 6758 : 253 - 0xfd
      13'h1A67: dout <= 8'b11111001; // 6759 : 249 - 0xf9
      13'h1A68: dout <= 8'b00000000; // 6760 :   0 - 0x0
      13'h1A69: dout <= 8'b00000000; // 6761 :   0 - 0x0
      13'h1A6A: dout <= 8'b00000000; // 6762 :   0 - 0x0
      13'h1A6B: dout <= 8'b01110000; // 6763 : 112 - 0x70
      13'h1A6C: dout <= 8'b00000000; // 6764 :   0 - 0x0
      13'h1A6D: dout <= 8'b01010000; // 6765 :  80 - 0x50
      13'h1A6E: dout <= 8'b01010010; // 6766 :  82 - 0x52
      13'h1A6F: dout <= 8'b00000110; // 6767 :   6 - 0x6
      13'h1A70: dout <= 8'b00000011; // 6768 :   3 - 0x3 -- Background 0xa7
      13'h1A71: dout <= 8'b11100101; // 6769 : 229 - 0xe5
      13'h1A72: dout <= 8'b11110010; // 6770 : 242 - 0xf2
      13'h1A73: dout <= 8'b11100110; // 6771 : 230 - 0xe6
      13'h1A74: dout <= 8'b11001010; // 6772 : 202 - 0xca
      13'h1A75: dout <= 8'b00010100; // 6773 :  20 - 0x14
      13'h1A76: dout <= 8'b00111000; // 6774 :  56 - 0x38
      13'h1A77: dout <= 8'b11100000; // 6775 : 224 - 0xe0
      13'h1A78: dout <= 8'b11111100; // 6776 : 252 - 0xfc
      13'h1A79: dout <= 8'b00011010; // 6777 :  26 - 0x1a
      13'h1A7A: dout <= 8'b11101100; // 6778 : 236 - 0xec
      13'h1A7B: dout <= 8'b11011000; // 6779 : 216 - 0xd8
      13'h1A7C: dout <= 8'b00110100; // 6780 :  52 - 0x34
      13'h1A7D: dout <= 8'b11101000; // 6781 : 232 - 0xe8
      13'h1A7E: dout <= 8'b11000000; // 6782 : 192 - 0xc0
      13'h1A7F: dout <= 8'b00000000; // 6783 :   0 - 0x0
      13'h1A80: dout <= 8'b00000000; // 6784 :   0 - 0x0 -- Background 0xa8
      13'h1A81: dout <= 8'b00001111; // 6785 :  15 - 0xf
      13'h1A82: dout <= 8'b00011111; // 6786 :  31 - 0x1f
      13'h1A83: dout <= 8'b00110001; // 6787 :  49 - 0x31
      13'h1A84: dout <= 8'b00111111; // 6788 :  63 - 0x3f
      13'h1A85: dout <= 8'b01111111; // 6789 : 127 - 0x7f
      13'h1A86: dout <= 8'b11111111; // 6790 : 255 - 0xff
      13'h1A87: dout <= 8'b11011111; // 6791 : 223 - 0xdf
      13'h1A88: dout <= 8'b00000000; // 6792 :   0 - 0x0
      13'h1A89: dout <= 8'b00000000; // 6793 :   0 - 0x0
      13'h1A8A: dout <= 8'b00000000; // 6794 :   0 - 0x0
      13'h1A8B: dout <= 8'b00001110; // 6795 :  14 - 0xe
      13'h1A8C: dout <= 8'b00000000; // 6796 :   0 - 0x0
      13'h1A8D: dout <= 8'b00001110; // 6797 :  14 - 0xe
      13'h1A8E: dout <= 8'b01001010; // 6798 :  74 - 0x4a
      13'h1A8F: dout <= 8'b01100000; // 6799 :  96 - 0x60
      13'h1A90: dout <= 8'b11000000; // 6800 : 192 - 0xc0 -- Background 0xa9
      13'h1A91: dout <= 8'b11000011; // 6801 : 195 - 0xc3
      13'h1A92: dout <= 8'b11000111; // 6802 : 199 - 0xc7
      13'h1A93: dout <= 8'b11001111; // 6803 : 207 - 0xcf
      13'h1A94: dout <= 8'b11000111; // 6804 : 199 - 0xc7
      13'h1A95: dout <= 8'b11000000; // 6805 : 192 - 0xc0
      13'h1A96: dout <= 8'b11100000; // 6806 : 224 - 0xe0
      13'h1A97: dout <= 8'b11111111; // 6807 : 255 - 0xff
      13'h1A98: dout <= 8'b01111111; // 6808 : 127 - 0x7f
      13'h1A99: dout <= 8'b01111100; // 6809 : 124 - 0x7c
      13'h1A9A: dout <= 8'b01111011; // 6810 : 123 - 0x7b
      13'h1A9B: dout <= 8'b01110111; // 6811 : 119 - 0x77
      13'h1A9C: dout <= 8'b01111000; // 6812 : 120 - 0x78
      13'h1A9D: dout <= 8'b01111111; // 6813 : 127 - 0x7f
      13'h1A9E: dout <= 8'b01111111; // 6814 : 127 - 0x7f
      13'h1A9F: dout <= 8'b00000000; // 6815 :   0 - 0x0
      13'h1AA0: dout <= 8'b00000000; // 6816 :   0 - 0x0 -- Background 0xaa
      13'h1AA1: dout <= 8'b11110000; // 6817 : 240 - 0xf0
      13'h1AA2: dout <= 8'b11111000; // 6818 : 248 - 0xf8
      13'h1AA3: dout <= 8'b10001100; // 6819 : 140 - 0x8c
      13'h1AA4: dout <= 8'b11111100; // 6820 : 252 - 0xfc
      13'h1AA5: dout <= 8'b11111110; // 6821 : 254 - 0xfe
      13'h1AA6: dout <= 8'b11111101; // 6822 : 253 - 0xfd
      13'h1AA7: dout <= 8'b11111001; // 6823 : 249 - 0xf9
      13'h1AA8: dout <= 8'b00000000; // 6824 :   0 - 0x0
      13'h1AA9: dout <= 8'b00000000; // 6825 :   0 - 0x0
      13'h1AAA: dout <= 8'b00000000; // 6826 :   0 - 0x0
      13'h1AAB: dout <= 8'b01110000; // 6827 : 112 - 0x70
      13'h1AAC: dout <= 8'b00000000; // 6828 :   0 - 0x0
      13'h1AAD: dout <= 8'b01110000; // 6829 : 112 - 0x70
      13'h1AAE: dout <= 8'b01010010; // 6830 :  82 - 0x52
      13'h1AAF: dout <= 8'b00000110; // 6831 :   6 - 0x6
      13'h1AB0: dout <= 8'b00000011; // 6832 :   3 - 0x3 -- Background 0xab
      13'h1AB1: dout <= 8'b11000101; // 6833 : 197 - 0xc5
      13'h1AB2: dout <= 8'b11100011; // 6834 : 227 - 0xe3
      13'h1AB3: dout <= 8'b11110101; // 6835 : 245 - 0xf5
      13'h1AB4: dout <= 8'b11100011; // 6836 : 227 - 0xe3
      13'h1AB5: dout <= 8'b00000101; // 6837 :   5 - 0x5
      13'h1AB6: dout <= 8'b00001011; // 6838 :  11 - 0xb
      13'h1AB7: dout <= 8'b11111111; // 6839 : 255 - 0xff
      13'h1AB8: dout <= 8'b11111100; // 6840 : 252 - 0xfc
      13'h1AB9: dout <= 8'b00111010; // 6841 :  58 - 0x3a
      13'h1ABA: dout <= 8'b11011100; // 6842 : 220 - 0xdc
      13'h1ABB: dout <= 8'b11101010; // 6843 : 234 - 0xea
      13'h1ABC: dout <= 8'b00011100; // 6844 :  28 - 0x1c
      13'h1ABD: dout <= 8'b11111010; // 6845 : 250 - 0xfa
      13'h1ABE: dout <= 8'b11110100; // 6846 : 244 - 0xf4
      13'h1ABF: dout <= 8'b00000000; // 6847 :   0 - 0x0
      13'h1AC0: dout <= 8'b10000011; // 6848 : 131 - 0x83 -- Background 0xac
      13'h1AC1: dout <= 8'b10001100; // 6849 : 140 - 0x8c
      13'h1AC2: dout <= 8'b10010000; // 6850 : 144 - 0x90
      13'h1AC3: dout <= 8'b10010000; // 6851 : 144 - 0x90
      13'h1AC4: dout <= 8'b11100000; // 6852 : 224 - 0xe0
      13'h1AC5: dout <= 8'b10100000; // 6853 : 160 - 0xa0
      13'h1AC6: dout <= 8'b10101111; // 6854 : 175 - 0xaf
      13'h1AC7: dout <= 8'b01101111; // 6855 : 111 - 0x6f
      13'h1AC8: dout <= 8'b00000000; // 6856 :   0 - 0x0
      13'h1AC9: dout <= 8'b00000011; // 6857 :   3 - 0x3
      13'h1ACA: dout <= 8'b00001111; // 6858 :  15 - 0xf
      13'h1ACB: dout <= 8'b00001111; // 6859 :  15 - 0xf
      13'h1ACC: dout <= 8'b00011111; // 6860 :  31 - 0x1f
      13'h1ACD: dout <= 8'b01011111; // 6861 :  95 - 0x5f
      13'h1ACE: dout <= 8'b01010000; // 6862 :  80 - 0x50
      13'h1ACF: dout <= 8'b00010000; // 6863 :  16 - 0x10
      13'h1AD0: dout <= 8'b11111011; // 6864 : 251 - 0xfb -- Background 0xad
      13'h1AD1: dout <= 8'b00000101; // 6865 :   5 - 0x5
      13'h1AD2: dout <= 8'b00000101; // 6866 :   5 - 0x5
      13'h1AD3: dout <= 8'b00000101; // 6867 :   5 - 0x5
      13'h1AD4: dout <= 8'b01000101; // 6868 :  69 - 0x45
      13'h1AD5: dout <= 8'b01100101; // 6869 : 101 - 0x65
      13'h1AD6: dout <= 8'b11110101; // 6870 : 245 - 0xf5
      13'h1AD7: dout <= 8'b11111101; // 6871 : 253 - 0xfd
      13'h1AD8: dout <= 8'b00000000; // 6872 :   0 - 0x0
      13'h1AD9: dout <= 8'b11111010; // 6873 : 250 - 0xfa
      13'h1ADA: dout <= 8'b11111010; // 6874 : 250 - 0xfa
      13'h1ADB: dout <= 8'b11111010; // 6875 : 250 - 0xfa
      13'h1ADC: dout <= 8'b10111010; // 6876 : 186 - 0xba
      13'h1ADD: dout <= 8'b10011010; // 6877 : 154 - 0x9a
      13'h1ADE: dout <= 8'b00001010; // 6878 :  10 - 0xa
      13'h1ADF: dout <= 8'b00000010; // 6879 :   2 - 0x2
      13'h1AE0: dout <= 8'b10000011; // 6880 : 131 - 0x83 -- Background 0xae
      13'h1AE1: dout <= 8'b10001100; // 6881 : 140 - 0x8c
      13'h1AE2: dout <= 8'b10010000; // 6882 : 144 - 0x90
      13'h1AE3: dout <= 8'b10010000; // 6883 : 144 - 0x90
      13'h1AE4: dout <= 8'b11100000; // 6884 : 224 - 0xe0
      13'h1AE5: dout <= 8'b10100000; // 6885 : 160 - 0xa0
      13'h1AE6: dout <= 8'b10101111; // 6886 : 175 - 0xaf
      13'h1AE7: dout <= 8'b01101111; // 6887 : 111 - 0x6f
      13'h1AE8: dout <= 8'b00000000; // 6888 :   0 - 0x0
      13'h1AE9: dout <= 8'b00000011; // 6889 :   3 - 0x3
      13'h1AEA: dout <= 8'b00001111; // 6890 :  15 - 0xf
      13'h1AEB: dout <= 8'b00001111; // 6891 :  15 - 0xf
      13'h1AEC: dout <= 8'b00011111; // 6892 :  31 - 0x1f
      13'h1AED: dout <= 8'b01011111; // 6893 :  95 - 0x5f
      13'h1AEE: dout <= 8'b01010000; // 6894 :  80 - 0x50
      13'h1AEF: dout <= 8'b00010111; // 6895 :  23 - 0x17
      13'h1AF0: dout <= 8'b11111011; // 6896 : 251 - 0xfb -- Background 0xaf
      13'h1AF1: dout <= 8'b00000101; // 6897 :   5 - 0x5
      13'h1AF2: dout <= 8'b00000101; // 6898 :   5 - 0x5
      13'h1AF3: dout <= 8'b00000101; // 6899 :   5 - 0x5
      13'h1AF4: dout <= 8'b11000101; // 6900 : 197 - 0xc5
      13'h1AF5: dout <= 8'b11100101; // 6901 : 229 - 0xe5
      13'h1AF6: dout <= 8'b11110101; // 6902 : 245 - 0xf5
      13'h1AF7: dout <= 8'b11111101; // 6903 : 253 - 0xfd
      13'h1AF8: dout <= 8'b00000000; // 6904 :   0 - 0x0
      13'h1AF9: dout <= 8'b11111010; // 6905 : 250 - 0xfa
      13'h1AFA: dout <= 8'b11111010; // 6906 : 250 - 0xfa
      13'h1AFB: dout <= 8'b11111010; // 6907 : 250 - 0xfa
      13'h1AFC: dout <= 8'b00111010; // 6908 :  58 - 0x3a
      13'h1AFD: dout <= 8'b01011010; // 6909 :  90 - 0x5a
      13'h1AFE: dout <= 8'b01101010; // 6910 : 106 - 0x6a
      13'h1AFF: dout <= 8'b11110010; // 6911 : 242 - 0xf2
      13'h1B00: dout <= 8'b00000000; // 6912 :   0 - 0x0 -- Background 0xb0
      13'h1B01: dout <= 8'b00000011; // 6913 :   3 - 0x3
      13'h1B02: dout <= 8'b00001111; // 6914 :  15 - 0xf
      13'h1B03: dout <= 8'b00111111; // 6915 :  63 - 0x3f
      13'h1B04: dout <= 8'b01111111; // 6916 : 127 - 0x7f
      13'h1B05: dout <= 8'b01111111; // 6917 : 127 - 0x7f
      13'h1B06: dout <= 8'b11111111; // 6918 : 255 - 0xff
      13'h1B07: dout <= 8'b11111111; // 6919 : 255 - 0xff
      13'h1B08: dout <= 8'b00000000; // 6920 :   0 - 0x0
      13'h1B09: dout <= 8'b00000000; // 6921 :   0 - 0x0
      13'h1B0A: dout <= 8'b00000011; // 6922 :   3 - 0x3
      13'h1B0B: dout <= 8'b00001111; // 6923 :  15 - 0xf
      13'h1B0C: dout <= 8'b00111011; // 6924 :  59 - 0x3b
      13'h1B0D: dout <= 8'b00111111; // 6925 :  63 - 0x3f
      13'h1B0E: dout <= 8'b01101111; // 6926 : 111 - 0x6f
      13'h1B0F: dout <= 8'b01111101; // 6927 : 125 - 0x7d
      13'h1B10: dout <= 8'b11111111; // 6928 : 255 - 0xff -- Background 0xb1
      13'h1B11: dout <= 8'b10001111; // 6929 : 143 - 0x8f
      13'h1B12: dout <= 8'b10000000; // 6930 : 128 - 0x80
      13'h1B13: dout <= 8'b11110000; // 6931 : 240 - 0xf0
      13'h1B14: dout <= 8'b11111111; // 6932 : 255 - 0xff
      13'h1B15: dout <= 8'b11111111; // 6933 : 255 - 0xff
      13'h1B16: dout <= 8'b01111111; // 6934 : 127 - 0x7f
      13'h1B17: dout <= 8'b00001111; // 6935 :  15 - 0xf
      13'h1B18: dout <= 8'b00001111; // 6936 :  15 - 0xf
      13'h1B19: dout <= 8'b01110000; // 6937 : 112 - 0x70
      13'h1B1A: dout <= 8'b01111111; // 6938 : 127 - 0x7f
      13'h1B1B: dout <= 8'b00001111; // 6939 :  15 - 0xf
      13'h1B1C: dout <= 8'b01110000; // 6940 : 112 - 0x70
      13'h1B1D: dout <= 8'b01111111; // 6941 : 127 - 0x7f
      13'h1B1E: dout <= 8'b00001111; // 6942 :  15 - 0xf
      13'h1B1F: dout <= 8'b00000000; // 6943 :   0 - 0x0
      13'h1B20: dout <= 8'b00000000; // 6944 :   0 - 0x0 -- Background 0xb2
      13'h1B21: dout <= 8'b11000000; // 6945 : 192 - 0xc0
      13'h1B22: dout <= 8'b11110000; // 6946 : 240 - 0xf0
      13'h1B23: dout <= 8'b11111100; // 6947 : 252 - 0xfc
      13'h1B24: dout <= 8'b11111110; // 6948 : 254 - 0xfe
      13'h1B25: dout <= 8'b11111110; // 6949 : 254 - 0xfe
      13'h1B26: dout <= 8'b11111111; // 6950 : 255 - 0xff
      13'h1B27: dout <= 8'b11111111; // 6951 : 255 - 0xff
      13'h1B28: dout <= 8'b00000000; // 6952 :   0 - 0x0
      13'h1B29: dout <= 8'b00000000; // 6953 :   0 - 0x0
      13'h1B2A: dout <= 8'b11000000; // 6954 : 192 - 0xc0
      13'h1B2B: dout <= 8'b11110000; // 6955 : 240 - 0xf0
      13'h1B2C: dout <= 8'b10111100; // 6956 : 188 - 0xbc
      13'h1B2D: dout <= 8'b11110100; // 6957 : 244 - 0xf4
      13'h1B2E: dout <= 8'b11111110; // 6958 : 254 - 0xfe
      13'h1B2F: dout <= 8'b11011110; // 6959 : 222 - 0xde
      13'h1B30: dout <= 8'b11111111; // 6960 : 255 - 0xff -- Background 0xb3
      13'h1B31: dout <= 8'b11110001; // 6961 : 241 - 0xf1
      13'h1B32: dout <= 8'b00000001; // 6962 :   1 - 0x1
      13'h1B33: dout <= 8'b00001111; // 6963 :  15 - 0xf
      13'h1B34: dout <= 8'b11111111; // 6964 : 255 - 0xff
      13'h1B35: dout <= 8'b11111111; // 6965 : 255 - 0xff
      13'h1B36: dout <= 8'b11111110; // 6966 : 254 - 0xfe
      13'h1B37: dout <= 8'b11110000; // 6967 : 240 - 0xf0
      13'h1B38: dout <= 8'b11110000; // 6968 : 240 - 0xf0
      13'h1B39: dout <= 8'b00001110; // 6969 :  14 - 0xe
      13'h1B3A: dout <= 8'b11111110; // 6970 : 254 - 0xfe
      13'h1B3B: dout <= 8'b11110000; // 6971 : 240 - 0xf0
      13'h1B3C: dout <= 8'b00001110; // 6972 :  14 - 0xe
      13'h1B3D: dout <= 8'b11111110; // 6973 : 254 - 0xfe
      13'h1B3E: dout <= 8'b11110000; // 6974 : 240 - 0xf0
      13'h1B3F: dout <= 8'b00000000; // 6975 :   0 - 0x0
      13'h1B40: dout <= 8'b00000000; // 6976 :   0 - 0x0 -- Background 0xb4
      13'h1B41: dout <= 8'b00000011; // 6977 :   3 - 0x3
      13'h1B42: dout <= 8'b00001110; // 6978 :  14 - 0xe
      13'h1B43: dout <= 8'b00110101; // 6979 :  53 - 0x35
      13'h1B44: dout <= 8'b01101110; // 6980 : 110 - 0x6e
      13'h1B45: dout <= 8'b01010101; // 6981 :  85 - 0x55
      13'h1B46: dout <= 8'b10111010; // 6982 : 186 - 0xba
      13'h1B47: dout <= 8'b11010111; // 6983 : 215 - 0xd7
      13'h1B48: dout <= 8'b00000000; // 6984 :   0 - 0x0
      13'h1B49: dout <= 8'b00000000; // 6985 :   0 - 0x0
      13'h1B4A: dout <= 8'b00000011; // 6986 :   3 - 0x3
      13'h1B4B: dout <= 8'b00001111; // 6987 :  15 - 0xf
      13'h1B4C: dout <= 8'b00111011; // 6988 :  59 - 0x3b
      13'h1B4D: dout <= 8'b00111111; // 6989 :  63 - 0x3f
      13'h1B4E: dout <= 8'b01101111; // 6990 : 111 - 0x6f
      13'h1B4F: dout <= 8'b01111101; // 6991 : 125 - 0x7d
      13'h1B50: dout <= 8'b11111010; // 6992 : 250 - 0xfa -- Background 0xb5
      13'h1B51: dout <= 8'b10001111; // 6993 : 143 - 0x8f
      13'h1B52: dout <= 8'b10000000; // 6994 : 128 - 0x80
      13'h1B53: dout <= 8'b11110000; // 6995 : 240 - 0xf0
      13'h1B54: dout <= 8'b10101111; // 6996 : 175 - 0xaf
      13'h1B55: dout <= 8'b11010101; // 6997 : 213 - 0xd5
      13'h1B56: dout <= 8'b01111010; // 6998 : 122 - 0x7a
      13'h1B57: dout <= 8'b00001111; // 6999 :  15 - 0xf
      13'h1B58: dout <= 8'b00001111; // 7000 :  15 - 0xf
      13'h1B59: dout <= 8'b01110000; // 7001 : 112 - 0x70
      13'h1B5A: dout <= 8'b01111111; // 7002 : 127 - 0x7f
      13'h1B5B: dout <= 8'b00001111; // 7003 :  15 - 0xf
      13'h1B5C: dout <= 8'b01110000; // 7004 : 112 - 0x70
      13'h1B5D: dout <= 8'b01111111; // 7005 : 127 - 0x7f
      13'h1B5E: dout <= 8'b00001111; // 7006 :  15 - 0xf
      13'h1B5F: dout <= 8'b00000000; // 7007 :   0 - 0x0
      13'h1B60: dout <= 8'b00000000; // 7008 :   0 - 0x0 -- Background 0xb6
      13'h1B61: dout <= 8'b11000000; // 7009 : 192 - 0xc0
      13'h1B62: dout <= 8'b10110000; // 7010 : 176 - 0xb0
      13'h1B63: dout <= 8'b01011100; // 7011 :  92 - 0x5c
      13'h1B64: dout <= 8'b11101010; // 7012 : 234 - 0xea
      13'h1B65: dout <= 8'b01011110; // 7013 :  94 - 0x5e
      13'h1B66: dout <= 8'b10101011; // 7014 : 171 - 0xab
      13'h1B67: dout <= 8'b01110101; // 7015 : 117 - 0x75
      13'h1B68: dout <= 8'b00000000; // 7016 :   0 - 0x0
      13'h1B69: dout <= 8'b00000000; // 7017 :   0 - 0x0
      13'h1B6A: dout <= 8'b11000000; // 7018 : 192 - 0xc0
      13'h1B6B: dout <= 8'b11110000; // 7019 : 240 - 0xf0
      13'h1B6C: dout <= 8'b10111100; // 7020 : 188 - 0xbc
      13'h1B6D: dout <= 8'b11110100; // 7021 : 244 - 0xf4
      13'h1B6E: dout <= 8'b11111110; // 7022 : 254 - 0xfe
      13'h1B6F: dout <= 8'b11011110; // 7023 : 222 - 0xde
      13'h1B70: dout <= 8'b10101111; // 7024 : 175 - 0xaf -- Background 0xb7
      13'h1B71: dout <= 8'b11110001; // 7025 : 241 - 0xf1
      13'h1B72: dout <= 8'b00000001; // 7026 :   1 - 0x1
      13'h1B73: dout <= 8'b00001111; // 7027 :  15 - 0xf
      13'h1B74: dout <= 8'b11111011; // 7028 : 251 - 0xfb
      13'h1B75: dout <= 8'b01010101; // 7029 :  85 - 0x55
      13'h1B76: dout <= 8'b10101110; // 7030 : 174 - 0xae
      13'h1B77: dout <= 8'b11110000; // 7031 : 240 - 0xf0
      13'h1B78: dout <= 8'b11110000; // 7032 : 240 - 0xf0
      13'h1B79: dout <= 8'b00001110; // 7033 :  14 - 0xe
      13'h1B7A: dout <= 8'b11111110; // 7034 : 254 - 0xfe
      13'h1B7B: dout <= 8'b11110000; // 7035 : 240 - 0xf0
      13'h1B7C: dout <= 8'b00001110; // 7036 :  14 - 0xe
      13'h1B7D: dout <= 8'b11111110; // 7037 : 254 - 0xfe
      13'h1B7E: dout <= 8'b11110000; // 7038 : 240 - 0xf0
      13'h1B7F: dout <= 8'b00000000; // 7039 :   0 - 0x0
      13'h1B80: dout <= 8'b00000000; // 7040 :   0 - 0x0 -- Background 0xb8
      13'h1B81: dout <= 8'b00000011; // 7041 :   3 - 0x3
      13'h1B82: dout <= 8'b00001100; // 7042 :  12 - 0xc
      13'h1B83: dout <= 8'b00110000; // 7043 :  48 - 0x30
      13'h1B84: dout <= 8'b01000100; // 7044 :  68 - 0x44
      13'h1B85: dout <= 8'b01000000; // 7045 :  64 - 0x40
      13'h1B86: dout <= 8'b10010000; // 7046 : 144 - 0x90
      13'h1B87: dout <= 8'b10000010; // 7047 : 130 - 0x82
      13'h1B88: dout <= 8'b00000000; // 7048 :   0 - 0x0
      13'h1B89: dout <= 8'b00000000; // 7049 :   0 - 0x0
      13'h1B8A: dout <= 8'b00000011; // 7050 :   3 - 0x3
      13'h1B8B: dout <= 8'b00001111; // 7051 :  15 - 0xf
      13'h1B8C: dout <= 8'b00111011; // 7052 :  59 - 0x3b
      13'h1B8D: dout <= 8'b00111111; // 7053 :  63 - 0x3f
      13'h1B8E: dout <= 8'b01101111; // 7054 : 111 - 0x6f
      13'h1B8F: dout <= 8'b01111101; // 7055 : 125 - 0x7d
      13'h1B90: dout <= 8'b11110000; // 7056 : 240 - 0xf0 -- Background 0xb9
      13'h1B91: dout <= 8'b11111111; // 7057 : 255 - 0xff
      13'h1B92: dout <= 8'b11111111; // 7058 : 255 - 0xff
      13'h1B93: dout <= 8'b11111111; // 7059 : 255 - 0xff
      13'h1B94: dout <= 8'b10001111; // 7060 : 143 - 0x8f
      13'h1B95: dout <= 8'b10000000; // 7061 : 128 - 0x80
      13'h1B96: dout <= 8'b01110000; // 7062 : 112 - 0x70
      13'h1B97: dout <= 8'b00001111; // 7063 :  15 - 0xf
      13'h1B98: dout <= 8'b00001111; // 7064 :  15 - 0xf
      13'h1B99: dout <= 8'b00100000; // 7065 :  32 - 0x20
      13'h1B9A: dout <= 8'b01010101; // 7066 :  85 - 0x55
      13'h1B9B: dout <= 8'b00001010; // 7067 :  10 - 0xa
      13'h1B9C: dout <= 8'b01110000; // 7068 : 112 - 0x70
      13'h1B9D: dout <= 8'b01111111; // 7069 : 127 - 0x7f
      13'h1B9E: dout <= 8'b00001111; // 7070 :  15 - 0xf
      13'h1B9F: dout <= 8'b00000000; // 7071 :   0 - 0x0
      13'h1BA0: dout <= 8'b00000000; // 7072 :   0 - 0x0 -- Background 0xba
      13'h1BA1: dout <= 8'b11000000; // 7073 : 192 - 0xc0
      13'h1BA2: dout <= 8'b00110000; // 7074 :  48 - 0x30
      13'h1BA3: dout <= 8'b00001100; // 7075 :  12 - 0xc
      13'h1BA4: dout <= 8'b01000010; // 7076 :  66 - 0x42
      13'h1BA5: dout <= 8'b00001010; // 7077 :  10 - 0xa
      13'h1BA6: dout <= 8'b00000001; // 7078 :   1 - 0x1
      13'h1BA7: dout <= 8'b00100001; // 7079 :  33 - 0x21
      13'h1BA8: dout <= 8'b00000000; // 7080 :   0 - 0x0
      13'h1BA9: dout <= 8'b00000000; // 7081 :   0 - 0x0
      13'h1BAA: dout <= 8'b11000000; // 7082 : 192 - 0xc0
      13'h1BAB: dout <= 8'b11110000; // 7083 : 240 - 0xf0
      13'h1BAC: dout <= 8'b10111100; // 7084 : 188 - 0xbc
      13'h1BAD: dout <= 8'b11110100; // 7085 : 244 - 0xf4
      13'h1BAE: dout <= 8'b11111110; // 7086 : 254 - 0xfe
      13'h1BAF: dout <= 8'b11011110; // 7087 : 222 - 0xde
      13'h1BB0: dout <= 8'b00001111; // 7088 :  15 - 0xf -- Background 0xbb
      13'h1BB1: dout <= 8'b11111111; // 7089 : 255 - 0xff
      13'h1BB2: dout <= 8'b11111111; // 7090 : 255 - 0xff
      13'h1BB3: dout <= 8'b11111111; // 7091 : 255 - 0xff
      13'h1BB4: dout <= 8'b11110001; // 7092 : 241 - 0xf1
      13'h1BB5: dout <= 8'b00000001; // 7093 :   1 - 0x1
      13'h1BB6: dout <= 8'b00001110; // 7094 :  14 - 0xe
      13'h1BB7: dout <= 8'b11110000; // 7095 : 240 - 0xf0
      13'h1BB8: dout <= 8'b11110000; // 7096 : 240 - 0xf0
      13'h1BB9: dout <= 8'b00001010; // 7097 :  10 - 0xa
      13'h1BBA: dout <= 8'b01010100; // 7098 :  84 - 0x54
      13'h1BBB: dout <= 8'b10100000; // 7099 : 160 - 0xa0
      13'h1BBC: dout <= 8'b00001110; // 7100 :  14 - 0xe
      13'h1BBD: dout <= 8'b11111110; // 7101 : 254 - 0xfe
      13'h1BBE: dout <= 8'b11110000; // 7102 : 240 - 0xf0
      13'h1BBF: dout <= 8'b00000000; // 7103 :   0 - 0x0
      13'h1BC0: dout <= 8'b11110011; // 7104 : 243 - 0xf3 -- Background 0xbc
      13'h1BC1: dout <= 8'b11111111; // 7105 : 255 - 0xff
      13'h1BC2: dout <= 8'b11000100; // 7106 : 196 - 0xc4
      13'h1BC3: dout <= 8'b11000000; // 7107 : 192 - 0xc0
      13'h1BC4: dout <= 8'b01000000; // 7108 :  64 - 0x40
      13'h1BC5: dout <= 8'b01100011; // 7109 :  99 - 0x63
      13'h1BC6: dout <= 8'b11000111; // 7110 : 199 - 0xc7
      13'h1BC7: dout <= 8'b11000110; // 7111 : 198 - 0xc6
      13'h1BC8: dout <= 8'b00000000; // 7112 :   0 - 0x0
      13'h1BC9: dout <= 8'b01110011; // 7113 : 115 - 0x73
      13'h1BCA: dout <= 8'b01111011; // 7114 : 123 - 0x7b
      13'h1BCB: dout <= 8'b01111111; // 7115 : 127 - 0x7f
      13'h1BCC: dout <= 8'b00111111; // 7116 :  63 - 0x3f
      13'h1BCD: dout <= 8'b00011100; // 7117 :  28 - 0x1c
      13'h1BCE: dout <= 8'b01111011; // 7118 : 123 - 0x7b
      13'h1BCF: dout <= 8'b01111011; // 7119 : 123 - 0x7b
      13'h1BD0: dout <= 8'b11000110; // 7120 : 198 - 0xc6 -- Background 0xbd
      13'h1BD1: dout <= 8'b11000110; // 7121 : 198 - 0xc6
      13'h1BD2: dout <= 8'b01100011; // 7122 :  99 - 0x63
      13'h1BD3: dout <= 8'b01000000; // 7123 :  64 - 0x40
      13'h1BD4: dout <= 8'b11000000; // 7124 : 192 - 0xc0
      13'h1BD5: dout <= 8'b11000100; // 7125 : 196 - 0xc4
      13'h1BD6: dout <= 8'b11001100; // 7126 : 204 - 0xcc
      13'h1BD7: dout <= 8'b11110011; // 7127 : 243 - 0xf3
      13'h1BD8: dout <= 8'b01111011; // 7128 : 123 - 0x7b
      13'h1BD9: dout <= 8'b01111011; // 7129 : 123 - 0x7b
      13'h1BDA: dout <= 8'b00011100; // 7130 :  28 - 0x1c
      13'h1BDB: dout <= 8'b00111111; // 7131 :  63 - 0x3f
      13'h1BDC: dout <= 8'b01111111; // 7132 : 127 - 0x7f
      13'h1BDD: dout <= 8'b01111011; // 7133 : 123 - 0x7b
      13'h1BDE: dout <= 8'b01110011; // 7134 : 115 - 0x73
      13'h1BDF: dout <= 8'b00000000; // 7135 :   0 - 0x0
      13'h1BE0: dout <= 8'b11001111; // 7136 : 207 - 0xcf -- Background 0xbe
      13'h1BE1: dout <= 8'b11111111; // 7137 : 255 - 0xff
      13'h1BE2: dout <= 8'b00100001; // 7138 :  33 - 0x21
      13'h1BE3: dout <= 8'b00000001; // 7139 :   1 - 0x1
      13'h1BE4: dout <= 8'b00000010; // 7140 :   2 - 0x2
      13'h1BE5: dout <= 8'b11000110; // 7141 : 198 - 0xc6
      13'h1BE6: dout <= 8'b11100001; // 7142 : 225 - 0xe1
      13'h1BE7: dout <= 8'b00100001; // 7143 :  33 - 0x21
      13'h1BE8: dout <= 8'b00000000; // 7144 :   0 - 0x0
      13'h1BE9: dout <= 8'b11001110; // 7145 : 206 - 0xce
      13'h1BEA: dout <= 8'b11011110; // 7146 : 222 - 0xde
      13'h1BEB: dout <= 8'b11111110; // 7147 : 254 - 0xfe
      13'h1BEC: dout <= 8'b11111100; // 7148 : 252 - 0xfc
      13'h1BED: dout <= 8'b00111000; // 7149 :  56 - 0x38
      13'h1BEE: dout <= 8'b11011110; // 7150 : 222 - 0xde
      13'h1BEF: dout <= 8'b11011110; // 7151 : 222 - 0xde
      13'h1BF0: dout <= 8'b00100001; // 7152 :  33 - 0x21 -- Background 0xbf
      13'h1BF1: dout <= 8'b00100001; // 7153 :  33 - 0x21
      13'h1BF2: dout <= 8'b11000110; // 7154 : 198 - 0xc6
      13'h1BF3: dout <= 8'b00000010; // 7155 :   2 - 0x2
      13'h1BF4: dout <= 8'b00000001; // 7156 :   1 - 0x1
      13'h1BF5: dout <= 8'b00100001; // 7157 :  33 - 0x21
      13'h1BF6: dout <= 8'b00110001; // 7158 :  49 - 0x31
      13'h1BF7: dout <= 8'b11001111; // 7159 : 207 - 0xcf
      13'h1BF8: dout <= 8'b11011110; // 7160 : 222 - 0xde
      13'h1BF9: dout <= 8'b11011110; // 7161 : 222 - 0xde
      13'h1BFA: dout <= 8'b00111000; // 7162 :  56 - 0x38
      13'h1BFB: dout <= 8'b11111100; // 7163 : 252 - 0xfc
      13'h1BFC: dout <= 8'b11111110; // 7164 : 254 - 0xfe
      13'h1BFD: dout <= 8'b11011110; // 7165 : 222 - 0xde
      13'h1BFE: dout <= 8'b11001110; // 7166 : 206 - 0xce
      13'h1BFF: dout <= 8'b00000000; // 7167 :   0 - 0x0
      13'h1C00: dout <= 8'b00000000; // 7168 :   0 - 0x0 -- Background 0xc0
      13'h1C01: dout <= 8'b01010000; // 7169 :  80 - 0x50
      13'h1C02: dout <= 8'b10110011; // 7170 : 179 - 0xb3
      13'h1C03: dout <= 8'b10010111; // 7171 : 151 - 0x97
      13'h1C04: dout <= 8'b10011111; // 7172 : 159 - 0x9f
      13'h1C05: dout <= 8'b01101111; // 7173 : 111 - 0x6f
      13'h1C06: dout <= 8'b00011111; // 7174 :  31 - 0x1f
      13'h1C07: dout <= 8'b00011111; // 7175 :  31 - 0x1f
      13'h1C08: dout <= 8'b00000000; // 7176 :   0 - 0x0
      13'h1C09: dout <= 8'b00000000; // 7177 :   0 - 0x0
      13'h1C0A: dout <= 8'b01000000; // 7178 :  64 - 0x40
      13'h1C0B: dout <= 8'b01100000; // 7179 :  96 - 0x60
      13'h1C0C: dout <= 8'b01100001; // 7180 :  97 - 0x61
      13'h1C0D: dout <= 8'b00000010; // 7181 :   2 - 0x2
      13'h1C0E: dout <= 8'b00000010; // 7182 :   2 - 0x2
      13'h1C0F: dout <= 8'b00000111; // 7183 :   7 - 0x7
      13'h1C10: dout <= 8'b00011111; // 7184 :  31 - 0x1f -- Background 0xc1
      13'h1C11: dout <= 8'b00011111; // 7185 :  31 - 0x1f
      13'h1C12: dout <= 8'b00001111; // 7186 :  15 - 0xf
      13'h1C13: dout <= 8'b00000111; // 7187 :   7 - 0x7
      13'h1C14: dout <= 8'b00011101; // 7188 :  29 - 0x1d
      13'h1C15: dout <= 8'b00101100; // 7189 :  44 - 0x2c
      13'h1C16: dout <= 8'b01010100; // 7190 :  84 - 0x54
      13'h1C17: dout <= 8'b01111100; // 7191 : 124 - 0x7c
      13'h1C18: dout <= 8'b00000111; // 7192 :   7 - 0x7
      13'h1C19: dout <= 8'b00000100; // 7193 :   4 - 0x4
      13'h1C1A: dout <= 8'b00000111; // 7194 :   7 - 0x7
      13'h1C1B: dout <= 8'b00000001; // 7195 :   1 - 0x1
      13'h1C1C: dout <= 8'b00000000; // 7196 :   0 - 0x0
      13'h1C1D: dout <= 8'b00010000; // 7197 :  16 - 0x10
      13'h1C1E: dout <= 8'b00101000; // 7198 :  40 - 0x28
      13'h1C1F: dout <= 8'b00000000; // 7199 :   0 - 0x0
      13'h1C20: dout <= 8'b00000000; // 7200 :   0 - 0x0 -- Background 0xc2
      13'h1C21: dout <= 8'b00001010; // 7201 :  10 - 0xa
      13'h1C22: dout <= 8'b11001101; // 7202 : 205 - 0xcd
      13'h1C23: dout <= 8'b11101001; // 7203 : 233 - 0xe9
      13'h1C24: dout <= 8'b11111001; // 7204 : 249 - 0xf9
      13'h1C25: dout <= 8'b11110110; // 7205 : 246 - 0xf6
      13'h1C26: dout <= 8'b11110000; // 7206 : 240 - 0xf0
      13'h1C27: dout <= 8'b11111000; // 7207 : 248 - 0xf8
      13'h1C28: dout <= 8'b00000000; // 7208 :   0 - 0x0
      13'h1C29: dout <= 8'b00000000; // 7209 :   0 - 0x0
      13'h1C2A: dout <= 8'b00000010; // 7210 :   2 - 0x2
      13'h1C2B: dout <= 8'b00000110; // 7211 :   6 - 0x6
      13'h1C2C: dout <= 8'b11100110; // 7212 : 230 - 0xe6
      13'h1C2D: dout <= 8'b10100000; // 7213 : 160 - 0xa0
      13'h1C2E: dout <= 8'b10100000; // 7214 : 160 - 0xa0
      13'h1C2F: dout <= 8'b11110000; // 7215 : 240 - 0xf0
      13'h1C30: dout <= 8'b11111000; // 7216 : 248 - 0xf8 -- Background 0xc3
      13'h1C31: dout <= 8'b11111000; // 7217 : 248 - 0xf8
      13'h1C32: dout <= 8'b11110000; // 7218 : 240 - 0xf0
      13'h1C33: dout <= 8'b11000000; // 7219 : 192 - 0xc0
      13'h1C34: dout <= 8'b10111000; // 7220 : 184 - 0xb8
      13'h1C35: dout <= 8'b00110100; // 7221 :  52 - 0x34
      13'h1C36: dout <= 8'b00101010; // 7222 :  42 - 0x2a
      13'h1C37: dout <= 8'b00111110; // 7223 :  62 - 0x3e
      13'h1C38: dout <= 8'b11110000; // 7224 : 240 - 0xf0
      13'h1C39: dout <= 8'b00110000; // 7225 :  48 - 0x30
      13'h1C3A: dout <= 8'b11000000; // 7226 : 192 - 0xc0
      13'h1C3B: dout <= 8'b10000000; // 7227 : 128 - 0x80
      13'h1C3C: dout <= 8'b00000000; // 7228 :   0 - 0x0
      13'h1C3D: dout <= 8'b00001000; // 7229 :   8 - 0x8
      13'h1C3E: dout <= 8'b00010100; // 7230 :  20 - 0x14
      13'h1C3F: dout <= 8'b00000000; // 7231 :   0 - 0x0
      13'h1C40: dout <= 8'b00000101; // 7232 :   5 - 0x5 -- Background 0xc4
      13'h1C41: dout <= 8'b00001010; // 7233 :  10 - 0xa
      13'h1C42: dout <= 8'b00001000; // 7234 :   8 - 0x8
      13'h1C43: dout <= 8'b00001111; // 7235 :  15 - 0xf
      13'h1C44: dout <= 8'b00000001; // 7236 :   1 - 0x1
      13'h1C45: dout <= 8'b00000011; // 7237 :   3 - 0x3
      13'h1C46: dout <= 8'b00000111; // 7238 :   7 - 0x7
      13'h1C47: dout <= 8'b00001111; // 7239 :  15 - 0xf
      13'h1C48: dout <= 8'b00000000; // 7240 :   0 - 0x0
      13'h1C49: dout <= 8'b00000101; // 7241 :   5 - 0x5
      13'h1C4A: dout <= 8'b00000111; // 7242 :   7 - 0x7
      13'h1C4B: dout <= 8'b00000000; // 7243 :   0 - 0x0
      13'h1C4C: dout <= 8'b00000000; // 7244 :   0 - 0x0
      13'h1C4D: dout <= 8'b00000000; // 7245 :   0 - 0x0
      13'h1C4E: dout <= 8'b00000000; // 7246 :   0 - 0x0
      13'h1C4F: dout <= 8'b00000001; // 7247 :   1 - 0x1
      13'h1C50: dout <= 8'b00001111; // 7248 :  15 - 0xf -- Background 0xc5
      13'h1C51: dout <= 8'b11101111; // 7249 : 239 - 0xef
      13'h1C52: dout <= 8'b11011111; // 7250 : 223 - 0xdf
      13'h1C53: dout <= 8'b10101111; // 7251 : 175 - 0xaf
      13'h1C54: dout <= 8'b01100111; // 7252 : 103 - 0x67
      13'h1C55: dout <= 8'b00001101; // 7253 :  13 - 0xd
      13'h1C56: dout <= 8'b00001010; // 7254 :  10 - 0xa
      13'h1C57: dout <= 8'b00000111; // 7255 :   7 - 0x7
      13'h1C58: dout <= 8'b00000010; // 7256 :   2 - 0x2
      13'h1C59: dout <= 8'b00000111; // 7257 :   7 - 0x7
      13'h1C5A: dout <= 8'b00100111; // 7258 :  39 - 0x27
      13'h1C5B: dout <= 8'b01010011; // 7259 :  83 - 0x53
      13'h1C5C: dout <= 8'b00000000; // 7260 :   0 - 0x0
      13'h1C5D: dout <= 8'b00000010; // 7261 :   2 - 0x2
      13'h1C5E: dout <= 8'b00000101; // 7262 :   5 - 0x5
      13'h1C5F: dout <= 8'b00000000; // 7263 :   0 - 0x0
      13'h1C60: dout <= 8'b00000000; // 7264 :   0 - 0x0 -- Background 0xc6
      13'h1C61: dout <= 8'b10000000; // 7265 : 128 - 0x80
      13'h1C62: dout <= 8'b10000000; // 7266 : 128 - 0x80
      13'h1C63: dout <= 8'b11110000; // 7267 : 240 - 0xf0
      13'h1C64: dout <= 8'b11111000; // 7268 : 248 - 0xf8
      13'h1C65: dout <= 8'b11111100; // 7269 : 252 - 0xfc
      13'h1C66: dout <= 8'b11111100; // 7270 : 252 - 0xfc
      13'h1C67: dout <= 8'b11111100; // 7271 : 252 - 0xfc
      13'h1C68: dout <= 8'b00000000; // 7272 :   0 - 0x0
      13'h1C69: dout <= 8'b00000000; // 7273 :   0 - 0x0
      13'h1C6A: dout <= 8'b00000000; // 7274 :   0 - 0x0
      13'h1C6B: dout <= 8'b00000000; // 7275 :   0 - 0x0
      13'h1C6C: dout <= 8'b00000000; // 7276 :   0 - 0x0
      13'h1C6D: dout <= 8'b01100000; // 7277 :  96 - 0x60
      13'h1C6E: dout <= 8'b11011000; // 7278 : 216 - 0xd8
      13'h1C6F: dout <= 8'b10110000; // 7279 : 176 - 0xb0
      13'h1C70: dout <= 8'b11111100; // 7280 : 252 - 0xfc -- Background 0xc7
      13'h1C71: dout <= 8'b11111110; // 7281 : 254 - 0xfe
      13'h1C72: dout <= 8'b11111001; // 7282 : 249 - 0xf9
      13'h1C73: dout <= 8'b11111010; // 7283 : 250 - 0xfa
      13'h1C74: dout <= 8'b11101001; // 7284 : 233 - 0xe9
      13'h1C75: dout <= 8'b00001110; // 7285 :  14 - 0xe
      13'h1C76: dout <= 8'b10000000; // 7286 : 128 - 0x80
      13'h1C77: dout <= 8'b00000000; // 7287 :   0 - 0x0
      13'h1C78: dout <= 8'b11101000; // 7288 : 232 - 0xe8
      13'h1C79: dout <= 8'b01111000; // 7289 : 120 - 0x78
      13'h1C7A: dout <= 8'b10110110; // 7290 : 182 - 0xb6
      13'h1C7B: dout <= 8'b11100100; // 7291 : 228 - 0xe4
      13'h1C7C: dout <= 8'b00000110; // 7292 :   6 - 0x6
      13'h1C7D: dout <= 8'b00000000; // 7293 :   0 - 0x0
      13'h1C7E: dout <= 8'b00000000; // 7294 :   0 - 0x0
      13'h1C7F: dout <= 8'b00000000; // 7295 :   0 - 0x0
      13'h1C80: dout <= 8'b00000000; // 7296 :   0 - 0x0 -- Background 0xc8
      13'h1C81: dout <= 8'b11000000; // 7297 : 192 - 0xc0
      13'h1C82: dout <= 8'b10100000; // 7298 : 160 - 0xa0
      13'h1C83: dout <= 8'b11010011; // 7299 : 211 - 0xd3
      13'h1C84: dout <= 8'b10110111; // 7300 : 183 - 0xb7
      13'h1C85: dout <= 8'b11111111; // 7301 : 255 - 0xff
      13'h1C86: dout <= 8'b00001111; // 7302 :  15 - 0xf
      13'h1C87: dout <= 8'b00011111; // 7303 :  31 - 0x1f
      13'h1C88: dout <= 8'b00000000; // 7304 :   0 - 0x0
      13'h1C89: dout <= 8'b00000000; // 7305 :   0 - 0x0
      13'h1C8A: dout <= 8'b01000000; // 7306 :  64 - 0x40
      13'h1C8B: dout <= 8'b00100000; // 7307 :  32 - 0x20
      13'h1C8C: dout <= 8'b01000000; // 7308 :  64 - 0x40
      13'h1C8D: dout <= 8'b00000111; // 7309 :   7 - 0x7
      13'h1C8E: dout <= 8'b00000101; // 7310 :   5 - 0x5
      13'h1C8F: dout <= 8'b00001101; // 7311 :  13 - 0xd
      13'h1C90: dout <= 8'b00011111; // 7312 :  31 - 0x1f -- Background 0xc9
      13'h1C91: dout <= 8'b00001111; // 7313 :  15 - 0xf
      13'h1C92: dout <= 8'b11110111; // 7314 : 247 - 0xf7
      13'h1C93: dout <= 8'b10110111; // 7315 : 183 - 0xb7
      13'h1C94: dout <= 8'b11010011; // 7316 : 211 - 0xd3
      13'h1C95: dout <= 8'b10100000; // 7317 : 160 - 0xa0
      13'h1C96: dout <= 8'b11000000; // 7318 : 192 - 0xc0
      13'h1C97: dout <= 8'b00000000; // 7319 :   0 - 0x0
      13'h1C98: dout <= 8'b00001101; // 7320 :  13 - 0xd
      13'h1C99: dout <= 8'b00000101; // 7321 :   5 - 0x5
      13'h1C9A: dout <= 8'b00000011; // 7322 :   3 - 0x3
      13'h1C9B: dout <= 8'b01000011; // 7323 :  67 - 0x43
      13'h1C9C: dout <= 8'b00100000; // 7324 :  32 - 0x20
      13'h1C9D: dout <= 8'b01000000; // 7325 :  64 - 0x40
      13'h1C9E: dout <= 8'b00000000; // 7326 :   0 - 0x0
      13'h1C9F: dout <= 8'b00000000; // 7327 :   0 - 0x0
      13'h1CA0: dout <= 8'b00011100; // 7328 :  28 - 0x1c -- Background 0xca
      13'h1CA1: dout <= 8'b00100010; // 7329 :  34 - 0x22
      13'h1CA2: dout <= 8'b00100100; // 7330 :  36 - 0x24
      13'h1CA3: dout <= 8'b11011110; // 7331 : 222 - 0xde
      13'h1CA4: dout <= 8'b11110000; // 7332 : 240 - 0xf0
      13'h1CA5: dout <= 8'b11111000; // 7333 : 248 - 0xf8
      13'h1CA6: dout <= 8'b11111100; // 7334 : 252 - 0xfc
      13'h1CA7: dout <= 8'b11111100; // 7335 : 252 - 0xfc
      13'h1CA8: dout <= 8'b00000000; // 7336 :   0 - 0x0
      13'h1CA9: dout <= 8'b00011100; // 7337 :  28 - 0x1c
      13'h1CAA: dout <= 8'b00011000; // 7338 :  24 - 0x18
      13'h1CAB: dout <= 8'b00000000; // 7339 :   0 - 0x0
      13'h1CAC: dout <= 8'b00000000; // 7340 :   0 - 0x0
      13'h1CAD: dout <= 8'b10000000; // 7341 : 128 - 0x80
      13'h1CAE: dout <= 8'b11100000; // 7342 : 224 - 0xe0
      13'h1CAF: dout <= 8'b10010000; // 7343 : 144 - 0x90
      13'h1CB0: dout <= 8'b11111100; // 7344 : 252 - 0xfc -- Background 0xcb
      13'h1CB1: dout <= 8'b11111100; // 7345 : 252 - 0xfc
      13'h1CB2: dout <= 8'b11111000; // 7346 : 248 - 0xf8
      13'h1CB3: dout <= 8'b11110000; // 7347 : 240 - 0xf0
      13'h1CB4: dout <= 8'b10011110; // 7348 : 158 - 0x9e
      13'h1CB5: dout <= 8'b00100100; // 7349 :  36 - 0x24
      13'h1CB6: dout <= 8'b00100010; // 7350 :  34 - 0x22
      13'h1CB7: dout <= 8'b00011100; // 7351 :  28 - 0x1c
      13'h1CB8: dout <= 8'b11110000; // 7352 : 240 - 0xf0
      13'h1CB9: dout <= 8'b10010000; // 7353 : 144 - 0x90
      13'h1CBA: dout <= 8'b11110000; // 7354 : 240 - 0xf0
      13'h1CBB: dout <= 8'b10000000; // 7355 : 128 - 0x80
      13'h1CBC: dout <= 8'b00000000; // 7356 :   0 - 0x0
      13'h1CBD: dout <= 8'b00011000; // 7357 :  24 - 0x18
      13'h1CBE: dout <= 8'b00011100; // 7358 :  28 - 0x1c
      13'h1CBF: dout <= 8'b00000000; // 7359 :   0 - 0x0
      13'h1CC0: dout <= 8'b00001110; // 7360 :  14 - 0xe -- Background 0xcc
      13'h1CC1: dout <= 8'b00010110; // 7361 :  22 - 0x16
      13'h1CC2: dout <= 8'b00011010; // 7362 :  26 - 0x1a
      13'h1CC3: dout <= 8'b00000100; // 7363 :   4 - 0x4
      13'h1CC4: dout <= 8'b01101111; // 7364 : 111 - 0x6f
      13'h1CC5: dout <= 8'b10111111; // 7365 : 191 - 0xbf
      13'h1CC6: dout <= 8'b11011111; // 7366 : 223 - 0xdf
      13'h1CC7: dout <= 8'b10111111; // 7367 : 191 - 0xbf
      13'h1CC8: dout <= 8'b00000000; // 7368 :   0 - 0x0
      13'h1CC9: dout <= 8'b00001000; // 7369 :   8 - 0x8
      13'h1CCA: dout <= 8'b00000100; // 7370 :   4 - 0x4
      13'h1CCB: dout <= 8'b00001000; // 7371 :   8 - 0x8
      13'h1CCC: dout <= 8'b00000000; // 7372 :   0 - 0x0
      13'h1CCD: dout <= 8'b01000110; // 7373 :  70 - 0x46
      13'h1CCE: dout <= 8'b00101111; // 7374 :  47 - 0x2f
      13'h1CCF: dout <= 8'b01001110; // 7375 :  78 - 0x4e
      13'h1CD0: dout <= 8'b01011111; // 7376 :  95 - 0x5f -- Background 0xcd
      13'h1CD1: dout <= 8'b00011111; // 7377 :  31 - 0x1f
      13'h1CD2: dout <= 8'b00011111; // 7378 :  31 - 0x1f
      13'h1CD3: dout <= 8'b00001111; // 7379 :  15 - 0xf
      13'h1CD4: dout <= 8'b00111111; // 7380 :  63 - 0x3f
      13'h1CD5: dout <= 8'b00100011; // 7381 :  35 - 0x23
      13'h1CD6: dout <= 8'b00101010; // 7382 :  42 - 0x2a
      13'h1CD7: dout <= 8'b00010100; // 7383 :  20 - 0x14
      13'h1CD8: dout <= 8'b00001101; // 7384 :  13 - 0xd
      13'h1CD9: dout <= 8'b00001011; // 7385 :  11 - 0xb
      13'h1CDA: dout <= 8'b00001111; // 7386 :  15 - 0xf
      13'h1CDB: dout <= 8'b00000110; // 7387 :   6 - 0x6
      13'h1CDC: dout <= 8'b00000011; // 7388 :   3 - 0x3
      13'h1CDD: dout <= 8'b00011100; // 7389 :  28 - 0x1c
      13'h1CDE: dout <= 8'b00010100; // 7390 :  20 - 0x14
      13'h1CDF: dout <= 8'b00000000; // 7391 :   0 - 0x0
      13'h1CE0: dout <= 8'b00000000; // 7392 :   0 - 0x0 -- Background 0xce
      13'h1CE1: dout <= 8'b00000000; // 7393 :   0 - 0x0
      13'h1CE2: dout <= 8'b00000000; // 7394 :   0 - 0x0
      13'h1CE3: dout <= 8'b00000000; // 7395 :   0 - 0x0
      13'h1CE4: dout <= 8'b10001110; // 7396 : 142 - 0x8e
      13'h1CE5: dout <= 8'b11001001; // 7397 : 201 - 0xc9
      13'h1CE6: dout <= 8'b11101010; // 7398 : 234 - 0xea
      13'h1CE7: dout <= 8'b11111001; // 7399 : 249 - 0xf9
      13'h1CE8: dout <= 8'b00000000; // 7400 :   0 - 0x0
      13'h1CE9: dout <= 8'b00000000; // 7401 :   0 - 0x0
      13'h1CEA: dout <= 8'b00000000; // 7402 :   0 - 0x0
      13'h1CEB: dout <= 8'b00000000; // 7403 :   0 - 0x0
      13'h1CEC: dout <= 8'b00000000; // 7404 :   0 - 0x0
      13'h1CED: dout <= 8'b00000110; // 7405 :   6 - 0x6
      13'h1CEE: dout <= 8'b00000100; // 7406 :   4 - 0x4
      13'h1CEF: dout <= 8'b10000110; // 7407 : 134 - 0x86
      13'h1CF0: dout <= 8'b11111110; // 7408 : 254 - 0xfe -- Background 0xcf
      13'h1CF1: dout <= 8'b11111000; // 7409 : 248 - 0xf8
      13'h1CF2: dout <= 8'b11111000; // 7410 : 248 - 0xf8
      13'h1CF3: dout <= 8'b11111000; // 7411 : 248 - 0xf8
      13'h1CF4: dout <= 8'b11110000; // 7412 : 240 - 0xf0
      13'h1CF5: dout <= 8'b11100000; // 7413 : 224 - 0xe0
      13'h1CF6: dout <= 8'b00000000; // 7414 :   0 - 0x0
      13'h1CF7: dout <= 8'b00000000; // 7415 :   0 - 0x0
      13'h1CF8: dout <= 8'b11000000; // 7416 : 192 - 0xc0
      13'h1CF9: dout <= 8'b01100000; // 7417 :  96 - 0x60
      13'h1CFA: dout <= 8'b10100000; // 7418 : 160 - 0xa0
      13'h1CFB: dout <= 8'b11000000; // 7419 : 192 - 0xc0
      13'h1CFC: dout <= 8'b01000000; // 7420 :  64 - 0x40
      13'h1CFD: dout <= 8'b00000000; // 7421 :   0 - 0x0
      13'h1CFE: dout <= 8'b00000000; // 7422 :   0 - 0x0
      13'h1CFF: dout <= 8'b00000000; // 7423 :   0 - 0x0
      13'h1D00: dout <= 8'b00000000; // 7424 :   0 - 0x0 -- Background 0xd0
      13'h1D01: dout <= 8'b00000000; // 7425 :   0 - 0x0
      13'h1D02: dout <= 8'b00000100; // 7426 :   4 - 0x4
      13'h1D03: dout <= 8'b00100110; // 7427 :  38 - 0x26
      13'h1D04: dout <= 8'b00101011; // 7428 :  43 - 0x2b
      13'h1D05: dout <= 8'b01110001; // 7429 : 113 - 0x71
      13'h1D06: dout <= 8'b01000000; // 7430 :  64 - 0x40
      13'h1D07: dout <= 8'b01000111; // 7431 :  71 - 0x47
      13'h1D08: dout <= 8'b00000000; // 7432 :   0 - 0x0
      13'h1D09: dout <= 8'b00000000; // 7433 :   0 - 0x0
      13'h1D0A: dout <= 8'b00000000; // 7434 :   0 - 0x0
      13'h1D0B: dout <= 8'b00000000; // 7435 :   0 - 0x0
      13'h1D0C: dout <= 8'b00000100; // 7436 :   4 - 0x4
      13'h1D0D: dout <= 8'b00001110; // 7437 :  14 - 0xe
      13'h1D0E: dout <= 8'b00111111; // 7438 :  63 - 0x3f
      13'h1D0F: dout <= 8'b00111001; // 7439 :  57 - 0x39
      13'h1D10: dout <= 8'b10001111; // 7440 : 143 - 0x8f -- Background 0xd1
      13'h1D11: dout <= 8'b10001111; // 7441 : 143 - 0x8f
      13'h1D12: dout <= 8'b01001111; // 7442 :  79 - 0x4f
      13'h1D13: dout <= 8'b01001111; // 7443 :  79 - 0x4f
      13'h1D14: dout <= 8'b00111111; // 7444 :  63 - 0x3f
      13'h1D15: dout <= 8'b00010011; // 7445 :  19 - 0x13
      13'h1D16: dout <= 8'b00010001; // 7446 :  17 - 0x11
      13'h1D17: dout <= 8'b00011111; // 7447 :  31 - 0x1f
      13'h1D18: dout <= 8'b01110000; // 7448 : 112 - 0x70
      13'h1D19: dout <= 8'b01111000; // 7449 : 120 - 0x78
      13'h1D1A: dout <= 8'b00111111; // 7450 :  63 - 0x3f
      13'h1D1B: dout <= 8'b00111111; // 7451 :  63 - 0x3f
      13'h1D1C: dout <= 8'b00000011; // 7452 :   3 - 0x3
      13'h1D1D: dout <= 8'b00001100; // 7453 :  12 - 0xc
      13'h1D1E: dout <= 8'b00001110; // 7454 :  14 - 0xe
      13'h1D1F: dout <= 8'b00000000; // 7455 :   0 - 0x0
      13'h1D20: dout <= 8'b00000000; // 7456 :   0 - 0x0 -- Background 0xd2
      13'h1D21: dout <= 8'b10000000; // 7457 : 128 - 0x80
      13'h1D22: dout <= 8'b11001000; // 7458 : 200 - 0xc8
      13'h1D23: dout <= 8'b11010100; // 7459 : 212 - 0xd4
      13'h1D24: dout <= 8'b00100100; // 7460 :  36 - 0x24
      13'h1D25: dout <= 8'b00000010; // 7461 :   2 - 0x2
      13'h1D26: dout <= 8'b00000010; // 7462 :   2 - 0x2
      13'h1D27: dout <= 8'b11110010; // 7463 : 242 - 0xf2
      13'h1D28: dout <= 8'b00000000; // 7464 :   0 - 0x0
      13'h1D29: dout <= 8'b00000000; // 7465 :   0 - 0x0
      13'h1D2A: dout <= 8'b00000000; // 7466 :   0 - 0x0
      13'h1D2B: dout <= 8'b00001000; // 7467 :   8 - 0x8
      13'h1D2C: dout <= 8'b11011000; // 7468 : 216 - 0xd8
      13'h1D2D: dout <= 8'b11111100; // 7469 : 252 - 0xfc
      13'h1D2E: dout <= 8'b11111100; // 7470 : 252 - 0xfc
      13'h1D2F: dout <= 8'b10011100; // 7471 : 156 - 0x9c
      13'h1D30: dout <= 8'b11110010; // 7472 : 242 - 0xf2 -- Background 0xd3
      13'h1D31: dout <= 8'b11110010; // 7473 : 242 - 0xf2
      13'h1D32: dout <= 8'b11110100; // 7474 : 244 - 0xf4
      13'h1D33: dout <= 8'b11110100; // 7475 : 244 - 0xf4
      13'h1D34: dout <= 8'b11110100; // 7476 : 244 - 0xf4
      13'h1D35: dout <= 8'b11001000; // 7477 : 200 - 0xc8
      13'h1D36: dout <= 8'b01000100; // 7478 :  68 - 0x44
      13'h1D37: dout <= 8'b01111100; // 7479 : 124 - 0x7c
      13'h1D38: dout <= 8'b00001100; // 7480 :  12 - 0xc
      13'h1D39: dout <= 8'b10011100; // 7481 : 156 - 0x9c
      13'h1D3A: dout <= 8'b11111000; // 7482 : 248 - 0xf8
      13'h1D3B: dout <= 8'b01111000; // 7483 : 120 - 0x78
      13'h1D3C: dout <= 8'b10001000; // 7484 : 136 - 0x88
      13'h1D3D: dout <= 8'b00110000; // 7485 :  48 - 0x30
      13'h1D3E: dout <= 8'b00111000; // 7486 :  56 - 0x38
      13'h1D3F: dout <= 8'b00000000; // 7487 :   0 - 0x0
      13'h1D40: dout <= 8'b00000000; // 7488 :   0 - 0x0 -- Background 0xd4
      13'h1D41: dout <= 8'b00000000; // 7489 :   0 - 0x0
      13'h1D42: dout <= 8'b00000000; // 7490 :   0 - 0x0
      13'h1D43: dout <= 8'b00001001; // 7491 :   9 - 0x9
      13'h1D44: dout <= 8'b00011010; // 7492 :  26 - 0x1a
      13'h1D45: dout <= 8'b00010100; // 7493 :  20 - 0x14
      13'h1D46: dout <= 8'b00100000; // 7494 :  32 - 0x20
      13'h1D47: dout <= 8'b01000111; // 7495 :  71 - 0x47
      13'h1D48: dout <= 8'b00000000; // 7496 :   0 - 0x0
      13'h1D49: dout <= 8'b00000000; // 7497 :   0 - 0x0
      13'h1D4A: dout <= 8'b00000000; // 7498 :   0 - 0x0
      13'h1D4B: dout <= 8'b00000000; // 7499 :   0 - 0x0
      13'h1D4C: dout <= 8'b00000001; // 7500 :   1 - 0x1
      13'h1D4D: dout <= 8'b00001011; // 7501 :  11 - 0xb
      13'h1D4E: dout <= 8'b00011111; // 7502 :  31 - 0x1f
      13'h1D4F: dout <= 8'b00111001; // 7503 :  57 - 0x39
      13'h1D50: dout <= 8'b10001111; // 7504 : 143 - 0x8f -- Background 0xd5
      13'h1D51: dout <= 8'b10001111; // 7505 : 143 - 0x8f
      13'h1D52: dout <= 8'b01001111; // 7506 :  79 - 0x4f
      13'h1D53: dout <= 8'b01001111; // 7507 :  79 - 0x4f
      13'h1D54: dout <= 8'b00111111; // 7508 :  63 - 0x3f
      13'h1D55: dout <= 8'b01000111; // 7509 :  71 - 0x47
      13'h1D56: dout <= 8'b00100010; // 7510 :  34 - 0x22
      13'h1D57: dout <= 8'b00011100; // 7511 :  28 - 0x1c
      13'h1D58: dout <= 8'b01110000; // 7512 : 112 - 0x70
      13'h1D59: dout <= 8'b01111000; // 7513 : 120 - 0x78
      13'h1D5A: dout <= 8'b00111111; // 7514 :  63 - 0x3f
      13'h1D5B: dout <= 8'b00111111; // 7515 :  63 - 0x3f
      13'h1D5C: dout <= 8'b00000011; // 7516 :   3 - 0x3
      13'h1D5D: dout <= 8'b00111000; // 7517 :  56 - 0x38
      13'h1D5E: dout <= 8'b00011100; // 7518 :  28 - 0x1c
      13'h1D5F: dout <= 8'b00000000; // 7519 :   0 - 0x0
      13'h1D60: dout <= 8'b00000000; // 7520 :   0 - 0x0 -- Background 0xd6
      13'h1D61: dout <= 8'b01000000; // 7521 :  64 - 0x40
      13'h1D62: dout <= 8'b11000000; // 7522 : 192 - 0xc0
      13'h1D63: dout <= 8'b00101100; // 7523 :  44 - 0x2c
      13'h1D64: dout <= 8'b00110100; // 7524 :  52 - 0x34
      13'h1D65: dout <= 8'b00000100; // 7525 :   4 - 0x4
      13'h1D66: dout <= 8'b00000010; // 7526 :   2 - 0x2
      13'h1D67: dout <= 8'b11110010; // 7527 : 242 - 0xf2
      13'h1D68: dout <= 8'b00000000; // 7528 :   0 - 0x0
      13'h1D69: dout <= 8'b00000000; // 7529 :   0 - 0x0
      13'h1D6A: dout <= 8'b00000000; // 7530 :   0 - 0x0
      13'h1D6B: dout <= 8'b11000000; // 7531 : 192 - 0xc0
      13'h1D6C: dout <= 8'b11001000; // 7532 : 200 - 0xc8
      13'h1D6D: dout <= 8'b11111000; // 7533 : 248 - 0xf8
      13'h1D6E: dout <= 8'b11111100; // 7534 : 252 - 0xfc
      13'h1D6F: dout <= 8'b10011100; // 7535 : 156 - 0x9c
      13'h1D70: dout <= 8'b11110010; // 7536 : 242 - 0xf2 -- Background 0xd7
      13'h1D71: dout <= 8'b11110010; // 7537 : 242 - 0xf2
      13'h1D72: dout <= 8'b11110100; // 7538 : 244 - 0xf4
      13'h1D73: dout <= 8'b11110111; // 7539 : 247 - 0xf7
      13'h1D74: dout <= 8'b11111101; // 7540 : 253 - 0xfd
      13'h1D75: dout <= 8'b11100001; // 7541 : 225 - 0xe1
      13'h1D76: dout <= 8'b00010010; // 7542 :  18 - 0x12
      13'h1D77: dout <= 8'b00001100; // 7543 :  12 - 0xc
      13'h1D78: dout <= 8'b00001100; // 7544 :  12 - 0xc
      13'h1D79: dout <= 8'b10011100; // 7545 : 156 - 0x9c
      13'h1D7A: dout <= 8'b11111000; // 7546 : 248 - 0xf8
      13'h1D7B: dout <= 8'b01111000; // 7547 : 120 - 0x78
      13'h1D7C: dout <= 8'b11100010; // 7548 : 226 - 0xe2
      13'h1D7D: dout <= 8'b00011110; // 7549 :  30 - 0x1e
      13'h1D7E: dout <= 8'b00001100; // 7550 :  12 - 0xc
      13'h1D7F: dout <= 8'b00000000; // 7551 :   0 - 0x0
      13'h1D80: dout <= 8'b01111000; // 7552 : 120 - 0x78 -- Background 0xd8
      13'h1D81: dout <= 8'b01001110; // 7553 :  78 - 0x4e
      13'h1D82: dout <= 8'b11000010; // 7554 : 194 - 0xc2
      13'h1D83: dout <= 8'b10011010; // 7555 : 154 - 0x9a
      13'h1D84: dout <= 8'b10011011; // 7556 : 155 - 0x9b
      13'h1D85: dout <= 8'b11011001; // 7557 : 217 - 0xd9
      13'h1D86: dout <= 8'b01100011; // 7558 :  99 - 0x63
      13'h1D87: dout <= 8'b00111110; // 7559 :  62 - 0x3e
      13'h1D88: dout <= 8'b00000000; // 7560 :   0 - 0x0
      13'h1D89: dout <= 8'b00110000; // 7561 :  48 - 0x30
      13'h1D8A: dout <= 8'b00111100; // 7562 :  60 - 0x3c
      13'h1D8B: dout <= 8'b01111100; // 7563 : 124 - 0x7c
      13'h1D8C: dout <= 8'b01111100; // 7564 : 124 - 0x7c
      13'h1D8D: dout <= 8'b00111110; // 7565 :  62 - 0x3e
      13'h1D8E: dout <= 8'b00011100; // 7566 :  28 - 0x1c
      13'h1D8F: dout <= 8'b00000000; // 7567 :   0 - 0x0
      13'h1D90: dout <= 8'b00011110; // 7568 :  30 - 0x1e -- Background 0xd9
      13'h1D91: dout <= 8'b01110001; // 7569 : 113 - 0x71
      13'h1D92: dout <= 8'b01001001; // 7570 :  73 - 0x49
      13'h1D93: dout <= 8'b10111001; // 7571 : 185 - 0xb9
      13'h1D94: dout <= 8'b10011101; // 7572 : 157 - 0x9d
      13'h1D95: dout <= 8'b01010010; // 7573 :  82 - 0x52
      13'h1D96: dout <= 8'b01110010; // 7574 : 114 - 0x72
      13'h1D97: dout <= 8'b00011110; // 7575 :  30 - 0x1e
      13'h1D98: dout <= 8'b00000000; // 7576 :   0 - 0x0
      13'h1D99: dout <= 8'b00001110; // 7577 :  14 - 0xe
      13'h1D9A: dout <= 8'b00111110; // 7578 :  62 - 0x3e
      13'h1D9B: dout <= 8'b01111110; // 7579 : 126 - 0x7e
      13'h1D9C: dout <= 8'b01111110; // 7580 : 126 - 0x7e
      13'h1D9D: dout <= 8'b00111100; // 7581 :  60 - 0x3c
      13'h1D9E: dout <= 8'b00001100; // 7582 :  12 - 0xc
      13'h1D9F: dout <= 8'b00000000; // 7583 :   0 - 0x0
      13'h1DA0: dout <= 8'b01100000; // 7584 :  96 - 0x60 -- Background 0xda
      13'h1DA1: dout <= 8'b01011110; // 7585 :  94 - 0x5e
      13'h1DA2: dout <= 8'b10001001; // 7586 : 137 - 0x89
      13'h1DA3: dout <= 8'b10111101; // 7587 : 189 - 0xbd
      13'h1DA4: dout <= 8'b10011101; // 7588 : 157 - 0x9d
      13'h1DA5: dout <= 8'b11010011; // 7589 : 211 - 0xd3
      13'h1DA6: dout <= 8'b01000110; // 7590 :  70 - 0x46
      13'h1DA7: dout <= 8'b01111100; // 7591 : 124 - 0x7c
      13'h1DA8: dout <= 8'b00000000; // 7592 :   0 - 0x0
      13'h1DA9: dout <= 8'b00100000; // 7593 :  32 - 0x20
      13'h1DAA: dout <= 8'b01111110; // 7594 : 126 - 0x7e
      13'h1DAB: dout <= 8'b01111110; // 7595 : 126 - 0x7e
      13'h1DAC: dout <= 8'b01111110; // 7596 : 126 - 0x7e
      13'h1DAD: dout <= 8'b00111100; // 7597 :  60 - 0x3c
      13'h1DAE: dout <= 8'b00111000; // 7598 :  56 - 0x38
      13'h1DAF: dout <= 8'b00000000; // 7599 :   0 - 0x0
      13'h1DB0: dout <= 8'b00011110; // 7600 :  30 - 0x1e -- Background 0xdb
      13'h1DB1: dout <= 8'b00100011; // 7601 :  35 - 0x23
      13'h1DB2: dout <= 8'b01001001; // 7602 :  73 - 0x49
      13'h1DB3: dout <= 8'b10111101; // 7603 : 189 - 0xbd
      13'h1DB4: dout <= 8'b10011001; // 7604 : 153 - 0x99
      13'h1DB5: dout <= 8'b01000011; // 7605 :  67 - 0x43
      13'h1DB6: dout <= 8'b01101110; // 7606 : 110 - 0x6e
      13'h1DB7: dout <= 8'b00011000; // 7607 :  24 - 0x18
      13'h1DB8: dout <= 8'b00000000; // 7608 :   0 - 0x0
      13'h1DB9: dout <= 8'b00011100; // 7609 :  28 - 0x1c
      13'h1DBA: dout <= 8'b00111110; // 7610 :  62 - 0x3e
      13'h1DBB: dout <= 8'b01111110; // 7611 : 126 - 0x7e
      13'h1DBC: dout <= 8'b01111110; // 7612 : 126 - 0x7e
      13'h1DBD: dout <= 8'b00111100; // 7613 :  60 - 0x3c
      13'h1DBE: dout <= 8'b00010000; // 7614 :  16 - 0x10
      13'h1DBF: dout <= 8'b00000000; // 7615 :   0 - 0x0
      13'h1DC0: dout <= 8'b00000000; // 7616 :   0 - 0x0 -- Background 0xdc
      13'h1DC1: dout <= 8'b00000000; // 7617 :   0 - 0x0
      13'h1DC2: dout <= 8'b00000001; // 7618 :   1 - 0x1
      13'h1DC3: dout <= 8'b00000010; // 7619 :   2 - 0x2
      13'h1DC4: dout <= 8'b00000100; // 7620 :   4 - 0x4
      13'h1DC5: dout <= 8'b00000010; // 7621 :   2 - 0x2
      13'h1DC6: dout <= 8'b00011110; // 7622 :  30 - 0x1e
      13'h1DC7: dout <= 8'b00010000; // 7623 :  16 - 0x10
      13'h1DC8: dout <= 8'b00000000; // 7624 :   0 - 0x0
      13'h1DC9: dout <= 8'b00000000; // 7625 :   0 - 0x0
      13'h1DCA: dout <= 8'b00000000; // 7626 :   0 - 0x0
      13'h1DCB: dout <= 8'b00000001; // 7627 :   1 - 0x1
      13'h1DCC: dout <= 8'b00000011; // 7628 :   3 - 0x3
      13'h1DCD: dout <= 8'b00000001; // 7629 :   1 - 0x1
      13'h1DCE: dout <= 8'b00000001; // 7630 :   1 - 0x1
      13'h1DCF: dout <= 8'b00001111; // 7631 :  15 - 0xf
      13'h1DD0: dout <= 8'b00001000; // 7632 :   8 - 0x8 -- Background 0xdd
      13'h1DD1: dout <= 8'b00001101; // 7633 :  13 - 0xd
      13'h1DD2: dout <= 8'b00111010; // 7634 :  58 - 0x3a
      13'h1DD3: dout <= 8'b00100101; // 7635 :  37 - 0x25
      13'h1DD4: dout <= 8'b00011011; // 7636 :  27 - 0x1b
      13'h1DD5: dout <= 8'b00001111; // 7637 :  15 - 0xf
      13'h1DD6: dout <= 8'b00000111; // 7638 :   7 - 0x7
      13'h1DD7: dout <= 8'b00000011; // 7639 :   3 - 0x3
      13'h1DD8: dout <= 8'b00000111; // 7640 :   7 - 0x7
      13'h1DD9: dout <= 8'b00000111; // 7641 :   7 - 0x7
      13'h1DDA: dout <= 8'b00000111; // 7642 :   7 - 0x7
      13'h1DDB: dout <= 8'b00011111; // 7643 :  31 - 0x1f
      13'h1DDC: dout <= 8'b00001111; // 7644 :  15 - 0xf
      13'h1DDD: dout <= 8'b00000111; // 7645 :   7 - 0x7
      13'h1DDE: dout <= 8'b00000011; // 7646 :   3 - 0x3
      13'h1DDF: dout <= 8'b00000000; // 7647 :   0 - 0x0
      13'h1DE0: dout <= 8'b00000000; // 7648 :   0 - 0x0 -- Background 0xde
      13'h1DE1: dout <= 8'b00000000; // 7649 :   0 - 0x0
      13'h1DE2: dout <= 8'b00000000; // 7650 :   0 - 0x0
      13'h1DE3: dout <= 8'b11000000; // 7651 : 192 - 0xc0
      13'h1DE4: dout <= 8'b01000000; // 7652 :  64 - 0x40
      13'h1DE5: dout <= 8'b01011000; // 7653 :  88 - 0x58
      13'h1DE6: dout <= 8'b01101000; // 7654 : 104 - 0x68
      13'h1DE7: dout <= 8'b00001000; // 7655 :   8 - 0x8
      13'h1DE8: dout <= 8'b00000000; // 7656 :   0 - 0x0
      13'h1DE9: dout <= 8'b00000000; // 7657 :   0 - 0x0
      13'h1DEA: dout <= 8'b00000000; // 7658 :   0 - 0x0
      13'h1DEB: dout <= 8'b00000000; // 7659 :   0 - 0x0
      13'h1DEC: dout <= 8'b10000000; // 7660 : 128 - 0x80
      13'h1DED: dout <= 8'b10000000; // 7661 : 128 - 0x80
      13'h1DEE: dout <= 8'b10010000; // 7662 : 144 - 0x90
      13'h1DEF: dout <= 8'b11110000; // 7663 : 240 - 0xf0
      13'h1DF0: dout <= 8'b00010000; // 7664 :  16 - 0x10 -- Background 0xdf
      13'h1DF1: dout <= 8'b01011100; // 7665 :  92 - 0x5c
      13'h1DF2: dout <= 8'b10101000; // 7666 : 168 - 0xa8
      13'h1DF3: dout <= 8'b11011000; // 7667 : 216 - 0xd8
      13'h1DF4: dout <= 8'b10111000; // 7668 : 184 - 0xb8
      13'h1DF5: dout <= 8'b11110000; // 7669 : 240 - 0xf0
      13'h1DF6: dout <= 8'b11100000; // 7670 : 224 - 0xe0
      13'h1DF7: dout <= 8'b11000000; // 7671 : 192 - 0xc0
      13'h1DF8: dout <= 8'b11100000; // 7672 : 224 - 0xe0
      13'h1DF9: dout <= 8'b11100000; // 7673 : 224 - 0xe0
      13'h1DFA: dout <= 8'b11110000; // 7674 : 240 - 0xf0
      13'h1DFB: dout <= 8'b11110000; // 7675 : 240 - 0xf0
      13'h1DFC: dout <= 8'b11100000; // 7676 : 224 - 0xe0
      13'h1DFD: dout <= 8'b11000000; // 7677 : 192 - 0xc0
      13'h1DFE: dout <= 8'b11000000; // 7678 : 192 - 0xc0
      13'h1DFF: dout <= 8'b00000000; // 7679 :   0 - 0x0
      13'h1E00: dout <= 8'b00000000; // 7680 :   0 - 0x0 -- Background 0xe0
      13'h1E01: dout <= 8'b00000000; // 7681 :   0 - 0x0
      13'h1E02: dout <= 8'b00000000; // 7682 :   0 - 0x0
      13'h1E03: dout <= 8'b00010011; // 7683 :  19 - 0x13
      13'h1E04: dout <= 8'b00010011; // 7684 :  19 - 0x13
      13'h1E05: dout <= 8'b00110111; // 7685 :  55 - 0x37
      13'h1E06: dout <= 8'b00110111; // 7686 :  55 - 0x37
      13'h1E07: dout <= 8'b00000111; // 7687 :   7 - 0x7
      13'h1E08: dout <= 8'b00001111; // 7688 :  15 - 0xf
      13'h1E09: dout <= 8'b00011111; // 7689 :  31 - 0x1f
      13'h1E0A: dout <= 8'b00011111; // 7690 :  31 - 0x1f
      13'h1E0B: dout <= 8'b00111111; // 7691 :  63 - 0x3f
      13'h1E0C: dout <= 8'b01111111; // 7692 : 127 - 0x7f
      13'h1E0D: dout <= 8'b11111111; // 7693 : 255 - 0xff
      13'h1E0E: dout <= 8'b11111111; // 7694 : 255 - 0xff
      13'h1E0F: dout <= 8'b11111111; // 7695 : 255 - 0xff
      13'h1E10: dout <= 8'b00000111; // 7696 :   7 - 0x7 -- Background 0xe1
      13'h1E11: dout <= 8'b00000100; // 7697 :   4 - 0x4
      13'h1E12: dout <= 8'b00000000; // 7698 :   0 - 0x0
      13'h1E13: dout <= 8'b00000000; // 7699 :   0 - 0x0
      13'h1E14: dout <= 8'b00000000; // 7700 :   0 - 0x0
      13'h1E15: dout <= 8'b00100000; // 7701 :  32 - 0x20
      13'h1E16: dout <= 8'b01110000; // 7702 : 112 - 0x70
      13'h1E17: dout <= 8'b11111000; // 7703 : 248 - 0xf8
      13'h1E18: dout <= 8'b11111111; // 7704 : 255 - 0xff
      13'h1E19: dout <= 8'b11111111; // 7705 : 255 - 0xff
      13'h1E1A: dout <= 8'b01111111; // 7706 : 127 - 0x7f
      13'h1E1B: dout <= 8'b00111111; // 7707 :  63 - 0x3f
      13'h1E1C: dout <= 8'b00111111; // 7708 :  63 - 0x3f
      13'h1E1D: dout <= 8'b00011111; // 7709 :  31 - 0x1f
      13'h1E1E: dout <= 8'b00001111; // 7710 :  15 - 0xf
      13'h1E1F: dout <= 8'b00000111; // 7711 :   7 - 0x7
      13'h1E20: dout <= 8'b00000000; // 7712 :   0 - 0x0 -- Background 0xe2
      13'h1E21: dout <= 8'b00000000; // 7713 :   0 - 0x0
      13'h1E22: dout <= 8'b00000000; // 7714 :   0 - 0x0
      13'h1E23: dout <= 8'b11111000; // 7715 : 248 - 0xf8
      13'h1E24: dout <= 8'b11111100; // 7716 : 252 - 0xfc
      13'h1E25: dout <= 8'b11111100; // 7717 : 252 - 0xfc
      13'h1E26: dout <= 8'b11111100; // 7718 : 252 - 0xfc
      13'h1E27: dout <= 8'b11111101; // 7719 : 253 - 0xfd
      13'h1E28: dout <= 8'b11111110; // 7720 : 254 - 0xfe
      13'h1E29: dout <= 8'b11111111; // 7721 : 255 - 0xff
      13'h1E2A: dout <= 8'b11111111; // 7722 : 255 - 0xff
      13'h1E2B: dout <= 8'b00001111; // 7723 :  15 - 0xf
      13'h1E2C: dout <= 8'b10111111; // 7724 : 191 - 0xbf
      13'h1E2D: dout <= 8'b10100011; // 7725 : 163 - 0xa3
      13'h1E2E: dout <= 8'b11110111; // 7726 : 247 - 0xf7
      13'h1E2F: dout <= 8'b11110111; // 7727 : 247 - 0xf7
      13'h1E30: dout <= 8'b11111100; // 7728 : 252 - 0xfc -- Background 0xe3
      13'h1E31: dout <= 8'b00011100; // 7729 :  28 - 0x1c
      13'h1E32: dout <= 8'b11000000; // 7730 : 192 - 0xc0
      13'h1E33: dout <= 8'b11100000; // 7731 : 224 - 0xe0
      13'h1E34: dout <= 8'b00000000; // 7732 :   0 - 0x0
      13'h1E35: dout <= 8'b00000000; // 7733 :   0 - 0x0
      13'h1E36: dout <= 8'b00000110; // 7734 :   6 - 0x6
      13'h1E37: dout <= 8'b00001111; // 7735 :  15 - 0xf
      13'h1E38: dout <= 8'b11111111; // 7736 : 255 - 0xff
      13'h1E39: dout <= 8'b11111111; // 7737 : 255 - 0xff
      13'h1E3A: dout <= 8'b00111111; // 7738 :  63 - 0x3f
      13'h1E3B: dout <= 8'b00011111; // 7739 :  31 - 0x1f
      13'h1E3C: dout <= 8'b11111110; // 7740 : 254 - 0xfe
      13'h1E3D: dout <= 8'b11111100; // 7741 : 252 - 0xfc
      13'h1E3E: dout <= 8'b11111000; // 7742 : 248 - 0xf8
      13'h1E3F: dout <= 8'b11110000; // 7743 : 240 - 0xf0
      13'h1E40: dout <= 8'b00000000; // 7744 :   0 - 0x0 -- Background 0xe4
      13'h1E41: dout <= 8'b00000000; // 7745 :   0 - 0x0
      13'h1E42: dout <= 8'b00000000; // 7746 :   0 - 0x0
      13'h1E43: dout <= 8'b00010011; // 7747 :  19 - 0x13
      13'h1E44: dout <= 8'b00010011; // 7748 :  19 - 0x13
      13'h1E45: dout <= 8'b00110111; // 7749 :  55 - 0x37
      13'h1E46: dout <= 8'b00110111; // 7750 :  55 - 0x37
      13'h1E47: dout <= 8'b00000111; // 7751 :   7 - 0x7
      13'h1E48: dout <= 8'b00001111; // 7752 :  15 - 0xf
      13'h1E49: dout <= 8'b00011111; // 7753 :  31 - 0x1f
      13'h1E4A: dout <= 8'b00011111; // 7754 :  31 - 0x1f
      13'h1E4B: dout <= 8'b00111111; // 7755 :  63 - 0x3f
      13'h1E4C: dout <= 8'b01111111; // 7756 : 127 - 0x7f
      13'h1E4D: dout <= 8'b11111111; // 7757 : 255 - 0xff
      13'h1E4E: dout <= 8'b11111111; // 7758 : 255 - 0xff
      13'h1E4F: dout <= 8'b11111111; // 7759 : 255 - 0xff
      13'h1E50: dout <= 8'b00000111; // 7760 :   7 - 0x7 -- Background 0xe5
      13'h1E51: dout <= 8'b00000100; // 7761 :   4 - 0x4
      13'h1E52: dout <= 8'b00000001; // 7762 :   1 - 0x1
      13'h1E53: dout <= 8'b00000000; // 7763 :   0 - 0x0
      13'h1E54: dout <= 8'b00000000; // 7764 :   0 - 0x0
      13'h1E55: dout <= 8'b00100000; // 7765 :  32 - 0x20
      13'h1E56: dout <= 8'b01110000; // 7766 : 112 - 0x70
      13'h1E57: dout <= 8'b11111000; // 7767 : 248 - 0xf8
      13'h1E58: dout <= 8'b11111111; // 7768 : 255 - 0xff
      13'h1E59: dout <= 8'b11111111; // 7769 : 255 - 0xff
      13'h1E5A: dout <= 8'b01111110; // 7770 : 126 - 0x7e
      13'h1E5B: dout <= 8'b00111111; // 7771 :  63 - 0x3f
      13'h1E5C: dout <= 8'b00111111; // 7772 :  63 - 0x3f
      13'h1E5D: dout <= 8'b00011111; // 7773 :  31 - 0x1f
      13'h1E5E: dout <= 8'b00001111; // 7774 :  15 - 0xf
      13'h1E5F: dout <= 8'b00000111; // 7775 :   7 - 0x7
      13'h1E60: dout <= 8'b00000000; // 7776 :   0 - 0x0 -- Background 0xe6
      13'h1E61: dout <= 8'b00000000; // 7777 :   0 - 0x0
      13'h1E62: dout <= 8'b00000000; // 7778 :   0 - 0x0
      13'h1E63: dout <= 8'b11111100; // 7779 : 252 - 0xfc
      13'h1E64: dout <= 8'b11111100; // 7780 : 252 - 0xfc
      13'h1E65: dout <= 8'b11111100; // 7781 : 252 - 0xfc
      13'h1E66: dout <= 8'b11111100; // 7782 : 252 - 0xfc
      13'h1E67: dout <= 8'b11111101; // 7783 : 253 - 0xfd
      13'h1E68: dout <= 8'b11111110; // 7784 : 254 - 0xfe
      13'h1E69: dout <= 8'b11111111; // 7785 : 255 - 0xff
      13'h1E6A: dout <= 8'b11111111; // 7786 : 255 - 0xff
      13'h1E6B: dout <= 8'b11100011; // 7787 : 227 - 0xe3
      13'h1E6C: dout <= 8'b00010111; // 7788 :  23 - 0x17
      13'h1E6D: dout <= 8'b10110111; // 7789 : 183 - 0xb7
      13'h1E6E: dout <= 8'b10111111; // 7790 : 191 - 0xbf
      13'h1E6F: dout <= 8'b11111111; // 7791 : 255 - 0xff
      13'h1E70: dout <= 8'b11111100; // 7792 : 252 - 0xfc -- Background 0xe7
      13'h1E71: dout <= 8'b00001100; // 7793 :  12 - 0xc
      13'h1E72: dout <= 8'b11000000; // 7794 : 192 - 0xc0
      13'h1E73: dout <= 8'b11110000; // 7795 : 240 - 0xf0
      13'h1E74: dout <= 8'b11110000; // 7796 : 240 - 0xf0
      13'h1E75: dout <= 8'b00000000; // 7797 :   0 - 0x0
      13'h1E76: dout <= 8'b00000110; // 7798 :   6 - 0x6
      13'h1E77: dout <= 8'b00001111; // 7799 :  15 - 0xf
      13'h1E78: dout <= 8'b11111111; // 7800 : 255 - 0xff
      13'h1E79: dout <= 8'b11111111; // 7801 : 255 - 0xff
      13'h1E7A: dout <= 8'b00111111; // 7802 :  63 - 0x3f
      13'h1E7B: dout <= 8'b00001111; // 7803 :  15 - 0xf
      13'h1E7C: dout <= 8'b00001110; // 7804 :  14 - 0xe
      13'h1E7D: dout <= 8'b11111100; // 7805 : 252 - 0xfc
      13'h1E7E: dout <= 8'b11111000; // 7806 : 248 - 0xf8
      13'h1E7F: dout <= 8'b11110000; // 7807 : 240 - 0xf0
      13'h1E80: dout <= 8'b11111111; // 7808 : 255 - 0xff -- Background 0xe8
      13'h1E81: dout <= 8'b11111111; // 7809 : 255 - 0xff
      13'h1E82: dout <= 8'b01111111; // 7810 : 127 - 0x7f
      13'h1E83: dout <= 8'b01111111; // 7811 : 127 - 0x7f
      13'h1E84: dout <= 8'b01111111; // 7812 : 127 - 0x7f
      13'h1E85: dout <= 8'b00111111; // 7813 :  63 - 0x3f
      13'h1E86: dout <= 8'b00111111; // 7814 :  63 - 0x3f
      13'h1E87: dout <= 8'b00111111; // 7815 :  63 - 0x3f
      13'h1E88: dout <= 8'b00000000; // 7816 :   0 - 0x0
      13'h1E89: dout <= 8'b00000101; // 7817 :   5 - 0x5
      13'h1E8A: dout <= 8'b00000111; // 7818 :   7 - 0x7
      13'h1E8B: dout <= 8'b00000011; // 7819 :   3 - 0x3
      13'h1E8C: dout <= 8'b00000000; // 7820 :   0 - 0x0
      13'h1E8D: dout <= 8'b00000000; // 7821 :   0 - 0x0
      13'h1E8E: dout <= 8'b00000000; // 7822 :   0 - 0x0
      13'h1E8F: dout <= 8'b00000000; // 7823 :   0 - 0x0
      13'h1E90: dout <= 8'b00111100; // 7824 :  60 - 0x3c -- Background 0xe9
      13'h1E91: dout <= 8'b00111110; // 7825 :  62 - 0x3e
      13'h1E92: dout <= 8'b00011111; // 7826 :  31 - 0x1f
      13'h1E93: dout <= 8'b00001111; // 7827 :  15 - 0xf
      13'h1E94: dout <= 8'b00000111; // 7828 :   7 - 0x7
      13'h1E95: dout <= 8'b00000000; // 7829 :   0 - 0x0
      13'h1E96: dout <= 8'b00000000; // 7830 :   0 - 0x0
      13'h1E97: dout <= 8'b00000000; // 7831 :   0 - 0x0
      13'h1E98: dout <= 8'b00000000; // 7832 :   0 - 0x0
      13'h1E99: dout <= 8'b00000000; // 7833 :   0 - 0x0
      13'h1E9A: dout <= 8'b00000000; // 7834 :   0 - 0x0
      13'h1E9B: dout <= 8'b00000000; // 7835 :   0 - 0x0
      13'h1E9C: dout <= 8'b00000000; // 7836 :   0 - 0x0
      13'h1E9D: dout <= 8'b00000000; // 7837 :   0 - 0x0
      13'h1E9E: dout <= 8'b00000000; // 7838 :   0 - 0x0
      13'h1E9F: dout <= 8'b00000000; // 7839 :   0 - 0x0
      13'h1EA0: dout <= 8'b11111111; // 7840 : 255 - 0xff -- Background 0xea
      13'h1EA1: dout <= 8'b11111110; // 7841 : 254 - 0xfe
      13'h1EA2: dout <= 8'b11111110; // 7842 : 254 - 0xfe
      13'h1EA3: dout <= 8'b11111100; // 7843 : 252 - 0xfc
      13'h1EA4: dout <= 8'b11111000; // 7844 : 248 - 0xf8
      13'h1EA5: dout <= 8'b11110000; // 7845 : 240 - 0xf0
      13'h1EA6: dout <= 8'b10110000; // 7846 : 176 - 0xb0
      13'h1EA7: dout <= 8'b00111001; // 7847 :  57 - 0x39
      13'h1EA8: dout <= 8'b00000011; // 7848 :   3 - 0x3
      13'h1EA9: dout <= 8'b10011110; // 7849 : 158 - 0x9e
      13'h1EAA: dout <= 8'b00001110; // 7850 :  14 - 0xe
      13'h1EAB: dout <= 8'b00000000; // 7851 :   0 - 0x0
      13'h1EAC: dout <= 8'b00000000; // 7852 :   0 - 0x0
      13'h1EAD: dout <= 8'b00000000; // 7853 :   0 - 0x0
      13'h1EAE: dout <= 8'b00000000; // 7854 :   0 - 0x0
      13'h1EAF: dout <= 8'b00000000; // 7855 :   0 - 0x0
      13'h1EB0: dout <= 8'b00011111; // 7856 :  31 - 0x1f -- Background 0xeb
      13'h1EB1: dout <= 8'b11001111; // 7857 : 207 - 0xcf
      13'h1EB2: dout <= 8'b11000110; // 7858 : 198 - 0xc6
      13'h1EB3: dout <= 8'b10000000; // 7859 : 128 - 0x80
      13'h1EB4: dout <= 8'b00000000; // 7860 :   0 - 0x0
      13'h1EB5: dout <= 8'b00000000; // 7861 :   0 - 0x0
      13'h1EB6: dout <= 8'b00000000; // 7862 :   0 - 0x0
      13'h1EB7: dout <= 8'b00000000; // 7863 :   0 - 0x0
      13'h1EB8: dout <= 8'b00000000; // 7864 :   0 - 0x0
      13'h1EB9: dout <= 8'b00000000; // 7865 :   0 - 0x0
      13'h1EBA: dout <= 8'b00000000; // 7866 :   0 - 0x0
      13'h1EBB: dout <= 8'b00000000; // 7867 :   0 - 0x0
      13'h1EBC: dout <= 8'b00000000; // 7868 :   0 - 0x0
      13'h1EBD: dout <= 8'b00000000; // 7869 :   0 - 0x0
      13'h1EBE: dout <= 8'b00000000; // 7870 :   0 - 0x0
      13'h1EBF: dout <= 8'b00000000; // 7871 :   0 - 0x0
      13'h1EC0: dout <= 8'b00000000; // 7872 :   0 - 0x0 -- Background 0xec
      13'h1EC1: dout <= 8'b00000000; // 7873 :   0 - 0x0
      13'h1EC2: dout <= 8'b00000000; // 7874 :   0 - 0x0
      13'h1EC3: dout <= 8'b00000000; // 7875 :   0 - 0x0
      13'h1EC4: dout <= 8'b00000000; // 7876 :   0 - 0x0
      13'h1EC5: dout <= 8'b00000000; // 7877 :   0 - 0x0
      13'h1EC6: dout <= 8'b00001100; // 7878 :  12 - 0xc
      13'h1EC7: dout <= 8'b00001100; // 7879 :  12 - 0xc
      13'h1EC8: dout <= 8'b00000000; // 7880 :   0 - 0x0
      13'h1EC9: dout <= 8'b00000000; // 7881 :   0 - 0x0
      13'h1ECA: dout <= 8'b00000000; // 7882 :   0 - 0x0
      13'h1ECB: dout <= 8'b00000000; // 7883 :   0 - 0x0
      13'h1ECC: dout <= 8'b00000100; // 7884 :   4 - 0x4
      13'h1ECD: dout <= 8'b00001110; // 7885 :  14 - 0xe
      13'h1ECE: dout <= 8'b00001111; // 7886 :  15 - 0xf
      13'h1ECF: dout <= 8'b00001011; // 7887 :  11 - 0xb
      13'h1ED0: dout <= 8'b00110000; // 7888 :  48 - 0x30 -- Background 0xed
      13'h1ED1: dout <= 8'b01000011; // 7889 :  67 - 0x43
      13'h1ED2: dout <= 8'b01000000; // 7890 :  64 - 0x40
      13'h1ED3: dout <= 8'b01100000; // 7891 :  96 - 0x60
      13'h1ED4: dout <= 8'b00000011; // 7892 :   3 - 0x3
      13'h1ED5: dout <= 8'b00000000; // 7893 :   0 - 0x0
      13'h1ED6: dout <= 8'b01111111; // 7894 : 127 - 0x7f
      13'h1ED7: dout <= 8'b00000000; // 7895 :   0 - 0x0
      13'h1ED8: dout <= 8'b00001111; // 7896 :  15 - 0xf
      13'h1ED9: dout <= 8'b00001100; // 7897 :  12 - 0xc
      13'h1EDA: dout <= 8'b00001111; // 7898 :  15 - 0xf
      13'h1EDB: dout <= 8'b00001111; // 7899 :  15 - 0xf
      13'h1EDC: dout <= 8'b00000000; // 7900 :   0 - 0x0
      13'h1EDD: dout <= 8'b01111111; // 7901 : 127 - 0x7f
      13'h1EDE: dout <= 8'b11010101; // 7902 : 213 - 0xd5
      13'h1EDF: dout <= 8'b01111111; // 7903 : 127 - 0x7f
      13'h1EE0: dout <= 8'b00000000; // 7904 :   0 - 0x0 -- Background 0xee
      13'h1EE1: dout <= 8'b00000000; // 7905 :   0 - 0x0
      13'h1EE2: dout <= 8'b00000000; // 7906 :   0 - 0x0
      13'h1EE3: dout <= 8'b00000000; // 7907 :   0 - 0x0
      13'h1EE4: dout <= 8'b00000000; // 7908 :   0 - 0x0
      13'h1EE5: dout <= 8'b00000000; // 7909 :   0 - 0x0
      13'h1EE6: dout <= 8'b00110000; // 7910 :  48 - 0x30
      13'h1EE7: dout <= 8'b00110000; // 7911 :  48 - 0x30
      13'h1EE8: dout <= 8'b00000000; // 7912 :   0 - 0x0
      13'h1EE9: dout <= 8'b00000000; // 7913 :   0 - 0x0
      13'h1EEA: dout <= 8'b00000000; // 7914 :   0 - 0x0
      13'h1EEB: dout <= 8'b00000000; // 7915 :   0 - 0x0
      13'h1EEC: dout <= 8'b00100000; // 7916 :  32 - 0x20
      13'h1EED: dout <= 8'b01110000; // 7917 : 112 - 0x70
      13'h1EEE: dout <= 8'b11110000; // 7918 : 240 - 0xf0
      13'h1EEF: dout <= 8'b11100000; // 7919 : 224 - 0xe0
      13'h1EF0: dout <= 8'b00001110; // 7920 :  14 - 0xe -- Background 0xef
      13'h1EF1: dout <= 8'b11001011; // 7921 : 203 - 0xcb
      13'h1EF2: dout <= 8'b00000000; // 7922 :   0 - 0x0
      13'h1EF3: dout <= 8'b00000000; // 7923 :   0 - 0x0
      13'h1EF4: dout <= 8'b11000000; // 7924 : 192 - 0xc0
      13'h1EF5: dout <= 8'b00000000; // 7925 :   0 - 0x0
      13'h1EF6: dout <= 8'b11111110; // 7926 : 254 - 0xfe
      13'h1EF7: dout <= 8'b00000000; // 7927 :   0 - 0x0
      13'h1EF8: dout <= 8'b11110000; // 7928 : 240 - 0xf0
      13'h1EF9: dout <= 8'b00110000; // 7929 :  48 - 0x30
      13'h1EFA: dout <= 8'b11110000; // 7930 : 240 - 0xf0
      13'h1EFB: dout <= 8'b11110000; // 7931 : 240 - 0xf0
      13'h1EFC: dout <= 8'b00000000; // 7932 :   0 - 0x0
      13'h1EFD: dout <= 8'b11111110; // 7933 : 254 - 0xfe
      13'h1EFE: dout <= 8'b01010101; // 7934 :  85 - 0x55
      13'h1EFF: dout <= 8'b11111110; // 7935 : 254 - 0xfe
      13'h1F00: dout <= 8'b00000000; // 7936 :   0 - 0x0 -- Background 0xf0
      13'h1F01: dout <= 8'b00000000; // 7937 :   0 - 0x0
      13'h1F02: dout <= 8'b00000000; // 7938 :   0 - 0x0
      13'h1F03: dout <= 8'b00000000; // 7939 :   0 - 0x0
      13'h1F04: dout <= 8'b00000000; // 7940 :   0 - 0x0
      13'h1F05: dout <= 8'b00000000; // 7941 :   0 - 0x0
      13'h1F06: dout <= 8'b00001100; // 7942 :  12 - 0xc
      13'h1F07: dout <= 8'b00001100; // 7943 :  12 - 0xc
      13'h1F08: dout <= 8'b00000000; // 7944 :   0 - 0x0
      13'h1F09: dout <= 8'b00000000; // 7945 :   0 - 0x0
      13'h1F0A: dout <= 8'b00000000; // 7946 :   0 - 0x0
      13'h1F0B: dout <= 8'b00000000; // 7947 :   0 - 0x0
      13'h1F0C: dout <= 8'b00000100; // 7948 :   4 - 0x4
      13'h1F0D: dout <= 8'b00001110; // 7949 :  14 - 0xe
      13'h1F0E: dout <= 8'b00001111; // 7950 :  15 - 0xf
      13'h1F0F: dout <= 8'b00001011; // 7951 :  11 - 0xb
      13'h1F10: dout <= 8'b00110000; // 7952 :  48 - 0x30 -- Background 0xf1
      13'h1F11: dout <= 8'b00100011; // 7953 :  35 - 0x23
      13'h1F12: dout <= 8'b00100000; // 7954 :  32 - 0x20
      13'h1F13: dout <= 8'b01100000; // 7955 :  96 - 0x60
      13'h1F14: dout <= 8'b00000011; // 7956 :   3 - 0x3
      13'h1F15: dout <= 8'b00000000; // 7957 :   0 - 0x0
      13'h1F16: dout <= 8'b01111111; // 7958 : 127 - 0x7f
      13'h1F17: dout <= 8'b00000000; // 7959 :   0 - 0x0
      13'h1F18: dout <= 8'b00001111; // 7960 :  15 - 0xf
      13'h1F19: dout <= 8'b00001100; // 7961 :  12 - 0xc
      13'h1F1A: dout <= 8'b00001111; // 7962 :  15 - 0xf
      13'h1F1B: dout <= 8'b00001111; // 7963 :  15 - 0xf
      13'h1F1C: dout <= 8'b00000000; // 7964 :   0 - 0x0
      13'h1F1D: dout <= 8'b01111111; // 7965 : 127 - 0x7f
      13'h1F1E: dout <= 8'b10101010; // 7966 : 170 - 0xaa
      13'h1F1F: dout <= 8'b01111111; // 7967 : 127 - 0x7f
      13'h1F20: dout <= 8'b00000000; // 7968 :   0 - 0x0 -- Background 0xf2
      13'h1F21: dout <= 8'b00000000; // 7969 :   0 - 0x0
      13'h1F22: dout <= 8'b00000000; // 7970 :   0 - 0x0
      13'h1F23: dout <= 8'b00000000; // 7971 :   0 - 0x0
      13'h1F24: dout <= 8'b00000000; // 7972 :   0 - 0x0
      13'h1F25: dout <= 8'b00000000; // 7973 :   0 - 0x0
      13'h1F26: dout <= 8'b00110000; // 7974 :  48 - 0x30
      13'h1F27: dout <= 8'b00110000; // 7975 :  48 - 0x30
      13'h1F28: dout <= 8'b00000000; // 7976 :   0 - 0x0
      13'h1F29: dout <= 8'b00000000; // 7977 :   0 - 0x0
      13'h1F2A: dout <= 8'b00000000; // 7978 :   0 - 0x0
      13'h1F2B: dout <= 8'b00000000; // 7979 :   0 - 0x0
      13'h1F2C: dout <= 8'b00100000; // 7980 :  32 - 0x20
      13'h1F2D: dout <= 8'b01110000; // 7981 : 112 - 0x70
      13'h1F2E: dout <= 8'b11110000; // 7982 : 240 - 0xf0
      13'h1F2F: dout <= 8'b11100000; // 7983 : 224 - 0xe0
      13'h1F30: dout <= 8'b00001001; // 7984 :   9 - 0x9 -- Background 0xf3
      13'h1F31: dout <= 8'b11001111; // 7985 : 207 - 0xcf
      13'h1F32: dout <= 8'b00000000; // 7986 :   0 - 0x0
      13'h1F33: dout <= 8'b00000000; // 7987 :   0 - 0x0
      13'h1F34: dout <= 8'b11000000; // 7988 : 192 - 0xc0
      13'h1F35: dout <= 8'b00000000; // 7989 :   0 - 0x0
      13'h1F36: dout <= 8'b11111110; // 7990 : 254 - 0xfe
      13'h1F37: dout <= 8'b00000000; // 7991 :   0 - 0x0
      13'h1F38: dout <= 8'b11110000; // 7992 : 240 - 0xf0
      13'h1F39: dout <= 8'b00110000; // 7993 :  48 - 0x30
      13'h1F3A: dout <= 8'b11110000; // 7994 : 240 - 0xf0
      13'h1F3B: dout <= 8'b11110000; // 7995 : 240 - 0xf0
      13'h1F3C: dout <= 8'b00000000; // 7996 :   0 - 0x0
      13'h1F3D: dout <= 8'b11111110; // 7997 : 254 - 0xfe
      13'h1F3E: dout <= 8'b10101011; // 7998 : 171 - 0xab
      13'h1F3F: dout <= 8'b11111110; // 7999 : 254 - 0xfe
      13'h1F40: dout <= 8'b00111111; // 8000 :  63 - 0x3f -- Background 0xf4
      13'h1F41: dout <= 8'b00110101; // 8001 :  53 - 0x35
      13'h1F42: dout <= 8'b00011010; // 8002 :  26 - 0x1a
      13'h1F43: dout <= 8'b00001101; // 8003 :  13 - 0xd
      13'h1F44: dout <= 8'b00001010; // 8004 :  10 - 0xa
      13'h1F45: dout <= 8'b00001101; // 8005 :  13 - 0xd
      13'h1F46: dout <= 8'b00001000; // 8006 :   8 - 0x8
      13'h1F47: dout <= 8'b00111000; // 8007 :  56 - 0x38
      13'h1F48: dout <= 8'b00000000; // 8008 :   0 - 0x0
      13'h1F49: dout <= 8'b00010101; // 8009 :  21 - 0x15
      13'h1F4A: dout <= 8'b00001010; // 8010 :  10 - 0xa
      13'h1F4B: dout <= 8'b00000101; // 8011 :   5 - 0x5
      13'h1F4C: dout <= 8'b00000010; // 8012 :   2 - 0x2
      13'h1F4D: dout <= 8'b00000101; // 8013 :   5 - 0x5
      13'h1F4E: dout <= 8'b00000111; // 8014 :   7 - 0x7
      13'h1F4F: dout <= 8'b00000111; // 8015 :   7 - 0x7
      13'h1F50: dout <= 8'b01110011; // 8016 : 115 - 0x73 -- Background 0xf5
      13'h1F51: dout <= 8'b11000100; // 8017 : 196 - 0xc4
      13'h1F52: dout <= 8'b11000100; // 8018 : 196 - 0xc4
      13'h1F53: dout <= 8'b11000000; // 8019 : 192 - 0xc0
      13'h1F54: dout <= 8'b11000001; // 8020 : 193 - 0xc1
      13'h1F55: dout <= 8'b11000000; // 8021 : 192 - 0xc0
      13'h1F56: dout <= 8'b01100001; // 8022 :  97 - 0x61
      13'h1F57: dout <= 8'b00111111; // 8023 :  63 - 0x3f
      13'h1F58: dout <= 8'b00111100; // 8024 :  60 - 0x3c
      13'h1F59: dout <= 8'b01111011; // 8025 : 123 - 0x7b
      13'h1F5A: dout <= 8'b01111011; // 8026 : 123 - 0x7b
      13'h1F5B: dout <= 8'b01111111; // 8027 : 127 - 0x7f
      13'h1F5C: dout <= 8'b01111110; // 8028 : 126 - 0x7e
      13'h1F5D: dout <= 8'b01111111; // 8029 : 127 - 0x7f
      13'h1F5E: dout <= 8'b00111110; // 8030 :  62 - 0x3e
      13'h1F5F: dout <= 8'b00000000; // 8031 :   0 - 0x0
      13'h1F60: dout <= 8'b11111100; // 8032 : 252 - 0xfc -- Background 0xf6
      13'h1F61: dout <= 8'b01010100; // 8033 :  84 - 0x54
      13'h1F62: dout <= 8'b10101000; // 8034 : 168 - 0xa8
      13'h1F63: dout <= 8'b01010000; // 8035 :  80 - 0x50
      13'h1F64: dout <= 8'b10110000; // 8036 : 176 - 0xb0
      13'h1F65: dout <= 8'b01010000; // 8037 :  80 - 0x50
      13'h1F66: dout <= 8'b10010000; // 8038 : 144 - 0x90
      13'h1F67: dout <= 8'b00011100; // 8039 :  28 - 0x1c
      13'h1F68: dout <= 8'b00000000; // 8040 :   0 - 0x0
      13'h1F69: dout <= 8'b01010000; // 8041 :  80 - 0x50
      13'h1F6A: dout <= 8'b10100000; // 8042 : 160 - 0xa0
      13'h1F6B: dout <= 8'b01000000; // 8043 :  64 - 0x40
      13'h1F6C: dout <= 8'b10100000; // 8044 : 160 - 0xa0
      13'h1F6D: dout <= 8'b01000000; // 8045 :  64 - 0x40
      13'h1F6E: dout <= 8'b11100000; // 8046 : 224 - 0xe0
      13'h1F6F: dout <= 8'b11100000; // 8047 : 224 - 0xe0
      13'h1F70: dout <= 8'b10000110; // 8048 : 134 - 0x86 -- Background 0xf7
      13'h1F71: dout <= 8'b01000010; // 8049 :  66 - 0x42
      13'h1F72: dout <= 8'b01000111; // 8050 :  71 - 0x47
      13'h1F73: dout <= 8'b01000001; // 8051 :  65 - 0x41
      13'h1F74: dout <= 8'b10000011; // 8052 : 131 - 0x83
      13'h1F75: dout <= 8'b00000001; // 8053 :   1 - 0x1
      13'h1F76: dout <= 8'b10000110; // 8054 : 134 - 0x86
      13'h1F77: dout <= 8'b11111100; // 8055 : 252 - 0xfc
      13'h1F78: dout <= 8'b01111000; // 8056 : 120 - 0x78
      13'h1F79: dout <= 8'b10111100; // 8057 : 188 - 0xbc
      13'h1F7A: dout <= 8'b10111000; // 8058 : 184 - 0xb8
      13'h1F7B: dout <= 8'b10111110; // 8059 : 190 - 0xbe
      13'h1F7C: dout <= 8'b01111100; // 8060 : 124 - 0x7c
      13'h1F7D: dout <= 8'b11111110; // 8061 : 254 - 0xfe
      13'h1F7E: dout <= 8'b01111000; // 8062 : 120 - 0x78
      13'h1F7F: dout <= 8'b00000000; // 8063 :   0 - 0x0
      13'h1F80: dout <= 8'b11100100; // 8064 : 228 - 0xe4 -- Background 0xf8
      13'h1F81: dout <= 8'b11100100; // 8065 : 228 - 0xe4
      13'h1F82: dout <= 8'b11101111; // 8066 : 239 - 0xef
      13'h1F83: dout <= 8'b11101111; // 8067 : 239 - 0xef
      13'h1F84: dout <= 8'b11111111; // 8068 : 255 - 0xff
      13'h1F85: dout <= 8'b11111111; // 8069 : 255 - 0xff
      13'h1F86: dout <= 8'b01111111; // 8070 : 127 - 0x7f
      13'h1F87: dout <= 8'b01111111; // 8071 : 127 - 0x7f
      13'h1F88: dout <= 8'b00000011; // 8072 :   3 - 0x3
      13'h1F89: dout <= 8'b00000011; // 8073 :   3 - 0x3
      13'h1F8A: dout <= 8'b00000000; // 8074 :   0 - 0x0
      13'h1F8B: dout <= 8'b00000011; // 8075 :   3 - 0x3
      13'h1F8C: dout <= 8'b00000111; // 8076 :   7 - 0x7
      13'h1F8D: dout <= 8'b00000110; // 8077 :   6 - 0x6
      13'h1F8E: dout <= 8'b00000111; // 8078 :   7 - 0x7
      13'h1F8F: dout <= 8'b00000000; // 8079 :   0 - 0x0
      13'h1F90: dout <= 8'b00111111; // 8080 :  63 - 0x3f -- Background 0xf9
      13'h1F91: dout <= 8'b01111111; // 8081 : 127 - 0x7f
      13'h1F92: dout <= 8'b01111111; // 8082 : 127 - 0x7f
      13'h1F93: dout <= 8'b11111111; // 8083 : 255 - 0xff
      13'h1F94: dout <= 8'b11111111; // 8084 : 255 - 0xff
      13'h1F95: dout <= 8'b11111111; // 8085 : 255 - 0xff
      13'h1F96: dout <= 8'b11111111; // 8086 : 255 - 0xff
      13'h1F97: dout <= 8'b11111111; // 8087 : 255 - 0xff
      13'h1F98: dout <= 8'b00000000; // 8088 :   0 - 0x0
      13'h1F99: dout <= 8'b00011111; // 8089 :  31 - 0x1f
      13'h1F9A: dout <= 8'b00011111; // 8090 :  31 - 0x1f
      13'h1F9B: dout <= 8'b00001111; // 8091 :  15 - 0xf
      13'h1F9C: dout <= 8'b00000011; // 8092 :   3 - 0x3
      13'h1F9D: dout <= 8'b00000000; // 8093 :   0 - 0x0
      13'h1F9E: dout <= 8'b00000000; // 8094 :   0 - 0x0
      13'h1F9F: dout <= 8'b00000000; // 8095 :   0 - 0x0
      13'h1FA0: dout <= 8'b00010011; // 8096 :  19 - 0x13 -- Background 0xfa
      13'h1FA1: dout <= 8'b00010011; // 8097 :  19 - 0x13
      13'h1FA2: dout <= 8'b11111011; // 8098 : 251 - 0xfb
      13'h1FA3: dout <= 8'b11111011; // 8099 : 251 - 0xfb
      13'h1FA4: dout <= 8'b11111111; // 8100 : 255 - 0xff
      13'h1FA5: dout <= 8'b11111111; // 8101 : 255 - 0xff
      13'h1FA6: dout <= 8'b11111110; // 8102 : 254 - 0xfe
      13'h1FA7: dout <= 8'b11111110; // 8103 : 254 - 0xfe
      13'h1FA8: dout <= 8'b11100000; // 8104 : 224 - 0xe0
      13'h1FA9: dout <= 8'b11100000; // 8105 : 224 - 0xe0
      13'h1FAA: dout <= 8'b00000000; // 8106 :   0 - 0x0
      13'h1FAB: dout <= 8'b00110000; // 8107 :  48 - 0x30
      13'h1FAC: dout <= 8'b01110000; // 8108 : 112 - 0x70
      13'h1FAD: dout <= 8'b01100000; // 8109 :  96 - 0x60
      13'h1FAE: dout <= 8'b01110000; // 8110 : 112 - 0x70
      13'h1FAF: dout <= 8'b00000000; // 8111 :   0 - 0x0
      13'h1FB0: dout <= 8'b11111110; // 8112 : 254 - 0xfe -- Background 0xfb
      13'h1FB1: dout <= 8'b11111111; // 8113 : 255 - 0xff
      13'h1FB2: dout <= 8'b11111111; // 8114 : 255 - 0xff
      13'h1FB3: dout <= 8'b11111111; // 8115 : 255 - 0xff
      13'h1FB4: dout <= 8'b11111111; // 8116 : 255 - 0xff
      13'h1FB5: dout <= 8'b11111111; // 8117 : 255 - 0xff
      13'h1FB6: dout <= 8'b11111111; // 8118 : 255 - 0xff
      13'h1FB7: dout <= 8'b11111111; // 8119 : 255 - 0xff
      13'h1FB8: dout <= 8'b00000000; // 8120 :   0 - 0x0
      13'h1FB9: dout <= 8'b11111000; // 8121 : 248 - 0xf8
      13'h1FBA: dout <= 8'b11111000; // 8122 : 248 - 0xf8
      13'h1FBB: dout <= 8'b11110000; // 8123 : 240 - 0xf0
      13'h1FBC: dout <= 8'b11000000; // 8124 : 192 - 0xc0
      13'h1FBD: dout <= 8'b00000000; // 8125 :   0 - 0x0
      13'h1FBE: dout <= 8'b00000000; // 8126 :   0 - 0x0
      13'h1FBF: dout <= 8'b00000000; // 8127 :   0 - 0x0
      13'h1FC0: dout <= 8'b00000000; // 8128 :   0 - 0x0 -- Background 0xfc
      13'h1FC1: dout <= 8'b00000000; // 8129 :   0 - 0x0
      13'h1FC2: dout <= 8'b01111100; // 8130 : 124 - 0x7c
      13'h1FC3: dout <= 8'b11111110; // 8131 : 254 - 0xfe
      13'h1FC4: dout <= 8'b11111110; // 8132 : 254 - 0xfe
      13'h1FC5: dout <= 8'b01111100; // 8133 : 124 - 0x7c
      13'h1FC6: dout <= 8'b01000100; // 8134 :  68 - 0x44
      13'h1FC7: dout <= 8'b10000010; // 8135 : 130 - 0x82
      13'h1FC8: dout <= 8'b00111000; // 8136 :  56 - 0x38
      13'h1FC9: dout <= 8'b00111000; // 8137 :  56 - 0x38
      13'h1FCA: dout <= 8'b00000000; // 8138 :   0 - 0x0
      13'h1FCB: dout <= 8'b01111100; // 8139 : 124 - 0x7c
      13'h1FCC: dout <= 8'b00000000; // 8140 :   0 - 0x0
      13'h1FCD: dout <= 8'b00111000; // 8141 :  56 - 0x38
      13'h1FCE: dout <= 8'b00111000; // 8142 :  56 - 0x38
      13'h1FCF: dout <= 8'b01111100; // 8143 : 124 - 0x7c
      13'h1FD0: dout <= 8'b10000010; // 8144 : 130 - 0x82 -- Background 0xfd
      13'h1FD1: dout <= 8'b10000010; // 8145 : 130 - 0x82
      13'h1FD2: dout <= 8'b10000010; // 8146 : 130 - 0x82
      13'h1FD3: dout <= 8'b11000110; // 8147 : 198 - 0xc6
      13'h1FD4: dout <= 8'b11111110; // 8148 : 254 - 0xfe
      13'h1FD5: dout <= 8'b11111110; // 8149 : 254 - 0xfe
      13'h1FD6: dout <= 8'b10111010; // 8150 : 186 - 0xba
      13'h1FD7: dout <= 8'b01111100; // 8151 : 124 - 0x7c
      13'h1FD8: dout <= 8'b01111100; // 8152 : 124 - 0x7c
      13'h1FD9: dout <= 8'b01111100; // 8153 : 124 - 0x7c
      13'h1FDA: dout <= 8'b01111100; // 8154 : 124 - 0x7c
      13'h1FDB: dout <= 8'b00111000; // 8155 :  56 - 0x38
      13'h1FDC: dout <= 8'b00000000; // 8156 :   0 - 0x0
      13'h1FDD: dout <= 8'b01111100; // 8157 : 124 - 0x7c
      13'h1FDE: dout <= 8'b01111100; // 8158 : 124 - 0x7c
      13'h1FDF: dout <= 8'b00000000; // 8159 :   0 - 0x0
      13'h1FE0: dout <= 8'b00000000; // 8160 :   0 - 0x0 -- Background 0xfe
      13'h1FE1: dout <= 8'b00011001; // 8161 :  25 - 0x19
      13'h1FE2: dout <= 8'b00111110; // 8162 :  62 - 0x3e
      13'h1FE3: dout <= 8'b00111100; // 8163 :  60 - 0x3c
      13'h1FE4: dout <= 8'b00111100; // 8164 :  60 - 0x3c
      13'h1FE5: dout <= 8'b00111100; // 8165 :  60 - 0x3c
      13'h1FE6: dout <= 8'b00111110; // 8166 :  62 - 0x3e
      13'h1FE7: dout <= 8'b00011001; // 8167 :  25 - 0x19
      13'h1FE8: dout <= 8'b00000000; // 8168 :   0 - 0x0
      13'h1FE9: dout <= 8'b00000000; // 8169 :   0 - 0x0
      13'h1FEA: dout <= 8'b00010001; // 8170 :  17 - 0x11
      13'h1FEB: dout <= 8'b11010111; // 8171 : 215 - 0xd7
      13'h1FEC: dout <= 8'b11010111; // 8172 : 215 - 0xd7
      13'h1FED: dout <= 8'b11010111; // 8173 : 215 - 0xd7
      13'h1FEE: dout <= 8'b00010001; // 8174 :  17 - 0x11
      13'h1FEF: dout <= 8'b00000000; // 8175 :   0 - 0x0
      13'h1FF0: dout <= 8'b00000000; // 8176 :   0 - 0x0 -- Background 0xff
      13'h1FF1: dout <= 8'b11111110; // 8177 : 254 - 0xfe
      13'h1FF2: dout <= 8'b00011101; // 8178 :  29 - 0x1d
      13'h1FF3: dout <= 8'b00001111; // 8179 :  15 - 0xf
      13'h1FF4: dout <= 8'b00001111; // 8180 :  15 - 0xf
      13'h1FF5: dout <= 8'b00001111; // 8181 :  15 - 0xf
      13'h1FF6: dout <= 8'b00011101; // 8182 :  29 - 0x1d
      13'h1FF7: dout <= 8'b11111110; // 8183 : 254 - 0xfe
      13'h1FF8: dout <= 8'b00000000; // 8184 :   0 - 0x0
      13'h1FF9: dout <= 8'b00000000; // 8185 :   0 - 0x0
      13'h1FFA: dout <= 8'b11100110; // 8186 : 230 - 0xe6
      13'h1FFB: dout <= 8'b11110110; // 8187 : 246 - 0xf6
      13'h1FFC: dout <= 8'b11110110; // 8188 : 246 - 0xf6
      13'h1FFD: dout <= 8'b11110110; // 8189 : 246 - 0xf6
      13'h1FFE: dout <= 8'b11100110; // 8190 : 230 - 0xe6
      13'h1FFF: dout <= 8'b00000000; // 8191 :   0 - 0x0
    endcase
  end

endmodule
