//- Autcmatically generated verilog ROM from a NES memory file----
//-   NAME TABLE
// https://wiki.nesdev.com/w/index.php/PPU_nametables
//- Only the first Name Table: 1KiB


//-  Original memory dump file name: pacman_ntable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_NTABLE_PACMAN_00
  (
     //input     clk,   // clock
     input      [10-1:0] addr,  //1024 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
     //----- Name Table 0---------
      10'h0: dout  = 8'b00100000; //    0 :  32 - 0x20 -- line 0x0
      10'h1: dout  = 8'b00100000; //    1 :  32 - 0x20
      10'h2: dout  = 8'b00100000; //    2 :  32 - 0x20
      10'h3: dout  = 8'b00100000; //    3 :  32 - 0x20
      10'h4: dout  = 8'b00100000; //    4 :  32 - 0x20
      10'h5: dout  = 8'b00100000; //    5 :  32 - 0x20
      10'h6: dout  = 8'b00100000; //    6 :  32 - 0x20
      10'h7: dout  = 8'b00100000; //    7 :  32 - 0x20
      10'h8: dout  = 8'b00100000; //    8 :  32 - 0x20
      10'h9: dout  = 8'b00100000; //    9 :  32 - 0x20
      10'hA: dout  = 8'b00100000; //   10 :  32 - 0x20
      10'hB: dout  = 8'b00100000; //   11 :  32 - 0x20
      10'hC: dout  = 8'b00100000; //   12 :  32 - 0x20
      10'hD: dout  = 8'b00100000; //   13 :  32 - 0x20
      10'hE: dout  = 8'b00100000; //   14 :  32 - 0x20
      10'hF: dout  = 8'b00100000; //   15 :  32 - 0x20
      10'h10: dout  = 8'b00100000; //   16 :  32 - 0x20
      10'h11: dout  = 8'b00100000; //   17 :  32 - 0x20
      10'h12: dout  = 8'b00100000; //   18 :  32 - 0x20
      10'h13: dout  = 8'b00100000; //   19 :  32 - 0x20
      10'h14: dout  = 8'b00100000; //   20 :  32 - 0x20
      10'h15: dout  = 8'b00100000; //   21 :  32 - 0x20
      10'h16: dout  = 8'b00100000; //   22 :  32 - 0x20
      10'h17: dout  = 8'b00100000; //   23 :  32 - 0x20
      10'h18: dout  = 8'b00100000; //   24 :  32 - 0x20
      10'h19: dout  = 8'b00100000; //   25 :  32 - 0x20
      10'h1A: dout  = 8'b00100000; //   26 :  32 - 0x20
      10'h1B: dout  = 8'b00100000; //   27 :  32 - 0x20
      10'h1C: dout  = 8'b00100000; //   28 :  32 - 0x20
      10'h1D: dout  = 8'b00100000; //   29 :  32 - 0x20
      10'h1E: dout  = 8'b00100000; //   30 :  32 - 0x20
      10'h1F: dout  = 8'b00100000; //   31 :  32 - 0x20
      10'h20: dout  = 8'b00100000; //   32 :  32 - 0x20 -- line 0x1
      10'h21: dout  = 8'b00100000; //   33 :  32 - 0x20
      10'h22: dout  = 8'b00100000; //   34 :  32 - 0x20
      10'h23: dout  = 8'b00100000; //   35 :  32 - 0x20
      10'h24: dout  = 8'b00100000; //   36 :  32 - 0x20
      10'h25: dout  = 8'b00100000; //   37 :  32 - 0x20
      10'h26: dout  = 8'b00100000; //   38 :  32 - 0x20
      10'h27: dout  = 8'b00100000; //   39 :  32 - 0x20
      10'h28: dout  = 8'b00100000; //   40 :  32 - 0x20
      10'h29: dout  = 8'b00100000; //   41 :  32 - 0x20
      10'h2A: dout  = 8'b00100000; //   42 :  32 - 0x20
      10'h2B: dout  = 8'b00100000; //   43 :  32 - 0x20
      10'h2C: dout  = 8'b00100000; //   44 :  32 - 0x20
      10'h2D: dout  = 8'b00100000; //   45 :  32 - 0x20
      10'h2E: dout  = 8'b00100000; //   46 :  32 - 0x20
      10'h2F: dout  = 8'b00100000; //   47 :  32 - 0x20
      10'h30: dout  = 8'b00100000; //   48 :  32 - 0x20
      10'h31: dout  = 8'b00100000; //   49 :  32 - 0x20
      10'h32: dout  = 8'b00100000; //   50 :  32 - 0x20
      10'h33: dout  = 8'b00100000; //   51 :  32 - 0x20
      10'h34: dout  = 8'b00100000; //   52 :  32 - 0x20
      10'h35: dout  = 8'b00100000; //   53 :  32 - 0x20
      10'h36: dout  = 8'b00100000; //   54 :  32 - 0x20
      10'h37: dout  = 8'b00100000; //   55 :  32 - 0x20
      10'h38: dout  = 8'b00100000; //   56 :  32 - 0x20
      10'h39: dout  = 8'b00100000; //   57 :  32 - 0x20
      10'h3A: dout  = 8'b00100000; //   58 :  32 - 0x20
      10'h3B: dout  = 8'b00100000; //   59 :  32 - 0x20
      10'h3C: dout  = 8'b00100000; //   60 :  32 - 0x20
      10'h3D: dout  = 8'b00100000; //   61 :  32 - 0x20
      10'h3E: dout  = 8'b00100000; //   62 :  32 - 0x20
      10'h3F: dout  = 8'b00100000; //   63 :  32 - 0x20
      10'h40: dout  = 8'b00101101; //   64 :  45 - 0x2d -- line 0x2
      10'h41: dout  = 8'b00011111; //   65 :  31 - 0x1f
      10'h42: dout  = 8'b00010000; //   66 :  16 - 0x10
      10'h43: dout  = 8'b00010000; //   67 :  16 - 0x10
      10'h44: dout  = 8'b00010000; //   68 :  16 - 0x10
      10'h45: dout  = 8'b00010000; //   69 :  16 - 0x10
      10'h46: dout  = 8'b00010000; //   70 :  16 - 0x10
      10'h47: dout  = 8'b00010000; //   71 :  16 - 0x10
      10'h48: dout  = 8'b00010000; //   72 :  16 - 0x10
      10'h49: dout  = 8'b00010000; //   73 :  16 - 0x10
      10'h4A: dout  = 8'b00010000; //   74 :  16 - 0x10
      10'h4B: dout  = 8'b00010011; //   75 :  19 - 0x13
      10'h4C: dout  = 8'b00010000; //   76 :  16 - 0x10
      10'h4D: dout  = 8'b00010000; //   77 :  16 - 0x10
      10'h4E: dout  = 8'b00010000; //   78 :  16 - 0x10
      10'h4F: dout  = 8'b00010000; //   79 :  16 - 0x10
      10'h50: dout  = 8'b00010000; //   80 :  16 - 0x10
      10'h51: dout  = 8'b00010000; //   81 :  16 - 0x10
      10'h52: dout  = 8'b00010000; //   82 :  16 - 0x10
      10'h53: dout  = 8'b00010000; //   83 :  16 - 0x10
      10'h54: dout  = 8'b00010000; //   84 :  16 - 0x10
      10'h55: dout  = 8'b00011101; //   85 :  29 - 0x1d
      10'h56: dout  = 8'b00100000; //   86 :  32 - 0x20
      10'h57: dout  = 8'b00100000; //   87 :  32 - 0x20
      10'h58: dout  = 8'b00100000; //   88 :  32 - 0x20
      10'h59: dout  = 8'b00100000; //   89 :  32 - 0x20
      10'h5A: dout  = 8'b00100000; //   90 :  32 - 0x20
      10'h5B: dout  = 8'b00100000; //   91 :  32 - 0x20
      10'h5C: dout  = 8'b00100000; //   92 :  32 - 0x20
      10'h5D: dout  = 8'b00100000; //   93 :  32 - 0x20
      10'h5E: dout  = 8'b00100000; //   94 :  32 - 0x20
      10'h5F: dout  = 8'b00100000; //   95 :  32 - 0x20
      10'h60: dout  = 8'b00101101; //   96 :  45 - 0x2d -- line 0x3
      10'h61: dout  = 8'b00010001; //   97 :  17 - 0x11
      10'h62: dout  = 8'b00000011; //   98 :   3 - 0x3
      10'h63: dout  = 8'b00000011; //   99 :   3 - 0x3
      10'h64: dout  = 8'b00000011; //  100 :   3 - 0x3
      10'h65: dout  = 8'b00000011; //  101 :   3 - 0x3
      10'h66: dout  = 8'b00000011; //  102 :   3 - 0x3
      10'h67: dout  = 8'b00000011; //  103 :   3 - 0x3
      10'h68: dout  = 8'b00000011; //  104 :   3 - 0x3
      10'h69: dout  = 8'b00000011; //  105 :   3 - 0x3
      10'h6A: dout  = 8'b00000011; //  106 :   3 - 0x3
      10'h6B: dout  = 8'b00010001; //  107 :  17 - 0x11
      10'h6C: dout  = 8'b00000011; //  108 :   3 - 0x3
      10'h6D: dout  = 8'b00000011; //  109 :   3 - 0x3
      10'h6E: dout  = 8'b00000011; //  110 :   3 - 0x3
      10'h6F: dout  = 8'b00000011; //  111 :   3 - 0x3
      10'h70: dout  = 8'b00000011; //  112 :   3 - 0x3
      10'h71: dout  = 8'b00000011; //  113 :   3 - 0x3
      10'h72: dout  = 8'b00000011; //  114 :   3 - 0x3
      10'h73: dout  = 8'b00000011; //  115 :   3 - 0x3
      10'h74: dout  = 8'b00000011; //  116 :   3 - 0x3
      10'h75: dout  = 8'b00010001; //  117 :  17 - 0x11
      10'h76: dout  = 8'b10110100; //  118 : 180 - 0xb4
      10'h77: dout  = 8'b10110101; //  119 : 181 - 0xb5
      10'h78: dout  = 8'b10110110; //  120 : 182 - 0xb6
      10'h79: dout  = 8'b10110111; //  121 : 183 - 0xb7
      10'h7A: dout  = 8'b10111000; //  122 : 184 - 0xb8
      10'h7B: dout  = 8'b10111001; //  123 : 185 - 0xb9
      10'h7C: dout  = 8'b10111010; //  124 : 186 - 0xba
      10'h7D: dout  = 8'b10111011; //  125 : 187 - 0xbb
      10'h7E: dout  = 8'b00100000; //  126 :  32 - 0x20
      10'h7F: dout  = 8'b00100000; //  127 :  32 - 0x20
      10'h80: dout  = 8'b00101101; //  128 :  45 - 0x2d -- line 0x4
      10'h81: dout  = 8'b00010001; //  129 :  17 - 0x11
      10'h82: dout  = 8'b00000011; //  130 :   3 - 0x3
      10'h83: dout  = 8'b00011111; //  131 :  31 - 0x1f
      10'h84: dout  = 8'b00010000; //  132 :  16 - 0x10
      10'h85: dout  = 8'b00011101; //  133 :  29 - 0x1d
      10'h86: dout  = 8'b00000011; //  134 :   3 - 0x3
      10'h87: dout  = 8'b00011111; //  135 :  31 - 0x1f
      10'h88: dout  = 8'b00010000; //  136 :  16 - 0x10
      10'h89: dout  = 8'b00011101; //  137 :  29 - 0x1d
      10'h8A: dout  = 8'b00000011; //  138 :   3 - 0x3
      10'h8B: dout  = 8'b00010001; //  139 :  17 - 0x11
      10'h8C: dout  = 8'b00000011; //  140 :   3 - 0x3
      10'h8D: dout  = 8'b00011111; //  141 :  31 - 0x1f
      10'h8E: dout  = 8'b00010000; //  142 :  16 - 0x10
      10'h8F: dout  = 8'b00011101; //  143 :  29 - 0x1d
      10'h90: dout  = 8'b00000011; //  144 :   3 - 0x3
      10'h91: dout  = 8'b00011111; //  145 :  31 - 0x1f
      10'h92: dout  = 8'b00010000; //  146 :  16 - 0x10
      10'h93: dout  = 8'b00011101; //  147 :  29 - 0x1d
      10'h94: dout  = 8'b00000011; //  148 :   3 - 0x3
      10'h95: dout  = 8'b00010001; //  149 :  17 - 0x11
      10'h96: dout  = 8'b00100000; //  150 :  32 - 0x20
      10'h97: dout  = 8'b00100000; //  151 :  32 - 0x20
      10'h98: dout  = 8'b00100000; //  152 :  32 - 0x20
      10'h99: dout  = 8'b00100000; //  153 :  32 - 0x20
      10'h9A: dout  = 8'b00100000; //  154 :  32 - 0x20
      10'h9B: dout  = 8'b00100000; //  155 :  32 - 0x20
      10'h9C: dout  = 8'b00100000; //  156 :  32 - 0x20
      10'h9D: dout  = 8'b00100000; //  157 :  32 - 0x20
      10'h9E: dout  = 8'b00100000; //  158 :  32 - 0x20
      10'h9F: dout  = 8'b00100000; //  159 :  32 - 0x20
      10'hA0: dout  = 8'b00101101; //  160 :  45 - 0x2d -- line 0x5
      10'hA1: dout  = 8'b00010001; //  161 :  17 - 0x11
      10'hA2: dout  = 8'b00000001; //  162 :   1 - 0x1
      10'hA3: dout  = 8'b00010001; //  163 :  17 - 0x11
      10'hA4: dout  = 8'b00100000; //  164 :  32 - 0x20
      10'hA5: dout  = 8'b00010001; //  165 :  17 - 0x11
      10'hA6: dout  = 8'b00000011; //  166 :   3 - 0x3
      10'hA7: dout  = 8'b00010001; //  167 :  17 - 0x11
      10'hA8: dout  = 8'b00100000; //  168 :  32 - 0x20
      10'hA9: dout  = 8'b00010001; //  169 :  17 - 0x11
      10'hAA: dout  = 8'b00000011; //  170 :   3 - 0x3
      10'hAB: dout  = 8'b00010001; //  171 :  17 - 0x11
      10'hAC: dout  = 8'b00000011; //  172 :   3 - 0x3
      10'hAD: dout  = 8'b00010001; //  173 :  17 - 0x11
      10'hAE: dout  = 8'b00100000; //  174 :  32 - 0x20
      10'hAF: dout  = 8'b00010001; //  175 :  17 - 0x11
      10'hB0: dout  = 8'b00000011; //  176 :   3 - 0x3
      10'hB1: dout  = 8'b00010001; //  177 :  17 - 0x11
      10'hB2: dout  = 8'b00100000; //  178 :  32 - 0x20
      10'hB3: dout  = 8'b00010001; //  179 :  17 - 0x11
      10'hB4: dout  = 8'b00000001; //  180 :   1 - 0x1
      10'hB5: dout  = 8'b00010001; //  181 :  17 - 0x11
      10'hB6: dout  = 8'b00100000; //  182 :  32 - 0x20
      10'hB7: dout  = 8'b00100000; //  183 :  32 - 0x20
      10'hB8: dout  = 8'b00110001; //  184 :  49 - 0x31
      10'hB9: dout  = 8'b00110000; //  185 :  48 - 0x30
      10'hBA: dout  = 8'b00110000; //  186 :  48 - 0x30
      10'hBB: dout  = 8'b00110000; //  187 :  48 - 0x30
      10'hBC: dout  = 8'b00110000; //  188 :  48 - 0x30
      10'hBD: dout  = 8'b00100000; //  189 :  32 - 0x20
      10'hBE: dout  = 8'b00100000; //  190 :  32 - 0x20
      10'hBF: dout  = 8'b00100000; //  191 :  32 - 0x20
      10'hC0: dout  = 8'b00101101; //  192 :  45 - 0x2d -- line 0x6
      10'hC1: dout  = 8'b00010001; //  193 :  17 - 0x11
      10'hC2: dout  = 8'b00000011; //  194 :   3 - 0x3
      10'hC3: dout  = 8'b00011110; //  195 :  30 - 0x1e
      10'hC4: dout  = 8'b00010000; //  196 :  16 - 0x10
      10'hC5: dout  = 8'b00011100; //  197 :  28 - 0x1c
      10'hC6: dout  = 8'b00000011; //  198 :   3 - 0x3
      10'hC7: dout  = 8'b00011110; //  199 :  30 - 0x1e
      10'hC8: dout  = 8'b00010000; //  200 :  16 - 0x10
      10'hC9: dout  = 8'b00011100; //  201 :  28 - 0x1c
      10'hCA: dout  = 8'b00000011; //  202 :   3 - 0x3
      10'hCB: dout  = 8'b00011010; //  203 :  26 - 0x1a
      10'hCC: dout  = 8'b00000011; //  204 :   3 - 0x3
      10'hCD: dout  = 8'b00011110; //  205 :  30 - 0x1e
      10'hCE: dout  = 8'b00010000; //  206 :  16 - 0x10
      10'hCF: dout  = 8'b00011100; //  207 :  28 - 0x1c
      10'hD0: dout  = 8'b00000011; //  208 :   3 - 0x3
      10'hD1: dout  = 8'b00011110; //  209 :  30 - 0x1e
      10'hD2: dout  = 8'b00010000; //  210 :  16 - 0x10
      10'hD3: dout  = 8'b00011100; //  211 :  28 - 0x1c
      10'hD4: dout  = 8'b00000011; //  212 :   3 - 0x3
      10'hD5: dout  = 8'b00010001; //  213 :  17 - 0x11
      10'hD6: dout  = 8'b00100000; //  214 :  32 - 0x20
      10'hD7: dout  = 8'b00100000; //  215 :  32 - 0x20
      10'hD8: dout  = 8'b00100000; //  216 :  32 - 0x20
      10'hD9: dout  = 8'b00100000; //  217 :  32 - 0x20
      10'hDA: dout  = 8'b00100000; //  218 :  32 - 0x20
      10'hDB: dout  = 8'b00100000; //  219 :  32 - 0x20
      10'hDC: dout  = 8'b00100000; //  220 :  32 - 0x20
      10'hDD: dout  = 8'b00100000; //  221 :  32 - 0x20
      10'hDE: dout  = 8'b00100000; //  222 :  32 - 0x20
      10'hDF: dout  = 8'b00100000; //  223 :  32 - 0x20
      10'hE0: dout  = 8'b00101101; //  224 :  45 - 0x2d -- line 0x7
      10'hE1: dout  = 8'b00010001; //  225 :  17 - 0x11
      10'hE2: dout  = 8'b00000011; //  226 :   3 - 0x3
      10'hE3: dout  = 8'b00000011; //  227 :   3 - 0x3
      10'hE4: dout  = 8'b00000011; //  228 :   3 - 0x3
      10'hE5: dout  = 8'b00000011; //  229 :   3 - 0x3
      10'hE6: dout  = 8'b00000011; //  230 :   3 - 0x3
      10'hE7: dout  = 8'b00000011; //  231 :   3 - 0x3
      10'hE8: dout  = 8'b00000011; //  232 :   3 - 0x3
      10'hE9: dout  = 8'b00000011; //  233 :   3 - 0x3
      10'hEA: dout  = 8'b00000011; //  234 :   3 - 0x3
      10'hEB: dout  = 8'b00000011; //  235 :   3 - 0x3
      10'hEC: dout  = 8'b00000011; //  236 :   3 - 0x3
      10'hED: dout  = 8'b00000011; //  237 :   3 - 0x3
      10'hEE: dout  = 8'b00000011; //  238 :   3 - 0x3
      10'hEF: dout  = 8'b00000011; //  239 :   3 - 0x3
      10'hF0: dout  = 8'b00000011; //  240 :   3 - 0x3
      10'hF1: dout  = 8'b00000011; //  241 :   3 - 0x3
      10'hF2: dout  = 8'b00000011; //  242 :   3 - 0x3
      10'hF3: dout  = 8'b00000011; //  243 :   3 - 0x3
      10'hF4: dout  = 8'b00000011; //  244 :   3 - 0x3
      10'hF5: dout  = 8'b00010001; //  245 :  17 - 0x11
      10'hF6: dout  = 8'b00100000; //  246 :  32 - 0x20
      10'hF7: dout  = 8'b00100000; //  247 :  32 - 0x20
      10'hF8: dout  = 8'b00100000; //  248 :  32 - 0x20
      10'hF9: dout  = 8'b00100000; //  249 :  32 - 0x20
      10'hFA: dout  = 8'b00100000; //  250 :  32 - 0x20
      10'hFB: dout  = 8'b00100000; //  251 :  32 - 0x20
      10'hFC: dout  = 8'b00100000; //  252 :  32 - 0x20
      10'hFD: dout  = 8'b00100000; //  253 :  32 - 0x20
      10'hFE: dout  = 8'b00100000; //  254 :  32 - 0x20
      10'hFF: dout  = 8'b00100000; //  255 :  32 - 0x20
      10'h100: dout  = 8'b00101101; //  256 :  45 - 0x2d -- line 0x8
      10'h101: dout  = 8'b00010001; //  257 :  17 - 0x11
      10'h102: dout  = 8'b00000011; //  258 :   3 - 0x3
      10'h103: dout  = 8'b00011111; //  259 :  31 - 0x1f
      10'h104: dout  = 8'b00010000; //  260 :  16 - 0x10
      10'h105: dout  = 8'b00011101; //  261 :  29 - 0x1d
      10'h106: dout  = 8'b00000011; //  262 :   3 - 0x3
      10'h107: dout  = 8'b00011011; //  263 :  27 - 0x1b
      10'h108: dout  = 8'b00000011; //  264 :   3 - 0x3
      10'h109: dout  = 8'b00011111; //  265 :  31 - 0x1f
      10'h10A: dout  = 8'b00010000; //  266 :  16 - 0x10
      10'h10B: dout  = 8'b00010000; //  267 :  16 - 0x10
      10'h10C: dout  = 8'b00010000; //  268 :  16 - 0x10
      10'h10D: dout  = 8'b00011101; //  269 :  29 - 0x1d
      10'h10E: dout  = 8'b00000011; //  270 :   3 - 0x3
      10'h10F: dout  = 8'b00011011; //  271 :  27 - 0x1b
      10'h110: dout  = 8'b00000011; //  272 :   3 - 0x3
      10'h111: dout  = 8'b00011111; //  273 :  31 - 0x1f
      10'h112: dout  = 8'b00010000; //  274 :  16 - 0x10
      10'h113: dout  = 8'b00011101; //  275 :  29 - 0x1d
      10'h114: dout  = 8'b00000011; //  276 :   3 - 0x3
      10'h115: dout  = 8'b00010001; //  277 :  17 - 0x11
      10'h116: dout  = 8'b00100000; //  278 :  32 - 0x20
      10'h117: dout  = 8'b00100000; //  279 :  32 - 0x20
      10'h118: dout  = 8'b00100000; //  280 :  32 - 0x20
      10'h119: dout  = 8'b00100000; //  281 :  32 - 0x20
      10'h11A: dout  = 8'b00100000; //  282 :  32 - 0x20
      10'h11B: dout  = 8'b00100000; //  283 :  32 - 0x20
      10'h11C: dout  = 8'b00100000; //  284 :  32 - 0x20
      10'h11D: dout  = 8'b00100000; //  285 :  32 - 0x20
      10'h11E: dout  = 8'b00100000; //  286 :  32 - 0x20
      10'h11F: dout  = 8'b00100000; //  287 :  32 - 0x20
      10'h120: dout  = 8'b00101101; //  288 :  45 - 0x2d -- line 0x9
      10'h121: dout  = 8'b00010001; //  289 :  17 - 0x11
      10'h122: dout  = 8'b00000011; //  290 :   3 - 0x3
      10'h123: dout  = 8'b00011110; //  291 :  30 - 0x1e
      10'h124: dout  = 8'b00010000; //  292 :  16 - 0x10
      10'h125: dout  = 8'b00011100; //  293 :  28 - 0x1c
      10'h126: dout  = 8'b00000011; //  294 :   3 - 0x3
      10'h127: dout  = 8'b00010001; //  295 :  17 - 0x11
      10'h128: dout  = 8'b00000011; //  296 :   3 - 0x3
      10'h129: dout  = 8'b00011110; //  297 :  30 - 0x1e
      10'h12A: dout  = 8'b00010000; //  298 :  16 - 0x10
      10'h12B: dout  = 8'b00010011; //  299 :  19 - 0x13
      10'h12C: dout  = 8'b00010000; //  300 :  16 - 0x10
      10'h12D: dout  = 8'b00011100; //  301 :  28 - 0x1c
      10'h12E: dout  = 8'b00000011; //  302 :   3 - 0x3
      10'h12F: dout  = 8'b00010001; //  303 :  17 - 0x11
      10'h130: dout  = 8'b00000011; //  304 :   3 - 0x3
      10'h131: dout  = 8'b00011110; //  305 :  30 - 0x1e
      10'h132: dout  = 8'b00010000; //  306 :  16 - 0x10
      10'h133: dout  = 8'b00011100; //  307 :  28 - 0x1c
      10'h134: dout  = 8'b00000011; //  308 :   3 - 0x3
      10'h135: dout  = 8'b00010001; //  309 :  17 - 0x11
      10'h136: dout  = 8'b00100000; //  310 :  32 - 0x20
      10'h137: dout  = 8'b00100000; //  311 :  32 - 0x20
      10'h138: dout  = 8'b00100000; //  312 :  32 - 0x20
      10'h139: dout  = 8'b00100000; //  313 :  32 - 0x20
      10'h13A: dout  = 8'b00100000; //  314 :  32 - 0x20
      10'h13B: dout  = 8'b00110000; //  315 :  48 - 0x30
      10'h13C: dout  = 8'b00110000; //  316 :  48 - 0x30
      10'h13D: dout  = 8'b00100000; //  317 :  32 - 0x20
      10'h13E: dout  = 8'b00100000; //  318 :  32 - 0x20
      10'h13F: dout  = 8'b00100000; //  319 :  32 - 0x20
      10'h140: dout  = 8'b00101101; //  320 :  45 - 0x2d -- line 0xa
      10'h141: dout  = 8'b00010001; //  321 :  17 - 0x11
      10'h142: dout  = 8'b00000011; //  322 :   3 - 0x3
      10'h143: dout  = 8'b00000011; //  323 :   3 - 0x3
      10'h144: dout  = 8'b00000011; //  324 :   3 - 0x3
      10'h145: dout  = 8'b00000011; //  325 :   3 - 0x3
      10'h146: dout  = 8'b00000011; //  326 :   3 - 0x3
      10'h147: dout  = 8'b00010001; //  327 :  17 - 0x11
      10'h148: dout  = 8'b00000011; //  328 :   3 - 0x3
      10'h149: dout  = 8'b00000011; //  329 :   3 - 0x3
      10'h14A: dout  = 8'b00000011; //  330 :   3 - 0x3
      10'h14B: dout  = 8'b00010001; //  331 :  17 - 0x11
      10'h14C: dout  = 8'b00000011; //  332 :   3 - 0x3
      10'h14D: dout  = 8'b00000011; //  333 :   3 - 0x3
      10'h14E: dout  = 8'b00000011; //  334 :   3 - 0x3
      10'h14F: dout  = 8'b00010001; //  335 :  17 - 0x11
      10'h150: dout  = 8'b00000011; //  336 :   3 - 0x3
      10'h151: dout  = 8'b00000011; //  337 :   3 - 0x3
      10'h152: dout  = 8'b00000011; //  338 :   3 - 0x3
      10'h153: dout  = 8'b00000011; //  339 :   3 - 0x3
      10'h154: dout  = 8'b00000011; //  340 :   3 - 0x3
      10'h155: dout  = 8'b00010001; //  341 :  17 - 0x11
      10'h156: dout  = 8'b00100000; //  342 :  32 - 0x20
      10'h157: dout  = 8'b00100000; //  343 :  32 - 0x20
      10'h158: dout  = 8'b00100000; //  344 :  32 - 0x20
      10'h159: dout  = 8'b00100000; //  345 :  32 - 0x20
      10'h15A: dout  = 8'b00100000; //  346 :  32 - 0x20
      10'h15B: dout  = 8'b00100000; //  347 :  32 - 0x20
      10'h15C: dout  = 8'b00100000; //  348 :  32 - 0x20
      10'h15D: dout  = 8'b00100000; //  349 :  32 - 0x20
      10'h15E: dout  = 8'b00100000; //  350 :  32 - 0x20
      10'h15F: dout  = 8'b00100000; //  351 :  32 - 0x20
      10'h160: dout  = 8'b00101101; //  352 :  45 - 0x2d -- line 0xb
      10'h161: dout  = 8'b00011110; //  353 :  30 - 0x1e
      10'h162: dout  = 8'b00010000; //  354 :  16 - 0x10
      10'h163: dout  = 8'b00010000; //  355 :  16 - 0x10
      10'h164: dout  = 8'b00010000; //  356 :  16 - 0x10
      10'h165: dout  = 8'b00011101; //  357 :  29 - 0x1d
      10'h166: dout  = 8'b00000011; //  358 :   3 - 0x3
      10'h167: dout  = 8'b00010101; //  359 :  21 - 0x15
      10'h168: dout  = 8'b00010000; //  360 :  16 - 0x10
      10'h169: dout  = 8'b00011000; //  361 :  24 - 0x18
      10'h16A: dout  = 8'b00001000; //  362 :   8 - 0x8
      10'h16B: dout  = 8'b00011010; //  363 :  26 - 0x1a
      10'h16C: dout  = 8'b00001000; //  364 :   8 - 0x8
      10'h16D: dout  = 8'b00011001; //  365 :  25 - 0x19
      10'h16E: dout  = 8'b00010000; //  366 :  16 - 0x10
      10'h16F: dout  = 8'b00010100; //  367 :  20 - 0x14
      10'h170: dout  = 8'b00000011; //  368 :   3 - 0x3
      10'h171: dout  = 8'b00011111; //  369 :  31 - 0x1f
      10'h172: dout  = 8'b00010000; //  370 :  16 - 0x10
      10'h173: dout  = 8'b00010000; //  371 :  16 - 0x10
      10'h174: dout  = 8'b00010000; //  372 :  16 - 0x10
      10'h175: dout  = 8'b00011100; //  373 :  28 - 0x1c
      10'h176: dout  = 8'b00100000; //  374 :  32 - 0x20
      10'h177: dout  = 8'b00100000; //  375 :  32 - 0x20
      10'h178: dout  = 8'b00100000; //  376 :  32 - 0x20
      10'h179: dout  = 8'b00100000; //  377 :  32 - 0x20
      10'h17A: dout  = 8'b00100000; //  378 :  32 - 0x20
      10'h17B: dout  = 8'b00100000; //  379 :  32 - 0x20
      10'h17C: dout  = 8'b00100000; //  380 :  32 - 0x20
      10'h17D: dout  = 8'b00100000; //  381 :  32 - 0x20
      10'h17E: dout  = 8'b00100000; //  382 :  32 - 0x20
      10'h17F: dout  = 8'b00100000; //  383 :  32 - 0x20
      10'h180: dout  = 8'b00101101; //  384 :  45 - 0x2d -- line 0xc
      10'h181: dout  = 8'b00100000; //  385 :  32 - 0x20
      10'h182: dout  = 8'b00100000; //  386 :  32 - 0x20
      10'h183: dout  = 8'b00100000; //  387 :  32 - 0x20
      10'h184: dout  = 8'b00100000; //  388 :  32 - 0x20
      10'h185: dout  = 8'b00010001; //  389 :  17 - 0x11
      10'h186: dout  = 8'b00000011; //  390 :   3 - 0x3
      10'h187: dout  = 8'b00010001; //  391 :  17 - 0x11
      10'h188: dout  = 8'b00000000; //  392 :   0 - 0x0
      10'h189: dout  = 8'b00000000; //  393 :   0 - 0x0
      10'h18A: dout  = 8'b00000000; //  394 :   0 - 0x0
      10'h18B: dout  = 8'b00000000; //  395 :   0 - 0x0
      10'h18C: dout  = 8'b00000000; //  396 :   0 - 0x0
      10'h18D: dout  = 8'b00000000; //  397 :   0 - 0x0
      10'h18E: dout  = 8'b00000000; //  398 :   0 - 0x0
      10'h18F: dout  = 8'b00010001; //  399 :  17 - 0x11
      10'h190: dout  = 8'b00000011; //  400 :   3 - 0x3
      10'h191: dout  = 8'b00010001; //  401 :  17 - 0x11
      10'h192: dout  = 8'b00100000; //  402 :  32 - 0x20
      10'h193: dout  = 8'b00100000; //  403 :  32 - 0x20
      10'h194: dout  = 8'b00100000; //  404 :  32 - 0x20
      10'h195: dout  = 8'b00100000; //  405 :  32 - 0x20
      10'h196: dout  = 8'b00100000; //  406 :  32 - 0x20
      10'h197: dout  = 8'b00100000; //  407 :  32 - 0x20
      10'h198: dout  = 8'b00100000; //  408 :  32 - 0x20
      10'h199: dout  = 8'b00100000; //  409 :  32 - 0x20
      10'h19A: dout  = 8'b00100000; //  410 :  32 - 0x20
      10'h19B: dout  = 8'b00100000; //  411 :  32 - 0x20
      10'h19C: dout  = 8'b00100000; //  412 :  32 - 0x20
      10'h19D: dout  = 8'b00100000; //  413 :  32 - 0x20
      10'h19E: dout  = 8'b00100000; //  414 :  32 - 0x20
      10'h19F: dout  = 8'b00100000; //  415 :  32 - 0x20
      10'h1A0: dout  = 8'b00101101; //  416 :  45 - 0x2d -- line 0xd
      10'h1A1: dout  = 8'b00100000; //  417 :  32 - 0x20
      10'h1A2: dout  = 8'b00100000; //  418 :  32 - 0x20
      10'h1A3: dout  = 8'b00100000; //  419 :  32 - 0x20
      10'h1A4: dout  = 8'b00100000; //  420 :  32 - 0x20
      10'h1A5: dout  = 8'b00010001; //  421 :  17 - 0x11
      10'h1A6: dout  = 8'b00000011; //  422 :   3 - 0x3
      10'h1A7: dout  = 8'b00010001; //  423 :  17 - 0x11
      10'h1A8: dout  = 8'b00000000; //  424 :   0 - 0x0
      10'h1A9: dout  = 8'b00011111; //  425 :  31 - 0x1f
      10'h1AA: dout  = 8'b00010111; //  426 :  23 - 0x17
      10'h1AB: dout  = 8'b00101100; //  427 :  44 - 0x2c
      10'h1AC: dout  = 8'b00010110; //  428 :  22 - 0x16
      10'h1AD: dout  = 8'b00011101; //  429 :  29 - 0x1d
      10'h1AE: dout  = 8'b00000000; //  430 :   0 - 0x0
      10'h1AF: dout  = 8'b00010001; //  431 :  17 - 0x11
      10'h1B0: dout  = 8'b00000011; //  432 :   3 - 0x3
      10'h1B1: dout  = 8'b00010001; //  433 :  17 - 0x11
      10'h1B2: dout  = 8'b00100000; //  434 :  32 - 0x20
      10'h1B3: dout  = 8'b00100000; //  435 :  32 - 0x20
      10'h1B4: dout  = 8'b00100000; //  436 :  32 - 0x20
      10'h1B5: dout  = 8'b00100000; //  437 :  32 - 0x20
      10'h1B6: dout  = 8'b00100000; //  438 :  32 - 0x20
      10'h1B7: dout  = 8'b00100000; //  439 :  32 - 0x20
      10'h1B8: dout  = 8'b00100000; //  440 :  32 - 0x20
      10'h1B9: dout  = 8'b00100000; //  441 :  32 - 0x20
      10'h1BA: dout  = 8'b00100000; //  442 :  32 - 0x20
      10'h1BB: dout  = 8'b00100000; //  443 :  32 - 0x20
      10'h1BC: dout  = 8'b00100000; //  444 :  32 - 0x20
      10'h1BD: dout  = 8'b00100000; //  445 :  32 - 0x20
      10'h1BE: dout  = 8'b00100000; //  446 :  32 - 0x20
      10'h1BF: dout  = 8'b00100000; //  447 :  32 - 0x20
      10'h1C0: dout  = 8'b00101101; //  448 :  45 - 0x2d -- line 0xe
      10'h1C1: dout  = 8'b00100010; //  449 :  34 - 0x22
      10'h1C2: dout  = 8'b00010000; //  450 :  16 - 0x10
      10'h1C3: dout  = 8'b00010000; //  451 :  16 - 0x10
      10'h1C4: dout  = 8'b00010000; //  452 :  16 - 0x10
      10'h1C5: dout  = 8'b00011100; //  453 :  28 - 0x1c
      10'h1C6: dout  = 8'b00000011; //  454 :   3 - 0x3
      10'h1C7: dout  = 8'b00011010; //  455 :  26 - 0x1a
      10'h1C8: dout  = 8'b00000000; //  456 :   0 - 0x0
      10'h1C9: dout  = 8'b00010001; //  457 :  17 - 0x11
      10'h1CA: dout  = 8'b00000000; //  458 :   0 - 0x0
      10'h1CB: dout  = 8'b00000000; //  459 :   0 - 0x0
      10'h1CC: dout  = 8'b00000000; //  460 :   0 - 0x0
      10'h1CD: dout  = 8'b00010001; //  461 :  17 - 0x11
      10'h1CE: dout  = 8'b00000000; //  462 :   0 - 0x0
      10'h1CF: dout  = 8'b00011010; //  463 :  26 - 0x1a
      10'h1D0: dout  = 8'b00000011; //  464 :   3 - 0x3
      10'h1D1: dout  = 8'b00011110; //  465 :  30 - 0x1e
      10'h1D2: dout  = 8'b00010000; //  466 :  16 - 0x10
      10'h1D3: dout  = 8'b00010000; //  467 :  16 - 0x10
      10'h1D4: dout  = 8'b00010000; //  468 :  16 - 0x10
      10'h1D5: dout  = 8'b00100001; //  469 :  33 - 0x21
      10'h1D6: dout  = 8'b00101101; //  470 :  45 - 0x2d
      10'h1D7: dout  = 8'b00101101; //  471 :  45 - 0x2d
      10'h1D8: dout  = 8'b00101101; //  472 :  45 - 0x2d
      10'h1D9: dout  = 8'b00101101; //  473 :  45 - 0x2d
      10'h1DA: dout  = 8'b00101101; //  474 :  45 - 0x2d
      10'h1DB: dout  = 8'b00101101; //  475 :  45 - 0x2d
      10'h1DC: dout  = 8'b00101101; //  476 :  45 - 0x2d
      10'h1DD: dout  = 8'b00101101; //  477 :  45 - 0x2d
      10'h1DE: dout  = 8'b00100000; //  478 :  32 - 0x20
      10'h1DF: dout  = 8'b00100000; //  479 :  32 - 0x20
      10'h1E0: dout  = 8'b00000100; //  480 :   4 - 0x4 -- line 0xf
      10'h1E1: dout  = 8'b00000110; //  481 :   6 - 0x6
      10'h1E2: dout  = 8'b00000000; //  482 :   0 - 0x0
      10'h1E3: dout  = 8'b00000000; //  483 :   0 - 0x0
      10'h1E4: dout  = 8'b00000000; //  484 :   0 - 0x0
      10'h1E5: dout  = 8'b00000000; //  485 :   0 - 0x0
      10'h1E6: dout  = 8'b00000011; //  486 :   3 - 0x3
      10'h1E7: dout  = 8'b00000000; //  487 :   0 - 0x0
      10'h1E8: dout  = 8'b00000000; //  488 :   0 - 0x0
      10'h1E9: dout  = 8'b00010001; //  489 :  17 - 0x11
      10'h1EA: dout  = 8'b00000000; //  490 :   0 - 0x0
      10'h1EB: dout  = 8'b00000000; //  491 :   0 - 0x0
      10'h1EC: dout  = 8'b00000000; //  492 :   0 - 0x0
      10'h1ED: dout  = 8'b00010001; //  493 :  17 - 0x11
      10'h1EE: dout  = 8'b00000000; //  494 :   0 - 0x0
      10'h1EF: dout  = 8'b00000000; //  495 :   0 - 0x0
      10'h1F0: dout  = 8'b00000011; //  496 :   3 - 0x3
      10'h1F1: dout  = 8'b00000000; //  497 :   0 - 0x0
      10'h1F2: dout  = 8'b00000000; //  498 :   0 - 0x0
      10'h1F3: dout  = 8'b00000000; //  499 :   0 - 0x0
      10'h1F4: dout  = 8'b00000000; //  500 :   0 - 0x0
      10'h1F5: dout  = 8'b00000101; //  501 :   5 - 0x5
      10'h1F6: dout  = 8'b00000100; //  502 :   4 - 0x4
      10'h1F7: dout  = 8'b00000100; //  503 :   4 - 0x4
      10'h1F8: dout  = 8'b00000100; //  504 :   4 - 0x4
      10'h1F9: dout  = 8'b00000100; //  505 :   4 - 0x4
      10'h1FA: dout  = 8'b00000100; //  506 :   4 - 0x4
      10'h1FB: dout  = 8'b00000100; //  507 :   4 - 0x4
      10'h1FC: dout  = 8'b00000100; //  508 :   4 - 0x4
      10'h1FD: dout  = 8'b00000100; //  509 :   4 - 0x4
      10'h1FE: dout  = 8'b00100000; //  510 :  32 - 0x20
      10'h1FF: dout  = 8'b00100000; //  511 :  32 - 0x20
      10'h200: dout  = 8'b00101101; //  512 :  45 - 0x2d -- line 0x10
      10'h201: dout  = 8'b00100010; //  513 :  34 - 0x22
      10'h202: dout  = 8'b00010000; //  514 :  16 - 0x10
      10'h203: dout  = 8'b00010000; //  515 :  16 - 0x10
      10'h204: dout  = 8'b00010000; //  516 :  16 - 0x10
      10'h205: dout  = 8'b00011101; //  517 :  29 - 0x1d
      10'h206: dout  = 8'b00000011; //  518 :   3 - 0x3
      10'h207: dout  = 8'b00011011; //  519 :  27 - 0x1b
      10'h208: dout  = 8'b00000000; //  520 :   0 - 0x0
      10'h209: dout  = 8'b00011110; //  521 :  30 - 0x1e
      10'h20A: dout  = 8'b00010000; //  522 :  16 - 0x10
      10'h20B: dout  = 8'b00010000; //  523 :  16 - 0x10
      10'h20C: dout  = 8'b00010000; //  524 :  16 - 0x10
      10'h20D: dout  = 8'b00011100; //  525 :  28 - 0x1c
      10'h20E: dout  = 8'b00000000; //  526 :   0 - 0x0
      10'h20F: dout  = 8'b00011011; //  527 :  27 - 0x1b
      10'h210: dout  = 8'b00000011; //  528 :   3 - 0x3
      10'h211: dout  = 8'b00011111; //  529 :  31 - 0x1f
      10'h212: dout  = 8'b00010000; //  530 :  16 - 0x10
      10'h213: dout  = 8'b00010000; //  531 :  16 - 0x10
      10'h214: dout  = 8'b00010000; //  532 :  16 - 0x10
      10'h215: dout  = 8'b00100001; //  533 :  33 - 0x21
      10'h216: dout  = 8'b00101101; //  534 :  45 - 0x2d
      10'h217: dout  = 8'b00101101; //  535 :  45 - 0x2d
      10'h218: dout  = 8'b00101101; //  536 :  45 - 0x2d
      10'h219: dout  = 8'b00101101; //  537 :  45 - 0x2d
      10'h21A: dout  = 8'b00101101; //  538 :  45 - 0x2d
      10'h21B: dout  = 8'b00101101; //  539 :  45 - 0x2d
      10'h21C: dout  = 8'b00101101; //  540 :  45 - 0x2d
      10'h21D: dout  = 8'b00101101; //  541 :  45 - 0x2d
      10'h21E: dout  = 8'b00100000; //  542 :  32 - 0x20
      10'h21F: dout  = 8'b00100000; //  543 :  32 - 0x20
      10'h220: dout  = 8'b00101101; //  544 :  45 - 0x2d -- line 0x11
      10'h221: dout  = 8'b00100000; //  545 :  32 - 0x20
      10'h222: dout  = 8'b00100000; //  546 :  32 - 0x20
      10'h223: dout  = 8'b00100000; //  547 :  32 - 0x20
      10'h224: dout  = 8'b00100000; //  548 :  32 - 0x20
      10'h225: dout  = 8'b00010001; //  549 :  17 - 0x11
      10'h226: dout  = 8'b00000011; //  550 :   3 - 0x3
      10'h227: dout  = 8'b00010001; //  551 :  17 - 0x11
      10'h228: dout  = 8'b00000000; //  552 :   0 - 0x0
      10'h229: dout  = 8'b00000000; //  553 :   0 - 0x0
      10'h22A: dout  = 8'b00000000; //  554 :   0 - 0x0
      10'h22B: dout  = 8'b00000000; //  555 :   0 - 0x0
      10'h22C: dout  = 8'b00000000; //  556 :   0 - 0x0
      10'h22D: dout  = 8'b00000000; //  557 :   0 - 0x0
      10'h22E: dout  = 8'b00000000; //  558 :   0 - 0x0
      10'h22F: dout  = 8'b00010001; //  559 :  17 - 0x11
      10'h230: dout  = 8'b00000011; //  560 :   3 - 0x3
      10'h231: dout  = 8'b00010001; //  561 :  17 - 0x11
      10'h232: dout  = 8'b00100000; //  562 :  32 - 0x20
      10'h233: dout  = 8'b00100000; //  563 :  32 - 0x20
      10'h234: dout  = 8'b00100000; //  564 :  32 - 0x20
      10'h235: dout  = 8'b00100000; //  565 :  32 - 0x20
      10'h236: dout  = 8'b00100000; //  566 :  32 - 0x20
      10'h237: dout  = 8'b00100000; //  567 :  32 - 0x20
      10'h238: dout  = 8'b00100000; //  568 :  32 - 0x20
      10'h239: dout  = 8'b00100000; //  569 :  32 - 0x20
      10'h23A: dout  = 8'b00100000; //  570 :  32 - 0x20
      10'h23B: dout  = 8'b00100000; //  571 :  32 - 0x20
      10'h23C: dout  = 8'b00100000; //  572 :  32 - 0x20
      10'h23D: dout  = 8'b00100000; //  573 :  32 - 0x20
      10'h23E: dout  = 8'b00100000; //  574 :  32 - 0x20
      10'h23F: dout  = 8'b00100000; //  575 :  32 - 0x20
      10'h240: dout  = 8'b00101101; //  576 :  45 - 0x2d -- line 0x12
      10'h241: dout  = 8'b00100000; //  577 :  32 - 0x20
      10'h242: dout  = 8'b00100000; //  578 :  32 - 0x20
      10'h243: dout  = 8'b00100000; //  579 :  32 - 0x20
      10'h244: dout  = 8'b00100000; //  580 :  32 - 0x20
      10'h245: dout  = 8'b00010001; //  581 :  17 - 0x11
      10'h246: dout  = 8'b00000011; //  582 :   3 - 0x3
      10'h247: dout  = 8'b00010001; //  583 :  17 - 0x11
      10'h248: dout  = 8'b00000000; //  584 :   0 - 0x0
      10'h249: dout  = 8'b00011111; //  585 :  31 - 0x1f
      10'h24A: dout  = 8'b00010000; //  586 :  16 - 0x10
      10'h24B: dout  = 8'b00010000; //  587 :  16 - 0x10
      10'h24C: dout  = 8'b00010000; //  588 :  16 - 0x10
      10'h24D: dout  = 8'b00011101; //  589 :  29 - 0x1d
      10'h24E: dout  = 8'b00000000; //  590 :   0 - 0x0
      10'h24F: dout  = 8'b00010001; //  591 :  17 - 0x11
      10'h250: dout  = 8'b00000011; //  592 :   3 - 0x3
      10'h251: dout  = 8'b00010001; //  593 :  17 - 0x11
      10'h252: dout  = 8'b00100000; //  594 :  32 - 0x20
      10'h253: dout  = 8'b00100000; //  595 :  32 - 0x20
      10'h254: dout  = 8'b00100000; //  596 :  32 - 0x20
      10'h255: dout  = 8'b00100000; //  597 :  32 - 0x20
      10'h256: dout  = 8'b01100000; //  598 :  96 - 0x60
      10'h257: dout  = 8'b01100001; //  599 :  97 - 0x61
      10'h258: dout  = 8'b00100000; //  600 :  32 - 0x20
      10'h259: dout  = 8'b00100000; //  601 :  32 - 0x20
      10'h25A: dout  = 8'b00100000; //  602 :  32 - 0x20
      10'h25B: dout  = 8'b00100000; //  603 :  32 - 0x20
      10'h25C: dout  = 8'b00101101; //  604 :  45 - 0x2d
      10'h25D: dout  = 8'b00101101; //  605 :  45 - 0x2d
      10'h25E: dout  = 8'b00100000; //  606 :  32 - 0x20
      10'h25F: dout  = 8'b00100000; //  607 :  32 - 0x20
      10'h260: dout  = 8'b00101101; //  608 :  45 - 0x2d -- line 0x13
      10'h261: dout  = 8'b00011111; //  609 :  31 - 0x1f
      10'h262: dout  = 8'b00010000; //  610 :  16 - 0x10
      10'h263: dout  = 8'b00010000; //  611 :  16 - 0x10
      10'h264: dout  = 8'b00010000; //  612 :  16 - 0x10
      10'h265: dout  = 8'b00011100; //  613 :  28 - 0x1c
      10'h266: dout  = 8'b00000011; //  614 :   3 - 0x3
      10'h267: dout  = 8'b00011010; //  615 :  26 - 0x1a
      10'h268: dout  = 8'b00000000; //  616 :   0 - 0x0
      10'h269: dout  = 8'b00011110; //  617 :  30 - 0x1e
      10'h26A: dout  = 8'b00010000; //  618 :  16 - 0x10
      10'h26B: dout  = 8'b00010011; //  619 :  19 - 0x13
      10'h26C: dout  = 8'b00010000; //  620 :  16 - 0x10
      10'h26D: dout  = 8'b00011100; //  621 :  28 - 0x1c
      10'h26E: dout  = 8'b00000000; //  622 :   0 - 0x0
      10'h26F: dout  = 8'b00011010; //  623 :  26 - 0x1a
      10'h270: dout  = 8'b00000011; //  624 :   3 - 0x3
      10'h271: dout  = 8'b00011110; //  625 :  30 - 0x1e
      10'h272: dout  = 8'b00010000; //  626 :  16 - 0x10
      10'h273: dout  = 8'b00010000; //  627 :  16 - 0x10
      10'h274: dout  = 8'b00010000; //  628 :  16 - 0x10
      10'h275: dout  = 8'b00011101; //  629 :  29 - 0x1d
      10'h276: dout  = 8'b01100010; //  630 :  98 - 0x62
      10'h277: dout  = 8'b01100011; //  631 :  99 - 0x63
      10'h278: dout  = 8'b00100000; //  632 :  32 - 0x20
      10'h279: dout  = 8'b00100000; //  633 :  32 - 0x20
      10'h27A: dout  = 8'b00100000; //  634 :  32 - 0x20
      10'h27B: dout  = 8'b00100000; //  635 :  32 - 0x20
      10'h27C: dout  = 8'b00101101; //  636 :  45 - 0x2d
      10'h27D: dout  = 8'b00101101; //  637 :  45 - 0x2d
      10'h27E: dout  = 8'b00100000; //  638 :  32 - 0x20
      10'h27F: dout  = 8'b00100000; //  639 :  32 - 0x20
      10'h280: dout  = 8'b00101101; //  640 :  45 - 0x2d -- line 0x14
      10'h281: dout  = 8'b00010001; //  641 :  17 - 0x11
      10'h282: dout  = 8'b00000011; //  642 :   3 - 0x3
      10'h283: dout  = 8'b00000011; //  643 :   3 - 0x3
      10'h284: dout  = 8'b00000011; //  644 :   3 - 0x3
      10'h285: dout  = 8'b00000011; //  645 :   3 - 0x3
      10'h286: dout  = 8'b00000011; //  646 :   3 - 0x3
      10'h287: dout  = 8'b00000011; //  647 :   3 - 0x3
      10'h288: dout  = 8'b00000011; //  648 :   3 - 0x3
      10'h289: dout  = 8'b00000011; //  649 :   3 - 0x3
      10'h28A: dout  = 8'b00000011; //  650 :   3 - 0x3
      10'h28B: dout  = 8'b00010001; //  651 :  17 - 0x11
      10'h28C: dout  = 8'b00000011; //  652 :   3 - 0x3
      10'h28D: dout  = 8'b00000011; //  653 :   3 - 0x3
      10'h28E: dout  = 8'b00000011; //  654 :   3 - 0x3
      10'h28F: dout  = 8'b00000011; //  655 :   3 - 0x3
      10'h290: dout  = 8'b00000011; //  656 :   3 - 0x3
      10'h291: dout  = 8'b00000011; //  657 :   3 - 0x3
      10'h292: dout  = 8'b00000011; //  658 :   3 - 0x3
      10'h293: dout  = 8'b00000011; //  659 :   3 - 0x3
      10'h294: dout  = 8'b00000011; //  660 :   3 - 0x3
      10'h295: dout  = 8'b00010001; //  661 :  17 - 0x11
      10'h296: dout  = 8'b00100000; //  662 :  32 - 0x20
      10'h297: dout  = 8'b00100000; //  663 :  32 - 0x20
      10'h298: dout  = 8'b00100000; //  664 :  32 - 0x20
      10'h299: dout  = 8'b00100000; //  665 :  32 - 0x20
      10'h29A: dout  = 8'b00100000; //  666 :  32 - 0x20
      10'h29B: dout  = 8'b00100000; //  667 :  32 - 0x20
      10'h29C: dout  = 8'b00101101; //  668 :  45 - 0x2d
      10'h29D: dout  = 8'b00101101; //  669 :  45 - 0x2d
      10'h29E: dout  = 8'b00100000; //  670 :  32 - 0x20
      10'h29F: dout  = 8'b00100000; //  671 :  32 - 0x20
      10'h2A0: dout  = 8'b00101101; //  672 :  45 - 0x2d -- line 0x15
      10'h2A1: dout  = 8'b00010001; //  673 :  17 - 0x11
      10'h2A2: dout  = 8'b00000011; //  674 :   3 - 0x3
      10'h2A3: dout  = 8'b00011001; //  675 :  25 - 0x19
      10'h2A4: dout  = 8'b00010000; //  676 :  16 - 0x10
      10'h2A5: dout  = 8'b00011101; //  677 :  29 - 0x1d
      10'h2A6: dout  = 8'b00000011; //  678 :   3 - 0x3
      10'h2A7: dout  = 8'b00011001; //  679 :  25 - 0x19
      10'h2A8: dout  = 8'b00010000; //  680 :  16 - 0x10
      10'h2A9: dout  = 8'b00011000; //  681 :  24 - 0x18
      10'h2AA: dout  = 8'b00001001; //  682 :   9 - 0x9
      10'h2AB: dout  = 8'b00011010; //  683 :  26 - 0x1a
      10'h2AC: dout  = 8'b00001001; //  684 :   9 - 0x9
      10'h2AD: dout  = 8'b00011001; //  685 :  25 - 0x19
      10'h2AE: dout  = 8'b00010000; //  686 :  16 - 0x10
      10'h2AF: dout  = 8'b00011000; //  687 :  24 - 0x18
      10'h2B0: dout  = 8'b00000011; //  688 :   3 - 0x3
      10'h2B1: dout  = 8'b00011111; //  689 :  31 - 0x1f
      10'h2B2: dout  = 8'b00010000; //  690 :  16 - 0x10
      10'h2B3: dout  = 8'b00011000; //  691 :  24 - 0x18
      10'h2B4: dout  = 8'b00000011; //  692 :   3 - 0x3
      10'h2B5: dout  = 8'b00010001; //  693 :  17 - 0x11
      10'h2B6: dout  = 8'b00100000; //  694 :  32 - 0x20
      10'h2B7: dout  = 8'b00100000; //  695 :  32 - 0x20
      10'h2B8: dout  = 8'b00100000; //  696 :  32 - 0x20
      10'h2B9: dout  = 8'b00100000; //  697 :  32 - 0x20
      10'h2BA: dout  = 8'b00100000; //  698 :  32 - 0x20
      10'h2BB: dout  = 8'b00100000; //  699 :  32 - 0x20
      10'h2BC: dout  = 8'b00101101; //  700 :  45 - 0x2d
      10'h2BD: dout  = 8'b00101101; //  701 :  45 - 0x2d
      10'h2BE: dout  = 8'b00100000; //  702 :  32 - 0x20
      10'h2BF: dout  = 8'b00100000; //  703 :  32 - 0x20
      10'h2C0: dout  = 8'b00101101; //  704 :  45 - 0x2d -- line 0x16
      10'h2C1: dout  = 8'b00010001; //  705 :  17 - 0x11
      10'h2C2: dout  = 8'b00000001; //  706 :   1 - 0x1
      10'h2C3: dout  = 8'b00000011; //  707 :   3 - 0x3
      10'h2C4: dout  = 8'b00000011; //  708 :   3 - 0x3
      10'h2C5: dout  = 8'b00010001; //  709 :  17 - 0x11
      10'h2C6: dout  = 8'b00000011; //  710 :   3 - 0x3
      10'h2C7: dout  = 8'b00000011; //  711 :   3 - 0x3
      10'h2C8: dout  = 8'b00000011; //  712 :   3 - 0x3
      10'h2C9: dout  = 8'b00000011; //  713 :   3 - 0x3
      10'h2CA: dout  = 8'b00000011; //  714 :   3 - 0x3
      10'h2CB: dout  = 8'b00000000; //  715 :   0 - 0x0
      10'h2CC: dout  = 8'b00000011; //  716 :   3 - 0x3
      10'h2CD: dout  = 8'b00000011; //  717 :   3 - 0x3
      10'h2CE: dout  = 8'b00000011; //  718 :   3 - 0x3
      10'h2CF: dout  = 8'b00000011; //  719 :   3 - 0x3
      10'h2D0: dout  = 8'b00000011; //  720 :   3 - 0x3
      10'h2D1: dout  = 8'b00010001; //  721 :  17 - 0x11
      10'h2D2: dout  = 8'b00000011; //  722 :   3 - 0x3
      10'h2D3: dout  = 8'b00000011; //  723 :   3 - 0x3
      10'h2D4: dout  = 8'b00000001; //  724 :   1 - 0x1
      10'h2D5: dout  = 8'b00010001; //  725 :  17 - 0x11
      10'h2D6: dout  = 8'b00100000; //  726 :  32 - 0x20
      10'h2D7: dout  = 8'b00100000; //  727 :  32 - 0x20
      10'h2D8: dout  = 8'b00100000; //  728 :  32 - 0x20
      10'h2D9: dout  = 8'b00100000; //  729 :  32 - 0x20
      10'h2DA: dout  = 8'b00100000; //  730 :  32 - 0x20
      10'h2DB: dout  = 8'b00100000; //  731 :  32 - 0x20
      10'h2DC: dout  = 8'b00101101; //  732 :  45 - 0x2d
      10'h2DD: dout  = 8'b00101101; //  733 :  45 - 0x2d
      10'h2DE: dout  = 8'b00100000; //  734 :  32 - 0x20
      10'h2DF: dout  = 8'b00100000; //  735 :  32 - 0x20
      10'h2E0: dout  = 8'b00101101; //  736 :  45 - 0x2d -- line 0x17
      10'h2E1: dout  = 8'b00010101; //  737 :  21 - 0x15
      10'h2E2: dout  = 8'b00010000; //  738 :  16 - 0x10
      10'h2E3: dout  = 8'b00011101; //  739 :  29 - 0x1d
      10'h2E4: dout  = 8'b00000011; //  740 :   3 - 0x3
      10'h2E5: dout  = 8'b00010001; //  741 :  17 - 0x11
      10'h2E6: dout  = 8'b00000011; //  742 :   3 - 0x3
      10'h2E7: dout  = 8'b00011011; //  743 :  27 - 0x1b
      10'h2E8: dout  = 8'b00000011; //  744 :   3 - 0x3
      10'h2E9: dout  = 8'b00011111; //  745 :  31 - 0x1f
      10'h2EA: dout  = 8'b00010000; //  746 :  16 - 0x10
      10'h2EB: dout  = 8'b00010000; //  747 :  16 - 0x10
      10'h2EC: dout  = 8'b00010000; //  748 :  16 - 0x10
      10'h2ED: dout  = 8'b00011101; //  749 :  29 - 0x1d
      10'h2EE: dout  = 8'b00000011; //  750 :   3 - 0x3
      10'h2EF: dout  = 8'b00011011; //  751 :  27 - 0x1b
      10'h2F0: dout  = 8'b00000011; //  752 :   3 - 0x3
      10'h2F1: dout  = 8'b00010001; //  753 :  17 - 0x11
      10'h2F2: dout  = 8'b00000011; //  754 :   3 - 0x3
      10'h2F3: dout  = 8'b00011111; //  755 :  31 - 0x1f
      10'h2F4: dout  = 8'b00010000; //  756 :  16 - 0x10
      10'h2F5: dout  = 8'b00010100; //  757 :  20 - 0x14
      10'h2F6: dout  = 8'b00100000; //  758 :  32 - 0x20
      10'h2F7: dout  = 8'b00100000; //  759 :  32 - 0x20
      10'h2F8: dout  = 8'b00100000; //  760 :  32 - 0x20
      10'h2F9: dout  = 8'b00100000; //  761 :  32 - 0x20
      10'h2FA: dout  = 8'b00100000; //  762 :  32 - 0x20
      10'h2FB: dout  = 8'b00100000; //  763 :  32 - 0x20
      10'h2FC: dout  = 8'b00101101; //  764 :  45 - 0x2d
      10'h2FD: dout  = 8'b00101101; //  765 :  45 - 0x2d
      10'h2FE: dout  = 8'b00100000; //  766 :  32 - 0x20
      10'h2FF: dout  = 8'b00100000; //  767 :  32 - 0x20
      10'h300: dout  = 8'b00101101; //  768 :  45 - 0x2d -- line 0x18
      10'h301: dout  = 8'b00010101; //  769 :  21 - 0x15
      10'h302: dout  = 8'b00010000; //  770 :  16 - 0x10
      10'h303: dout  = 8'b00011100; //  771 :  28 - 0x1c
      10'h304: dout  = 8'b00000011; //  772 :   3 - 0x3
      10'h305: dout  = 8'b00011010; //  773 :  26 - 0x1a
      10'h306: dout  = 8'b00000011; //  774 :   3 - 0x3
      10'h307: dout  = 8'b00010001; //  775 :  17 - 0x11
      10'h308: dout  = 8'b00000011; //  776 :   3 - 0x3
      10'h309: dout  = 8'b00011110; //  777 :  30 - 0x1e
      10'h30A: dout  = 8'b00010000; //  778 :  16 - 0x10
      10'h30B: dout  = 8'b00010011; //  779 :  19 - 0x13
      10'h30C: dout  = 8'b00010000; //  780 :  16 - 0x10
      10'h30D: dout  = 8'b00011100; //  781 :  28 - 0x1c
      10'h30E: dout  = 8'b00000011; //  782 :   3 - 0x3
      10'h30F: dout  = 8'b00010001; //  783 :  17 - 0x11
      10'h310: dout  = 8'b00000011; //  784 :   3 - 0x3
      10'h311: dout  = 8'b00011010; //  785 :  26 - 0x1a
      10'h312: dout  = 8'b00000011; //  786 :   3 - 0x3
      10'h313: dout  = 8'b00011110; //  787 :  30 - 0x1e
      10'h314: dout  = 8'b00010000; //  788 :  16 - 0x10
      10'h315: dout  = 8'b00010100; //  789 :  20 - 0x14
      10'h316: dout  = 8'b00100000; //  790 :  32 - 0x20
      10'h317: dout  = 8'b00111100; //  791 :  60 - 0x3c
      10'h318: dout  = 8'b00111101; //  792 :  61 - 0x3d
      10'h319: dout  = 8'b00111100; //  793 :  60 - 0x3c
      10'h31A: dout  = 8'b00111101; //  794 :  61 - 0x3d
      10'h31B: dout  = 8'b00101101; //  795 :  45 - 0x2d
      10'h31C: dout  = 8'b00101101; //  796 :  45 - 0x2d
      10'h31D: dout  = 8'b00101101; //  797 :  45 - 0x2d
      10'h31E: dout  = 8'b00100000; //  798 :  32 - 0x20
      10'h31F: dout  = 8'b00100000; //  799 :  32 - 0x20
      10'h320: dout  = 8'b00101101; //  800 :  45 - 0x2d -- line 0x19
      10'h321: dout  = 8'b00010001; //  801 :  17 - 0x11
      10'h322: dout  = 8'b00000011; //  802 :   3 - 0x3
      10'h323: dout  = 8'b00000011; //  803 :   3 - 0x3
      10'h324: dout  = 8'b00000011; //  804 :   3 - 0x3
      10'h325: dout  = 8'b00000011; //  805 :   3 - 0x3
      10'h326: dout  = 8'b00000011; //  806 :   3 - 0x3
      10'h327: dout  = 8'b00010001; //  807 :  17 - 0x11
      10'h328: dout  = 8'b00000011; //  808 :   3 - 0x3
      10'h329: dout  = 8'b00000011; //  809 :   3 - 0x3
      10'h32A: dout  = 8'b00000011; //  810 :   3 - 0x3
      10'h32B: dout  = 8'b00010001; //  811 :  17 - 0x11
      10'h32C: dout  = 8'b00000011; //  812 :   3 - 0x3
      10'h32D: dout  = 8'b00000011; //  813 :   3 - 0x3
      10'h32E: dout  = 8'b00000011; //  814 :   3 - 0x3
      10'h32F: dout  = 8'b00010001; //  815 :  17 - 0x11
      10'h330: dout  = 8'b00000011; //  816 :   3 - 0x3
      10'h331: dout  = 8'b00000011; //  817 :   3 - 0x3
      10'h332: dout  = 8'b00000011; //  818 :   3 - 0x3
      10'h333: dout  = 8'b00000011; //  819 :   3 - 0x3
      10'h334: dout  = 8'b00000011; //  820 :   3 - 0x3
      10'h335: dout  = 8'b00010001; //  821 :  17 - 0x11
      10'h336: dout  = 8'b00100000; //  822 :  32 - 0x20
      10'h337: dout  = 8'b00111110; //  823 :  62 - 0x3e
      10'h338: dout  = 8'b00111111; //  824 :  63 - 0x3f
      10'h339: dout  = 8'b00111110; //  825 :  62 - 0x3e
      10'h33A: dout  = 8'b00111111; //  826 :  63 - 0x3f
      10'h33B: dout  = 8'b00101101; //  827 :  45 - 0x2d
      10'h33C: dout  = 8'b00101101; //  828 :  45 - 0x2d
      10'h33D: dout  = 8'b00101101; //  829 :  45 - 0x2d
      10'h33E: dout  = 8'b00100000; //  830 :  32 - 0x20
      10'h33F: dout  = 8'b00100000; //  831 :  32 - 0x20
      10'h340: dout  = 8'b00101101; //  832 :  45 - 0x2d -- line 0x1a
      10'h341: dout  = 8'b00010001; //  833 :  17 - 0x11
      10'h342: dout  = 8'b00000011; //  834 :   3 - 0x3
      10'h343: dout  = 8'b00011001; //  835 :  25 - 0x19
      10'h344: dout  = 8'b00010000; //  836 :  16 - 0x10
      10'h345: dout  = 8'b00010000; //  837 :  16 - 0x10
      10'h346: dout  = 8'b00010000; //  838 :  16 - 0x10
      10'h347: dout  = 8'b00010010; //  839 :  18 - 0x12
      10'h348: dout  = 8'b00010000; //  840 :  16 - 0x10
      10'h349: dout  = 8'b00011000; //  841 :  24 - 0x18
      10'h34A: dout  = 8'b00000011; //  842 :   3 - 0x3
      10'h34B: dout  = 8'b00011010; //  843 :  26 - 0x1a
      10'h34C: dout  = 8'b00000011; //  844 :   3 - 0x3
      10'h34D: dout  = 8'b00011001; //  845 :  25 - 0x19
      10'h34E: dout  = 8'b00010000; //  846 :  16 - 0x10
      10'h34F: dout  = 8'b00010010; //  847 :  18 - 0x12
      10'h350: dout  = 8'b00010000; //  848 :  16 - 0x10
      10'h351: dout  = 8'b00010000; //  849 :  16 - 0x10
      10'h352: dout  = 8'b00010000; //  850 :  16 - 0x10
      10'h353: dout  = 8'b00011000; //  851 :  24 - 0x18
      10'h354: dout  = 8'b00000011; //  852 :   3 - 0x3
      10'h355: dout  = 8'b00010001; //  853 :  17 - 0x11
      10'h356: dout  = 8'b00100000; //  854 :  32 - 0x20
      10'h357: dout  = 8'b00100000; //  855 :  32 - 0x20
      10'h358: dout  = 8'b00100000; //  856 :  32 - 0x20
      10'h359: dout  = 8'b00100000; //  857 :  32 - 0x20
      10'h35A: dout  = 8'b00100000; //  858 :  32 - 0x20
      10'h35B: dout  = 8'b00100000; //  859 :  32 - 0x20
      10'h35C: dout  = 8'b00101101; //  860 :  45 - 0x2d
      10'h35D: dout  = 8'b00101101; //  861 :  45 - 0x2d
      10'h35E: dout  = 8'b00100000; //  862 :  32 - 0x20
      10'h35F: dout  = 8'b00100000; //  863 :  32 - 0x20
      10'h360: dout  = 8'b00101101; //  864 :  45 - 0x2d -- line 0x1b
      10'h361: dout  = 8'b00010001; //  865 :  17 - 0x11
      10'h362: dout  = 8'b00000011; //  866 :   3 - 0x3
      10'h363: dout  = 8'b00000011; //  867 :   3 - 0x3
      10'h364: dout  = 8'b00000011; //  868 :   3 - 0x3
      10'h365: dout  = 8'b00000011; //  869 :   3 - 0x3
      10'h366: dout  = 8'b00000011; //  870 :   3 - 0x3
      10'h367: dout  = 8'b00000011; //  871 :   3 - 0x3
      10'h368: dout  = 8'b00000011; //  872 :   3 - 0x3
      10'h369: dout  = 8'b00000011; //  873 :   3 - 0x3
      10'h36A: dout  = 8'b00000011; //  874 :   3 - 0x3
      10'h36B: dout  = 8'b00000011; //  875 :   3 - 0x3
      10'h36C: dout  = 8'b00000011; //  876 :   3 - 0x3
      10'h36D: dout  = 8'b00000011; //  877 :   3 - 0x3
      10'h36E: dout  = 8'b00000011; //  878 :   3 - 0x3
      10'h36F: dout  = 8'b00000011; //  879 :   3 - 0x3
      10'h370: dout  = 8'b00000011; //  880 :   3 - 0x3
      10'h371: dout  = 8'b00000011; //  881 :   3 - 0x3
      10'h372: dout  = 8'b00000011; //  882 :   3 - 0x3
      10'h373: dout  = 8'b00000011; //  883 :   3 - 0x3
      10'h374: dout  = 8'b00000011; //  884 :   3 - 0x3
      10'h375: dout  = 8'b00010001; //  885 :  17 - 0x11
      10'h376: dout  = 8'b00100000; //  886 :  32 - 0x20
      10'h377: dout  = 8'b00100000; //  887 :  32 - 0x20
      10'h378: dout  = 8'b00100000; //  888 :  32 - 0x20
      10'h379: dout  = 8'b00100000; //  889 :  32 - 0x20
      10'h37A: dout  = 8'b00100000; //  890 :  32 - 0x20
      10'h37B: dout  = 8'b00100000; //  891 :  32 - 0x20
      10'h37C: dout  = 8'b00101101; //  892 :  45 - 0x2d
      10'h37D: dout  = 8'b00101101; //  893 :  45 - 0x2d
      10'h37E: dout  = 8'b00100000; //  894 :  32 - 0x20
      10'h37F: dout  = 8'b00100000; //  895 :  32 - 0x20
      10'h380: dout  = 8'b00101101; //  896 :  45 - 0x2d -- line 0x1c
      10'h381: dout  = 8'b00011110; //  897 :  30 - 0x1e
      10'h382: dout  = 8'b00010000; //  898 :  16 - 0x10
      10'h383: dout  = 8'b00010000; //  899 :  16 - 0x10
      10'h384: dout  = 8'b00010000; //  900 :  16 - 0x10
      10'h385: dout  = 8'b00010000; //  901 :  16 - 0x10
      10'h386: dout  = 8'b00010000; //  902 :  16 - 0x10
      10'h387: dout  = 8'b00010000; //  903 :  16 - 0x10
      10'h388: dout  = 8'b00010000; //  904 :  16 - 0x10
      10'h389: dout  = 8'b00010000; //  905 :  16 - 0x10
      10'h38A: dout  = 8'b00010000; //  906 :  16 - 0x10
      10'h38B: dout  = 8'b00010000; //  907 :  16 - 0x10
      10'h38C: dout  = 8'b00010000; //  908 :  16 - 0x10
      10'h38D: dout  = 8'b00010000; //  909 :  16 - 0x10
      10'h38E: dout  = 8'b00010000; //  910 :  16 - 0x10
      10'h38F: dout  = 8'b00010000; //  911 :  16 - 0x10
      10'h390: dout  = 8'b00010000; //  912 :  16 - 0x10
      10'h391: dout  = 8'b00010000; //  913 :  16 - 0x10
      10'h392: dout  = 8'b00010000; //  914 :  16 - 0x10
      10'h393: dout  = 8'b00010000; //  915 :  16 - 0x10
      10'h394: dout  = 8'b00010000; //  916 :  16 - 0x10
      10'h395: dout  = 8'b00011100; //  917 :  28 - 0x1c
      10'h396: dout  = 8'b00100000; //  918 :  32 - 0x20
      10'h397: dout  = 8'b00100000; //  919 :  32 - 0x20
      10'h398: dout  = 8'b00100000; //  920 :  32 - 0x20
      10'h399: dout  = 8'b00100000; //  921 :  32 - 0x20
      10'h39A: dout  = 8'b00100000; //  922 :  32 - 0x20
      10'h39B: dout  = 8'b00100000; //  923 :  32 - 0x20
      10'h39C: dout  = 8'b00100000; //  924 :  32 - 0x20
      10'h39D: dout  = 8'b00100000; //  925 :  32 - 0x20
      10'h39E: dout  = 8'b00100000; //  926 :  32 - 0x20
      10'h39F: dout  = 8'b00100000; //  927 :  32 - 0x20
      10'h3A0: dout  = 8'b00100000; //  928 :  32 - 0x20 -- line 0x1d
      10'h3A1: dout  = 8'b00100000; //  929 :  32 - 0x20
      10'h3A2: dout  = 8'b00100000; //  930 :  32 - 0x20
      10'h3A3: dout  = 8'b00100000; //  931 :  32 - 0x20
      10'h3A4: dout  = 8'b00100000; //  932 :  32 - 0x20
      10'h3A5: dout  = 8'b00100000; //  933 :  32 - 0x20
      10'h3A6: dout  = 8'b00100000; //  934 :  32 - 0x20
      10'h3A7: dout  = 8'b00100000; //  935 :  32 - 0x20
      10'h3A8: dout  = 8'b00100000; //  936 :  32 - 0x20
      10'h3A9: dout  = 8'b00100000; //  937 :  32 - 0x20
      10'h3AA: dout  = 8'b00100000; //  938 :  32 - 0x20
      10'h3AB: dout  = 8'b00100000; //  939 :  32 - 0x20
      10'h3AC: dout  = 8'b00100000; //  940 :  32 - 0x20
      10'h3AD: dout  = 8'b00100000; //  941 :  32 - 0x20
      10'h3AE: dout  = 8'b00100000; //  942 :  32 - 0x20
      10'h3AF: dout  = 8'b00100000; //  943 :  32 - 0x20
      10'h3B0: dout  = 8'b00100000; //  944 :  32 - 0x20
      10'h3B1: dout  = 8'b00100000; //  945 :  32 - 0x20
      10'h3B2: dout  = 8'b00100000; //  946 :  32 - 0x20
      10'h3B3: dout  = 8'b00100000; //  947 :  32 - 0x20
      10'h3B4: dout  = 8'b00100000; //  948 :  32 - 0x20
      10'h3B5: dout  = 8'b00100000; //  949 :  32 - 0x20
      10'h3B6: dout  = 8'b00100000; //  950 :  32 - 0x20
      10'h3B7: dout  = 8'b00100000; //  951 :  32 - 0x20
      10'h3B8: dout  = 8'b00100000; //  952 :  32 - 0x20
      10'h3B9: dout  = 8'b00100000; //  953 :  32 - 0x20
      10'h3BA: dout  = 8'b00100000; //  954 :  32 - 0x20
      10'h3BB: dout  = 8'b00100000; //  955 :  32 - 0x20
      10'h3BC: dout  = 8'b00100000; //  956 :  32 - 0x20
      10'h3BD: dout  = 8'b00100000; //  957 :  32 - 0x20
      10'h3BE: dout  = 8'b00100000; //  958 :  32 - 0x20
      10'h3BF: dout  = 8'b00100000; //  959 :  32 - 0x20
        //-- Attribute Table 0----
      10'h3C0: dout  = 8'b01010101; //  960 :  85 - 0x55
      10'h3C1: dout  = 8'b01010101; //  961 :  85 - 0x55
      10'h3C2: dout  = 8'b01010101; //  962 :  85 - 0x55
      10'h3C3: dout  = 8'b01010101; //  963 :  85 - 0x55
      10'h3C4: dout  = 8'b01010101; //  964 :  85 - 0x55
      10'h3C5: dout  = 8'b00010001; //  965 :  17 - 0x11
      10'h3C6: dout  = 8'b00000000; //  966 :   0 - 0x0
      10'h3C7: dout  = 8'b00000000; //  967 :   0 - 0x0
      10'h3C8: dout  = 8'b01010101; //  968 :  85 - 0x55
      10'h3C9: dout  = 8'b01010101; //  969 :  85 - 0x55
      10'h3CA: dout  = 8'b01010101; //  970 :  85 - 0x55
      10'h3CB: dout  = 8'b01010101; //  971 :  85 - 0x55
      10'h3CC: dout  = 8'b01010101; //  972 :  85 - 0x55
      10'h3CD: dout  = 8'b00010001; //  973 :  17 - 0x11
      10'h3CE: dout  = 8'b00000000; //  974 :   0 - 0x0
      10'h3CF: dout  = 8'b00000000; //  975 :   0 - 0x0
      10'h3D0: dout  = 8'b01010101; //  976 :  85 - 0x55
      10'h3D1: dout  = 8'b01010101; //  977 :  85 - 0x55
      10'h3D2: dout  = 8'b01010101; //  978 :  85 - 0x55
      10'h3D3: dout  = 8'b01010101; //  979 :  85 - 0x55
      10'h3D4: dout  = 8'b01010101; //  980 :  85 - 0x55
      10'h3D5: dout  = 8'b00010001; //  981 :  17 - 0x11
      10'h3D6: dout  = 8'b00000000; //  982 :   0 - 0x0
      10'h3D7: dout  = 8'b00000000; //  983 :   0 - 0x0
      10'h3D8: dout  = 8'b01010101; //  984 :  85 - 0x55
      10'h3D9: dout  = 8'b01010101; //  985 :  85 - 0x55
      10'h3DA: dout  = 8'b01010101; //  986 :  85 - 0x55
      10'h3DB: dout  = 8'b01010101; //  987 :  85 - 0x55
      10'h3DC: dout  = 8'b01010101; //  988 :  85 - 0x55
      10'h3DD: dout  = 8'b01010001; //  989 :  81 - 0x51
      10'h3DE: dout  = 8'b01010000; //  990 :  80 - 0x50
      10'h3DF: dout  = 8'b01010000; //  991 :  80 - 0x50
      10'h3E0: dout  = 8'b01010101; //  992 :  85 - 0x55
      10'h3E1: dout  = 8'b01010101; //  993 :  85 - 0x55
      10'h3E2: dout  = 8'b01010101; //  994 :  85 - 0x55
      10'h3E3: dout  = 8'b01010101; //  995 :  85 - 0x55
      10'h3E4: dout  = 8'b01010101; //  996 :  85 - 0x55
      10'h3E5: dout  = 8'b10010101; //  997 : 149 - 0x95
      10'h3E6: dout  = 8'b00000101; //  998 :   5 - 0x5
      10'h3E7: dout  = 8'b00000101; //  999 :   5 - 0x5
      10'h3E8: dout  = 8'b01010101; // 1000 :  85 - 0x55
      10'h3E9: dout  = 8'b01010101; // 1001 :  85 - 0x55
      10'h3EA: dout  = 8'b01010101; // 1002 :  85 - 0x55
      10'h3EB: dout  = 8'b01010101; // 1003 :  85 - 0x55
      10'h3EC: dout  = 8'b01010101; // 1004 :  85 - 0x55
      10'h3ED: dout  = 8'b00010001; // 1005 :  17 - 0x11
      10'h3EE: dout  = 8'b00000000; // 1006 :   0 - 0x0
      10'h3EF: dout  = 8'b00000000; // 1007 :   0 - 0x0
      10'h3F0: dout  = 8'b01010101; // 1008 :  85 - 0x55
      10'h3F1: dout  = 8'b01010101; // 1009 :  85 - 0x55
      10'h3F2: dout  = 8'b01010101; // 1010 :  85 - 0x55
      10'h3F3: dout  = 8'b01010101; // 1011 :  85 - 0x55
      10'h3F4: dout  = 8'b01010101; // 1012 :  85 - 0x55
      10'h3F5: dout  = 8'b01010101; // 1013 :  85 - 0x55
      10'h3F6: dout  = 8'b01010101; // 1014 :  85 - 0x55
      10'h3F7: dout  = 8'b01010101; // 1015 :  85 - 0x55
      10'h3F8: dout  = 8'b01010101; // 1016 :  85 - 0x55
      10'h3F9: dout  = 8'b01010101; // 1017 :  85 - 0x55
      10'h3FA: dout  = 8'b01010101; // 1018 :  85 - 0x55
      10'h3FB: dout  = 8'b01010101; // 1019 :  85 - 0x55
      10'h3FC: dout  = 8'b01010101; // 1020 :  85 - 0x55
      10'h3FD: dout  = 8'b01010101; // 1021 :  85 - 0x55
      10'h3FE: dout  = 8'b01010101; // 1022 :  85 - 0x55
      10'h3FF: dout  = 8'b01010101; // 1023 :  85 - 0x55
    endcase
  end

endmodule
