---   Sprites Pattern table COLOR PLANE 1
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
--- Autcmatically generated VHDL ROM from a NES memory file----


---  Original memory dump file name: smario_traspas_patron.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_MARIO_TRASPAS_SPR_PLN1 is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(11-1 downto 0);  --2048 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_MARIO_TRASPAS_SPR_PLN1;

architecture BEHAVIORAL of ROM_PTABLE_MARIO_TRASPAS_SPR_PLN1 is
  signal addr_int  : natural range 0 to 2**11-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Sprite pattern Table COLOR PLANE 1
    "00000000", --    0 -  0x0  :    0 - 0x0 -- Sprite 0x0
    "00000000", --    1 -  0x1  :    0 - 0x0
    "00000000", --    2 -  0x2  :    0 - 0x0
    "00000000", --    3 -  0x3  :    0 - 0x0
    "00011111", --    4 -  0x4  :   31 - 0x1f
    "00111111", --    5 -  0x5  :   63 - 0x3f
    "00111111", --    6 -  0x6  :   63 - 0x3f
    "01111111", --    7 -  0x7  :  127 - 0x7f
    "00000000", --    8 -  0x8  :    0 - 0x0 -- Sprite 0x1
    "00100000", --    9 -  0x9  :   32 - 0x20
    "01100000", --   10 -  0xa  :   96 - 0x60
    "00000000", --   11 -  0xb  :    0 - 0x0
    "11110000", --   12 -  0xc  :  240 - 0xf0
    "11111100", --   13 -  0xd  :  252 - 0xfc
    "11111110", --   14 -  0xe  :  254 - 0xfe
    "11111110", --   15 -  0xf  :  254 - 0xfe
    "01111111", --   16 - 0x10  :  127 - 0x7f -- Sprite 0x2
    "01111111", --   17 - 0x11  :  127 - 0x7f
    "00011111", --   18 - 0x12  :   31 - 0x1f
    "00000111", --   19 - 0x13  :    7 - 0x7
    "00000000", --   20 - 0x14  :    0 - 0x0
    "00011110", --   21 - 0x15  :   30 - 0x1e
    "00111111", --   22 - 0x16  :   63 - 0x3f
    "01111111", --   23 - 0x17  :  127 - 0x7f
    "11111100", --   24 - 0x18  :  252 - 0xfc -- Sprite 0x3
    "11111100", --   25 - 0x19  :  252 - 0xfc
    "11111000", --   26 - 0x1a  :  248 - 0xf8
    "11000000", --   27 - 0x1b  :  192 - 0xc0
    "11000010", --   28 - 0x1c  :  194 - 0xc2
    "01100111", --   29 - 0x1d  :  103 - 0x67
    "00101111", --   30 - 0x1e  :   47 - 0x2f
    "00110111", --   31 - 0x1f  :   55 - 0x37
    "01111111", --   32 - 0x20  :  127 - 0x7f -- Sprite 0x4
    "01111110", --   33 - 0x21  :  126 - 0x7e
    "11111100", --   34 - 0x22  :  252 - 0xfc
    "11110000", --   35 - 0x23  :  240 - 0xf0
    "11111000", --   36 - 0x24  :  248 - 0xf8
    "11111000", --   37 - 0x25  :  248 - 0xf8
    "11110000", --   38 - 0x26  :  240 - 0xf0
    "01110000", --   39 - 0x27  :  112 - 0x70
    "00110111", --   40 - 0x28  :   55 - 0x37 -- Sprite 0x5
    "00110110", --   41 - 0x29  :   54 - 0x36
    "01011100", --   42 - 0x2a  :   92 - 0x5c
    "00000000", --   43 - 0x2b  :    0 - 0x0
    "00000000", --   44 - 0x2c  :    0 - 0x0
    "00000001", --   45 - 0x2d  :    1 - 0x1
    "00000011", --   46 - 0x2e  :    3 - 0x3
    "00011111", --   47 - 0x2f  :   31 - 0x1f
    "00001000", --   48 - 0x30  :    8 - 0x8 -- Sprite 0x6
    "00100100", --   49 - 0x31  :   36 - 0x24
    "11100011", --   50 - 0x32  :  227 - 0xe3
    "11110000", --   51 - 0x33  :  240 - 0xf0
    "11111000", --   52 - 0x34  :  248 - 0xf8
    "01110000", --   53 - 0x35  :  112 - 0x70
    "01110000", --   54 - 0x36  :  112 - 0x70
    "00111000", --   55 - 0x37  :   56 - 0x38
    "00011111", --   56 - 0x38  :   31 - 0x1f -- Sprite 0x7
    "00011111", --   57 - 0x39  :   31 - 0x1f
    "00011111", --   58 - 0x3a  :   31 - 0x1f
    "00011111", --   59 - 0x3b  :   31 - 0x1f
    "00000000", --   60 - 0x3c  :    0 - 0x0
    "00000000", --   61 - 0x3d  :    0 - 0x0
    "00000000", --   62 - 0x3e  :    0 - 0x0
    "00000000", --   63 - 0x3f  :    0 - 0x0
    "00000000", --   64 - 0x40  :    0 - 0x0 -- Sprite 0x8
    "00000000", --   65 - 0x41  :    0 - 0x0
    "00000000", --   66 - 0x42  :    0 - 0x0
    "00000000", --   67 - 0x43  :    0 - 0x0
    "00000000", --   68 - 0x44  :    0 - 0x0
    "00000000", --   69 - 0x45  :    0 - 0x0
    "00001111", --   70 - 0x46  :   15 - 0xf
    "00011111", --   71 - 0x47  :   31 - 0x1f
    "00000000", --   72 - 0x48  :    0 - 0x0 -- Sprite 0x9
    "00000000", --   73 - 0x49  :    0 - 0x0
    "00000000", --   74 - 0x4a  :    0 - 0x0
    "00010000", --   75 - 0x4b  :   16 - 0x10
    "00110000", --   76 - 0x4c  :   48 - 0x30
    "00000000", --   77 - 0x4d  :    0 - 0x0
    "11111000", --   78 - 0x4e  :  248 - 0xf8
    "11111110", --   79 - 0x4f  :  254 - 0xfe
    "00011111", --   80 - 0x50  :   31 - 0x1f -- Sprite 0xa
    "00111111", --   81 - 0x51  :   63 - 0x3f
    "00111111", --   82 - 0x52  :   63 - 0x3f
    "00011111", --   83 - 0x53  :   31 - 0x1f
    "00000111", --   84 - 0x54  :    7 - 0x7
    "00001000", --   85 - 0x55  :    8 - 0x8
    "00010111", --   86 - 0x56  :   23 - 0x17
    "00010111", --   87 - 0x57  :   23 - 0x17
    "11111111", --   88 - 0x58  :  255 - 0xff -- Sprite 0xb
    "11111111", --   89 - 0x59  :  255 - 0xff
    "11111110", --   90 - 0x5a  :  254 - 0xfe
    "11111110", --   91 - 0x5b  :  254 - 0xfe
    "11111100", --   92 - 0x5c  :  252 - 0xfc
    "11100000", --   93 - 0x5d  :  224 - 0xe0
    "01000000", --   94 - 0x5e  :   64 - 0x40
    "10100000", --   95 - 0x5f  :  160 - 0xa0
    "00110111", --   96 - 0x60  :   55 - 0x37 -- Sprite 0xc
    "00100111", --   97 - 0x61  :   39 - 0x27
    "00100011", --   98 - 0x62  :   35 - 0x23
    "00000011", --   99 - 0x63  :    3 - 0x3
    "00000001", --  100 - 0x64  :    1 - 0x1
    "00000000", --  101 - 0x65  :    0 - 0x0
    "00000000", --  102 - 0x66  :    0 - 0x0
    "00000000", --  103 - 0x67  :    0 - 0x0
    "11001100", --  104 - 0x68  :  204 - 0xcc -- Sprite 0xd
    "11111111", --  105 - 0x69  :  255 - 0xff
    "11111111", --  106 - 0x6a  :  255 - 0xff
    "11111111", --  107 - 0x6b  :  255 - 0xff
    "11111111", --  108 - 0x6c  :  255 - 0xff
    "01110000", --  109 - 0x6d  :  112 - 0x70
    "00000000", --  110 - 0x6e  :    0 - 0x0
    "00001000", --  111 - 0x6f  :    8 - 0x8
    "11110000", --  112 - 0x70  :  240 - 0xf0 -- Sprite 0xe
    "11110000", --  113 - 0x71  :  240 - 0xf0
    "11110000", --  114 - 0x72  :  240 - 0xf0
    "11110000", --  115 - 0x73  :  240 - 0xf0
    "11110000", --  116 - 0x74  :  240 - 0xf0
    "11000000", --  117 - 0x75  :  192 - 0xc0
    "10000000", --  118 - 0x76  :  128 - 0x80
    "00000000", --  119 - 0x77  :    0 - 0x0
    "00010000", --  120 - 0x78  :   16 - 0x10 -- Sprite 0xf
    "01100000", --  121 - 0x79  :   96 - 0x60
    "10000000", --  122 - 0x7a  :  128 - 0x80
    "00000000", --  123 - 0x7b  :    0 - 0x0
    "01111000", --  124 - 0x7c  :  120 - 0x78
    "01111000", --  125 - 0x7d  :  120 - 0x78
    "01111110", --  126 - 0x7e  :  126 - 0x7e
    "01111110", --  127 - 0x7f  :  126 - 0x7e
    "00000000", --  128 - 0x80  :    0 - 0x0 -- Sprite 0x10
    "00000000", --  129 - 0x81  :    0 - 0x0
    "00000000", --  130 - 0x82  :    0 - 0x0
    "00000000", --  131 - 0x83  :    0 - 0x0
    "00000000", --  132 - 0x84  :    0 - 0x0
    "00011111", --  133 - 0x85  :   31 - 0x1f
    "00111111", --  134 - 0x86  :   63 - 0x3f
    "00111111", --  135 - 0x87  :   63 - 0x3f
    "00000000", --  136 - 0x88  :    0 - 0x0 -- Sprite 0x11
    "00000000", --  137 - 0x89  :    0 - 0x0
    "00100000", --  138 - 0x8a  :   32 - 0x20
    "01100000", --  139 - 0x8b  :   96 - 0x60
    "00000000", --  140 - 0x8c  :    0 - 0x0
    "11110000", --  141 - 0x8d  :  240 - 0xf0
    "11111100", --  142 - 0x8e  :  252 - 0xfc
    "11111110", --  143 - 0x8f  :  254 - 0xfe
    "01111111", --  144 - 0x90  :  127 - 0x7f -- Sprite 0x12
    "01111111", --  145 - 0x91  :  127 - 0x7f
    "00111111", --  146 - 0x92  :   63 - 0x3f
    "00011111", --  147 - 0x93  :   31 - 0x1f
    "00000000", --  148 - 0x94  :    0 - 0x0
    "00010110", --  149 - 0x95  :   22 - 0x16
    "00101111", --  150 - 0x96  :   47 - 0x2f
    "00101111", --  151 - 0x97  :   47 - 0x2f
    "11111110", --  152 - 0x98  :  254 - 0xfe -- Sprite 0x13
    "11111100", --  153 - 0x99  :  252 - 0xfc
    "11111100", --  154 - 0x9a  :  252 - 0xfc
    "11111000", --  155 - 0x9b  :  248 - 0xf8
    "11000000", --  156 - 0x9c  :  192 - 0xc0
    "01100000", --  157 - 0x9d  :   96 - 0x60
    "00100000", --  158 - 0x9e  :   32 - 0x20
    "00110000", --  159 - 0x9f  :   48 - 0x30
    "00101111", --  160 - 0xa0  :   47 - 0x2f -- Sprite 0x14
    "00101111", --  161 - 0xa1  :   47 - 0x2f
    "00101111", --  162 - 0xa2  :   47 - 0x2f
    "00001111", --  163 - 0xa3  :   15 - 0xf
    "00000111", --  164 - 0xa4  :    7 - 0x7
    "00000011", --  165 - 0xa5  :    3 - 0x3
    "00000000", --  166 - 0xa6  :    0 - 0x0
    "00000000", --  167 - 0xa7  :    0 - 0x0
    "00010000", --  168 - 0xa8  :   16 - 0x10 -- Sprite 0x15
    "11110000", --  169 - 0xa9  :  240 - 0xf0
    "11110000", --  170 - 0xaa  :  240 - 0xf0
    "11110000", --  171 - 0xab  :  240 - 0xf0
    "11110000", --  172 - 0xac  :  240 - 0xf0
    "11100000", --  173 - 0xad  :  224 - 0xe0
    "11000000", --  174 - 0xae  :  192 - 0xc0
    "11100000", --  175 - 0xaf  :  224 - 0xe0
    "00000001", --  176 - 0xb0  :    1 - 0x1 -- Sprite 0x16
    "00000011", --  177 - 0xb1  :    3 - 0x3
    "00000001", --  178 - 0xb2  :    1 - 0x1
    "00000100", --  179 - 0xb3  :    4 - 0x4
    "00000111", --  180 - 0xb4  :    7 - 0x7
    "00001111", --  181 - 0xb5  :   15 - 0xf
    "00001111", --  182 - 0xb6  :   15 - 0xf
    "00000011", --  183 - 0xb7  :    3 - 0x3
    "11111000", --  184 - 0xb8  :  248 - 0xf8 -- Sprite 0x17
    "11110000", --  185 - 0xb9  :  240 - 0xf0
    "11100000", --  186 - 0xba  :  224 - 0xe0
    "01110000", --  187 - 0xbb  :  112 - 0x70
    "10110000", --  188 - 0xbc  :  176 - 0xb0
    "10000000", --  189 - 0xbd  :  128 - 0x80
    "11100000", --  190 - 0xbe  :  224 - 0xe0
    "11100000", --  191 - 0xbf  :  224 - 0xe0
    "00000000", --  192 - 0xc0  :    0 - 0x0 -- Sprite 0x18
    "00110000", --  193 - 0xc1  :   48 - 0x30
    "01110000", --  194 - 0xc2  :  112 - 0x70
    "01111111", --  195 - 0xc3  :  127 - 0x7f
    "11111111", --  196 - 0xc4  :  255 - 0xff
    "11111111", --  197 - 0xc5  :  255 - 0xff
    "11110111", --  198 - 0xc6  :  247 - 0xf7
    "11110011", --  199 - 0xc7  :  243 - 0xf3
    "00000000", --  200 - 0xc8  :    0 - 0x0 -- Sprite 0x19
    "00011000", --  201 - 0xc9  :   24 - 0x18
    "00010000", --  202 - 0xca  :   16 - 0x10
    "00000000", --  203 - 0xcb  :    0 - 0x0
    "11111000", --  204 - 0xcc  :  248 - 0xf8
    "11111000", --  205 - 0xcd  :  248 - 0xf8
    "11111110", --  206 - 0xce  :  254 - 0xfe
    "11111111", --  207 - 0xcf  :  255 - 0xff
    "11100111", --  208 - 0xd0  :  231 - 0xe7 -- Sprite 0x1a
    "00001111", --  209 - 0xd1  :   15 - 0xf
    "00001111", --  210 - 0xd2  :   15 - 0xf
    "00011111", --  211 - 0xd3  :   31 - 0x1f
    "00011111", --  212 - 0xd4  :   31 - 0x1f
    "00011111", --  213 - 0xd5  :   31 - 0x1f
    "00001111", --  214 - 0xd6  :   15 - 0xf
    "00000111", --  215 - 0xd7  :    7 - 0x7
    "11111111", --  216 - 0xd8  :  255 - 0xff -- Sprite 0x1b
    "11111110", --  217 - 0xd9  :  254 - 0xfe
    "11111100", --  218 - 0xda  :  252 - 0xfc
    "11000110", --  219 - 0xdb  :  198 - 0xc6
    "10001110", --  220 - 0xdc  :  142 - 0x8e
    "11101110", --  221 - 0xdd  :  238 - 0xee
    "11111111", --  222 - 0xde  :  255 - 0xff
    "11111111", --  223 - 0xdf  :  255 - 0xff
    "00000011", --  224 - 0xe0  :    3 - 0x3 -- Sprite 0x1c
    "00000000", --  225 - 0xe1  :    0 - 0x0
    "00000000", --  226 - 0xe2  :    0 - 0x0
    "00001110", --  227 - 0xe3  :   14 - 0xe
    "00000111", --  228 - 0xe4  :    7 - 0x7
    "00111111", --  229 - 0xe5  :   63 - 0x3f
    "00111111", --  230 - 0xe6  :   63 - 0x3f
    "00111111", --  231 - 0xe7  :   63 - 0x3f
    "11111111", --  232 - 0xe8  :  255 - 0xff -- Sprite 0x1d
    "01111111", --  233 - 0xe9  :  127 - 0x7f
    "00111111", --  234 - 0xea  :   63 - 0x3f
    "00001110", --  235 - 0xeb  :   14 - 0xe
    "11000000", --  236 - 0xec  :  192 - 0xc0
    "11000000", --  237 - 0xed  :  192 - 0xc0
    "11100000", --  238 - 0xee  :  224 - 0xe0
    "11100000", --  239 - 0xef  :  224 - 0xe0
    "00000000", --  240 - 0xf0  :    0 - 0x0 -- Sprite 0x1e
    "10000000", --  241 - 0xf1  :  128 - 0x80
    "11001000", --  242 - 0xf2  :  200 - 0xc8
    "11111110", --  243 - 0xf3  :  254 - 0xfe
    "01111111", --  244 - 0xf4  :  127 - 0x7f
    "00111111", --  245 - 0xf5  :   63 - 0x3f
    "00011110", --  246 - 0xf6  :   30 - 0x1e
    "00001110", --  247 - 0xf7  :   14 - 0xe
    "11100000", --  248 - 0xf8  :  224 - 0xe0 -- Sprite 0x1f
    "00000000", --  249 - 0xf9  :    0 - 0x0
    "00000000", --  250 - 0xfa  :    0 - 0x0
    "00000000", --  251 - 0xfb  :    0 - 0x0
    "00000000", --  252 - 0xfc  :    0 - 0x0
    "00000000", --  253 - 0xfd  :    0 - 0x0
    "00000000", --  254 - 0xfe  :    0 - 0x0
    "00000000", --  255 - 0xff  :    0 - 0x0
    "00000000", --  256 - 0x100  :    0 - 0x0 -- Sprite 0x20
    "00000000", --  257 - 0x101  :    0 - 0x0
    "00000000", --  258 - 0x102  :    0 - 0x0
    "00000000", --  259 - 0x103  :    0 - 0x0
    "00000000", --  260 - 0x104  :    0 - 0x0
    "00000000", --  261 - 0x105  :    0 - 0x0
    "00011111", --  262 - 0x106  :   31 - 0x1f
    "00111111", --  263 - 0x107  :   63 - 0x3f
    "00001110", --  264 - 0x108  :   14 - 0xe -- Sprite 0x21
    "00011111", --  265 - 0x109  :   31 - 0x1f
    "00011111", --  266 - 0x10a  :   31 - 0x1f
    "00011111", --  267 - 0x10b  :   31 - 0x1f
    "00011111", --  268 - 0x10c  :   31 - 0x1f
    "00000011", --  269 - 0x10d  :    3 - 0x3
    "11111111", --  270 - 0x10e  :  255 - 0xff
    "11111111", --  271 - 0x10f  :  255 - 0xff
    "00111111", --  272 - 0x110  :   63 - 0x3f -- Sprite 0x22
    "00111111", --  273 - 0x111  :   63 - 0x3f
    "01111111", --  274 - 0x112  :  127 - 0x7f
    "01111111", --  275 - 0x113  :  127 - 0x7f
    "00011111", --  276 - 0x114  :   31 - 0x1f
    "00000000", --  277 - 0x115  :    0 - 0x0
    "01111110", --  278 - 0x116  :  126 - 0x7e
    "11111111", --  279 - 0x117  :  255 - 0xff
    "11111111", --  280 - 0x118  :  255 - 0xff -- Sprite 0x23
    "11111111", --  281 - 0x119  :  255 - 0xff
    "11111110", --  282 - 0x11a  :  254 - 0xfe
    "11111110", --  283 - 0x11b  :  254 - 0xfe
    "11111110", --  284 - 0x11c  :  254 - 0xfe
    "11011110", --  285 - 0x11d  :  222 - 0xde
    "01011100", --  286 - 0x11e  :   92 - 0x5c
    "01101100", --  287 - 0x11f  :  108 - 0x6c
    "11111111", --  288 - 0x120  :  255 - 0xff -- Sprite 0x24
    "11111111", --  289 - 0x121  :  255 - 0xff
    "11111110", --  290 - 0x122  :  254 - 0xfe
    "11111100", --  291 - 0x123  :  252 - 0xfc
    "11111000", --  292 - 0x124  :  248 - 0xf8
    "10110000", --  293 - 0x125  :  176 - 0xb0
    "01100000", --  294 - 0x126  :   96 - 0x60
    "00000000", --  295 - 0x127  :    0 - 0x0
    "00101000", --  296 - 0x128  :   40 - 0x28 -- Sprite 0x25
    "00110000", --  297 - 0x129  :   48 - 0x30
    "00011000", --  298 - 0x12a  :   24 - 0x18
    "01000000", --  299 - 0x12b  :   64 - 0x40
    "00000000", --  300 - 0x12c  :    0 - 0x0
    "00000001", --  301 - 0x12d  :    1 - 0x1
    "00000011", --  302 - 0x12e  :    3 - 0x3
    "00001111", --  303 - 0x12f  :   15 - 0xf
    "00010000", --  304 - 0x130  :   16 - 0x10 -- Sprite 0x26
    "11101100", --  305 - 0x131  :  236 - 0xec
    "11100011", --  306 - 0x132  :  227 - 0xe3
    "11100000", --  307 - 0x133  :  224 - 0xe0
    "11100000", --  308 - 0x134  :  224 - 0xe0
    "11100000", --  309 - 0x135  :  224 - 0xe0
    "11000000", --  310 - 0x136  :  192 - 0xc0
    "10000000", --  311 - 0x137  :  128 - 0x80
    "00001111", --  312 - 0x138  :   15 - 0xf -- Sprite 0x27
    "00001111", --  313 - 0x139  :   15 - 0xf
    "00001111", --  314 - 0x13a  :   15 - 0xf
    "00001111", --  315 - 0x13b  :   15 - 0xf
    "00000000", --  316 - 0x13c  :    0 - 0x0
    "00000000", --  317 - 0x13d  :    0 - 0x0
    "00000000", --  318 - 0x13e  :    0 - 0x0
    "00000000", --  319 - 0x13f  :    0 - 0x0
    "00011111", --  320 - 0x140  :   31 - 0x1f -- Sprite 0x28
    "00111111", --  321 - 0x141  :   63 - 0x3f
    "00111111", --  322 - 0x142  :   63 - 0x3f
    "00011111", --  323 - 0x143  :   31 - 0x1f
    "00000111", --  324 - 0x144  :    7 - 0x7
    "00001001", --  325 - 0x145  :    9 - 0x9
    "00010011", --  326 - 0x146  :   19 - 0x13
    "00010111", --  327 - 0x147  :   23 - 0x17
    "11111111", --  328 - 0x148  :  255 - 0xff -- Sprite 0x29
    "11111111", --  329 - 0x149  :  255 - 0xff
    "11111110", --  330 - 0x14a  :  254 - 0xfe
    "11111111", --  331 - 0x14b  :  255 - 0xff
    "11111110", --  332 - 0x14c  :  254 - 0xfe
    "11111100", --  333 - 0x14d  :  252 - 0xfc
    "11111000", --  334 - 0x14e  :  248 - 0xf8
    "11100000", --  335 - 0x14f  :  224 - 0xe0
    "00010111", --  336 - 0x150  :   23 - 0x17 -- Sprite 0x2a
    "00010111", --  337 - 0x151  :   23 - 0x17
    "00000011", --  338 - 0x152  :    3 - 0x3
    "00000000", --  339 - 0x153  :    0 - 0x0
    "00000000", --  340 - 0x154  :    0 - 0x0
    "00000000", --  341 - 0x155  :    0 - 0x0
    "00000000", --  342 - 0x156  :    0 - 0x0
    "00000000", --  343 - 0x157  :    0 - 0x0
    "11010000", --  344 - 0x158  :  208 - 0xd0 -- Sprite 0x2b
    "10010000", --  345 - 0x159  :  144 - 0x90
    "00011000", --  346 - 0x15a  :   24 - 0x18
    "00001000", --  347 - 0x15b  :    8 - 0x8
    "01000000", --  348 - 0x15c  :   64 - 0x40
    "00000000", --  349 - 0x15d  :    0 - 0x0
    "00000000", --  350 - 0x15e  :    0 - 0x0
    "00000000", --  351 - 0x15f  :    0 - 0x0
    "00110000", --  352 - 0x160  :   48 - 0x30 -- Sprite 0x2c
    "11110000", --  353 - 0x161  :  240 - 0xf0
    "11110000", --  354 - 0x162  :  240 - 0xf0
    "11110001", --  355 - 0x163  :  241 - 0xf1
    "11110110", --  356 - 0x164  :  246 - 0xf6
    "11000110", --  357 - 0x165  :  198 - 0xc6
    "10000100", --  358 - 0x166  :  132 - 0x84
    "00000000", --  359 - 0x167  :    0 - 0x0
    "00000000", --  360 - 0x168  :    0 - 0x0 -- Sprite 0x2d
    "00000000", --  361 - 0x169  :    0 - 0x0
    "00000000", --  362 - 0x16a  :    0 - 0x0
    "00000000", --  363 - 0x16b  :    0 - 0x0
    "00000000", --  364 - 0x16c  :    0 - 0x0
    "00000000", --  365 - 0x16d  :    0 - 0x0
    "00000000", --  366 - 0x16e  :    0 - 0x0
    "00000000", --  367 - 0x16f  :    0 - 0x0
    "00011111", --  368 - 0x170  :   31 - 0x1f -- Sprite 0x2e
    "00011111", --  369 - 0x171  :   31 - 0x1f
    "00111111", --  370 - 0x172  :   63 - 0x3f
    "00111110", --  371 - 0x173  :   62 - 0x3e
    "01111100", --  372 - 0x174  :  124 - 0x7c
    "01111000", --  373 - 0x175  :  120 - 0x78
    "11110000", --  374 - 0x176  :  240 - 0xf0
    "11100000", --  375 - 0x177  :  224 - 0xe0
    "10110000", --  376 - 0x178  :  176 - 0xb0 -- Sprite 0x2f
    "10010000", --  377 - 0x179  :  144 - 0x90
    "00011000", --  378 - 0x17a  :   24 - 0x18
    "00001000", --  379 - 0x17b  :    8 - 0x8
    "01000000", --  380 - 0x17c  :   64 - 0x40
    "00000000", --  381 - 0x17d  :    0 - 0x0
    "00000000", --  382 - 0x17e  :    0 - 0x0
    "00000000", --  383 - 0x17f  :    0 - 0x0
    "11000000", --  384 - 0x180  :  192 - 0xc0 -- Sprite 0x30
    "11100000", --  385 - 0x181  :  224 - 0xe0
    "11111100", --  386 - 0x182  :  252 - 0xfc
    "11111110", --  387 - 0x183  :  254 - 0xfe
    "11111111", --  388 - 0x184  :  255 - 0xff
    "01111111", --  389 - 0x185  :  127 - 0x7f
    "00000011", --  390 - 0x186  :    3 - 0x3
    "00000000", --  391 - 0x187  :    0 - 0x0
    "00000000", --  392 - 0x188  :    0 - 0x0 -- Sprite 0x31
    "00000000", --  393 - 0x189  :    0 - 0x0
    "00010000", --  394 - 0x18a  :   16 - 0x10
    "00111000", --  395 - 0x18b  :   56 - 0x38
    "00111110", --  396 - 0x18c  :   62 - 0x3e
    "00111100", --  397 - 0x18d  :   60 - 0x3c
    "00111000", --  398 - 0x18e  :   56 - 0x38
    "00011000", --  399 - 0x18f  :   24 - 0x18
    "00000000", --  400 - 0x190  :    0 - 0x0 -- Sprite 0x32
    "00000000", --  401 - 0x191  :    0 - 0x0
    "00000000", --  402 - 0x192  :    0 - 0x0
    "00000111", --  403 - 0x193  :    7 - 0x7
    "00001111", --  404 - 0x194  :   15 - 0xf
    "00001111", --  405 - 0x195  :   15 - 0xf
    "00001111", --  406 - 0x196  :   15 - 0xf
    "00000011", --  407 - 0x197  :    3 - 0x3
    "00000000", --  408 - 0x198  :    0 - 0x0 -- Sprite 0x33
    "00000000", --  409 - 0x199  :    0 - 0x0
    "00000000", --  410 - 0x19a  :    0 - 0x0
    "11110000", --  411 - 0x19b  :  240 - 0xf0
    "11111100", --  412 - 0x19c  :  252 - 0xfc
    "11111110", --  413 - 0x19d  :  254 - 0xfe
    "11111100", --  414 - 0x19e  :  252 - 0xfc
    "11111000", --  415 - 0x19f  :  248 - 0xf8
    "00000111", --  416 - 0x1a0  :    7 - 0x7 -- Sprite 0x34
    "00001111", --  417 - 0x1a1  :   15 - 0xf
    "00011011", --  418 - 0x1a2  :   27 - 0x1b
    "00011000", --  419 - 0x1a3  :   24 - 0x18
    "00010000", --  420 - 0x1a4  :   16 - 0x10
    "00110000", --  421 - 0x1a5  :   48 - 0x30
    "00100001", --  422 - 0x1a6  :   33 - 0x21
    "00000001", --  423 - 0x1a7  :    1 - 0x1
    "10101000", --  424 - 0x1a8  :  168 - 0xa8 -- Sprite 0x35
    "11111100", --  425 - 0x1a9  :  252 - 0xfc
    "11111000", --  426 - 0x1aa  :  248 - 0xf8
    "00000000", --  427 - 0x1ab  :    0 - 0x0
    "00000000", --  428 - 0x1ac  :    0 - 0x0
    "00000000", --  429 - 0x1ad  :    0 - 0x0
    "11000000", --  430 - 0x1ae  :  192 - 0xc0
    "11100000", --  431 - 0x1af  :  224 - 0xe0
    "00000000", --  432 - 0x1b0  :    0 - 0x0 -- Sprite 0x36
    "00000000", --  433 - 0x1b1  :    0 - 0x0
    "00001111", --  434 - 0x1b2  :   15 - 0xf
    "00011111", --  435 - 0x1b3  :   31 - 0x1f
    "00011111", --  436 - 0x1b4  :   31 - 0x1f
    "00011111", --  437 - 0x1b5  :   31 - 0x1f
    "00000111", --  438 - 0x1b6  :    7 - 0x7
    "00111100", --  439 - 0x1b7  :   60 - 0x3c
    "00000000", --  440 - 0x1b8  :    0 - 0x0 -- Sprite 0x37
    "00000000", --  441 - 0x1b9  :    0 - 0x0
    "11100000", --  442 - 0x1ba  :  224 - 0xe0
    "11111000", --  443 - 0x1bb  :  248 - 0xf8
    "11111100", --  444 - 0x1bc  :  252 - 0xfc
    "11111000", --  445 - 0x1bd  :  248 - 0xf8
    "11110000", --  446 - 0x1be  :  240 - 0xf0
    "11000000", --  447 - 0x1bf  :  192 - 0xc0
    "11111100", --  448 - 0x1c0  :  252 - 0xfc -- Sprite 0x38
    "11101101", --  449 - 0x1c1  :  237 - 0xed
    "11000000", --  450 - 0x1c2  :  192 - 0xc0
    "00000000", --  451 - 0x1c3  :    0 - 0x0
    "00000000", --  452 - 0x1c4  :    0 - 0x0
    "01100000", --  453 - 0x1c5  :   96 - 0x60
    "01110000", --  454 - 0x1c6  :  112 - 0x70
    "00111000", --  455 - 0x1c7  :   56 - 0x38
    "01111110", --  456 - 0x1c8  :  126 - 0x7e -- Sprite 0x39
    "00011110", --  457 - 0x1c9  :   30 - 0x1e
    "00000100", --  458 - 0x1ca  :    4 - 0x4
    "00001100", --  459 - 0x1cb  :   12 - 0xc
    "00001100", --  460 - 0x1cc  :   12 - 0xc
    "00001100", --  461 - 0x1cd  :   12 - 0xc
    "00000000", --  462 - 0x1ce  :    0 - 0x0
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "00000000", --  464 - 0x1d0  :    0 - 0x0 -- Sprite 0x3a
    "00000000", --  465 - 0x1d1  :    0 - 0x0
    "00001111", --  466 - 0x1d2  :   15 - 0xf
    "00011111", --  467 - 0x1d3  :   31 - 0x1f
    "00011111", --  468 - 0x1d4  :   31 - 0x1f
    "00011111", --  469 - 0x1d5  :   31 - 0x1f
    "00000111", --  470 - 0x1d6  :    7 - 0x7
    "00001101", --  471 - 0x1d7  :   13 - 0xd
    "00011110", --  472 - 0x1d8  :   30 - 0x1e -- Sprite 0x3b
    "00011100", --  473 - 0x1d9  :   28 - 0x1c
    "00011110", --  474 - 0x1da  :   30 - 0x1e
    "00001111", --  475 - 0x1db  :   15 - 0xf
    "00000111", --  476 - 0x1dc  :    7 - 0x7
    "00000000", --  477 - 0x1dd  :    0 - 0x0
    "00000111", --  478 - 0x1de  :    7 - 0x7
    "00000111", --  479 - 0x1df  :    7 - 0x7
    "01100000", --  480 - 0x1e0  :   96 - 0x60 -- Sprite 0x3c
    "10010000", --  481 - 0x1e1  :  144 - 0x90
    "00000000", --  482 - 0x1e2  :    0 - 0x0
    "10000000", --  483 - 0x1e3  :  128 - 0x80
    "00000000", --  484 - 0x1e4  :    0 - 0x0
    "11100000", --  485 - 0x1e5  :  224 - 0xe0
    "11110000", --  486 - 0x1e6  :  240 - 0xf0
    "10000000", --  487 - 0x1e7  :  128 - 0x80
    "00000000", --  488 - 0x1e8  :    0 - 0x0 -- Sprite 0x3d
    "00010000", --  489 - 0x1e9  :   16 - 0x10
    "00111111", --  490 - 0x1ea  :   63 - 0x3f
    "01111111", --  491 - 0x1eb  :  127 - 0x7f
    "01111111", --  492 - 0x1ec  :  127 - 0x7f
    "00111111", --  493 - 0x1ed  :   63 - 0x3f
    "00000011", --  494 - 0x1ee  :    3 - 0x3
    "00001111", --  495 - 0x1ef  :   15 - 0xf
    "00000000", --  496 - 0x1f0  :    0 - 0x0 -- Sprite 0x3e
    "00000000", --  497 - 0x1f1  :    0 - 0x0
    "11100000", --  498 - 0x1f2  :  224 - 0xe0
    "11111000", --  499 - 0x1f3  :  248 - 0xf8
    "11111100", --  500 - 0x1f4  :  252 - 0xfc
    "11111000", --  501 - 0x1f5  :  248 - 0xf8
    "10110000", --  502 - 0x1f6  :  176 - 0xb0
    "00111000", --  503 - 0x1f7  :   56 - 0x38
    "00011111", --  504 - 0x1f8  :   31 - 0x1f -- Sprite 0x3f
    "00000111", --  505 - 0x1f9  :    7 - 0x7
    "00000000", --  506 - 0x1fa  :    0 - 0x0
    "00001110", --  507 - 0x1fb  :   14 - 0xe
    "00001111", --  508 - 0x1fc  :   15 - 0xf
    "01010011", --  509 - 0x1fd  :   83 - 0x53
    "01111100", --  510 - 0x1fe  :  124 - 0x7c
    "00111100", --  511 - 0x1ff  :   60 - 0x3c
    "11111000", --  512 - 0x200  :  248 - 0xf8 -- Sprite 0x40
    "11111000", --  513 - 0x201  :  248 - 0xf8
    "11110000", --  514 - 0x202  :  240 - 0xf0
    "00000000", --  515 - 0x203  :    0 - 0x0
    "00000000", --  516 - 0x204  :    0 - 0x0
    "10000000", --  517 - 0x205  :  128 - 0x80
    "00000000", --  518 - 0x206  :    0 - 0x0
    "00000000", --  519 - 0x207  :    0 - 0x0
    "00000111", --  520 - 0x208  :    7 - 0x7 -- Sprite 0x41
    "00000111", --  521 - 0x209  :    7 - 0x7
    "00000011", --  522 - 0x20a  :    3 - 0x3
    "11110111", --  523 - 0x20b  :  247 - 0xf7
    "11111111", --  524 - 0x20c  :  255 - 0xff
    "11111111", --  525 - 0x20d  :  255 - 0xff
    "11111110", --  526 - 0x20e  :  254 - 0xfe
    "11111100", --  527 - 0x20f  :  252 - 0xfc
    "00111110", --  528 - 0x210  :   62 - 0x3e -- Sprite 0x42
    "01111111", --  529 - 0x211  :  127 - 0x7f
    "11111111", --  530 - 0x212  :  255 - 0xff
    "11100010", --  531 - 0x213  :  226 - 0xe2
    "01010000", --  532 - 0x214  :   80 - 0x50
    "00111000", --  533 - 0x215  :   56 - 0x38
    "01110000", --  534 - 0x216  :  112 - 0x70
    "01000000", --  535 - 0x217  :   64 - 0x40
    "11101000", --  536 - 0x218  :  232 - 0xe8 -- Sprite 0x43
    "01110001", --  537 - 0x219  :  113 - 0x71
    "00000001", --  538 - 0x21a  :    1 - 0x1
    "01001011", --  539 - 0x21b  :   75 - 0x4b
    "00000011", --  540 - 0x21c  :    3 - 0x3
    "00000011", --  541 - 0x21d  :    3 - 0x3
    "00000000", --  542 - 0x21e  :    0 - 0x0
    "00000000", --  543 - 0x21f  :    0 - 0x0
    "00000101", --  544 - 0x220  :    5 - 0x5 -- Sprite 0x44
    "00000011", --  545 - 0x221  :    3 - 0x3
    "00000001", --  546 - 0x222  :    1 - 0x1
    "00110000", --  547 - 0x223  :   48 - 0x30
    "00110000", --  548 - 0x224  :   48 - 0x30
    "00110000", --  549 - 0x225  :   48 - 0x30
    "00100110", --  550 - 0x226  :   38 - 0x26
    "00000100", --  551 - 0x227  :    4 - 0x4
    "11111110", --  552 - 0x228  :  254 - 0xfe -- Sprite 0x45
    "11111100", --  553 - 0x229  :  252 - 0xfc
    "11100000", --  554 - 0x22a  :  224 - 0xe0
    "00000000", --  555 - 0x22b  :    0 - 0x0
    "00000000", --  556 - 0x22c  :    0 - 0x0
    "00000000", --  557 - 0x22d  :    0 - 0x0
    "00000000", --  558 - 0x22e  :    0 - 0x0
    "00000000", --  559 - 0x22f  :    0 - 0x0
    "00000101", --  560 - 0x230  :    5 - 0x5 -- Sprite 0x46
    "00000011", --  561 - 0x231  :    3 - 0x3
    "00000001", --  562 - 0x232  :    1 - 0x1
    "00010000", --  563 - 0x233  :   16 - 0x10
    "00110000", --  564 - 0x234  :   48 - 0x30
    "00001100", --  565 - 0x235  :   12 - 0xc
    "00011100", --  566 - 0x236  :   28 - 0x1c
    "00011000", --  567 - 0x237  :   24 - 0x18
    "11000000", --  568 - 0x238  :  192 - 0xc0 -- Sprite 0x47
    "11100000", --  569 - 0x239  :  224 - 0xe0
    "11110000", --  570 - 0x23a  :  240 - 0xf0
    "01111000", --  571 - 0x23b  :  120 - 0x78
    "00011000", --  572 - 0x23c  :   24 - 0x18
    "00001000", --  573 - 0x23d  :    8 - 0x8
    "00000000", --  574 - 0x23e  :    0 - 0x0
    "00000000", --  575 - 0x23f  :    0 - 0x0
    "00000111", --  576 - 0x240  :    7 - 0x7 -- Sprite 0x48
    "00001111", --  577 - 0x241  :   15 - 0xf
    "00111110", --  578 - 0x242  :   62 - 0x3e
    "01111100", --  579 - 0x243  :  124 - 0x7c
    "00110000", --  580 - 0x244  :   48 - 0x30
    "00001100", --  581 - 0x245  :   12 - 0xc
    "00011100", --  582 - 0x246  :   28 - 0x1c
    "00011000", --  583 - 0x247  :   24 - 0x18
    "01100000", --  584 - 0x248  :   96 - 0x60 -- Sprite 0x49
    "01100000", --  585 - 0x249  :   96 - 0x60
    "01100000", --  586 - 0x24a  :   96 - 0x60
    "10000000", --  587 - 0x24b  :  128 - 0x80
    "00000000", --  588 - 0x24c  :    0 - 0x0
    "00000000", --  589 - 0x24d  :    0 - 0x0
    "00000000", --  590 - 0x24e  :    0 - 0x0
    "00000000", --  591 - 0x24f  :    0 - 0x0
    "01110011", --  592 - 0x250  :  115 - 0x73 -- Sprite 0x4a
    "11110011", --  593 - 0x251  :  243 - 0xf3
    "11110000", --  594 - 0x252  :  240 - 0xf0
    "11110100", --  595 - 0x253  :  244 - 0xf4
    "11110000", --  596 - 0x254  :  240 - 0xf0
    "11110000", --  597 - 0x255  :  240 - 0xf0
    "01110000", --  598 - 0x256  :  112 - 0x70
    "01100000", --  599 - 0x257  :   96 - 0x60
    "00000000", --  600 - 0x258  :    0 - 0x0 -- Sprite 0x4b
    "00000000", --  601 - 0x259  :    0 - 0x0
    "00000000", --  602 - 0x25a  :    0 - 0x0
    "00000000", --  603 - 0x25b  :    0 - 0x0
    "00111100", --  604 - 0x25c  :   60 - 0x3c
    "00111100", --  605 - 0x25d  :   60 - 0x3c
    "11111100", --  606 - 0x25e  :  252 - 0xfc
    "11111100", --  607 - 0x25f  :  252 - 0xfc
    "01111111", --  608 - 0x260  :  127 - 0x7f -- Sprite 0x4c
    "01111111", --  609 - 0x261  :  127 - 0x7f
    "00011111", --  610 - 0x262  :   31 - 0x1f
    "00000111", --  611 - 0x263  :    7 - 0x7
    "00001011", --  612 - 0x264  :   11 - 0xb
    "00011011", --  613 - 0x265  :   27 - 0x1b
    "00111011", --  614 - 0x266  :   59 - 0x3b
    "01111011", --  615 - 0x267  :  123 - 0x7b
    "11111100", --  616 - 0x268  :  252 - 0xfc -- Sprite 0x4d
    "11111100", --  617 - 0x269  :  252 - 0xfc
    "11111000", --  618 - 0x26a  :  248 - 0xf8
    "11100000", --  619 - 0x26b  :  224 - 0xe0
    "11010000", --  620 - 0x26c  :  208 - 0xd0
    "11011000", --  621 - 0x26d  :  216 - 0xd8
    "11011100", --  622 - 0x26e  :  220 - 0xdc
    "11011110", --  623 - 0x26f  :  222 - 0xde
    "11000100", --  624 - 0x270  :  196 - 0xc4 -- Sprite 0x4e
    "11100000", --  625 - 0x271  :  224 - 0xe0
    "11100000", --  626 - 0x272  :  224 - 0xe0
    "01000000", --  627 - 0x273  :   64 - 0x40
    "00000000", --  628 - 0x274  :    0 - 0x0
    "00111100", --  629 - 0x275  :   60 - 0x3c
    "00111100", --  630 - 0x276  :   60 - 0x3c
    "01111100", --  631 - 0x277  :  124 - 0x7c
    "00011101", --  632 - 0x278  :   29 - 0x1d -- Sprite 0x4f
    "00111100", --  633 - 0x279  :   60 - 0x3c
    "00111010", --  634 - 0x27a  :   58 - 0x3a
    "00111000", --  635 - 0x27b  :   56 - 0x38
    "00110000", --  636 - 0x27c  :   48 - 0x30
    "00000000", --  637 - 0x27d  :    0 - 0x0
    "00011100", --  638 - 0x27e  :   28 - 0x1c
    "00111100", --  639 - 0x27f  :   60 - 0x3c
    "00100010", --  640 - 0x280  :   34 - 0x22 -- Sprite 0x50
    "01010101", --  641 - 0x281  :   85 - 0x55
    "01010101", --  642 - 0x282  :   85 - 0x55
    "01010101", --  643 - 0x283  :   85 - 0x55
    "01010101", --  644 - 0x284  :   85 - 0x55
    "01010101", --  645 - 0x285  :   85 - 0x55
    "01110111", --  646 - 0x286  :  119 - 0x77
    "00100010", --  647 - 0x287  :   34 - 0x22
    "00000000", --  648 - 0x288  :    0 - 0x0 -- Sprite 0x51
    "00000000", --  649 - 0x289  :    0 - 0x0
    "00000000", --  650 - 0x28a  :    0 - 0x0
    "00000000", --  651 - 0x28b  :    0 - 0x0
    "00000000", --  652 - 0x28c  :    0 - 0x0
    "00000000", --  653 - 0x28d  :    0 - 0x0
    "00000000", --  654 - 0x28e  :    0 - 0x0
    "00000000", --  655 - 0x28f  :    0 - 0x0
    "00000000", --  656 - 0x290  :    0 - 0x0 -- Sprite 0x52
    "00000000", --  657 - 0x291  :    0 - 0x0
    "11001111", --  658 - 0x292  :  207 - 0xcf
    "00000111", --  659 - 0x293  :    7 - 0x7
    "01111111", --  660 - 0x294  :  127 - 0x7f
    "00000000", --  661 - 0x295  :    0 - 0x0
    "00000000", --  662 - 0x296  :    0 - 0x0
    "00000000", --  663 - 0x297  :    0 - 0x0
    "00000000", --  664 - 0x298  :    0 - 0x0 -- Sprite 0x53
    "00000000", --  665 - 0x299  :    0 - 0x0
    "00111100", --  666 - 0x29a  :   60 - 0x3c
    "11111100", --  667 - 0x29b  :  252 - 0xfc
    "11111110", --  668 - 0x29c  :  254 - 0xfe
    "11100000", --  669 - 0x29d  :  224 - 0xe0
    "00000000", --  670 - 0x29e  :    0 - 0x0
    "00000000", --  671 - 0x29f  :    0 - 0x0
    "01000000", --  672 - 0x2a0  :   64 - 0x40 -- Sprite 0x54
    "11100000", --  673 - 0x2a1  :  224 - 0xe0
    "01000000", --  674 - 0x2a2  :   64 - 0x40
    "00111111", --  675 - 0x2a3  :   63 - 0x3f
    "00111110", --  676 - 0x2a4  :   62 - 0x3e
    "00111110", --  677 - 0x2a5  :   62 - 0x3e
    "00110000", --  678 - 0x2a6  :   48 - 0x30
    "00111000", --  679 - 0x2a7  :   56 - 0x38
    "00000000", --  680 - 0x2a8  :    0 - 0x0 -- Sprite 0x55
    "00000000", --  681 - 0x2a9  :    0 - 0x0
    "00000000", --  682 - 0x2aa  :    0 - 0x0
    "11111000", --  683 - 0x2ab  :  248 - 0xf8
    "11111000", --  684 - 0x2ac  :  248 - 0xf8
    "11111000", --  685 - 0x2ad  :  248 - 0xf8
    "00011000", --  686 - 0x2ae  :   24 - 0x18
    "00111000", --  687 - 0x2af  :   56 - 0x38
    "00111100", --  688 - 0x2b0  :   60 - 0x3c -- Sprite 0x56
    "00111001", --  689 - 0x2b1  :   57 - 0x39
    "00111011", --  690 - 0x2b2  :   59 - 0x3b
    "00111111", --  691 - 0x2b3  :   63 - 0x3f
    "00000000", --  692 - 0x2b4  :    0 - 0x0
    "00000000", --  693 - 0x2b5  :    0 - 0x0
    "00000000", --  694 - 0x2b6  :    0 - 0x0
    "00000000", --  695 - 0x2b7  :    0 - 0x0
    "01111000", --  696 - 0x2b8  :  120 - 0x78 -- Sprite 0x57
    "00111000", --  697 - 0x2b9  :   56 - 0x38
    "10111000", --  698 - 0x2ba  :  184 - 0xb8
    "11111000", --  699 - 0x2bb  :  248 - 0xf8
    "00000000", --  700 - 0x2bc  :    0 - 0x0
    "00000000", --  701 - 0x2bd  :    0 - 0x0
    "00000000", --  702 - 0x2be  :    0 - 0x0
    "00000000", --  703 - 0x2bf  :    0 - 0x0
    "00111111", --  704 - 0x2c0  :   63 - 0x3f -- Sprite 0x58
    "00111111", --  705 - 0x2c1  :   63 - 0x3f
    "00001111", --  706 - 0x2c2  :   15 - 0xf
    "01110111", --  707 - 0x2c3  :  119 - 0x77
    "01110111", --  708 - 0x2c4  :  119 - 0x77
    "11110111", --  709 - 0x2c5  :  247 - 0xf7
    "11110111", --  710 - 0x2c6  :  247 - 0xf7
    "11110111", --  711 - 0x2c7  :  247 - 0xf7
    "11111111", --  712 - 0x2c8  :  255 - 0xff -- Sprite 0x59
    "11111110", --  713 - 0x2c9  :  254 - 0xfe
    "11111110", --  714 - 0x2ca  :  254 - 0xfe
    "11111110", --  715 - 0x2cb  :  254 - 0xfe
    "11111010", --  716 - 0x2cc  :  250 - 0xfa
    "11111010", --  717 - 0x2cd  :  250 - 0xfa
    "11110011", --  718 - 0x2ce  :  243 - 0xf3
    "11100111", --  719 - 0x2cf  :  231 - 0xe7
    "11110000", --  720 - 0x2d0  :  240 - 0xf0 -- Sprite 0x5a
    "11111000", --  721 - 0x2d1  :  248 - 0xf8
    "11111100", --  722 - 0x2d2  :  252 - 0xfc
    "01111100", --  723 - 0x2d3  :  124 - 0x7c
    "01111000", --  724 - 0x2d4  :  120 - 0x78
    "00111000", --  725 - 0x2d5  :   56 - 0x38
    "00111100", --  726 - 0x2d6  :   60 - 0x3c
    "11111100", --  727 - 0x2d7  :  252 - 0xfc
    "11111111", --  728 - 0x2d8  :  255 - 0xff -- Sprite 0x5b
    "00000000", --  729 - 0x2d9  :    0 - 0x0
    "11000011", --  730 - 0x2da  :  195 - 0xc3
    "10000001", --  731 - 0x2db  :  129 - 0x81
    "10000001", --  732 - 0x2dc  :  129 - 0x81
    "11000011", --  733 - 0x2dd  :  195 - 0xc3
    "11111111", --  734 - 0x2de  :  255 - 0xff
    "00000000", --  735 - 0x2df  :    0 - 0x0
    "00000000", --  736 - 0x2e0  :    0 - 0x0 -- Sprite 0x5c
    "00000000", --  737 - 0x2e1  :    0 - 0x0
    "00000000", --  738 - 0x2e2  :    0 - 0x0
    "00000000", --  739 - 0x2e3  :    0 - 0x0
    "00000000", --  740 - 0x2e4  :    0 - 0x0
    "00000000", --  741 - 0x2e5  :    0 - 0x0
    "00000000", --  742 - 0x2e6  :    0 - 0x0
    "00000000", --  743 - 0x2e7  :    0 - 0x0
    "00000000", --  744 - 0x2e8  :    0 - 0x0 -- Sprite 0x5d
    "00001011", --  745 - 0x2e9  :   11 - 0xb
    "00011111", --  746 - 0x2ea  :   31 - 0x1f
    "00011111", --  747 - 0x2eb  :   31 - 0x1f
    "00011110", --  748 - 0x2ec  :   30 - 0x1e
    "00111110", --  749 - 0x2ed  :   62 - 0x3e
    "00001100", --  750 - 0x2ee  :   12 - 0xc
    "00000100", --  751 - 0x2ef  :    4 - 0x4
    "00000000", --  752 - 0x2f0  :    0 - 0x0 -- Sprite 0x5e
    "00000000", --  753 - 0x2f1  :    0 - 0x0
    "00000000", --  754 - 0x2f2  :    0 - 0x0
    "00000000", --  755 - 0x2f3  :    0 - 0x0
    "00000000", --  756 - 0x2f4  :    0 - 0x0
    "00000000", --  757 - 0x2f5  :    0 - 0x0
    "00000000", --  758 - 0x2f6  :    0 - 0x0
    "00000000", --  759 - 0x2f7  :    0 - 0x0
    "00000011", --  760 - 0x2f8  :    3 - 0x3 -- Sprite 0x5f
    "00001111", --  761 - 0x2f9  :   15 - 0xf
    "00001111", --  762 - 0x2fa  :   15 - 0xf
    "00001111", --  763 - 0x2fb  :   15 - 0xf
    "00001111", --  764 - 0x2fc  :   15 - 0xf
    "00000000", --  765 - 0x2fd  :    0 - 0x0
    "00000000", --  766 - 0x2fe  :    0 - 0x0
    "00000000", --  767 - 0x2ff  :    0 - 0x0
    "00000000", --  768 - 0x300  :    0 - 0x0 -- Sprite 0x60
    "00011000", --  769 - 0x301  :   24 - 0x18
    "00111100", --  770 - 0x302  :   60 - 0x3c
    "01111110", --  771 - 0x303  :  126 - 0x7e
    "01110110", --  772 - 0x304  :  118 - 0x76
    "11111011", --  773 - 0x305  :  251 - 0xfb
    "11111011", --  774 - 0x306  :  251 - 0xfb
    "11111011", --  775 - 0x307  :  251 - 0xfb
    "00000000", --  776 - 0x308  :    0 - 0x0 -- Sprite 0x61
    "00010000", --  777 - 0x309  :   16 - 0x10
    "00010000", --  778 - 0x30a  :   16 - 0x10
    "00100000", --  779 - 0x30b  :   32 - 0x20
    "00100000", --  780 - 0x30c  :   32 - 0x20
    "00100000", --  781 - 0x30d  :   32 - 0x20
    "00100000", --  782 - 0x30e  :   32 - 0x20
    "00100000", --  783 - 0x30f  :   32 - 0x20
    "00000000", --  784 - 0x310  :    0 - 0x0 -- Sprite 0x62
    "00001000", --  785 - 0x311  :    8 - 0x8
    "00001000", --  786 - 0x312  :    8 - 0x8
    "00001000", --  787 - 0x313  :    8 - 0x8
    "00001000", --  788 - 0x314  :    8 - 0x8
    "00001000", --  789 - 0x315  :    8 - 0x8
    "00001000", --  790 - 0x316  :    8 - 0x8
    "00001000", --  791 - 0x317  :    8 - 0x8
    "00000000", --  792 - 0x318  :    0 - 0x0 -- Sprite 0x63
    "00010000", --  793 - 0x319  :   16 - 0x10
    "00010000", --  794 - 0x31a  :   16 - 0x10
    "00111000", --  795 - 0x31b  :   56 - 0x38
    "00111000", --  796 - 0x31c  :   56 - 0x38
    "00111000", --  797 - 0x31d  :   56 - 0x38
    "00111000", --  798 - 0x31e  :   56 - 0x38
    "00111000", --  799 - 0x31f  :   56 - 0x38
    "00000000", --  800 - 0x320  :    0 - 0x0 -- Sprite 0x64
    "00011000", --  801 - 0x321  :   24 - 0x18
    "00111100", --  802 - 0x322  :   60 - 0x3c
    "00001110", --  803 - 0x323  :   14 - 0xe
    "00001110", --  804 - 0x324  :   14 - 0xe
    "00000100", --  805 - 0x325  :    4 - 0x4
    "00000000", --  806 - 0x326  :    0 - 0x0
    "00000000", --  807 - 0x327  :    0 - 0x0
    "00000000", --  808 - 0x328  :    0 - 0x0 -- Sprite 0x65
    "00000000", --  809 - 0x329  :    0 - 0x0
    "00000100", --  810 - 0x32a  :    4 - 0x4
    "00000110", --  811 - 0x32b  :    6 - 0x6
    "00011110", --  812 - 0x32c  :   30 - 0x1e
    "00111100", --  813 - 0x32d  :   60 - 0x3c
    "00011000", --  814 - 0x32e  :   24 - 0x18
    "00000000", --  815 - 0x32f  :    0 - 0x0
    "00000000", --  816 - 0x330  :    0 - 0x0 -- Sprite 0x66
    "00000000", --  817 - 0x331  :    0 - 0x0
    "00000001", --  818 - 0x332  :    1 - 0x1
    "00001010", --  819 - 0x333  :   10 - 0xa
    "00010111", --  820 - 0x334  :   23 - 0x17
    "00001111", --  821 - 0x335  :   15 - 0xf
    "00101111", --  822 - 0x336  :   47 - 0x2f
    "00011111", --  823 - 0x337  :   31 - 0x1f
    "00000000", --  824 - 0x338  :    0 - 0x0 -- Sprite 0x67
    "00000000", --  825 - 0x339  :    0 - 0x0
    "00000000", --  826 - 0x33a  :    0 - 0x0
    "00000000", --  827 - 0x33b  :    0 - 0x0
    "00000101", --  828 - 0x33c  :    5 - 0x5
    "00000111", --  829 - 0x33d  :    7 - 0x7
    "00001111", --  830 - 0x33e  :   15 - 0xf
    "00000111", --  831 - 0x33f  :    7 - 0x7
    "00000000", --  832 - 0x340  :    0 - 0x0 -- Sprite 0x68
    "00000000", --  833 - 0x341  :    0 - 0x0
    "00000000", --  834 - 0x342  :    0 - 0x0
    "00000000", --  835 - 0x343  :    0 - 0x0
    "00000000", --  836 - 0x344  :    0 - 0x0
    "00000000", --  837 - 0x345  :    0 - 0x0
    "00000001", --  838 - 0x346  :    1 - 0x1
    "00000011", --  839 - 0x347  :    3 - 0x3
    "00000000", --  840 - 0x348  :    0 - 0x0 -- Sprite 0x69
    "01100000", --  841 - 0x349  :   96 - 0x60
    "11110000", --  842 - 0x34a  :  240 - 0xf0
    "11111000", --  843 - 0x34b  :  248 - 0xf8
    "01111100", --  844 - 0x34c  :  124 - 0x7c
    "00111110", --  845 - 0x34d  :   62 - 0x3e
    "01111110", --  846 - 0x34e  :  126 - 0x7e
    "01111111", --  847 - 0x34f  :  127 - 0x7f
    "00111111", --  848 - 0x350  :   63 - 0x3f -- Sprite 0x6a
    "01011111", --  849 - 0x351  :   95 - 0x5f
    "01111111", --  850 - 0x352  :  127 - 0x7f
    "00111110", --  851 - 0x353  :   62 - 0x3e
    "00001110", --  852 - 0x354  :   14 - 0xe
    "00001010", --  853 - 0x355  :   10 - 0xa
    "01010001", --  854 - 0x356  :   81 - 0x51
    "00100000", --  855 - 0x357  :   32 - 0x20
    "00000000", --  856 - 0x358  :    0 - 0x0 -- Sprite 0x6b
    "00000000", --  857 - 0x359  :    0 - 0x0
    "00000000", --  858 - 0x35a  :    0 - 0x0
    "00000000", --  859 - 0x35b  :    0 - 0x0
    "00000000", --  860 - 0x35c  :    0 - 0x0
    "00000000", --  861 - 0x35d  :    0 - 0x0
    "00001110", --  862 - 0x35e  :   14 - 0xe
    "00011111", --  863 - 0x35f  :   31 - 0x1f
    "00111111", --  864 - 0x360  :   63 - 0x3f -- Sprite 0x6c
    "01111111", --  865 - 0x361  :  127 - 0x7f
    "01111111", --  866 - 0x362  :  127 - 0x7f
    "11111110", --  867 - 0x363  :  254 - 0xfe
    "11101100", --  868 - 0x364  :  236 - 0xec
    "11001010", --  869 - 0x365  :  202 - 0xca
    "01010001", --  870 - 0x366  :   81 - 0x51
    "00100000", --  871 - 0x367  :   32 - 0x20
    "00000000", --  872 - 0x368  :    0 - 0x0 -- Sprite 0x6d
    "01000000", --  873 - 0x369  :   64 - 0x40
    "01100011", --  874 - 0x36a  :   99 - 0x63
    "01110111", --  875 - 0x36b  :  119 - 0x77
    "01111100", --  876 - 0x36c  :  124 - 0x7c
    "00111000", --  877 - 0x36d  :   56 - 0x38
    "11111000", --  878 - 0x36e  :  248 - 0xf8
    "11100100", --  879 - 0x36f  :  228 - 0xe4
    "00000000", --  880 - 0x370  :    0 - 0x0 -- Sprite 0x6e
    "00000000", --  881 - 0x371  :    0 - 0x0
    "00000011", --  882 - 0x372  :    3 - 0x3
    "00000111", --  883 - 0x373  :    7 - 0x7
    "00001100", --  884 - 0x374  :   12 - 0xc
    "00011000", --  885 - 0x375  :   24 - 0x18
    "11111000", --  886 - 0x376  :  248 - 0xf8
    "11100100", --  887 - 0x377  :  228 - 0xe4
    "00000011", --  888 - 0x378  :    3 - 0x3 -- Sprite 0x6f
    "01000100", --  889 - 0x379  :   68 - 0x44
    "00101000", --  890 - 0x37a  :   40 - 0x28
    "00010000", --  891 - 0x37b  :   16 - 0x10
    "00001000", --  892 - 0x37c  :    8 - 0x8
    "00000100", --  893 - 0x37d  :    4 - 0x4
    "00000011", --  894 - 0x37e  :    3 - 0x3
    "00000100", --  895 - 0x37f  :    4 - 0x4
    "00000011", --  896 - 0x380  :    3 - 0x3 -- Sprite 0x70
    "00000111", --  897 - 0x381  :    7 - 0x7
    "00001111", --  898 - 0x382  :   15 - 0xf
    "00011111", --  899 - 0x383  :   31 - 0x1f
    "00100111", --  900 - 0x384  :   39 - 0x27
    "01111011", --  901 - 0x385  :  123 - 0x7b
    "01111000", --  902 - 0x386  :  120 - 0x78
    "11111011", --  903 - 0x387  :  251 - 0xfb
    "11000000", --  904 - 0x388  :  192 - 0xc0 -- Sprite 0x71
    "11100000", --  905 - 0x389  :  224 - 0xe0
    "11110000", --  906 - 0x38a  :  240 - 0xf0
    "11111000", --  907 - 0x38b  :  248 - 0xf8
    "11100100", --  908 - 0x38c  :  228 - 0xe4
    "11011110", --  909 - 0x38d  :  222 - 0xde
    "00011110", --  910 - 0x38e  :   30 - 0x1e
    "11011111", --  911 - 0x38f  :  223 - 0xdf
    "11111111", --  912 - 0x390  :  255 - 0xff -- Sprite 0x72
    "11111111", --  913 - 0x391  :  255 - 0xff
    "01111111", --  914 - 0x392  :  127 - 0x7f
    "00001111", --  915 - 0x393  :   15 - 0xf
    "00001111", --  916 - 0x394  :   15 - 0xf
    "00000111", --  917 - 0x395  :    7 - 0x7
    "00000011", --  918 - 0x396  :    3 - 0x3
    "00000000", --  919 - 0x397  :    0 - 0x0
    "11111111", --  920 - 0x398  :  255 - 0xff -- Sprite 0x73
    "11111111", --  921 - 0x399  :  255 - 0xff
    "11111110", --  922 - 0x39a  :  254 - 0xfe
    "11110000", --  923 - 0x39b  :  240 - 0xf0
    "11110000", --  924 - 0x39c  :  240 - 0xf0
    "11000000", --  925 - 0x39d  :  192 - 0xc0
    "10000000", --  926 - 0x39e  :  128 - 0x80
    "00000000", --  927 - 0x39f  :    0 - 0x0
    "00000000", --  928 - 0x3a0  :    0 - 0x0 -- Sprite 0x74
    "00000000", --  929 - 0x3a1  :    0 - 0x0
    "00011000", --  930 - 0x3a2  :   24 - 0x18
    "00100100", --  931 - 0x3a3  :   36 - 0x24
    "00100100", --  932 - 0x3a4  :   36 - 0x24
    "00011000", --  933 - 0x3a5  :   24 - 0x18
    "00000000", --  934 - 0x3a6  :    0 - 0x0
    "00000000", --  935 - 0x3a7  :    0 - 0x0
    "00111100", --  936 - 0x3a8  :   60 - 0x3c -- Sprite 0x75
    "01111110", --  937 - 0x3a9  :  126 - 0x7e
    "11111111", --  938 - 0x3aa  :  255 - 0xff
    "11111111", --  939 - 0x3ab  :  255 - 0xff
    "11111111", --  940 - 0x3ac  :  255 - 0xff
    "11111111", --  941 - 0x3ad  :  255 - 0xff
    "01111110", --  942 - 0x3ae  :  126 - 0x7e
    "00111100", --  943 - 0x3af  :   60 - 0x3c
    "00000011", --  944 - 0x3b0  :    3 - 0x3 -- Sprite 0x76
    "00000111", --  945 - 0x3b1  :    7 - 0x7
    "00001111", --  946 - 0x3b2  :   15 - 0xf
    "00011111", --  947 - 0x3b3  :   31 - 0x1f
    "00111111", --  948 - 0x3b4  :   63 - 0x3f
    "01100011", --  949 - 0x3b5  :   99 - 0x63
    "01000001", --  950 - 0x3b6  :   65 - 0x41
    "11000001", --  951 - 0x3b7  :  193 - 0xc1
    "11000000", --  952 - 0x3b8  :  192 - 0xc0 -- Sprite 0x77
    "10000000", --  953 - 0x3b9  :  128 - 0x80
    "00000000", --  954 - 0x3ba  :    0 - 0x0
    "00000000", --  955 - 0x3bb  :    0 - 0x0
    "10001100", --  956 - 0x3bc  :  140 - 0x8c
    "11111110", --  957 - 0x3bd  :  254 - 0xfe
    "11111110", --  958 - 0x3be  :  254 - 0xfe
    "11110011", --  959 - 0x3bf  :  243 - 0xf3
    "11000001", --  960 - 0x3c0  :  193 - 0xc1 -- Sprite 0x78
    "11100011", --  961 - 0x3c1  :  227 - 0xe3
    "11111111", --  962 - 0x3c2  :  255 - 0xff
    "01000111", --  963 - 0x3c3  :   71 - 0x47
    "00001111", --  964 - 0x3c4  :   15 - 0xf
    "00001111", --  965 - 0x3c5  :   15 - 0xf
    "00001111", --  966 - 0x3c6  :   15 - 0xf
    "00000111", --  967 - 0x3c7  :    7 - 0x7
    "11110001", --  968 - 0x3c8  :  241 - 0xf1 -- Sprite 0x79
    "11111001", --  969 - 0x3c9  :  249 - 0xf9
    "11111111", --  970 - 0x3ca  :  255 - 0xff
    "11100010", --  971 - 0x3cb  :  226 - 0xe2
    "11110000", --  972 - 0x3cc  :  240 - 0xf0
    "11110000", --  973 - 0x3cd  :  240 - 0xf0
    "11110000", --  974 - 0x3ce  :  240 - 0xf0
    "11100000", --  975 - 0x3cf  :  224 - 0xe0
    "00010110", --  976 - 0x3d0  :   22 - 0x16 -- Sprite 0x7a
    "00011111", --  977 - 0x3d1  :   31 - 0x1f
    "00000000", --  978 - 0x3d2  :    0 - 0x0
    "00000000", --  979 - 0x3d3  :    0 - 0x0
    "00000101", --  980 - 0x3d4  :    5 - 0x5
    "00001101", --  981 - 0x3d5  :   13 - 0xd
    "00111111", --  982 - 0x3d6  :   63 - 0x3f
    "00011111", --  983 - 0x3d7  :   31 - 0x1f
    "10000000", --  984 - 0x3d8  :  128 - 0x80 -- Sprite 0x7b
    "10000000", --  985 - 0x3d9  :  128 - 0x80
    "00000000", --  986 - 0x3da  :    0 - 0x0
    "00000000", --  987 - 0x3db  :    0 - 0x0
    "00000000", --  988 - 0x3dc  :    0 - 0x0
    "10100000", --  989 - 0x3dd  :  160 - 0xa0
    "10100000", --  990 - 0x3de  :  160 - 0xa0
    "11100000", --  991 - 0x3df  :  224 - 0xe0
    "00000000", --  992 - 0x3e0  :    0 - 0x0 -- Sprite 0x7c
    "00000100", --  993 - 0x3e1  :    4 - 0x4
    "01001110", --  994 - 0x3e2  :   78 - 0x4e
    "10001100", --  995 - 0x3e3  :  140 - 0x8c
    "00001100", --  996 - 0x3e4  :   12 - 0xc
    "01111111", --  997 - 0x3e5  :  127 - 0x7f
    "11111111", --  998 - 0x3e6  :  255 - 0xff
    "11111111", --  999 - 0x3e7  :  255 - 0xff
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0 -- Sprite 0x7d
    "00000000", -- 1001 - 0x3e9  :    0 - 0x0
    "00000000", -- 1002 - 0x3ea  :    0 - 0x0
    "00000000", -- 1003 - 0x3eb  :    0 - 0x0
    "00000000", -- 1004 - 0x3ec  :    0 - 0x0
    "00000000", -- 1005 - 0x3ed  :    0 - 0x0
    "00000001", -- 1006 - 0x3ee  :    1 - 0x1
    "00000001", -- 1007 - 0x3ef  :    1 - 0x1
    "11111111", -- 1008 - 0x3f0  :  255 - 0xff -- Sprite 0x7e
    "01111111", -- 1009 - 0x3f1  :  127 - 0x7f
    "00111111", -- 1010 - 0x3f2  :   63 - 0x3f
    "00011111", -- 1011 - 0x3f3  :   31 - 0x1f
    "00001111", -- 1012 - 0x3f4  :   15 - 0xf
    "00000111", -- 1013 - 0x3f5  :    7 - 0x7
    "00000011", -- 1014 - 0x3f6  :    3 - 0x3
    "00000001", -- 1015 - 0x3f7  :    1 - 0x1
    "11111111", -- 1016 - 0x3f8  :  255 - 0xff -- Sprite 0x7f
    "10000011", -- 1017 - 0x3f9  :  131 - 0x83
    "00101001", -- 1018 - 0x3fa  :   41 - 0x29
    "01101101", -- 1019 - 0x3fb  :  109 - 0x6d
    "01000101", -- 1020 - 0x3fc  :   69 - 0x45
    "00010001", -- 1021 - 0x3fd  :   17 - 0x11
    "00000001", -- 1022 - 0x3fe  :    1 - 0x1
    "11000111", -- 1023 - 0x3ff  :  199 - 0xc7
    "00001000", -- 1024 - 0x400  :    8 - 0x8 -- Sprite 0x80
    "00001000", -- 1025 - 0x401  :    8 - 0x8
    "00000010", -- 1026 - 0x402  :    2 - 0x2
    "00011111", -- 1027 - 0x403  :   31 - 0x1f
    "00100010", -- 1028 - 0x404  :   34 - 0x22
    "00000010", -- 1029 - 0x405  :    2 - 0x2
    "00000010", -- 1030 - 0x406  :    2 - 0x2
    "00000000", -- 1031 - 0x407  :    0 - 0x0
    "00001000", -- 1032 - 0x408  :    8 - 0x8 -- Sprite 0x81
    "00001000", -- 1033 - 0x409  :    8 - 0x8
    "00001000", -- 1034 - 0x40a  :    8 - 0x8
    "00001000", -- 1035 - 0x40b  :    8 - 0x8
    "00001000", -- 1036 - 0x40c  :    8 - 0x8
    "00001000", -- 1037 - 0x40d  :    8 - 0x8
    "00001000", -- 1038 - 0x40e  :    8 - 0x8
    "00001000", -- 1039 - 0x40f  :    8 - 0x8
    "00010000", -- 1040 - 0x410  :   16 - 0x10 -- Sprite 0x82
    "00011110", -- 1041 - 0x411  :   30 - 0x1e
    "00010000", -- 1042 - 0x412  :   16 - 0x10
    "01010000", -- 1043 - 0x413  :   80 - 0x50
    "00010000", -- 1044 - 0x414  :   16 - 0x10
    "00001000", -- 1045 - 0x415  :    8 - 0x8
    "00000000", -- 1046 - 0x416  :    0 - 0x0
    "00000000", -- 1047 - 0x417  :    0 - 0x0
    "00000000", -- 1048 - 0x418  :    0 - 0x0 -- Sprite 0x83
    "00000000", -- 1049 - 0x419  :    0 - 0x0
    "00000000", -- 1050 - 0x41a  :    0 - 0x0
    "11111110", -- 1051 - 0x41b  :  254 - 0xfe
    "00000000", -- 1052 - 0x41c  :    0 - 0x0
    "00000000", -- 1053 - 0x41d  :    0 - 0x0
    "00000000", -- 1054 - 0x41e  :    0 - 0x0
    "00000000", -- 1055 - 0x41f  :    0 - 0x0
    "00011100", -- 1056 - 0x420  :   28 - 0x1c -- Sprite 0x84
    "00101010", -- 1057 - 0x421  :   42 - 0x2a
    "01110111", -- 1058 - 0x422  :  119 - 0x77
    "11101110", -- 1059 - 0x423  :  238 - 0xee
    "11011101", -- 1060 - 0x424  :  221 - 0xdd
    "10101010", -- 1061 - 0x425  :  170 - 0xaa
    "01110100", -- 1062 - 0x426  :  116 - 0x74
    "00101000", -- 1063 - 0x427  :   40 - 0x28
    "11111111", -- 1064 - 0x428  :  255 - 0xff -- Sprite 0x85
    "11111110", -- 1065 - 0x429  :  254 - 0xfe
    "11111110", -- 1066 - 0x42a  :  254 - 0xfe
    "00000000", -- 1067 - 0x42b  :    0 - 0x0
    "11101111", -- 1068 - 0x42c  :  239 - 0xef
    "11101111", -- 1069 - 0x42d  :  239 - 0xef
    "11101111", -- 1070 - 0x42e  :  239 - 0xef
    "00000000", -- 1071 - 0x42f  :    0 - 0x0
    "11111110", -- 1072 - 0x430  :  254 - 0xfe -- Sprite 0x86
    "11111110", -- 1073 - 0x431  :  254 - 0xfe
    "11111110", -- 1074 - 0x432  :  254 - 0xfe
    "00000000", -- 1075 - 0x433  :    0 - 0x0
    "11101111", -- 1076 - 0x434  :  239 - 0xef
    "11101111", -- 1077 - 0x435  :  239 - 0xef
    "11101111", -- 1078 - 0x436  :  239 - 0xef
    "00000000", -- 1079 - 0x437  :    0 - 0x0
    "00000000", -- 1080 - 0x438  :    0 - 0x0 -- Sprite 0x87
    "01111111", -- 1081 - 0x439  :  127 - 0x7f
    "01011111", -- 1082 - 0x43a  :   95 - 0x5f
    "01111111", -- 1083 - 0x43b  :  127 - 0x7f
    "01111111", -- 1084 - 0x43c  :  127 - 0x7f
    "01111111", -- 1085 - 0x43d  :  127 - 0x7f
    "01111111", -- 1086 - 0x43e  :  127 - 0x7f
    "01111111", -- 1087 - 0x43f  :  127 - 0x7f
    "10111000", -- 1088 - 0x440  :  184 - 0xb8 -- Sprite 0x88
    "10011110", -- 1089 - 0x441  :  158 - 0x9e
    "10000000", -- 1090 - 0x442  :  128 - 0x80
    "11000000", -- 1091 - 0x443  :  192 - 0xc0
    "11100000", -- 1092 - 0x444  :  224 - 0xe0
    "11110000", -- 1093 - 0x445  :  240 - 0xf0
    "11111000", -- 1094 - 0x446  :  248 - 0xf8
    "01111100", -- 1095 - 0x447  :  124 - 0x7c
    "00000000", -- 1096 - 0x448  :    0 - 0x0 -- Sprite 0x89
    "00100011", -- 1097 - 0x449  :   35 - 0x23
    "01010111", -- 1098 - 0x44a  :   87 - 0x57
    "01001111", -- 1099 - 0x44b  :   79 - 0x4f
    "01010111", -- 1100 - 0x44c  :   87 - 0x57
    "00100111", -- 1101 - 0x44d  :   39 - 0x27
    "11000011", -- 1102 - 0x44e  :  195 - 0xc3
    "00100001", -- 1103 - 0x44f  :   33 - 0x21
    "00000000", -- 1104 - 0x450  :    0 - 0x0 -- Sprite 0x8a
    "00110000", -- 1105 - 0x451  :   48 - 0x30
    "01110000", -- 1106 - 0x452  :  112 - 0x70
    "01110000", -- 1107 - 0x453  :  112 - 0x70
    "11110000", -- 1108 - 0x454  :  240 - 0xf0
    "11100000", -- 1109 - 0x455  :  224 - 0xe0
    "11000000", -- 1110 - 0x456  :  192 - 0xc0
    "00000000", -- 1111 - 0x457  :    0 - 0x0
    "00010011", -- 1112 - 0x458  :   19 - 0x13 -- Sprite 0x8b
    "00001111", -- 1113 - 0x459  :   15 - 0xf
    "00011110", -- 1114 - 0x45a  :   30 - 0x1e
    "11110000", -- 1115 - 0x45b  :  240 - 0xf0
    "11111100", -- 1116 - 0x45c  :  252 - 0xfc
    "11111000", -- 1117 - 0x45d  :  248 - 0xf8
    "11110000", -- 1118 - 0x45e  :  240 - 0xf0
    "11100000", -- 1119 - 0x45f  :  224 - 0xe0
    "10111110", -- 1120 - 0x460  :  190 - 0xbe -- Sprite 0x8c
    "10010000", -- 1121 - 0x461  :  144 - 0x90
    "10000000", -- 1122 - 0x462  :  128 - 0x80
    "11000000", -- 1123 - 0x463  :  192 - 0xc0
    "11000000", -- 1124 - 0x464  :  192 - 0xc0
    "10000000", -- 1125 - 0x465  :  128 - 0x80
    "00000000", -- 1126 - 0x466  :    0 - 0x0
    "00000000", -- 1127 - 0x467  :    0 - 0x0
    "00000001", -- 1128 - 0x468  :    1 - 0x1 -- Sprite 0x8d
    "00000001", -- 1129 - 0x469  :    1 - 0x1
    "00000011", -- 1130 - 0x46a  :    3 - 0x3
    "00000011", -- 1131 - 0x46b  :    3 - 0x3
    "00000111", -- 1132 - 0x46c  :    7 - 0x7
    "01111111", -- 1133 - 0x46d  :  127 - 0x7f
    "01111101", -- 1134 - 0x46e  :  125 - 0x7d
    "00111101", -- 1135 - 0x46f  :   61 - 0x3d
    "00000110", -- 1136 - 0x470  :    6 - 0x6 -- Sprite 0x8e
    "00000100", -- 1137 - 0x471  :    4 - 0x4
    "00110000", -- 1138 - 0x472  :   48 - 0x30
    "00100011", -- 1139 - 0x473  :   35 - 0x23
    "00000110", -- 1140 - 0x474  :    6 - 0x6
    "01100100", -- 1141 - 0x475  :  100 - 0x64
    "01100000", -- 1142 - 0x476  :   96 - 0x60
    "00000000", -- 1143 - 0x477  :    0 - 0x0
    "00000000", -- 1144 - 0x478  :    0 - 0x0 -- Sprite 0x8f
    "01100000", -- 1145 - 0x479  :   96 - 0x60
    "01100000", -- 1146 - 0x47a  :   96 - 0x60
    "00000000", -- 1147 - 0x47b  :    0 - 0x0
    "00100000", -- 1148 - 0x47c  :   32 - 0x20
    "00110000", -- 1149 - 0x47d  :   48 - 0x30
    "00000100", -- 1150 - 0x47e  :    4 - 0x4
    "00000110", -- 1151 - 0x47f  :    6 - 0x6
    "00000000", -- 1152 - 0x480  :    0 - 0x0 -- Sprite 0x90
    "00000001", -- 1153 - 0x481  :    1 - 0x1
    "00000001", -- 1154 - 0x482  :    1 - 0x1
    "00000000", -- 1155 - 0x483  :    0 - 0x0
    "00000000", -- 1156 - 0x484  :    0 - 0x0
    "00000000", -- 1157 - 0x485  :    0 - 0x0
    "00000000", -- 1158 - 0x486  :    0 - 0x0
    "00000000", -- 1159 - 0x487  :    0 - 0x0
    "11111110", -- 1160 - 0x488  :  254 - 0xfe -- Sprite 0x91
    "11111111", -- 1161 - 0x489  :  255 - 0xff
    "11111111", -- 1162 - 0x48a  :  255 - 0xff
    "01000000", -- 1163 - 0x48b  :   64 - 0x40
    "00000001", -- 1164 - 0x48c  :    1 - 0x1
    "00000011", -- 1165 - 0x48d  :    3 - 0x3
    "00000011", -- 1166 - 0x48e  :    3 - 0x3
    "00000011", -- 1167 - 0x48f  :    3 - 0x3
    "00000001", -- 1168 - 0x490  :    1 - 0x1 -- Sprite 0x92
    "00000001", -- 1169 - 0x491  :    1 - 0x1
    "00000000", -- 1170 - 0x492  :    0 - 0x0
    "00000000", -- 1171 - 0x493  :    0 - 0x0
    "00000000", -- 1172 - 0x494  :    0 - 0x0
    "00000000", -- 1173 - 0x495  :    0 - 0x0
    "00000000", -- 1174 - 0x496  :    0 - 0x0
    "00000000", -- 1175 - 0x497  :    0 - 0x0
    "11100000", -- 1176 - 0x498  :  224 - 0xe0 -- Sprite 0x93
    "11111110", -- 1177 - 0x499  :  254 - 0xfe
    "11111111", -- 1178 - 0x49a  :  255 - 0xff
    "01111111", -- 1179 - 0x49b  :  127 - 0x7f
    "00000011", -- 1180 - 0x49c  :    3 - 0x3
    "00000010", -- 1181 - 0x49d  :    2 - 0x2
    "00000000", -- 1182 - 0x49e  :    0 - 0x0
    "00000000", -- 1183 - 0x49f  :    0 - 0x0
    "00000001", -- 1184 - 0x4a0  :    1 - 0x1 -- Sprite 0x94
    "00001101", -- 1185 - 0x4a1  :   13 - 0xd
    "00001000", -- 1186 - 0x4a2  :    8 - 0x8
    "00000000", -- 1187 - 0x4a3  :    0 - 0x0
    "00110110", -- 1188 - 0x4a4  :   54 - 0x36
    "00101100", -- 1189 - 0x4a5  :   44 - 0x2c
    "00001000", -- 1190 - 0x4a6  :    8 - 0x8
    "01100000", -- 1191 - 0x4a7  :   96 - 0x60
    "01100000", -- 1192 - 0x4a8  :   96 - 0x60 -- Sprite 0x95
    "00000000", -- 1193 - 0x4a9  :    0 - 0x0
    "00100000", -- 1194 - 0x4aa  :   32 - 0x20
    "00110000", -- 1195 - 0x4ab  :   48 - 0x30
    "00000000", -- 1196 - 0x4ac  :    0 - 0x0
    "00001000", -- 1197 - 0x4ad  :    8 - 0x8
    "00001101", -- 1198 - 0x4ae  :   13 - 0xd
    "00000001", -- 1199 - 0x4af  :    1 - 0x1
    "00000001", -- 1200 - 0x4b0  :    1 - 0x1 -- Sprite 0x96
    "00000001", -- 1201 - 0x4b1  :    1 - 0x1
    "00000011", -- 1202 - 0x4b2  :    3 - 0x3
    "01000011", -- 1203 - 0x4b3  :   67 - 0x43
    "01100111", -- 1204 - 0x4b4  :  103 - 0x67
    "01110111", -- 1205 - 0x4b5  :  119 - 0x77
    "01111011", -- 1206 - 0x4b6  :  123 - 0x7b
    "01111000", -- 1207 - 0x4b7  :  120 - 0x78
    "00000000", -- 1208 - 0x4b8  :    0 - 0x0 -- Sprite 0x97
    "00000000", -- 1209 - 0x4b9  :    0 - 0x0
    "10000000", -- 1210 - 0x4ba  :  128 - 0x80
    "10000100", -- 1211 - 0x4bb  :  132 - 0x84
    "11001100", -- 1212 - 0x4bc  :  204 - 0xcc
    "11011100", -- 1213 - 0x4bd  :  220 - 0xdc
    "10111100", -- 1214 - 0x4be  :  188 - 0xbc
    "00111100", -- 1215 - 0x4bf  :   60 - 0x3c
    "00110011", -- 1216 - 0x4c0  :   51 - 0x33 -- Sprite 0x98
    "00000111", -- 1217 - 0x4c1  :    7 - 0x7
    "00000111", -- 1218 - 0x4c2  :    7 - 0x7
    "11100011", -- 1219 - 0x4c3  :  227 - 0xe3
    "00111000", -- 1220 - 0x4c4  :   56 - 0x38
    "00111111", -- 1221 - 0x4c5  :   63 - 0x3f
    "00011100", -- 1222 - 0x4c6  :   28 - 0x1c
    "00001100", -- 1223 - 0x4c7  :   12 - 0xc
    "10011000", -- 1224 - 0x4c8  :  152 - 0x98 -- Sprite 0x99
    "11000111", -- 1225 - 0x4c9  :  199 - 0xc7
    "11001000", -- 1226 - 0x4ca  :  200 - 0xc8
    "10010010", -- 1227 - 0x4cb  :  146 - 0x92
    "00110000", -- 1228 - 0x4cc  :   48 - 0x30
    "11111000", -- 1229 - 0x4cd  :  248 - 0xf8
    "01110000", -- 1230 - 0x4ce  :  112 - 0x70
    "01100000", -- 1231 - 0x4cf  :   96 - 0x60
    "00000000", -- 1232 - 0x4d0  :    0 - 0x0 -- Sprite 0x9a
    "00000001", -- 1233 - 0x4d1  :    1 - 0x1
    "00000001", -- 1234 - 0x4d2  :    1 - 0x1
    "00000011", -- 1235 - 0x4d3  :    3 - 0x3
    "01000011", -- 1236 - 0x4d4  :   67 - 0x43
    "01100111", -- 1237 - 0x4d5  :  103 - 0x67
    "01110111", -- 1238 - 0x4d6  :  119 - 0x77
    "01111011", -- 1239 - 0x4d7  :  123 - 0x7b
    "00000000", -- 1240 - 0x4d8  :    0 - 0x0 -- Sprite 0x9b
    "00000000", -- 1241 - 0x4d9  :    0 - 0x0
    "00000000", -- 1242 - 0x4da  :    0 - 0x0
    "10000000", -- 1243 - 0x4db  :  128 - 0x80
    "10000100", -- 1244 - 0x4dc  :  132 - 0x84
    "11001100", -- 1245 - 0x4dd  :  204 - 0xcc
    "11011100", -- 1246 - 0x4de  :  220 - 0xdc
    "10111100", -- 1247 - 0x4df  :  188 - 0xbc
    "01111000", -- 1248 - 0x4e0  :  120 - 0x78 -- Sprite 0x9c
    "00110011", -- 1249 - 0x4e1  :   51 - 0x33
    "00000111", -- 1250 - 0x4e2  :    7 - 0x7
    "00000111", -- 1251 - 0x4e3  :    7 - 0x7
    "11100011", -- 1252 - 0x4e4  :  227 - 0xe3
    "00111000", -- 1253 - 0x4e5  :   56 - 0x38
    "01111111", -- 1254 - 0x4e6  :  127 - 0x7f
    "11110000", -- 1255 - 0x4e7  :  240 - 0xf0
    "00111100", -- 1256 - 0x4e8  :   60 - 0x3c -- Sprite 0x9d
    "10011000", -- 1257 - 0x4e9  :  152 - 0x98
    "11000111", -- 1258 - 0x4ea  :  199 - 0xc7
    "11001000", -- 1259 - 0x4eb  :  200 - 0xc8
    "10010010", -- 1260 - 0x4ec  :  146 - 0x92
    "00110000", -- 1261 - 0x4ed  :   48 - 0x30
    "11111000", -- 1262 - 0x4ee  :  248 - 0xf8
    "00111100", -- 1263 - 0x4ef  :   60 - 0x3c
    "00000000", -- 1264 - 0x4f0  :    0 - 0x0 -- Sprite 0x9e
    "00010000", -- 1265 - 0x4f1  :   16 - 0x10
    "01111111", -- 1266 - 0x4f2  :  127 - 0x7f
    "01111111", -- 1267 - 0x4f3  :  127 - 0x7f
    "01111111", -- 1268 - 0x4f4  :  127 - 0x7f
    "00011111", -- 1269 - 0x4f5  :   31 - 0x1f
    "00001111", -- 1270 - 0x4f6  :   15 - 0xf
    "00001111", -- 1271 - 0x4f7  :   15 - 0xf
    "00000011", -- 1272 - 0x4f8  :    3 - 0x3 -- Sprite 0x9f
    "00110011", -- 1273 - 0x4f9  :   51 - 0x33
    "00111001", -- 1274 - 0x4fa  :   57 - 0x39
    "00111010", -- 1275 - 0x4fb  :   58 - 0x3a
    "00111000", -- 1276 - 0x4fc  :   56 - 0x38
    "00011000", -- 1277 - 0x4fd  :   24 - 0x18
    "00000000", -- 1278 - 0x4fe  :    0 - 0x0
    "00000000", -- 1279 - 0x4ff  :    0 - 0x0
    "00010000", -- 1280 - 0x500  :   16 - 0x10 -- Sprite 0xa0
    "00111000", -- 1281 - 0x501  :   56 - 0x38
    "00111100", -- 1282 - 0x502  :   60 - 0x3c
    "01110100", -- 1283 - 0x503  :  116 - 0x74
    "01110110", -- 1284 - 0x504  :  118 - 0x76
    "01110110", -- 1285 - 0x505  :  118 - 0x76
    "01111110", -- 1286 - 0x506  :  126 - 0x7e
    "01111101", -- 1287 - 0x507  :  125 - 0x7d
    "00000000", -- 1288 - 0x508  :    0 - 0x0 -- Sprite 0xa1
    "00000000", -- 1289 - 0x509  :    0 - 0x0
    "00010001", -- 1290 - 0x50a  :   17 - 0x11
    "00001010", -- 1291 - 0x50b  :   10 - 0xa
    "00110100", -- 1292 - 0x50c  :   52 - 0x34
    "00101010", -- 1293 - 0x50d  :   42 - 0x2a
    "01010001", -- 1294 - 0x50e  :   81 - 0x51
    "00100000", -- 1295 - 0x50f  :   32 - 0x20
    "01111111", -- 1296 - 0x510  :  127 - 0x7f -- Sprite 0xa2
    "01100111", -- 1297 - 0x511  :  103 - 0x67
    "01100011", -- 1298 - 0x512  :   99 - 0x63
    "01110000", -- 1299 - 0x513  :  112 - 0x70
    "00111000", -- 1300 - 0x514  :   56 - 0x38
    "00111110", -- 1301 - 0x515  :   62 - 0x3e
    "01111100", -- 1302 - 0x516  :  124 - 0x7c
    "10111000", -- 1303 - 0x517  :  184 - 0xb8
    "01010001", -- 1304 - 0x518  :   81 - 0x51 -- Sprite 0xa3
    "00001010", -- 1305 - 0x519  :   10 - 0xa
    "00000100", -- 1306 - 0x51a  :    4 - 0x4
    "11101010", -- 1307 - 0x51b  :  234 - 0xea
    "01111001", -- 1308 - 0x51c  :  121 - 0x79
    "01111111", -- 1309 - 0x51d  :  127 - 0x7f
    "01110000", -- 1310 - 0x51e  :  112 - 0x70
    "00111001", -- 1311 - 0x51f  :   57 - 0x39
    "01011000", -- 1312 - 0x520  :   88 - 0x58 -- Sprite 0xa4
    "00111000", -- 1313 - 0x521  :   56 - 0x38
    "00010000", -- 1314 - 0x522  :   16 - 0x10
    "00110000", -- 1315 - 0x523  :   48 - 0x30
    "11110000", -- 1316 - 0x524  :  240 - 0xf0
    "11110000", -- 1317 - 0x525  :  240 - 0xf0
    "11100000", -- 1318 - 0x526  :  224 - 0xe0
    "11000000", -- 1319 - 0x527  :  192 - 0xc0
    "00000000", -- 1320 - 0x528  :    0 - 0x0 -- Sprite 0xa5
    "00001000", -- 1321 - 0x529  :    8 - 0x8
    "00011100", -- 1322 - 0x52a  :   28 - 0x1c
    "00111100", -- 1323 - 0x52b  :   60 - 0x3c
    "01111010", -- 1324 - 0x52c  :  122 - 0x7a
    "01111010", -- 1325 - 0x52d  :  122 - 0x7a
    "01111010", -- 1326 - 0x52e  :  122 - 0x7a
    "01111110", -- 1327 - 0x52f  :  126 - 0x7e
    "00000000", -- 1328 - 0x530  :    0 - 0x0 -- Sprite 0xa6
    "00000000", -- 1329 - 0x531  :    0 - 0x0
    "00000000", -- 1330 - 0x532  :    0 - 0x0
    "00010001", -- 1331 - 0x533  :   17 - 0x11
    "00001010", -- 1332 - 0x534  :   10 - 0xa
    "00110100", -- 1333 - 0x535  :   52 - 0x34
    "00101010", -- 1334 - 0x536  :   42 - 0x2a
    "01010001", -- 1335 - 0x537  :   81 - 0x51
    "01111111", -- 1336 - 0x538  :  127 - 0x7f -- Sprite 0xa7
    "01111101", -- 1337 - 0x539  :  125 - 0x7d
    "00111111", -- 1338 - 0x53a  :   63 - 0x3f
    "00110111", -- 1339 - 0x53b  :   55 - 0x37
    "00110011", -- 1340 - 0x53c  :   51 - 0x33
    "00111011", -- 1341 - 0x53d  :   59 - 0x3b
    "00111010", -- 1342 - 0x53e  :   58 - 0x3a
    "01111000", -- 1343 - 0x53f  :  120 - 0x78
    "00100000", -- 1344 - 0x540  :   32 - 0x20 -- Sprite 0xa8
    "01010001", -- 1345 - 0x541  :   81 - 0x51
    "00001010", -- 1346 - 0x542  :   10 - 0xa
    "00000100", -- 1347 - 0x543  :    4 - 0x4
    "11101010", -- 1348 - 0x544  :  234 - 0xea
    "00111001", -- 1349 - 0x545  :   57 - 0x39
    "01111111", -- 1350 - 0x546  :  127 - 0x7f
    "11110000", -- 1351 - 0x547  :  240 - 0xf0
    "10111100", -- 1352 - 0x548  :  188 - 0xbc -- Sprite 0xa9
    "01011000", -- 1353 - 0x549  :   88 - 0x58
    "00111000", -- 1354 - 0x54a  :   56 - 0x38
    "00010000", -- 1355 - 0x54b  :   16 - 0x10
    "00110000", -- 1356 - 0x54c  :   48 - 0x30
    "11111000", -- 1357 - 0x54d  :  248 - 0xf8
    "11111100", -- 1358 - 0x54e  :  252 - 0xfc
    "00111110", -- 1359 - 0x54f  :   62 - 0x3e
    "00000000", -- 1360 - 0x550  :    0 - 0x0 -- Sprite 0xaa
    "00000000", -- 1361 - 0x551  :    0 - 0x0
    "00000000", -- 1362 - 0x552  :    0 - 0x0
    "00000110", -- 1363 - 0x553  :    6 - 0x6
    "00001110", -- 1364 - 0x554  :   14 - 0xe
    "00001100", -- 1365 - 0x555  :   12 - 0xc
    "00000000", -- 1366 - 0x556  :    0 - 0x0
    "00000000", -- 1367 - 0x557  :    0 - 0x0
    "00000000", -- 1368 - 0x558  :    0 - 0x0 -- Sprite 0xab
    "00000000", -- 1369 - 0x559  :    0 - 0x0
    "00000000", -- 1370 - 0x55a  :    0 - 0x0
    "00000000", -- 1371 - 0x55b  :    0 - 0x0
    "00000000", -- 1372 - 0x55c  :    0 - 0x0
    "00000000", -- 1373 - 0x55d  :    0 - 0x0
    "00001111", -- 1374 - 0x55e  :   15 - 0xf
    "00011000", -- 1375 - 0x55f  :   24 - 0x18
    "00000000", -- 1376 - 0x560  :    0 - 0x0 -- Sprite 0xac
    "00000000", -- 1377 - 0x561  :    0 - 0x0
    "00000000", -- 1378 - 0x562  :    0 - 0x0
    "00000000", -- 1379 - 0x563  :    0 - 0x0
    "11111000", -- 1380 - 0x564  :  248 - 0xf8
    "00111110", -- 1381 - 0x565  :   62 - 0x3e
    "00111011", -- 1382 - 0x566  :   59 - 0x3b
    "00011000", -- 1383 - 0x567  :   24 - 0x18
    "00010000", -- 1384 - 0x568  :   16 - 0x10 -- Sprite 0xad
    "00010100", -- 1385 - 0x569  :   20 - 0x14
    "00010000", -- 1386 - 0x56a  :   16 - 0x10
    "00010000", -- 1387 - 0x56b  :   16 - 0x10
    "00111000", -- 1388 - 0x56c  :   56 - 0x38
    "01111000", -- 1389 - 0x56d  :  120 - 0x78
    "11111000", -- 1390 - 0x56e  :  248 - 0xf8
    "00110000", -- 1391 - 0x56f  :   48 - 0x30
    "00000000", -- 1392 - 0x570  :    0 - 0x0 -- Sprite 0xae
    "00000000", -- 1393 - 0x571  :    0 - 0x0
    "00000000", -- 1394 - 0x572  :    0 - 0x0
    "00000000", -- 1395 - 0x573  :    0 - 0x0
    "00000110", -- 1396 - 0x574  :    6 - 0x6
    "00001110", -- 1397 - 0x575  :   14 - 0xe
    "00001100", -- 1398 - 0x576  :   12 - 0xc
    "00000000", -- 1399 - 0x577  :    0 - 0x0
    "00000000", -- 1400 - 0x578  :    0 - 0x0 -- Sprite 0xaf
    "00000000", -- 1401 - 0x579  :    0 - 0x0
    "00000000", -- 1402 - 0x57a  :    0 - 0x0
    "00000000", -- 1403 - 0x57b  :    0 - 0x0
    "00000000", -- 1404 - 0x57c  :    0 - 0x0
    "00000000", -- 1405 - 0x57d  :    0 - 0x0
    "00000000", -- 1406 - 0x57e  :    0 - 0x0
    "00001111", -- 1407 - 0x57f  :   15 - 0xf
    "00000000", -- 1408 - 0x580  :    0 - 0x0 -- Sprite 0xb0
    "00000000", -- 1409 - 0x581  :    0 - 0x0
    "00000000", -- 1410 - 0x582  :    0 - 0x0
    "00000000", -- 1411 - 0x583  :    0 - 0x0
    "00000000", -- 1412 - 0x584  :    0 - 0x0
    "11111000", -- 1413 - 0x585  :  248 - 0xf8
    "01111110", -- 1414 - 0x586  :  126 - 0x7e
    "11110011", -- 1415 - 0x587  :  243 - 0xf3
    "00011000", -- 1416 - 0x588  :   24 - 0x18 -- Sprite 0xb1
    "00010000", -- 1417 - 0x589  :   16 - 0x10
    "00010100", -- 1418 - 0x58a  :   20 - 0x14
    "00010000", -- 1419 - 0x58b  :   16 - 0x10
    "00010000", -- 1420 - 0x58c  :   16 - 0x10
    "00111000", -- 1421 - 0x58d  :   56 - 0x38
    "01111100", -- 1422 - 0x58e  :  124 - 0x7c
    "11011110", -- 1423 - 0x58f  :  222 - 0xde
    "00000000", -- 1424 - 0x590  :    0 - 0x0 -- Sprite 0xb2
    "00001101", -- 1425 - 0x591  :   13 - 0xd
    "00011110", -- 1426 - 0x592  :   30 - 0x1e
    "00011110", -- 1427 - 0x593  :   30 - 0x1e
    "00011110", -- 1428 - 0x594  :   30 - 0x1e
    "00011111", -- 1429 - 0x595  :   31 - 0x1f
    "00001111", -- 1430 - 0x596  :   15 - 0xf
    "00000111", -- 1431 - 0x597  :    7 - 0x7
    "01111000", -- 1432 - 0x598  :  120 - 0x78 -- Sprite 0xb3
    "11110000", -- 1433 - 0x599  :  240 - 0xf0
    "00000000", -- 1434 - 0x59a  :    0 - 0x0
    "00011010", -- 1435 - 0x59b  :   26 - 0x1a
    "00111111", -- 1436 - 0x59c  :   63 - 0x3f
    "00110101", -- 1437 - 0x59d  :   53 - 0x35
    "00110101", -- 1438 - 0x59e  :   53 - 0x35
    "00111111", -- 1439 - 0x59f  :   63 - 0x3f
    "00000000", -- 1440 - 0x5a0  :    0 - 0x0 -- Sprite 0xb4
    "00000000", -- 1441 - 0x5a1  :    0 - 0x0
    "10000000", -- 1442 - 0x5a2  :  128 - 0x80
    "11100000", -- 1443 - 0x5a3  :  224 - 0xe0
    "11100000", -- 1444 - 0x5a4  :  224 - 0xe0
    "01110000", -- 1445 - 0x5a5  :  112 - 0x70
    "01110011", -- 1446 - 0x5a6  :  115 - 0x73
    "00100001", -- 1447 - 0x5a7  :   33 - 0x21
    "00011010", -- 1448 - 0x5a8  :   26 - 0x1a -- Sprite 0xb5
    "00000111", -- 1449 - 0x5a9  :    7 - 0x7
    "00001100", -- 1450 - 0x5aa  :   12 - 0xc
    "00011000", -- 1451 - 0x5ab  :   24 - 0x18
    "01111000", -- 1452 - 0x5ac  :  120 - 0x78
    "11111110", -- 1453 - 0x5ad  :  254 - 0xfe
    "11111100", -- 1454 - 0x5ae  :  252 - 0xfc
    "11110000", -- 1455 - 0x5af  :  240 - 0xf0
    "00000000", -- 1456 - 0x5b0  :    0 - 0x0 -- Sprite 0xb6
    "00000001", -- 1457 - 0x5b1  :    1 - 0x1
    "00000010", -- 1458 - 0x5b2  :    2 - 0x2
    "00000000", -- 1459 - 0x5b3  :    0 - 0x0
    "00111000", -- 1460 - 0x5b4  :   56 - 0x38
    "01111100", -- 1461 - 0x5b5  :  124 - 0x7c
    "01111110", -- 1462 - 0x5b6  :  126 - 0x7e
    "00111111", -- 1463 - 0x5b7  :   63 - 0x3f
    "00111111", -- 1464 - 0x5b8  :   63 - 0x3f -- Sprite 0xb7
    "01000000", -- 1465 - 0x5b9  :   64 - 0x40
    "01100000", -- 1466 - 0x5ba  :   96 - 0x60
    "01100000", -- 1467 - 0x5bb  :   96 - 0x60
    "00100000", -- 1468 - 0x5bc  :   32 - 0x20
    "00110000", -- 1469 - 0x5bd  :   48 - 0x30
    "00010011", -- 1470 - 0x5be  :   19 - 0x13
    "00000001", -- 1471 - 0x5bf  :    1 - 0x1
    "11000000", -- 1472 - 0x5c0  :  192 - 0xc0 -- Sprite 0xb8
    "11100000", -- 1473 - 0x5c1  :  224 - 0xe0
    "00110000", -- 1474 - 0x5c2  :   48 - 0x30
    "11010000", -- 1475 - 0x5c3  :  208 - 0xd0
    "11010000", -- 1476 - 0x5c4  :  208 - 0xd0
    "11010000", -- 1477 - 0x5c5  :  208 - 0xd0
    "11010000", -- 1478 - 0x5c6  :  208 - 0xd0
    "00000000", -- 1479 - 0x5c7  :    0 - 0x0
    "00000111", -- 1480 - 0x5c8  :    7 - 0x7 -- Sprite 0xb9
    "00001111", -- 1481 - 0x5c9  :   15 - 0xf
    "00000010", -- 1482 - 0x5ca  :    2 - 0x2
    "00011101", -- 1483 - 0x5cb  :   29 - 0x1d
    "00011111", -- 1484 - 0x5cc  :   31 - 0x1f
    "00011010", -- 1485 - 0x5cd  :   26 - 0x1a
    "00011010", -- 1486 - 0x5ce  :   26 - 0x1a
    "00000010", -- 1487 - 0x5cf  :    2 - 0x2
    "00111000", -- 1488 - 0x5d0  :   56 - 0x38 -- Sprite 0xba
    "01111100", -- 1489 - 0x5d1  :  124 - 0x7c
    "11111100", -- 1490 - 0x5d2  :  252 - 0xfc
    "11111100", -- 1491 - 0x5d3  :  252 - 0xfc
    "11111100", -- 1492 - 0x5d4  :  252 - 0xfc
    "11111110", -- 1493 - 0x5d5  :  254 - 0xfe
    "10111110", -- 1494 - 0x5d6  :  190 - 0xbe
    "10111110", -- 1495 - 0x5d7  :  190 - 0xbe
    "00011100", -- 1496 - 0x5d8  :   28 - 0x1c -- Sprite 0xbb
    "00111110", -- 1497 - 0x5d9  :   62 - 0x3e
    "00111111", -- 1498 - 0x5da  :   63 - 0x3f
    "00111111", -- 1499 - 0x5db  :   63 - 0x3f
    "00111111", -- 1500 - 0x5dc  :   63 - 0x3f
    "01111111", -- 1501 - 0x5dd  :  127 - 0x7f
    "01111101", -- 1502 - 0x5de  :  125 - 0x7d
    "01111101", -- 1503 - 0x5df  :  125 - 0x7d
    "01111101", -- 1504 - 0x5e0  :  125 - 0x7d -- Sprite 0xbc
    "01111111", -- 1505 - 0x5e1  :  127 - 0x7f
    "01011111", -- 1506 - 0x5e2  :   95 - 0x5f
    "00111011", -- 1507 - 0x5e3  :   59 - 0x3b
    "00111100", -- 1508 - 0x5e4  :   60 - 0x3c
    "00111111", -- 1509 - 0x5e5  :   63 - 0x3f
    "00011110", -- 1510 - 0x5e6  :   30 - 0x1e
    "00000000", -- 1511 - 0x5e7  :    0 - 0x0
    "00011100", -- 1512 - 0x5e8  :   28 - 0x1c -- Sprite 0xbd
    "00111110", -- 1513 - 0x5e9  :   62 - 0x3e
    "00111111", -- 1514 - 0x5ea  :   63 - 0x3f
    "00011111", -- 1515 - 0x5eb  :   31 - 0x1f
    "00111111", -- 1516 - 0x5ec  :   63 - 0x3f
    "01111111", -- 1517 - 0x5ed  :  127 - 0x7f
    "01111101", -- 1518 - 0x5ee  :  125 - 0x7d
    "01111101", -- 1519 - 0x5ef  :  125 - 0x7d
    "00000000", -- 1520 - 0x5f0  :    0 - 0x0 -- Sprite 0xbe
    "00000000", -- 1521 - 0x5f1  :    0 - 0x0
    "00000000", -- 1522 - 0x5f2  :    0 - 0x0
    "01100000", -- 1523 - 0x5f3  :   96 - 0x60
    "01100010", -- 1524 - 0x5f4  :   98 - 0x62
    "01100101", -- 1525 - 0x5f5  :  101 - 0x65
    "00111111", -- 1526 - 0x5f6  :   63 - 0x3f
    "00011111", -- 1527 - 0x5f7  :   31 - 0x1f
    "01110000", -- 1528 - 0x5f8  :  112 - 0x70 -- Sprite 0xbf
    "00111100", -- 1529 - 0x5f9  :   60 - 0x3c
    "00111100", -- 1530 - 0x5fa  :   60 - 0x3c
    "00011000", -- 1531 - 0x5fb  :   24 - 0x18
    "00000000", -- 1532 - 0x5fc  :    0 - 0x0
    "00000000", -- 1533 - 0x5fd  :    0 - 0x0
    "00000010", -- 1534 - 0x5fe  :    2 - 0x2
    "00000111", -- 1535 - 0x5ff  :    7 - 0x7
    "11001111", -- 1536 - 0x600  :  207 - 0xcf -- Sprite 0xc0
    "01111010", -- 1537 - 0x601  :  122 - 0x7a
    "01011010", -- 1538 - 0x602  :   90 - 0x5a
    "00010000", -- 1539 - 0x603  :   16 - 0x10
    "00000000", -- 1540 - 0x604  :    0 - 0x0
    "00000000", -- 1541 - 0x605  :    0 - 0x0
    "11000000", -- 1542 - 0x606  :  192 - 0xc0
    "10000000", -- 1543 - 0x607  :  128 - 0x80
    "10000101", -- 1544 - 0x608  :  133 - 0x85 -- Sprite 0xc1
    "10000100", -- 1545 - 0x609  :  132 - 0x84
    "10000110", -- 1546 - 0x60a  :  134 - 0x86
    "11000110", -- 1547 - 0x60b  :  198 - 0xc6
    "11100111", -- 1548 - 0x60c  :  231 - 0xe7
    "01110011", -- 1549 - 0x60d  :  115 - 0x73
    "01110011", -- 1550 - 0x60e  :  115 - 0x73
    "11100001", -- 1551 - 0x60f  :  225 - 0xe1
    "10000000", -- 1552 - 0x610  :  128 - 0x80 -- Sprite 0xc2
    "01001110", -- 1553 - 0x611  :   78 - 0x4e
    "01110111", -- 1554 - 0x612  :  119 - 0x77
    "11110011", -- 1555 - 0x613  :  243 - 0xf3
    "11111011", -- 1556 - 0x614  :  251 - 0xfb
    "11111001", -- 1557 - 0x615  :  249 - 0xf9
    "11111010", -- 1558 - 0x616  :  250 - 0xfa
    "01111000", -- 1559 - 0x617  :  120 - 0x78
    "00010001", -- 1560 - 0x618  :   17 - 0x11 -- Sprite 0xc3
    "00111001", -- 1561 - 0x619  :   57 - 0x39
    "01111101", -- 1562 - 0x61a  :  125 - 0x7d
    "00111001", -- 1563 - 0x61b  :   57 - 0x39
    "00000000", -- 1564 - 0x61c  :    0 - 0x0
    "00000000", -- 1565 - 0x61d  :    0 - 0x0
    "11100000", -- 1566 - 0x61e  :  224 - 0xe0
    "11100111", -- 1567 - 0x61f  :  231 - 0xe7
    "00000000", -- 1568 - 0x620  :    0 - 0x0 -- Sprite 0xc4
    "00000000", -- 1569 - 0x621  :    0 - 0x0
    "00000111", -- 1570 - 0x622  :    7 - 0x7
    "00000111", -- 1571 - 0x623  :    7 - 0x7
    "00010110", -- 1572 - 0x624  :   22 - 0x16
    "00010000", -- 1573 - 0x625  :   16 - 0x10
    "00000000", -- 1574 - 0x626  :    0 - 0x0
    "00111000", -- 1575 - 0x627  :   56 - 0x38
    "11001111", -- 1576 - 0x628  :  207 - 0xcf -- Sprite 0xc5
    "00011111", -- 1577 - 0x629  :   31 - 0x1f
    "00010111", -- 1578 - 0x62a  :   23 - 0x17
    "00010000", -- 1579 - 0x62b  :   16 - 0x10
    "00110011", -- 1580 - 0x62c  :   51 - 0x33
    "00110000", -- 1581 - 0x62d  :   48 - 0x30
    "00110000", -- 1582 - 0x62e  :   48 - 0x30
    "00100000", -- 1583 - 0x62f  :   32 - 0x20
    "00111000", -- 1584 - 0x630  :   56 - 0x38 -- Sprite 0xc6
    "00110000", -- 1585 - 0x631  :   48 - 0x30
    "01000000", -- 1586 - 0x632  :   64 - 0x40
    "11000111", -- 1587 - 0x633  :  199 - 0xc7
    "00000111", -- 1588 - 0x634  :    7 - 0x7
    "01100110", -- 1589 - 0x635  :  102 - 0x66
    "11100000", -- 1590 - 0x636  :  224 - 0xe0
    "01101100", -- 1591 - 0x637  :  108 - 0x6c
    "01100000", -- 1592 - 0x638  :   96 - 0x60 -- Sprite 0xc7
    "11000000", -- 1593 - 0x639  :  192 - 0xc0
    "10000000", -- 1594 - 0x63a  :  128 - 0x80
    "00000100", -- 1595 - 0x63b  :    4 - 0x4
    "10011110", -- 1596 - 0x63c  :  158 - 0x9e
    "11111111", -- 1597 - 0x63d  :  255 - 0xff
    "11110000", -- 1598 - 0x63e  :  240 - 0xf0
    "11111000", -- 1599 - 0x63f  :  248 - 0xf8
    "00100100", -- 1600 - 0x640  :   36 - 0x24 -- Sprite 0xc8
    "00000001", -- 1601 - 0x641  :    1 - 0x1
    "00000111", -- 1602 - 0x642  :    7 - 0x7
    "11111110", -- 1603 - 0x643  :  254 - 0xfe
    "11111111", -- 1604 - 0x644  :  255 - 0xff
    "01111111", -- 1605 - 0x645  :  127 - 0x7f
    "00111111", -- 1606 - 0x646  :   63 - 0x3f
    "01111111", -- 1607 - 0x647  :  127 - 0x7f
    "11001111", -- 1608 - 0x648  :  207 - 0xcf -- Sprite 0xc9
    "01111010", -- 1609 - 0x649  :  122 - 0x7a
    "00001010", -- 1610 - 0x64a  :   10 - 0xa
    "11111110", -- 1611 - 0x64b  :  254 - 0xfe
    "11111100", -- 1612 - 0x64c  :  252 - 0xfc
    "00000000", -- 1613 - 0x64d  :    0 - 0x0
    "00000000", -- 1614 - 0x64e  :    0 - 0x0
    "00000000", -- 1615 - 0x64f  :    0 - 0x0
    "10000101", -- 1616 - 0x650  :  133 - 0x85 -- Sprite 0xca
    "10000110", -- 1617 - 0x651  :  134 - 0x86
    "10000011", -- 1618 - 0x652  :  131 - 0x83
    "11000011", -- 1619 - 0x653  :  195 - 0xc3
    "11100001", -- 1620 - 0x654  :  225 - 0xe1
    "01110000", -- 1621 - 0x655  :  112 - 0x70
    "01110000", -- 1622 - 0x656  :  112 - 0x70
    "11100000", -- 1623 - 0x657  :  224 - 0xe0
    "01100000", -- 1624 - 0x658  :   96 - 0x60 -- Sprite 0xcb
    "11000000", -- 1625 - 0x659  :  192 - 0xc0
    "10000000", -- 1626 - 0x65a  :  128 - 0x80
    "00000000", -- 1627 - 0x65b  :    0 - 0x0
    "10011000", -- 1628 - 0x65c  :  152 - 0x98
    "11111100", -- 1629 - 0x65d  :  252 - 0xfc
    "11111110", -- 1630 - 0x65e  :  254 - 0xfe
    "11111111", -- 1631 - 0x65f  :  255 - 0xff
    "00100100", -- 1632 - 0x660  :   36 - 0x24 -- Sprite 0xcc
    "00000000", -- 1633 - 0x661  :    0 - 0x0
    "00000111", -- 1634 - 0x662  :    7 - 0x7
    "11111110", -- 1635 - 0x663  :  254 - 0xfe
    "11111111", -- 1636 - 0x664  :  255 - 0xff
    "01111111", -- 1637 - 0x665  :  127 - 0x7f
    "11111111", -- 1638 - 0x666  :  255 - 0xff
    "00000011", -- 1639 - 0x667  :    3 - 0x3
    "00000011", -- 1640 - 0x668  :    3 - 0x3 -- Sprite 0xcd
    "00001111", -- 1641 - 0x669  :   15 - 0xf
    "00100011", -- 1642 - 0x66a  :   35 - 0x23
    "01100010", -- 1643 - 0x66b  :   98 - 0x62
    "01100100", -- 1644 - 0x66c  :  100 - 0x64
    "00111100", -- 1645 - 0x66d  :   60 - 0x3c
    "00011100", -- 1646 - 0x66e  :   28 - 0x1c
    "00011110", -- 1647 - 0x66f  :   30 - 0x1e
    "00011111", -- 1648 - 0x670  :   31 - 0x1f -- Sprite 0xce
    "00111101", -- 1649 - 0x671  :   61 - 0x3d
    "01101101", -- 1650 - 0x672  :  109 - 0x6d
    "01001111", -- 1651 - 0x673  :   79 - 0x4f
    "11101110", -- 1652 - 0x674  :  238 - 0xee
    "11110011", -- 1653 - 0x675  :  243 - 0xf3
    "00100000", -- 1654 - 0x676  :   32 - 0x20
    "00000011", -- 1655 - 0x677  :    3 - 0x3
    "00000111", -- 1656 - 0x678  :    7 - 0x7 -- Sprite 0xcf
    "00000111", -- 1657 - 0x679  :    7 - 0x7
    "00011111", -- 1658 - 0x67a  :   31 - 0x1f
    "00111111", -- 1659 - 0x67b  :   63 - 0x3f
    "00001111", -- 1660 - 0x67c  :   15 - 0xf
    "01000111", -- 1661 - 0x67d  :   71 - 0x47
    "00000011", -- 1662 - 0x67e  :    3 - 0x3
    "00000000", -- 1663 - 0x67f  :    0 - 0x0
    "00000000", -- 1664 - 0x680  :    0 - 0x0 -- Sprite 0xd0
    "00000000", -- 1665 - 0x681  :    0 - 0x0
    "00000011", -- 1666 - 0x682  :    3 - 0x3
    "00000111", -- 1667 - 0x683  :    7 - 0x7
    "00001111", -- 1668 - 0x684  :   15 - 0xf
    "00001111", -- 1669 - 0x685  :   15 - 0xf
    "00011111", -- 1670 - 0x686  :   31 - 0x1f
    "00011111", -- 1671 - 0x687  :   31 - 0x1f
    "00000000", -- 1672 - 0x688  :    0 - 0x0 -- Sprite 0xd1
    "00100011", -- 1673 - 0x689  :   35 - 0x23
    "01010111", -- 1674 - 0x68a  :   87 - 0x57
    "01001111", -- 1675 - 0x68b  :   79 - 0x4f
    "01010111", -- 1676 - 0x68c  :   87 - 0x57
    "00101111", -- 1677 - 0x68d  :   47 - 0x2f
    "11011111", -- 1678 - 0x68e  :  223 - 0xdf
    "00100001", -- 1679 - 0x68f  :   33 - 0x21
    "00000000", -- 1680 - 0x690  :    0 - 0x0 -- Sprite 0xd2
    "00000000", -- 1681 - 0x691  :    0 - 0x0
    "00000000", -- 1682 - 0x692  :    0 - 0x0
    "00000000", -- 1683 - 0x693  :    0 - 0x0
    "10000000", -- 1684 - 0x694  :  128 - 0x80
    "10000000", -- 1685 - 0x695  :  128 - 0x80
    "00000000", -- 1686 - 0x696  :    0 - 0x0
    "00000000", -- 1687 - 0x697  :    0 - 0x0
    "00100011", -- 1688 - 0x698  :   35 - 0x23 -- Sprite 0xd3
    "00001111", -- 1689 - 0x699  :   15 - 0xf
    "00011110", -- 1690 - 0x69a  :   30 - 0x1e
    "11110000", -- 1691 - 0x69b  :  240 - 0xf0
    "00011100", -- 1692 - 0x69c  :   28 - 0x1c
    "00111111", -- 1693 - 0x69d  :   63 - 0x3f
    "00011111", -- 1694 - 0x69e  :   31 - 0x1f
    "00011110", -- 1695 - 0x69f  :   30 - 0x1e
    "00000000", -- 1696 - 0x6a0  :    0 - 0x0 -- Sprite 0xd4
    "10000000", -- 1697 - 0x6a1  :  128 - 0x80
    "00011000", -- 1698 - 0x6a2  :   24 - 0x18
    "00110000", -- 1699 - 0x6a3  :   48 - 0x30
    "00110100", -- 1700 - 0x6a4  :   52 - 0x34
    "11111110", -- 1701 - 0x6a5  :  254 - 0xfe
    "11111110", -- 1702 - 0x6a6  :  254 - 0xfe
    "11111110", -- 1703 - 0x6a7  :  254 - 0xfe
    "00000000", -- 1704 - 0x6a8  :    0 - 0x0 -- Sprite 0xd5
    "00000000", -- 1705 - 0x6a9  :    0 - 0x0
    "00000001", -- 1706 - 0x6aa  :    1 - 0x1
    "00000100", -- 1707 - 0x6ab  :    4 - 0x4
    "00000110", -- 1708 - 0x6ac  :    6 - 0x6
    "00000110", -- 1709 - 0x6ad  :    6 - 0x6
    "00000111", -- 1710 - 0x6ae  :    7 - 0x7
    "00000111", -- 1711 - 0x6af  :    7 - 0x7
    "00001111", -- 1712 - 0x6b0  :   15 - 0xf -- Sprite 0xd6
    "00111111", -- 1713 - 0x6b1  :   63 - 0x3f
    "01111111", -- 1714 - 0x6b2  :  127 - 0x7f
    "11111000", -- 1715 - 0x6b3  :  248 - 0xf8
    "11111000", -- 1716 - 0x6b4  :  248 - 0xf8
    "01111111", -- 1717 - 0x6b5  :  127 - 0x7f
    "00111111", -- 1718 - 0x6b6  :   63 - 0x3f
    "00001111", -- 1719 - 0x6b7  :   15 - 0xf
    "00011111", -- 1720 - 0x6b8  :   31 - 0x1f -- Sprite 0xd7
    "00011111", -- 1721 - 0x6b9  :   31 - 0x1f
    "00011111", -- 1722 - 0x6ba  :   31 - 0x1f
    "00001011", -- 1723 - 0x6bb  :   11 - 0xb
    "00000001", -- 1724 - 0x6bc  :    1 - 0x1
    "00000001", -- 1725 - 0x6bd  :    1 - 0x1
    "00000000", -- 1726 - 0x6be  :    0 - 0x0
    "00000000", -- 1727 - 0x6bf  :    0 - 0x0
    "00000011", -- 1728 - 0x6c0  :    3 - 0x3 -- Sprite 0xd8
    "00011111", -- 1729 - 0x6c1  :   31 - 0x1f
    "00111111", -- 1730 - 0x6c2  :   63 - 0x3f
    "00111111", -- 1731 - 0x6c3  :   63 - 0x3f
    "01111000", -- 1732 - 0x6c4  :  120 - 0x78
    "00000000", -- 1733 - 0x6c5  :    0 - 0x0
    "00000011", -- 1734 - 0x6c6  :    3 - 0x3
    "11111111", -- 1735 - 0x6c7  :  255 - 0xff
    "00000000", -- 1736 - 0x6c8  :    0 - 0x0 -- Sprite 0xd9
    "00000000", -- 1737 - 0x6c9  :    0 - 0x0
    "00000000", -- 1738 - 0x6ca  :    0 - 0x0
    "00000000", -- 1739 - 0x6cb  :    0 - 0x0
    "00000000", -- 1740 - 0x6cc  :    0 - 0x0
    "00000000", -- 1741 - 0x6cd  :    0 - 0x0
    "00000000", -- 1742 - 0x6ce  :    0 - 0x0
    "00000000", -- 1743 - 0x6cf  :    0 - 0x0
    "00100011", -- 1744 - 0x6d0  :   35 - 0x23 -- Sprite 0xda
    "00100111", -- 1745 - 0x6d1  :   39 - 0x27
    "00011111", -- 1746 - 0x6d2  :   31 - 0x1f
    "00000111", -- 1747 - 0x6d3  :    7 - 0x7
    "00001111", -- 1748 - 0x6d4  :   15 - 0xf
    "00011111", -- 1749 - 0x6d5  :   31 - 0x1f
    "01111111", -- 1750 - 0x6d6  :  127 - 0x7f
    "00111111", -- 1751 - 0x6d7  :   63 - 0x3f
    "11100000", -- 1752 - 0x6d8  :  224 - 0xe0 -- Sprite 0xdb
    "10000000", -- 1753 - 0x6d9  :  128 - 0x80
    "10000000", -- 1754 - 0x6da  :  128 - 0x80
    "01000000", -- 1755 - 0x6db  :   64 - 0x40
    "11100000", -- 1756 - 0x6dc  :  224 - 0xe0
    "11100000", -- 1757 - 0x6dd  :  224 - 0xe0
    "11100000", -- 1758 - 0x6de  :  224 - 0xe0
    "11000000", -- 1759 - 0x6df  :  192 - 0xc0
    "00000011", -- 1760 - 0x6e0  :    3 - 0x3 -- Sprite 0xdc
    "00000111", -- 1761 - 0x6e1  :    7 - 0x7
    "00001111", -- 1762 - 0x6e2  :   15 - 0xf
    "00011111", -- 1763 - 0x6e3  :   31 - 0x1f
    "00111111", -- 1764 - 0x6e4  :   63 - 0x3f
    "01111111", -- 1765 - 0x6e5  :  127 - 0x7f
    "11111111", -- 1766 - 0x6e6  :  255 - 0xff
    "00011111", -- 1767 - 0x6e7  :   31 - 0x1f
    "00011111", -- 1768 - 0x6e8  :   31 - 0x1f -- Sprite 0xdd
    "00010000", -- 1769 - 0x6e9  :   16 - 0x10
    "00001100", -- 1770 - 0x6ea  :   12 - 0xc
    "00010010", -- 1771 - 0x6eb  :   18 - 0x12
    "00010010", -- 1772 - 0x6ec  :   18 - 0x12
    "00101100", -- 1773 - 0x6ed  :   44 - 0x2c
    "00111111", -- 1774 - 0x6ee  :   63 - 0x3f
    "00111111", -- 1775 - 0x6ef  :   63 - 0x3f
    "00110111", -- 1776 - 0x6f0  :   55 - 0x37 -- Sprite 0xde
    "00110110", -- 1777 - 0x6f1  :   54 - 0x36
    "00110110", -- 1778 - 0x6f2  :   54 - 0x36
    "00110110", -- 1779 - 0x6f3  :   54 - 0x36
    "00010110", -- 1780 - 0x6f4  :   22 - 0x16
    "00010110", -- 1781 - 0x6f5  :   22 - 0x16
    "00010010", -- 1782 - 0x6f6  :   18 - 0x12
    "00000010", -- 1783 - 0x6f7  :    2 - 0x2
    "00010000", -- 1784 - 0x6f8  :   16 - 0x10 -- Sprite 0xdf
    "01111110", -- 1785 - 0x6f9  :  126 - 0x7e
    "11111111", -- 1786 - 0x6fa  :  255 - 0xff
    "11111111", -- 1787 - 0x6fb  :  255 - 0xff
    "11110110", -- 1788 - 0x6fc  :  246 - 0xf6
    "01110110", -- 1789 - 0x6fd  :  118 - 0x76
    "00111010", -- 1790 - 0x6fe  :   58 - 0x3a
    "00011010", -- 1791 - 0x6ff  :   26 - 0x1a
    "00000000", -- 1792 - 0x700  :    0 - 0x0 -- Sprite 0xe0
    "00000000", -- 1793 - 0x701  :    0 - 0x0
    "00111000", -- 1794 - 0x702  :   56 - 0x38
    "00000100", -- 1795 - 0x703  :    4 - 0x4
    "00000000", -- 1796 - 0x704  :    0 - 0x0
    "00000000", -- 1797 - 0x705  :    0 - 0x0
    "00000000", -- 1798 - 0x706  :    0 - 0x0
    "00000000", -- 1799 - 0x707  :    0 - 0x0
    "00000000", -- 1800 - 0x708  :    0 - 0x0 -- Sprite 0xe1
    "00000000", -- 1801 - 0x709  :    0 - 0x0
    "00000000", -- 1802 - 0x70a  :    0 - 0x0
    "00111000", -- 1803 - 0x70b  :   56 - 0x38
    "01000000", -- 1804 - 0x70c  :   64 - 0x40
    "00000000", -- 1805 - 0x70d  :    0 - 0x0
    "00000000", -- 1806 - 0x70e  :    0 - 0x0
    "00000000", -- 1807 - 0x70f  :    0 - 0x0
    "11111100", -- 1808 - 0x710  :  252 - 0xfc -- Sprite 0xe2
    "10100000", -- 1809 - 0x711  :  160 - 0xa0
    "10000000", -- 1810 - 0x712  :  128 - 0x80
    "10000000", -- 1811 - 0x713  :  128 - 0x80
    "00000000", -- 1812 - 0x714  :    0 - 0x0
    "00000000", -- 1813 - 0x715  :    0 - 0x0
    "00000000", -- 1814 - 0x716  :    0 - 0x0
    "00000000", -- 1815 - 0x717  :    0 - 0x0
    "00000111", -- 1816 - 0x718  :    7 - 0x7 -- Sprite 0xe3
    "00100111", -- 1817 - 0x719  :   39 - 0x27
    "01010111", -- 1818 - 0x71a  :   87 - 0x57
    "01001111", -- 1819 - 0x71b  :   79 - 0x4f
    "01010111", -- 1820 - 0x71c  :   87 - 0x57
    "00100111", -- 1821 - 0x71d  :   39 - 0x27
    "11000001", -- 1822 - 0x71e  :  193 - 0xc1
    "00100001", -- 1823 - 0x71f  :   33 - 0x21
    "00011101", -- 1824 - 0x720  :   29 - 0x1d -- Sprite 0xe4
    "00001111", -- 1825 - 0x721  :   15 - 0xf
    "00001111", -- 1826 - 0x722  :   15 - 0xf
    "00011111", -- 1827 - 0x723  :   31 - 0x1f
    "00011111", -- 1828 - 0x724  :   31 - 0x1f
    "00011110", -- 1829 - 0x725  :   30 - 0x1e
    "00111000", -- 1830 - 0x726  :   56 - 0x38
    "00110000", -- 1831 - 0x727  :   48 - 0x30
    "00000000", -- 1832 - 0x728  :    0 - 0x0 -- Sprite 0xe5
    "00000000", -- 1833 - 0x729  :    0 - 0x0
    "00111000", -- 1834 - 0x72a  :   56 - 0x38
    "00010000", -- 1835 - 0x72b  :   16 - 0x10
    "01001100", -- 1836 - 0x72c  :   76 - 0x4c
    "00011000", -- 1837 - 0x72d  :   24 - 0x18
    "10000110", -- 1838 - 0x72e  :  134 - 0x86
    "00100100", -- 1839 - 0x72f  :   36 - 0x24
    "00000000", -- 1840 - 0x730  :    0 - 0x0 -- Sprite 0xe6
    "01000010", -- 1841 - 0x731  :   66 - 0x42
    "00001010", -- 1842 - 0x732  :   10 - 0xa
    "01000000", -- 1843 - 0x733  :   64 - 0x40
    "00010000", -- 1844 - 0x734  :   16 - 0x10
    "00000010", -- 1845 - 0x735  :    2 - 0x2
    "00001000", -- 1846 - 0x736  :    8 - 0x8
    "00000010", -- 1847 - 0x737  :    2 - 0x2
    "00000000", -- 1848 - 0x738  :    0 - 0x0 -- Sprite 0xe7
    "00000000", -- 1849 - 0x739  :    0 - 0x0
    "10000000", -- 1850 - 0x73a  :  128 - 0x80
    "01000000", -- 1851 - 0x73b  :   64 - 0x40
    "00001000", -- 1852 - 0x73c  :    8 - 0x8
    "00001100", -- 1853 - 0x73d  :   12 - 0xc
    "00001010", -- 1854 - 0x73e  :   10 - 0xa
    "10000100", -- 1855 - 0x73f  :  132 - 0x84
    "00000000", -- 1856 - 0x740  :    0 - 0x0 -- Sprite 0xe8
    "00000000", -- 1857 - 0x741  :    0 - 0x0
    "11001111", -- 1858 - 0x742  :  207 - 0xcf
    "00100000", -- 1859 - 0x743  :   32 - 0x20
    "00100000", -- 1860 - 0x744  :   32 - 0x20
    "00100000", -- 1861 - 0x745  :   32 - 0x20
    "00100110", -- 1862 - 0x746  :   38 - 0x26
    "00101110", -- 1863 - 0x747  :   46 - 0x2e
    "11100000", -- 1864 - 0x748  :  224 - 0xe0 -- Sprite 0xe9
    "11100000", -- 1865 - 0x749  :  224 - 0xe0
    "11000000", -- 1866 - 0x74a  :  192 - 0xc0
    "00000000", -- 1867 - 0x74b  :    0 - 0x0
    "00000000", -- 1868 - 0x74c  :    0 - 0x0
    "00000000", -- 1869 - 0x74d  :    0 - 0x0
    "00000000", -- 1870 - 0x74e  :    0 - 0x0
    "00000000", -- 1871 - 0x74f  :    0 - 0x0
    "00101111", -- 1872 - 0x750  :   47 - 0x2f -- Sprite 0xea
    "00100011", -- 1873 - 0x751  :   35 - 0x23
    "00100001", -- 1874 - 0x752  :   33 - 0x21
    "00100000", -- 1875 - 0x753  :   32 - 0x20
    "00100000", -- 1876 - 0x754  :   32 - 0x20
    "00000000", -- 1877 - 0x755  :    0 - 0x0
    "00000000", -- 1878 - 0x756  :    0 - 0x0
    "00000000", -- 1879 - 0x757  :    0 - 0x0
    "11000001", -- 1880 - 0x758  :  193 - 0xc1 -- Sprite 0xeb
    "10110001", -- 1881 - 0x759  :  177 - 0xb1
    "01011001", -- 1882 - 0x75a  :   89 - 0x59
    "01101101", -- 1883 - 0x75b  :  109 - 0x6d
    "00110101", -- 1884 - 0x75c  :   53 - 0x35
    "00111011", -- 1885 - 0x75d  :   59 - 0x3b
    "00011111", -- 1886 - 0x75e  :   31 - 0x1f
    "00000011", -- 1887 - 0x75f  :    3 - 0x3
    "00000000", -- 1888 - 0x760  :    0 - 0x0 -- Sprite 0xec
    "00000010", -- 1889 - 0x761  :    2 - 0x2
    "00000000", -- 1890 - 0x762  :    0 - 0x0
    "00001000", -- 1891 - 0x763  :    8 - 0x8
    "00000010", -- 1892 - 0x764  :    2 - 0x2
    "00000000", -- 1893 - 0x765  :    0 - 0x0
    "00101000", -- 1894 - 0x766  :   40 - 0x28
    "00000000", -- 1895 - 0x767  :    0 - 0x0
    "00000100", -- 1896 - 0x768  :    4 - 0x4 -- Sprite 0xed
    "00010000", -- 1897 - 0x769  :   16 - 0x10
    "00000010", -- 1898 - 0x76a  :    2 - 0x2
    "00010000", -- 1899 - 0x76b  :   16 - 0x10
    "00000100", -- 1900 - 0x76c  :    4 - 0x4
    "00000000", -- 1901 - 0x76d  :    0 - 0x0
    "00001010", -- 1902 - 0x76e  :   10 - 0xa
    "00000000", -- 1903 - 0x76f  :    0 - 0x0
    "11000001", -- 1904 - 0x770  :  193 - 0xc1 -- Sprite 0xee
    "10110001", -- 1905 - 0x771  :  177 - 0xb1
    "01011001", -- 1906 - 0x772  :   89 - 0x59
    "01101101", -- 1907 - 0x773  :  109 - 0x6d
    "00110101", -- 1908 - 0x774  :   53 - 0x35
    "00111011", -- 1909 - 0x775  :   59 - 0x3b
    "00011111", -- 1910 - 0x776  :   31 - 0x1f
    "00000011", -- 1911 - 0x777  :    3 - 0x3
    "00000000", -- 1912 - 0x778  :    0 - 0x0 -- Sprite 0xef
    "00001111", -- 1913 - 0x779  :   15 - 0xf
    "00011111", -- 1914 - 0x77a  :   31 - 0x1f
    "11111111", -- 1915 - 0x77b  :  255 - 0xff
    "11111100", -- 1916 - 0x77c  :  252 - 0xfc
    "01100011", -- 1917 - 0x77d  :   99 - 0x63
    "00011111", -- 1918 - 0x77e  :   31 - 0x1f
    "00000011", -- 1919 - 0x77f  :    3 - 0x3
    "00000000", -- 1920 - 0x780  :    0 - 0x0 -- Sprite 0xf0
    "00000000", -- 1921 - 0x781  :    0 - 0x0
    "11111110", -- 1922 - 0x782  :  254 - 0xfe
    "11000110", -- 1923 - 0x783  :  198 - 0xc6
    "11000110", -- 1924 - 0x784  :  198 - 0xc6
    "11111110", -- 1925 - 0x785  :  254 - 0xfe
    "00000000", -- 1926 - 0x786  :    0 - 0x0
    "00000000", -- 1927 - 0x787  :    0 - 0x0
    "00000000", -- 1928 - 0x788  :    0 - 0x0 -- Sprite 0xf1
    "00000000", -- 1929 - 0x789  :    0 - 0x0
    "00000110", -- 1930 - 0x78a  :    6 - 0x6
    "00000110", -- 1931 - 0x78b  :    6 - 0x6
    "00001100", -- 1932 - 0x78c  :   12 - 0xc
    "00011000", -- 1933 - 0x78d  :   24 - 0x18
    "01110000", -- 1934 - 0x78e  :  112 - 0x70
    "01100000", -- 1935 - 0x78f  :   96 - 0x60
    "00000000", -- 1936 - 0x790  :    0 - 0x0 -- Sprite 0xf2
    "00000000", -- 1937 - 0x791  :    0 - 0x0
    "00000110", -- 1938 - 0x792  :    6 - 0x6
    "00000110", -- 1939 - 0x793  :    6 - 0x6
    "00000100", -- 1940 - 0x794  :    4 - 0x4
    "00000100", -- 1941 - 0x795  :    4 - 0x4
    "00001000", -- 1942 - 0x796  :    8 - 0x8
    "00001000", -- 1943 - 0x797  :    8 - 0x8
    "00001000", -- 1944 - 0x798  :    8 - 0x8 -- Sprite 0xf3
    "00010000", -- 1945 - 0x799  :   16 - 0x10
    "00110000", -- 1946 - 0x79a  :   48 - 0x30
    "00110000", -- 1947 - 0x79b  :   48 - 0x30
    "00110000", -- 1948 - 0x79c  :   48 - 0x30
    "00110000", -- 1949 - 0x79d  :   48 - 0x30
    "00010000", -- 1950 - 0x79e  :   16 - 0x10
    "00001000", -- 1951 - 0x79f  :    8 - 0x8
    "00000000", -- 1952 - 0x7a0  :    0 - 0x0 -- Sprite 0xf4
    "00000000", -- 1953 - 0x7a1  :    0 - 0x0
    "00000001", -- 1954 - 0x7a2  :    1 - 0x1
    "00000011", -- 1955 - 0x7a3  :    3 - 0x3
    "00000001", -- 1956 - 0x7a4  :    1 - 0x1
    "00000000", -- 1957 - 0x7a5  :    0 - 0x0
    "00000000", -- 1958 - 0x7a6  :    0 - 0x0
    "00000000", -- 1959 - 0x7a7  :    0 - 0x0
    "00000011", -- 1960 - 0x7a8  :    3 - 0x3 -- Sprite 0xf5
    "00001110", -- 1961 - 0x7a9  :   14 - 0xe
    "11111000", -- 1962 - 0x7aa  :  248 - 0xf8
    "00000000", -- 1963 - 0x7ab  :    0 - 0x0
    "00000000", -- 1964 - 0x7ac  :    0 - 0x0
    "00000000", -- 1965 - 0x7ad  :    0 - 0x0
    "00000000", -- 1966 - 0x7ae  :    0 - 0x0
    "00000000", -- 1967 - 0x7af  :    0 - 0x0
    "00100010", -- 1968 - 0x7b0  :   34 - 0x22 -- Sprite 0xf6
    "01100101", -- 1969 - 0x7b1  :  101 - 0x65
    "00100101", -- 1970 - 0x7b2  :   37 - 0x25
    "00100101", -- 1971 - 0x7b3  :   37 - 0x25
    "00100101", -- 1972 - 0x7b4  :   37 - 0x25
    "00100101", -- 1973 - 0x7b5  :   37 - 0x25
    "01110111", -- 1974 - 0x7b6  :  119 - 0x77
    "01110010", -- 1975 - 0x7b7  :  114 - 0x72
    "01100010", -- 1976 - 0x7b8  :   98 - 0x62 -- Sprite 0xf7
    "10010101", -- 1977 - 0x7b9  :  149 - 0x95
    "00010101", -- 1978 - 0x7ba  :   21 - 0x15
    "00100101", -- 1979 - 0x7bb  :   37 - 0x25
    "01000101", -- 1980 - 0x7bc  :   69 - 0x45
    "10000101", -- 1981 - 0x7bd  :  133 - 0x85
    "11110111", -- 1982 - 0x7be  :  247 - 0xf7
    "11110010", -- 1983 - 0x7bf  :  242 - 0xf2
    "10100010", -- 1984 - 0x7c0  :  162 - 0xa2 -- Sprite 0xf8
    "10100101", -- 1985 - 0x7c1  :  165 - 0xa5
    "10100101", -- 1986 - 0x7c2  :  165 - 0xa5
    "10100101", -- 1987 - 0x7c3  :  165 - 0xa5
    "11110101", -- 1988 - 0x7c4  :  245 - 0xf5
    "11110101", -- 1989 - 0x7c5  :  245 - 0xf5
    "00100111", -- 1990 - 0x7c6  :   39 - 0x27
    "00100010", -- 1991 - 0x7c7  :   34 - 0x22
    "11110010", -- 1992 - 0x7c8  :  242 - 0xf2 -- Sprite 0xf9
    "10000101", -- 1993 - 0x7c9  :  133 - 0x85
    "10000101", -- 1994 - 0x7ca  :  133 - 0x85
    "11100101", -- 1995 - 0x7cb  :  229 - 0xe5
    "00010101", -- 1996 - 0x7cc  :   21 - 0x15
    "00010101", -- 1997 - 0x7cd  :   21 - 0x15
    "11110111", -- 1998 - 0x7ce  :  247 - 0xf7
    "11100010", -- 1999 - 0x7cf  :  226 - 0xe2
    "01100010", -- 2000 - 0x7d0  :   98 - 0x62 -- Sprite 0xfa
    "10010101", -- 2001 - 0x7d1  :  149 - 0x95
    "01010101", -- 2002 - 0x7d2  :   85 - 0x55
    "01100101", -- 2003 - 0x7d3  :  101 - 0x65
    "10110101", -- 2004 - 0x7d4  :  181 - 0xb5
    "10010101", -- 2005 - 0x7d5  :  149 - 0x95
    "10010111", -- 2006 - 0x7d6  :  151 - 0x97
    "01100010", -- 2007 - 0x7d7  :   98 - 0x62
    "00100000", -- 2008 - 0x7d8  :   32 - 0x20 -- Sprite 0xfb
    "01010000", -- 2009 - 0x7d9  :   80 - 0x50
    "01010000", -- 2010 - 0x7da  :   80 - 0x50
    "01010000", -- 2011 - 0x7db  :   80 - 0x50
    "01010000", -- 2012 - 0x7dc  :   80 - 0x50
    "01010000", -- 2013 - 0x7dd  :   80 - 0x50
    "01110000", -- 2014 - 0x7de  :  112 - 0x70
    "00100000", -- 2015 - 0x7df  :   32 - 0x20
    "00000000", -- 2016 - 0x7e0  :    0 - 0x0 -- Sprite 0xfc
    "00000000", -- 2017 - 0x7e1  :    0 - 0x0
    "00000000", -- 2018 - 0x7e2  :    0 - 0x0
    "00000000", -- 2019 - 0x7e3  :    0 - 0x0
    "00000000", -- 2020 - 0x7e4  :    0 - 0x0
    "00000000", -- 2021 - 0x7e5  :    0 - 0x0
    "00000000", -- 2022 - 0x7e6  :    0 - 0x0
    "00000000", -- 2023 - 0x7e7  :    0 - 0x0
    "01100110", -- 2024 - 0x7e8  :  102 - 0x66 -- Sprite 0xfd
    "11100110", -- 2025 - 0x7e9  :  230 - 0xe6
    "01100110", -- 2026 - 0x7ea  :  102 - 0x66
    "01100110", -- 2027 - 0x7eb  :  102 - 0x66
    "01100110", -- 2028 - 0x7ec  :  102 - 0x66
    "01100111", -- 2029 - 0x7ed  :  103 - 0x67
    "11110011", -- 2030 - 0x7ee  :  243 - 0xf3
    "00000000", -- 2031 - 0x7ef  :    0 - 0x0
    "01011110", -- 2032 - 0x7f0  :   94 - 0x5e -- Sprite 0xfe
    "01011001", -- 2033 - 0x7f1  :   89 - 0x59
    "01011001", -- 2034 - 0x7f2  :   89 - 0x59
    "01011001", -- 2035 - 0x7f3  :   89 - 0x59
    "01011110", -- 2036 - 0x7f4  :   94 - 0x5e
    "11011000", -- 2037 - 0x7f5  :  216 - 0xd8
    "10011000", -- 2038 - 0x7f6  :  152 - 0x98
    "00000000", -- 2039 - 0x7f7  :    0 - 0x0
    "00000000", -- 2040 - 0x7f8  :    0 - 0x0 -- Sprite 0xff
    "00000000", -- 2041 - 0x7f9  :    0 - 0x0
    "00000000", -- 2042 - 0x7fa  :    0 - 0x0
    "00000000", -- 2043 - 0x7fb  :    0 - 0x0
    "00000000", -- 2044 - 0x7fc  :    0 - 0x0
    "00000100", -- 2045 - 0x7fd  :    4 - 0x4
    "00001000", -- 2046 - 0x7fe  :    8 - 0x8
    "00000000"  -- 2047 - 0x7ff  :    0 - 0x0
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
