//- Autcmatically generated verilog ROM from a NES memory file----
//-   PATTERN TABLE
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


//-  Original memory dump file name: donkeykong_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_PTABLE_DONKEYKONG
  (
     //input     clk,   // clock
     input      [13-1:0] addr,  //8192 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Pattern Table 0---------
      13'h0: dout  = 8'b00000000; //    0 :   0 - 0x0 -- Sprite 0x0
      13'h1: dout  = 8'b00000011; //    1 :   3 - 0x3
      13'h2: dout  = 8'b00000111; //    2 :   7 - 0x7
      13'h3: dout  = 8'b00000111; //    3 :   7 - 0x7
      13'h4: dout  = 8'b00001001; //    4 :   9 - 0x9
      13'h5: dout  = 8'b00001001; //    5 :   9 - 0x9
      13'h6: dout  = 8'b00011100; //    6 :  28 - 0x1c
      13'h7: dout  = 8'b00000000; //    7 :   0 - 0x0
      13'h8: dout  = 8'b00000000; //    8 :   0 - 0x0
      13'h9: dout  = 8'b00000011; //    9 :   3 - 0x3
      13'hA: dout  = 8'b00000111; //   10 :   7 - 0x7
      13'hB: dout  = 8'b00000000; //   11 :   0 - 0x0
      13'hC: dout  = 8'b00000110; //   12 :   6 - 0x6
      13'hD: dout  = 8'b00000110; //   13 :   6 - 0x6
      13'hE: dout  = 8'b00000011; //   14 :   3 - 0x3
      13'hF: dout  = 8'b00000011; //   15 :   3 - 0x3
      13'h10: dout  = 8'b00001111; //   16 :  15 - 0xf -- Sprite 0x1
      13'h11: dout  = 8'b00001111; //   17 :  15 - 0xf
      13'h12: dout  = 8'b00001111; //   18 :  15 - 0xf
      13'h13: dout  = 8'b11111111; //   19 : 255 - 0xff
      13'h14: dout  = 8'b11111111; //   20 : 255 - 0xff
      13'h15: dout  = 8'b11111100; //   21 : 252 - 0xfc
      13'h16: dout  = 8'b10000001; //   22 : 129 - 0x81
      13'h17: dout  = 8'b00000001; //   23 :   1 - 0x1
      13'h18: dout  = 8'b00000000; //   24 :   0 - 0x0
      13'h19: dout  = 8'b00010000; //   25 :  16 - 0x10
      13'h1A: dout  = 8'b00111100; //   26 :  60 - 0x3c
      13'h1B: dout  = 8'b00111111; //   27 :  63 - 0x3f
      13'h1C: dout  = 8'b00111111; //   28 :  63 - 0x3f
      13'h1D: dout  = 8'b00111100; //   29 :  60 - 0x3c
      13'h1E: dout  = 8'b00000000; //   30 :   0 - 0x0
      13'h1F: dout  = 8'b00000000; //   31 :   0 - 0x0
      13'h20: dout  = 8'b00000000; //   32 :   0 - 0x0 -- Sprite 0x2
      13'h21: dout  = 8'b11000000; //   33 : 192 - 0xc0
      13'h22: dout  = 8'b11111000; //   34 : 248 - 0xf8
      13'h23: dout  = 8'b10000000; //   35 : 128 - 0x80
      13'h24: dout  = 8'b00100000; //   36 :  32 - 0x20
      13'h25: dout  = 8'b10010000; //   37 : 144 - 0x90
      13'h26: dout  = 8'b00111100; //   38 :  60 - 0x3c
      13'h27: dout  = 8'b00000000; //   39 :   0 - 0x0
      13'h28: dout  = 8'b00000000; //   40 :   0 - 0x0
      13'h29: dout  = 8'b11000000; //   41 : 192 - 0xc0
      13'h2A: dout  = 8'b11111000; //   42 : 248 - 0xf8
      13'h2B: dout  = 8'b01100000; //   43 :  96 - 0x60
      13'h2C: dout  = 8'b11011100; //   44 : 220 - 0xdc
      13'h2D: dout  = 8'b01101110; //   45 : 110 - 0x6e
      13'h2E: dout  = 8'b11000000; //   46 : 192 - 0xc0
      13'h2F: dout  = 8'b11111000; //   47 : 248 - 0xf8
      13'h30: dout  = 8'b11000000; //   48 : 192 - 0xc0 -- Sprite 0x3
      13'h31: dout  = 8'b11000000; //   49 : 192 - 0xc0
      13'h32: dout  = 8'b11000000; //   50 : 192 - 0xc0
      13'h33: dout  = 8'b11110000; //   51 : 240 - 0xf0
      13'h34: dout  = 8'b11110000; //   52 : 240 - 0xf0
      13'h35: dout  = 8'b11100000; //   53 : 224 - 0xe0
      13'h36: dout  = 8'b11000000; //   54 : 192 - 0xc0
      13'h37: dout  = 8'b11100000; //   55 : 224 - 0xe0
      13'h38: dout  = 8'b01010000; //   56 :  80 - 0x50
      13'h39: dout  = 8'b00111000; //   57 :  56 - 0x38
      13'h3A: dout  = 8'b00110000; //   58 :  48 - 0x30
      13'h3B: dout  = 8'b11110000; //   59 : 240 - 0xf0
      13'h3C: dout  = 8'b11110000; //   60 : 240 - 0xf0
      13'h3D: dout  = 8'b11100000; //   61 : 224 - 0xe0
      13'h3E: dout  = 8'b00000000; //   62 :   0 - 0x0
      13'h3F: dout  = 8'b00000000; //   63 :   0 - 0x0
      13'h40: dout  = 8'b00000111; //   64 :   7 - 0x7 -- Sprite 0x4
      13'h41: dout  = 8'b00001111; //   65 :  15 - 0xf
      13'h42: dout  = 8'b00001111; //   66 :  15 - 0xf
      13'h43: dout  = 8'b00010010; //   67 :  18 - 0x12
      13'h44: dout  = 8'b00010011; //   68 :  19 - 0x13
      13'h45: dout  = 8'b00111000; //   69 :  56 - 0x38
      13'h46: dout  = 8'b00000000; //   70 :   0 - 0x0
      13'h47: dout  = 8'b00001111; //   71 :  15 - 0xf
      13'h48: dout  = 8'b00000111; //   72 :   7 - 0x7
      13'h49: dout  = 8'b00001111; //   73 :  15 - 0xf
      13'h4A: dout  = 8'b00000000; //   74 :   0 - 0x0
      13'h4B: dout  = 8'b00001101; //   75 :  13 - 0xd
      13'h4C: dout  = 8'b00001100; //   76 :  12 - 0xc
      13'h4D: dout  = 8'b00000111; //   77 :   7 - 0x7
      13'h4E: dout  = 8'b00000111; //   78 :   7 - 0x7
      13'h4F: dout  = 8'b00000000; //   79 :   0 - 0x0
      13'h50: dout  = 8'b00011111; //   80 :  31 - 0x1f -- Sprite 0x5
      13'h51: dout  = 8'b00011111; //   81 :  31 - 0x1f
      13'h52: dout  = 8'b00011111; //   82 :  31 - 0x1f
      13'h53: dout  = 8'b00011000; //   83 :  24 - 0x18
      13'h54: dout  = 8'b00011001; //   84 :  25 - 0x19
      13'h55: dout  = 8'b00011110; //   85 :  30 - 0x1e
      13'h56: dout  = 8'b00011100; //   86 :  28 - 0x1c
      13'h57: dout  = 8'b00011110; //   87 :  30 - 0x1e
      13'h58: dout  = 8'b00000001; //   88 :   1 - 0x1
      13'h59: dout  = 8'b00000011; //   89 :   3 - 0x3
      13'h5A: dout  = 8'b00000001; //   90 :   1 - 0x1
      13'h5B: dout  = 8'b00010111; //   91 :  23 - 0x17
      13'h5C: dout  = 8'b00011111; //   92 :  31 - 0x1f
      13'h5D: dout  = 8'b00011110; //   93 :  30 - 0x1e
      13'h5E: dout  = 8'b00000000; //   94 :   0 - 0x0
      13'h5F: dout  = 8'b00000000; //   95 :   0 - 0x0
      13'h60: dout  = 8'b10000000; //   96 : 128 - 0x80 -- Sprite 0x6
      13'h61: dout  = 8'b11110000; //   97 : 240 - 0xf0
      13'h62: dout  = 8'b00000000; //   98 :   0 - 0x0
      13'h63: dout  = 8'b01000000; //   99 :  64 - 0x40
      13'h64: dout  = 8'b00100000; //  100 :  32 - 0x20
      13'h65: dout  = 8'b01111000; //  101 : 120 - 0x78
      13'h66: dout  = 8'b00000000; //  102 :   0 - 0x0
      13'h67: dout  = 8'b11000000; //  103 : 192 - 0xc0
      13'h68: dout  = 8'b10000000; //  104 : 128 - 0x80
      13'h69: dout  = 8'b11110000; //  105 : 240 - 0xf0
      13'h6A: dout  = 8'b11000000; //  106 : 192 - 0xc0
      13'h6B: dout  = 8'b10111000; //  107 : 184 - 0xb8
      13'h6C: dout  = 8'b11011100; //  108 : 220 - 0xdc
      13'h6D: dout  = 8'b10000000; //  109 : 128 - 0x80
      13'h6E: dout  = 8'b11110000; //  110 : 240 - 0xf0
      13'h6F: dout  = 8'b00000000; //  111 :   0 - 0x0
      13'h70: dout  = 8'b11100000; //  112 : 224 - 0xe0 -- Sprite 0x7
      13'h71: dout  = 8'b01100000; //  113 :  96 - 0x60
      13'h72: dout  = 8'b11110000; //  114 : 240 - 0xf0
      13'h73: dout  = 8'b11110000; //  115 : 240 - 0xf0
      13'h74: dout  = 8'b11110000; //  116 : 240 - 0xf0
      13'h75: dout  = 8'b11100000; //  117 : 224 - 0xe0
      13'h76: dout  = 8'b11100000; //  118 : 224 - 0xe0
      13'h77: dout  = 8'b11110000; //  119 : 240 - 0xf0
      13'h78: dout  = 8'b10000000; //  120 : 128 - 0x80
      13'h79: dout  = 8'b11100000; //  121 : 224 - 0xe0
      13'h7A: dout  = 8'b11110000; //  122 : 240 - 0xf0
      13'h7B: dout  = 8'b11110000; //  123 : 240 - 0xf0
      13'h7C: dout  = 8'b11110000; //  124 : 240 - 0xf0
      13'h7D: dout  = 8'b11100000; //  125 : 224 - 0xe0
      13'h7E: dout  = 8'b00000000; //  126 :   0 - 0x0
      13'h7F: dout  = 8'b00000000; //  127 :   0 - 0x0
      13'h80: dout  = 8'b00000111; //  128 :   7 - 0x7 -- Sprite 0x8
      13'h81: dout  = 8'b00001111; //  129 :  15 - 0xf
      13'h82: dout  = 8'b00001111; //  130 :  15 - 0xf
      13'h83: dout  = 8'b00010010; //  131 :  18 - 0x12
      13'h84: dout  = 8'b00010011; //  132 :  19 - 0x13
      13'h85: dout  = 8'b00111000; //  133 :  56 - 0x38
      13'h86: dout  = 8'b00000000; //  134 :   0 - 0x0
      13'h87: dout  = 8'b00111111; //  135 :  63 - 0x3f
      13'h88: dout  = 8'b00000111; //  136 :   7 - 0x7
      13'h89: dout  = 8'b00001111; //  137 :  15 - 0xf
      13'h8A: dout  = 8'b00000000; //  138 :   0 - 0x0
      13'h8B: dout  = 8'b00001101; //  139 :  13 - 0xd
      13'h8C: dout  = 8'b00001100; //  140 :  12 - 0xc
      13'h8D: dout  = 8'b00000111; //  141 :   7 - 0x7
      13'h8E: dout  = 8'b00000111; //  142 :   7 - 0x7
      13'h8F: dout  = 8'b00000011; //  143 :   3 - 0x3
      13'h90: dout  = 8'b00111111; //  144 :  63 - 0x3f -- Sprite 0x9
      13'h91: dout  = 8'b00001110; //  145 :  14 - 0xe
      13'h92: dout  = 8'b00001111; //  146 :  15 - 0xf
      13'h93: dout  = 8'b00011111; //  147 :  31 - 0x1f
      13'h94: dout  = 8'b00111111; //  148 :  63 - 0x3f
      13'h95: dout  = 8'b01111100; //  149 : 124 - 0x7c
      13'h96: dout  = 8'b01110000; //  150 : 112 - 0x70
      13'h97: dout  = 8'b00111000; //  151 :  56 - 0x38
      13'h98: dout  = 8'b11000011; //  152 : 195 - 0xc3
      13'h99: dout  = 8'b11100011; //  153 : 227 - 0xe3
      13'h9A: dout  = 8'b11001111; //  154 : 207 - 0xcf
      13'h9B: dout  = 8'b00011111; //  155 :  31 - 0x1f
      13'h9C: dout  = 8'b00111111; //  156 :  63 - 0x3f
      13'h9D: dout  = 8'b00001100; //  157 :  12 - 0xc
      13'h9E: dout  = 8'b00000000; //  158 :   0 - 0x0
      13'h9F: dout  = 8'b00000000; //  159 :   0 - 0x0
      13'hA0: dout  = 8'b10000000; //  160 : 128 - 0x80 -- Sprite 0xa
      13'hA1: dout  = 8'b11110000; //  161 : 240 - 0xf0
      13'hA2: dout  = 8'b00000000; //  162 :   0 - 0x0
      13'hA3: dout  = 8'b01000000; //  163 :  64 - 0x40
      13'hA4: dout  = 8'b00100000; //  164 :  32 - 0x20
      13'hA5: dout  = 8'b01111000; //  165 : 120 - 0x78
      13'hA6: dout  = 8'b00000000; //  166 :   0 - 0x0
      13'hA7: dout  = 8'b11000000; //  167 : 192 - 0xc0
      13'hA8: dout  = 8'b10000000; //  168 : 128 - 0x80
      13'hA9: dout  = 8'b11110000; //  169 : 240 - 0xf0
      13'hAA: dout  = 8'b11000000; //  170 : 192 - 0xc0
      13'hAB: dout  = 8'b10111000; //  171 : 184 - 0xb8
      13'hAC: dout  = 8'b11011100; //  172 : 220 - 0xdc
      13'hAD: dout  = 8'b10000000; //  173 : 128 - 0x80
      13'hAE: dout  = 8'b11110000; //  174 : 240 - 0xf0
      13'hAF: dout  = 8'b00000110; //  175 :   6 - 0x6
      13'hB0: dout  = 8'b11110000; //  176 : 240 - 0xf0 -- Sprite 0xb
      13'hB1: dout  = 8'b11111000; //  177 : 248 - 0xf8
      13'hB2: dout  = 8'b11100100; //  178 : 228 - 0xe4
      13'hB3: dout  = 8'b11111100; //  179 : 252 - 0xfc
      13'hB4: dout  = 8'b11111100; //  180 : 252 - 0xfc
      13'hB5: dout  = 8'b01111100; //  181 : 124 - 0x7c
      13'hB6: dout  = 8'b00000000; //  182 :   0 - 0x0
      13'hB7: dout  = 8'b00000000; //  183 :   0 - 0x0
      13'hB8: dout  = 8'b10001110; //  184 : 142 - 0x8e
      13'hB9: dout  = 8'b11100110; //  185 : 230 - 0xe6
      13'hBA: dout  = 8'b11100000; //  186 : 224 - 0xe0
      13'hBB: dout  = 8'b11110000; //  187 : 240 - 0xf0
      13'hBC: dout  = 8'b11110000; //  188 : 240 - 0xf0
      13'hBD: dout  = 8'b01110000; //  189 : 112 - 0x70
      13'hBE: dout  = 8'b00000000; //  190 :   0 - 0x0
      13'hBF: dout  = 8'b00000000; //  191 :   0 - 0x0
      13'hC0: dout  = 8'b00000000; //  192 :   0 - 0x0 -- Sprite 0xc
      13'hC1: dout  = 8'b00000010; //  193 :   2 - 0x2
      13'hC2: dout  = 8'b00000110; //  194 :   6 - 0x6
      13'hC3: dout  = 8'b00000111; //  195 :   7 - 0x7
      13'hC4: dout  = 8'b00001001; //  196 :   9 - 0x9
      13'hC5: dout  = 8'b00001001; //  197 :   9 - 0x9
      13'hC6: dout  = 8'b00011101; //  198 :  29 - 0x1d
      13'hC7: dout  = 8'b00000011; //  199 :   3 - 0x3
      13'hC8: dout  = 8'b00000001; //  200 :   1 - 0x1
      13'hC9: dout  = 8'b00000011; //  201 :   3 - 0x3
      13'hCA: dout  = 8'b00000111; //  202 :   7 - 0x7
      13'hCB: dout  = 8'b00000000; //  203 :   0 - 0x0
      13'hCC: dout  = 8'b00000110; //  204 :   6 - 0x6
      13'hCD: dout  = 8'b00000110; //  205 :   6 - 0x6
      13'hCE: dout  = 8'b00000010; //  206 :   2 - 0x2
      13'hCF: dout  = 8'b00000000; //  207 :   0 - 0x0
      13'hD0: dout  = 8'b00001111; //  208 :  15 - 0xf -- Sprite 0xd
      13'hD1: dout  = 8'b00001111; //  209 :  15 - 0xf
      13'hD2: dout  = 8'b00001111; //  210 :  15 - 0xf
      13'hD3: dout  = 8'b11111111; //  211 : 255 - 0xff
      13'hD4: dout  = 8'b11111111; //  212 : 255 - 0xff
      13'hD5: dout  = 8'b11111100; //  213 : 252 - 0xfc
      13'hD6: dout  = 8'b10000001; //  214 : 129 - 0x81
      13'hD7: dout  = 8'b00000001; //  215 :   1 - 0x1
      13'hD8: dout  = 8'b00000000; //  216 :   0 - 0x0
      13'hD9: dout  = 8'b00000000; //  217 :   0 - 0x0
      13'hDA: dout  = 8'b00001100; //  218 :  12 - 0xc
      13'hDB: dout  = 8'b00111111; //  219 :  63 - 0x3f
      13'hDC: dout  = 8'b00111111; //  220 :  63 - 0x3f
      13'hDD: dout  = 8'b00111100; //  221 :  60 - 0x3c
      13'hDE: dout  = 8'b00000000; //  222 :   0 - 0x0
      13'hDF: dout  = 8'b00000000; //  223 :   0 - 0x0
      13'hE0: dout  = 8'b00000000; //  224 :   0 - 0x0 -- Sprite 0xe
      13'hE1: dout  = 8'b00000000; //  225 :   0 - 0x0
      13'hE2: dout  = 8'b00111000; //  226 :  56 - 0x38
      13'hE3: dout  = 8'b11000000; //  227 : 192 - 0xc0
      13'hE4: dout  = 8'b11100000; //  228 : 224 - 0xe0
      13'hE5: dout  = 8'b11010000; //  229 : 208 - 0xd0
      13'hE6: dout  = 8'b11111100; //  230 : 252 - 0xfc
      13'hE7: dout  = 8'b11000000; //  231 : 192 - 0xc0
      13'hE8: dout  = 8'b11000000; //  232 : 192 - 0xc0
      13'hE9: dout  = 8'b11000000; //  233 : 192 - 0xc0
      13'hEA: dout  = 8'b11111000; //  234 : 248 - 0xf8
      13'hEB: dout  = 8'b00100000; //  235 :  32 - 0x20
      13'hEC: dout  = 8'b00011100; //  236 :  28 - 0x1c
      13'hED: dout  = 8'b00101110; //  237 :  46 - 0x2e
      13'hEE: dout  = 8'b00000000; //  238 :   0 - 0x0
      13'hEF: dout  = 8'b00111000; //  239 :  56 - 0x38
      13'hF0: dout  = 8'b11100000; //  240 : 224 - 0xe0 -- Sprite 0xf
      13'hF1: dout  = 8'b11100000; //  241 : 224 - 0xe0
      13'hF2: dout  = 8'b10110000; //  242 : 176 - 0xb0
      13'hF3: dout  = 8'b11110000; //  243 : 240 - 0xf0
      13'hF4: dout  = 8'b11110000; //  244 : 240 - 0xf0
      13'hF5: dout  = 8'b11100000; //  245 : 224 - 0xe0
      13'hF6: dout  = 8'b11000000; //  246 : 192 - 0xc0
      13'hF7: dout  = 8'b11100000; //  247 : 224 - 0xe0
      13'hF8: dout  = 8'b00000000; //  248 :   0 - 0x0
      13'hF9: dout  = 8'b01100000; //  249 :  96 - 0x60
      13'hFA: dout  = 8'b11110000; //  250 : 240 - 0xf0
      13'hFB: dout  = 8'b11110000; //  251 : 240 - 0xf0
      13'hFC: dout  = 8'b11110000; //  252 : 240 - 0xf0
      13'hFD: dout  = 8'b11100000; //  253 : 224 - 0xe0
      13'hFE: dout  = 8'b00000000; //  254 :   0 - 0x0
      13'hFF: dout  = 8'b00000000; //  255 :   0 - 0x0
      13'h100: dout  = 8'b00000000; //  256 :   0 - 0x0 -- Sprite 0x10
      13'h101: dout  = 8'b00000011; //  257 :   3 - 0x3
      13'h102: dout  = 8'b00000111; //  258 :   7 - 0x7
      13'h103: dout  = 8'b00000111; //  259 :   7 - 0x7
      13'h104: dout  = 8'b00001001; //  260 :   9 - 0x9
      13'h105: dout  = 8'b00001001; //  261 :   9 - 0x9
      13'h106: dout  = 8'b00011100; //  262 :  28 - 0x1c
      13'h107: dout  = 8'b00000000; //  263 :   0 - 0x0
      13'h108: dout  = 8'b00000000; //  264 :   0 - 0x0
      13'h109: dout  = 8'b00000011; //  265 :   3 - 0x3
      13'h10A: dout  = 8'b00000111; //  266 :   7 - 0x7
      13'h10B: dout  = 8'b00000000; //  267 :   0 - 0x0
      13'h10C: dout  = 8'b00000110; //  268 :   6 - 0x6
      13'h10D: dout  = 8'b00000110; //  269 :   6 - 0x6
      13'h10E: dout  = 8'b00000011; //  270 :   3 - 0x3
      13'h10F: dout  = 8'b00000011; //  271 :   3 - 0x3
      13'h110: dout  = 8'b00001111; //  272 :  15 - 0xf -- Sprite 0x11
      13'h111: dout  = 8'b00001111; //  273 :  15 - 0xf
      13'h112: dout  = 8'b00001111; //  274 :  15 - 0xf
      13'h113: dout  = 8'b11111111; //  275 : 255 - 0xff
      13'h114: dout  = 8'b11111111; //  276 : 255 - 0xff
      13'h115: dout  = 8'b11111100; //  277 : 252 - 0xfc
      13'h116: dout  = 8'b10000001; //  278 : 129 - 0x81
      13'h117: dout  = 8'b00000001; //  279 :   1 - 0x1
      13'h118: dout  = 8'b00000000; //  280 :   0 - 0x0
      13'h119: dout  = 8'b00000000; //  281 :   0 - 0x0
      13'h11A: dout  = 8'b00001100; //  282 :  12 - 0xc
      13'h11B: dout  = 8'b00111111; //  283 :  63 - 0x3f
      13'h11C: dout  = 8'b00111111; //  284 :  63 - 0x3f
      13'h11D: dout  = 8'b00111100; //  285 :  60 - 0x3c
      13'h11E: dout  = 8'b00000000; //  286 :   0 - 0x0
      13'h11F: dout  = 8'b00000000; //  287 :   0 - 0x0
      13'h120: dout  = 8'b00000000; //  288 :   0 - 0x0 -- Sprite 0x12
      13'h121: dout  = 8'b11000000; //  289 : 192 - 0xc0
      13'h122: dout  = 8'b11111000; //  290 : 248 - 0xf8
      13'h123: dout  = 8'b10000000; //  291 : 128 - 0x80
      13'h124: dout  = 8'b00100000; //  292 :  32 - 0x20
      13'h125: dout  = 8'b10010000; //  293 : 144 - 0x90
      13'h126: dout  = 8'b00111100; //  294 :  60 - 0x3c
      13'h127: dout  = 8'b00000000; //  295 :   0 - 0x0
      13'h128: dout  = 8'b00000000; //  296 :   0 - 0x0
      13'h129: dout  = 8'b11000000; //  297 : 192 - 0xc0
      13'h12A: dout  = 8'b11111000; //  298 : 248 - 0xf8
      13'h12B: dout  = 8'b01100000; //  299 :  96 - 0x60
      13'h12C: dout  = 8'b11011100; //  300 : 220 - 0xdc
      13'h12D: dout  = 8'b01101110; //  301 : 110 - 0x6e
      13'h12E: dout  = 8'b11000000; //  302 : 192 - 0xc0
      13'h12F: dout  = 8'b11111000; //  303 : 248 - 0xf8
      13'h130: dout  = 8'b11100000; //  304 : 224 - 0xe0 -- Sprite 0x13
      13'h131: dout  = 8'b11110000; //  305 : 240 - 0xf0
      13'h132: dout  = 8'b11110000; //  306 : 240 - 0xf0
      13'h133: dout  = 8'b11110000; //  307 : 240 - 0xf0
      13'h134: dout  = 8'b11110000; //  308 : 240 - 0xf0
      13'h135: dout  = 8'b11100000; //  309 : 224 - 0xe0
      13'h136: dout  = 8'b11000000; //  310 : 192 - 0xc0
      13'h137: dout  = 8'b11100000; //  311 : 224 - 0xe0
      13'h138: dout  = 8'b01000111; //  312 :  71 - 0x47
      13'h139: dout  = 8'b00001111; //  313 :  15 - 0xf
      13'h13A: dout  = 8'b00001110; //  314 :  14 - 0xe
      13'h13B: dout  = 8'b11110000; //  315 : 240 - 0xf0
      13'h13C: dout  = 8'b11110000; //  316 : 240 - 0xf0
      13'h13D: dout  = 8'b11100000; //  317 : 224 - 0xe0
      13'h13E: dout  = 8'b00000000; //  318 :   0 - 0x0
      13'h13F: dout  = 8'b00000000; //  319 :   0 - 0x0
      13'h140: dout  = 8'b00000100; //  320 :   4 - 0x4 -- Sprite 0x14
      13'h141: dout  = 8'b00001100; //  321 :  12 - 0xc
      13'h142: dout  = 8'b00001100; //  322 :  12 - 0xc
      13'h143: dout  = 8'b00010011; //  323 :  19 - 0x13
      13'h144: dout  = 8'b00010011; //  324 :  19 - 0x13
      13'h145: dout  = 8'b00111011; //  325 :  59 - 0x3b
      13'h146: dout  = 8'b00000111; //  326 :   7 - 0x7
      13'h147: dout  = 8'b00001111; //  327 :  15 - 0xf
      13'h148: dout  = 8'b00000111; //  328 :   7 - 0x7
      13'h149: dout  = 8'b00001111; //  329 :  15 - 0xf
      13'h14A: dout  = 8'b00000011; //  330 :   3 - 0x3
      13'h14B: dout  = 8'b00001100; //  331 :  12 - 0xc
      13'h14C: dout  = 8'b00001100; //  332 :  12 - 0xc
      13'h14D: dout  = 8'b00000100; //  333 :   4 - 0x4
      13'h14E: dout  = 8'b00000000; //  334 :   0 - 0x0
      13'h14F: dout  = 8'b00000000; //  335 :   0 - 0x0
      13'h150: dout  = 8'b00001111; //  336 :  15 - 0xf -- Sprite 0x15
      13'h151: dout  = 8'b00001111; //  337 :  15 - 0xf
      13'h152: dout  = 8'b00001111; //  338 :  15 - 0xf
      13'h153: dout  = 8'b00011111; //  339 :  31 - 0x1f
      13'h154: dout  = 8'b00011111; //  340 :  31 - 0x1f
      13'h155: dout  = 8'b00011110; //  341 :  30 - 0x1e
      13'h156: dout  = 8'b00011100; //  342 :  28 - 0x1c
      13'h157: dout  = 8'b00011110; //  343 :  30 - 0x1e
      13'h158: dout  = 8'b00000000; //  344 :   0 - 0x0
      13'h159: dout  = 8'b00000001; //  345 :   1 - 0x1
      13'h15A: dout  = 8'b00001111; //  346 :  15 - 0xf
      13'h15B: dout  = 8'b00011111; //  347 :  31 - 0x1f
      13'h15C: dout  = 8'b00011111; //  348 :  31 - 0x1f
      13'h15D: dout  = 8'b00011110; //  349 :  30 - 0x1e
      13'h15E: dout  = 8'b00000000; //  350 :   0 - 0x0
      13'h15F: dout  = 8'b00000000; //  351 :   0 - 0x0
      13'h160: dout  = 8'b00000000; //  352 :   0 - 0x0 -- Sprite 0x16
      13'h161: dout  = 8'b01110000; //  353 : 112 - 0x70
      13'h162: dout  = 8'b00000000; //  354 :   0 - 0x0
      13'h163: dout  = 8'b11000000; //  355 : 192 - 0xc0
      13'h164: dout  = 8'b10100000; //  356 : 160 - 0xa0
      13'h165: dout  = 8'b11111000; //  357 : 248 - 0xf8
      13'h166: dout  = 8'b10000000; //  358 : 128 - 0x80
      13'h167: dout  = 8'b11000000; //  359 : 192 - 0xc0
      13'h168: dout  = 8'b10000000; //  360 : 128 - 0x80
      13'h169: dout  = 8'b11110000; //  361 : 240 - 0xf0
      13'h16A: dout  = 8'b11000000; //  362 : 192 - 0xc0
      13'h16B: dout  = 8'b00111000; //  363 :  56 - 0x38
      13'h16C: dout  = 8'b01011100; //  364 :  92 - 0x5c
      13'h16D: dout  = 8'b00000000; //  365 :   0 - 0x0
      13'h16E: dout  = 8'b01110000; //  366 : 112 - 0x70
      13'h16F: dout  = 8'b01000000; //  367 :  64 - 0x40
      13'h170: dout  = 8'b11100000; //  368 : 224 - 0xe0 -- Sprite 0x17
      13'h171: dout  = 8'b01100000; //  369 :  96 - 0x60
      13'h172: dout  = 8'b11110000; //  370 : 240 - 0xf0
      13'h173: dout  = 8'b11110000; //  371 : 240 - 0xf0
      13'h174: dout  = 8'b11110000; //  372 : 240 - 0xf0
      13'h175: dout  = 8'b11100000; //  373 : 224 - 0xe0
      13'h176: dout  = 8'b11100000; //  374 : 224 - 0xe0
      13'h177: dout  = 8'b11110000; //  375 : 240 - 0xf0
      13'h178: dout  = 8'b11000000; //  376 : 192 - 0xc0
      13'h179: dout  = 8'b11100000; //  377 : 224 - 0xe0
      13'h17A: dout  = 8'b11110000; //  378 : 240 - 0xf0
      13'h17B: dout  = 8'b11110000; //  379 : 240 - 0xf0
      13'h17C: dout  = 8'b11110000; //  380 : 240 - 0xf0
      13'h17D: dout  = 8'b11100000; //  381 : 224 - 0xe0
      13'h17E: dout  = 8'b00000000; //  382 :   0 - 0x0
      13'h17F: dout  = 8'b00000000; //  383 :   0 - 0x0
      13'h180: dout  = 8'b00000111; //  384 :   7 - 0x7 -- Sprite 0x18
      13'h181: dout  = 8'b00001111; //  385 :  15 - 0xf
      13'h182: dout  = 8'b00001111; //  386 :  15 - 0xf
      13'h183: dout  = 8'b00010010; //  387 :  18 - 0x12
      13'h184: dout  = 8'b00010011; //  388 :  19 - 0x13
      13'h185: dout  = 8'b00111000; //  389 :  56 - 0x38
      13'h186: dout  = 8'b00000000; //  390 :   0 - 0x0
      13'h187: dout  = 8'b00001111; //  391 :  15 - 0xf
      13'h188: dout  = 8'b00000111; //  392 :   7 - 0x7
      13'h189: dout  = 8'b00001111; //  393 :  15 - 0xf
      13'h18A: dout  = 8'b00000000; //  394 :   0 - 0x0
      13'h18B: dout  = 8'b00001101; //  395 :  13 - 0xd
      13'h18C: dout  = 8'b00001100; //  396 :  12 - 0xc
      13'h18D: dout  = 8'b00000111; //  397 :   7 - 0x7
      13'h18E: dout  = 8'b00000111; //  398 :   7 - 0x7
      13'h18F: dout  = 8'b00000001; //  399 :   1 - 0x1
      13'h190: dout  = 8'b00011111; //  400 :  31 - 0x1f -- Sprite 0x19
      13'h191: dout  = 8'b00011111; //  401 :  31 - 0x1f
      13'h192: dout  = 8'b00011111; //  402 :  31 - 0x1f
      13'h193: dout  = 8'b00011111; //  403 :  31 - 0x1f
      13'h194: dout  = 8'b00011111; //  404 :  31 - 0x1f
      13'h195: dout  = 8'b00011110; //  405 :  30 - 0x1e
      13'h196: dout  = 8'b00011100; //  406 :  28 - 0x1c
      13'h197: dout  = 8'b00011110; //  407 :  30 - 0x1e
      13'h198: dout  = 8'b00000000; //  408 :   0 - 0x0
      13'h199: dout  = 8'b00000000; //  409 :   0 - 0x0
      13'h19A: dout  = 8'b00010011; //  410 :  19 - 0x13
      13'h19B: dout  = 8'b00011111; //  411 :  31 - 0x1f
      13'h19C: dout  = 8'b00011111; //  412 :  31 - 0x1f
      13'h19D: dout  = 8'b00011110; //  413 :  30 - 0x1e
      13'h19E: dout  = 8'b00000000; //  414 :   0 - 0x0
      13'h19F: dout  = 8'b00000000; //  415 :   0 - 0x0
      13'h1A0: dout  = 8'b10000000; //  416 : 128 - 0x80 -- Sprite 0x1a
      13'h1A1: dout  = 8'b11110000; //  417 : 240 - 0xf0
      13'h1A2: dout  = 8'b00000000; //  418 :   0 - 0x0
      13'h1A3: dout  = 8'b01000000; //  419 :  64 - 0x40
      13'h1A4: dout  = 8'b00100000; //  420 :  32 - 0x20
      13'h1A5: dout  = 8'b01111000; //  421 : 120 - 0x78
      13'h1A6: dout  = 8'b00000000; //  422 :   0 - 0x0
      13'h1A7: dout  = 8'b11000000; //  423 : 192 - 0xc0
      13'h1A8: dout  = 8'b10000000; //  424 : 128 - 0x80
      13'h1A9: dout  = 8'b11110000; //  425 : 240 - 0xf0
      13'h1AA: dout  = 8'b11000000; //  426 : 192 - 0xc0
      13'h1AB: dout  = 8'b10111000; //  427 : 184 - 0xb8
      13'h1AC: dout  = 8'b11011100; //  428 : 220 - 0xdc
      13'h1AD: dout  = 8'b10000000; //  429 : 128 - 0x80
      13'h1AE: dout  = 8'b11110000; //  430 : 240 - 0xf0
      13'h1AF: dout  = 8'b10000000; //  431 : 128 - 0x80
      13'h1B0: dout  = 8'b11111000; //  432 : 248 - 0xf8 -- Sprite 0x1b
      13'h1B1: dout  = 8'b11111000; //  433 : 248 - 0xf8
      13'h1B2: dout  = 8'b11110000; //  434 : 240 - 0xf0
      13'h1B3: dout  = 8'b11110000; //  435 : 240 - 0xf0
      13'h1B4: dout  = 8'b11110000; //  436 : 240 - 0xf0
      13'h1B5: dout  = 8'b11100000; //  437 : 224 - 0xe0
      13'h1B6: dout  = 8'b11100000; //  438 : 224 - 0xe0
      13'h1B7: dout  = 8'b11110000; //  439 : 240 - 0xf0
      13'h1B8: dout  = 8'b00000111; //  440 :   7 - 0x7
      13'h1B9: dout  = 8'b00000111; //  441 :   7 - 0x7
      13'h1BA: dout  = 8'b11111110; //  442 : 254 - 0xfe
      13'h1BB: dout  = 8'b11110000; //  443 : 240 - 0xf0
      13'h1BC: dout  = 8'b11110000; //  444 : 240 - 0xf0
      13'h1BD: dout  = 8'b11100000; //  445 : 224 - 0xe0
      13'h1BE: dout  = 8'b00000000; //  446 :   0 - 0x0
      13'h1BF: dout  = 8'b00000000; //  447 :   0 - 0x0
      13'h1C0: dout  = 8'b00000100; //  448 :   4 - 0x4 -- Sprite 0x1c
      13'h1C1: dout  = 8'b00001100; //  449 :  12 - 0xc
      13'h1C2: dout  = 8'b00001100; //  450 :  12 - 0xc
      13'h1C3: dout  = 8'b00010011; //  451 :  19 - 0x13
      13'h1C4: dout  = 8'b00010011; //  452 :  19 - 0x13
      13'h1C5: dout  = 8'b00111111; //  453 :  63 - 0x3f
      13'h1C6: dout  = 8'b00000111; //  454 :   7 - 0x7
      13'h1C7: dout  = 8'b00001111; //  455 :  15 - 0xf
      13'h1C8: dout  = 8'b00000111; //  456 :   7 - 0x7
      13'h1C9: dout  = 8'b00001111; //  457 :  15 - 0xf
      13'h1CA: dout  = 8'b00000011; //  458 :   3 - 0x3
      13'h1CB: dout  = 8'b00001100; //  459 :  12 - 0xc
      13'h1CC: dout  = 8'b00001100; //  460 :  12 - 0xc
      13'h1CD: dout  = 8'b00000000; //  461 :   0 - 0x0
      13'h1CE: dout  = 8'b00000000; //  462 :   0 - 0x0
      13'h1CF: dout  = 8'b00000000; //  463 :   0 - 0x0
      13'h1D0: dout  = 8'b00001111; //  464 :  15 - 0xf -- Sprite 0x1d
      13'h1D1: dout  = 8'b00001111; //  465 :  15 - 0xf
      13'h1D2: dout  = 8'b00001111; //  466 :  15 - 0xf
      13'h1D3: dout  = 8'b00011111; //  467 :  31 - 0x1f
      13'h1D4: dout  = 8'b00111111; //  468 :  63 - 0x3f
      13'h1D5: dout  = 8'b01111100; //  469 : 124 - 0x7c
      13'h1D6: dout  = 8'b01110000; //  470 : 112 - 0x70
      13'h1D7: dout  = 8'b00111000; //  471 :  56 - 0x38
      13'h1D8: dout  = 8'b00000001; //  472 :   1 - 0x1
      13'h1D9: dout  = 8'b00000001; //  473 :   1 - 0x1
      13'h1DA: dout  = 8'b00001111; //  474 :  15 - 0xf
      13'h1DB: dout  = 8'b00011111; //  475 :  31 - 0x1f
      13'h1DC: dout  = 8'b00111111; //  476 :  63 - 0x3f
      13'h1DD: dout  = 8'b00011100; //  477 :  28 - 0x1c
      13'h1DE: dout  = 8'b00000000; //  478 :   0 - 0x0
      13'h1DF: dout  = 8'b00000000; //  479 :   0 - 0x0
      13'h1E0: dout  = 8'b00000000; //  480 :   0 - 0x0 -- Sprite 0x1e
      13'h1E1: dout  = 8'b01110000; //  481 : 112 - 0x70
      13'h1E2: dout  = 8'b00000000; //  482 :   0 - 0x0
      13'h1E3: dout  = 8'b11000000; //  483 : 192 - 0xc0
      13'h1E4: dout  = 8'b10100000; //  484 : 160 - 0xa0
      13'h1E5: dout  = 8'b11111000; //  485 : 248 - 0xf8
      13'h1E6: dout  = 8'b10000000; //  486 : 128 - 0x80
      13'h1E7: dout  = 8'b11000000; //  487 : 192 - 0xc0
      13'h1E8: dout  = 8'b10000000; //  488 : 128 - 0x80
      13'h1E9: dout  = 8'b11110000; //  489 : 240 - 0xf0
      13'h1EA: dout  = 8'b11000000; //  490 : 192 - 0xc0
      13'h1EB: dout  = 8'b00111000; //  491 :  56 - 0x38
      13'h1EC: dout  = 8'b01011100; //  492 :  92 - 0x5c
      13'h1ED: dout  = 8'b00000000; //  493 :   0 - 0x0
      13'h1EE: dout  = 8'b01110000; //  494 : 112 - 0x70
      13'h1EF: dout  = 8'b01000000; //  495 :  64 - 0x40
      13'h1F0: dout  = 8'b11000000; //  496 : 192 - 0xc0 -- Sprite 0x1f
      13'h1F1: dout  = 8'b01100000; //  497 :  96 - 0x60
      13'h1F2: dout  = 8'b11100100; //  498 : 228 - 0xe4
      13'h1F3: dout  = 8'b11111100; //  499 : 252 - 0xfc
      13'h1F4: dout  = 8'b11111100; //  500 : 252 - 0xfc
      13'h1F5: dout  = 8'b01111100; //  501 : 124 - 0x7c
      13'h1F6: dout  = 8'b00000000; //  502 :   0 - 0x0
      13'h1F7: dout  = 8'b00000000; //  503 :   0 - 0x0
      13'h1F8: dout  = 8'b11000000; //  504 : 192 - 0xc0
      13'h1F9: dout  = 8'b11100000; //  505 : 224 - 0xe0
      13'h1FA: dout  = 8'b11100000; //  506 : 224 - 0xe0
      13'h1FB: dout  = 8'b11110000; //  507 : 240 - 0xf0
      13'h1FC: dout  = 8'b11110000; //  508 : 240 - 0xf0
      13'h1FD: dout  = 8'b01110000; //  509 : 112 - 0x70
      13'h1FE: dout  = 8'b00000000; //  510 :   0 - 0x0
      13'h1FF: dout  = 8'b00000000; //  511 :   0 - 0x0
      13'h200: dout  = 8'b00000111; //  512 :   7 - 0x7 -- Sprite 0x20
      13'h201: dout  = 8'b00001111; //  513 :  15 - 0xf
      13'h202: dout  = 8'b00001111; //  514 :  15 - 0xf
      13'h203: dout  = 8'b00010010; //  515 :  18 - 0x12
      13'h204: dout  = 8'b00010011; //  516 :  19 - 0x13
      13'h205: dout  = 8'b00111000; //  517 :  56 - 0x38
      13'h206: dout  = 8'b00000000; //  518 :   0 - 0x0
      13'h207: dout  = 8'b00000111; //  519 :   7 - 0x7
      13'h208: dout  = 8'b00000111; //  520 :   7 - 0x7
      13'h209: dout  = 8'b00001111; //  521 :  15 - 0xf
      13'h20A: dout  = 8'b00000000; //  522 :   0 - 0x0
      13'h20B: dout  = 8'b00001101; //  523 :  13 - 0xd
      13'h20C: dout  = 8'b00001100; //  524 :  12 - 0xc
      13'h20D: dout  = 8'b00000111; //  525 :   7 - 0x7
      13'h20E: dout  = 8'b00000111; //  526 :   7 - 0x7
      13'h20F: dout  = 8'b00000001; //  527 :   1 - 0x1
      13'h210: dout  = 8'b00001111; //  528 :  15 - 0xf -- Sprite 0x21
      13'h211: dout  = 8'b00001111; //  529 :  15 - 0xf
      13'h212: dout  = 8'b00001111; //  530 :  15 - 0xf
      13'h213: dout  = 8'b00011111; //  531 :  31 - 0x1f
      13'h214: dout  = 8'b00111111; //  532 :  63 - 0x3f
      13'h215: dout  = 8'b01111100; //  533 : 124 - 0x7c
      13'h216: dout  = 8'b01110000; //  534 : 112 - 0x70
      13'h217: dout  = 8'b00111000; //  535 :  56 - 0x38
      13'h218: dout  = 8'b00000000; //  536 :   0 - 0x0
      13'h219: dout  = 8'b00000000; //  537 :   0 - 0x0
      13'h21A: dout  = 8'b00001001; //  538 :   9 - 0x9
      13'h21B: dout  = 8'b00011111; //  539 :  31 - 0x1f
      13'h21C: dout  = 8'b00111111; //  540 :  63 - 0x3f
      13'h21D: dout  = 8'b00011100; //  541 :  28 - 0x1c
      13'h21E: dout  = 8'b00000000; //  542 :   0 - 0x0
      13'h21F: dout  = 8'b00000000; //  543 :   0 - 0x0
      13'h220: dout  = 8'b10000000; //  544 : 128 - 0x80 -- Sprite 0x22
      13'h221: dout  = 8'b11110000; //  545 : 240 - 0xf0
      13'h222: dout  = 8'b00000000; //  546 :   0 - 0x0
      13'h223: dout  = 8'b01000000; //  547 :  64 - 0x40
      13'h224: dout  = 8'b00100000; //  548 :  32 - 0x20
      13'h225: dout  = 8'b01111000; //  549 : 120 - 0x78
      13'h226: dout  = 8'b00000000; //  550 :   0 - 0x0
      13'h227: dout  = 8'b11000000; //  551 : 192 - 0xc0
      13'h228: dout  = 8'b10000000; //  552 : 128 - 0x80
      13'h229: dout  = 8'b11110000; //  553 : 240 - 0xf0
      13'h22A: dout  = 8'b11000000; //  554 : 192 - 0xc0
      13'h22B: dout  = 8'b10111000; //  555 : 184 - 0xb8
      13'h22C: dout  = 8'b11011100; //  556 : 220 - 0xdc
      13'h22D: dout  = 8'b10000000; //  557 : 128 - 0x80
      13'h22E: dout  = 8'b11110000; //  558 : 240 - 0xf0
      13'h22F: dout  = 8'b10000000; //  559 : 128 - 0x80
      13'h230: dout  = 8'b11111000; //  560 : 248 - 0xf8 -- Sprite 0x23
      13'h231: dout  = 8'b11111000; //  561 : 248 - 0xf8
      13'h232: dout  = 8'b11100000; //  562 : 224 - 0xe0
      13'h233: dout  = 8'b11111100; //  563 : 252 - 0xfc
      13'h234: dout  = 8'b11111100; //  564 : 252 - 0xfc
      13'h235: dout  = 8'b01111100; //  565 : 124 - 0x7c
      13'h236: dout  = 8'b00000000; //  566 :   0 - 0x0
      13'h237: dout  = 8'b00000000; //  567 :   0 - 0x0
      13'h238: dout  = 8'b00000111; //  568 :   7 - 0x7
      13'h239: dout  = 8'b00000111; //  569 :   7 - 0x7
      13'h23A: dout  = 8'b11101110; //  570 : 238 - 0xee
      13'h23B: dout  = 8'b11110000; //  571 : 240 - 0xf0
      13'h23C: dout  = 8'b11110000; //  572 : 240 - 0xf0
      13'h23D: dout  = 8'b01110000; //  573 : 112 - 0x70
      13'h23E: dout  = 8'b00000000; //  574 :   0 - 0x0
      13'h23F: dout  = 8'b00000000; //  575 :   0 - 0x0
      13'h240: dout  = 8'b00000000; //  576 :   0 - 0x0 -- Sprite 0x24
      13'h241: dout  = 8'b00000111; //  577 :   7 - 0x7
      13'h242: dout  = 8'b00000111; //  578 :   7 - 0x7
      13'h243: dout  = 8'b00001111; //  579 :  15 - 0xf
      13'h244: dout  = 8'b00001111; //  580 :  15 - 0xf
      13'h245: dout  = 8'b00111000; //  581 :  56 - 0x38
      13'h246: dout  = 8'b01111111; //  582 : 127 - 0x7f
      13'h247: dout  = 8'b01111111; //  583 : 127 - 0x7f
      13'h248: dout  = 8'b00000000; //  584 :   0 - 0x0
      13'h249: dout  = 8'b00000111; //  585 :   7 - 0x7
      13'h24A: dout  = 8'b00000011; //  586 :   3 - 0x3
      13'h24B: dout  = 8'b00000000; //  587 :   0 - 0x0
      13'h24C: dout  = 8'b00000000; //  588 :   0 - 0x0
      13'h24D: dout  = 8'b00000111; //  589 :   7 - 0x7
      13'h24E: dout  = 8'b00000100; //  590 :   4 - 0x4
      13'h24F: dout  = 8'b00000100; //  591 :   4 - 0x4
      13'h250: dout  = 8'b00011111; //  592 :  31 - 0x1f -- Sprite 0x25
      13'h251: dout  = 8'b00011111; //  593 :  31 - 0x1f
      13'h252: dout  = 8'b00011111; //  594 :  31 - 0x1f
      13'h253: dout  = 8'b00011111; //  595 :  31 - 0x1f
      13'h254: dout  = 8'b00001111; //  596 :  15 - 0xf
      13'h255: dout  = 8'b00001111; //  597 :  15 - 0xf
      13'h256: dout  = 8'b00001111; //  598 :  15 - 0xf
      13'h257: dout  = 8'b00000111; //  599 :   7 - 0x7
      13'h258: dout  = 8'b00011110; //  600 :  30 - 0x1e
      13'h259: dout  = 8'b00011111; //  601 :  31 - 0x1f
      13'h25A: dout  = 8'b00011111; //  602 :  31 - 0x1f
      13'h25B: dout  = 8'b00011111; //  603 :  31 - 0x1f
      13'h25C: dout  = 8'b00001111; //  604 :  15 - 0xf
      13'h25D: dout  = 8'b00001000; //  605 :   8 - 0x8
      13'h25E: dout  = 8'b00000000; //  606 :   0 - 0x0
      13'h25F: dout  = 8'b00000000; //  607 :   0 - 0x0
      13'h260: dout  = 8'b00000000; //  608 :   0 - 0x0 -- Sprite 0x26
      13'h261: dout  = 8'b11100000; //  609 : 224 - 0xe0
      13'h262: dout  = 8'b11111000; //  610 : 248 - 0xf8
      13'h263: dout  = 8'b11111100; //  611 : 252 - 0xfc
      13'h264: dout  = 8'b11111100; //  612 : 252 - 0xfc
      13'h265: dout  = 8'b00011100; //  613 :  28 - 0x1c
      13'h266: dout  = 8'b11111000; //  614 : 248 - 0xf8
      13'h267: dout  = 8'b11111000; //  615 : 248 - 0xf8
      13'h268: dout  = 8'b00111000; //  616 :  56 - 0x38
      13'h269: dout  = 8'b11111000; //  617 : 248 - 0xf8
      13'h26A: dout  = 8'b11000000; //  618 : 192 - 0xc0
      13'h26B: dout  = 8'b00000000; //  619 :   0 - 0x0
      13'h26C: dout  = 8'b00000000; //  620 :   0 - 0x0
      13'h26D: dout  = 8'b11100000; //  621 : 224 - 0xe0
      13'h26E: dout  = 8'b00100000; //  622 :  32 - 0x20
      13'h26F: dout  = 8'b00100000; //  623 :  32 - 0x20
      13'h270: dout  = 8'b11111000; //  624 : 248 - 0xf8 -- Sprite 0x27
      13'h271: dout  = 8'b11111100; //  625 : 252 - 0xfc
      13'h272: dout  = 8'b11111100; //  626 : 252 - 0xfc
      13'h273: dout  = 8'b11111000; //  627 : 248 - 0xf8
      13'h274: dout  = 8'b01111000; //  628 : 120 - 0x78
      13'h275: dout  = 8'b10000000; //  629 : 128 - 0x80
      13'h276: dout  = 8'b11000000; //  630 : 192 - 0xc0
      13'h277: dout  = 8'b11000000; //  631 : 192 - 0xc0
      13'h278: dout  = 8'b01111000; //  632 : 120 - 0x78
      13'h279: dout  = 8'b11111100; //  633 : 252 - 0xfc
      13'h27A: dout  = 8'b11111100; //  634 : 252 - 0xfc
      13'h27B: dout  = 8'b11111000; //  635 : 248 - 0xf8
      13'h27C: dout  = 8'b00000000; //  636 :   0 - 0x0
      13'h27D: dout  = 8'b10000000; //  637 : 128 - 0x80
      13'h27E: dout  = 8'b00000000; //  638 :   0 - 0x0
      13'h27F: dout  = 8'b00000000; //  639 :   0 - 0x0
      13'h280: dout  = 8'b00000000; //  640 :   0 - 0x0 -- Sprite 0x28
      13'h281: dout  = 8'b00000011; //  641 :   3 - 0x3
      13'h282: dout  = 8'b00000111; //  642 :   7 - 0x7
      13'h283: dout  = 8'b00000111; //  643 :   7 - 0x7
      13'h284: dout  = 8'b00001001; //  644 :   9 - 0x9
      13'h285: dout  = 8'b00001001; //  645 :   9 - 0x9
      13'h286: dout  = 8'b00011100; //  646 :  28 - 0x1c
      13'h287: dout  = 8'b00000000; //  647 :   0 - 0x0
      13'h288: dout  = 8'b00000000; //  648 :   0 - 0x0
      13'h289: dout  = 8'b00000011; //  649 :   3 - 0x3
      13'h28A: dout  = 8'b00000111; //  650 :   7 - 0x7
      13'h28B: dout  = 8'b00000000; //  651 :   0 - 0x0
      13'h28C: dout  = 8'b00000110; //  652 :   6 - 0x6
      13'h28D: dout  = 8'b00000110; //  653 :   6 - 0x6
      13'h28E: dout  = 8'b00000011; //  654 :   3 - 0x3
      13'h28F: dout  = 8'b01100011; //  655 :  99 - 0x63
      13'h290: dout  = 8'b00011111; //  656 :  31 - 0x1f -- Sprite 0x29
      13'h291: dout  = 8'b00001111; //  657 :  15 - 0xf
      13'h292: dout  = 8'b00000111; //  658 :   7 - 0x7
      13'h293: dout  = 8'b00110111; //  659 :  55 - 0x37
      13'h294: dout  = 8'b01111111; //  660 : 127 - 0x7f
      13'h295: dout  = 8'b11011111; //  661 : 223 - 0xdf
      13'h296: dout  = 8'b00001111; //  662 :  15 - 0xf
      13'h297: dout  = 8'b00000110; //  663 :   6 - 0x6
      13'h298: dout  = 8'b11100000; //  664 : 224 - 0xe0
      13'h299: dout  = 8'b00100001; //  665 :  33 - 0x21
      13'h29A: dout  = 8'b00000001; //  666 :   1 - 0x1
      13'h29B: dout  = 8'b00000111; //  667 :   7 - 0x7
      13'h29C: dout  = 8'b00000111; //  668 :   7 - 0x7
      13'h29D: dout  = 8'b00011111; //  669 :  31 - 0x1f
      13'h29E: dout  = 8'b00001111; //  670 :  15 - 0xf
      13'h29F: dout  = 8'b00000110; //  671 :   6 - 0x6
      13'h2A0: dout  = 8'b00000000; //  672 :   0 - 0x0 -- Sprite 0x2a
      13'h2A1: dout  = 8'b11000000; //  673 : 192 - 0xc0
      13'h2A2: dout  = 8'b11111000; //  674 : 248 - 0xf8
      13'h2A3: dout  = 8'b10000000; //  675 : 128 - 0x80
      13'h2A4: dout  = 8'b00100000; //  676 :  32 - 0x20
      13'h2A5: dout  = 8'b10010000; //  677 : 144 - 0x90
      13'h2A6: dout  = 8'b00111100; //  678 :  60 - 0x3c
      13'h2A7: dout  = 8'b00000000; //  679 :   0 - 0x0
      13'h2A8: dout  = 8'b00000000; //  680 :   0 - 0x0
      13'h2A9: dout  = 8'b11000000; //  681 : 192 - 0xc0
      13'h2AA: dout  = 8'b11111000; //  682 : 248 - 0xf8
      13'h2AB: dout  = 8'b01100000; //  683 :  96 - 0x60
      13'h2AC: dout  = 8'b11011100; //  684 : 220 - 0xdc
      13'h2AD: dout  = 8'b01101110; //  685 : 110 - 0x6e
      13'h2AE: dout  = 8'b11000000; //  686 : 192 - 0xc0
      13'h2AF: dout  = 8'b11111011; //  687 : 251 - 0xfb
      13'h2B0: dout  = 8'b11100100; //  688 : 228 - 0xe4 -- Sprite 0x2b
      13'h2B1: dout  = 8'b11111110; //  689 : 254 - 0xfe
      13'h2B2: dout  = 8'b01110000; //  690 : 112 - 0x70
      13'h2B3: dout  = 8'b11110001; //  691 : 241 - 0xf1
      13'h2B4: dout  = 8'b11111111; //  692 : 255 - 0xff
      13'h2B5: dout  = 8'b11111111; //  693 : 255 - 0xff
      13'h2B6: dout  = 8'b00000000; //  694 :   0 - 0x0
      13'h2B7: dout  = 8'b00000000; //  695 :   0 - 0x0
      13'h2B8: dout  = 8'b10000011; //  696 : 131 - 0x83
      13'h2B9: dout  = 8'b11000000; //  697 : 192 - 0xc0
      13'h2BA: dout  = 8'b11110000; //  698 : 240 - 0xf0
      13'h2BB: dout  = 8'b11110000; //  699 : 240 - 0xf0
      13'h2BC: dout  = 8'b11111100; //  700 : 252 - 0xfc
      13'h2BD: dout  = 8'b11111100; //  701 : 252 - 0xfc
      13'h2BE: dout  = 8'b00000000; //  702 :   0 - 0x0
      13'h2BF: dout  = 8'b00000000; //  703 :   0 - 0x0
      13'h2C0: dout  = 8'b00000111; //  704 :   7 - 0x7 -- Sprite 0x2c
      13'h2C1: dout  = 8'b00001111; //  705 :  15 - 0xf
      13'h2C2: dout  = 8'b00001111; //  706 :  15 - 0xf
      13'h2C3: dout  = 8'b00010010; //  707 :  18 - 0x12
      13'h2C4: dout  = 8'b00010011; //  708 :  19 - 0x13
      13'h2C5: dout  = 8'b00111000; //  709 :  56 - 0x38
      13'h2C6: dout  = 8'b01110000; //  710 : 112 - 0x70
      13'h2C7: dout  = 8'b11111111; //  711 : 255 - 0xff
      13'h2C8: dout  = 8'b00000111; //  712 :   7 - 0x7
      13'h2C9: dout  = 8'b00001111; //  713 :  15 - 0xf
      13'h2CA: dout  = 8'b00000000; //  714 :   0 - 0x0
      13'h2CB: dout  = 8'b00001101; //  715 :  13 - 0xd
      13'h2CC: dout  = 8'b00001100; //  716 :  12 - 0xc
      13'h2CD: dout  = 8'b00000111; //  717 :   7 - 0x7
      13'h2CE: dout  = 8'b00001111; //  718 :  15 - 0xf
      13'h2CF: dout  = 8'b00000010; //  719 :   2 - 0x2
      13'h2D0: dout  = 8'b11011111; //  720 : 223 - 0xdf -- Sprite 0x2d
      13'h2D1: dout  = 8'b00011110; //  721 :  30 - 0x1e
      13'h2D2: dout  = 8'b00011111; //  722 :  31 - 0x1f
      13'h2D3: dout  = 8'b00011111; //  723 :  31 - 0x1f
      13'h2D4: dout  = 8'b00011111; //  724 :  31 - 0x1f
      13'h2D5: dout  = 8'b00001111; //  725 :  15 - 0xf
      13'h2D6: dout  = 8'b00000111; //  726 :   7 - 0x7
      13'h2D7: dout  = 8'b00000001; //  727 :   1 - 0x1
      13'h2D8: dout  = 8'b00000001; //  728 :   1 - 0x1
      13'h2D9: dout  = 8'b11110011; //  729 : 243 - 0xf3
      13'h2DA: dout  = 8'b01011111; //  730 :  95 - 0x5f
      13'h2DB: dout  = 8'b00011111; //  731 :  31 - 0x1f
      13'h2DC: dout  = 8'b00011111; //  732 :  31 - 0x1f
      13'h2DD: dout  = 8'b01001111; //  733 :  79 - 0x4f
      13'h2DE: dout  = 8'b00110111; //  734 :  55 - 0x37
      13'h2DF: dout  = 8'b11000000; //  735 : 192 - 0xc0
      13'h2E0: dout  = 8'b10000000; //  736 : 128 - 0x80 -- Sprite 0x2e
      13'h2E1: dout  = 8'b11110000; //  737 : 240 - 0xf0
      13'h2E2: dout  = 8'b00000000; //  738 :   0 - 0x0
      13'h2E3: dout  = 8'b01000000; //  739 :  64 - 0x40
      13'h2E4: dout  = 8'b00100000; //  740 :  32 - 0x20
      13'h2E5: dout  = 8'b01111000; //  741 : 120 - 0x78
      13'h2E6: dout  = 8'b00000000; //  742 :   0 - 0x0
      13'h2E7: dout  = 8'b11111100; //  743 : 252 - 0xfc
      13'h2E8: dout  = 8'b10000000; //  744 : 128 - 0x80
      13'h2E9: dout  = 8'b11110000; //  745 : 240 - 0xf0
      13'h2EA: dout  = 8'b11000000; //  746 : 192 - 0xc0
      13'h2EB: dout  = 8'b10111000; //  747 : 184 - 0xb8
      13'h2EC: dout  = 8'b11011100; //  748 : 220 - 0xdc
      13'h2ED: dout  = 8'b10000000; //  749 : 128 - 0x80
      13'h2EE: dout  = 8'b11110000; //  750 : 240 - 0xf0
      13'h2EF: dout  = 8'b00000000; //  751 :   0 - 0x0
      13'h2F0: dout  = 8'b11110000; //  752 : 240 - 0xf0 -- Sprite 0x2f
      13'h2F1: dout  = 8'b11100000; //  753 : 224 - 0xe0
      13'h2F2: dout  = 8'b11100000; //  754 : 224 - 0xe0
      13'h2F3: dout  = 8'b11110000; //  755 : 240 - 0xf0
      13'h2F4: dout  = 8'b11111010; //  756 : 250 - 0xfa
      13'h2F5: dout  = 8'b11111110; //  757 : 254 - 0xfe
      13'h2F6: dout  = 8'b11111100; //  758 : 252 - 0xfc
      13'h2F7: dout  = 8'b11011000; //  759 : 216 - 0xd8
      13'h2F8: dout  = 8'b10001111; //  760 : 143 - 0x8f
      13'h2F9: dout  = 8'b11100111; //  761 : 231 - 0xe7
      13'h2FA: dout  = 8'b11100000; //  762 : 224 - 0xe0
      13'h2FB: dout  = 8'b11110000; //  763 : 240 - 0xf0
      13'h2FC: dout  = 8'b11001000; //  764 : 200 - 0xc8
      13'h2FD: dout  = 8'b10001000; //  765 : 136 - 0x88
      13'h2FE: dout  = 8'b00010000; //  766 :  16 - 0x10
      13'h2FF: dout  = 8'b00000000; //  767 :   0 - 0x0
      13'h300: dout  = 8'b00000000; //  768 :   0 - 0x0 -- Sprite 0x30
      13'h301: dout  = 8'b00000000; //  769 :   0 - 0x0
      13'h302: dout  = 8'b00000111; //  770 :   7 - 0x7
      13'h303: dout  = 8'b00001000; //  771 :   8 - 0x8
      13'h304: dout  = 8'b00010000; //  772 :  16 - 0x10
      13'h305: dout  = 8'b00100000; //  773 :  32 - 0x20
      13'h306: dout  = 8'b01000000; //  774 :  64 - 0x40
      13'h307: dout  = 8'b01000000; //  775 :  64 - 0x40
      13'h308: dout  = 8'b00000000; //  776 :   0 - 0x0
      13'h309: dout  = 8'b00000000; //  777 :   0 - 0x0
      13'h30A: dout  = 8'b00000000; //  778 :   0 - 0x0
      13'h30B: dout  = 8'b00000111; //  779 :   7 - 0x7
      13'h30C: dout  = 8'b00001000; //  780 :   8 - 0x8
      13'h30D: dout  = 8'b00010000; //  781 :  16 - 0x10
      13'h30E: dout  = 8'b00100000; //  782 :  32 - 0x20
      13'h30F: dout  = 8'b00100000; //  783 :  32 - 0x20
      13'h310: dout  = 8'b01000000; //  784 :  64 - 0x40 -- Sprite 0x31
      13'h311: dout  = 8'b01000000; //  785 :  64 - 0x40
      13'h312: dout  = 8'b00100000; //  786 :  32 - 0x20
      13'h313: dout  = 8'b00010000; //  787 :  16 - 0x10
      13'h314: dout  = 8'b00001000; //  788 :   8 - 0x8
      13'h315: dout  = 8'b00000111; //  789 :   7 - 0x7
      13'h316: dout  = 8'b00000000; //  790 :   0 - 0x0
      13'h317: dout  = 8'b00000000; //  791 :   0 - 0x0
      13'h318: dout  = 8'b00100000; //  792 :  32 - 0x20
      13'h319: dout  = 8'b00100000; //  793 :  32 - 0x20
      13'h31A: dout  = 8'b00010000; //  794 :  16 - 0x10
      13'h31B: dout  = 8'b00001000; //  795 :   8 - 0x8
      13'h31C: dout  = 8'b00000111; //  796 :   7 - 0x7
      13'h31D: dout  = 8'b00000000; //  797 :   0 - 0x0
      13'h31E: dout  = 8'b00000000; //  798 :   0 - 0x0
      13'h31F: dout  = 8'b00000000; //  799 :   0 - 0x0
      13'h320: dout  = 8'b00000000; //  800 :   0 - 0x0 -- Sprite 0x32
      13'h321: dout  = 8'b00000000; //  801 :   0 - 0x0
      13'h322: dout  = 8'b11100000; //  802 : 224 - 0xe0
      13'h323: dout  = 8'b00010000; //  803 :  16 - 0x10
      13'h324: dout  = 8'b00001000; //  804 :   8 - 0x8
      13'h325: dout  = 8'b00000100; //  805 :   4 - 0x4
      13'h326: dout  = 8'b00000010; //  806 :   2 - 0x2
      13'h327: dout  = 8'b00000010; //  807 :   2 - 0x2
      13'h328: dout  = 8'b00000000; //  808 :   0 - 0x0
      13'h329: dout  = 8'b00000000; //  809 :   0 - 0x0
      13'h32A: dout  = 8'b00000000; //  810 :   0 - 0x0
      13'h32B: dout  = 8'b11100000; //  811 : 224 - 0xe0
      13'h32C: dout  = 8'b00010000; //  812 :  16 - 0x10
      13'h32D: dout  = 8'b00001000; //  813 :   8 - 0x8
      13'h32E: dout  = 8'b00000100; //  814 :   4 - 0x4
      13'h32F: dout  = 8'b00000100; //  815 :   4 - 0x4
      13'h330: dout  = 8'b00000010; //  816 :   2 - 0x2 -- Sprite 0x33
      13'h331: dout  = 8'b00000010; //  817 :   2 - 0x2
      13'h332: dout  = 8'b00000100; //  818 :   4 - 0x4
      13'h333: dout  = 8'b00001000; //  819 :   8 - 0x8
      13'h334: dout  = 8'b00010000; //  820 :  16 - 0x10
      13'h335: dout  = 8'b11100000; //  821 : 224 - 0xe0
      13'h336: dout  = 8'b00000000; //  822 :   0 - 0x0
      13'h337: dout  = 8'b00000000; //  823 :   0 - 0x0
      13'h338: dout  = 8'b00000100; //  824 :   4 - 0x4
      13'h339: dout  = 8'b00000100; //  825 :   4 - 0x4
      13'h33A: dout  = 8'b00001000; //  826 :   8 - 0x8
      13'h33B: dout  = 8'b00010000; //  827 :  16 - 0x10
      13'h33C: dout  = 8'b11100000; //  828 : 224 - 0xe0
      13'h33D: dout  = 8'b00000000; //  829 :   0 - 0x0
      13'h33E: dout  = 8'b00000000; //  830 :   0 - 0x0
      13'h33F: dout  = 8'b00000000; //  831 :   0 - 0x0
      13'h340: dout  = 8'b00000000; //  832 :   0 - 0x0 -- Sprite 0x34
      13'h341: dout  = 8'b00000000; //  833 :   0 - 0x0
      13'h342: dout  = 8'b00000000; //  834 :   0 - 0x0
      13'h343: dout  = 8'b00000000; //  835 :   0 - 0x0
      13'h344: dout  = 8'b00000011; //  836 :   3 - 0x3
      13'h345: dout  = 8'b00000100; //  837 :   4 - 0x4
      13'h346: dout  = 8'b00001000; //  838 :   8 - 0x8
      13'h347: dout  = 8'b00010000; //  839 :  16 - 0x10
      13'h348: dout  = 8'b00000000; //  840 :   0 - 0x0
      13'h349: dout  = 8'b00000000; //  841 :   0 - 0x0
      13'h34A: dout  = 8'b00000000; //  842 :   0 - 0x0
      13'h34B: dout  = 8'b00000000; //  843 :   0 - 0x0
      13'h34C: dout  = 8'b00000000; //  844 :   0 - 0x0
      13'h34D: dout  = 8'b00000011; //  845 :   3 - 0x3
      13'h34E: dout  = 8'b00000100; //  846 :   4 - 0x4
      13'h34F: dout  = 8'b00001000; //  847 :   8 - 0x8
      13'h350: dout  = 8'b00010000; //  848 :  16 - 0x10 -- Sprite 0x35
      13'h351: dout  = 8'b00001000; //  849 :   8 - 0x8
      13'h352: dout  = 8'b00000100; //  850 :   4 - 0x4
      13'h353: dout  = 8'b00000011; //  851 :   3 - 0x3
      13'h354: dout  = 8'b00000000; //  852 :   0 - 0x0
      13'h355: dout  = 8'b00000000; //  853 :   0 - 0x0
      13'h356: dout  = 8'b00000000; //  854 :   0 - 0x0
      13'h357: dout  = 8'b00000000; //  855 :   0 - 0x0
      13'h358: dout  = 8'b00001000; //  856 :   8 - 0x8
      13'h359: dout  = 8'b00000100; //  857 :   4 - 0x4
      13'h35A: dout  = 8'b00000011; //  858 :   3 - 0x3
      13'h35B: dout  = 8'b00000000; //  859 :   0 - 0x0
      13'h35C: dout  = 8'b00000000; //  860 :   0 - 0x0
      13'h35D: dout  = 8'b00000000; //  861 :   0 - 0x0
      13'h35E: dout  = 8'b00000000; //  862 :   0 - 0x0
      13'h35F: dout  = 8'b00000000; //  863 :   0 - 0x0
      13'h360: dout  = 8'b00000000; //  864 :   0 - 0x0 -- Sprite 0x36
      13'h361: dout  = 8'b00000000; //  865 :   0 - 0x0
      13'h362: dout  = 8'b00000000; //  866 :   0 - 0x0
      13'h363: dout  = 8'b00000000; //  867 :   0 - 0x0
      13'h364: dout  = 8'b11000000; //  868 : 192 - 0xc0
      13'h365: dout  = 8'b00100000; //  869 :  32 - 0x20
      13'h366: dout  = 8'b00010000; //  870 :  16 - 0x10
      13'h367: dout  = 8'b00001000; //  871 :   8 - 0x8
      13'h368: dout  = 8'b00000000; //  872 :   0 - 0x0
      13'h369: dout  = 8'b00000000; //  873 :   0 - 0x0
      13'h36A: dout  = 8'b00000000; //  874 :   0 - 0x0
      13'h36B: dout  = 8'b00000000; //  875 :   0 - 0x0
      13'h36C: dout  = 8'b00000000; //  876 :   0 - 0x0
      13'h36D: dout  = 8'b11000000; //  877 : 192 - 0xc0
      13'h36E: dout  = 8'b00100000; //  878 :  32 - 0x20
      13'h36F: dout  = 8'b00010000; //  879 :  16 - 0x10
      13'h370: dout  = 8'b00001000; //  880 :   8 - 0x8 -- Sprite 0x37
      13'h371: dout  = 8'b00010000; //  881 :  16 - 0x10
      13'h372: dout  = 8'b00100000; //  882 :  32 - 0x20
      13'h373: dout  = 8'b11000000; //  883 : 192 - 0xc0
      13'h374: dout  = 8'b00000000; //  884 :   0 - 0x0
      13'h375: dout  = 8'b00000000; //  885 :   0 - 0x0
      13'h376: dout  = 8'b00000000; //  886 :   0 - 0x0
      13'h377: dout  = 8'b00000000; //  887 :   0 - 0x0
      13'h378: dout  = 8'b00010000; //  888 :  16 - 0x10
      13'h379: dout  = 8'b00100000; //  889 :  32 - 0x20
      13'h37A: dout  = 8'b11000000; //  890 : 192 - 0xc0
      13'h37B: dout  = 8'b00000000; //  891 :   0 - 0x0
      13'h37C: dout  = 8'b00000000; //  892 :   0 - 0x0
      13'h37D: dout  = 8'b00000000; //  893 :   0 - 0x0
      13'h37E: dout  = 8'b00000000; //  894 :   0 - 0x0
      13'h37F: dout  = 8'b00000000; //  895 :   0 - 0x0
      13'h380: dout  = 8'b00000000; //  896 :   0 - 0x0 -- Sprite 0x38
      13'h381: dout  = 8'b00000000; //  897 :   0 - 0x0
      13'h382: dout  = 8'b00000000; //  898 :   0 - 0x0
      13'h383: dout  = 8'b00000000; //  899 :   0 - 0x0
      13'h384: dout  = 8'b00000000; //  900 :   0 - 0x0
      13'h385: dout  = 8'b00000000; //  901 :   0 - 0x0
      13'h386: dout  = 8'b00000000; //  902 :   0 - 0x0
      13'h387: dout  = 8'b00000001; //  903 :   1 - 0x1
      13'h388: dout  = 8'b00000000; //  904 :   0 - 0x0
      13'h389: dout  = 8'b00000000; //  905 :   0 - 0x0
      13'h38A: dout  = 8'b00000000; //  906 :   0 - 0x0
      13'h38B: dout  = 8'b00000000; //  907 :   0 - 0x0
      13'h38C: dout  = 8'b00000000; //  908 :   0 - 0x0
      13'h38D: dout  = 8'b00000000; //  909 :   0 - 0x0
      13'h38E: dout  = 8'b00000000; //  910 :   0 - 0x0
      13'h38F: dout  = 8'b00000000; //  911 :   0 - 0x0
      13'h390: dout  = 8'b00000010; //  912 :   2 - 0x2 -- Sprite 0x39
      13'h391: dout  = 8'b00000001; //  913 :   1 - 0x1
      13'h392: dout  = 8'b00000000; //  914 :   0 - 0x0
      13'h393: dout  = 8'b00000000; //  915 :   0 - 0x0
      13'h394: dout  = 8'b00000000; //  916 :   0 - 0x0
      13'h395: dout  = 8'b00000000; //  917 :   0 - 0x0
      13'h396: dout  = 8'b00000000; //  918 :   0 - 0x0
      13'h397: dout  = 8'b00000000; //  919 :   0 - 0x0
      13'h398: dout  = 8'b00000001; //  920 :   1 - 0x1
      13'h399: dout  = 8'b00000000; //  921 :   0 - 0x0
      13'h39A: dout  = 8'b00000000; //  922 :   0 - 0x0
      13'h39B: dout  = 8'b00000000; //  923 :   0 - 0x0
      13'h39C: dout  = 8'b00000000; //  924 :   0 - 0x0
      13'h39D: dout  = 8'b00000000; //  925 :   0 - 0x0
      13'h39E: dout  = 8'b00000000; //  926 :   0 - 0x0
      13'h39F: dout  = 8'b00000000; //  927 :   0 - 0x0
      13'h3A0: dout  = 8'b00000000; //  928 :   0 - 0x0 -- Sprite 0x3a
      13'h3A1: dout  = 8'b00000000; //  929 :   0 - 0x0
      13'h3A2: dout  = 8'b00000000; //  930 :   0 - 0x0
      13'h3A3: dout  = 8'b00000000; //  931 :   0 - 0x0
      13'h3A4: dout  = 8'b00000000; //  932 :   0 - 0x0
      13'h3A5: dout  = 8'b00000000; //  933 :   0 - 0x0
      13'h3A6: dout  = 8'b00000000; //  934 :   0 - 0x0
      13'h3A7: dout  = 8'b00000000; //  935 :   0 - 0x0
      13'h3A8: dout  = 8'b00000000; //  936 :   0 - 0x0
      13'h3A9: dout  = 8'b00000000; //  937 :   0 - 0x0
      13'h3AA: dout  = 8'b00000000; //  938 :   0 - 0x0
      13'h3AB: dout  = 8'b00000000; //  939 :   0 - 0x0
      13'h3AC: dout  = 8'b00000000; //  940 :   0 - 0x0
      13'h3AD: dout  = 8'b00000000; //  941 :   0 - 0x0
      13'h3AE: dout  = 8'b00000000; //  942 :   0 - 0x0
      13'h3AF: dout  = 8'b00000000; //  943 :   0 - 0x0
      13'h3B0: dout  = 8'b10000000; //  944 : 128 - 0x80 -- Sprite 0x3b
      13'h3B1: dout  = 8'b00000000; //  945 :   0 - 0x0
      13'h3B2: dout  = 8'b00000000; //  946 :   0 - 0x0
      13'h3B3: dout  = 8'b00000000; //  947 :   0 - 0x0
      13'h3B4: dout  = 8'b00000000; //  948 :   0 - 0x0
      13'h3B5: dout  = 8'b00000000; //  949 :   0 - 0x0
      13'h3B6: dout  = 8'b00000000; //  950 :   0 - 0x0
      13'h3B7: dout  = 8'b00000000; //  951 :   0 - 0x0
      13'h3B8: dout  = 8'b00000000; //  952 :   0 - 0x0
      13'h3B9: dout  = 8'b00000000; //  953 :   0 - 0x0
      13'h3BA: dout  = 8'b00000000; //  954 :   0 - 0x0
      13'h3BB: dout  = 8'b00000000; //  955 :   0 - 0x0
      13'h3BC: dout  = 8'b00000000; //  956 :   0 - 0x0
      13'h3BD: dout  = 8'b00000000; //  957 :   0 - 0x0
      13'h3BE: dout  = 8'b00000000; //  958 :   0 - 0x0
      13'h3BF: dout  = 8'b00000000; //  959 :   0 - 0x0
      13'h3C0: dout  = 8'b00000000; //  960 :   0 - 0x0 -- Sprite 0x3c
      13'h3C1: dout  = 8'b00000000; //  961 :   0 - 0x0
      13'h3C2: dout  = 8'b00000000; //  962 :   0 - 0x0
      13'h3C3: dout  = 8'b00000001; //  963 :   1 - 0x1
      13'h3C4: dout  = 8'b00100001; //  964 :  33 - 0x21
      13'h3C5: dout  = 8'b00010000; //  965 :  16 - 0x10
      13'h3C6: dout  = 8'b00000000; //  966 :   0 - 0x0
      13'h3C7: dout  = 8'b00000000; //  967 :   0 - 0x0
      13'h3C8: dout  = 8'b00000000; //  968 :   0 - 0x0
      13'h3C9: dout  = 8'b00000001; //  969 :   1 - 0x1
      13'h3CA: dout  = 8'b00000001; //  970 :   1 - 0x1
      13'h3CB: dout  = 8'b01000000; //  971 :  64 - 0x40
      13'h3CC: dout  = 8'b00000000; //  972 :   0 - 0x0
      13'h3CD: dout  = 8'b00000000; //  973 :   0 - 0x0
      13'h3CE: dout  = 8'b00000000; //  974 :   0 - 0x0
      13'h3CF: dout  = 8'b00000000; //  975 :   0 - 0x0
      13'h3D0: dout  = 8'b01100000; //  976 :  96 - 0x60 -- Sprite 0x3d
      13'h3D1: dout  = 8'b00000000; //  977 :   0 - 0x0
      13'h3D2: dout  = 8'b00000000; //  978 :   0 - 0x0
      13'h3D3: dout  = 8'b00010000; //  979 :  16 - 0x10
      13'h3D4: dout  = 8'b00100001; //  980 :  33 - 0x21
      13'h3D5: dout  = 8'b00000001; //  981 :   1 - 0x1
      13'h3D6: dout  = 8'b00000000; //  982 :   0 - 0x0
      13'h3D7: dout  = 8'b00000000; //  983 :   0 - 0x0
      13'h3D8: dout  = 8'b10000000; //  984 : 128 - 0x80
      13'h3D9: dout  = 8'b00000000; //  985 :   0 - 0x0
      13'h3DA: dout  = 8'b00000000; //  986 :   0 - 0x0
      13'h3DB: dout  = 8'b00000000; //  987 :   0 - 0x0
      13'h3DC: dout  = 8'b00000000; //  988 :   0 - 0x0
      13'h3DD: dout  = 8'b01000000; //  989 :  64 - 0x40
      13'h3DE: dout  = 8'b00000001; //  990 :   1 - 0x1
      13'h3DF: dout  = 8'b00000001; //  991 :   1 - 0x1
      13'h3E0: dout  = 8'b00000000; //  992 :   0 - 0x0 -- Sprite 0x3e
      13'h3E1: dout  = 8'b00000000; //  993 :   0 - 0x0
      13'h3E2: dout  = 8'b00000000; //  994 :   0 - 0x0
      13'h3E3: dout  = 8'b00000000; //  995 :   0 - 0x0
      13'h3E4: dout  = 8'b00001000; //  996 :   8 - 0x8
      13'h3E5: dout  = 8'b00010000; //  997 :  16 - 0x10
      13'h3E6: dout  = 8'b00000000; //  998 :   0 - 0x0
      13'h3E7: dout  = 8'b00000000; //  999 :   0 - 0x0
      13'h3E8: dout  = 8'b00000000; // 1000 :   0 - 0x0
      13'h3E9: dout  = 8'b00000000; // 1001 :   0 - 0x0
      13'h3EA: dout  = 8'b00000000; // 1002 :   0 - 0x0
      13'h3EB: dout  = 8'b00000100; // 1003 :   4 - 0x4
      13'h3EC: dout  = 8'b00000000; // 1004 :   0 - 0x0
      13'h3ED: dout  = 8'b00000000; // 1005 :   0 - 0x0
      13'h3EE: dout  = 8'b00000000; // 1006 :   0 - 0x0
      13'h3EF: dout  = 8'b00000000; // 1007 :   0 - 0x0
      13'h3F0: dout  = 8'b00001100; // 1008 :  12 - 0xc -- Sprite 0x3f
      13'h3F1: dout  = 8'b00000000; // 1009 :   0 - 0x0
      13'h3F2: dout  = 8'b00000000; // 1010 :   0 - 0x0
      13'h3F3: dout  = 8'b00010000; // 1011 :  16 - 0x10
      13'h3F4: dout  = 8'b00001000; // 1012 :   8 - 0x8
      13'h3F5: dout  = 8'b00000000; // 1013 :   0 - 0x0
      13'h3F6: dout  = 8'b00000000; // 1014 :   0 - 0x0
      13'h3F7: dout  = 8'b00000000; // 1015 :   0 - 0x0
      13'h3F8: dout  = 8'b00000010; // 1016 :   2 - 0x2
      13'h3F9: dout  = 8'b00000000; // 1017 :   0 - 0x0
      13'h3FA: dout  = 8'b00000000; // 1018 :   0 - 0x0
      13'h3FB: dout  = 8'b00000000; // 1019 :   0 - 0x0
      13'h3FC: dout  = 8'b00000000; // 1020 :   0 - 0x0
      13'h3FD: dout  = 8'b00000100; // 1021 :   4 - 0x4
      13'h3FE: dout  = 8'b00000000; // 1022 :   0 - 0x0
      13'h3FF: dout  = 8'b00000000; // 1023 :   0 - 0x0
      13'h400: dout  = 8'b00000100; // 1024 :   4 - 0x4 -- Sprite 0x40
      13'h401: dout  = 8'b00000010; // 1025 :   2 - 0x2
      13'h402: dout  = 8'b00000001; // 1026 :   1 - 0x1
      13'h403: dout  = 8'b00000000; // 1027 :   0 - 0x0
      13'h404: dout  = 8'b00000000; // 1028 :   0 - 0x0
      13'h405: dout  = 8'b00000000; // 1029 :   0 - 0x0
      13'h406: dout  = 8'b00000000; // 1030 :   0 - 0x0
      13'h407: dout  = 8'b00000000; // 1031 :   0 - 0x0
      13'h408: dout  = 8'b00001111; // 1032 :  15 - 0xf
      13'h409: dout  = 8'b00000111; // 1033 :   7 - 0x7
      13'h40A: dout  = 8'b00000011; // 1034 :   3 - 0x3
      13'h40B: dout  = 8'b00000000; // 1035 :   0 - 0x0
      13'h40C: dout  = 8'b00000000; // 1036 :   0 - 0x0
      13'h40D: dout  = 8'b00000001; // 1037 :   1 - 0x1
      13'h40E: dout  = 8'b00000001; // 1038 :   1 - 0x1
      13'h40F: dout  = 8'b00000001; // 1039 :   1 - 0x1
      13'h410: dout  = 8'b00000000; // 1040 :   0 - 0x0 -- Sprite 0x41
      13'h411: dout  = 8'b00000000; // 1041 :   0 - 0x0
      13'h412: dout  = 8'b00000000; // 1042 :   0 - 0x0
      13'h413: dout  = 8'b00000000; // 1043 :   0 - 0x0
      13'h414: dout  = 8'b00000000; // 1044 :   0 - 0x0
      13'h415: dout  = 8'b00000000; // 1045 :   0 - 0x0
      13'h416: dout  = 8'b00000001; // 1046 :   1 - 0x1
      13'h417: dout  = 8'b00000011; // 1047 :   3 - 0x3
      13'h418: dout  = 8'b00000000; // 1048 :   0 - 0x0
      13'h419: dout  = 8'b00000000; // 1049 :   0 - 0x0
      13'h41A: dout  = 8'b00000000; // 1050 :   0 - 0x0
      13'h41B: dout  = 8'b00000000; // 1051 :   0 - 0x0
      13'h41C: dout  = 8'b00000000; // 1052 :   0 - 0x0
      13'h41D: dout  = 8'b00000000; // 1053 :   0 - 0x0
      13'h41E: dout  = 8'b00000001; // 1054 :   1 - 0x1
      13'h41F: dout  = 8'b00000011; // 1055 :   3 - 0x3
      13'h420: dout  = 8'b00000111; // 1056 :   7 - 0x7 -- Sprite 0x42
      13'h421: dout  = 8'b00000111; // 1057 :   7 - 0x7
      13'h422: dout  = 8'b00000111; // 1058 :   7 - 0x7
      13'h423: dout  = 8'b00000011; // 1059 :   3 - 0x3
      13'h424: dout  = 8'b00000001; // 1060 :   1 - 0x1
      13'h425: dout  = 8'b00000000; // 1061 :   0 - 0x0
      13'h426: dout  = 8'b00000000; // 1062 :   0 - 0x0
      13'h427: dout  = 8'b00000000; // 1063 :   0 - 0x0
      13'h428: dout  = 8'b00000111; // 1064 :   7 - 0x7
      13'h429: dout  = 8'b00000111; // 1065 :   7 - 0x7
      13'h42A: dout  = 8'b00000111; // 1066 :   7 - 0x7
      13'h42B: dout  = 8'b00000111; // 1067 :   7 - 0x7
      13'h42C: dout  = 8'b00000011; // 1068 :   3 - 0x3
      13'h42D: dout  = 8'b00000001; // 1069 :   1 - 0x1
      13'h42E: dout  = 8'b00000000; // 1070 :   0 - 0x0
      13'h42F: dout  = 8'b00000000; // 1071 :   0 - 0x0
      13'h430: dout  = 8'b00000000; // 1072 :   0 - 0x0 -- Sprite 0x43
      13'h431: dout  = 8'b00000000; // 1073 :   0 - 0x0
      13'h432: dout  = 8'b00000000; // 1074 :   0 - 0x0
      13'h433: dout  = 8'b00000000; // 1075 :   0 - 0x0
      13'h434: dout  = 8'b00000000; // 1076 :   0 - 0x0
      13'h435: dout  = 8'b00000000; // 1077 :   0 - 0x0
      13'h436: dout  = 8'b00000000; // 1078 :   0 - 0x0
      13'h437: dout  = 8'b00000000; // 1079 :   0 - 0x0
      13'h438: dout  = 8'b00000000; // 1080 :   0 - 0x0
      13'h439: dout  = 8'b00000000; // 1081 :   0 - 0x0
      13'h43A: dout  = 8'b00000000; // 1082 :   0 - 0x0
      13'h43B: dout  = 8'b00000000; // 1083 :   0 - 0x0
      13'h43C: dout  = 8'b00000000; // 1084 :   0 - 0x0
      13'h43D: dout  = 8'b00000000; // 1085 :   0 - 0x0
      13'h43E: dout  = 8'b00000000; // 1086 :   0 - 0x0
      13'h43F: dout  = 8'b00000000; // 1087 :   0 - 0x0
      13'h440: dout  = 8'b00000000; // 1088 :   0 - 0x0 -- Sprite 0x44
      13'h441: dout  = 8'b01000010; // 1089 :  66 - 0x42
      13'h442: dout  = 8'b00111001; // 1090 :  57 - 0x39
      13'h443: dout  = 8'b11111111; // 1091 : 255 - 0xff
      13'h444: dout  = 8'b11111111; // 1092 : 255 - 0xff
      13'h445: dout  = 8'b11111111; // 1093 : 255 - 0xff
      13'h446: dout  = 8'b11111111; // 1094 : 255 - 0xff
      13'h447: dout  = 8'b11111111; // 1095 : 255 - 0xff
      13'h448: dout  = 8'b11111111; // 1096 : 255 - 0xff
      13'h449: dout  = 8'b11111111; // 1097 : 255 - 0xff
      13'h44A: dout  = 8'b11111111; // 1098 : 255 - 0xff
      13'h44B: dout  = 8'b11111111; // 1099 : 255 - 0xff
      13'h44C: dout  = 8'b11111111; // 1100 : 255 - 0xff
      13'h44D: dout  = 8'b11111111; // 1101 : 255 - 0xff
      13'h44E: dout  = 8'b11111111; // 1102 : 255 - 0xff
      13'h44F: dout  = 8'b11111111; // 1103 : 255 - 0xff
      13'h450: dout  = 8'b01111111; // 1104 : 127 - 0x7f -- Sprite 0x45
      13'h451: dout  = 8'b00111111; // 1105 :  63 - 0x3f
      13'h452: dout  = 8'b00011111; // 1106 :  31 - 0x1f
      13'h453: dout  = 8'b00001111; // 1107 :  15 - 0xf
      13'h454: dout  = 8'b00011111; // 1108 :  31 - 0x1f
      13'h455: dout  = 8'b11111111; // 1109 : 255 - 0xff
      13'h456: dout  = 8'b11111111; // 1110 : 255 - 0xff
      13'h457: dout  = 8'b11111111; // 1111 : 255 - 0xff
      13'h458: dout  = 8'b11111111; // 1112 : 255 - 0xff
      13'h459: dout  = 8'b01111111; // 1113 : 127 - 0x7f
      13'h45A: dout  = 8'b00111111; // 1114 :  63 - 0x3f
      13'h45B: dout  = 8'b00011111; // 1115 :  31 - 0x1f
      13'h45C: dout  = 8'b00011111; // 1116 :  31 - 0x1f
      13'h45D: dout  = 8'b11111111; // 1117 : 255 - 0xff
      13'h45E: dout  = 8'b11111111; // 1118 : 255 - 0xff
      13'h45F: dout  = 8'b11111111; // 1119 : 255 - 0xff
      13'h460: dout  = 8'b11111000; // 1120 : 248 - 0xf8 -- Sprite 0x46
      13'h461: dout  = 8'b11110111; // 1121 : 247 - 0xf7
      13'h462: dout  = 8'b11101111; // 1122 : 239 - 0xef
      13'h463: dout  = 8'b11111111; // 1123 : 255 - 0xff
      13'h464: dout  = 8'b11111111; // 1124 : 255 - 0xff
      13'h465: dout  = 8'b11111110; // 1125 : 254 - 0xfe
      13'h466: dout  = 8'b01111110; // 1126 : 126 - 0x7e
      13'h467: dout  = 8'b00111110; // 1127 :  62 - 0x3e
      13'h468: dout  = 8'b11111111; // 1128 : 255 - 0xff
      13'h469: dout  = 8'b11111111; // 1129 : 255 - 0xff
      13'h46A: dout  = 8'b11111111; // 1130 : 255 - 0xff
      13'h46B: dout  = 8'b11111111; // 1131 : 255 - 0xff
      13'h46C: dout  = 8'b11111111; // 1132 : 255 - 0xff
      13'h46D: dout  = 8'b11111111; // 1133 : 255 - 0xff
      13'h46E: dout  = 8'b11111111; // 1134 : 255 - 0xff
      13'h46F: dout  = 8'b01111111; // 1135 : 127 - 0x7f
      13'h470: dout  = 8'b00000111; // 1136 :   7 - 0x7 -- Sprite 0x47
      13'h471: dout  = 8'b00000000; // 1137 :   0 - 0x0
      13'h472: dout  = 8'b00000000; // 1138 :   0 - 0x0
      13'h473: dout  = 8'b00000000; // 1139 :   0 - 0x0
      13'h474: dout  = 8'b00000000; // 1140 :   0 - 0x0
      13'h475: dout  = 8'b00000000; // 1141 :   0 - 0x0
      13'h476: dout  = 8'b00000000; // 1142 :   0 - 0x0
      13'h477: dout  = 8'b00000000; // 1143 :   0 - 0x0
      13'h478: dout  = 8'b00000111; // 1144 :   7 - 0x7
      13'h479: dout  = 8'b00000011; // 1145 :   3 - 0x3
      13'h47A: dout  = 8'b00000011; // 1146 :   3 - 0x3
      13'h47B: dout  = 8'b00000001; // 1147 :   1 - 0x1
      13'h47C: dout  = 8'b00000000; // 1148 :   0 - 0x0
      13'h47D: dout  = 8'b00000000; // 1149 :   0 - 0x0
      13'h47E: dout  = 8'b00000000; // 1150 :   0 - 0x0
      13'h47F: dout  = 8'b00000000; // 1151 :   0 - 0x0
      13'h480: dout  = 8'b00000000; // 1152 :   0 - 0x0 -- Sprite 0x48
      13'h481: dout  = 8'b00000000; // 1153 :   0 - 0x0
      13'h482: dout  = 8'b00000000; // 1154 :   0 - 0x0
      13'h483: dout  = 8'b11000000; // 1155 : 192 - 0xc0
      13'h484: dout  = 8'b11100000; // 1156 : 224 - 0xe0
      13'h485: dout  = 8'b11110000; // 1157 : 240 - 0xf0
      13'h486: dout  = 8'b11011011; // 1158 : 219 - 0xdb
      13'h487: dout  = 8'b11110110; // 1159 : 246 - 0xf6
      13'h488: dout  = 8'b00000000; // 1160 :   0 - 0x0
      13'h489: dout  = 8'b10000000; // 1161 : 128 - 0x80
      13'h48A: dout  = 8'b10000000; // 1162 : 128 - 0x80
      13'h48B: dout  = 8'b11000000; // 1163 : 192 - 0xc0
      13'h48C: dout  = 8'b11100000; // 1164 : 224 - 0xe0
      13'h48D: dout  = 8'b11110000; // 1165 : 240 - 0xf0
      13'h48E: dout  = 8'b11111111; // 1166 : 255 - 0xff
      13'h48F: dout  = 8'b11111111; // 1167 : 255 - 0xff
      13'h490: dout  = 8'b11001011; // 1168 : 203 - 0xcb -- Sprite 0x49
      13'h491: dout  = 8'b11100000; // 1169 : 224 - 0xe0
      13'h492: dout  = 8'b11000100; // 1170 : 196 - 0xc4
      13'h493: dout  = 8'b00000010; // 1171 :   2 - 0x2
      13'h494: dout  = 8'b11010001; // 1172 : 209 - 0xd1
      13'h495: dout  = 8'b11100001; // 1173 : 225 - 0xe1
      13'h496: dout  = 8'b11010001; // 1174 : 209 - 0xd1
      13'h497: dout  = 8'b10000011; // 1175 : 131 - 0x83
      13'h498: dout  = 8'b11111111; // 1176 : 255 - 0xff
      13'h499: dout  = 8'b11111111; // 1177 : 255 - 0xff
      13'h49A: dout  = 8'b11111111; // 1178 : 255 - 0xff
      13'h49B: dout  = 8'b11111111; // 1179 : 255 - 0xff
      13'h49C: dout  = 8'b11111111; // 1180 : 255 - 0xff
      13'h49D: dout  = 8'b11111111; // 1181 : 255 - 0xff
      13'h49E: dout  = 8'b11111111; // 1182 : 255 - 0xff
      13'h49F: dout  = 8'b11111111; // 1183 : 255 - 0xff
      13'h4A0: dout  = 8'b00001111; // 1184 :  15 - 0xf -- Sprite 0x4a
      13'h4A1: dout  = 8'b11111111; // 1185 : 255 - 0xff
      13'h4A2: dout  = 8'b11100000; // 1186 : 224 - 0xe0
      13'h4A3: dout  = 8'b10001111; // 1187 : 143 - 0x8f
      13'h4A4: dout  = 8'b01101110; // 1188 : 110 - 0x6e
      13'h4A5: dout  = 8'b01000100; // 1189 :  68 - 0x44
      13'h4A6: dout  = 8'b11101110; // 1190 : 238 - 0xee
      13'h4A7: dout  = 8'b01100000; // 1191 :  96 - 0x60
      13'h4A8: dout  = 8'b11111111; // 1192 : 255 - 0xff
      13'h4A9: dout  = 8'b11111111; // 1193 : 255 - 0xff
      13'h4AA: dout  = 8'b11111111; // 1194 : 255 - 0xff
      13'h4AB: dout  = 8'b11110000; // 1195 : 240 - 0xf0
      13'h4AC: dout  = 8'b10000000; // 1196 : 128 - 0x80
      13'h4AD: dout  = 8'b00000000; // 1197 :   0 - 0x0
      13'h4AE: dout  = 8'b00000000; // 1198 :   0 - 0x0
      13'h4AF: dout  = 8'b10011111; // 1199 : 159 - 0x9f
      13'h4B0: dout  = 8'b10000011; // 1200 : 131 - 0x83 -- Sprite 0x4b
      13'h4B1: dout  = 8'b11100000; // 1201 : 224 - 0xe0
      13'h4B2: dout  = 8'b11100100; // 1202 : 228 - 0xe4
      13'h4B3: dout  = 8'b11000110; // 1203 : 198 - 0xc6
      13'h4B4: dout  = 8'b01100001; // 1204 :  97 - 0x61
      13'h4B5: dout  = 8'b00110011; // 1205 :  51 - 0x33
      13'h4B6: dout  = 8'b00011111; // 1206 :  31 - 0x1f
      13'h4B7: dout  = 8'b00001111; // 1207 :  15 - 0xf
      13'h4B8: dout  = 8'b11111111; // 1208 : 255 - 0xff
      13'h4B9: dout  = 8'b11111111; // 1209 : 255 - 0xff
      13'h4BA: dout  = 8'b11111001; // 1210 : 249 - 0xf9
      13'h4BB: dout  = 8'b11111001; // 1211 : 249 - 0xf9
      13'h4BC: dout  = 8'b01111111; // 1212 : 127 - 0x7f
      13'h4BD: dout  = 8'b00111111; // 1213 :  63 - 0x3f
      13'h4BE: dout  = 8'b00011111; // 1214 :  31 - 0x1f
      13'h4BF: dout  = 8'b00001111; // 1215 :  15 - 0xf
      13'h4C0: dout  = 8'b00000000; // 1216 :   0 - 0x0 -- Sprite 0x4c
      13'h4C1: dout  = 8'b00000000; // 1217 :   0 - 0x0
      13'h4C2: dout  = 8'b00000000; // 1218 :   0 - 0x0
      13'h4C3: dout  = 8'b00000011; // 1219 :   3 - 0x3
      13'h4C4: dout  = 8'b00000111; // 1220 :   7 - 0x7
      13'h4C5: dout  = 8'b00001111; // 1221 :  15 - 0xf
      13'h4C6: dout  = 8'b01011011; // 1222 :  91 - 0x5b
      13'h4C7: dout  = 8'b10100111; // 1223 : 167 - 0xa7
      13'h4C8: dout  = 8'b00000000; // 1224 :   0 - 0x0
      13'h4C9: dout  = 8'b00000001; // 1225 :   1 - 0x1
      13'h4CA: dout  = 8'b00000001; // 1226 :   1 - 0x1
      13'h4CB: dout  = 8'b00000011; // 1227 :   3 - 0x3
      13'h4CC: dout  = 8'b00000111; // 1228 :   7 - 0x7
      13'h4CD: dout  = 8'b00001111; // 1229 :  15 - 0xf
      13'h4CE: dout  = 8'b11111111; // 1230 : 255 - 0xff
      13'h4CF: dout  = 8'b11111111; // 1231 : 255 - 0xff
      13'h4D0: dout  = 8'b01110011; // 1232 : 115 - 0x73 -- Sprite 0x4d
      13'h4D1: dout  = 8'b00000111; // 1233 :   7 - 0x7
      13'h4D2: dout  = 8'b00100111; // 1234 :  39 - 0x27
      13'h4D3: dout  = 8'b01000000; // 1235 :  64 - 0x40
      13'h4D4: dout  = 8'b10001011; // 1236 : 139 - 0x8b
      13'h4D5: dout  = 8'b10000111; // 1237 : 135 - 0x87
      13'h4D6: dout  = 8'b10001011; // 1238 : 139 - 0x8b
      13'h4D7: dout  = 8'b11000001; // 1239 : 193 - 0xc1
      13'h4D8: dout  = 8'b11111111; // 1240 : 255 - 0xff
      13'h4D9: dout  = 8'b11111111; // 1241 : 255 - 0xff
      13'h4DA: dout  = 8'b11111111; // 1242 : 255 - 0xff
      13'h4DB: dout  = 8'b11111111; // 1243 : 255 - 0xff
      13'h4DC: dout  = 8'b11111111; // 1244 : 255 - 0xff
      13'h4DD: dout  = 8'b11111111; // 1245 : 255 - 0xff
      13'h4DE: dout  = 8'b11111111; // 1246 : 255 - 0xff
      13'h4DF: dout  = 8'b11111111; // 1247 : 255 - 0xff
      13'h4E0: dout  = 8'b11110000; // 1248 : 240 - 0xf0 -- Sprite 0x4e
      13'h4E1: dout  = 8'b11111111; // 1249 : 255 - 0xff
      13'h4E2: dout  = 8'b00001111; // 1250 :  15 - 0xf
      13'h4E3: dout  = 8'b11100001; // 1251 : 225 - 0xe1
      13'h4E4: dout  = 8'b11101100; // 1252 : 236 - 0xec
      13'h4E5: dout  = 8'b01000100; // 1253 :  68 - 0x44
      13'h4E6: dout  = 8'b11101110; // 1254 : 238 - 0xee
      13'h4E7: dout  = 8'b00001100; // 1255 :  12 - 0xc
      13'h4E8: dout  = 8'b11111111; // 1256 : 255 - 0xff
      13'h4E9: dout  = 8'b11111111; // 1257 : 255 - 0xff
      13'h4EA: dout  = 8'b11111111; // 1258 : 255 - 0xff
      13'h4EB: dout  = 8'b00011111; // 1259 :  31 - 0x1f
      13'h4EC: dout  = 8'b00000011; // 1260 :   3 - 0x3
      13'h4ED: dout  = 8'b00000001; // 1261 :   1 - 0x1
      13'h4EE: dout  = 8'b00000001; // 1262 :   1 - 0x1
      13'h4EF: dout  = 8'b11110011; // 1263 : 243 - 0xf3
      13'h4F0: dout  = 8'b10000000; // 1264 : 128 - 0x80 -- Sprite 0x4f
      13'h4F1: dout  = 8'b00001110; // 1265 :  14 - 0xe
      13'h4F2: dout  = 8'b01001110; // 1266 :  78 - 0x4e
      13'h4F3: dout  = 8'b11000110; // 1267 : 198 - 0xc6
      13'h4F4: dout  = 8'b00001100; // 1268 :  12 - 0xc
      13'h4F5: dout  = 8'b10011000; // 1269 : 152 - 0x98
      13'h4F6: dout  = 8'b11110000; // 1270 : 240 - 0xf0
      13'h4F7: dout  = 8'b11100000; // 1271 : 224 - 0xe0
      13'h4F8: dout  = 8'b11111111; // 1272 : 255 - 0xff
      13'h4F9: dout  = 8'b11111111; // 1273 : 255 - 0xff
      13'h4FA: dout  = 8'b00111111; // 1274 :  63 - 0x3f
      13'h4FB: dout  = 8'b00111111; // 1275 :  63 - 0x3f
      13'h4FC: dout  = 8'b11111100; // 1276 : 252 - 0xfc
      13'h4FD: dout  = 8'b11111000; // 1277 : 248 - 0xf8
      13'h4FE: dout  = 8'b11110000; // 1278 : 240 - 0xf0
      13'h4FF: dout  = 8'b11100000; // 1279 : 224 - 0xe0
      13'h500: dout  = 8'b00000000; // 1280 :   0 - 0x0 -- Sprite 0x50
      13'h501: dout  = 8'b01000010; // 1281 :  66 - 0x42
      13'h502: dout  = 8'b10011100; // 1282 : 156 - 0x9c
      13'h503: dout  = 8'b11111111; // 1283 : 255 - 0xff
      13'h504: dout  = 8'b11111111; // 1284 : 255 - 0xff
      13'h505: dout  = 8'b11111111; // 1285 : 255 - 0xff
      13'h506: dout  = 8'b11111111; // 1286 : 255 - 0xff
      13'h507: dout  = 8'b11111111; // 1287 : 255 - 0xff
      13'h508: dout  = 8'b11111111; // 1288 : 255 - 0xff
      13'h509: dout  = 8'b11111111; // 1289 : 255 - 0xff
      13'h50A: dout  = 8'b11111111; // 1290 : 255 - 0xff
      13'h50B: dout  = 8'b11111111; // 1291 : 255 - 0xff
      13'h50C: dout  = 8'b11111111; // 1292 : 255 - 0xff
      13'h50D: dout  = 8'b11111111; // 1293 : 255 - 0xff
      13'h50E: dout  = 8'b11111111; // 1294 : 255 - 0xff
      13'h50F: dout  = 8'b11111111; // 1295 : 255 - 0xff
      13'h510: dout  = 8'b11111110; // 1296 : 254 - 0xfe -- Sprite 0x51
      13'h511: dout  = 8'b11111100; // 1297 : 252 - 0xfc
      13'h512: dout  = 8'b11111000; // 1298 : 248 - 0xf8
      13'h513: dout  = 8'b11110000; // 1299 : 240 - 0xf0
      13'h514: dout  = 8'b11111000; // 1300 : 248 - 0xf8
      13'h515: dout  = 8'b11111111; // 1301 : 255 - 0xff
      13'h516: dout  = 8'b11111111; // 1302 : 255 - 0xff
      13'h517: dout  = 8'b11111111; // 1303 : 255 - 0xff
      13'h518: dout  = 8'b11111111; // 1304 : 255 - 0xff
      13'h519: dout  = 8'b11111110; // 1305 : 254 - 0xfe
      13'h51A: dout  = 8'b11111100; // 1306 : 252 - 0xfc
      13'h51B: dout  = 8'b11111000; // 1307 : 248 - 0xf8
      13'h51C: dout  = 8'b11111000; // 1308 : 248 - 0xf8
      13'h51D: dout  = 8'b11111111; // 1309 : 255 - 0xff
      13'h51E: dout  = 8'b11111111; // 1310 : 255 - 0xff
      13'h51F: dout  = 8'b11111111; // 1311 : 255 - 0xff
      13'h520: dout  = 8'b00011111; // 1312 :  31 - 0x1f -- Sprite 0x52
      13'h521: dout  = 8'b11101111; // 1313 : 239 - 0xef
      13'h522: dout  = 8'b11110111; // 1314 : 247 - 0xf7
      13'h523: dout  = 8'b11111111; // 1315 : 255 - 0xff
      13'h524: dout  = 8'b11111111; // 1316 : 255 - 0xff
      13'h525: dout  = 8'b11111110; // 1317 : 254 - 0xfe
      13'h526: dout  = 8'b01111100; // 1318 : 124 - 0x7c
      13'h527: dout  = 8'b01110000; // 1319 : 112 - 0x70
      13'h528: dout  = 8'b11111111; // 1320 : 255 - 0xff
      13'h529: dout  = 8'b11111111; // 1321 : 255 - 0xff
      13'h52A: dout  = 8'b11111111; // 1322 : 255 - 0xff
      13'h52B: dout  = 8'b11111111; // 1323 : 255 - 0xff
      13'h52C: dout  = 8'b11111111; // 1324 : 255 - 0xff
      13'h52D: dout  = 8'b11111111; // 1325 : 255 - 0xff
      13'h52E: dout  = 8'b11111110; // 1326 : 254 - 0xfe
      13'h52F: dout  = 8'b11111100; // 1327 : 252 - 0xfc
      13'h530: dout  = 8'b11100000; // 1328 : 224 - 0xe0 -- Sprite 0x53
      13'h531: dout  = 8'b00000000; // 1329 :   0 - 0x0
      13'h532: dout  = 8'b00000000; // 1330 :   0 - 0x0
      13'h533: dout  = 8'b00000000; // 1331 :   0 - 0x0
      13'h534: dout  = 8'b00000000; // 1332 :   0 - 0x0
      13'h535: dout  = 8'b00000000; // 1333 :   0 - 0x0
      13'h536: dout  = 8'b00000000; // 1334 :   0 - 0x0
      13'h537: dout  = 8'b00000000; // 1335 :   0 - 0x0
      13'h538: dout  = 8'b11100000; // 1336 : 224 - 0xe0
      13'h539: dout  = 8'b10000000; // 1337 : 128 - 0x80
      13'h53A: dout  = 8'b10000000; // 1338 : 128 - 0x80
      13'h53B: dout  = 8'b00000000; // 1339 :   0 - 0x0
      13'h53C: dout  = 8'b00000000; // 1340 :   0 - 0x0
      13'h53D: dout  = 8'b00000000; // 1341 :   0 - 0x0
      13'h53E: dout  = 8'b00000000; // 1342 :   0 - 0x0
      13'h53F: dout  = 8'b00000000; // 1343 :   0 - 0x0
      13'h540: dout  = 8'b00100000; // 1344 :  32 - 0x20 -- Sprite 0x54
      13'h541: dout  = 8'b01000000; // 1345 :  64 - 0x40
      13'h542: dout  = 8'b10000000; // 1346 : 128 - 0x80
      13'h543: dout  = 8'b00000000; // 1347 :   0 - 0x0
      13'h544: dout  = 8'b00000000; // 1348 :   0 - 0x0
      13'h545: dout  = 8'b00000000; // 1349 :   0 - 0x0
      13'h546: dout  = 8'b00000000; // 1350 :   0 - 0x0
      13'h547: dout  = 8'b00000000; // 1351 :   0 - 0x0
      13'h548: dout  = 8'b11110000; // 1352 : 240 - 0xf0
      13'h549: dout  = 8'b11100000; // 1353 : 224 - 0xe0
      13'h54A: dout  = 8'b11000000; // 1354 : 192 - 0xc0
      13'h54B: dout  = 8'b00000000; // 1355 :   0 - 0x0
      13'h54C: dout  = 8'b00000000; // 1356 :   0 - 0x0
      13'h54D: dout  = 8'b10000000; // 1357 : 128 - 0x80
      13'h54E: dout  = 8'b10000000; // 1358 : 128 - 0x80
      13'h54F: dout  = 8'b10000000; // 1359 : 128 - 0x80
      13'h550: dout  = 8'b00000000; // 1360 :   0 - 0x0 -- Sprite 0x55
      13'h551: dout  = 8'b00000000; // 1361 :   0 - 0x0
      13'h552: dout  = 8'b00000000; // 1362 :   0 - 0x0
      13'h553: dout  = 8'b00000000; // 1363 :   0 - 0x0
      13'h554: dout  = 8'b00000000; // 1364 :   0 - 0x0
      13'h555: dout  = 8'b00000000; // 1365 :   0 - 0x0
      13'h556: dout  = 8'b10000000; // 1366 : 128 - 0x80
      13'h557: dout  = 8'b11000000; // 1367 : 192 - 0xc0
      13'h558: dout  = 8'b00000000; // 1368 :   0 - 0x0
      13'h559: dout  = 8'b00000000; // 1369 :   0 - 0x0
      13'h55A: dout  = 8'b00000000; // 1370 :   0 - 0x0
      13'h55B: dout  = 8'b00000000; // 1371 :   0 - 0x0
      13'h55C: dout  = 8'b00000000; // 1372 :   0 - 0x0
      13'h55D: dout  = 8'b00000000; // 1373 :   0 - 0x0
      13'h55E: dout  = 8'b10000000; // 1374 : 128 - 0x80
      13'h55F: dout  = 8'b11000000; // 1375 : 192 - 0xc0
      13'h560: dout  = 8'b11100000; // 1376 : 224 - 0xe0 -- Sprite 0x56
      13'h561: dout  = 8'b11100000; // 1377 : 224 - 0xe0
      13'h562: dout  = 8'b11100000; // 1378 : 224 - 0xe0
      13'h563: dout  = 8'b11000000; // 1379 : 192 - 0xc0
      13'h564: dout  = 8'b10000000; // 1380 : 128 - 0x80
      13'h565: dout  = 8'b00000000; // 1381 :   0 - 0x0
      13'h566: dout  = 8'b00000000; // 1382 :   0 - 0x0
      13'h567: dout  = 8'b00000000; // 1383 :   0 - 0x0
      13'h568: dout  = 8'b11100000; // 1384 : 224 - 0xe0
      13'h569: dout  = 8'b11100000; // 1385 : 224 - 0xe0
      13'h56A: dout  = 8'b11100000; // 1386 : 224 - 0xe0
      13'h56B: dout  = 8'b11100000; // 1387 : 224 - 0xe0
      13'h56C: dout  = 8'b11000000; // 1388 : 192 - 0xc0
      13'h56D: dout  = 8'b10000000; // 1389 : 128 - 0x80
      13'h56E: dout  = 8'b00000000; // 1390 :   0 - 0x0
      13'h56F: dout  = 8'b00000000; // 1391 :   0 - 0x0
      13'h570: dout  = 8'b00000000; // 1392 :   0 - 0x0 -- Sprite 0x57
      13'h571: dout  = 8'b00000000; // 1393 :   0 - 0x0
      13'h572: dout  = 8'b00000000; // 1394 :   0 - 0x0
      13'h573: dout  = 8'b00000000; // 1395 :   0 - 0x0
      13'h574: dout  = 8'b00000000; // 1396 :   0 - 0x0
      13'h575: dout  = 8'b00000000; // 1397 :   0 - 0x0
      13'h576: dout  = 8'b00000000; // 1398 :   0 - 0x0
      13'h577: dout  = 8'b00000000; // 1399 :   0 - 0x0
      13'h578: dout  = 8'b00000000; // 1400 :   0 - 0x0
      13'h579: dout  = 8'b00000000; // 1401 :   0 - 0x0
      13'h57A: dout  = 8'b00000000; // 1402 :   0 - 0x0
      13'h57B: dout  = 8'b00000000; // 1403 :   0 - 0x0
      13'h57C: dout  = 8'b00000000; // 1404 :   0 - 0x0
      13'h57D: dout  = 8'b00000000; // 1405 :   0 - 0x0
      13'h57E: dout  = 8'b00000000; // 1406 :   0 - 0x0
      13'h57F: dout  = 8'b00000000; // 1407 :   0 - 0x0
      13'h580: dout  = 8'b11111111; // 1408 : 255 - 0xff -- Sprite 0x58
      13'h581: dout  = 8'b11111111; // 1409 : 255 - 0xff
      13'h582: dout  = 8'b11111111; // 1410 : 255 - 0xff
      13'h583: dout  = 8'b11111111; // 1411 : 255 - 0xff
      13'h584: dout  = 8'b11111111; // 1412 : 255 - 0xff
      13'h585: dout  = 8'b11111111; // 1413 : 255 - 0xff
      13'h586: dout  = 8'b11111111; // 1414 : 255 - 0xff
      13'h587: dout  = 8'b11111111; // 1415 : 255 - 0xff
      13'h588: dout  = 8'b11111111; // 1416 : 255 - 0xff
      13'h589: dout  = 8'b11111111; // 1417 : 255 - 0xff
      13'h58A: dout  = 8'b11111111; // 1418 : 255 - 0xff
      13'h58B: dout  = 8'b11111111; // 1419 : 255 - 0xff
      13'h58C: dout  = 8'b11111111; // 1420 : 255 - 0xff
      13'h58D: dout  = 8'b11111111; // 1421 : 255 - 0xff
      13'h58E: dout  = 8'b11111111; // 1422 : 255 - 0xff
      13'h58F: dout  = 8'b11111111; // 1423 : 255 - 0xff
      13'h590: dout  = 8'b11111111; // 1424 : 255 - 0xff -- Sprite 0x59
      13'h591: dout  = 8'b11111111; // 1425 : 255 - 0xff
      13'h592: dout  = 8'b11111111; // 1426 : 255 - 0xff
      13'h593: dout  = 8'b11111111; // 1427 : 255 - 0xff
      13'h594: dout  = 8'b11111111; // 1428 : 255 - 0xff
      13'h595: dout  = 8'b11111111; // 1429 : 255 - 0xff
      13'h596: dout  = 8'b11111111; // 1430 : 255 - 0xff
      13'h597: dout  = 8'b11111111; // 1431 : 255 - 0xff
      13'h598: dout  = 8'b11111111; // 1432 : 255 - 0xff
      13'h599: dout  = 8'b11111111; // 1433 : 255 - 0xff
      13'h59A: dout  = 8'b11111111; // 1434 : 255 - 0xff
      13'h59B: dout  = 8'b11111111; // 1435 : 255 - 0xff
      13'h59C: dout  = 8'b11111111; // 1436 : 255 - 0xff
      13'h59D: dout  = 8'b11111111; // 1437 : 255 - 0xff
      13'h59E: dout  = 8'b11111111; // 1438 : 255 - 0xff
      13'h59F: dout  = 8'b11111111; // 1439 : 255 - 0xff
      13'h5A0: dout  = 8'b11111111; // 1440 : 255 - 0xff -- Sprite 0x5a
      13'h5A1: dout  = 8'b11111111; // 1441 : 255 - 0xff
      13'h5A2: dout  = 8'b11111111; // 1442 : 255 - 0xff
      13'h5A3: dout  = 8'b11111111; // 1443 : 255 - 0xff
      13'h5A4: dout  = 8'b11111111; // 1444 : 255 - 0xff
      13'h5A5: dout  = 8'b11111111; // 1445 : 255 - 0xff
      13'h5A6: dout  = 8'b11111111; // 1446 : 255 - 0xff
      13'h5A7: dout  = 8'b11111111; // 1447 : 255 - 0xff
      13'h5A8: dout  = 8'b11111111; // 1448 : 255 - 0xff
      13'h5A9: dout  = 8'b11111111; // 1449 : 255 - 0xff
      13'h5AA: dout  = 8'b11111111; // 1450 : 255 - 0xff
      13'h5AB: dout  = 8'b11111111; // 1451 : 255 - 0xff
      13'h5AC: dout  = 8'b11111111; // 1452 : 255 - 0xff
      13'h5AD: dout  = 8'b11111111; // 1453 : 255 - 0xff
      13'h5AE: dout  = 8'b11111111; // 1454 : 255 - 0xff
      13'h5AF: dout  = 8'b11111111; // 1455 : 255 - 0xff
      13'h5B0: dout  = 8'b11111111; // 1456 : 255 - 0xff -- Sprite 0x5b
      13'h5B1: dout  = 8'b11111111; // 1457 : 255 - 0xff
      13'h5B2: dout  = 8'b11111111; // 1458 : 255 - 0xff
      13'h5B3: dout  = 8'b11111111; // 1459 : 255 - 0xff
      13'h5B4: dout  = 8'b11111111; // 1460 : 255 - 0xff
      13'h5B5: dout  = 8'b11111111; // 1461 : 255 - 0xff
      13'h5B6: dout  = 8'b11111111; // 1462 : 255 - 0xff
      13'h5B7: dout  = 8'b11111111; // 1463 : 255 - 0xff
      13'h5B8: dout  = 8'b11111111; // 1464 : 255 - 0xff
      13'h5B9: dout  = 8'b11111111; // 1465 : 255 - 0xff
      13'h5BA: dout  = 8'b11111111; // 1466 : 255 - 0xff
      13'h5BB: dout  = 8'b11111111; // 1467 : 255 - 0xff
      13'h5BC: dout  = 8'b11111111; // 1468 : 255 - 0xff
      13'h5BD: dout  = 8'b11111111; // 1469 : 255 - 0xff
      13'h5BE: dout  = 8'b11111111; // 1470 : 255 - 0xff
      13'h5BF: dout  = 8'b11111111; // 1471 : 255 - 0xff
      13'h5C0: dout  = 8'b11111111; // 1472 : 255 - 0xff -- Sprite 0x5c
      13'h5C1: dout  = 8'b11111111; // 1473 : 255 - 0xff
      13'h5C2: dout  = 8'b11111111; // 1474 : 255 - 0xff
      13'h5C3: dout  = 8'b11111111; // 1475 : 255 - 0xff
      13'h5C4: dout  = 8'b11111111; // 1476 : 255 - 0xff
      13'h5C5: dout  = 8'b11111111; // 1477 : 255 - 0xff
      13'h5C6: dout  = 8'b11111111; // 1478 : 255 - 0xff
      13'h5C7: dout  = 8'b11111111; // 1479 : 255 - 0xff
      13'h5C8: dout  = 8'b11111111; // 1480 : 255 - 0xff
      13'h5C9: dout  = 8'b11111111; // 1481 : 255 - 0xff
      13'h5CA: dout  = 8'b11111111; // 1482 : 255 - 0xff
      13'h5CB: dout  = 8'b11111111; // 1483 : 255 - 0xff
      13'h5CC: dout  = 8'b11111111; // 1484 : 255 - 0xff
      13'h5CD: dout  = 8'b11111111; // 1485 : 255 - 0xff
      13'h5CE: dout  = 8'b11111111; // 1486 : 255 - 0xff
      13'h5CF: dout  = 8'b11111111; // 1487 : 255 - 0xff
      13'h5D0: dout  = 8'b11111111; // 1488 : 255 - 0xff -- Sprite 0x5d
      13'h5D1: dout  = 8'b11111111; // 1489 : 255 - 0xff
      13'h5D2: dout  = 8'b11111111; // 1490 : 255 - 0xff
      13'h5D3: dout  = 8'b11111111; // 1491 : 255 - 0xff
      13'h5D4: dout  = 8'b11111111; // 1492 : 255 - 0xff
      13'h5D5: dout  = 8'b11111111; // 1493 : 255 - 0xff
      13'h5D6: dout  = 8'b11111111; // 1494 : 255 - 0xff
      13'h5D7: dout  = 8'b11111111; // 1495 : 255 - 0xff
      13'h5D8: dout  = 8'b11111111; // 1496 : 255 - 0xff
      13'h5D9: dout  = 8'b11111111; // 1497 : 255 - 0xff
      13'h5DA: dout  = 8'b11111111; // 1498 : 255 - 0xff
      13'h5DB: dout  = 8'b11111111; // 1499 : 255 - 0xff
      13'h5DC: dout  = 8'b11111111; // 1500 : 255 - 0xff
      13'h5DD: dout  = 8'b11111111; // 1501 : 255 - 0xff
      13'h5DE: dout  = 8'b11111111; // 1502 : 255 - 0xff
      13'h5DF: dout  = 8'b11111111; // 1503 : 255 - 0xff
      13'h5E0: dout  = 8'b11111111; // 1504 : 255 - 0xff -- Sprite 0x5e
      13'h5E1: dout  = 8'b11111111; // 1505 : 255 - 0xff
      13'h5E2: dout  = 8'b11111111; // 1506 : 255 - 0xff
      13'h5E3: dout  = 8'b11111111; // 1507 : 255 - 0xff
      13'h5E4: dout  = 8'b11111111; // 1508 : 255 - 0xff
      13'h5E5: dout  = 8'b11111111; // 1509 : 255 - 0xff
      13'h5E6: dout  = 8'b11111111; // 1510 : 255 - 0xff
      13'h5E7: dout  = 8'b11111111; // 1511 : 255 - 0xff
      13'h5E8: dout  = 8'b11111111; // 1512 : 255 - 0xff
      13'h5E9: dout  = 8'b11111111; // 1513 : 255 - 0xff
      13'h5EA: dout  = 8'b11111111; // 1514 : 255 - 0xff
      13'h5EB: dout  = 8'b11111111; // 1515 : 255 - 0xff
      13'h5EC: dout  = 8'b11111111; // 1516 : 255 - 0xff
      13'h5ED: dout  = 8'b11111111; // 1517 : 255 - 0xff
      13'h5EE: dout  = 8'b11111111; // 1518 : 255 - 0xff
      13'h5EF: dout  = 8'b11111111; // 1519 : 255 - 0xff
      13'h5F0: dout  = 8'b11111111; // 1520 : 255 - 0xff -- Sprite 0x5f
      13'h5F1: dout  = 8'b11111111; // 1521 : 255 - 0xff
      13'h5F2: dout  = 8'b11111111; // 1522 : 255 - 0xff
      13'h5F3: dout  = 8'b11111111; // 1523 : 255 - 0xff
      13'h5F4: dout  = 8'b11111111; // 1524 : 255 - 0xff
      13'h5F5: dout  = 8'b11111111; // 1525 : 255 - 0xff
      13'h5F6: dout  = 8'b11111111; // 1526 : 255 - 0xff
      13'h5F7: dout  = 8'b11111111; // 1527 : 255 - 0xff
      13'h5F8: dout  = 8'b11111111; // 1528 : 255 - 0xff
      13'h5F9: dout  = 8'b11111111; // 1529 : 255 - 0xff
      13'h5FA: dout  = 8'b11111111; // 1530 : 255 - 0xff
      13'h5FB: dout  = 8'b11111111; // 1531 : 255 - 0xff
      13'h5FC: dout  = 8'b11111111; // 1532 : 255 - 0xff
      13'h5FD: dout  = 8'b11111111; // 1533 : 255 - 0xff
      13'h5FE: dout  = 8'b11111111; // 1534 : 255 - 0xff
      13'h5FF: dout  = 8'b11111111; // 1535 : 255 - 0xff
      13'h600: dout  = 8'b00000000; // 1536 :   0 - 0x0 -- Sprite 0x60
      13'h601: dout  = 8'b00000000; // 1537 :   0 - 0x0
      13'h602: dout  = 8'b00011111; // 1538 :  31 - 0x1f
      13'h603: dout  = 8'b00111111; // 1539 :  63 - 0x3f
      13'h604: dout  = 8'b00111111; // 1540 :  63 - 0x3f
      13'h605: dout  = 8'b01111111; // 1541 : 127 - 0x7f
      13'h606: dout  = 8'b01111111; // 1542 : 127 - 0x7f
      13'h607: dout  = 8'b01111111; // 1543 : 127 - 0x7f
      13'h608: dout  = 8'b00000000; // 1544 :   0 - 0x0
      13'h609: dout  = 8'b00001111; // 1545 :  15 - 0xf
      13'h60A: dout  = 8'b00101000; // 1546 :  40 - 0x28
      13'h60B: dout  = 8'b01011100; // 1547 :  92 - 0x5c
      13'h60C: dout  = 8'b00111111; // 1548 :  63 - 0x3f
      13'h60D: dout  = 8'b01111111; // 1549 : 127 - 0x7f
      13'h60E: dout  = 8'b01111111; // 1550 : 127 - 0x7f
      13'h60F: dout  = 8'b01111111; // 1551 : 127 - 0x7f
      13'h610: dout  = 8'b01111111; // 1552 : 127 - 0x7f -- Sprite 0x61
      13'h611: dout  = 8'b00111110; // 1553 :  62 - 0x3e
      13'h612: dout  = 8'b00011111; // 1554 :  31 - 0x1f
      13'h613: dout  = 8'b00011111; // 1555 :  31 - 0x1f
      13'h614: dout  = 8'b00001111; // 1556 :  15 - 0xf
      13'h615: dout  = 8'b00001111; // 1557 :  15 - 0xf
      13'h616: dout  = 8'b00001111; // 1558 :  15 - 0xf
      13'h617: dout  = 8'b00000111; // 1559 :   7 - 0x7
      13'h618: dout  = 8'b01111111; // 1560 : 127 - 0x7f
      13'h619: dout  = 8'b00111110; // 1561 :  62 - 0x3e
      13'h61A: dout  = 8'b00011111; // 1562 :  31 - 0x1f
      13'h61B: dout  = 8'b00011111; // 1563 :  31 - 0x1f
      13'h61C: dout  = 8'b00001000; // 1564 :   8 - 0x8
      13'h61D: dout  = 8'b00000000; // 1565 :   0 - 0x0
      13'h61E: dout  = 8'b00000000; // 1566 :   0 - 0x0
      13'h61F: dout  = 8'b00000000; // 1567 :   0 - 0x0
      13'h620: dout  = 8'b00000000; // 1568 :   0 - 0x0 -- Sprite 0x62
      13'h621: dout  = 8'b01100000; // 1569 :  96 - 0x60
      13'h622: dout  = 8'b11110000; // 1570 : 240 - 0xf0
      13'h623: dout  = 8'b11111000; // 1571 : 248 - 0xf8
      13'h624: dout  = 8'b11111000; // 1572 : 248 - 0xf8
      13'h625: dout  = 8'b11111000; // 1573 : 248 - 0xf8
      13'h626: dout  = 8'b11111100; // 1574 : 252 - 0xfc
      13'h627: dout  = 8'b11111100; // 1575 : 252 - 0xfc
      13'h628: dout  = 8'b00000000; // 1576 :   0 - 0x0
      13'h629: dout  = 8'b10000000; // 1577 : 128 - 0x80
      13'h62A: dout  = 8'b01000000; // 1578 :  64 - 0x40
      13'h62B: dout  = 8'b11000100; // 1579 : 196 - 0xc4
      13'h62C: dout  = 8'b11110110; // 1580 : 246 - 0xf6
      13'h62D: dout  = 8'b11111110; // 1581 : 254 - 0xfe
      13'h62E: dout  = 8'b11111100; // 1582 : 252 - 0xfc
      13'h62F: dout  = 8'b11111100; // 1583 : 252 - 0xfc
      13'h630: dout  = 8'b11111000; // 1584 : 248 - 0xf8 -- Sprite 0x63
      13'h631: dout  = 8'b11110000; // 1585 : 240 - 0xf0
      13'h632: dout  = 8'b11110000; // 1586 : 240 - 0xf0
      13'h633: dout  = 8'b11100000; // 1587 : 224 - 0xe0
      13'h634: dout  = 8'b10000000; // 1588 : 128 - 0x80
      13'h635: dout  = 8'b10000000; // 1589 : 128 - 0x80
      13'h636: dout  = 8'b11000000; // 1590 : 192 - 0xc0
      13'h637: dout  = 8'b11000000; // 1591 : 192 - 0xc0
      13'h638: dout  = 8'b11111000; // 1592 : 248 - 0xf8
      13'h639: dout  = 8'b11110000; // 1593 : 240 - 0xf0
      13'h63A: dout  = 8'b00000000; // 1594 :   0 - 0x0
      13'h63B: dout  = 8'b00000000; // 1595 :   0 - 0x0
      13'h63C: dout  = 8'b10000000; // 1596 : 128 - 0x80
      13'h63D: dout  = 8'b00000000; // 1597 :   0 - 0x0
      13'h63E: dout  = 8'b00000000; // 1598 :   0 - 0x0
      13'h63F: dout  = 8'b00000000; // 1599 :   0 - 0x0
      13'h640: dout  = 8'b00000000; // 1600 :   0 - 0x0 -- Sprite 0x64
      13'h641: dout  = 8'b00011111; // 1601 :  31 - 0x1f
      13'h642: dout  = 8'b00111111; // 1602 :  63 - 0x3f
      13'h643: dout  = 8'b01111111; // 1603 : 127 - 0x7f
      13'h644: dout  = 8'b11111111; // 1604 : 255 - 0xff
      13'h645: dout  = 8'b11111111; // 1605 : 255 - 0xff
      13'h646: dout  = 8'b00111110; // 1606 :  62 - 0x3e
      13'h647: dout  = 8'b00001111; // 1607 :  15 - 0xf
      13'h648: dout  = 8'b00000000; // 1608 :   0 - 0x0
      13'h649: dout  = 8'b00011100; // 1609 :  28 - 0x1c
      13'h64A: dout  = 8'b00111111; // 1610 :  63 - 0x3f
      13'h64B: dout  = 8'b01111111; // 1611 : 127 - 0x7f
      13'h64C: dout  = 8'b11111111; // 1612 : 255 - 0xff
      13'h64D: dout  = 8'b11111111; // 1613 : 255 - 0xff
      13'h64E: dout  = 8'b00111110; // 1614 :  62 - 0x3e
      13'h64F: dout  = 8'b01110000; // 1615 : 112 - 0x70
      13'h650: dout  = 8'b00000000; // 1616 :   0 - 0x0 -- Sprite 0x65
      13'h651: dout  = 8'b00000000; // 1617 :   0 - 0x0
      13'h652: dout  = 8'b00000000; // 1618 :   0 - 0x0
      13'h653: dout  = 8'b00000001; // 1619 :   1 - 0x1
      13'h654: dout  = 8'b00000000; // 1620 :   0 - 0x0
      13'h655: dout  = 8'b00000000; // 1621 :   0 - 0x0
      13'h656: dout  = 8'b00000000; // 1622 :   0 - 0x0
      13'h657: dout  = 8'b00000000; // 1623 :   0 - 0x0
      13'h658: dout  = 8'b00000000; // 1624 :   0 - 0x0
      13'h659: dout  = 8'b00000000; // 1625 :   0 - 0x0
      13'h65A: dout  = 8'b00000000; // 1626 :   0 - 0x0
      13'h65B: dout  = 8'b00000000; // 1627 :   0 - 0x0
      13'h65C: dout  = 8'b00000000; // 1628 :   0 - 0x0
      13'h65D: dout  = 8'b00000000; // 1629 :   0 - 0x0
      13'h65E: dout  = 8'b00000000; // 1630 :   0 - 0x0
      13'h65F: dout  = 8'b00000000; // 1631 :   0 - 0x0
      13'h660: dout  = 8'b00000000; // 1632 :   0 - 0x0 -- Sprite 0x66
      13'h661: dout  = 8'b11100000; // 1633 : 224 - 0xe0
      13'h662: dout  = 8'b11110000; // 1634 : 240 - 0xf0
      13'h663: dout  = 8'b11111100; // 1635 : 252 - 0xfc
      13'h664: dout  = 8'b11111110; // 1636 : 254 - 0xfe
      13'h665: dout  = 8'b11111110; // 1637 : 254 - 0xfe
      13'h666: dout  = 8'b11111111; // 1638 : 255 - 0xff
      13'h667: dout  = 8'b11111100; // 1639 : 252 - 0xfc
      13'h668: dout  = 8'b00000000; // 1640 :   0 - 0x0
      13'h669: dout  = 8'b01100000; // 1641 :  96 - 0x60
      13'h66A: dout  = 8'b11110000; // 1642 : 240 - 0xf0
      13'h66B: dout  = 8'b11111000; // 1643 : 248 - 0xf8
      13'h66C: dout  = 8'b11111100; // 1644 : 252 - 0xfc
      13'h66D: dout  = 8'b11111100; // 1645 : 252 - 0xfc
      13'h66E: dout  = 8'b11111100; // 1646 : 252 - 0xfc
      13'h66F: dout  = 8'b11111111; // 1647 : 255 - 0xff
      13'h670: dout  = 8'b01111100; // 1648 : 124 - 0x7c -- Sprite 0x67
      13'h671: dout  = 8'b11111100; // 1649 : 252 - 0xfc
      13'h672: dout  = 8'b11111000; // 1650 : 248 - 0xf8
      13'h673: dout  = 8'b11110000; // 1651 : 240 - 0xf0
      13'h674: dout  = 8'b11100000; // 1652 : 224 - 0xe0
      13'h675: dout  = 8'b00000000; // 1653 :   0 - 0x0
      13'h676: dout  = 8'b00000000; // 1654 :   0 - 0x0
      13'h677: dout  = 8'b00000000; // 1655 :   0 - 0x0
      13'h678: dout  = 8'b01111100; // 1656 : 124 - 0x7c
      13'h679: dout  = 8'b11111100; // 1657 : 252 - 0xfc
      13'h67A: dout  = 8'b10001000; // 1658 : 136 - 0x88
      13'h67B: dout  = 8'b00000000; // 1659 :   0 - 0x0
      13'h67C: dout  = 8'b00000000; // 1660 :   0 - 0x0
      13'h67D: dout  = 8'b00000000; // 1661 :   0 - 0x0
      13'h67E: dout  = 8'b00000000; // 1662 :   0 - 0x0
      13'h67F: dout  = 8'b00000000; // 1663 :   0 - 0x0
      13'h680: dout  = 8'b00000000; // 1664 :   0 - 0x0 -- Sprite 0x68
      13'h681: dout  = 8'b00000111; // 1665 :   7 - 0x7
      13'h682: dout  = 8'b00000111; // 1666 :   7 - 0x7
      13'h683: dout  = 8'b00001111; // 1667 :  15 - 0xf
      13'h684: dout  = 8'b00001111; // 1668 :  15 - 0xf
      13'h685: dout  = 8'b00000000; // 1669 :   0 - 0x0
      13'h686: dout  = 8'b00011111; // 1670 :  31 - 0x1f
      13'h687: dout  = 8'b00111111; // 1671 :  63 - 0x3f
      13'h688: dout  = 8'b00000000; // 1672 :   0 - 0x0
      13'h689: dout  = 8'b00000111; // 1673 :   7 - 0x7
      13'h68A: dout  = 8'b00000011; // 1674 :   3 - 0x3
      13'h68B: dout  = 8'b00000000; // 1675 :   0 - 0x0
      13'h68C: dout  = 8'b00000000; // 1676 :   0 - 0x0
      13'h68D: dout  = 8'b00000111; // 1677 :   7 - 0x7
      13'h68E: dout  = 8'b00000100; // 1678 :   4 - 0x4
      13'h68F: dout  = 8'b00000100; // 1679 :   4 - 0x4
      13'h690: dout  = 8'b01111111; // 1680 : 127 - 0x7f -- Sprite 0x69
      13'h691: dout  = 8'b01111111; // 1681 : 127 - 0x7f
      13'h692: dout  = 8'b00011111; // 1682 :  31 - 0x1f
      13'h693: dout  = 8'b00011111; // 1683 :  31 - 0x1f
      13'h694: dout  = 8'b00011111; // 1684 :  31 - 0x1f
      13'h695: dout  = 8'b00011110; // 1685 :  30 - 0x1e
      13'h696: dout  = 8'b00001111; // 1686 :  15 - 0xf
      13'h697: dout  = 8'b00011111; // 1687 :  31 - 0x1f
      13'h698: dout  = 8'b00001100; // 1688 :  12 - 0xc
      13'h699: dout  = 8'b10011110; // 1689 : 158 - 0x9e
      13'h69A: dout  = 8'b11111111; // 1690 : 255 - 0xff
      13'h69B: dout  = 8'b00011111; // 1691 :  31 - 0x1f
      13'h69C: dout  = 8'b00011111; // 1692 :  31 - 0x1f
      13'h69D: dout  = 8'b00011110; // 1693 :  30 - 0x1e
      13'h69E: dout  = 8'b00001111; // 1694 :  15 - 0xf
      13'h69F: dout  = 8'b00000000; // 1695 :   0 - 0x0
      13'h6A0: dout  = 8'b00000000; // 1696 :   0 - 0x0 -- Sprite 0x6a
      13'h6A1: dout  = 8'b11100000; // 1697 : 224 - 0xe0
      13'h6A2: dout  = 8'b11100000; // 1698 : 224 - 0xe0
      13'h6A3: dout  = 8'b11110000; // 1699 : 240 - 0xf0
      13'h6A4: dout  = 8'b11110000; // 1700 : 240 - 0xf0
      13'h6A5: dout  = 8'b00000000; // 1701 :   0 - 0x0
      13'h6A6: dout  = 8'b11111000; // 1702 : 248 - 0xf8
      13'h6A7: dout  = 8'b11111100; // 1703 : 252 - 0xfc
      13'h6A8: dout  = 8'b00000000; // 1704 :   0 - 0x0
      13'h6A9: dout  = 8'b11100000; // 1705 : 224 - 0xe0
      13'h6AA: dout  = 8'b11000000; // 1706 : 192 - 0xc0
      13'h6AB: dout  = 8'b00000000; // 1707 :   0 - 0x0
      13'h6AC: dout  = 8'b00000000; // 1708 :   0 - 0x0
      13'h6AD: dout  = 8'b11100000; // 1709 : 224 - 0xe0
      13'h6AE: dout  = 8'b00100000; // 1710 :  32 - 0x20
      13'h6AF: dout  = 8'b00100000; // 1711 :  32 - 0x20
      13'h6B0: dout  = 8'b11111110; // 1712 : 254 - 0xfe -- Sprite 0x6b
      13'h6B1: dout  = 8'b11111110; // 1713 : 254 - 0xfe
      13'h6B2: dout  = 8'b11111000; // 1714 : 248 - 0xf8
      13'h6B3: dout  = 8'b11111000; // 1715 : 248 - 0xf8
      13'h6B4: dout  = 8'b11111000; // 1716 : 248 - 0xf8
      13'h6B5: dout  = 8'b01111000; // 1717 : 120 - 0x78
      13'h6B6: dout  = 8'b11110000; // 1718 : 240 - 0xf0
      13'h6B7: dout  = 8'b11111000; // 1719 : 248 - 0xf8
      13'h6B8: dout  = 8'b00110000; // 1720 :  48 - 0x30
      13'h6B9: dout  = 8'b01111001; // 1721 : 121 - 0x79
      13'h6BA: dout  = 8'b11111111; // 1722 : 255 - 0xff
      13'h6BB: dout  = 8'b11111000; // 1723 : 248 - 0xf8
      13'h6BC: dout  = 8'b11111000; // 1724 : 248 - 0xf8
      13'h6BD: dout  = 8'b01111000; // 1725 : 120 - 0x78
      13'h6BE: dout  = 8'b11110000; // 1726 : 240 - 0xf0
      13'h6BF: dout  = 8'b00000000; // 1727 :   0 - 0x0
      13'h6C0: dout  = 8'b00000011; // 1728 :   3 - 0x3 -- Sprite 0x6c
      13'h6C1: dout  = 8'b00000111; // 1729 :   7 - 0x7
      13'h6C2: dout  = 8'b00000101; // 1730 :   5 - 0x5
      13'h6C3: dout  = 8'b00001000; // 1731 :   8 - 0x8
      13'h6C4: dout  = 8'b00011011; // 1732 :  27 - 0x1b
      13'h6C5: dout  = 8'b00011001; // 1733 :  25 - 0x19
      13'h6C6: dout  = 8'b00000101; // 1734 :   5 - 0x5
      13'h6C7: dout  = 8'b00111111; // 1735 :  63 - 0x3f
      13'h6C8: dout  = 8'b00000011; // 1736 :   3 - 0x3
      13'h6C9: dout  = 8'b00000111; // 1737 :   7 - 0x7
      13'h6CA: dout  = 8'b00000010; // 1738 :   2 - 0x2
      13'h6CB: dout  = 8'b00000111; // 1739 :   7 - 0x7
      13'h6CC: dout  = 8'b00000100; // 1740 :   4 - 0x4
      13'h6CD: dout  = 8'b01000110; // 1741 :  70 - 0x46
      13'h6CE: dout  = 8'b11100011; // 1742 : 227 - 0xe3
      13'h6CF: dout  = 8'b11000010; // 1743 : 194 - 0xc2
      13'h6D0: dout  = 8'b00111111; // 1744 :  63 - 0x3f -- Sprite 0x6d
      13'h6D1: dout  = 8'b00001111; // 1745 :  15 - 0xf
      13'h6D2: dout  = 8'b00000101; // 1746 :   5 - 0x5
      13'h6D3: dout  = 8'b00110111; // 1747 :  55 - 0x37
      13'h6D4: dout  = 8'b00111111; // 1748 :  63 - 0x3f
      13'h6D5: dout  = 8'b00111111; // 1749 :  63 - 0x3f
      13'h6D6: dout  = 8'b00111110; // 1750 :  62 - 0x3e
      13'h6D7: dout  = 8'b00011100; // 1751 :  28 - 0x1c
      13'h6D8: dout  = 8'b01000010; // 1752 :  66 - 0x42
      13'h6D9: dout  = 8'b00000111; // 1753 :   7 - 0x7
      13'h6DA: dout  = 8'b00000111; // 1754 :   7 - 0x7
      13'h6DB: dout  = 8'b00000111; // 1755 :   7 - 0x7
      13'h6DC: dout  = 8'b00000111; // 1756 :   7 - 0x7
      13'h6DD: dout  = 8'b00000011; // 1757 :   3 - 0x3
      13'h6DE: dout  = 8'b00000010; // 1758 :   2 - 0x2
      13'h6DF: dout  = 8'b00000000; // 1759 :   0 - 0x0
      13'h6E0: dout  = 8'b11100000; // 1760 : 224 - 0xe0 -- Sprite 0x6e
      13'h6E1: dout  = 8'b11110000; // 1761 : 240 - 0xf0
      13'h6E2: dout  = 8'b01010000; // 1762 :  80 - 0x50
      13'h6E3: dout  = 8'b00001000; // 1763 :   8 - 0x8
      13'h6E4: dout  = 8'b01101100; // 1764 : 108 - 0x6c
      13'h6E5: dout  = 8'b11001100; // 1765 : 204 - 0xcc
      13'h6E6: dout  = 8'b11010000; // 1766 : 208 - 0xd0
      13'h6E7: dout  = 8'b11111110; // 1767 : 254 - 0xfe
      13'h6E8: dout  = 8'b11100000; // 1768 : 224 - 0xe0
      13'h6E9: dout  = 8'b11110000; // 1769 : 240 - 0xf0
      13'h6EA: dout  = 8'b10100000; // 1770 : 160 - 0xa0
      13'h6EB: dout  = 8'b11110000; // 1771 : 240 - 0xf0
      13'h6EC: dout  = 8'b10010000; // 1772 : 144 - 0x90
      13'h6ED: dout  = 8'b00110010; // 1773 :  50 - 0x32
      13'h6EE: dout  = 8'b11100011; // 1774 : 227 - 0xe3
      13'h6EF: dout  = 8'b00100001; // 1775 :  33 - 0x21
      13'h6F0: dout  = 8'b11111110; // 1776 : 254 - 0xfe -- Sprite 0x6f
      13'h6F1: dout  = 8'b11111000; // 1777 : 248 - 0xf8
      13'h6F2: dout  = 8'b11010000; // 1778 : 208 - 0xd0
      13'h6F3: dout  = 8'b11111011; // 1779 : 251 - 0xfb
      13'h6F4: dout  = 8'b11111111; // 1780 : 255 - 0xff
      13'h6F5: dout  = 8'b11111111; // 1781 : 255 - 0xff
      13'h6F6: dout  = 8'b00111110; // 1782 :  62 - 0x3e
      13'h6F7: dout  = 8'b00001100; // 1783 :  12 - 0xc
      13'h6F8: dout  = 8'b00100000; // 1784 :  32 - 0x20
      13'h6F9: dout  = 8'b01110000; // 1785 : 112 - 0x70
      13'h6FA: dout  = 8'b11110000; // 1786 : 240 - 0xf0
      13'h6FB: dout  = 8'b11111000; // 1787 : 248 - 0xf8
      13'h6FC: dout  = 8'b11111000; // 1788 : 248 - 0xf8
      13'h6FD: dout  = 8'b11110000; // 1789 : 240 - 0xf0
      13'h6FE: dout  = 8'b00110000; // 1790 :  48 - 0x30
      13'h6FF: dout  = 8'b00000000; // 1791 :   0 - 0x0
      13'h700: dout  = 8'b00000000; // 1792 :   0 - 0x0 -- Sprite 0x70
      13'h701: dout  = 8'b00000000; // 1793 :   0 - 0x0
      13'h702: dout  = 8'b01111001; // 1794 : 121 - 0x79
      13'h703: dout  = 8'b11111001; // 1795 : 249 - 0xf9
      13'h704: dout  = 8'b11110011; // 1796 : 243 - 0xf3
      13'h705: dout  = 8'b11111111; // 1797 : 255 - 0xff
      13'h706: dout  = 8'b01111011; // 1798 : 123 - 0x7b
      13'h707: dout  = 8'b00111111; // 1799 :  63 - 0x3f
      13'h708: dout  = 8'b00000000; // 1800 :   0 - 0x0
      13'h709: dout  = 8'b00000001; // 1801 :   1 - 0x1
      13'h70A: dout  = 8'b00000000; // 1802 :   0 - 0x0
      13'h70B: dout  = 8'b00000000; // 1803 :   0 - 0x0
      13'h70C: dout  = 8'b00000000; // 1804 :   0 - 0x0
      13'h70D: dout  = 8'b00011110; // 1805 :  30 - 0x1e
      13'h70E: dout  = 8'b01111111; // 1806 : 127 - 0x7f
      13'h70F: dout  = 8'b00111110; // 1807 :  62 - 0x3e
      13'h710: dout  = 8'b00111111; // 1808 :  63 - 0x3f -- Sprite 0x71
      13'h711: dout  = 8'b00111111; // 1809 :  63 - 0x3f
      13'h712: dout  = 8'b01111011; // 1810 : 123 - 0x7b
      13'h713: dout  = 8'b01111111; // 1811 : 127 - 0x7f
      13'h714: dout  = 8'b11111011; // 1812 : 251 - 0xfb
      13'h715: dout  = 8'b11110001; // 1813 : 241 - 0xf1
      13'h716: dout  = 8'b01111001; // 1814 : 121 - 0x79
      13'h717: dout  = 8'b00111000; // 1815 :  56 - 0x38
      13'h718: dout  = 8'b00111100; // 1816 :  60 - 0x3c
      13'h719: dout  = 8'b00111110; // 1817 :  62 - 0x3e
      13'h71A: dout  = 8'b01111111; // 1818 : 127 - 0x7f
      13'h71B: dout  = 8'b01111110; // 1819 : 126 - 0x7e
      13'h71C: dout  = 8'b00011000; // 1820 :  24 - 0x18
      13'h71D: dout  = 8'b00000000; // 1821 :   0 - 0x0
      13'h71E: dout  = 8'b00000000; // 1822 :   0 - 0x0
      13'h71F: dout  = 8'b00000000; // 1823 :   0 - 0x0
      13'h720: dout  = 8'b00000000; // 1824 :   0 - 0x0 -- Sprite 0x72
      13'h721: dout  = 8'b00000000; // 1825 :   0 - 0x0
      13'h722: dout  = 8'b10000000; // 1826 : 128 - 0x80
      13'h723: dout  = 8'b10110000; // 1827 : 176 - 0xb0
      13'h724: dout  = 8'b10111000; // 1828 : 184 - 0xb8
      13'h725: dout  = 8'b11000110; // 1829 : 198 - 0xc6
      13'h726: dout  = 8'b10010011; // 1830 : 147 - 0x93
      13'h727: dout  = 8'b11110111; // 1831 : 247 - 0xf7
      13'h728: dout  = 8'b11000000; // 1832 : 192 - 0xc0
      13'h729: dout  = 8'b11100000; // 1833 : 224 - 0xe0
      13'h72A: dout  = 8'b01000000; // 1834 :  64 - 0x40
      13'h72B: dout  = 8'b00000000; // 1835 :   0 - 0x0
      13'h72C: dout  = 8'b00000000; // 1836 :   0 - 0x0
      13'h72D: dout  = 8'b00111010; // 1837 :  58 - 0x3a
      13'h72E: dout  = 8'b11101111; // 1838 : 239 - 0xef
      13'h72F: dout  = 8'b01001011; // 1839 :  75 - 0x4b
      13'h730: dout  = 8'b11100011; // 1840 : 227 - 0xe3 -- Sprite 0x73
      13'h731: dout  = 8'b11110111; // 1841 : 247 - 0xf7
      13'h732: dout  = 8'b10010011; // 1842 : 147 - 0x93
      13'h733: dout  = 8'b11000110; // 1843 : 198 - 0xc6
      13'h734: dout  = 8'b10111000; // 1844 : 184 - 0xb8
      13'h735: dout  = 8'b10110000; // 1845 : 176 - 0xb0
      13'h736: dout  = 8'b10000000; // 1846 : 128 - 0x80
      13'h737: dout  = 8'b00000000; // 1847 :   0 - 0x0
      13'h738: dout  = 8'b01011111; // 1848 :  95 - 0x5f
      13'h739: dout  = 8'b01001011; // 1849 :  75 - 0x4b
      13'h73A: dout  = 8'b11101111; // 1850 : 239 - 0xef
      13'h73B: dout  = 8'b00111010; // 1851 :  58 - 0x3a
      13'h73C: dout  = 8'b00000000; // 1852 :   0 - 0x0
      13'h73D: dout  = 8'b00000000; // 1853 :   0 - 0x0
      13'h73E: dout  = 8'b01100000; // 1854 :  96 - 0x60
      13'h73F: dout  = 8'b11000000; // 1855 : 192 - 0xc0
      13'h740: dout  = 8'b00110000; // 1856 :  48 - 0x30 -- Sprite 0x74
      13'h741: dout  = 8'b01111100; // 1857 : 124 - 0x7c
      13'h742: dout  = 8'b11111111; // 1858 : 255 - 0xff
      13'h743: dout  = 8'b11111111; // 1859 : 255 - 0xff
      13'h744: dout  = 8'b11011111; // 1860 : 223 - 0xdf
      13'h745: dout  = 8'b00001011; // 1861 :  11 - 0xb
      13'h746: dout  = 8'b00011111; // 1862 :  31 - 0x1f
      13'h747: dout  = 8'b01111111; // 1863 : 127 - 0x7f
      13'h748: dout  = 8'b00000000; // 1864 :   0 - 0x0
      13'h749: dout  = 8'b00001100; // 1865 :  12 - 0xc
      13'h74A: dout  = 8'b00001111; // 1866 :  15 - 0xf
      13'h74B: dout  = 8'b00011111; // 1867 :  31 - 0x1f
      13'h74C: dout  = 8'b00011111; // 1868 :  31 - 0x1f
      13'h74D: dout  = 8'b00001111; // 1869 :  15 - 0xf
      13'h74E: dout  = 8'b00001110; // 1870 :  14 - 0xe
      13'h74F: dout  = 8'b00000100; // 1871 :   4 - 0x4
      13'h750: dout  = 8'b01111111; // 1872 : 127 - 0x7f -- Sprite 0x75
      13'h751: dout  = 8'b00001011; // 1873 :  11 - 0xb
      13'h752: dout  = 8'b00110011; // 1874 :  51 - 0x33
      13'h753: dout  = 8'b00110110; // 1875 :  54 - 0x36
      13'h754: dout  = 8'b00010000; // 1876 :  16 - 0x10
      13'h755: dout  = 8'b00001010; // 1877 :  10 - 0xa
      13'h756: dout  = 8'b00001111; // 1878 :  15 - 0xf
      13'h757: dout  = 8'b00000111; // 1879 :   7 - 0x7
      13'h758: dout  = 8'b10000100; // 1880 : 132 - 0x84
      13'h759: dout  = 8'b11000111; // 1881 : 199 - 0xc7
      13'h75A: dout  = 8'b01001100; // 1882 :  76 - 0x4c
      13'h75B: dout  = 8'b00001001; // 1883 :   9 - 0x9
      13'h75C: dout  = 8'b00001111; // 1884 :  15 - 0xf
      13'h75D: dout  = 8'b00000101; // 1885 :   5 - 0x5
      13'h75E: dout  = 8'b00001111; // 1886 :  15 - 0xf
      13'h75F: dout  = 8'b00000111; // 1887 :   7 - 0x7
      13'h760: dout  = 8'b00111000; // 1888 :  56 - 0x38 -- Sprite 0x76
      13'h761: dout  = 8'b01111100; // 1889 : 124 - 0x7c
      13'h762: dout  = 8'b11111100; // 1890 : 252 - 0xfc
      13'h763: dout  = 8'b11111100; // 1891 : 252 - 0xfc
      13'h764: dout  = 8'b11101100; // 1892 : 236 - 0xec
      13'h765: dout  = 8'b10100000; // 1893 : 160 - 0xa0
      13'h766: dout  = 8'b11110000; // 1894 : 240 - 0xf0
      13'h767: dout  = 8'b11111100; // 1895 : 252 - 0xfc
      13'h768: dout  = 8'b00000000; // 1896 :   0 - 0x0
      13'h769: dout  = 8'b01000000; // 1897 :  64 - 0x40
      13'h76A: dout  = 8'b11000000; // 1898 : 192 - 0xc0
      13'h76B: dout  = 8'b11100000; // 1899 : 224 - 0xe0
      13'h76C: dout  = 8'b11100000; // 1900 : 224 - 0xe0
      13'h76D: dout  = 8'b11100000; // 1901 : 224 - 0xe0
      13'h76E: dout  = 8'b11100000; // 1902 : 224 - 0xe0
      13'h76F: dout  = 8'b01000010; // 1903 :  66 - 0x42
      13'h770: dout  = 8'b11111100; // 1904 : 252 - 0xfc -- Sprite 0x77
      13'h771: dout  = 8'b10100000; // 1905 : 160 - 0xa0
      13'h772: dout  = 8'b10011000; // 1906 : 152 - 0x98
      13'h773: dout  = 8'b11011000; // 1907 : 216 - 0xd8
      13'h774: dout  = 8'b00010000; // 1908 :  16 - 0x10
      13'h775: dout  = 8'b10100000; // 1909 : 160 - 0xa0
      13'h776: dout  = 8'b11100000; // 1910 : 224 - 0xe0
      13'h777: dout  = 8'b11000000; // 1911 : 192 - 0xc0
      13'h778: dout  = 8'b01000011; // 1912 :  67 - 0x43
      13'h779: dout  = 8'b11000111; // 1913 : 199 - 0xc7
      13'h77A: dout  = 8'b01100010; // 1914 :  98 - 0x62
      13'h77B: dout  = 8'b00100000; // 1915 :  32 - 0x20
      13'h77C: dout  = 8'b11100000; // 1916 : 224 - 0xe0
      13'h77D: dout  = 8'b01000000; // 1917 :  64 - 0x40
      13'h77E: dout  = 8'b11100000; // 1918 : 224 - 0xe0
      13'h77F: dout  = 8'b11000000; // 1919 : 192 - 0xc0
      13'h780: dout  = 8'b00000000; // 1920 :   0 - 0x0 -- Sprite 0x78
      13'h781: dout  = 8'b00000001; // 1921 :   1 - 0x1
      13'h782: dout  = 8'b00001101; // 1922 :  13 - 0xd
      13'h783: dout  = 8'b00011101; // 1923 :  29 - 0x1d
      13'h784: dout  = 8'b01100011; // 1924 :  99 - 0x63
      13'h785: dout  = 8'b11001001; // 1925 : 201 - 0xc9
      13'h786: dout  = 8'b11101111; // 1926 : 239 - 0xef
      13'h787: dout  = 8'b11000111; // 1927 : 199 - 0xc7
      13'h788: dout  = 8'b00000011; // 1928 :   3 - 0x3
      13'h789: dout  = 8'b00000100; // 1929 :   4 - 0x4
      13'h78A: dout  = 8'b00000000; // 1930 :   0 - 0x0
      13'h78B: dout  = 8'b00000000; // 1931 :   0 - 0x0
      13'h78C: dout  = 8'b01011100; // 1932 :  92 - 0x5c
      13'h78D: dout  = 8'b11110111; // 1933 : 247 - 0xf7
      13'h78E: dout  = 8'b11010010; // 1934 : 210 - 0xd2
      13'h78F: dout  = 8'b11111010; // 1935 : 250 - 0xfa
      13'h790: dout  = 8'b11101111; // 1936 : 239 - 0xef -- Sprite 0x79
      13'h791: dout  = 8'b11001001; // 1937 : 201 - 0xc9
      13'h792: dout  = 8'b01100011; // 1938 :  99 - 0x63
      13'h793: dout  = 8'b00011101; // 1939 :  29 - 0x1d
      13'h794: dout  = 8'b00001101; // 1940 :  13 - 0xd
      13'h795: dout  = 8'b00000001; // 1941 :   1 - 0x1
      13'h796: dout  = 8'b00000000; // 1942 :   0 - 0x0
      13'h797: dout  = 8'b00000000; // 1943 :   0 - 0x0
      13'h798: dout  = 8'b11010010; // 1944 : 210 - 0xd2
      13'h799: dout  = 8'b11110111; // 1945 : 247 - 0xf7
      13'h79A: dout  = 8'b01011100; // 1946 :  92 - 0x5c
      13'h79B: dout  = 8'b00000000; // 1947 :   0 - 0x0
      13'h79C: dout  = 8'b00000000; // 1948 :   0 - 0x0
      13'h79D: dout  = 8'b00000010; // 1949 :   2 - 0x2
      13'h79E: dout  = 8'b00000111; // 1950 :   7 - 0x7
      13'h79F: dout  = 8'b00000011; // 1951 :   3 - 0x3
      13'h7A0: dout  = 8'b00011100; // 1952 :  28 - 0x1c -- Sprite 0x7a
      13'h7A1: dout  = 8'b10011110; // 1953 : 158 - 0x9e
      13'h7A2: dout  = 8'b10001111; // 1954 : 143 - 0x8f
      13'h7A3: dout  = 8'b11011111; // 1955 : 223 - 0xdf
      13'h7A4: dout  = 8'b11111110; // 1956 : 254 - 0xfe
      13'h7A5: dout  = 8'b11011110; // 1957 : 222 - 0xde
      13'h7A6: dout  = 8'b11111100; // 1958 : 252 - 0xfc
      13'h7A7: dout  = 8'b11111100; // 1959 : 252 - 0xfc
      13'h7A8: dout  = 8'b00000000; // 1960 :   0 - 0x0
      13'h7A9: dout  = 8'b00000000; // 1961 :   0 - 0x0
      13'h7AA: dout  = 8'b00000000; // 1962 :   0 - 0x0
      13'h7AB: dout  = 8'b00011000; // 1963 :  24 - 0x18
      13'h7AC: dout  = 8'b01111110; // 1964 : 126 - 0x7e
      13'h7AD: dout  = 8'b11111110; // 1965 : 254 - 0xfe
      13'h7AE: dout  = 8'b01111100; // 1966 : 124 - 0x7c
      13'h7AF: dout  = 8'b00111100; // 1967 :  60 - 0x3c
      13'h7B0: dout  = 8'b11111100; // 1968 : 252 - 0xfc -- Sprite 0x7b
      13'h7B1: dout  = 8'b11011110; // 1969 : 222 - 0xde
      13'h7B2: dout  = 8'b11111111; // 1970 : 255 - 0xff
      13'h7B3: dout  = 8'b11001111; // 1971 : 207 - 0xcf
      13'h7B4: dout  = 8'b10011111; // 1972 : 159 - 0x9f
      13'h7B5: dout  = 8'b10011110; // 1973 : 158 - 0x9e
      13'h7B6: dout  = 8'b00000000; // 1974 :   0 - 0x0
      13'h7B7: dout  = 8'b00000000; // 1975 :   0 - 0x0
      13'h7B8: dout  = 8'b01111100; // 1976 : 124 - 0x7c
      13'h7B9: dout  = 8'b11111110; // 1977 : 254 - 0xfe
      13'h7BA: dout  = 8'b01111000; // 1978 : 120 - 0x78
      13'h7BB: dout  = 8'b00000000; // 1979 :   0 - 0x0
      13'h7BC: dout  = 8'b00000000; // 1980 :   0 - 0x0
      13'h7BD: dout  = 8'b00000000; // 1981 :   0 - 0x0
      13'h7BE: dout  = 8'b10000000; // 1982 : 128 - 0x80
      13'h7BF: dout  = 8'b00000000; // 1983 :   0 - 0x0
      13'h7C0: dout  = 8'b00000000; // 1984 :   0 - 0x0 -- Sprite 0x7c
      13'h7C1: dout  = 8'b00000000; // 1985 :   0 - 0x0
      13'h7C2: dout  = 8'b00000000; // 1986 :   0 - 0x0
      13'h7C3: dout  = 8'b00000000; // 1987 :   0 - 0x0
      13'h7C4: dout  = 8'b00011110; // 1988 :  30 - 0x1e
      13'h7C5: dout  = 8'b00111111; // 1989 :  63 - 0x3f
      13'h7C6: dout  = 8'b01111101; // 1990 : 125 - 0x7d
      13'h7C7: dout  = 8'b01111000; // 1991 : 120 - 0x78
      13'h7C8: dout  = 8'b00000000; // 1992 :   0 - 0x0
      13'h7C9: dout  = 8'b00000000; // 1993 :   0 - 0x0
      13'h7CA: dout  = 8'b00000001; // 1994 :   1 - 0x1
      13'h7CB: dout  = 8'b00000000; // 1995 :   0 - 0x0
      13'h7CC: dout  = 8'b00000000; // 1996 :   0 - 0x0
      13'h7CD: dout  = 8'b00100000; // 1997 :  32 - 0x20
      13'h7CE: dout  = 8'b01111100; // 1998 : 124 - 0x7c
      13'h7CF: dout  = 8'b01111000; // 1999 : 120 - 0x78
      13'h7D0: dout  = 8'b01111100; // 2000 : 124 - 0x7c -- Sprite 0x7d
      13'h7D1: dout  = 8'b11111011; // 2001 : 251 - 0xfb
      13'h7D2: dout  = 8'b11111111; // 2002 : 255 - 0xff
      13'h7D3: dout  = 8'b11111111; // 2003 : 255 - 0xff
      13'h7D4: dout  = 8'b01011111; // 2004 :  95 - 0x5f
      13'h7D5: dout  = 8'b00011111; // 2005 :  31 - 0x1f
      13'h7D6: dout  = 8'b00011111; // 2006 :  31 - 0x1f
      13'h7D7: dout  = 8'b00011111; // 2007 :  31 - 0x1f
      13'h7D8: dout  = 8'b01111100; // 2008 : 124 - 0x7c
      13'h7D9: dout  = 8'b11111110; // 2009 : 254 - 0xfe
      13'h7DA: dout  = 8'b11111111; // 2010 : 255 - 0xff
      13'h7DB: dout  = 8'b11111110; // 2011 : 254 - 0xfe
      13'h7DC: dout  = 8'b01111100; // 2012 : 124 - 0x7c
      13'h7DD: dout  = 8'b01100000; // 2013 :  96 - 0x60
      13'h7DE: dout  = 8'b11100000; // 2014 : 224 - 0xe0
      13'h7DF: dout  = 8'b11100001; // 2015 : 225 - 0xe1
      13'h7E0: dout  = 8'b00000000; // 2016 :   0 - 0x0 -- Sprite 0x7e
      13'h7E1: dout  = 8'b00000000; // 2017 :   0 - 0x0
      13'h7E2: dout  = 8'b00000000; // 2018 :   0 - 0x0
      13'h7E3: dout  = 8'b00000000; // 2019 :   0 - 0x0
      13'h7E4: dout  = 8'b00000000; // 2020 :   0 - 0x0
      13'h7E5: dout  = 8'b10000000; // 2021 : 128 - 0x80
      13'h7E6: dout  = 8'b10000000; // 2022 : 128 - 0x80
      13'h7E7: dout  = 8'b00000000; // 2023 :   0 - 0x0
      13'h7E8: dout  = 8'b01111100; // 2024 : 124 - 0x7c
      13'h7E9: dout  = 8'b10000010; // 2025 : 130 - 0x82
      13'h7EA: dout  = 8'b00000001; // 2026 :   1 - 0x1
      13'h7EB: dout  = 8'b10000010; // 2027 : 130 - 0x82
      13'h7EC: dout  = 8'b01111100; // 2028 : 124 - 0x7c
      13'h7ED: dout  = 8'b00000000; // 2029 :   0 - 0x0
      13'h7EE: dout  = 8'b00000000; // 2030 :   0 - 0x0
      13'h7EF: dout  = 8'b00000000; // 2031 :   0 - 0x0
      13'h7F0: dout  = 8'b00000000; // 2032 :   0 - 0x0 -- Sprite 0x7f
      13'h7F1: dout  = 8'b00100001; // 2033 :  33 - 0x21
      13'h7F2: dout  = 8'b10100010; // 2034 : 162 - 0xa2
      13'h7F3: dout  = 8'b10100011; // 2035 : 163 - 0xa3
      13'h7F4: dout  = 8'b10110011; // 2036 : 179 - 0xb3
      13'h7F5: dout  = 8'b10001111; // 2037 : 143 - 0x8f
      13'h7F6: dout  = 8'b00100111; // 2038 :  39 - 0x27
      13'h7F7: dout  = 8'b11111110; // 2039 : 254 - 0xfe
      13'h7F8: dout  = 8'b00010000; // 2040 :  16 - 0x10
      13'h7F9: dout  = 8'b00011001; // 2041 :  25 - 0x19
      13'h7FA: dout  = 8'b01011010; // 2042 :  90 - 0x5a
      13'h7FB: dout  = 8'b11011111; // 2043 : 223 - 0xdf
      13'h7FC: dout  = 8'b01001111; // 2044 :  79 - 0x4f
      13'h7FD: dout  = 8'b01110011; // 2045 : 115 - 0x73
      13'h7FE: dout  = 8'b11011011; // 2046 : 219 - 0xdb
      13'h7FF: dout  = 8'b00000010; // 2047 :   2 - 0x2
      13'h800: dout  = 8'b00000000; // 2048 :   0 - 0x0 -- Sprite 0x80
      13'h801: dout  = 8'b00000000; // 2049 :   0 - 0x0
      13'h802: dout  = 8'b00000000; // 2050 :   0 - 0x0
      13'h803: dout  = 8'b00000000; // 2051 :   0 - 0x0
      13'h804: dout  = 8'b00000011; // 2052 :   3 - 0x3
      13'h805: dout  = 8'b00001111; // 2053 :  15 - 0xf
      13'h806: dout  = 8'b00011111; // 2054 :  31 - 0x1f
      13'h807: dout  = 8'b00011111; // 2055 :  31 - 0x1f
      13'h808: dout  = 8'b00000000; // 2056 :   0 - 0x0
      13'h809: dout  = 8'b00000000; // 2057 :   0 - 0x0
      13'h80A: dout  = 8'b00000000; // 2058 :   0 - 0x0
      13'h80B: dout  = 8'b00000011; // 2059 :   3 - 0x3
      13'h80C: dout  = 8'b00001100; // 2060 :  12 - 0xc
      13'h80D: dout  = 8'b00010000; // 2061 :  16 - 0x10
      13'h80E: dout  = 8'b00100010; // 2062 :  34 - 0x22
      13'h80F: dout  = 8'b00100000; // 2063 :  32 - 0x20
      13'h810: dout  = 8'b00011111; // 2064 :  31 - 0x1f -- Sprite 0x81
      13'h811: dout  = 8'b00011111; // 2065 :  31 - 0x1f
      13'h812: dout  = 8'b00001111; // 2066 :  15 - 0xf
      13'h813: dout  = 8'b00000011; // 2067 :   3 - 0x3
      13'h814: dout  = 8'b00000000; // 2068 :   0 - 0x0
      13'h815: dout  = 8'b00000000; // 2069 :   0 - 0x0
      13'h816: dout  = 8'b00000000; // 2070 :   0 - 0x0
      13'h817: dout  = 8'b00000000; // 2071 :   0 - 0x0
      13'h818: dout  = 8'b00100001; // 2072 :  33 - 0x21
      13'h819: dout  = 8'b00100011; // 2073 :  35 - 0x23
      13'h81A: dout  = 8'b00010000; // 2074 :  16 - 0x10
      13'h81B: dout  = 8'b00001100; // 2075 :  12 - 0xc
      13'h81C: dout  = 8'b00000011; // 2076 :   3 - 0x3
      13'h81D: dout  = 8'b00000000; // 2077 :   0 - 0x0
      13'h81E: dout  = 8'b00000000; // 2078 :   0 - 0x0
      13'h81F: dout  = 8'b00000000; // 2079 :   0 - 0x0
      13'h820: dout  = 8'b00000000; // 2080 :   0 - 0x0 -- Sprite 0x82
      13'h821: dout  = 8'b00000000; // 2081 :   0 - 0x0
      13'h822: dout  = 8'b00000000; // 2082 :   0 - 0x0
      13'h823: dout  = 8'b00000000; // 2083 :   0 - 0x0
      13'h824: dout  = 8'b11000000; // 2084 : 192 - 0xc0
      13'h825: dout  = 8'b11110000; // 2085 : 240 - 0xf0
      13'h826: dout  = 8'b11111000; // 2086 : 248 - 0xf8
      13'h827: dout  = 8'b11111000; // 2087 : 248 - 0xf8
      13'h828: dout  = 8'b00000000; // 2088 :   0 - 0x0
      13'h829: dout  = 8'b00000000; // 2089 :   0 - 0x0
      13'h82A: dout  = 8'b00000000; // 2090 :   0 - 0x0
      13'h82B: dout  = 8'b11000000; // 2091 : 192 - 0xc0
      13'h82C: dout  = 8'b00110000; // 2092 :  48 - 0x30
      13'h82D: dout  = 8'b00001000; // 2093 :   8 - 0x8
      13'h82E: dout  = 8'b01100100; // 2094 : 100 - 0x64
      13'h82F: dout  = 8'b11000100; // 2095 : 196 - 0xc4
      13'h830: dout  = 8'b11111000; // 2096 : 248 - 0xf8 -- Sprite 0x83
      13'h831: dout  = 8'b11111000; // 2097 : 248 - 0xf8
      13'h832: dout  = 8'b11110000; // 2098 : 240 - 0xf0
      13'h833: dout  = 8'b11000000; // 2099 : 192 - 0xc0
      13'h834: dout  = 8'b00000000; // 2100 :   0 - 0x0
      13'h835: dout  = 8'b00000000; // 2101 :   0 - 0x0
      13'h836: dout  = 8'b00000000; // 2102 :   0 - 0x0
      13'h837: dout  = 8'b00000000; // 2103 :   0 - 0x0
      13'h838: dout  = 8'b10000100; // 2104 : 132 - 0x84
      13'h839: dout  = 8'b00000100; // 2105 :   4 - 0x4
      13'h83A: dout  = 8'b00001000; // 2106 :   8 - 0x8
      13'h83B: dout  = 8'b00110000; // 2107 :  48 - 0x30
      13'h83C: dout  = 8'b11000000; // 2108 : 192 - 0xc0
      13'h83D: dout  = 8'b00000000; // 2109 :   0 - 0x0
      13'h83E: dout  = 8'b00000000; // 2110 :   0 - 0x0
      13'h83F: dout  = 8'b00000000; // 2111 :   0 - 0x0
      13'h840: dout  = 8'b00000000; // 2112 :   0 - 0x0 -- Sprite 0x84
      13'h841: dout  = 8'b00000000; // 2113 :   0 - 0x0
      13'h842: dout  = 8'b00000000; // 2114 :   0 - 0x0
      13'h843: dout  = 8'b00000000; // 2115 :   0 - 0x0
      13'h844: dout  = 8'b00000011; // 2116 :   3 - 0x3
      13'h845: dout  = 8'b00001111; // 2117 :  15 - 0xf
      13'h846: dout  = 8'b00011111; // 2118 :  31 - 0x1f
      13'h847: dout  = 8'b00011111; // 2119 :  31 - 0x1f
      13'h848: dout  = 8'b00000000; // 2120 :   0 - 0x0
      13'h849: dout  = 8'b00000000; // 2121 :   0 - 0x0
      13'h84A: dout  = 8'b00000000; // 2122 :   0 - 0x0
      13'h84B: dout  = 8'b00000011; // 2123 :   3 - 0x3
      13'h84C: dout  = 8'b00001100; // 2124 :  12 - 0xc
      13'h84D: dout  = 8'b00010000; // 2125 :  16 - 0x10
      13'h84E: dout  = 8'b00100110; // 2126 :  38 - 0x26
      13'h84F: dout  = 8'b00100011; // 2127 :  35 - 0x23
      13'h850: dout  = 8'b00011111; // 2128 :  31 - 0x1f -- Sprite 0x85
      13'h851: dout  = 8'b00011111; // 2129 :  31 - 0x1f
      13'h852: dout  = 8'b00001111; // 2130 :  15 - 0xf
      13'h853: dout  = 8'b00000011; // 2131 :   3 - 0x3
      13'h854: dout  = 8'b00000000; // 2132 :   0 - 0x0
      13'h855: dout  = 8'b00000000; // 2133 :   0 - 0x0
      13'h856: dout  = 8'b00000000; // 2134 :   0 - 0x0
      13'h857: dout  = 8'b00000000; // 2135 :   0 - 0x0
      13'h858: dout  = 8'b00100001; // 2136 :  33 - 0x21
      13'h859: dout  = 8'b00100000; // 2137 :  32 - 0x20
      13'h85A: dout  = 8'b00010000; // 2138 :  16 - 0x10
      13'h85B: dout  = 8'b00001100; // 2139 :  12 - 0xc
      13'h85C: dout  = 8'b00000011; // 2140 :   3 - 0x3
      13'h85D: dout  = 8'b00000000; // 2141 :   0 - 0x0
      13'h85E: dout  = 8'b00000000; // 2142 :   0 - 0x0
      13'h85F: dout  = 8'b00000000; // 2143 :   0 - 0x0
      13'h860: dout  = 8'b00000000; // 2144 :   0 - 0x0 -- Sprite 0x86
      13'h861: dout  = 8'b00000000; // 2145 :   0 - 0x0
      13'h862: dout  = 8'b00000000; // 2146 :   0 - 0x0
      13'h863: dout  = 8'b00000000; // 2147 :   0 - 0x0
      13'h864: dout  = 8'b11000000; // 2148 : 192 - 0xc0
      13'h865: dout  = 8'b11110000; // 2149 : 240 - 0xf0
      13'h866: dout  = 8'b11111000; // 2150 : 248 - 0xf8
      13'h867: dout  = 8'b11111000; // 2151 : 248 - 0xf8
      13'h868: dout  = 8'b00000000; // 2152 :   0 - 0x0
      13'h869: dout  = 8'b00000000; // 2153 :   0 - 0x0
      13'h86A: dout  = 8'b00000000; // 2154 :   0 - 0x0
      13'h86B: dout  = 8'b11000000; // 2155 : 192 - 0xc0
      13'h86C: dout  = 8'b00110000; // 2156 :  48 - 0x30
      13'h86D: dout  = 8'b00001000; // 2157 :   8 - 0x8
      13'h86E: dout  = 8'b01000100; // 2158 :  68 - 0x44
      13'h86F: dout  = 8'b00000100; // 2159 :   4 - 0x4
      13'h870: dout  = 8'b11111000; // 2160 : 248 - 0xf8 -- Sprite 0x87
      13'h871: dout  = 8'b11111000; // 2161 : 248 - 0xf8
      13'h872: dout  = 8'b11110000; // 2162 : 240 - 0xf0
      13'h873: dout  = 8'b11000000; // 2163 : 192 - 0xc0
      13'h874: dout  = 8'b00000000; // 2164 :   0 - 0x0
      13'h875: dout  = 8'b00000000; // 2165 :   0 - 0x0
      13'h876: dout  = 8'b00000000; // 2166 :   0 - 0x0
      13'h877: dout  = 8'b00000000; // 2167 :   0 - 0x0
      13'h878: dout  = 8'b10000100; // 2168 : 132 - 0x84
      13'h879: dout  = 8'b11000100; // 2169 : 196 - 0xc4
      13'h87A: dout  = 8'b00001000; // 2170 :   8 - 0x8
      13'h87B: dout  = 8'b00110000; // 2171 :  48 - 0x30
      13'h87C: dout  = 8'b11000000; // 2172 : 192 - 0xc0
      13'h87D: dout  = 8'b00000000; // 2173 :   0 - 0x0
      13'h87E: dout  = 8'b00000000; // 2174 :   0 - 0x0
      13'h87F: dout  = 8'b00000000; // 2175 :   0 - 0x0
      13'h880: dout  = 8'b00000000; // 2176 :   0 - 0x0 -- Sprite 0x88
      13'h881: dout  = 8'b00000000; // 2177 :   0 - 0x0
      13'h882: dout  = 8'b00000000; // 2178 :   0 - 0x0
      13'h883: dout  = 8'b00000000; // 2179 :   0 - 0x0
      13'h884: dout  = 8'b00000011; // 2180 :   3 - 0x3
      13'h885: dout  = 8'b00001111; // 2181 :  15 - 0xf
      13'h886: dout  = 8'b00011111; // 2182 :  31 - 0x1f
      13'h887: dout  = 8'b00011111; // 2183 :  31 - 0x1f
      13'h888: dout  = 8'b00000000; // 2184 :   0 - 0x0
      13'h889: dout  = 8'b00000000; // 2185 :   0 - 0x0
      13'h88A: dout  = 8'b00000000; // 2186 :   0 - 0x0
      13'h88B: dout  = 8'b00000011; // 2187 :   3 - 0x3
      13'h88C: dout  = 8'b00001100; // 2188 :  12 - 0xc
      13'h88D: dout  = 8'b00010000; // 2189 :  16 - 0x10
      13'h88E: dout  = 8'b00100000; // 2190 :  32 - 0x20
      13'h88F: dout  = 8'b00100001; // 2191 :  33 - 0x21
      13'h890: dout  = 8'b00011111; // 2192 :  31 - 0x1f -- Sprite 0x89
      13'h891: dout  = 8'b00011111; // 2193 :  31 - 0x1f
      13'h892: dout  = 8'b00001111; // 2194 :  15 - 0xf
      13'h893: dout  = 8'b00000011; // 2195 :   3 - 0x3
      13'h894: dout  = 8'b00000000; // 2196 :   0 - 0x0
      13'h895: dout  = 8'b00000000; // 2197 :   0 - 0x0
      13'h896: dout  = 8'b00000000; // 2198 :   0 - 0x0
      13'h897: dout  = 8'b00000000; // 2199 :   0 - 0x0
      13'h898: dout  = 8'b00100011; // 2200 :  35 - 0x23
      13'h899: dout  = 8'b00100110; // 2201 :  38 - 0x26
      13'h89A: dout  = 8'b00010000; // 2202 :  16 - 0x10
      13'h89B: dout  = 8'b00001100; // 2203 :  12 - 0xc
      13'h89C: dout  = 8'b00000011; // 2204 :   3 - 0x3
      13'h89D: dout  = 8'b00000000; // 2205 :   0 - 0x0
      13'h89E: dout  = 8'b00000000; // 2206 :   0 - 0x0
      13'h89F: dout  = 8'b00000000; // 2207 :   0 - 0x0
      13'h8A0: dout  = 8'b00000000; // 2208 :   0 - 0x0 -- Sprite 0x8a
      13'h8A1: dout  = 8'b00000000; // 2209 :   0 - 0x0
      13'h8A2: dout  = 8'b00000000; // 2210 :   0 - 0x0
      13'h8A3: dout  = 8'b00000000; // 2211 :   0 - 0x0
      13'h8A4: dout  = 8'b11000000; // 2212 : 192 - 0xc0
      13'h8A5: dout  = 8'b11110000; // 2213 : 240 - 0xf0
      13'h8A6: dout  = 8'b11111000; // 2214 : 248 - 0xf8
      13'h8A7: dout  = 8'b11111000; // 2215 : 248 - 0xf8
      13'h8A8: dout  = 8'b00000000; // 2216 :   0 - 0x0
      13'h8A9: dout  = 8'b00000000; // 2217 :   0 - 0x0
      13'h8AA: dout  = 8'b00000000; // 2218 :   0 - 0x0
      13'h8AB: dout  = 8'b11000000; // 2219 : 192 - 0xc0
      13'h8AC: dout  = 8'b00110000; // 2220 :  48 - 0x30
      13'h8AD: dout  = 8'b00001000; // 2221 :   8 - 0x8
      13'h8AE: dout  = 8'b11000100; // 2222 : 196 - 0xc4
      13'h8AF: dout  = 8'b10000100; // 2223 : 132 - 0x84
      13'h8B0: dout  = 8'b11111000; // 2224 : 248 - 0xf8 -- Sprite 0x8b
      13'h8B1: dout  = 8'b11111000; // 2225 : 248 - 0xf8
      13'h8B2: dout  = 8'b11110000; // 2226 : 240 - 0xf0
      13'h8B3: dout  = 8'b11000000; // 2227 : 192 - 0xc0
      13'h8B4: dout  = 8'b00000000; // 2228 :   0 - 0x0
      13'h8B5: dout  = 8'b00000000; // 2229 :   0 - 0x0
      13'h8B6: dout  = 8'b00000000; // 2230 :   0 - 0x0
      13'h8B7: dout  = 8'b00000000; // 2231 :   0 - 0x0
      13'h8B8: dout  = 8'b00000100; // 2232 :   4 - 0x4
      13'h8B9: dout  = 8'b01000100; // 2233 :  68 - 0x44
      13'h8BA: dout  = 8'b00001000; // 2234 :   8 - 0x8
      13'h8BB: dout  = 8'b00110000; // 2235 :  48 - 0x30
      13'h8BC: dout  = 8'b11000000; // 2236 : 192 - 0xc0
      13'h8BD: dout  = 8'b00000000; // 2237 :   0 - 0x0
      13'h8BE: dout  = 8'b00000000; // 2238 :   0 - 0x0
      13'h8BF: dout  = 8'b00000000; // 2239 :   0 - 0x0
      13'h8C0: dout  = 8'b00000000; // 2240 :   0 - 0x0 -- Sprite 0x8c
      13'h8C1: dout  = 8'b00000000; // 2241 :   0 - 0x0
      13'h8C2: dout  = 8'b00000000; // 2242 :   0 - 0x0
      13'h8C3: dout  = 8'b00000000; // 2243 :   0 - 0x0
      13'h8C4: dout  = 8'b00000011; // 2244 :   3 - 0x3
      13'h8C5: dout  = 8'b00001111; // 2245 :  15 - 0xf
      13'h8C6: dout  = 8'b00011111; // 2246 :  31 - 0x1f
      13'h8C7: dout  = 8'b00011111; // 2247 :  31 - 0x1f
      13'h8C8: dout  = 8'b00000000; // 2248 :   0 - 0x0
      13'h8C9: dout  = 8'b00000000; // 2249 :   0 - 0x0
      13'h8CA: dout  = 8'b00000000; // 2250 :   0 - 0x0
      13'h8CB: dout  = 8'b00000011; // 2251 :   3 - 0x3
      13'h8CC: dout  = 8'b00001100; // 2252 :  12 - 0xc
      13'h8CD: dout  = 8'b00010000; // 2253 :  16 - 0x10
      13'h8CE: dout  = 8'b00100011; // 2254 :  35 - 0x23
      13'h8CF: dout  = 8'b00100001; // 2255 :  33 - 0x21
      13'h8D0: dout  = 8'b00011111; // 2256 :  31 - 0x1f -- Sprite 0x8d
      13'h8D1: dout  = 8'b00011111; // 2257 :  31 - 0x1f
      13'h8D2: dout  = 8'b00001111; // 2258 :  15 - 0xf
      13'h8D3: dout  = 8'b00000011; // 2259 :   3 - 0x3
      13'h8D4: dout  = 8'b00000000; // 2260 :   0 - 0x0
      13'h8D5: dout  = 8'b00000000; // 2261 :   0 - 0x0
      13'h8D6: dout  = 8'b00000000; // 2262 :   0 - 0x0
      13'h8D7: dout  = 8'b00000000; // 2263 :   0 - 0x0
      13'h8D8: dout  = 8'b00100000; // 2264 :  32 - 0x20
      13'h8D9: dout  = 8'b00100010; // 2265 :  34 - 0x22
      13'h8DA: dout  = 8'b00010000; // 2266 :  16 - 0x10
      13'h8DB: dout  = 8'b00001100; // 2267 :  12 - 0xc
      13'h8DC: dout  = 8'b00000011; // 2268 :   3 - 0x3
      13'h8DD: dout  = 8'b00000000; // 2269 :   0 - 0x0
      13'h8DE: dout  = 8'b00000000; // 2270 :   0 - 0x0
      13'h8DF: dout  = 8'b00000000; // 2271 :   0 - 0x0
      13'h8E0: dout  = 8'b00000000; // 2272 :   0 - 0x0 -- Sprite 0x8e
      13'h8E1: dout  = 8'b00000000; // 2273 :   0 - 0x0
      13'h8E2: dout  = 8'b00000000; // 2274 :   0 - 0x0
      13'h8E3: dout  = 8'b00000000; // 2275 :   0 - 0x0
      13'h8E4: dout  = 8'b11000000; // 2276 : 192 - 0xc0
      13'h8E5: dout  = 8'b11110000; // 2277 : 240 - 0xf0
      13'h8E6: dout  = 8'b11111000; // 2278 : 248 - 0xf8
      13'h8E7: dout  = 8'b11111000; // 2279 : 248 - 0xf8
      13'h8E8: dout  = 8'b00000000; // 2280 :   0 - 0x0
      13'h8E9: dout  = 8'b00000000; // 2281 :   0 - 0x0
      13'h8EA: dout  = 8'b00000000; // 2282 :   0 - 0x0
      13'h8EB: dout  = 8'b11000000; // 2283 : 192 - 0xc0
      13'h8EC: dout  = 8'b00110000; // 2284 :  48 - 0x30
      13'h8ED: dout  = 8'b00001000; // 2285 :   8 - 0x8
      13'h8EE: dout  = 8'b00000100; // 2286 :   4 - 0x4
      13'h8EF: dout  = 8'b10000100; // 2287 : 132 - 0x84
      13'h8F0: dout  = 8'b11111000; // 2288 : 248 - 0xf8 -- Sprite 0x8f
      13'h8F1: dout  = 8'b11111000; // 2289 : 248 - 0xf8
      13'h8F2: dout  = 8'b11110000; // 2290 : 240 - 0xf0
      13'h8F3: dout  = 8'b11000000; // 2291 : 192 - 0xc0
      13'h8F4: dout  = 8'b00000000; // 2292 :   0 - 0x0
      13'h8F5: dout  = 8'b00000000; // 2293 :   0 - 0x0
      13'h8F6: dout  = 8'b00000000; // 2294 :   0 - 0x0
      13'h8F7: dout  = 8'b00000000; // 2295 :   0 - 0x0
      13'h8F8: dout  = 8'b11000100; // 2296 : 196 - 0xc4
      13'h8F9: dout  = 8'b01100100; // 2297 : 100 - 0x64
      13'h8FA: dout  = 8'b00001000; // 2298 :   8 - 0x8
      13'h8FB: dout  = 8'b00110000; // 2299 :  48 - 0x30
      13'h8FC: dout  = 8'b11000000; // 2300 : 192 - 0xc0
      13'h8FD: dout  = 8'b00000000; // 2301 :   0 - 0x0
      13'h8FE: dout  = 8'b00000000; // 2302 :   0 - 0x0
      13'h8FF: dout  = 8'b00000000; // 2303 :   0 - 0x0
      13'h900: dout  = 8'b00000000; // 2304 :   0 - 0x0 -- Sprite 0x90
      13'h901: dout  = 8'b00000000; // 2305 :   0 - 0x0
      13'h902: dout  = 8'b00000000; // 2306 :   0 - 0x0
      13'h903: dout  = 8'b00001111; // 2307 :  15 - 0xf
      13'h904: dout  = 8'b00110000; // 2308 :  48 - 0x30
      13'h905: dout  = 8'b01100000; // 2309 :  96 - 0x60
      13'h906: dout  = 8'b00111111; // 2310 :  63 - 0x3f
      13'h907: dout  = 8'b01111111; // 2311 : 127 - 0x7f
      13'h908: dout  = 8'b00000000; // 2312 :   0 - 0x0
      13'h909: dout  = 8'b00000000; // 2313 :   0 - 0x0
      13'h90A: dout  = 8'b00000000; // 2314 :   0 - 0x0
      13'h90B: dout  = 8'b00000000; // 2315 :   0 - 0x0
      13'h90C: dout  = 8'b00101111; // 2316 :  47 - 0x2f
      13'h90D: dout  = 8'b00111111; // 2317 :  63 - 0x3f
      13'h90E: dout  = 8'b01100000; // 2318 :  96 - 0x60
      13'h90F: dout  = 8'b00100000; // 2319 :  32 - 0x20
      13'h910: dout  = 8'b01111111; // 2320 : 127 - 0x7f -- Sprite 0x91
      13'h911: dout  = 8'b00111111; // 2321 :  63 - 0x3f
      13'h912: dout  = 8'b01100000; // 2322 :  96 - 0x60
      13'h913: dout  = 8'b00110000; // 2323 :  48 - 0x30
      13'h914: dout  = 8'b00001111; // 2324 :  15 - 0xf
      13'h915: dout  = 8'b00000000; // 2325 :   0 - 0x0
      13'h916: dout  = 8'b00000000; // 2326 :   0 - 0x0
      13'h917: dout  = 8'b00000000; // 2327 :   0 - 0x0
      13'h918: dout  = 8'b00100000; // 2328 :  32 - 0x20
      13'h919: dout  = 8'b01100000; // 2329 :  96 - 0x60
      13'h91A: dout  = 8'b00111111; // 2330 :  63 - 0x3f
      13'h91B: dout  = 8'b00101111; // 2331 :  47 - 0x2f
      13'h91C: dout  = 8'b00000000; // 2332 :   0 - 0x0
      13'h91D: dout  = 8'b00000000; // 2333 :   0 - 0x0
      13'h91E: dout  = 8'b00000000; // 2334 :   0 - 0x0
      13'h91F: dout  = 8'b00000000; // 2335 :   0 - 0x0
      13'h920: dout  = 8'b00000000; // 2336 :   0 - 0x0 -- Sprite 0x92
      13'h921: dout  = 8'b00000000; // 2337 :   0 - 0x0
      13'h922: dout  = 8'b00000000; // 2338 :   0 - 0x0
      13'h923: dout  = 8'b11111000; // 2339 : 248 - 0xf8
      13'h924: dout  = 8'b00000110; // 2340 :   6 - 0x6
      13'h925: dout  = 8'b00000011; // 2341 :   3 - 0x3
      13'h926: dout  = 8'b11111110; // 2342 : 254 - 0xfe
      13'h927: dout  = 8'b11111111; // 2343 : 255 - 0xff
      13'h928: dout  = 8'b00000000; // 2344 :   0 - 0x0
      13'h929: dout  = 8'b00000000; // 2345 :   0 - 0x0
      13'h92A: dout  = 8'b00000000; // 2346 :   0 - 0x0
      13'h92B: dout  = 8'b00000000; // 2347 :   0 - 0x0
      13'h92C: dout  = 8'b11111010; // 2348 : 250 - 0xfa
      13'h92D: dout  = 8'b11111110; // 2349 : 254 - 0xfe
      13'h92E: dout  = 8'b00000011; // 2350 :   3 - 0x3
      13'h92F: dout  = 8'b00000010; // 2351 :   2 - 0x2
      13'h930: dout  = 8'b11111111; // 2352 : 255 - 0xff -- Sprite 0x93
      13'h931: dout  = 8'b11111110; // 2353 : 254 - 0xfe
      13'h932: dout  = 8'b00000011; // 2354 :   3 - 0x3
      13'h933: dout  = 8'b00000110; // 2355 :   6 - 0x6
      13'h934: dout  = 8'b11111000; // 2356 : 248 - 0xf8
      13'h935: dout  = 8'b00000000; // 2357 :   0 - 0x0
      13'h936: dout  = 8'b00000000; // 2358 :   0 - 0x0
      13'h937: dout  = 8'b00000000; // 2359 :   0 - 0x0
      13'h938: dout  = 8'b00000010; // 2360 :   2 - 0x2
      13'h939: dout  = 8'b00000011; // 2361 :   3 - 0x3
      13'h93A: dout  = 8'b11111110; // 2362 : 254 - 0xfe
      13'h93B: dout  = 8'b11111010; // 2363 : 250 - 0xfa
      13'h93C: dout  = 8'b00000000; // 2364 :   0 - 0x0
      13'h93D: dout  = 8'b00000000; // 2365 :   0 - 0x0
      13'h93E: dout  = 8'b00000000; // 2366 :   0 - 0x0
      13'h93F: dout  = 8'b00000000; // 2367 :   0 - 0x0
      13'h940: dout  = 8'b00000000; // 2368 :   0 - 0x0 -- Sprite 0x94
      13'h941: dout  = 8'b00000000; // 2369 :   0 - 0x0
      13'h942: dout  = 8'b00000000; // 2370 :   0 - 0x0
      13'h943: dout  = 8'b00000000; // 2371 :   0 - 0x0
      13'h944: dout  = 8'b00101111; // 2372 :  47 - 0x2f
      13'h945: dout  = 8'b00111111; // 2373 :  63 - 0x3f
      13'h946: dout  = 8'b01100000; // 2374 :  96 - 0x60
      13'h947: dout  = 8'b00100000; // 2375 :  32 - 0x20
      13'h948: dout  = 8'b00000000; // 2376 :   0 - 0x0
      13'h949: dout  = 8'b00000000; // 2377 :   0 - 0x0
      13'h94A: dout  = 8'b00000000; // 2378 :   0 - 0x0
      13'h94B: dout  = 8'b00001111; // 2379 :  15 - 0xf
      13'h94C: dout  = 8'b00110000; // 2380 :  48 - 0x30
      13'h94D: dout  = 8'b01100000; // 2381 :  96 - 0x60
      13'h94E: dout  = 8'b00111111; // 2382 :  63 - 0x3f
      13'h94F: dout  = 8'b01111111; // 2383 : 127 - 0x7f
      13'h950: dout  = 8'b00100000; // 2384 :  32 - 0x20 -- Sprite 0x95
      13'h951: dout  = 8'b01100000; // 2385 :  96 - 0x60
      13'h952: dout  = 8'b00111111; // 2386 :  63 - 0x3f
      13'h953: dout  = 8'b00101111; // 2387 :  47 - 0x2f
      13'h954: dout  = 8'b00000000; // 2388 :   0 - 0x0
      13'h955: dout  = 8'b00000000; // 2389 :   0 - 0x0
      13'h956: dout  = 8'b00000000; // 2390 :   0 - 0x0
      13'h957: dout  = 8'b00000000; // 2391 :   0 - 0x0
      13'h958: dout  = 8'b01111111; // 2392 : 127 - 0x7f
      13'h959: dout  = 8'b00111111; // 2393 :  63 - 0x3f
      13'h95A: dout  = 8'b01100000; // 2394 :  96 - 0x60
      13'h95B: dout  = 8'b00110000; // 2395 :  48 - 0x30
      13'h95C: dout  = 8'b00001111; // 2396 :  15 - 0xf
      13'h95D: dout  = 8'b00000000; // 2397 :   0 - 0x0
      13'h95E: dout  = 8'b00000000; // 2398 :   0 - 0x0
      13'h95F: dout  = 8'b00000000; // 2399 :   0 - 0x0
      13'h960: dout  = 8'b00000000; // 2400 :   0 - 0x0 -- Sprite 0x96
      13'h961: dout  = 8'b00000000; // 2401 :   0 - 0x0
      13'h962: dout  = 8'b00000000; // 2402 :   0 - 0x0
      13'h963: dout  = 8'b00000000; // 2403 :   0 - 0x0
      13'h964: dout  = 8'b11111010; // 2404 : 250 - 0xfa
      13'h965: dout  = 8'b11111110; // 2405 : 254 - 0xfe
      13'h966: dout  = 8'b00000011; // 2406 :   3 - 0x3
      13'h967: dout  = 8'b00000010; // 2407 :   2 - 0x2
      13'h968: dout  = 8'b00000000; // 2408 :   0 - 0x0
      13'h969: dout  = 8'b00000000; // 2409 :   0 - 0x0
      13'h96A: dout  = 8'b00000000; // 2410 :   0 - 0x0
      13'h96B: dout  = 8'b11111000; // 2411 : 248 - 0xf8
      13'h96C: dout  = 8'b00000110; // 2412 :   6 - 0x6
      13'h96D: dout  = 8'b00000011; // 2413 :   3 - 0x3
      13'h96E: dout  = 8'b11111110; // 2414 : 254 - 0xfe
      13'h96F: dout  = 8'b11111111; // 2415 : 255 - 0xff
      13'h970: dout  = 8'b00000010; // 2416 :   2 - 0x2 -- Sprite 0x97
      13'h971: dout  = 8'b00000011; // 2417 :   3 - 0x3
      13'h972: dout  = 8'b11111110; // 2418 : 254 - 0xfe
      13'h973: dout  = 8'b11111010; // 2419 : 250 - 0xfa
      13'h974: dout  = 8'b00000000; // 2420 :   0 - 0x0
      13'h975: dout  = 8'b00000000; // 2421 :   0 - 0x0
      13'h976: dout  = 8'b00000000; // 2422 :   0 - 0x0
      13'h977: dout  = 8'b00000000; // 2423 :   0 - 0x0
      13'h978: dout  = 8'b11111111; // 2424 : 255 - 0xff
      13'h979: dout  = 8'b11111110; // 2425 : 254 - 0xfe
      13'h97A: dout  = 8'b00000011; // 2426 :   3 - 0x3
      13'h97B: dout  = 8'b00000110; // 2427 :   6 - 0x6
      13'h97C: dout  = 8'b11111000; // 2428 : 248 - 0xf8
      13'h97D: dout  = 8'b00000000; // 2429 :   0 - 0x0
      13'h97E: dout  = 8'b00000000; // 2430 :   0 - 0x0
      13'h97F: dout  = 8'b00000000; // 2431 :   0 - 0x0
      13'h980: dout  = 8'b00000000; // 2432 :   0 - 0x0 -- Sprite 0x98
      13'h981: dout  = 8'b01000100; // 2433 :  68 - 0x44
      13'h982: dout  = 8'b00000000; // 2434 :   0 - 0x0
      13'h983: dout  = 8'b01000001; // 2435 :  65 - 0x41
      13'h984: dout  = 8'b00100000; // 2436 :  32 - 0x20
      13'h985: dout  = 8'b01001011; // 2437 :  75 - 0x4b
      13'h986: dout  = 8'b00100111; // 2438 :  39 - 0x27
      13'h987: dout  = 8'b00011111; // 2439 :  31 - 0x1f
      13'h988: dout  = 8'b00000000; // 2440 :   0 - 0x0
      13'h989: dout  = 8'b00000000; // 2441 :   0 - 0x0
      13'h98A: dout  = 8'b00000000; // 2442 :   0 - 0x0
      13'h98B: dout  = 8'b01000000; // 2443 :  64 - 0x40
      13'h98C: dout  = 8'b00100000; // 2444 :  32 - 0x20
      13'h98D: dout  = 8'b00000000; // 2445 :   0 - 0x0
      13'h98E: dout  = 8'b00000000; // 2446 :   0 - 0x0
      13'h98F: dout  = 8'b00000001; // 2447 :   1 - 0x1
      13'h990: dout  = 8'b00001111; // 2448 :  15 - 0xf -- Sprite 0x99
      13'h991: dout  = 8'b00011110; // 2449 :  30 - 0x1e
      13'h992: dout  = 8'b00011111; // 2450 :  31 - 0x1f
      13'h993: dout  = 8'b00011111; // 2451 :  31 - 0x1f
      13'h994: dout  = 8'b00011111; // 2452 :  31 - 0x1f
      13'h995: dout  = 8'b00001111; // 2453 :  15 - 0xf
      13'h996: dout  = 8'b00001111; // 2454 :  15 - 0xf
      13'h997: dout  = 8'b00000011; // 2455 :   3 - 0x3
      13'h998: dout  = 8'b00000011; // 2456 :   3 - 0x3
      13'h999: dout  = 8'b00000111; // 2457 :   7 - 0x7
      13'h99A: dout  = 8'b00000110; // 2458 :   6 - 0x6
      13'h99B: dout  = 8'b00000110; // 2459 :   6 - 0x6
      13'h99C: dout  = 8'b00000111; // 2460 :   7 - 0x7
      13'h99D: dout  = 8'b00000011; // 2461 :   3 - 0x3
      13'h99E: dout  = 8'b00000000; // 2462 :   0 - 0x0
      13'h99F: dout  = 8'b00000000; // 2463 :   0 - 0x0
      13'h9A0: dout  = 8'b00000000; // 2464 :   0 - 0x0 -- Sprite 0x9a
      13'h9A1: dout  = 8'b00100000; // 2465 :  32 - 0x20
      13'h9A2: dout  = 8'b01010000; // 2466 :  80 - 0x50
      13'h9A3: dout  = 8'b00100000; // 2467 :  32 - 0x20
      13'h9A4: dout  = 8'b01100000; // 2468 :  96 - 0x60
      13'h9A5: dout  = 8'b01001000; // 2469 :  72 - 0x48
      13'h9A6: dout  = 8'b11100000; // 2470 : 224 - 0xe0
      13'h9A7: dout  = 8'b11110000; // 2471 : 240 - 0xf0
      13'h9A8: dout  = 8'b00000000; // 2472 :   0 - 0x0
      13'h9A9: dout  = 8'b00000000; // 2473 :   0 - 0x0
      13'h9AA: dout  = 8'b01000000; // 2474 :  64 - 0x40
      13'h9AB: dout  = 8'b00000000; // 2475 :   0 - 0x0
      13'h9AC: dout  = 8'b00000000; // 2476 :   0 - 0x0
      13'h9AD: dout  = 8'b00001000; // 2477 :   8 - 0x8
      13'h9AE: dout  = 8'b00000000; // 2478 :   0 - 0x0
      13'h9AF: dout  = 8'b01000000; // 2479 :  64 - 0x40
      13'h9B0: dout  = 8'b11111000; // 2480 : 248 - 0xf8 -- Sprite 0x9b
      13'h9B1: dout  = 8'b01111000; // 2481 : 120 - 0x78
      13'h9B2: dout  = 8'b00111100; // 2482 :  60 - 0x3c
      13'h9B3: dout  = 8'b00111100; // 2483 :  60 - 0x3c
      13'h9B4: dout  = 8'b00111100; // 2484 :  60 - 0x3c
      13'h9B5: dout  = 8'b11111100; // 2485 : 252 - 0xfc
      13'h9B6: dout  = 8'b11111000; // 2486 : 248 - 0xf8
      13'h9B7: dout  = 8'b11100000; // 2487 : 224 - 0xe0
      13'h9B8: dout  = 8'b11100000; // 2488 : 224 - 0xe0
      13'h9B9: dout  = 8'b11110000; // 2489 : 240 - 0xf0
      13'h9BA: dout  = 8'b11010000; // 2490 : 208 - 0xd0
      13'h9BB: dout  = 8'b11010000; // 2491 : 208 - 0xd0
      13'h9BC: dout  = 8'b11110000; // 2492 : 240 - 0xf0
      13'h9BD: dout  = 8'b11100000; // 2493 : 224 - 0xe0
      13'h9BE: dout  = 8'b00000000; // 2494 :   0 - 0x0
      13'h9BF: dout  = 8'b00000000; // 2495 :   0 - 0x0
      13'h9C0: dout  = 8'b00010000; // 2496 :  16 - 0x10 -- Sprite 0x9c
      13'h9C1: dout  = 8'b00000001; // 2497 :   1 - 0x1
      13'h9C2: dout  = 8'b00101010; // 2498 :  42 - 0x2a
      13'h9C3: dout  = 8'b00001100; // 2499 :  12 - 0xc
      13'h9C4: dout  = 8'b10100110; // 2500 : 166 - 0xa6
      13'h9C5: dout  = 8'b00010111; // 2501 :  23 - 0x17
      13'h9C6: dout  = 8'b00011111; // 2502 :  31 - 0x1f
      13'h9C7: dout  = 8'b00011111; // 2503 :  31 - 0x1f
      13'h9C8: dout  = 8'b00000000; // 2504 :   0 - 0x0
      13'h9C9: dout  = 8'b00000000; // 2505 :   0 - 0x0
      13'h9CA: dout  = 8'b00000010; // 2506 :   2 - 0x2
      13'h9CB: dout  = 8'b00000000; // 2507 :   0 - 0x0
      13'h9CC: dout  = 8'b10000000; // 2508 : 128 - 0x80
      13'h9CD: dout  = 8'b00000000; // 2509 :   0 - 0x0
      13'h9CE: dout  = 8'b00000011; // 2510 :   3 - 0x3
      13'h9CF: dout  = 8'b00000111; // 2511 :   7 - 0x7
      13'h9D0: dout  = 8'b01011110; // 2512 :  94 - 0x5e -- Sprite 0x9d
      13'h9D1: dout  = 8'b00111100; // 2513 :  60 - 0x3c
      13'h9D2: dout  = 8'b00111101; // 2514 :  61 - 0x3d
      13'h9D3: dout  = 8'b00111101; // 2515 :  61 - 0x3d
      13'h9D4: dout  = 8'b00111110; // 2516 :  62 - 0x3e
      13'h9D5: dout  = 8'b00011111; // 2517 :  31 - 0x1f
      13'h9D6: dout  = 8'b00001111; // 2518 :  15 - 0xf
      13'h9D7: dout  = 8'b00000111; // 2519 :   7 - 0x7
      13'h9D8: dout  = 8'b00000111; // 2520 :   7 - 0x7
      13'h9D9: dout  = 8'b00001111; // 2521 :  15 - 0xf
      13'h9DA: dout  = 8'b00001110; // 2522 :  14 - 0xe
      13'h9DB: dout  = 8'b00001110; // 2523 :  14 - 0xe
      13'h9DC: dout  = 8'b00001111; // 2524 :  15 - 0xf
      13'h9DD: dout  = 8'b00000111; // 2525 :   7 - 0x7
      13'h9DE: dout  = 8'b00000011; // 2526 :   3 - 0x3
      13'h9DF: dout  = 8'b00000000; // 2527 :   0 - 0x0
      13'h9E0: dout  = 8'b00000000; // 2528 :   0 - 0x0 -- Sprite 0x9e
      13'h9E1: dout  = 8'b00000000; // 2529 :   0 - 0x0
      13'h9E2: dout  = 8'b10000000; // 2530 : 128 - 0x80
      13'h9E3: dout  = 8'b11001000; // 2531 : 200 - 0xc8
      13'h9E4: dout  = 8'b01100000; // 2532 :  96 - 0x60
      13'h9E5: dout  = 8'b11100000; // 2533 : 224 - 0xe0
      13'h9E6: dout  = 8'b11110100; // 2534 : 244 - 0xf4
      13'h9E7: dout  = 8'b11111000; // 2535 : 248 - 0xf8
      13'h9E8: dout  = 8'b00000000; // 2536 :   0 - 0x0
      13'h9E9: dout  = 8'b00000000; // 2537 :   0 - 0x0
      13'h9EA: dout  = 8'b00000000; // 2538 :   0 - 0x0
      13'h9EB: dout  = 8'b00001000; // 2539 :   8 - 0x8
      13'h9EC: dout  = 8'b00000000; // 2540 :   0 - 0x0
      13'h9ED: dout  = 8'b10000000; // 2541 : 128 - 0x80
      13'h9EE: dout  = 8'b00100100; // 2542 :  36 - 0x24
      13'h9EF: dout  = 8'b11000000; // 2543 : 192 - 0xc0
      13'h9F0: dout  = 8'b01111100; // 2544 : 124 - 0x7c -- Sprite 0x9f
      13'h9F1: dout  = 8'b00011100; // 2545 :  28 - 0x1c
      13'h9F2: dout  = 8'b00101110; // 2546 :  46 - 0x2e
      13'h9F3: dout  = 8'b00101110; // 2547 :  46 - 0x2e
      13'h9F4: dout  = 8'b00011110; // 2548 :  30 - 0x1e
      13'h9F5: dout  = 8'b11111100; // 2549 : 252 - 0xfc
      13'h9F6: dout  = 8'b11111000; // 2550 : 248 - 0xf8
      13'h9F7: dout  = 8'b11100000; // 2551 : 224 - 0xe0
      13'h9F8: dout  = 8'b11110000; // 2552 : 240 - 0xf0
      13'h9F9: dout  = 8'b11111000; // 2553 : 248 - 0xf8
      13'h9FA: dout  = 8'b11011000; // 2554 : 216 - 0xd8
      13'h9FB: dout  = 8'b11011000; // 2555 : 216 - 0xd8
      13'h9FC: dout  = 8'b11111000; // 2556 : 248 - 0xf8
      13'h9FD: dout  = 8'b11110000; // 2557 : 240 - 0xf0
      13'h9FE: dout  = 8'b11000000; // 2558 : 192 - 0xc0
      13'h9FF: dout  = 8'b00000000; // 2559 :   0 - 0x0
      13'hA00: dout  = 8'b11111111; // 2560 : 255 - 0xff -- Sprite 0xa0
      13'hA01: dout  = 8'b11111111; // 2561 : 255 - 0xff
      13'hA02: dout  = 8'b00111000; // 2562 :  56 - 0x38
      13'hA03: dout  = 8'b01101100; // 2563 : 108 - 0x6c
      13'hA04: dout  = 8'b11000110; // 2564 : 198 - 0xc6
      13'hA05: dout  = 8'b10000011; // 2565 : 131 - 0x83
      13'hA06: dout  = 8'b11111111; // 2566 : 255 - 0xff
      13'hA07: dout  = 8'b11111111; // 2567 : 255 - 0xff
      13'hA08: dout  = 8'b11111111; // 2568 : 255 - 0xff
      13'hA09: dout  = 8'b11111111; // 2569 : 255 - 0xff
      13'hA0A: dout  = 8'b00111000; // 2570 :  56 - 0x38
      13'hA0B: dout  = 8'b01101100; // 2571 : 108 - 0x6c
      13'hA0C: dout  = 8'b11000110; // 2572 : 198 - 0xc6
      13'hA0D: dout  = 8'b10000011; // 2573 : 131 - 0x83
      13'hA0E: dout  = 8'b11111111; // 2574 : 255 - 0xff
      13'hA0F: dout  = 8'b11111111; // 2575 : 255 - 0xff
      13'hA10: dout  = 8'b11111111; // 2576 : 255 - 0xff -- Sprite 0xa1
      13'hA11: dout  = 8'b11111111; // 2577 : 255 - 0xff
      13'hA12: dout  = 8'b00111000; // 2578 :  56 - 0x38
      13'hA13: dout  = 8'b01101100; // 2579 : 108 - 0x6c
      13'hA14: dout  = 8'b11000110; // 2580 : 198 - 0xc6
      13'hA15: dout  = 8'b10000011; // 2581 : 131 - 0x83
      13'hA16: dout  = 8'b11111111; // 2582 : 255 - 0xff
      13'hA17: dout  = 8'b11111111; // 2583 : 255 - 0xff
      13'hA18: dout  = 8'b11111111; // 2584 : 255 - 0xff
      13'hA19: dout  = 8'b11111111; // 2585 : 255 - 0xff
      13'hA1A: dout  = 8'b00111000; // 2586 :  56 - 0x38
      13'hA1B: dout  = 8'b01101100; // 2587 : 108 - 0x6c
      13'hA1C: dout  = 8'b11000110; // 2588 : 198 - 0xc6
      13'hA1D: dout  = 8'b10000011; // 2589 : 131 - 0x83
      13'hA1E: dout  = 8'b11111111; // 2590 : 255 - 0xff
      13'hA1F: dout  = 8'b11111111; // 2591 : 255 - 0xff
      13'hA20: dout  = 8'b10010010; // 2592 : 146 - 0x92 -- Sprite 0xa2
      13'hA21: dout  = 8'b01010100; // 2593 :  84 - 0x54
      13'hA22: dout  = 8'b00111000; // 2594 :  56 - 0x38
      13'hA23: dout  = 8'b11111110; // 2595 : 254 - 0xfe
      13'hA24: dout  = 8'b00111000; // 2596 :  56 - 0x38
      13'hA25: dout  = 8'b01010100; // 2597 :  84 - 0x54
      13'hA26: dout  = 8'b10010010; // 2598 : 146 - 0x92
      13'hA27: dout  = 8'b00000000; // 2599 :   0 - 0x0
      13'hA28: dout  = 8'b00000000; // 2600 :   0 - 0x0
      13'hA29: dout  = 8'b00000000; // 2601 :   0 - 0x0
      13'hA2A: dout  = 8'b00000000; // 2602 :   0 - 0x0
      13'hA2B: dout  = 8'b00000000; // 2603 :   0 - 0x0
      13'hA2C: dout  = 8'b00000000; // 2604 :   0 - 0x0
      13'hA2D: dout  = 8'b00000000; // 2605 :   0 - 0x0
      13'hA2E: dout  = 8'b00000000; // 2606 :   0 - 0x0
      13'hA2F: dout  = 8'b00000000; // 2607 :   0 - 0x0
      13'hA30: dout  = 8'b11111111; // 2608 : 255 - 0xff -- Sprite 0xa3
      13'hA31: dout  = 8'b11111111; // 2609 : 255 - 0xff
      13'hA32: dout  = 8'b11111111; // 2610 : 255 - 0xff
      13'hA33: dout  = 8'b11111111; // 2611 : 255 - 0xff
      13'hA34: dout  = 8'b11111111; // 2612 : 255 - 0xff
      13'hA35: dout  = 8'b11111111; // 2613 : 255 - 0xff
      13'hA36: dout  = 8'b11111111; // 2614 : 255 - 0xff
      13'hA37: dout  = 8'b11111111; // 2615 : 255 - 0xff
      13'hA38: dout  = 8'b11111111; // 2616 : 255 - 0xff
      13'hA39: dout  = 8'b11111111; // 2617 : 255 - 0xff
      13'hA3A: dout  = 8'b11111111; // 2618 : 255 - 0xff
      13'hA3B: dout  = 8'b11111111; // 2619 : 255 - 0xff
      13'hA3C: dout  = 8'b11111111; // 2620 : 255 - 0xff
      13'hA3D: dout  = 8'b11111111; // 2621 : 255 - 0xff
      13'hA3E: dout  = 8'b11111111; // 2622 : 255 - 0xff
      13'hA3F: dout  = 8'b11111111; // 2623 : 255 - 0xff
      13'hA40: dout  = 8'b11111111; // 2624 : 255 - 0xff -- Sprite 0xa4
      13'hA41: dout  = 8'b11111111; // 2625 : 255 - 0xff
      13'hA42: dout  = 8'b11111111; // 2626 : 255 - 0xff
      13'hA43: dout  = 8'b11111111; // 2627 : 255 - 0xff
      13'hA44: dout  = 8'b11111111; // 2628 : 255 - 0xff
      13'hA45: dout  = 8'b11111111; // 2629 : 255 - 0xff
      13'hA46: dout  = 8'b11111111; // 2630 : 255 - 0xff
      13'hA47: dout  = 8'b11111111; // 2631 : 255 - 0xff
      13'hA48: dout  = 8'b11111111; // 2632 : 255 - 0xff
      13'hA49: dout  = 8'b11111111; // 2633 : 255 - 0xff
      13'hA4A: dout  = 8'b11111111; // 2634 : 255 - 0xff
      13'hA4B: dout  = 8'b11111111; // 2635 : 255 - 0xff
      13'hA4C: dout  = 8'b11111111; // 2636 : 255 - 0xff
      13'hA4D: dout  = 8'b11111111; // 2637 : 255 - 0xff
      13'hA4E: dout  = 8'b11111111; // 2638 : 255 - 0xff
      13'hA4F: dout  = 8'b11111111; // 2639 : 255 - 0xff
      13'hA50: dout  = 8'b11111111; // 2640 : 255 - 0xff -- Sprite 0xa5
      13'hA51: dout  = 8'b11111111; // 2641 : 255 - 0xff
      13'hA52: dout  = 8'b11111111; // 2642 : 255 - 0xff
      13'hA53: dout  = 8'b11111111; // 2643 : 255 - 0xff
      13'hA54: dout  = 8'b11111111; // 2644 : 255 - 0xff
      13'hA55: dout  = 8'b11111111; // 2645 : 255 - 0xff
      13'hA56: dout  = 8'b11111111; // 2646 : 255 - 0xff
      13'hA57: dout  = 8'b11111111; // 2647 : 255 - 0xff
      13'hA58: dout  = 8'b11111111; // 2648 : 255 - 0xff
      13'hA59: dout  = 8'b11111111; // 2649 : 255 - 0xff
      13'hA5A: dout  = 8'b11111111; // 2650 : 255 - 0xff
      13'hA5B: dout  = 8'b11111111; // 2651 : 255 - 0xff
      13'hA5C: dout  = 8'b11111111; // 2652 : 255 - 0xff
      13'hA5D: dout  = 8'b11111111; // 2653 : 255 - 0xff
      13'hA5E: dout  = 8'b11111111; // 2654 : 255 - 0xff
      13'hA5F: dout  = 8'b11111111; // 2655 : 255 - 0xff
      13'hA60: dout  = 8'b11111111; // 2656 : 255 - 0xff -- Sprite 0xa6
      13'hA61: dout  = 8'b11111111; // 2657 : 255 - 0xff
      13'hA62: dout  = 8'b11111111; // 2658 : 255 - 0xff
      13'hA63: dout  = 8'b11111111; // 2659 : 255 - 0xff
      13'hA64: dout  = 8'b11111111; // 2660 : 255 - 0xff
      13'hA65: dout  = 8'b11111111; // 2661 : 255 - 0xff
      13'hA66: dout  = 8'b11111111; // 2662 : 255 - 0xff
      13'hA67: dout  = 8'b11111111; // 2663 : 255 - 0xff
      13'hA68: dout  = 8'b11111111; // 2664 : 255 - 0xff
      13'hA69: dout  = 8'b11111111; // 2665 : 255 - 0xff
      13'hA6A: dout  = 8'b11111111; // 2666 : 255 - 0xff
      13'hA6B: dout  = 8'b11111111; // 2667 : 255 - 0xff
      13'hA6C: dout  = 8'b11111111; // 2668 : 255 - 0xff
      13'hA6D: dout  = 8'b11111111; // 2669 : 255 - 0xff
      13'hA6E: dout  = 8'b11111111; // 2670 : 255 - 0xff
      13'hA6F: dout  = 8'b11111111; // 2671 : 255 - 0xff
      13'hA70: dout  = 8'b11111111; // 2672 : 255 - 0xff -- Sprite 0xa7
      13'hA71: dout  = 8'b11111111; // 2673 : 255 - 0xff
      13'hA72: dout  = 8'b11111111; // 2674 : 255 - 0xff
      13'hA73: dout  = 8'b11111111; // 2675 : 255 - 0xff
      13'hA74: dout  = 8'b11111111; // 2676 : 255 - 0xff
      13'hA75: dout  = 8'b11111111; // 2677 : 255 - 0xff
      13'hA76: dout  = 8'b11111111; // 2678 : 255 - 0xff
      13'hA77: dout  = 8'b11111111; // 2679 : 255 - 0xff
      13'hA78: dout  = 8'b11111111; // 2680 : 255 - 0xff
      13'hA79: dout  = 8'b11111111; // 2681 : 255 - 0xff
      13'hA7A: dout  = 8'b11111111; // 2682 : 255 - 0xff
      13'hA7B: dout  = 8'b11111111; // 2683 : 255 - 0xff
      13'hA7C: dout  = 8'b11111111; // 2684 : 255 - 0xff
      13'hA7D: dout  = 8'b11111111; // 2685 : 255 - 0xff
      13'hA7E: dout  = 8'b11111111; // 2686 : 255 - 0xff
      13'hA7F: dout  = 8'b11111111; // 2687 : 255 - 0xff
      13'hA80: dout  = 8'b00000000; // 2688 :   0 - 0x0 -- Sprite 0xa8
      13'hA81: dout  = 8'b00000000; // 2689 :   0 - 0x0
      13'hA82: dout  = 8'b00000000; // 2690 :   0 - 0x0
      13'hA83: dout  = 8'b00000000; // 2691 :   0 - 0x0
      13'hA84: dout  = 8'b00000000; // 2692 :   0 - 0x0
      13'hA85: dout  = 8'b00100011; // 2693 :  35 - 0x23
      13'hA86: dout  = 8'b10010111; // 2694 : 151 - 0x97
      13'hA87: dout  = 8'b00101111; // 2695 :  47 - 0x2f
      13'hA88: dout  = 8'b00000000; // 2696 :   0 - 0x0
      13'hA89: dout  = 8'b00000000; // 2697 :   0 - 0x0
      13'hA8A: dout  = 8'b00000000; // 2698 :   0 - 0x0
      13'hA8B: dout  = 8'b00000000; // 2699 :   0 - 0x0
      13'hA8C: dout  = 8'b00000000; // 2700 :   0 - 0x0
      13'hA8D: dout  = 8'b00000000; // 2701 :   0 - 0x0
      13'hA8E: dout  = 8'b00000001; // 2702 :   1 - 0x1
      13'hA8F: dout  = 8'b00000011; // 2703 :   3 - 0x3
      13'hA90: dout  = 8'b01101110; // 2704 : 110 - 0x6e -- Sprite 0xa9
      13'hA91: dout  = 8'b11101111; // 2705 : 239 - 0xef
      13'hA92: dout  = 8'b11110111; // 2706 : 247 - 0xf7
      13'hA93: dout  = 8'b11111111; // 2707 : 255 - 0xff
      13'hA94: dout  = 8'b01111111; // 2708 : 127 - 0x7f
      13'hA95: dout  = 8'b00111111; // 2709 :  63 - 0x3f
      13'hA96: dout  = 8'b01011111; // 2710 :  95 - 0x5f
      13'hA97: dout  = 8'b00001111; // 2711 :  15 - 0xf
      13'hA98: dout  = 8'b00000111; // 2712 :   7 - 0x7
      13'hA99: dout  = 8'b00000111; // 2713 :   7 - 0x7
      13'hA9A: dout  = 8'b00000011; // 2714 :   3 - 0x3
      13'hA9B: dout  = 8'b00100111; // 2715 :  39 - 0x27
      13'hA9C: dout  = 8'b00011111; // 2716 :  31 - 0x1f
      13'hA9D: dout  = 8'b00000111; // 2717 :   7 - 0x7
      13'hA9E: dout  = 8'b00000000; // 2718 :   0 - 0x0
      13'hA9F: dout  = 8'b00000000; // 2719 :   0 - 0x0
      13'hAA0: dout  = 8'b00000000; // 2720 :   0 - 0x0 -- Sprite 0xaa
      13'hAA1: dout  = 8'b00000000; // 2721 :   0 - 0x0
      13'hAA2: dout  = 8'b00000000; // 2722 :   0 - 0x0
      13'hAA3: dout  = 8'b00000000; // 2723 :   0 - 0x0
      13'hAA4: dout  = 8'b11111000; // 2724 : 248 - 0xf8
      13'hAA5: dout  = 8'b11111100; // 2725 : 252 - 0xfc
      13'hAA6: dout  = 8'b11111110; // 2726 : 254 - 0xfe
      13'hAA7: dout  = 8'b01011110; // 2727 :  94 - 0x5e
      13'hAA8: dout  = 8'b00000000; // 2728 :   0 - 0x0
      13'hAA9: dout  = 8'b00000000; // 2729 :   0 - 0x0
      13'hAAA: dout  = 8'b00000000; // 2730 :   0 - 0x0
      13'hAAB: dout  = 8'b00000000; // 2731 :   0 - 0x0
      13'hAAC: dout  = 8'b00000000; // 2732 :   0 - 0x0
      13'hAAD: dout  = 8'b11110000; // 2733 : 240 - 0xf0
      13'hAAE: dout  = 8'b11111000; // 2734 : 248 - 0xf8
      13'hAAF: dout  = 8'b10101100; // 2735 : 172 - 0xac
      13'hAB0: dout  = 8'b01011110; // 2736 :  94 - 0x5e -- Sprite 0xab
      13'hAB1: dout  = 8'b00001100; // 2737 :  12 - 0xc
      13'hAB2: dout  = 8'b10011110; // 2738 : 158 - 0x9e
      13'hAB3: dout  = 8'b11111110; // 2739 : 254 - 0xfe
      13'hAB4: dout  = 8'b11111110; // 2740 : 254 - 0xfe
      13'hAB5: dout  = 8'b11111110; // 2741 : 254 - 0xfe
      13'hAB6: dout  = 8'b11111000; // 2742 : 248 - 0xf8
      13'hAB7: dout  = 8'b11000000; // 2743 : 192 - 0xc0
      13'hAB8: dout  = 8'b10101100; // 2744 : 172 - 0xac
      13'hAB9: dout  = 8'b11111000; // 2745 : 248 - 0xf8
      13'hABA: dout  = 8'b11111000; // 2746 : 248 - 0xf8
      13'hABB: dout  = 8'b11111000; // 2747 : 248 - 0xf8
      13'hABC: dout  = 8'b11110000; // 2748 : 240 - 0xf0
      13'hABD: dout  = 8'b11000000; // 2749 : 192 - 0xc0
      13'hABE: dout  = 8'b00000000; // 2750 :   0 - 0x0
      13'hABF: dout  = 8'b00000000; // 2751 :   0 - 0x0
      13'hAC0: dout  = 8'b00000000; // 2752 :   0 - 0x0 -- Sprite 0xac
      13'hAC1: dout  = 8'b00000000; // 2753 :   0 - 0x0
      13'hAC2: dout  = 8'b00000000; // 2754 :   0 - 0x0
      13'hAC3: dout  = 8'b00000000; // 2755 :   0 - 0x0
      13'hAC4: dout  = 8'b00000000; // 2756 :   0 - 0x0
      13'hAC5: dout  = 8'b00000011; // 2757 :   3 - 0x3
      13'hAC6: dout  = 8'b00000111; // 2758 :   7 - 0x7
      13'hAC7: dout  = 8'b00101111; // 2759 :  47 - 0x2f
      13'hAC8: dout  = 8'b00000000; // 2760 :   0 - 0x0
      13'hAC9: dout  = 8'b00000000; // 2761 :   0 - 0x0
      13'hACA: dout  = 8'b00000000; // 2762 :   0 - 0x0
      13'hACB: dout  = 8'b00000000; // 2763 :   0 - 0x0
      13'hACC: dout  = 8'b00000000; // 2764 :   0 - 0x0
      13'hACD: dout  = 8'b00000000; // 2765 :   0 - 0x0
      13'hACE: dout  = 8'b00000001; // 2766 :   1 - 0x1
      13'hACF: dout  = 8'b00000011; // 2767 :   3 - 0x3
      13'hAD0: dout  = 8'b01001110; // 2768 :  78 - 0x4e -- Sprite 0xad
      13'hAD1: dout  = 8'b01101110; // 2769 : 110 - 0x6e
      13'hAD2: dout  = 8'b11111110; // 2770 : 254 - 0xfe
      13'hAD3: dout  = 8'b01111111; // 2771 : 127 - 0x7f
      13'hAD4: dout  = 8'b00111111; // 2772 :  63 - 0x3f
      13'hAD5: dout  = 8'b00011111; // 2773 :  31 - 0x1f
      13'hAD6: dout  = 8'b00001111; // 2774 :  15 - 0xf
      13'hAD7: dout  = 8'b00000011; // 2775 :   3 - 0x3
      13'hAD8: dout  = 8'b00000111; // 2776 :   7 - 0x7
      13'hAD9: dout  = 8'b00000111; // 2777 :   7 - 0x7
      13'hADA: dout  = 8'b00000111; // 2778 :   7 - 0x7
      13'hADB: dout  = 8'b00100111; // 2779 :  39 - 0x27
      13'hADC: dout  = 8'b00011111; // 2780 :  31 - 0x1f
      13'hADD: dout  = 8'b00000111; // 2781 :   7 - 0x7
      13'hADE: dout  = 8'b00000001; // 2782 :   1 - 0x1
      13'hADF: dout  = 8'b00000000; // 2783 :   0 - 0x0
      13'hAE0: dout  = 8'b00000000; // 2784 :   0 - 0x0 -- Sprite 0xae
      13'hAE1: dout  = 8'b00000000; // 2785 :   0 - 0x0
      13'hAE2: dout  = 8'b00000000; // 2786 :   0 - 0x0
      13'hAE3: dout  = 8'b00000000; // 2787 :   0 - 0x0
      13'hAE4: dout  = 8'b11111000; // 2788 : 248 - 0xf8
      13'hAE5: dout  = 8'b11111100; // 2789 : 252 - 0xfc
      13'hAE6: dout  = 8'b11111110; // 2790 : 254 - 0xfe
      13'hAE7: dout  = 8'b01010110; // 2791 :  86 - 0x56
      13'hAE8: dout  = 8'b00000000; // 2792 :   0 - 0x0
      13'hAE9: dout  = 8'b00000000; // 2793 :   0 - 0x0
      13'hAEA: dout  = 8'b00000000; // 2794 :   0 - 0x0
      13'hAEB: dout  = 8'b00000000; // 2795 :   0 - 0x0
      13'hAEC: dout  = 8'b00000000; // 2796 :   0 - 0x0
      13'hAED: dout  = 8'b11110000; // 2797 : 240 - 0xf0
      13'hAEE: dout  = 8'b11111000; // 2798 : 248 - 0xf8
      13'hAEF: dout  = 8'b10101100; // 2799 : 172 - 0xac
      13'hAF0: dout  = 8'b01010110; // 2800 :  86 - 0x56 -- Sprite 0xaf
      13'hAF1: dout  = 8'b00001100; // 2801 :  12 - 0xc
      13'hAF2: dout  = 8'b00001110; // 2802 :  14 - 0xe
      13'hAF3: dout  = 8'b00011111; // 2803 :  31 - 0x1f
      13'hAF4: dout  = 8'b11111111; // 2804 : 255 - 0xff
      13'hAF5: dout  = 8'b11111111; // 2805 : 255 - 0xff
      13'hAF6: dout  = 8'b11111110; // 2806 : 254 - 0xfe
      13'hAF7: dout  = 8'b11111000; // 2807 : 248 - 0xf8
      13'hAF8: dout  = 8'b10101100; // 2808 : 172 - 0xac
      13'hAF9: dout  = 8'b11111000; // 2809 : 248 - 0xf8
      13'hAFA: dout  = 8'b11111000; // 2810 : 248 - 0xf8
      13'hAFB: dout  = 8'b11111100; // 2811 : 252 - 0xfc
      13'hAFC: dout  = 8'b11111100; // 2812 : 252 - 0xfc
      13'hAFD: dout  = 8'b11111000; // 2813 : 248 - 0xf8
      13'hAFE: dout  = 8'b11110000; // 2814 : 240 - 0xf0
      13'hAFF: dout  = 8'b00000000; // 2815 :   0 - 0x0
      13'hB00: dout  = 8'b11111111; // 2816 : 255 - 0xff -- Sprite 0xb0
      13'hB01: dout  = 8'b11111111; // 2817 : 255 - 0xff
      13'hB02: dout  = 8'b11111111; // 2818 : 255 - 0xff
      13'hB03: dout  = 8'b11111111; // 2819 : 255 - 0xff
      13'hB04: dout  = 8'b11111111; // 2820 : 255 - 0xff
      13'hB05: dout  = 8'b11111111; // 2821 : 255 - 0xff
      13'hB06: dout  = 8'b11111111; // 2822 : 255 - 0xff
      13'hB07: dout  = 8'b11111111; // 2823 : 255 - 0xff
      13'hB08: dout  = 8'b11111111; // 2824 : 255 - 0xff
      13'hB09: dout  = 8'b11111111; // 2825 : 255 - 0xff
      13'hB0A: dout  = 8'b11111111; // 2826 : 255 - 0xff
      13'hB0B: dout  = 8'b11111111; // 2827 : 255 - 0xff
      13'hB0C: dout  = 8'b11111111; // 2828 : 255 - 0xff
      13'hB0D: dout  = 8'b11111111; // 2829 : 255 - 0xff
      13'hB0E: dout  = 8'b11111111; // 2830 : 255 - 0xff
      13'hB0F: dout  = 8'b11111111; // 2831 : 255 - 0xff
      13'hB10: dout  = 8'b11111111; // 2832 : 255 - 0xff -- Sprite 0xb1
      13'hB11: dout  = 8'b11111111; // 2833 : 255 - 0xff
      13'hB12: dout  = 8'b11111111; // 2834 : 255 - 0xff
      13'hB13: dout  = 8'b11111111; // 2835 : 255 - 0xff
      13'hB14: dout  = 8'b11111111; // 2836 : 255 - 0xff
      13'hB15: dout  = 8'b11111111; // 2837 : 255 - 0xff
      13'hB16: dout  = 8'b11111111; // 2838 : 255 - 0xff
      13'hB17: dout  = 8'b11111111; // 2839 : 255 - 0xff
      13'hB18: dout  = 8'b11111111; // 2840 : 255 - 0xff
      13'hB19: dout  = 8'b11111111; // 2841 : 255 - 0xff
      13'hB1A: dout  = 8'b11111111; // 2842 : 255 - 0xff
      13'hB1B: dout  = 8'b11111111; // 2843 : 255 - 0xff
      13'hB1C: dout  = 8'b11111111; // 2844 : 255 - 0xff
      13'hB1D: dout  = 8'b11111111; // 2845 : 255 - 0xff
      13'hB1E: dout  = 8'b11111111; // 2846 : 255 - 0xff
      13'hB1F: dout  = 8'b11111111; // 2847 : 255 - 0xff
      13'hB20: dout  = 8'b11111111; // 2848 : 255 - 0xff -- Sprite 0xb2
      13'hB21: dout  = 8'b11111111; // 2849 : 255 - 0xff
      13'hB22: dout  = 8'b11111111; // 2850 : 255 - 0xff
      13'hB23: dout  = 8'b11111111; // 2851 : 255 - 0xff
      13'hB24: dout  = 8'b11111111; // 2852 : 255 - 0xff
      13'hB25: dout  = 8'b11111111; // 2853 : 255 - 0xff
      13'hB26: dout  = 8'b11111111; // 2854 : 255 - 0xff
      13'hB27: dout  = 8'b11111111; // 2855 : 255 - 0xff
      13'hB28: dout  = 8'b11111111; // 2856 : 255 - 0xff
      13'hB29: dout  = 8'b11111111; // 2857 : 255 - 0xff
      13'hB2A: dout  = 8'b11111111; // 2858 : 255 - 0xff
      13'hB2B: dout  = 8'b11111111; // 2859 : 255 - 0xff
      13'hB2C: dout  = 8'b11111111; // 2860 : 255 - 0xff
      13'hB2D: dout  = 8'b11111111; // 2861 : 255 - 0xff
      13'hB2E: dout  = 8'b11111111; // 2862 : 255 - 0xff
      13'hB2F: dout  = 8'b11111111; // 2863 : 255 - 0xff
      13'hB30: dout  = 8'b11111111; // 2864 : 255 - 0xff -- Sprite 0xb3
      13'hB31: dout  = 8'b11111111; // 2865 : 255 - 0xff
      13'hB32: dout  = 8'b11111111; // 2866 : 255 - 0xff
      13'hB33: dout  = 8'b11111111; // 2867 : 255 - 0xff
      13'hB34: dout  = 8'b11111111; // 2868 : 255 - 0xff
      13'hB35: dout  = 8'b11111111; // 2869 : 255 - 0xff
      13'hB36: dout  = 8'b11111111; // 2870 : 255 - 0xff
      13'hB37: dout  = 8'b11111111; // 2871 : 255 - 0xff
      13'hB38: dout  = 8'b11111111; // 2872 : 255 - 0xff
      13'hB39: dout  = 8'b11111111; // 2873 : 255 - 0xff
      13'hB3A: dout  = 8'b11111111; // 2874 : 255 - 0xff
      13'hB3B: dout  = 8'b11111111; // 2875 : 255 - 0xff
      13'hB3C: dout  = 8'b11111111; // 2876 : 255 - 0xff
      13'hB3D: dout  = 8'b11111111; // 2877 : 255 - 0xff
      13'hB3E: dout  = 8'b11111111; // 2878 : 255 - 0xff
      13'hB3F: dout  = 8'b11111111; // 2879 : 255 - 0xff
      13'hB40: dout  = 8'b11111111; // 2880 : 255 - 0xff -- Sprite 0xb4
      13'hB41: dout  = 8'b11111111; // 2881 : 255 - 0xff
      13'hB42: dout  = 8'b11111111; // 2882 : 255 - 0xff
      13'hB43: dout  = 8'b11111111; // 2883 : 255 - 0xff
      13'hB44: dout  = 8'b11111111; // 2884 : 255 - 0xff
      13'hB45: dout  = 8'b11111111; // 2885 : 255 - 0xff
      13'hB46: dout  = 8'b11111111; // 2886 : 255 - 0xff
      13'hB47: dout  = 8'b11111111; // 2887 : 255 - 0xff
      13'hB48: dout  = 8'b11111111; // 2888 : 255 - 0xff
      13'hB49: dout  = 8'b11111111; // 2889 : 255 - 0xff
      13'hB4A: dout  = 8'b11111111; // 2890 : 255 - 0xff
      13'hB4B: dout  = 8'b11111111; // 2891 : 255 - 0xff
      13'hB4C: dout  = 8'b11111111; // 2892 : 255 - 0xff
      13'hB4D: dout  = 8'b11111111; // 2893 : 255 - 0xff
      13'hB4E: dout  = 8'b11111111; // 2894 : 255 - 0xff
      13'hB4F: dout  = 8'b11111111; // 2895 : 255 - 0xff
      13'hB50: dout  = 8'b11111111; // 2896 : 255 - 0xff -- Sprite 0xb5
      13'hB51: dout  = 8'b11111111; // 2897 : 255 - 0xff
      13'hB52: dout  = 8'b11111111; // 2898 : 255 - 0xff
      13'hB53: dout  = 8'b11111111; // 2899 : 255 - 0xff
      13'hB54: dout  = 8'b11111111; // 2900 : 255 - 0xff
      13'hB55: dout  = 8'b11111111; // 2901 : 255 - 0xff
      13'hB56: dout  = 8'b11111111; // 2902 : 255 - 0xff
      13'hB57: dout  = 8'b11111111; // 2903 : 255 - 0xff
      13'hB58: dout  = 8'b11111111; // 2904 : 255 - 0xff
      13'hB59: dout  = 8'b11111111; // 2905 : 255 - 0xff
      13'hB5A: dout  = 8'b11111111; // 2906 : 255 - 0xff
      13'hB5B: dout  = 8'b11111111; // 2907 : 255 - 0xff
      13'hB5C: dout  = 8'b11111111; // 2908 : 255 - 0xff
      13'hB5D: dout  = 8'b11111111; // 2909 : 255 - 0xff
      13'hB5E: dout  = 8'b11111111; // 2910 : 255 - 0xff
      13'hB5F: dout  = 8'b11111111; // 2911 : 255 - 0xff
      13'hB60: dout  = 8'b11111111; // 2912 : 255 - 0xff -- Sprite 0xb6
      13'hB61: dout  = 8'b11111111; // 2913 : 255 - 0xff
      13'hB62: dout  = 8'b11111111; // 2914 : 255 - 0xff
      13'hB63: dout  = 8'b11111111; // 2915 : 255 - 0xff
      13'hB64: dout  = 8'b11111111; // 2916 : 255 - 0xff
      13'hB65: dout  = 8'b11111111; // 2917 : 255 - 0xff
      13'hB66: dout  = 8'b11111111; // 2918 : 255 - 0xff
      13'hB67: dout  = 8'b11111111; // 2919 : 255 - 0xff
      13'hB68: dout  = 8'b11111111; // 2920 : 255 - 0xff
      13'hB69: dout  = 8'b11111111; // 2921 : 255 - 0xff
      13'hB6A: dout  = 8'b11111111; // 2922 : 255 - 0xff
      13'hB6B: dout  = 8'b11111111; // 2923 : 255 - 0xff
      13'hB6C: dout  = 8'b11111111; // 2924 : 255 - 0xff
      13'hB6D: dout  = 8'b11111111; // 2925 : 255 - 0xff
      13'hB6E: dout  = 8'b11111111; // 2926 : 255 - 0xff
      13'hB6F: dout  = 8'b11111111; // 2927 : 255 - 0xff
      13'hB70: dout  = 8'b11111111; // 2928 : 255 - 0xff -- Sprite 0xb7
      13'hB71: dout  = 8'b11111111; // 2929 : 255 - 0xff
      13'hB72: dout  = 8'b11111111; // 2930 : 255 - 0xff
      13'hB73: dout  = 8'b11111111; // 2931 : 255 - 0xff
      13'hB74: dout  = 8'b11111111; // 2932 : 255 - 0xff
      13'hB75: dout  = 8'b11111111; // 2933 : 255 - 0xff
      13'hB76: dout  = 8'b11111111; // 2934 : 255 - 0xff
      13'hB77: dout  = 8'b11111111; // 2935 : 255 - 0xff
      13'hB78: dout  = 8'b11111111; // 2936 : 255 - 0xff
      13'hB79: dout  = 8'b11111111; // 2937 : 255 - 0xff
      13'hB7A: dout  = 8'b11111111; // 2938 : 255 - 0xff
      13'hB7B: dout  = 8'b11111111; // 2939 : 255 - 0xff
      13'hB7C: dout  = 8'b11111111; // 2940 : 255 - 0xff
      13'hB7D: dout  = 8'b11111111; // 2941 : 255 - 0xff
      13'hB7E: dout  = 8'b11111111; // 2942 : 255 - 0xff
      13'hB7F: dout  = 8'b11111111; // 2943 : 255 - 0xff
      13'hB80: dout  = 8'b00000000; // 2944 :   0 - 0x0 -- Sprite 0xb8
      13'hB81: dout  = 8'b00000111; // 2945 :   7 - 0x7
      13'hB82: dout  = 8'b00001000; // 2946 :   8 - 0x8
      13'hB83: dout  = 8'b00010000; // 2947 :  16 - 0x10
      13'hB84: dout  = 8'b00010000; // 2948 :  16 - 0x10
      13'hB85: dout  = 8'b00100000; // 2949 :  32 - 0x20
      13'hB86: dout  = 8'b00100000; // 2950 :  32 - 0x20
      13'hB87: dout  = 8'b00100000; // 2951 :  32 - 0x20
      13'hB88: dout  = 8'b00000000; // 2952 :   0 - 0x0
      13'hB89: dout  = 8'b00000111; // 2953 :   7 - 0x7
      13'hB8A: dout  = 8'b00001000; // 2954 :   8 - 0x8
      13'hB8B: dout  = 8'b00010000; // 2955 :  16 - 0x10
      13'hB8C: dout  = 8'b00010000; // 2956 :  16 - 0x10
      13'hB8D: dout  = 8'b00100000; // 2957 :  32 - 0x20
      13'hB8E: dout  = 8'b00100000; // 2958 :  32 - 0x20
      13'hB8F: dout  = 8'b00100000; // 2959 :  32 - 0x20
      13'hB90: dout  = 8'b00011111; // 2960 :  31 - 0x1f -- Sprite 0xb9
      13'hB91: dout  = 8'b00101111; // 2961 :  47 - 0x2f
      13'hB92: dout  = 8'b00110111; // 2962 :  55 - 0x37
      13'hB93: dout  = 8'b00111010; // 2963 :  58 - 0x3a
      13'hB94: dout  = 8'b00111101; // 2964 :  61 - 0x3d
      13'hB95: dout  = 8'b00111110; // 2965 :  62 - 0x3e
      13'hB96: dout  = 8'b00111111; // 2966 :  63 - 0x3f
      13'hB97: dout  = 8'b00000000; // 2967 :   0 - 0x0
      13'hB98: dout  = 8'b00011111; // 2968 :  31 - 0x1f
      13'hB99: dout  = 8'b00111111; // 2969 :  63 - 0x3f
      13'hB9A: dout  = 8'b00111111; // 2970 :  63 - 0x3f
      13'hB9B: dout  = 8'b00111111; // 2971 :  63 - 0x3f
      13'hB9C: dout  = 8'b00111110; // 2972 :  62 - 0x3e
      13'hB9D: dout  = 8'b00111111; // 2973 :  63 - 0x3f
      13'hB9E: dout  = 8'b00111111; // 2974 :  63 - 0x3f
      13'hB9F: dout  = 8'b00000000; // 2975 :   0 - 0x0
      13'hBA0: dout  = 8'b00000000; // 2976 :   0 - 0x0 -- Sprite 0xba
      13'hBA1: dout  = 8'b00000101; // 2977 :   5 - 0x5
      13'hBA2: dout  = 8'b00011001; // 2978 :  25 - 0x19
      13'hBA3: dout  = 8'b00110011; // 2979 :  51 - 0x33
      13'hBA4: dout  = 8'b01100011; // 2980 :  99 - 0x63
      13'hBA5: dout  = 8'b11000111; // 2981 : 199 - 0xc7
      13'hBA6: dout  = 8'b11000111; // 2982 : 199 - 0xc7
      13'hBA7: dout  = 8'b11000100; // 2983 : 196 - 0xc4
      13'hBA8: dout  = 8'b00000000; // 2984 :   0 - 0x0
      13'hBA9: dout  = 8'b00000111; // 2985 :   7 - 0x7
      13'hBAA: dout  = 8'b00011111; // 2986 :  31 - 0x1f
      13'hBAB: dout  = 8'b00111111; // 2987 :  63 - 0x3f
      13'hBAC: dout  = 8'b01111111; // 2988 : 127 - 0x7f
      13'hBAD: dout  = 8'b11111111; // 2989 : 255 - 0xff
      13'hBAE: dout  = 8'b11111111; // 2990 : 255 - 0xff
      13'hBAF: dout  = 8'b11011101; // 2991 : 221 - 0xdd
      13'hBB0: dout  = 8'b10000000; // 2992 : 128 - 0x80 -- Sprite 0xbb
      13'hBB1: dout  = 8'b00000000; // 2993 :   0 - 0x0
      13'hBB2: dout  = 8'b00000000; // 2994 :   0 - 0x0
      13'hBB3: dout  = 8'b00000000; // 2995 :   0 - 0x0
      13'hBB4: dout  = 8'b00000000; // 2996 :   0 - 0x0
      13'hBB5: dout  = 8'b00000011; // 2997 :   3 - 0x3
      13'hBB6: dout  = 8'b00000011; // 2998 :   3 - 0x3
      13'hBB7: dout  = 8'b00000000; // 2999 :   0 - 0x0
      13'hBB8: dout  = 8'b10001001; // 3000 : 137 - 0x89
      13'hBB9: dout  = 8'b00000001; // 3001 :   1 - 0x1
      13'hBBA: dout  = 8'b00000001; // 3002 :   1 - 0x1
      13'hBBB: dout  = 8'b00000001; // 3003 :   1 - 0x1
      13'hBBC: dout  = 8'b00000001; // 3004 :   1 - 0x1
      13'hBBD: dout  = 8'b00000000; // 3005 :   0 - 0x0
      13'hBBE: dout  = 8'b00000000; // 3006 :   0 - 0x0
      13'hBBF: dout  = 8'b00000000; // 3007 :   0 - 0x0
      13'hBC0: dout  = 8'b00000000; // 3008 :   0 - 0x0 -- Sprite 0xbc
      13'hBC1: dout  = 8'b00000000; // 3009 :   0 - 0x0
      13'hBC2: dout  = 8'b00000000; // 3010 :   0 - 0x0
      13'hBC3: dout  = 8'b00000000; // 3011 :   0 - 0x0
      13'hBC4: dout  = 8'b00000000; // 3012 :   0 - 0x0
      13'hBC5: dout  = 8'b00000000; // 3013 :   0 - 0x0
      13'hBC6: dout  = 8'b00000000; // 3014 :   0 - 0x0
      13'hBC7: dout  = 8'b00000000; // 3015 :   0 - 0x0
      13'hBC8: dout  = 8'b00000000; // 3016 :   0 - 0x0
      13'hBC9: dout  = 8'b00000000; // 3017 :   0 - 0x0
      13'hBCA: dout  = 8'b00000000; // 3018 :   0 - 0x0
      13'hBCB: dout  = 8'b00000000; // 3019 :   0 - 0x0
      13'hBCC: dout  = 8'b00000000; // 3020 :   0 - 0x0
      13'hBCD: dout  = 8'b00000000; // 3021 :   0 - 0x0
      13'hBCE: dout  = 8'b00000011; // 3022 :   3 - 0x3
      13'hBCF: dout  = 8'b00000111; // 3023 :   7 - 0x7
      13'hBD0: dout  = 8'b00000000; // 3024 :   0 - 0x0 -- Sprite 0xbd
      13'hBD1: dout  = 8'b00000000; // 3025 :   0 - 0x0
      13'hBD2: dout  = 8'b00001111; // 3026 :  15 - 0xf
      13'hBD3: dout  = 8'b00000000; // 3027 :   0 - 0x0
      13'hBD4: dout  = 8'b10000000; // 3028 : 128 - 0x80
      13'hBD5: dout  = 8'b01100011; // 3029 :  99 - 0x63
      13'hBD6: dout  = 8'b00011110; // 3030 :  30 - 0x1e
      13'hBD7: dout  = 8'b00000000; // 3031 :   0 - 0x0
      13'hBD8: dout  = 8'b00001111; // 3032 :  15 - 0xf
      13'hBD9: dout  = 8'b00001111; // 3033 :  15 - 0xf
      13'hBDA: dout  = 8'b00000000; // 3034 :   0 - 0x0
      13'hBDB: dout  = 8'b00011111; // 3035 :  31 - 0x1f
      13'hBDC: dout  = 8'b01111111; // 3036 : 127 - 0x7f
      13'hBDD: dout  = 8'b00011100; // 3037 :  28 - 0x1c
      13'hBDE: dout  = 8'b00000000; // 3038 :   0 - 0x0
      13'hBDF: dout  = 8'b00000000; // 3039 :   0 - 0x0
      13'hBE0: dout  = 8'b00000001; // 3040 :   1 - 0x1 -- Sprite 0xbe
      13'hBE1: dout  = 8'b00000011; // 3041 :   3 - 0x3
      13'hBE2: dout  = 8'b00011001; // 3042 :  25 - 0x19
      13'hBE3: dout  = 8'b00111100; // 3043 :  60 - 0x3c
      13'hBE4: dout  = 8'b00011001; // 3044 :  25 - 0x19
      13'hBE5: dout  = 8'b00100011; // 3045 :  35 - 0x23
      13'hBE6: dout  = 8'b01010001; // 3046 :  81 - 0x51
      13'hBE7: dout  = 8'b00100000; // 3047 :  32 - 0x20
      13'hBE8: dout  = 8'b00000001; // 3048 :   1 - 0x1
      13'hBE9: dout  = 8'b00000010; // 3049 :   2 - 0x2
      13'hBEA: dout  = 8'b00011001; // 3050 :  25 - 0x19
      13'hBEB: dout  = 8'b00100100; // 3051 :  36 - 0x24
      13'hBEC: dout  = 8'b00011001; // 3052 :  25 - 0x19
      13'hBED: dout  = 8'b00100010; // 3053 :  34 - 0x22
      13'hBEE: dout  = 8'b00010001; // 3054 :  17 - 0x11
      13'hBEF: dout  = 8'b00101100; // 3055 :  44 - 0x2c
      13'hBF0: dout  = 8'b00000000; // 3056 :   0 - 0x0 -- Sprite 0xbf
      13'hBF1: dout  = 8'b00000000; // 3057 :   0 - 0x0
      13'hBF2: dout  = 8'b00000000; // 3058 :   0 - 0x0
      13'hBF3: dout  = 8'b00000000; // 3059 :   0 - 0x0
      13'hBF4: dout  = 8'b00000000; // 3060 :   0 - 0x0
      13'hBF5: dout  = 8'b00000000; // 3061 :   0 - 0x0
      13'hBF6: dout  = 8'b00000000; // 3062 :   0 - 0x0
      13'hBF7: dout  = 8'b00000000; // 3063 :   0 - 0x0
      13'hBF8: dout  = 8'b00011111; // 3064 :  31 - 0x1f
      13'hBF9: dout  = 8'b00000111; // 3065 :   7 - 0x7
      13'hBFA: dout  = 8'b00000011; // 3066 :   3 - 0x3
      13'hBFB: dout  = 8'b00000011; // 3067 :   3 - 0x3
      13'hBFC: dout  = 8'b00000001; // 3068 :   1 - 0x1
      13'hBFD: dout  = 8'b00000001; // 3069 :   1 - 0x1
      13'hBFE: dout  = 8'b00000001; // 3070 :   1 - 0x1
      13'hBFF: dout  = 8'b00000000; // 3071 :   0 - 0x0
      13'hC00: dout  = 8'b00000000; // 3072 :   0 - 0x0 -- Sprite 0xc0
      13'hC01: dout  = 8'b00111111; // 3073 :  63 - 0x3f
      13'hC02: dout  = 8'b00011111; // 3074 :  31 - 0x1f
      13'hC03: dout  = 8'b00000000; // 3075 :   0 - 0x0
      13'hC04: dout  = 8'b00000001; // 3076 :   1 - 0x1
      13'hC05: dout  = 8'b00000000; // 3077 :   0 - 0x0
      13'hC06: dout  = 8'b00000001; // 3078 :   1 - 0x1
      13'hC07: dout  = 8'b00000000; // 3079 :   0 - 0x0
      13'hC08: dout  = 8'b00000000; // 3080 :   0 - 0x0
      13'hC09: dout  = 8'b00000000; // 3081 :   0 - 0x0
      13'hC0A: dout  = 8'b00000000; // 3082 :   0 - 0x0
      13'hC0B: dout  = 8'b00000001; // 3083 :   1 - 0x1
      13'hC0C: dout  = 8'b00000011; // 3084 :   3 - 0x3
      13'hC0D: dout  = 8'b00000111; // 3085 :   7 - 0x7
      13'hC0E: dout  = 8'b00001101; // 3086 :  13 - 0xd
      13'hC0F: dout  = 8'b00011001; // 3087 :  25 - 0x19
      13'hC10: dout  = 8'b00010001; // 3088 :  17 - 0x11 -- Sprite 0xc1
      13'hC11: dout  = 8'b00000000; // 3089 :   0 - 0x0
      13'hC12: dout  = 8'b00000001; // 3090 :   1 - 0x1
      13'hC13: dout  = 8'b00000000; // 3091 :   0 - 0x0
      13'hC14: dout  = 8'b00000001; // 3092 :   1 - 0x1
      13'hC15: dout  = 8'b00000000; // 3093 :   0 - 0x0
      13'hC16: dout  = 8'b00011111; // 3094 :  31 - 0x1f
      13'hC17: dout  = 8'b00111111; // 3095 :  63 - 0x3f
      13'hC18: dout  = 8'b00101001; // 3096 :  41 - 0x29
      13'hC19: dout  = 8'b00011001; // 3097 :  25 - 0x19
      13'hC1A: dout  = 8'b00001101; // 3098 :  13 - 0xd
      13'hC1B: dout  = 8'b00000111; // 3099 :   7 - 0x7
      13'hC1C: dout  = 8'b00000011; // 3100 :   3 - 0x3
      13'hC1D: dout  = 8'b00000001; // 3101 :   1 - 0x1
      13'hC1E: dout  = 8'b00000000; // 3102 :   0 - 0x0
      13'hC1F: dout  = 8'b00000000; // 3103 :   0 - 0x0
      13'hC20: dout  = 8'b00000000; // 3104 :   0 - 0x0 -- Sprite 0xc2
      13'hC21: dout  = 8'b11111100; // 3105 : 252 - 0xfc
      13'hC22: dout  = 8'b11111000; // 3106 : 248 - 0xf8
      13'hC23: dout  = 8'b00000000; // 3107 :   0 - 0x0
      13'hC24: dout  = 8'b10000000; // 3108 : 128 - 0x80
      13'hC25: dout  = 8'b00000000; // 3109 :   0 - 0x0
      13'hC26: dout  = 8'b10000000; // 3110 : 128 - 0x80
      13'hC27: dout  = 8'b00000000; // 3111 :   0 - 0x0
      13'hC28: dout  = 8'b00000000; // 3112 :   0 - 0x0
      13'hC29: dout  = 8'b00000000; // 3113 :   0 - 0x0
      13'hC2A: dout  = 8'b00000000; // 3114 :   0 - 0x0
      13'hC2B: dout  = 8'b10000000; // 3115 : 128 - 0x80
      13'hC2C: dout  = 8'b11000000; // 3116 : 192 - 0xc0
      13'hC2D: dout  = 8'b11100000; // 3117 : 224 - 0xe0
      13'hC2E: dout  = 8'b10110000; // 3118 : 176 - 0xb0
      13'hC2F: dout  = 8'b10011000; // 3119 : 152 - 0x98
      13'hC30: dout  = 8'b10001000; // 3120 : 136 - 0x88 -- Sprite 0xc3
      13'hC31: dout  = 8'b00000000; // 3121 :   0 - 0x0
      13'hC32: dout  = 8'b10000000; // 3122 : 128 - 0x80
      13'hC33: dout  = 8'b00000000; // 3123 :   0 - 0x0
      13'hC34: dout  = 8'b10000000; // 3124 : 128 - 0x80
      13'hC35: dout  = 8'b00000000; // 3125 :   0 - 0x0
      13'hC36: dout  = 8'b11111000; // 3126 : 248 - 0xf8
      13'hC37: dout  = 8'b11111100; // 3127 : 252 - 0xfc
      13'hC38: dout  = 8'b10010100; // 3128 : 148 - 0x94
      13'hC39: dout  = 8'b10011000; // 3129 : 152 - 0x98
      13'hC3A: dout  = 8'b10110000; // 3130 : 176 - 0xb0
      13'hC3B: dout  = 8'b11100000; // 3131 : 224 - 0xe0
      13'hC3C: dout  = 8'b11000000; // 3132 : 192 - 0xc0
      13'hC3D: dout  = 8'b10000000; // 3133 : 128 - 0x80
      13'hC3E: dout  = 8'b00000000; // 3134 :   0 - 0x0
      13'hC3F: dout  = 8'b00000000; // 3135 :   0 - 0x0
      13'hC40: dout  = 8'b00000000; // 3136 :   0 - 0x0 -- Sprite 0xc4
      13'hC41: dout  = 8'b00000000; // 3137 :   0 - 0x0
      13'hC42: dout  = 8'b00000000; // 3138 :   0 - 0x0
      13'hC43: dout  = 8'b00000000; // 3139 :   0 - 0x0
      13'hC44: dout  = 8'b00000000; // 3140 :   0 - 0x0
      13'hC45: dout  = 8'b00111111; // 3141 :  63 - 0x3f
      13'hC46: dout  = 8'b00011111; // 3142 :  31 - 0x1f
      13'hC47: dout  = 8'b00000000; // 3143 :   0 - 0x0
      13'hC48: dout  = 8'b00000000; // 3144 :   0 - 0x0
      13'hC49: dout  = 8'b00000000; // 3145 :   0 - 0x0
      13'hC4A: dout  = 8'b00000000; // 3146 :   0 - 0x0
      13'hC4B: dout  = 8'b00000000; // 3147 :   0 - 0x0
      13'hC4C: dout  = 8'b00000000; // 3148 :   0 - 0x0
      13'hC4D: dout  = 8'b00000000; // 3149 :   0 - 0x0
      13'hC4E: dout  = 8'b00000000; // 3150 :   0 - 0x0
      13'hC4F: dout  = 8'b00000001; // 3151 :   1 - 0x1
      13'hC50: dout  = 8'b00000001; // 3152 :   1 - 0x1 -- Sprite 0xc5
      13'hC51: dout  = 8'b00000001; // 3153 :   1 - 0x1
      13'hC52: dout  = 8'b01000001; // 3154 :  65 - 0x41
      13'hC53: dout  = 8'b00000001; // 3155 :   1 - 0x1
      13'hC54: dout  = 8'b00000001; // 3156 :   1 - 0x1
      13'hC55: dout  = 8'b00000000; // 3157 :   0 - 0x0
      13'hC56: dout  = 8'b00011111; // 3158 :  31 - 0x1f
      13'hC57: dout  = 8'b00111111; // 3159 :  63 - 0x3f
      13'hC58: dout  = 8'b00001111; // 3160 :  15 - 0xf
      13'hC59: dout  = 8'b01111001; // 3161 : 121 - 0x79
      13'hC5A: dout  = 8'b10100001; // 3162 : 161 - 0xa1
      13'hC5B: dout  = 8'b01111001; // 3163 : 121 - 0x79
      13'hC5C: dout  = 8'b00001111; // 3164 :  15 - 0xf
      13'hC5D: dout  = 8'b00000001; // 3165 :   1 - 0x1
      13'hC5E: dout  = 8'b00000000; // 3166 :   0 - 0x0
      13'hC5F: dout  = 8'b00000000; // 3167 :   0 - 0x0
      13'hC60: dout  = 8'b00000000; // 3168 :   0 - 0x0 -- Sprite 0xc6
      13'hC61: dout  = 8'b00000000; // 3169 :   0 - 0x0
      13'hC62: dout  = 8'b00000000; // 3170 :   0 - 0x0
      13'hC63: dout  = 8'b00000000; // 3171 :   0 - 0x0
      13'hC64: dout  = 8'b00000000; // 3172 :   0 - 0x0
      13'hC65: dout  = 8'b11111100; // 3173 : 252 - 0xfc
      13'hC66: dout  = 8'b11111000; // 3174 : 248 - 0xf8
      13'hC67: dout  = 8'b00000000; // 3175 :   0 - 0x0
      13'hC68: dout  = 8'b00000000; // 3176 :   0 - 0x0
      13'hC69: dout  = 8'b00000000; // 3177 :   0 - 0x0
      13'hC6A: dout  = 8'b00000000; // 3178 :   0 - 0x0
      13'hC6B: dout  = 8'b00000000; // 3179 :   0 - 0x0
      13'hC6C: dout  = 8'b00000000; // 3180 :   0 - 0x0
      13'hC6D: dout  = 8'b00000000; // 3181 :   0 - 0x0
      13'hC6E: dout  = 8'b00000000; // 3182 :   0 - 0x0
      13'hC6F: dout  = 8'b10000000; // 3183 : 128 - 0x80
      13'hC70: dout  = 8'b10000000; // 3184 : 128 - 0x80 -- Sprite 0xc7
      13'hC71: dout  = 8'b10000000; // 3185 : 128 - 0x80
      13'hC72: dout  = 8'b10000010; // 3186 : 130 - 0x82
      13'hC73: dout  = 8'b10000000; // 3187 : 128 - 0x80
      13'hC74: dout  = 8'b10000000; // 3188 : 128 - 0x80
      13'hC75: dout  = 8'b00000000; // 3189 :   0 - 0x0
      13'hC76: dout  = 8'b11111000; // 3190 : 248 - 0xf8
      13'hC77: dout  = 8'b11111100; // 3191 : 252 - 0xfc
      13'hC78: dout  = 8'b11110000; // 3192 : 240 - 0xf0
      13'hC79: dout  = 8'b10011110; // 3193 : 158 - 0x9e
      13'hC7A: dout  = 8'b10000101; // 3194 : 133 - 0x85
      13'hC7B: dout  = 8'b10011110; // 3195 : 158 - 0x9e
      13'hC7C: dout  = 8'b11110000; // 3196 : 240 - 0xf0
      13'hC7D: dout  = 8'b10000000; // 3197 : 128 - 0x80
      13'hC7E: dout  = 8'b00000000; // 3198 :   0 - 0x0
      13'hC7F: dout  = 8'b00000000; // 3199 :   0 - 0x0
      13'hC80: dout  = 8'b00000000; // 3200 :   0 - 0x0 -- Sprite 0xc8
      13'hC81: dout  = 8'b00000000; // 3201 :   0 - 0x0
      13'hC82: dout  = 8'b00000000; // 3202 :   0 - 0x0
      13'hC83: dout  = 8'b00011110; // 3203 :  30 - 0x1e
      13'hC84: dout  = 8'b00111111; // 3204 :  63 - 0x3f
      13'hC85: dout  = 8'b00111111; // 3205 :  63 - 0x3f
      13'hC86: dout  = 8'b00111111; // 3206 :  63 - 0x3f
      13'hC87: dout  = 8'b00111111; // 3207 :  63 - 0x3f
      13'hC88: dout  = 8'b00000000; // 3208 :   0 - 0x0
      13'hC89: dout  = 8'b00000000; // 3209 :   0 - 0x0
      13'hC8A: dout  = 8'b00000000; // 3210 :   0 - 0x0
      13'hC8B: dout  = 8'b00011110; // 3211 :  30 - 0x1e
      13'hC8C: dout  = 8'b00111111; // 3212 :  63 - 0x3f
      13'hC8D: dout  = 8'b00111111; // 3213 :  63 - 0x3f
      13'hC8E: dout  = 8'b00111111; // 3214 :  63 - 0x3f
      13'hC8F: dout  = 8'b00111111; // 3215 :  63 - 0x3f
      13'hC90: dout  = 8'b00011111; // 3216 :  31 - 0x1f -- Sprite 0xc9
      13'hC91: dout  = 8'b00001111; // 3217 :  15 - 0xf
      13'hC92: dout  = 8'b00000111; // 3218 :   7 - 0x7
      13'hC93: dout  = 8'b00000011; // 3219 :   3 - 0x3
      13'hC94: dout  = 8'b00000001; // 3220 :   1 - 0x1
      13'hC95: dout  = 8'b00000000; // 3221 :   0 - 0x0
      13'hC96: dout  = 8'b00000000; // 3222 :   0 - 0x0
      13'hC97: dout  = 8'b00000000; // 3223 :   0 - 0x0
      13'hC98: dout  = 8'b00011111; // 3224 :  31 - 0x1f
      13'hC99: dout  = 8'b00001111; // 3225 :  15 - 0xf
      13'hC9A: dout  = 8'b00000111; // 3226 :   7 - 0x7
      13'hC9B: dout  = 8'b00000011; // 3227 :   3 - 0x3
      13'hC9C: dout  = 8'b00000001; // 3228 :   1 - 0x1
      13'hC9D: dout  = 8'b00000000; // 3229 :   0 - 0x0
      13'hC9E: dout  = 8'b00000000; // 3230 :   0 - 0x0
      13'hC9F: dout  = 8'b00000000; // 3231 :   0 - 0x0
      13'hCA0: dout  = 8'b00000000; // 3232 :   0 - 0x0 -- Sprite 0xca
      13'hCA1: dout  = 8'b00000000; // 3233 :   0 - 0x0
      13'hCA2: dout  = 8'b00000000; // 3234 :   0 - 0x0
      13'hCA3: dout  = 8'b00111100; // 3235 :  60 - 0x3c
      13'hCA4: dout  = 8'b01111110; // 3236 : 126 - 0x7e
      13'hCA5: dout  = 8'b11111110; // 3237 : 254 - 0xfe
      13'hCA6: dout  = 8'b11111110; // 3238 : 254 - 0xfe
      13'hCA7: dout  = 8'b11111110; // 3239 : 254 - 0xfe
      13'hCA8: dout  = 8'b00000000; // 3240 :   0 - 0x0
      13'hCA9: dout  = 8'b00000000; // 3241 :   0 - 0x0
      13'hCAA: dout  = 8'b00000000; // 3242 :   0 - 0x0
      13'hCAB: dout  = 8'b00111100; // 3243 :  60 - 0x3c
      13'hCAC: dout  = 8'b01111110; // 3244 : 126 - 0x7e
      13'hCAD: dout  = 8'b11111110; // 3245 : 254 - 0xfe
      13'hCAE: dout  = 8'b11111110; // 3246 : 254 - 0xfe
      13'hCAF: dout  = 8'b11111110; // 3247 : 254 - 0xfe
      13'hCB0: dout  = 8'b11111100; // 3248 : 252 - 0xfc -- Sprite 0xcb
      13'hCB1: dout  = 8'b11111000; // 3249 : 248 - 0xf8
      13'hCB2: dout  = 8'b11110000; // 3250 : 240 - 0xf0
      13'hCB3: dout  = 8'b11100000; // 3251 : 224 - 0xe0
      13'hCB4: dout  = 8'b11000000; // 3252 : 192 - 0xc0
      13'hCB5: dout  = 8'b10000000; // 3253 : 128 - 0x80
      13'hCB6: dout  = 8'b00000000; // 3254 :   0 - 0x0
      13'hCB7: dout  = 8'b00000000; // 3255 :   0 - 0x0
      13'hCB8: dout  = 8'b11111100; // 3256 : 252 - 0xfc
      13'hCB9: dout  = 8'b11111000; // 3257 : 248 - 0xf8
      13'hCBA: dout  = 8'b11110000; // 3258 : 240 - 0xf0
      13'hCBB: dout  = 8'b11100000; // 3259 : 224 - 0xe0
      13'hCBC: dout  = 8'b11000000; // 3260 : 192 - 0xc0
      13'hCBD: dout  = 8'b10000000; // 3261 : 128 - 0x80
      13'hCBE: dout  = 8'b00000000; // 3262 :   0 - 0x0
      13'hCBF: dout  = 8'b00000000; // 3263 :   0 - 0x0
      13'hCC0: dout  = 8'b11111111; // 3264 : 255 - 0xff -- Sprite 0xcc
      13'hCC1: dout  = 8'b11111111; // 3265 : 255 - 0xff
      13'hCC2: dout  = 8'b11111111; // 3266 : 255 - 0xff
      13'hCC3: dout  = 8'b11111111; // 3267 : 255 - 0xff
      13'hCC4: dout  = 8'b11111111; // 3268 : 255 - 0xff
      13'hCC5: dout  = 8'b11111111; // 3269 : 255 - 0xff
      13'hCC6: dout  = 8'b11111111; // 3270 : 255 - 0xff
      13'hCC7: dout  = 8'b11111111; // 3271 : 255 - 0xff
      13'hCC8: dout  = 8'b11111111; // 3272 : 255 - 0xff
      13'hCC9: dout  = 8'b11111111; // 3273 : 255 - 0xff
      13'hCCA: dout  = 8'b11111111; // 3274 : 255 - 0xff
      13'hCCB: dout  = 8'b11111111; // 3275 : 255 - 0xff
      13'hCCC: dout  = 8'b11111111; // 3276 : 255 - 0xff
      13'hCCD: dout  = 8'b11111111; // 3277 : 255 - 0xff
      13'hCCE: dout  = 8'b11111111; // 3278 : 255 - 0xff
      13'hCCF: dout  = 8'b11111111; // 3279 : 255 - 0xff
      13'hCD0: dout  = 8'b11111111; // 3280 : 255 - 0xff -- Sprite 0xcd
      13'hCD1: dout  = 8'b11111111; // 3281 : 255 - 0xff
      13'hCD2: dout  = 8'b11111111; // 3282 : 255 - 0xff
      13'hCD3: dout  = 8'b11111111; // 3283 : 255 - 0xff
      13'hCD4: dout  = 8'b11111111; // 3284 : 255 - 0xff
      13'hCD5: dout  = 8'b11111111; // 3285 : 255 - 0xff
      13'hCD6: dout  = 8'b11111111; // 3286 : 255 - 0xff
      13'hCD7: dout  = 8'b11111111; // 3287 : 255 - 0xff
      13'hCD8: dout  = 8'b11111111; // 3288 : 255 - 0xff
      13'hCD9: dout  = 8'b11111111; // 3289 : 255 - 0xff
      13'hCDA: dout  = 8'b11111111; // 3290 : 255 - 0xff
      13'hCDB: dout  = 8'b11111111; // 3291 : 255 - 0xff
      13'hCDC: dout  = 8'b11111111; // 3292 : 255 - 0xff
      13'hCDD: dout  = 8'b11111111; // 3293 : 255 - 0xff
      13'hCDE: dout  = 8'b11111111; // 3294 : 255 - 0xff
      13'hCDF: dout  = 8'b11111111; // 3295 : 255 - 0xff
      13'hCE0: dout  = 8'b11111111; // 3296 : 255 - 0xff -- Sprite 0xce
      13'hCE1: dout  = 8'b11111111; // 3297 : 255 - 0xff
      13'hCE2: dout  = 8'b11111111; // 3298 : 255 - 0xff
      13'hCE3: dout  = 8'b11111111; // 3299 : 255 - 0xff
      13'hCE4: dout  = 8'b11111111; // 3300 : 255 - 0xff
      13'hCE5: dout  = 8'b11111111; // 3301 : 255 - 0xff
      13'hCE6: dout  = 8'b11111111; // 3302 : 255 - 0xff
      13'hCE7: dout  = 8'b11111111; // 3303 : 255 - 0xff
      13'hCE8: dout  = 8'b11111111; // 3304 : 255 - 0xff
      13'hCE9: dout  = 8'b11111111; // 3305 : 255 - 0xff
      13'hCEA: dout  = 8'b11111111; // 3306 : 255 - 0xff
      13'hCEB: dout  = 8'b11111111; // 3307 : 255 - 0xff
      13'hCEC: dout  = 8'b11111111; // 3308 : 255 - 0xff
      13'hCED: dout  = 8'b11111111; // 3309 : 255 - 0xff
      13'hCEE: dout  = 8'b11111111; // 3310 : 255 - 0xff
      13'hCEF: dout  = 8'b11111111; // 3311 : 255 - 0xff
      13'hCF0: dout  = 8'b11111111; // 3312 : 255 - 0xff -- Sprite 0xcf
      13'hCF1: dout  = 8'b11111111; // 3313 : 255 - 0xff
      13'hCF2: dout  = 8'b11111111; // 3314 : 255 - 0xff
      13'hCF3: dout  = 8'b11111111; // 3315 : 255 - 0xff
      13'hCF4: dout  = 8'b11111111; // 3316 : 255 - 0xff
      13'hCF5: dout  = 8'b11111111; // 3317 : 255 - 0xff
      13'hCF6: dout  = 8'b11111111; // 3318 : 255 - 0xff
      13'hCF7: dout  = 8'b11111111; // 3319 : 255 - 0xff
      13'hCF8: dout  = 8'b11111111; // 3320 : 255 - 0xff
      13'hCF9: dout  = 8'b11111111; // 3321 : 255 - 0xff
      13'hCFA: dout  = 8'b11111111; // 3322 : 255 - 0xff
      13'hCFB: dout  = 8'b11111111; // 3323 : 255 - 0xff
      13'hCFC: dout  = 8'b11111111; // 3324 : 255 - 0xff
      13'hCFD: dout  = 8'b11111111; // 3325 : 255 - 0xff
      13'hCFE: dout  = 8'b11111111; // 3326 : 255 - 0xff
      13'hCFF: dout  = 8'b11111111; // 3327 : 255 - 0xff
      13'hD00: dout  = 8'b00001000; // 3328 :   8 - 0x8 -- Sprite 0xd0
      13'hD01: dout  = 8'b00011001; // 3329 :  25 - 0x19
      13'hD02: dout  = 8'b00001001; // 3330 :   9 - 0x9
      13'hD03: dout  = 8'b00001001; // 3331 :   9 - 0x9
      13'hD04: dout  = 8'b00001001; // 3332 :   9 - 0x9
      13'hD05: dout  = 8'b00001001; // 3333 :   9 - 0x9
      13'hD06: dout  = 8'b00011100; // 3334 :  28 - 0x1c
      13'hD07: dout  = 8'b00000000; // 3335 :   0 - 0x0
      13'hD08: dout  = 8'b00000000; // 3336 :   0 - 0x0
      13'hD09: dout  = 8'b00000000; // 3337 :   0 - 0x0
      13'hD0A: dout  = 8'b00000000; // 3338 :   0 - 0x0
      13'hD0B: dout  = 8'b00000000; // 3339 :   0 - 0x0
      13'hD0C: dout  = 8'b00000000; // 3340 :   0 - 0x0
      13'hD0D: dout  = 8'b00000000; // 3341 :   0 - 0x0
      13'hD0E: dout  = 8'b00000000; // 3342 :   0 - 0x0
      13'hD0F: dout  = 8'b00000000; // 3343 :   0 - 0x0
      13'hD10: dout  = 8'b00111000; // 3344 :  56 - 0x38 -- Sprite 0xd1
      13'hD11: dout  = 8'b00000101; // 3345 :   5 - 0x5
      13'hD12: dout  = 8'b00000101; // 3346 :   5 - 0x5
      13'hD13: dout  = 8'b00011001; // 3347 :  25 - 0x19
      13'hD14: dout  = 8'b00000101; // 3348 :   5 - 0x5
      13'hD15: dout  = 8'b00000101; // 3349 :   5 - 0x5
      13'hD16: dout  = 8'b00111000; // 3350 :  56 - 0x38
      13'hD17: dout  = 8'b00000000; // 3351 :   0 - 0x0
      13'hD18: dout  = 8'b00000000; // 3352 :   0 - 0x0
      13'hD19: dout  = 8'b00000000; // 3353 :   0 - 0x0
      13'hD1A: dout  = 8'b00000000; // 3354 :   0 - 0x0
      13'hD1B: dout  = 8'b00000000; // 3355 :   0 - 0x0
      13'hD1C: dout  = 8'b00000000; // 3356 :   0 - 0x0
      13'hD1D: dout  = 8'b00000000; // 3357 :   0 - 0x0
      13'hD1E: dout  = 8'b00000000; // 3358 :   0 - 0x0
      13'hD1F: dout  = 8'b00000000; // 3359 :   0 - 0x0
      13'hD20: dout  = 8'b00111100; // 3360 :  60 - 0x3c -- Sprite 0xd2
      13'hD21: dout  = 8'b00100001; // 3361 :  33 - 0x21
      13'hD22: dout  = 8'b00100001; // 3362 :  33 - 0x21
      13'hD23: dout  = 8'b00111101; // 3363 :  61 - 0x3d
      13'hD24: dout  = 8'b00000101; // 3364 :   5 - 0x5
      13'hD25: dout  = 8'b00000101; // 3365 :   5 - 0x5
      13'hD26: dout  = 8'b00111000; // 3366 :  56 - 0x38
      13'hD27: dout  = 8'b00000000; // 3367 :   0 - 0x0
      13'hD28: dout  = 8'b00000000; // 3368 :   0 - 0x0
      13'hD29: dout  = 8'b00000000; // 3369 :   0 - 0x0
      13'hD2A: dout  = 8'b00000000; // 3370 :   0 - 0x0
      13'hD2B: dout  = 8'b00000000; // 3371 :   0 - 0x0
      13'hD2C: dout  = 8'b00000000; // 3372 :   0 - 0x0
      13'hD2D: dout  = 8'b00000000; // 3373 :   0 - 0x0
      13'hD2E: dout  = 8'b00000000; // 3374 :   0 - 0x0
      13'hD2F: dout  = 8'b00000000; // 3375 :   0 - 0x0
      13'hD30: dout  = 8'b00011000; // 3376 :  24 - 0x18 -- Sprite 0xd3
      13'hD31: dout  = 8'b00100101; // 3377 :  37 - 0x25
      13'hD32: dout  = 8'b00100101; // 3378 :  37 - 0x25
      13'hD33: dout  = 8'b00011001; // 3379 :  25 - 0x19
      13'hD34: dout  = 8'b00100101; // 3380 :  37 - 0x25
      13'hD35: dout  = 8'b00100101; // 3381 :  37 - 0x25
      13'hD36: dout  = 8'b00011000; // 3382 :  24 - 0x18
      13'hD37: dout  = 8'b00000000; // 3383 :   0 - 0x0
      13'hD38: dout  = 8'b00000000; // 3384 :   0 - 0x0
      13'hD39: dout  = 8'b00000000; // 3385 :   0 - 0x0
      13'hD3A: dout  = 8'b00000000; // 3386 :   0 - 0x0
      13'hD3B: dout  = 8'b00000000; // 3387 :   0 - 0x0
      13'hD3C: dout  = 8'b00000000; // 3388 :   0 - 0x0
      13'hD3D: dout  = 8'b00000000; // 3389 :   0 - 0x0
      13'hD3E: dout  = 8'b00000000; // 3390 :   0 - 0x0
      13'hD3F: dout  = 8'b00000000; // 3391 :   0 - 0x0
      13'hD40: dout  = 8'b11000110; // 3392 : 198 - 0xc6 -- Sprite 0xd4
      13'hD41: dout  = 8'b00101001; // 3393 :  41 - 0x29
      13'hD42: dout  = 8'b00101001; // 3394 :  41 - 0x29
      13'hD43: dout  = 8'b00101001; // 3395 :  41 - 0x29
      13'hD44: dout  = 8'b00101001; // 3396 :  41 - 0x29
      13'hD45: dout  = 8'b00101001; // 3397 :  41 - 0x29
      13'hD46: dout  = 8'b11000110; // 3398 : 198 - 0xc6
      13'hD47: dout  = 8'b00000000; // 3399 :   0 - 0x0
      13'hD48: dout  = 8'b00000000; // 3400 :   0 - 0x0
      13'hD49: dout  = 8'b00000000; // 3401 :   0 - 0x0
      13'hD4A: dout  = 8'b00000000; // 3402 :   0 - 0x0
      13'hD4B: dout  = 8'b00000000; // 3403 :   0 - 0x0
      13'hD4C: dout  = 8'b00000000; // 3404 :   0 - 0x0
      13'hD4D: dout  = 8'b00000000; // 3405 :   0 - 0x0
      13'hD4E: dout  = 8'b00000000; // 3406 :   0 - 0x0
      13'hD4F: dout  = 8'b00000000; // 3407 :   0 - 0x0
      13'hD50: dout  = 8'b00000000; // 3408 :   0 - 0x0 -- Sprite 0xd5
      13'hD51: dout  = 8'b00000000; // 3409 :   0 - 0x0
      13'hD52: dout  = 8'b00000000; // 3410 :   0 - 0x0
      13'hD53: dout  = 8'b00000000; // 3411 :   0 - 0x0
      13'hD54: dout  = 8'b00000000; // 3412 :   0 - 0x0
      13'hD55: dout  = 8'b00000000; // 3413 :   0 - 0x0
      13'hD56: dout  = 8'b00000000; // 3414 :   0 - 0x0
      13'hD57: dout  = 8'b00000000; // 3415 :   0 - 0x0
      13'hD58: dout  = 8'b00000000; // 3416 :   0 - 0x0
      13'hD59: dout  = 8'b00000000; // 3417 :   0 - 0x0
      13'hD5A: dout  = 8'b00000000; // 3418 :   0 - 0x0
      13'hD5B: dout  = 8'b00000001; // 3419 :   1 - 0x1
      13'hD5C: dout  = 8'b00000011; // 3420 :   3 - 0x3
      13'hD5D: dout  = 8'b01100011; // 3421 :  99 - 0x63
      13'hD5E: dout  = 8'b00110001; // 3422 :  49 - 0x31
      13'hD5F: dout  = 8'b00011111; // 3423 :  31 - 0x1f
      13'hD60: dout  = 8'b00000000; // 3424 :   0 - 0x0 -- Sprite 0xd6
      13'hD61: dout  = 8'b00000000; // 3425 :   0 - 0x0
      13'hD62: dout  = 8'b00000000; // 3426 :   0 - 0x0
      13'hD63: dout  = 8'b00000000; // 3427 :   0 - 0x0
      13'hD64: dout  = 8'b00111100; // 3428 :  60 - 0x3c
      13'hD65: dout  = 8'b10110110; // 3429 : 182 - 0xb6
      13'hD66: dout  = 8'b01111100; // 3430 : 124 - 0x7c
      13'hD67: dout  = 8'b11111000; // 3431 : 248 - 0xf8
      13'hD68: dout  = 8'b00000000; // 3432 :   0 - 0x0
      13'hD69: dout  = 8'b00000000; // 3433 :   0 - 0x0
      13'hD6A: dout  = 8'b11111100; // 3434 : 252 - 0xfc
      13'hD6B: dout  = 8'b11111110; // 3435 : 254 - 0xfe
      13'hD6C: dout  = 8'b11000000; // 3436 : 192 - 0xc0
      13'hD6D: dout  = 8'b01000000; // 3437 :  64 - 0x40
      13'hD6E: dout  = 8'b10000000; // 3438 : 128 - 0x80
      13'hD6F: dout  = 8'b00000000; // 3439 :   0 - 0x0
      13'hD70: dout  = 8'b00000011; // 3440 :   3 - 0x3 -- Sprite 0xd7
      13'hD71: dout  = 8'b00000011; // 3441 :   3 - 0x3
      13'hD72: dout  = 8'b00000011; // 3442 :   3 - 0x3
      13'hD73: dout  = 8'b00000111; // 3443 :   7 - 0x7
      13'hD74: dout  = 8'b00001100; // 3444 :  12 - 0xc
      13'hD75: dout  = 8'b00011011; // 3445 :  27 - 0x1b
      13'hD76: dout  = 8'b01110111; // 3446 : 119 - 0x77
      13'hD77: dout  = 8'b00000111; // 3447 :   7 - 0x7
      13'hD78: dout  = 8'b01111111; // 3448 : 127 - 0x7f
      13'hD79: dout  = 8'b00111111; // 3449 :  63 - 0x3f
      13'hD7A: dout  = 8'b01010011; // 3450 :  83 - 0x53
      13'hD7B: dout  = 8'b00000111; // 3451 :   7 - 0x7
      13'hD7C: dout  = 8'b00001100; // 3452 :  12 - 0xc
      13'hD7D: dout  = 8'b00011011; // 3453 :  27 - 0x1b
      13'hD7E: dout  = 8'b00000111; // 3454 :   7 - 0x7
      13'hD7F: dout  = 8'b00000111; // 3455 :   7 - 0x7
      13'hD80: dout  = 8'b00001111; // 3456 :  15 - 0xf -- Sprite 0xd8
      13'hD81: dout  = 8'b00001111; // 3457 :  15 - 0xf
      13'hD82: dout  = 8'b00011111; // 3458 :  31 - 0x1f
      13'hD83: dout  = 8'b00111111; // 3459 :  63 - 0x3f
      13'hD84: dout  = 8'b01111111; // 3460 : 127 - 0x7f
      13'hD85: dout  = 8'b00111111; // 3461 :  63 - 0x3f
      13'hD86: dout  = 8'b00000000; // 3462 :   0 - 0x0
      13'hD87: dout  = 8'b00000000; // 3463 :   0 - 0x0
      13'hD88: dout  = 8'b00001111; // 3464 :  15 - 0xf
      13'hD89: dout  = 8'b00001111; // 3465 :  15 - 0xf
      13'hD8A: dout  = 8'b00000011; // 3466 :   3 - 0x3
      13'hD8B: dout  = 8'b00111000; // 3467 :  56 - 0x38
      13'hD8C: dout  = 8'b00111111; // 3468 :  63 - 0x3f
      13'hD8D: dout  = 8'b00001110; // 3469 :  14 - 0xe
      13'hD8E: dout  = 8'b00011100; // 3470 :  28 - 0x1c
      13'hD8F: dout  = 8'b00001110; // 3471 :  14 - 0xe
      13'hD90: dout  = 8'b11100000; // 3472 : 224 - 0xe0 -- Sprite 0xd9
      13'hD91: dout  = 8'b11110000; // 3473 : 240 - 0xf0
      13'hD92: dout  = 8'b11110000; // 3474 : 240 - 0xf0
      13'hD93: dout  = 8'b11110000; // 3475 : 240 - 0xf0
      13'hD94: dout  = 8'b00011000; // 3476 :  24 - 0x18
      13'hD95: dout  = 8'b11111100; // 3477 : 252 - 0xfc
      13'hD96: dout  = 8'b11111100; // 3478 : 252 - 0xfc
      13'hD97: dout  = 8'b11111100; // 3479 : 252 - 0xfc
      13'hD98: dout  = 8'b00000000; // 3480 :   0 - 0x0
      13'hD99: dout  = 8'b10010000; // 3481 : 144 - 0x90
      13'hD9A: dout  = 8'b11110000; // 3482 : 240 - 0xf0
      13'hD9B: dout  = 8'b11110000; // 3483 : 240 - 0xf0
      13'hD9C: dout  = 8'b00011000; // 3484 :  24 - 0x18
      13'hD9D: dout  = 8'b11111100; // 3485 : 252 - 0xfc
      13'hD9E: dout  = 8'b11110000; // 3486 : 240 - 0xf0
      13'hD9F: dout  = 8'b11111000; // 3487 : 248 - 0xf8
      13'hDA0: dout  = 8'b11111000; // 3488 : 248 - 0xf8 -- Sprite 0xda
      13'hDA1: dout  = 8'b11111100; // 3489 : 252 - 0xfc
      13'hDA2: dout  = 8'b11111111; // 3490 : 255 - 0xff
      13'hDA3: dout  = 8'b11111111; // 3491 : 255 - 0xff
      13'hDA4: dout  = 8'b11111110; // 3492 : 254 - 0xfe
      13'hDA5: dout  = 8'b11110000; // 3493 : 240 - 0xf0
      13'hDA6: dout  = 8'b00000000; // 3494 :   0 - 0x0
      13'hDA7: dout  = 8'b00000000; // 3495 :   0 - 0x0
      13'hDA8: dout  = 8'b11111000; // 3496 : 248 - 0xf8
      13'hDA9: dout  = 8'b11110000; // 3497 : 240 - 0xf0
      13'hDAA: dout  = 8'b10000111; // 3498 : 135 - 0x87
      13'hDAB: dout  = 8'b00111101; // 3499 :  61 - 0x3d
      13'hDAC: dout  = 8'b11111110; // 3500 : 254 - 0xfe
      13'hDAD: dout  = 8'b00011100; // 3501 :  28 - 0x1c
      13'hDAE: dout  = 8'b00001000; // 3502 :   8 - 0x8
      13'hDAF: dout  = 8'b00000000; // 3503 :   0 - 0x0
      13'hDB0: dout  = 8'b00000011; // 3504 :   3 - 0x3 -- Sprite 0xdb
      13'hDB1: dout  = 8'b00000011; // 3505 :   3 - 0x3
      13'hDB2: dout  = 8'b00000011; // 3506 :   3 - 0x3
      13'hDB3: dout  = 8'b00000011; // 3507 :   3 - 0x3
      13'hDB4: dout  = 8'b00000001; // 3508 :   1 - 0x1
      13'hDB5: dout  = 8'b00000000; // 3509 :   0 - 0x0
      13'hDB6: dout  = 8'b00000111; // 3510 :   7 - 0x7
      13'hDB7: dout  = 8'b00011111; // 3511 :  31 - 0x1f
      13'hDB8: dout  = 8'b01111111; // 3512 : 127 - 0x7f
      13'hDB9: dout  = 8'b00111111; // 3513 :  63 - 0x3f
      13'hDBA: dout  = 8'b01010011; // 3514 :  83 - 0x53
      13'hDBB: dout  = 8'b00000011; // 3515 :   3 - 0x3
      13'hDBC: dout  = 8'b00000001; // 3516 :   1 - 0x1
      13'hDBD: dout  = 8'b00000000; // 3517 :   0 - 0x0
      13'hDBE: dout  = 8'b00000111; // 3518 :   7 - 0x7
      13'hDBF: dout  = 8'b00011111; // 3519 :  31 - 0x1f
      13'hDC0: dout  = 8'b11111111; // 3520 : 255 - 0xff -- Sprite 0xdc
      13'hDC1: dout  = 8'b11111111; // 3521 : 255 - 0xff
      13'hDC2: dout  = 8'b01111111; // 3522 : 127 - 0x7f
      13'hDC3: dout  = 8'b00111111; // 3523 :  63 - 0x3f
      13'hDC4: dout  = 8'b00001111; // 3524 :  15 - 0xf
      13'hDC5: dout  = 8'b00000011; // 3525 :   3 - 0x3
      13'hDC6: dout  = 8'b00000000; // 3526 :   0 - 0x0
      13'hDC7: dout  = 8'b00000000; // 3527 :   0 - 0x0
      13'hDC8: dout  = 8'b11001111; // 3528 : 207 - 0xcf
      13'hDC9: dout  = 8'b01100011; // 3529 :  99 - 0x63
      13'hDCA: dout  = 8'b00111000; // 3530 :  56 - 0x38
      13'hDCB: dout  = 8'b00111110; // 3531 :  62 - 0x3e
      13'hDCC: dout  = 8'b01111011; // 3532 : 123 - 0x7b
      13'hDCD: dout  = 8'b00110000; // 3533 :  48 - 0x30
      13'hDCE: dout  = 8'b00011000; // 3534 :  24 - 0x18
      13'hDCF: dout  = 8'b00000000; // 3535 :   0 - 0x0
      13'hDD0: dout  = 8'b11100000; // 3536 : 224 - 0xe0 -- Sprite 0xdd
      13'hDD1: dout  = 8'b11110000; // 3537 : 240 - 0xf0
      13'hDD2: dout  = 8'b11110000; // 3538 : 240 - 0xf0
      13'hDD3: dout  = 8'b11100000; // 3539 : 224 - 0xe0
      13'hDD4: dout  = 8'b11111110; // 3540 : 254 - 0xfe
      13'hDD5: dout  = 8'b00111100; // 3541 :  60 - 0x3c
      13'hDD6: dout  = 8'b11110000; // 3542 : 240 - 0xf0
      13'hDD7: dout  = 8'b11111100; // 3543 : 252 - 0xfc
      13'hDD8: dout  = 8'b00000000; // 3544 :   0 - 0x0
      13'hDD9: dout  = 8'b10010000; // 3545 : 144 - 0x90
      13'hDDA: dout  = 8'b11110000; // 3546 : 240 - 0xf0
      13'hDDB: dout  = 8'b11100000; // 3547 : 224 - 0xe0
      13'hDDC: dout  = 8'b11111000; // 3548 : 248 - 0xf8
      13'hDDD: dout  = 8'b00111000; // 3549 :  56 - 0x38
      13'hDDE: dout  = 8'b11110000; // 3550 : 240 - 0xf0
      13'hDDF: dout  = 8'b11110000; // 3551 : 240 - 0xf0
      13'hDE0: dout  = 8'b11111100; // 3552 : 252 - 0xfc -- Sprite 0xde
      13'hDE1: dout  = 8'b11111000; // 3553 : 248 - 0xf8
      13'hDE2: dout  = 8'b11111000; // 3554 : 248 - 0xf8
      13'hDE3: dout  = 8'b11111000; // 3555 : 248 - 0xf8
      13'hDE4: dout  = 8'b11111000; // 3556 : 248 - 0xf8
      13'hDE5: dout  = 8'b11111000; // 3557 : 248 - 0xf8
      13'hDE6: dout  = 8'b11111000; // 3558 : 248 - 0xf8
      13'hDE7: dout  = 8'b00000000; // 3559 :   0 - 0x0
      13'hDE8: dout  = 8'b11111000; // 3560 : 248 - 0xf8
      13'hDE9: dout  = 8'b11111000; // 3561 : 248 - 0xf8
      13'hDEA: dout  = 8'b11111000; // 3562 : 248 - 0xf8
      13'hDEB: dout  = 8'b00111000; // 3563 :  56 - 0x38
      13'hDEC: dout  = 8'b10000000; // 3564 : 128 - 0x80
      13'hDED: dout  = 8'b11111000; // 3565 : 248 - 0xf8
      13'hDEE: dout  = 8'b00000000; // 3566 :   0 - 0x0
      13'hDEF: dout  = 8'b01011100; // 3567 :  92 - 0x5c
      13'hDF0: dout  = 8'b11111111; // 3568 : 255 - 0xff -- Sprite 0xdf
      13'hDF1: dout  = 8'b11111111; // 3569 : 255 - 0xff
      13'hDF2: dout  = 8'b11111111; // 3570 : 255 - 0xff
      13'hDF3: dout  = 8'b11111111; // 3571 : 255 - 0xff
      13'hDF4: dout  = 8'b11111111; // 3572 : 255 - 0xff
      13'hDF5: dout  = 8'b11111111; // 3573 : 255 - 0xff
      13'hDF6: dout  = 8'b11111111; // 3574 : 255 - 0xff
      13'hDF7: dout  = 8'b11111111; // 3575 : 255 - 0xff
      13'hDF8: dout  = 8'b11111111; // 3576 : 255 - 0xff
      13'hDF9: dout  = 8'b11111111; // 3577 : 255 - 0xff
      13'hDFA: dout  = 8'b11111111; // 3578 : 255 - 0xff
      13'hDFB: dout  = 8'b11111111; // 3579 : 255 - 0xff
      13'hDFC: dout  = 8'b11111111; // 3580 : 255 - 0xff
      13'hDFD: dout  = 8'b11111111; // 3581 : 255 - 0xff
      13'hDFE: dout  = 8'b11111111; // 3582 : 255 - 0xff
      13'hDFF: dout  = 8'b11111111; // 3583 : 255 - 0xff
      13'hE00: dout  = 8'b11111111; // 3584 : 255 - 0xff -- Sprite 0xe0
      13'hE01: dout  = 8'b11111111; // 3585 : 255 - 0xff
      13'hE02: dout  = 8'b11111111; // 3586 : 255 - 0xff
      13'hE03: dout  = 8'b11111111; // 3587 : 255 - 0xff
      13'hE04: dout  = 8'b11111111; // 3588 : 255 - 0xff
      13'hE05: dout  = 8'b11111111; // 3589 : 255 - 0xff
      13'hE06: dout  = 8'b11111111; // 3590 : 255 - 0xff
      13'hE07: dout  = 8'b11111111; // 3591 : 255 - 0xff
      13'hE08: dout  = 8'b11111111; // 3592 : 255 - 0xff
      13'hE09: dout  = 8'b11111111; // 3593 : 255 - 0xff
      13'hE0A: dout  = 8'b11111111; // 3594 : 255 - 0xff
      13'hE0B: dout  = 8'b11111111; // 3595 : 255 - 0xff
      13'hE0C: dout  = 8'b11111111; // 3596 : 255 - 0xff
      13'hE0D: dout  = 8'b11111111; // 3597 : 255 - 0xff
      13'hE0E: dout  = 8'b11111111; // 3598 : 255 - 0xff
      13'hE0F: dout  = 8'b11111111; // 3599 : 255 - 0xff
      13'hE10: dout  = 8'b11111111; // 3600 : 255 - 0xff -- Sprite 0xe1
      13'hE11: dout  = 8'b11111111; // 3601 : 255 - 0xff
      13'hE12: dout  = 8'b11111111; // 3602 : 255 - 0xff
      13'hE13: dout  = 8'b11111111; // 3603 : 255 - 0xff
      13'hE14: dout  = 8'b11111111; // 3604 : 255 - 0xff
      13'hE15: dout  = 8'b11111111; // 3605 : 255 - 0xff
      13'hE16: dout  = 8'b11111111; // 3606 : 255 - 0xff
      13'hE17: dout  = 8'b11111111; // 3607 : 255 - 0xff
      13'hE18: dout  = 8'b11111111; // 3608 : 255 - 0xff
      13'hE19: dout  = 8'b11111111; // 3609 : 255 - 0xff
      13'hE1A: dout  = 8'b11111111; // 3610 : 255 - 0xff
      13'hE1B: dout  = 8'b11111111; // 3611 : 255 - 0xff
      13'hE1C: dout  = 8'b11111111; // 3612 : 255 - 0xff
      13'hE1D: dout  = 8'b11111111; // 3613 : 255 - 0xff
      13'hE1E: dout  = 8'b11111111; // 3614 : 255 - 0xff
      13'hE1F: dout  = 8'b11111111; // 3615 : 255 - 0xff
      13'hE20: dout  = 8'b11111111; // 3616 : 255 - 0xff -- Sprite 0xe2
      13'hE21: dout  = 8'b11111111; // 3617 : 255 - 0xff
      13'hE22: dout  = 8'b11111111; // 3618 : 255 - 0xff
      13'hE23: dout  = 8'b11111111; // 3619 : 255 - 0xff
      13'hE24: dout  = 8'b11111111; // 3620 : 255 - 0xff
      13'hE25: dout  = 8'b11111111; // 3621 : 255 - 0xff
      13'hE26: dout  = 8'b11111111; // 3622 : 255 - 0xff
      13'hE27: dout  = 8'b11111111; // 3623 : 255 - 0xff
      13'hE28: dout  = 8'b11111111; // 3624 : 255 - 0xff
      13'hE29: dout  = 8'b11111111; // 3625 : 255 - 0xff
      13'hE2A: dout  = 8'b11111111; // 3626 : 255 - 0xff
      13'hE2B: dout  = 8'b11111111; // 3627 : 255 - 0xff
      13'hE2C: dout  = 8'b11111111; // 3628 : 255 - 0xff
      13'hE2D: dout  = 8'b11111111; // 3629 : 255 - 0xff
      13'hE2E: dout  = 8'b11111111; // 3630 : 255 - 0xff
      13'hE2F: dout  = 8'b11111111; // 3631 : 255 - 0xff
      13'hE30: dout  = 8'b11111111; // 3632 : 255 - 0xff -- Sprite 0xe3
      13'hE31: dout  = 8'b11111111; // 3633 : 255 - 0xff
      13'hE32: dout  = 8'b11111111; // 3634 : 255 - 0xff
      13'hE33: dout  = 8'b11111111; // 3635 : 255 - 0xff
      13'hE34: dout  = 8'b11111111; // 3636 : 255 - 0xff
      13'hE35: dout  = 8'b11111111; // 3637 : 255 - 0xff
      13'hE36: dout  = 8'b11111111; // 3638 : 255 - 0xff
      13'hE37: dout  = 8'b11111111; // 3639 : 255 - 0xff
      13'hE38: dout  = 8'b11111111; // 3640 : 255 - 0xff
      13'hE39: dout  = 8'b11111111; // 3641 : 255 - 0xff
      13'hE3A: dout  = 8'b11111111; // 3642 : 255 - 0xff
      13'hE3B: dout  = 8'b11111111; // 3643 : 255 - 0xff
      13'hE3C: dout  = 8'b11111111; // 3644 : 255 - 0xff
      13'hE3D: dout  = 8'b11111111; // 3645 : 255 - 0xff
      13'hE3E: dout  = 8'b11111111; // 3646 : 255 - 0xff
      13'hE3F: dout  = 8'b11111111; // 3647 : 255 - 0xff
      13'hE40: dout  = 8'b11111111; // 3648 : 255 - 0xff -- Sprite 0xe4
      13'hE41: dout  = 8'b11111111; // 3649 : 255 - 0xff
      13'hE42: dout  = 8'b11111111; // 3650 : 255 - 0xff
      13'hE43: dout  = 8'b11111111; // 3651 : 255 - 0xff
      13'hE44: dout  = 8'b11111111; // 3652 : 255 - 0xff
      13'hE45: dout  = 8'b11111111; // 3653 : 255 - 0xff
      13'hE46: dout  = 8'b11111111; // 3654 : 255 - 0xff
      13'hE47: dout  = 8'b11111111; // 3655 : 255 - 0xff
      13'hE48: dout  = 8'b11111111; // 3656 : 255 - 0xff
      13'hE49: dout  = 8'b11111111; // 3657 : 255 - 0xff
      13'hE4A: dout  = 8'b11111111; // 3658 : 255 - 0xff
      13'hE4B: dout  = 8'b11111111; // 3659 : 255 - 0xff
      13'hE4C: dout  = 8'b11111111; // 3660 : 255 - 0xff
      13'hE4D: dout  = 8'b11111111; // 3661 : 255 - 0xff
      13'hE4E: dout  = 8'b11111111; // 3662 : 255 - 0xff
      13'hE4F: dout  = 8'b11111111; // 3663 : 255 - 0xff
      13'hE50: dout  = 8'b11111111; // 3664 : 255 - 0xff -- Sprite 0xe5
      13'hE51: dout  = 8'b11111111; // 3665 : 255 - 0xff
      13'hE52: dout  = 8'b11111111; // 3666 : 255 - 0xff
      13'hE53: dout  = 8'b11111111; // 3667 : 255 - 0xff
      13'hE54: dout  = 8'b11111111; // 3668 : 255 - 0xff
      13'hE55: dout  = 8'b11111111; // 3669 : 255 - 0xff
      13'hE56: dout  = 8'b11111111; // 3670 : 255 - 0xff
      13'hE57: dout  = 8'b11111111; // 3671 : 255 - 0xff
      13'hE58: dout  = 8'b11111111; // 3672 : 255 - 0xff
      13'hE59: dout  = 8'b11111111; // 3673 : 255 - 0xff
      13'hE5A: dout  = 8'b11111111; // 3674 : 255 - 0xff
      13'hE5B: dout  = 8'b11111111; // 3675 : 255 - 0xff
      13'hE5C: dout  = 8'b11111111; // 3676 : 255 - 0xff
      13'hE5D: dout  = 8'b11111111; // 3677 : 255 - 0xff
      13'hE5E: dout  = 8'b11111111; // 3678 : 255 - 0xff
      13'hE5F: dout  = 8'b11111111; // 3679 : 255 - 0xff
      13'hE60: dout  = 8'b11111111; // 3680 : 255 - 0xff -- Sprite 0xe6
      13'hE61: dout  = 8'b11111111; // 3681 : 255 - 0xff
      13'hE62: dout  = 8'b11111111; // 3682 : 255 - 0xff
      13'hE63: dout  = 8'b11111111; // 3683 : 255 - 0xff
      13'hE64: dout  = 8'b11111111; // 3684 : 255 - 0xff
      13'hE65: dout  = 8'b11111111; // 3685 : 255 - 0xff
      13'hE66: dout  = 8'b11111111; // 3686 : 255 - 0xff
      13'hE67: dout  = 8'b11111111; // 3687 : 255 - 0xff
      13'hE68: dout  = 8'b11111111; // 3688 : 255 - 0xff
      13'hE69: dout  = 8'b11111111; // 3689 : 255 - 0xff
      13'hE6A: dout  = 8'b11111111; // 3690 : 255 - 0xff
      13'hE6B: dout  = 8'b11111111; // 3691 : 255 - 0xff
      13'hE6C: dout  = 8'b11111111; // 3692 : 255 - 0xff
      13'hE6D: dout  = 8'b11111111; // 3693 : 255 - 0xff
      13'hE6E: dout  = 8'b11111111; // 3694 : 255 - 0xff
      13'hE6F: dout  = 8'b11111111; // 3695 : 255 - 0xff
      13'hE70: dout  = 8'b11111111; // 3696 : 255 - 0xff -- Sprite 0xe7
      13'hE71: dout  = 8'b11111111; // 3697 : 255 - 0xff
      13'hE72: dout  = 8'b11111111; // 3698 : 255 - 0xff
      13'hE73: dout  = 8'b11111111; // 3699 : 255 - 0xff
      13'hE74: dout  = 8'b11111111; // 3700 : 255 - 0xff
      13'hE75: dout  = 8'b11111111; // 3701 : 255 - 0xff
      13'hE76: dout  = 8'b11111111; // 3702 : 255 - 0xff
      13'hE77: dout  = 8'b11111111; // 3703 : 255 - 0xff
      13'hE78: dout  = 8'b11111111; // 3704 : 255 - 0xff
      13'hE79: dout  = 8'b11111111; // 3705 : 255 - 0xff
      13'hE7A: dout  = 8'b11111111; // 3706 : 255 - 0xff
      13'hE7B: dout  = 8'b11111111; // 3707 : 255 - 0xff
      13'hE7C: dout  = 8'b11111111; // 3708 : 255 - 0xff
      13'hE7D: dout  = 8'b11111111; // 3709 : 255 - 0xff
      13'hE7E: dout  = 8'b11111111; // 3710 : 255 - 0xff
      13'hE7F: dout  = 8'b11111111; // 3711 : 255 - 0xff
      13'hE80: dout  = 8'b11111111; // 3712 : 255 - 0xff -- Sprite 0xe8
      13'hE81: dout  = 8'b11111111; // 3713 : 255 - 0xff
      13'hE82: dout  = 8'b11111111; // 3714 : 255 - 0xff
      13'hE83: dout  = 8'b11111111; // 3715 : 255 - 0xff
      13'hE84: dout  = 8'b11111111; // 3716 : 255 - 0xff
      13'hE85: dout  = 8'b11111111; // 3717 : 255 - 0xff
      13'hE86: dout  = 8'b11111111; // 3718 : 255 - 0xff
      13'hE87: dout  = 8'b11111111; // 3719 : 255 - 0xff
      13'hE88: dout  = 8'b11111111; // 3720 : 255 - 0xff
      13'hE89: dout  = 8'b11111111; // 3721 : 255 - 0xff
      13'hE8A: dout  = 8'b11111111; // 3722 : 255 - 0xff
      13'hE8B: dout  = 8'b11111111; // 3723 : 255 - 0xff
      13'hE8C: dout  = 8'b11111111; // 3724 : 255 - 0xff
      13'hE8D: dout  = 8'b11111111; // 3725 : 255 - 0xff
      13'hE8E: dout  = 8'b11111111; // 3726 : 255 - 0xff
      13'hE8F: dout  = 8'b11111111; // 3727 : 255 - 0xff
      13'hE90: dout  = 8'b11111111; // 3728 : 255 - 0xff -- Sprite 0xe9
      13'hE91: dout  = 8'b11111111; // 3729 : 255 - 0xff
      13'hE92: dout  = 8'b11111111; // 3730 : 255 - 0xff
      13'hE93: dout  = 8'b11111111; // 3731 : 255 - 0xff
      13'hE94: dout  = 8'b11111111; // 3732 : 255 - 0xff
      13'hE95: dout  = 8'b11111111; // 3733 : 255 - 0xff
      13'hE96: dout  = 8'b11111111; // 3734 : 255 - 0xff
      13'hE97: dout  = 8'b11111111; // 3735 : 255 - 0xff
      13'hE98: dout  = 8'b11111111; // 3736 : 255 - 0xff
      13'hE99: dout  = 8'b11111111; // 3737 : 255 - 0xff
      13'hE9A: dout  = 8'b11111111; // 3738 : 255 - 0xff
      13'hE9B: dout  = 8'b11111111; // 3739 : 255 - 0xff
      13'hE9C: dout  = 8'b11111111; // 3740 : 255 - 0xff
      13'hE9D: dout  = 8'b11111111; // 3741 : 255 - 0xff
      13'hE9E: dout  = 8'b11111111; // 3742 : 255 - 0xff
      13'hE9F: dout  = 8'b11111111; // 3743 : 255 - 0xff
      13'hEA0: dout  = 8'b11111111; // 3744 : 255 - 0xff -- Sprite 0xea
      13'hEA1: dout  = 8'b11111111; // 3745 : 255 - 0xff
      13'hEA2: dout  = 8'b11111111; // 3746 : 255 - 0xff
      13'hEA3: dout  = 8'b11111111; // 3747 : 255 - 0xff
      13'hEA4: dout  = 8'b11111111; // 3748 : 255 - 0xff
      13'hEA5: dout  = 8'b11111111; // 3749 : 255 - 0xff
      13'hEA6: dout  = 8'b11111111; // 3750 : 255 - 0xff
      13'hEA7: dout  = 8'b11111111; // 3751 : 255 - 0xff
      13'hEA8: dout  = 8'b11111111; // 3752 : 255 - 0xff
      13'hEA9: dout  = 8'b11111111; // 3753 : 255 - 0xff
      13'hEAA: dout  = 8'b11111111; // 3754 : 255 - 0xff
      13'hEAB: dout  = 8'b11111111; // 3755 : 255 - 0xff
      13'hEAC: dout  = 8'b11111111; // 3756 : 255 - 0xff
      13'hEAD: dout  = 8'b11111111; // 3757 : 255 - 0xff
      13'hEAE: dout  = 8'b11111111; // 3758 : 255 - 0xff
      13'hEAF: dout  = 8'b11111111; // 3759 : 255 - 0xff
      13'hEB0: dout  = 8'b11111111; // 3760 : 255 - 0xff -- Sprite 0xeb
      13'hEB1: dout  = 8'b11111111; // 3761 : 255 - 0xff
      13'hEB2: dout  = 8'b11111111; // 3762 : 255 - 0xff
      13'hEB3: dout  = 8'b11111111; // 3763 : 255 - 0xff
      13'hEB4: dout  = 8'b11111111; // 3764 : 255 - 0xff
      13'hEB5: dout  = 8'b11111111; // 3765 : 255 - 0xff
      13'hEB6: dout  = 8'b11111111; // 3766 : 255 - 0xff
      13'hEB7: dout  = 8'b11111111; // 3767 : 255 - 0xff
      13'hEB8: dout  = 8'b11111111; // 3768 : 255 - 0xff
      13'hEB9: dout  = 8'b11111111; // 3769 : 255 - 0xff
      13'hEBA: dout  = 8'b11111111; // 3770 : 255 - 0xff
      13'hEBB: dout  = 8'b11111111; // 3771 : 255 - 0xff
      13'hEBC: dout  = 8'b11111111; // 3772 : 255 - 0xff
      13'hEBD: dout  = 8'b11111111; // 3773 : 255 - 0xff
      13'hEBE: dout  = 8'b11111111; // 3774 : 255 - 0xff
      13'hEBF: dout  = 8'b11111111; // 3775 : 255 - 0xff
      13'hEC0: dout  = 8'b00000000; // 3776 :   0 - 0x0 -- Sprite 0xec
      13'hEC1: dout  = 8'b00000001; // 3777 :   1 - 0x1
      13'hEC2: dout  = 8'b00000011; // 3778 :   3 - 0x3
      13'hEC3: dout  = 8'b00110011; // 3779 :  51 - 0x33
      13'hEC4: dout  = 8'b00011001; // 3780 :  25 - 0x19
      13'hEC5: dout  = 8'b00001111; // 3781 :  15 - 0xf
      13'hEC6: dout  = 8'b00111111; // 3782 :  63 - 0x3f
      13'hEC7: dout  = 8'b00011111; // 3783 :  31 - 0x1f
      13'hEC8: dout  = 8'b00000000; // 3784 :   0 - 0x0
      13'hEC9: dout  = 8'b00000001; // 3785 :   1 - 0x1
      13'hECA: dout  = 8'b00000011; // 3786 :   3 - 0x3
      13'hECB: dout  = 8'b00110011; // 3787 :  51 - 0x33
      13'hECC: dout  = 8'b00011001; // 3788 :  25 - 0x19
      13'hECD: dout  = 8'b00001111; // 3789 :  15 - 0xf
      13'hECE: dout  = 8'b00111111; // 3790 :  63 - 0x3f
      13'hECF: dout  = 8'b00011111; // 3791 :  31 - 0x1f
      13'hED0: dout  = 8'b00101011; // 3792 :  43 - 0x2b -- Sprite 0xed
      13'hED1: dout  = 8'b00000111; // 3793 :   7 - 0x7
      13'hED2: dout  = 8'b00000101; // 3794 :   5 - 0x5
      13'hED3: dout  = 8'b00001101; // 3795 :  13 - 0xd
      13'hED4: dout  = 8'b00001011; // 3796 :  11 - 0xb
      13'hED5: dout  = 8'b00011011; // 3797 :  27 - 0x1b
      13'hED6: dout  = 8'b00011011; // 3798 :  27 - 0x1b
      13'hED7: dout  = 8'b00111011; // 3799 :  59 - 0x3b
      13'hED8: dout  = 8'b00101011; // 3800 :  43 - 0x2b
      13'hED9: dout  = 8'b00000111; // 3801 :   7 - 0x7
      13'hEDA: dout  = 8'b00000101; // 3802 :   5 - 0x5
      13'hEDB: dout  = 8'b00001101; // 3803 :  13 - 0xd
      13'hEDC: dout  = 8'b00001011; // 3804 :  11 - 0xb
      13'hEDD: dout  = 8'b00011011; // 3805 :  27 - 0x1b
      13'hEDE: dout  = 8'b00011011; // 3806 :  27 - 0x1b
      13'hEDF: dout  = 8'b00000011; // 3807 :   3 - 0x3
      13'hEE0: dout  = 8'b00001001; // 3808 :   9 - 0x9 -- Sprite 0xee
      13'hEE1: dout  = 8'b00000000; // 3809 :   0 - 0x0
      13'hEE2: dout  = 8'b00000111; // 3810 :   7 - 0x7
      13'hEE3: dout  = 8'b00000111; // 3811 :   7 - 0x7
      13'hEE4: dout  = 8'b00001111; // 3812 :  15 - 0xf
      13'hEE5: dout  = 8'b00001101; // 3813 :  13 - 0xd
      13'hEE6: dout  = 8'b00000001; // 3814 :   1 - 0x1
      13'hEE7: dout  = 8'b00000000; // 3815 :   0 - 0x0
      13'hEE8: dout  = 8'b00000001; // 3816 :   1 - 0x1
      13'hEE9: dout  = 8'b00000000; // 3817 :   0 - 0x0
      13'hEEA: dout  = 8'b00000011; // 3818 :   3 - 0x3
      13'hEEB: dout  = 8'b00000101; // 3819 :   5 - 0x5
      13'hEEC: dout  = 8'b00001110; // 3820 :  14 - 0xe
      13'hEED: dout  = 8'b00001101; // 3821 :  13 - 0xd
      13'hEEE: dout  = 8'b00000001; // 3822 :   1 - 0x1
      13'hEEF: dout  = 8'b00000000; // 3823 :   0 - 0x0
      13'hEF0: dout  = 8'b11111000; // 3824 : 248 - 0xf8 -- Sprite 0xef
      13'hEF1: dout  = 8'b11111100; // 3825 : 252 - 0xfc
      13'hEF2: dout  = 8'b11111000; // 3826 : 248 - 0xf8
      13'hEF3: dout  = 8'b11101100; // 3827 : 236 - 0xec
      13'hEF4: dout  = 8'b11111000; // 3828 : 248 - 0xf8
      13'hEF5: dout  = 8'b11110000; // 3829 : 240 - 0xf0
      13'hEF6: dout  = 8'b11000000; // 3830 : 192 - 0xc0
      13'hEF7: dout  = 8'b11000000; // 3831 : 192 - 0xc0
      13'hEF8: dout  = 8'b11111000; // 3832 : 248 - 0xf8
      13'hEF9: dout  = 8'b11111100; // 3833 : 252 - 0xfc
      13'hEFA: dout  = 8'b11000000; // 3834 : 192 - 0xc0
      13'hEFB: dout  = 8'b01000000; // 3835 :  64 - 0x40
      13'hEFC: dout  = 8'b10000000; // 3836 : 128 - 0x80
      13'hEFD: dout  = 8'b10000000; // 3837 : 128 - 0x80
      13'hEFE: dout  = 8'b00000000; // 3838 :   0 - 0x0
      13'hEFF: dout  = 8'b10000000; // 3839 : 128 - 0x80
      13'hF00: dout  = 8'b11110000; // 3840 : 240 - 0xf0 -- Sprite 0xf0
      13'hF01: dout  = 8'b11111000; // 3841 : 248 - 0xf8
      13'hF02: dout  = 8'b11111000; // 3842 : 248 - 0xf8
      13'hF03: dout  = 8'b11101000; // 3843 : 232 - 0xe8
      13'hF04: dout  = 8'b11001100; // 3844 : 204 - 0xcc
      13'hF05: dout  = 8'b11100110; // 3845 : 230 - 0xe6
      13'hF06: dout  = 8'b11111011; // 3846 : 251 - 0xfb
      13'hF07: dout  = 8'b11111111; // 3847 : 255 - 0xff
      13'hF08: dout  = 8'b11010000; // 3848 : 208 - 0xd0
      13'hF09: dout  = 8'b11111000; // 3849 : 248 - 0xf8
      13'hF0A: dout  = 8'b11111000; // 3850 : 248 - 0xf8
      13'hF0B: dout  = 8'b11101000; // 3851 : 232 - 0xe8
      13'hF0C: dout  = 8'b11001100; // 3852 : 204 - 0xcc
      13'hF0D: dout  = 8'b11100110; // 3853 : 230 - 0xe6
      13'hF0E: dout  = 8'b11111000; // 3854 : 248 - 0xf8
      13'hF0F: dout  = 8'b11111110; // 3855 : 254 - 0xfe
      13'hF10: dout  = 8'b11111111; // 3856 : 255 - 0xff -- Sprite 0xf1
      13'hF11: dout  = 8'b11111110; // 3857 : 254 - 0xfe
      13'hF12: dout  = 8'b11111110; // 3858 : 254 - 0xfe
      13'hF13: dout  = 8'b11111110; // 3859 : 254 - 0xfe
      13'hF14: dout  = 8'b11111110; // 3860 : 254 - 0xfe
      13'hF15: dout  = 8'b10001111; // 3861 : 143 - 0x8f
      13'hF16: dout  = 8'b00000000; // 3862 :   0 - 0x0
      13'hF17: dout  = 8'b00000000; // 3863 :   0 - 0x0
      13'hF18: dout  = 8'b11111110; // 3864 : 254 - 0xfe
      13'hF19: dout  = 8'b11111110; // 3865 : 254 - 0xfe
      13'hF1A: dout  = 8'b00000110; // 3866 :   6 - 0x6
      13'hF1B: dout  = 8'b11111000; // 3867 : 248 - 0xf8
      13'hF1C: dout  = 8'b00001110; // 3868 :  14 - 0xe
      13'hF1D: dout  = 8'b10000000; // 3869 : 128 - 0x80
      13'hF1E: dout  = 8'b00000000; // 3870 :   0 - 0x0
      13'hF1F: dout  = 8'b00000000; // 3871 :   0 - 0x0
      13'hF20: dout  = 8'b00000001; // 3872 :   1 - 0x1 -- Sprite 0xf2
      13'hF21: dout  = 8'b00001111; // 3873 :  15 - 0xf
      13'hF22: dout  = 8'b00000000; // 3874 :   0 - 0x0
      13'hF23: dout  = 8'b00000000; // 3875 :   0 - 0x0
      13'hF24: dout  = 8'b00000100; // 3876 :   4 - 0x4
      13'hF25: dout  = 8'b00011110; // 3877 :  30 - 0x1e
      13'hF26: dout  = 8'b00000000; // 3878 :   0 - 0x0
      13'hF27: dout  = 8'b00000011; // 3879 :   3 - 0x3
      13'hF28: dout  = 8'b00000001; // 3880 :   1 - 0x1
      13'hF29: dout  = 8'b00001111; // 3881 :  15 - 0xf
      13'hF2A: dout  = 8'b00000111; // 3882 :   7 - 0x7
      13'hF2B: dout  = 8'b00011101; // 3883 :  29 - 0x1d
      13'hF2C: dout  = 8'b00111011; // 3884 :  59 - 0x3b
      13'hF2D: dout  = 8'b00000001; // 3885 :   1 - 0x1
      13'hF2E: dout  = 8'b00001111; // 3886 :  15 - 0xf
      13'hF2F: dout  = 8'b00000010; // 3887 :   2 - 0x2
      13'hF30: dout  = 8'b00000111; // 3888 :   7 - 0x7 -- Sprite 0xf3
      13'hF31: dout  = 8'b00001111; // 3889 :  15 - 0xf
      13'hF32: dout  = 8'b00011111; // 3890 :  31 - 0x1f
      13'hF33: dout  = 8'b00001111; // 3891 :  15 - 0xf
      13'hF34: dout  = 8'b00000111; // 3892 :   7 - 0x7
      13'hF35: dout  = 8'b00001111; // 3893 :  15 - 0xf
      13'hF36: dout  = 8'b00001111; // 3894 :  15 - 0xf
      13'hF37: dout  = 8'b00000011; // 3895 :   3 - 0x3
      13'hF38: dout  = 8'b00000010; // 3896 :   2 - 0x2
      13'hF39: dout  = 8'b00000011; // 3897 :   3 - 0x3
      13'hF3A: dout  = 8'b00000010; // 3898 :   2 - 0x2
      13'hF3B: dout  = 8'b01110111; // 3899 : 119 - 0x77
      13'hF3C: dout  = 8'b00010111; // 3900 :  23 - 0x17
      13'hF3D: dout  = 8'b00000001; // 3901 :   1 - 0x1
      13'hF3E: dout  = 8'b00000000; // 3902 :   0 - 0x0
      13'hF3F: dout  = 8'b00000000; // 3903 :   0 - 0x0
      13'hF40: dout  = 8'b11100000; // 3904 : 224 - 0xe0 -- Sprite 0xf4
      13'hF41: dout  = 8'b11110000; // 3905 : 240 - 0xf0
      13'hF42: dout  = 8'b11110000; // 3906 : 240 - 0xf0
      13'hF43: dout  = 8'b01001000; // 3907 :  72 - 0x48
      13'hF44: dout  = 8'b11001000; // 3908 : 200 - 0xc8
      13'hF45: dout  = 8'b10011100; // 3909 : 156 - 0x9c
      13'hF46: dout  = 8'b00000000; // 3910 :   0 - 0x0
      13'hF47: dout  = 8'b11110000; // 3911 : 240 - 0xf0
      13'hF48: dout  = 8'b11100000; // 3912 : 224 - 0xe0
      13'hF49: dout  = 8'b11110000; // 3913 : 240 - 0xf0
      13'hF4A: dout  = 8'b00000000; // 3914 :   0 - 0x0
      13'hF4B: dout  = 8'b10110000; // 3915 : 176 - 0xb0
      13'hF4C: dout  = 8'b00110000; // 3916 :  48 - 0x30
      13'hF4D: dout  = 8'b01100000; // 3917 :  96 - 0x60
      13'hF4E: dout  = 8'b11110000; // 3918 : 240 - 0xf0
      13'hF4F: dout  = 8'b00010000; // 3919 :  16 - 0x10
      13'hF50: dout  = 8'b11111000; // 3920 : 248 - 0xf8 -- Sprite 0xf5
      13'hF51: dout  = 8'b11111100; // 3921 : 252 - 0xfc
      13'hF52: dout  = 8'b11111100; // 3922 : 252 - 0xfc
      13'hF53: dout  = 8'b11111000; // 3923 : 248 - 0xf8
      13'hF54: dout  = 8'b11111000; // 3924 : 248 - 0xf8
      13'hF55: dout  = 8'b01111000; // 3925 : 120 - 0x78
      13'hF56: dout  = 8'b01110000; // 3926 : 112 - 0x70
      13'hF57: dout  = 8'b01100000; // 3927 :  96 - 0x60
      13'hF58: dout  = 8'b00110000; // 3928 :  48 - 0x30
      13'hF59: dout  = 8'b11110000; // 3929 : 240 - 0xf0
      13'hF5A: dout  = 8'b11010000; // 3930 : 208 - 0xd0
      13'hF5B: dout  = 8'b11111100; // 3931 : 252 - 0xfc
      13'hF5C: dout  = 8'b11111110; // 3932 : 254 - 0xfe
      13'hF5D: dout  = 8'b00001000; // 3933 :   8 - 0x8
      13'hF5E: dout  = 8'b00000000; // 3934 :   0 - 0x0
      13'hF5F: dout  = 8'b00000000; // 3935 :   0 - 0x0
      13'hF60: dout  = 8'b00000000; // 3936 :   0 - 0x0 -- Sprite 0xf6
      13'hF61: dout  = 8'b00000000; // 3937 :   0 - 0x0
      13'hF62: dout  = 8'b01111100; // 3938 : 124 - 0x7c
      13'hF63: dout  = 8'b10001010; // 3939 : 138 - 0x8a
      13'hF64: dout  = 8'b11111110; // 3940 : 254 - 0xfe
      13'hF65: dout  = 8'b11111110; // 3941 : 254 - 0xfe
      13'hF66: dout  = 8'b11111110; // 3942 : 254 - 0xfe
      13'hF67: dout  = 8'b11111110; // 3943 : 254 - 0xfe
      13'hF68: dout  = 8'b00000000; // 3944 :   0 - 0x0
      13'hF69: dout  = 8'b00010000; // 3945 :  16 - 0x10
      13'hF6A: dout  = 8'b00000000; // 3946 :   0 - 0x0
      13'hF6B: dout  = 8'b01110100; // 3947 : 116 - 0x74
      13'hF6C: dout  = 8'b00000000; // 3948 :   0 - 0x0
      13'hF6D: dout  = 8'b00000000; // 3949 :   0 - 0x0
      13'hF6E: dout  = 8'b00000000; // 3950 :   0 - 0x0
      13'hF6F: dout  = 8'b00000000; // 3951 :   0 - 0x0
      13'hF70: dout  = 8'b11111110; // 3952 : 254 - 0xfe -- Sprite 0xf7
      13'hF71: dout  = 8'b01111100; // 3953 : 124 - 0x7c
      13'hF72: dout  = 8'b00000000; // 3954 :   0 - 0x0
      13'hF73: dout  = 8'b00000000; // 3955 :   0 - 0x0
      13'hF74: dout  = 8'b00000000; // 3956 :   0 - 0x0
      13'hF75: dout  = 8'b00000000; // 3957 :   0 - 0x0
      13'hF76: dout  = 8'b00000000; // 3958 :   0 - 0x0
      13'hF77: dout  = 8'b00000000; // 3959 :   0 - 0x0
      13'hF78: dout  = 8'b00000000; // 3960 :   0 - 0x0
      13'hF79: dout  = 8'b00000000; // 3961 :   0 - 0x0
      13'hF7A: dout  = 8'b00010000; // 3962 :  16 - 0x10
      13'hF7B: dout  = 8'b00010000; // 3963 :  16 - 0x10
      13'hF7C: dout  = 8'b00010000; // 3964 :  16 - 0x10
      13'hF7D: dout  = 8'b00010000; // 3965 :  16 - 0x10
      13'hF7E: dout  = 8'b00010000; // 3966 :  16 - 0x10
      13'hF7F: dout  = 8'b00010000; // 3967 :  16 - 0x10
      13'hF80: dout  = 8'b00000111; // 3968 :   7 - 0x7 -- Sprite 0xf8
      13'hF81: dout  = 8'b00001011; // 3969 :  11 - 0xb
      13'hF82: dout  = 8'b00001111; // 3970 :  15 - 0xf
      13'hF83: dout  = 8'b00001011; // 3971 :  11 - 0xb
      13'hF84: dout  = 8'b00001011; // 3972 :  11 - 0xb
      13'hF85: dout  = 8'b00001011; // 3973 :  11 - 0xb
      13'hF86: dout  = 8'b00001011; // 3974 :  11 - 0xb
      13'hF87: dout  = 8'b00000111; // 3975 :   7 - 0x7
      13'hF88: dout  = 8'b00000000; // 3976 :   0 - 0x0
      13'hF89: dout  = 8'b00000100; // 3977 :   4 - 0x4
      13'hF8A: dout  = 8'b00000000; // 3978 :   0 - 0x0
      13'hF8B: dout  = 8'b00010100; // 3979 :  20 - 0x14
      13'hF8C: dout  = 8'b00000100; // 3980 :   4 - 0x4
      13'hF8D: dout  = 8'b00000100; // 3981 :   4 - 0x4
      13'hF8E: dout  = 8'b00000100; // 3982 :   4 - 0x4
      13'hF8F: dout  = 8'b00000000; // 3983 :   0 - 0x0
      13'hF90: dout  = 8'b11000000; // 3984 : 192 - 0xc0 -- Sprite 0xf9
      13'hF91: dout  = 8'b11100000; // 3985 : 224 - 0xe0
      13'hF92: dout  = 8'b11100000; // 3986 : 224 - 0xe0
      13'hF93: dout  = 8'b11100000; // 3987 : 224 - 0xe0
      13'hF94: dout  = 8'b11100000; // 3988 : 224 - 0xe0
      13'hF95: dout  = 8'b11100000; // 3989 : 224 - 0xe0
      13'hF96: dout  = 8'b11100000; // 3990 : 224 - 0xe0
      13'hF97: dout  = 8'b11000000; // 3991 : 192 - 0xc0
      13'hF98: dout  = 8'b00000000; // 3992 :   0 - 0x0
      13'hF99: dout  = 8'b00000000; // 3993 :   0 - 0x0
      13'hF9A: dout  = 8'b00000000; // 3994 :   0 - 0x0
      13'hF9B: dout  = 8'b00011111; // 3995 :  31 - 0x1f
      13'hF9C: dout  = 8'b00000000; // 3996 :   0 - 0x0
      13'hF9D: dout  = 8'b00000000; // 3997 :   0 - 0x0
      13'hF9E: dout  = 8'b00000000; // 3998 :   0 - 0x0
      13'hF9F: dout  = 8'b00000000; // 3999 :   0 - 0x0
      13'hFA0: dout  = 8'b00000011; // 4000 :   3 - 0x3 -- Sprite 0xfa
      13'hFA1: dout  = 8'b00000111; // 4001 :   7 - 0x7
      13'hFA2: dout  = 8'b00000111; // 4002 :   7 - 0x7
      13'hFA3: dout  = 8'b00000111; // 4003 :   7 - 0x7
      13'hFA4: dout  = 8'b00000111; // 4004 :   7 - 0x7
      13'hFA5: dout  = 8'b00000111; // 4005 :   7 - 0x7
      13'hFA6: dout  = 8'b00000111; // 4006 :   7 - 0x7
      13'hFA7: dout  = 8'b00000011; // 4007 :   3 - 0x3
      13'hFA8: dout  = 8'b00000000; // 4008 :   0 - 0x0
      13'hFA9: dout  = 8'b00000000; // 4009 :   0 - 0x0
      13'hFAA: dout  = 8'b00000000; // 4010 :   0 - 0x0
      13'hFAB: dout  = 8'b11111000; // 4011 : 248 - 0xf8
      13'hFAC: dout  = 8'b00000000; // 4012 :   0 - 0x0
      13'hFAD: dout  = 8'b00000000; // 4013 :   0 - 0x0
      13'hFAE: dout  = 8'b00000000; // 4014 :   0 - 0x0
      13'hFAF: dout  = 8'b00000000; // 4015 :   0 - 0x0
      13'hFB0: dout  = 8'b11100000; // 4016 : 224 - 0xe0 -- Sprite 0xfb
      13'hFB1: dout  = 8'b11010000; // 4017 : 208 - 0xd0
      13'hFB2: dout  = 8'b11010000; // 4018 : 208 - 0xd0
      13'hFB3: dout  = 8'b11010000; // 4019 : 208 - 0xd0
      13'hFB4: dout  = 8'b11010000; // 4020 : 208 - 0xd0
      13'hFB5: dout  = 8'b11110000; // 4021 : 240 - 0xf0
      13'hFB6: dout  = 8'b11010000; // 4022 : 208 - 0xd0
      13'hFB7: dout  = 8'b11100000; // 4023 : 224 - 0xe0
      13'hFB8: dout  = 8'b00000000; // 4024 :   0 - 0x0
      13'hFB9: dout  = 8'b00100000; // 4025 :  32 - 0x20
      13'hFBA: dout  = 8'b00100000; // 4026 :  32 - 0x20
      13'hFBB: dout  = 8'b00101000; // 4027 :  40 - 0x28
      13'hFBC: dout  = 8'b00100000; // 4028 :  32 - 0x20
      13'hFBD: dout  = 8'b00000000; // 4029 :   0 - 0x0
      13'hFBE: dout  = 8'b00100000; // 4030 :  32 - 0x20
      13'hFBF: dout  = 8'b00000000; // 4031 :   0 - 0x0
      13'hFC0: dout  = 8'b00000000; // 4032 :   0 - 0x0 -- Sprite 0xfc
      13'hFC1: dout  = 8'b00000001; // 4033 :   1 - 0x1
      13'hFC2: dout  = 8'b00010011; // 4034 :  19 - 0x13
      13'hFC3: dout  = 8'b00110111; // 4035 :  55 - 0x37
      13'hFC4: dout  = 8'b00111011; // 4036 :  59 - 0x3b
      13'hFC5: dout  = 8'b01110100; // 4037 : 116 - 0x74
      13'hFC6: dout  = 8'b01111010; // 4038 : 122 - 0x7a
      13'hFC7: dout  = 8'b00111110; // 4039 :  62 - 0x3e
      13'hFC8: dout  = 8'b00000000; // 4040 :   0 - 0x0
      13'hFC9: dout  = 8'b00000000; // 4041 :   0 - 0x0
      13'hFCA: dout  = 8'b00001000; // 4042 :   8 - 0x8
      13'hFCB: dout  = 8'b00100101; // 4043 :  37 - 0x25
      13'hFCC: dout  = 8'b00010010; // 4044 :  18 - 0x12
      13'hFCD: dout  = 8'b01010011; // 4045 :  83 - 0x53
      13'hFCE: dout  = 8'b00110011; // 4046 :  51 - 0x33
      13'hFCF: dout  = 8'b00111001; // 4047 :  57 - 0x39
      13'hFD0: dout  = 8'b11011000; // 4048 : 216 - 0xd8 -- Sprite 0xfd
      13'hFD1: dout  = 8'b10011000; // 4049 : 152 - 0x98
      13'hFD2: dout  = 8'b10101000; // 4050 : 168 - 0xa8
      13'hFD3: dout  = 8'b11011000; // 4051 : 216 - 0xd8
      13'hFD4: dout  = 8'b11011010; // 4052 : 218 - 0xda
      13'hFD5: dout  = 8'b01110100; // 4053 : 116 - 0x74
      13'hFD6: dout  = 8'b00101000; // 4054 :  40 - 0x28
      13'hFD7: dout  = 8'b11001000; // 4055 : 200 - 0xc8
      13'hFD8: dout  = 8'b00001000; // 4056 :   8 - 0x8
      13'hFD9: dout  = 8'b10000000; // 4057 : 128 - 0x80
      13'hFDA: dout  = 8'b00110000; // 4058 :  48 - 0x30
      13'hFDB: dout  = 8'b10011100; // 4059 : 156 - 0x9c
      13'hFDC: dout  = 8'b11001010; // 4060 : 202 - 0xca
      13'hFDD: dout  = 8'b10111000; // 4061 : 184 - 0xb8
      13'hFDE: dout  = 8'b10011000; // 4062 : 152 - 0x98
      13'hFDF: dout  = 8'b01111000; // 4063 : 120 - 0x78
      13'hFE0: dout  = 8'b00001000; // 4064 :   8 - 0x8 -- Sprite 0xfe
      13'hFE1: dout  = 8'b01011001; // 4065 :  89 - 0x59
      13'hFE2: dout  = 8'b00110000; // 4066 :  48 - 0x30
      13'hFE3: dout  = 8'b01110001; // 4067 : 113 - 0x71
      13'hFE4: dout  = 8'b01111001; // 4068 : 121 - 0x79
      13'hFE5: dout  = 8'b00101011; // 4069 :  43 - 0x2b
      13'hFE6: dout  = 8'b00110110; // 4070 :  54 - 0x36
      13'hFE7: dout  = 8'b00010110; // 4071 :  22 - 0x16
      13'hFE8: dout  = 8'b00000000; // 4072 :   0 - 0x0
      13'hFE9: dout  = 8'b00001000; // 4073 :   8 - 0x8
      13'hFEA: dout  = 8'b00000000; // 4074 :   0 - 0x0
      13'hFEB: dout  = 8'b01000000; // 4075 :  64 - 0x40
      13'hFEC: dout  = 8'b00000000; // 4076 :   0 - 0x0
      13'hFED: dout  = 8'b00110001; // 4077 :  49 - 0x31
      13'hFEE: dout  = 8'b00111101; // 4078 :  61 - 0x3d
      13'hFEF: dout  = 8'b00011001; // 4079 :  25 - 0x19
      13'hFF0: dout  = 8'b11000110; // 4080 : 198 - 0xc6 -- Sprite 0xff
      13'hFF1: dout  = 8'b11000100; // 4081 : 196 - 0xc4
      13'hFF2: dout  = 8'b11001100; // 4082 : 204 - 0xcc
      13'hFF3: dout  = 8'b11001100; // 4083 : 204 - 0xcc
      13'hFF4: dout  = 8'b10111000; // 4084 : 184 - 0xb8
      13'hFF5: dout  = 8'b01111100; // 4085 : 124 - 0x7c
      13'hFF6: dout  = 8'b11101100; // 4086 : 236 - 0xec
      13'hFF7: dout  = 8'b11001000; // 4087 : 200 - 0xc8
      13'hFF8: dout  = 8'b00000000; // 4088 :   0 - 0x0
      13'hFF9: dout  = 8'b10000000; // 4089 : 128 - 0x80
      13'hFFA: dout  = 8'b11000000; // 4090 : 192 - 0xc0
      13'hFFB: dout  = 8'b11000000; // 4091 : 192 - 0xc0
      13'hFFC: dout  = 8'b11000000; // 4092 : 192 - 0xc0
      13'hFFD: dout  = 8'b10001000; // 4093 : 136 - 0x88
      13'hFFE: dout  = 8'b10111000; // 4094 : 184 - 0xb8
      13'hFFF: dout  = 8'b10111000; // 4095 : 184 - 0xb8
          // Pattern Table 1---------
      13'h1000: dout  = 8'b00111000; // 4096 :  56 - 0x38 -- Background 0x0
      13'h1001: dout  = 8'b01001100; // 4097 :  76 - 0x4c
      13'h1002: dout  = 8'b11000110; // 4098 : 198 - 0xc6
      13'h1003: dout  = 8'b11000110; // 4099 : 198 - 0xc6
      13'h1004: dout  = 8'b11000110; // 4100 : 198 - 0xc6
      13'h1005: dout  = 8'b01100100; // 4101 : 100 - 0x64
      13'h1006: dout  = 8'b00111000; // 4102 :  56 - 0x38
      13'h1007: dout  = 8'b00000000; // 4103 :   0 - 0x0
      13'h1008: dout  = 8'b00000000; // 4104 :   0 - 0x0
      13'h1009: dout  = 8'b00000000; // 4105 :   0 - 0x0
      13'h100A: dout  = 8'b00000000; // 4106 :   0 - 0x0
      13'h100B: dout  = 8'b00000000; // 4107 :   0 - 0x0
      13'h100C: dout  = 8'b00000000; // 4108 :   0 - 0x0
      13'h100D: dout  = 8'b00000000; // 4109 :   0 - 0x0
      13'h100E: dout  = 8'b00000000; // 4110 :   0 - 0x0
      13'h100F: dout  = 8'b00000000; // 4111 :   0 - 0x0
      13'h1010: dout  = 8'b00011000; // 4112 :  24 - 0x18 -- Background 0x1
      13'h1011: dout  = 8'b00111000; // 4113 :  56 - 0x38
      13'h1012: dout  = 8'b00011000; // 4114 :  24 - 0x18
      13'h1013: dout  = 8'b00011000; // 4115 :  24 - 0x18
      13'h1014: dout  = 8'b00011000; // 4116 :  24 - 0x18
      13'h1015: dout  = 8'b00011000; // 4117 :  24 - 0x18
      13'h1016: dout  = 8'b01111110; // 4118 : 126 - 0x7e
      13'h1017: dout  = 8'b00000000; // 4119 :   0 - 0x0
      13'h1018: dout  = 8'b00000000; // 4120 :   0 - 0x0
      13'h1019: dout  = 8'b00000000; // 4121 :   0 - 0x0
      13'h101A: dout  = 8'b00000000; // 4122 :   0 - 0x0
      13'h101B: dout  = 8'b00000000; // 4123 :   0 - 0x0
      13'h101C: dout  = 8'b00000000; // 4124 :   0 - 0x0
      13'h101D: dout  = 8'b00000000; // 4125 :   0 - 0x0
      13'h101E: dout  = 8'b00000000; // 4126 :   0 - 0x0
      13'h101F: dout  = 8'b00000000; // 4127 :   0 - 0x0
      13'h1020: dout  = 8'b01111100; // 4128 : 124 - 0x7c -- Background 0x2
      13'h1021: dout  = 8'b11000110; // 4129 : 198 - 0xc6
      13'h1022: dout  = 8'b00001110; // 4130 :  14 - 0xe
      13'h1023: dout  = 8'b00111100; // 4131 :  60 - 0x3c
      13'h1024: dout  = 8'b01111000; // 4132 : 120 - 0x78
      13'h1025: dout  = 8'b11100000; // 4133 : 224 - 0xe0
      13'h1026: dout  = 8'b11111110; // 4134 : 254 - 0xfe
      13'h1027: dout  = 8'b00000000; // 4135 :   0 - 0x0
      13'h1028: dout  = 8'b00000000; // 4136 :   0 - 0x0
      13'h1029: dout  = 8'b00000000; // 4137 :   0 - 0x0
      13'h102A: dout  = 8'b00000000; // 4138 :   0 - 0x0
      13'h102B: dout  = 8'b00000000; // 4139 :   0 - 0x0
      13'h102C: dout  = 8'b00000000; // 4140 :   0 - 0x0
      13'h102D: dout  = 8'b00000000; // 4141 :   0 - 0x0
      13'h102E: dout  = 8'b00000000; // 4142 :   0 - 0x0
      13'h102F: dout  = 8'b00000000; // 4143 :   0 - 0x0
      13'h1030: dout  = 8'b01111110; // 4144 : 126 - 0x7e -- Background 0x3
      13'h1031: dout  = 8'b00001100; // 4145 :  12 - 0xc
      13'h1032: dout  = 8'b00011000; // 4146 :  24 - 0x18
      13'h1033: dout  = 8'b00111100; // 4147 :  60 - 0x3c
      13'h1034: dout  = 8'b00000110; // 4148 :   6 - 0x6
      13'h1035: dout  = 8'b11000110; // 4149 : 198 - 0xc6
      13'h1036: dout  = 8'b01111100; // 4150 : 124 - 0x7c
      13'h1037: dout  = 8'b00000000; // 4151 :   0 - 0x0
      13'h1038: dout  = 8'b00000000; // 4152 :   0 - 0x0
      13'h1039: dout  = 8'b00000000; // 4153 :   0 - 0x0
      13'h103A: dout  = 8'b00000000; // 4154 :   0 - 0x0
      13'h103B: dout  = 8'b00000000; // 4155 :   0 - 0x0
      13'h103C: dout  = 8'b00000000; // 4156 :   0 - 0x0
      13'h103D: dout  = 8'b00000000; // 4157 :   0 - 0x0
      13'h103E: dout  = 8'b00000000; // 4158 :   0 - 0x0
      13'h103F: dout  = 8'b00000000; // 4159 :   0 - 0x0
      13'h1040: dout  = 8'b00011100; // 4160 :  28 - 0x1c -- Background 0x4
      13'h1041: dout  = 8'b00111100; // 4161 :  60 - 0x3c
      13'h1042: dout  = 8'b01101100; // 4162 : 108 - 0x6c
      13'h1043: dout  = 8'b11001100; // 4163 : 204 - 0xcc
      13'h1044: dout  = 8'b11111110; // 4164 : 254 - 0xfe
      13'h1045: dout  = 8'b00001100; // 4165 :  12 - 0xc
      13'h1046: dout  = 8'b00001100; // 4166 :  12 - 0xc
      13'h1047: dout  = 8'b00000000; // 4167 :   0 - 0x0
      13'h1048: dout  = 8'b00000000; // 4168 :   0 - 0x0
      13'h1049: dout  = 8'b00000000; // 4169 :   0 - 0x0
      13'h104A: dout  = 8'b00000000; // 4170 :   0 - 0x0
      13'h104B: dout  = 8'b00000000; // 4171 :   0 - 0x0
      13'h104C: dout  = 8'b00000000; // 4172 :   0 - 0x0
      13'h104D: dout  = 8'b00000000; // 4173 :   0 - 0x0
      13'h104E: dout  = 8'b00000000; // 4174 :   0 - 0x0
      13'h104F: dout  = 8'b00000000; // 4175 :   0 - 0x0
      13'h1050: dout  = 8'b11111100; // 4176 : 252 - 0xfc -- Background 0x5
      13'h1051: dout  = 8'b11000000; // 4177 : 192 - 0xc0
      13'h1052: dout  = 8'b11111100; // 4178 : 252 - 0xfc
      13'h1053: dout  = 8'b00000110; // 4179 :   6 - 0x6
      13'h1054: dout  = 8'b00000110; // 4180 :   6 - 0x6
      13'h1055: dout  = 8'b11000110; // 4181 : 198 - 0xc6
      13'h1056: dout  = 8'b01111100; // 4182 : 124 - 0x7c
      13'h1057: dout  = 8'b00000000; // 4183 :   0 - 0x0
      13'h1058: dout  = 8'b00000000; // 4184 :   0 - 0x0
      13'h1059: dout  = 8'b00000000; // 4185 :   0 - 0x0
      13'h105A: dout  = 8'b00000000; // 4186 :   0 - 0x0
      13'h105B: dout  = 8'b00000000; // 4187 :   0 - 0x0
      13'h105C: dout  = 8'b00000000; // 4188 :   0 - 0x0
      13'h105D: dout  = 8'b00000000; // 4189 :   0 - 0x0
      13'h105E: dout  = 8'b00000000; // 4190 :   0 - 0x0
      13'h105F: dout  = 8'b00000000; // 4191 :   0 - 0x0
      13'h1060: dout  = 8'b00111100; // 4192 :  60 - 0x3c -- Background 0x6
      13'h1061: dout  = 8'b01100000; // 4193 :  96 - 0x60
      13'h1062: dout  = 8'b11000000; // 4194 : 192 - 0xc0
      13'h1063: dout  = 8'b11111100; // 4195 : 252 - 0xfc
      13'h1064: dout  = 8'b11000110; // 4196 : 198 - 0xc6
      13'h1065: dout  = 8'b11000110; // 4197 : 198 - 0xc6
      13'h1066: dout  = 8'b01111100; // 4198 : 124 - 0x7c
      13'h1067: dout  = 8'b00000000; // 4199 :   0 - 0x0
      13'h1068: dout  = 8'b00000000; // 4200 :   0 - 0x0
      13'h1069: dout  = 8'b00000000; // 4201 :   0 - 0x0
      13'h106A: dout  = 8'b00000000; // 4202 :   0 - 0x0
      13'h106B: dout  = 8'b00000000; // 4203 :   0 - 0x0
      13'h106C: dout  = 8'b00000000; // 4204 :   0 - 0x0
      13'h106D: dout  = 8'b00000000; // 4205 :   0 - 0x0
      13'h106E: dout  = 8'b00000000; // 4206 :   0 - 0x0
      13'h106F: dout  = 8'b00000000; // 4207 :   0 - 0x0
      13'h1070: dout  = 8'b11111110; // 4208 : 254 - 0xfe -- Background 0x7
      13'h1071: dout  = 8'b11000110; // 4209 : 198 - 0xc6
      13'h1072: dout  = 8'b00001100; // 4210 :  12 - 0xc
      13'h1073: dout  = 8'b00011000; // 4211 :  24 - 0x18
      13'h1074: dout  = 8'b00110000; // 4212 :  48 - 0x30
      13'h1075: dout  = 8'b00110000; // 4213 :  48 - 0x30
      13'h1076: dout  = 8'b00110000; // 4214 :  48 - 0x30
      13'h1077: dout  = 8'b00000000; // 4215 :   0 - 0x0
      13'h1078: dout  = 8'b00000000; // 4216 :   0 - 0x0
      13'h1079: dout  = 8'b00000000; // 4217 :   0 - 0x0
      13'h107A: dout  = 8'b00000000; // 4218 :   0 - 0x0
      13'h107B: dout  = 8'b00000000; // 4219 :   0 - 0x0
      13'h107C: dout  = 8'b00000000; // 4220 :   0 - 0x0
      13'h107D: dout  = 8'b00000000; // 4221 :   0 - 0x0
      13'h107E: dout  = 8'b00000000; // 4222 :   0 - 0x0
      13'h107F: dout  = 8'b00000000; // 4223 :   0 - 0x0
      13'h1080: dout  = 8'b01111000; // 4224 : 120 - 0x78 -- Background 0x8
      13'h1081: dout  = 8'b11000100; // 4225 : 196 - 0xc4
      13'h1082: dout  = 8'b11100100; // 4226 : 228 - 0xe4
      13'h1083: dout  = 8'b01111000; // 4227 : 120 - 0x78
      13'h1084: dout  = 8'b10000110; // 4228 : 134 - 0x86
      13'h1085: dout  = 8'b10000110; // 4229 : 134 - 0x86
      13'h1086: dout  = 8'b01111100; // 4230 : 124 - 0x7c
      13'h1087: dout  = 8'b00000000; // 4231 :   0 - 0x0
      13'h1088: dout  = 8'b00000000; // 4232 :   0 - 0x0
      13'h1089: dout  = 8'b00000000; // 4233 :   0 - 0x0
      13'h108A: dout  = 8'b00000000; // 4234 :   0 - 0x0
      13'h108B: dout  = 8'b00000000; // 4235 :   0 - 0x0
      13'h108C: dout  = 8'b00000000; // 4236 :   0 - 0x0
      13'h108D: dout  = 8'b00000000; // 4237 :   0 - 0x0
      13'h108E: dout  = 8'b00000000; // 4238 :   0 - 0x0
      13'h108F: dout  = 8'b00000000; // 4239 :   0 - 0x0
      13'h1090: dout  = 8'b01111100; // 4240 : 124 - 0x7c -- Background 0x9
      13'h1091: dout  = 8'b11000110; // 4241 : 198 - 0xc6
      13'h1092: dout  = 8'b11000110; // 4242 : 198 - 0xc6
      13'h1093: dout  = 8'b01111110; // 4243 : 126 - 0x7e
      13'h1094: dout  = 8'b00000110; // 4244 :   6 - 0x6
      13'h1095: dout  = 8'b00001100; // 4245 :  12 - 0xc
      13'h1096: dout  = 8'b01111000; // 4246 : 120 - 0x78
      13'h1097: dout  = 8'b00000000; // 4247 :   0 - 0x0
      13'h1098: dout  = 8'b00000000; // 4248 :   0 - 0x0
      13'h1099: dout  = 8'b00000000; // 4249 :   0 - 0x0
      13'h109A: dout  = 8'b00000000; // 4250 :   0 - 0x0
      13'h109B: dout  = 8'b00000000; // 4251 :   0 - 0x0
      13'h109C: dout  = 8'b00000000; // 4252 :   0 - 0x0
      13'h109D: dout  = 8'b00000000; // 4253 :   0 - 0x0
      13'h109E: dout  = 8'b00000000; // 4254 :   0 - 0x0
      13'h109F: dout  = 8'b00000000; // 4255 :   0 - 0x0
      13'h10A0: dout  = 8'b00111000; // 4256 :  56 - 0x38 -- Background 0xa
      13'h10A1: dout  = 8'b01101100; // 4257 : 108 - 0x6c
      13'h10A2: dout  = 8'b11000110; // 4258 : 198 - 0xc6
      13'h10A3: dout  = 8'b11000110; // 4259 : 198 - 0xc6
      13'h10A4: dout  = 8'b11111110; // 4260 : 254 - 0xfe
      13'h10A5: dout  = 8'b11000110; // 4261 : 198 - 0xc6
      13'h10A6: dout  = 8'b11000110; // 4262 : 198 - 0xc6
      13'h10A7: dout  = 8'b00000000; // 4263 :   0 - 0x0
      13'h10A8: dout  = 8'b00000000; // 4264 :   0 - 0x0
      13'h10A9: dout  = 8'b00000000; // 4265 :   0 - 0x0
      13'h10AA: dout  = 8'b00000000; // 4266 :   0 - 0x0
      13'h10AB: dout  = 8'b00000000; // 4267 :   0 - 0x0
      13'h10AC: dout  = 8'b00000000; // 4268 :   0 - 0x0
      13'h10AD: dout  = 8'b00000000; // 4269 :   0 - 0x0
      13'h10AE: dout  = 8'b00000000; // 4270 :   0 - 0x0
      13'h10AF: dout  = 8'b00000000; // 4271 :   0 - 0x0
      13'h10B0: dout  = 8'b11111100; // 4272 : 252 - 0xfc -- Background 0xb
      13'h10B1: dout  = 8'b11000110; // 4273 : 198 - 0xc6
      13'h10B2: dout  = 8'b11000110; // 4274 : 198 - 0xc6
      13'h10B3: dout  = 8'b11111100; // 4275 : 252 - 0xfc
      13'h10B4: dout  = 8'b11000110; // 4276 : 198 - 0xc6
      13'h10B5: dout  = 8'b11000110; // 4277 : 198 - 0xc6
      13'h10B6: dout  = 8'b11111100; // 4278 : 252 - 0xfc
      13'h10B7: dout  = 8'b00000000; // 4279 :   0 - 0x0
      13'h10B8: dout  = 8'b00000000; // 4280 :   0 - 0x0
      13'h10B9: dout  = 8'b00000000; // 4281 :   0 - 0x0
      13'h10BA: dout  = 8'b00000000; // 4282 :   0 - 0x0
      13'h10BB: dout  = 8'b00000000; // 4283 :   0 - 0x0
      13'h10BC: dout  = 8'b00000000; // 4284 :   0 - 0x0
      13'h10BD: dout  = 8'b00000000; // 4285 :   0 - 0x0
      13'h10BE: dout  = 8'b00000000; // 4286 :   0 - 0x0
      13'h10BF: dout  = 8'b00000000; // 4287 :   0 - 0x0
      13'h10C0: dout  = 8'b00111100; // 4288 :  60 - 0x3c -- Background 0xc
      13'h10C1: dout  = 8'b01100110; // 4289 : 102 - 0x66
      13'h10C2: dout  = 8'b11000000; // 4290 : 192 - 0xc0
      13'h10C3: dout  = 8'b11000000; // 4291 : 192 - 0xc0
      13'h10C4: dout  = 8'b11000000; // 4292 : 192 - 0xc0
      13'h10C5: dout  = 8'b01100110; // 4293 : 102 - 0x66
      13'h10C6: dout  = 8'b00111100; // 4294 :  60 - 0x3c
      13'h10C7: dout  = 8'b00000000; // 4295 :   0 - 0x0
      13'h10C8: dout  = 8'b00000000; // 4296 :   0 - 0x0
      13'h10C9: dout  = 8'b00000000; // 4297 :   0 - 0x0
      13'h10CA: dout  = 8'b00000000; // 4298 :   0 - 0x0
      13'h10CB: dout  = 8'b00000000; // 4299 :   0 - 0x0
      13'h10CC: dout  = 8'b00000000; // 4300 :   0 - 0x0
      13'h10CD: dout  = 8'b00000000; // 4301 :   0 - 0x0
      13'h10CE: dout  = 8'b00000000; // 4302 :   0 - 0x0
      13'h10CF: dout  = 8'b00000000; // 4303 :   0 - 0x0
      13'h10D0: dout  = 8'b11111000; // 4304 : 248 - 0xf8 -- Background 0xd
      13'h10D1: dout  = 8'b11001100; // 4305 : 204 - 0xcc
      13'h10D2: dout  = 8'b11000110; // 4306 : 198 - 0xc6
      13'h10D3: dout  = 8'b11000110; // 4307 : 198 - 0xc6
      13'h10D4: dout  = 8'b11000110; // 4308 : 198 - 0xc6
      13'h10D5: dout  = 8'b11001100; // 4309 : 204 - 0xcc
      13'h10D6: dout  = 8'b11111000; // 4310 : 248 - 0xf8
      13'h10D7: dout  = 8'b00000000; // 4311 :   0 - 0x0
      13'h10D8: dout  = 8'b00000000; // 4312 :   0 - 0x0
      13'h10D9: dout  = 8'b00000000; // 4313 :   0 - 0x0
      13'h10DA: dout  = 8'b00000000; // 4314 :   0 - 0x0
      13'h10DB: dout  = 8'b00000000; // 4315 :   0 - 0x0
      13'h10DC: dout  = 8'b00000000; // 4316 :   0 - 0x0
      13'h10DD: dout  = 8'b00000000; // 4317 :   0 - 0x0
      13'h10DE: dout  = 8'b00000000; // 4318 :   0 - 0x0
      13'h10DF: dout  = 8'b00000000; // 4319 :   0 - 0x0
      13'h10E0: dout  = 8'b11111110; // 4320 : 254 - 0xfe -- Background 0xe
      13'h10E1: dout  = 8'b11000000; // 4321 : 192 - 0xc0
      13'h10E2: dout  = 8'b11000000; // 4322 : 192 - 0xc0
      13'h10E3: dout  = 8'b11111100; // 4323 : 252 - 0xfc
      13'h10E4: dout  = 8'b11000000; // 4324 : 192 - 0xc0
      13'h10E5: dout  = 8'b11000000; // 4325 : 192 - 0xc0
      13'h10E6: dout  = 8'b11111110; // 4326 : 254 - 0xfe
      13'h10E7: dout  = 8'b00000000; // 4327 :   0 - 0x0
      13'h10E8: dout  = 8'b00000000; // 4328 :   0 - 0x0
      13'h10E9: dout  = 8'b00000000; // 4329 :   0 - 0x0
      13'h10EA: dout  = 8'b00000000; // 4330 :   0 - 0x0
      13'h10EB: dout  = 8'b00000000; // 4331 :   0 - 0x0
      13'h10EC: dout  = 8'b00000000; // 4332 :   0 - 0x0
      13'h10ED: dout  = 8'b00000000; // 4333 :   0 - 0x0
      13'h10EE: dout  = 8'b00000000; // 4334 :   0 - 0x0
      13'h10EF: dout  = 8'b00000000; // 4335 :   0 - 0x0
      13'h10F0: dout  = 8'b11111110; // 4336 : 254 - 0xfe -- Background 0xf
      13'h10F1: dout  = 8'b11000000; // 4337 : 192 - 0xc0
      13'h10F2: dout  = 8'b11000000; // 4338 : 192 - 0xc0
      13'h10F3: dout  = 8'b11111100; // 4339 : 252 - 0xfc
      13'h10F4: dout  = 8'b11000000; // 4340 : 192 - 0xc0
      13'h10F5: dout  = 8'b11000000; // 4341 : 192 - 0xc0
      13'h10F6: dout  = 8'b11000000; // 4342 : 192 - 0xc0
      13'h10F7: dout  = 8'b00000000; // 4343 :   0 - 0x0
      13'h10F8: dout  = 8'b00000000; // 4344 :   0 - 0x0
      13'h10F9: dout  = 8'b00000000; // 4345 :   0 - 0x0
      13'h10FA: dout  = 8'b00000000; // 4346 :   0 - 0x0
      13'h10FB: dout  = 8'b00000000; // 4347 :   0 - 0x0
      13'h10FC: dout  = 8'b00000000; // 4348 :   0 - 0x0
      13'h10FD: dout  = 8'b00000000; // 4349 :   0 - 0x0
      13'h10FE: dout  = 8'b00000000; // 4350 :   0 - 0x0
      13'h10FF: dout  = 8'b00000000; // 4351 :   0 - 0x0
      13'h1100: dout  = 8'b00111110; // 4352 :  62 - 0x3e -- Background 0x10
      13'h1101: dout  = 8'b01100000; // 4353 :  96 - 0x60
      13'h1102: dout  = 8'b11000000; // 4354 : 192 - 0xc0
      13'h1103: dout  = 8'b11011110; // 4355 : 222 - 0xde
      13'h1104: dout  = 8'b11000110; // 4356 : 198 - 0xc6
      13'h1105: dout  = 8'b01100110; // 4357 : 102 - 0x66
      13'h1106: dout  = 8'b01111110; // 4358 : 126 - 0x7e
      13'h1107: dout  = 8'b00000000; // 4359 :   0 - 0x0
      13'h1108: dout  = 8'b00000000; // 4360 :   0 - 0x0
      13'h1109: dout  = 8'b00000000; // 4361 :   0 - 0x0
      13'h110A: dout  = 8'b00000000; // 4362 :   0 - 0x0
      13'h110B: dout  = 8'b00000000; // 4363 :   0 - 0x0
      13'h110C: dout  = 8'b00000000; // 4364 :   0 - 0x0
      13'h110D: dout  = 8'b00000000; // 4365 :   0 - 0x0
      13'h110E: dout  = 8'b00000000; // 4366 :   0 - 0x0
      13'h110F: dout  = 8'b00000000; // 4367 :   0 - 0x0
      13'h1110: dout  = 8'b11000110; // 4368 : 198 - 0xc6 -- Background 0x11
      13'h1111: dout  = 8'b11000110; // 4369 : 198 - 0xc6
      13'h1112: dout  = 8'b11000110; // 4370 : 198 - 0xc6
      13'h1113: dout  = 8'b11111110; // 4371 : 254 - 0xfe
      13'h1114: dout  = 8'b11000110; // 4372 : 198 - 0xc6
      13'h1115: dout  = 8'b11000110; // 4373 : 198 - 0xc6
      13'h1116: dout  = 8'b11000110; // 4374 : 198 - 0xc6
      13'h1117: dout  = 8'b00000000; // 4375 :   0 - 0x0
      13'h1118: dout  = 8'b00000000; // 4376 :   0 - 0x0
      13'h1119: dout  = 8'b00000000; // 4377 :   0 - 0x0
      13'h111A: dout  = 8'b00000000; // 4378 :   0 - 0x0
      13'h111B: dout  = 8'b00000000; // 4379 :   0 - 0x0
      13'h111C: dout  = 8'b00000000; // 4380 :   0 - 0x0
      13'h111D: dout  = 8'b00000000; // 4381 :   0 - 0x0
      13'h111E: dout  = 8'b00000000; // 4382 :   0 - 0x0
      13'h111F: dout  = 8'b00000000; // 4383 :   0 - 0x0
      13'h1120: dout  = 8'b01111110; // 4384 : 126 - 0x7e -- Background 0x12
      13'h1121: dout  = 8'b00011000; // 4385 :  24 - 0x18
      13'h1122: dout  = 8'b00011000; // 4386 :  24 - 0x18
      13'h1123: dout  = 8'b00011000; // 4387 :  24 - 0x18
      13'h1124: dout  = 8'b00011000; // 4388 :  24 - 0x18
      13'h1125: dout  = 8'b00011000; // 4389 :  24 - 0x18
      13'h1126: dout  = 8'b01111110; // 4390 : 126 - 0x7e
      13'h1127: dout  = 8'b00000000; // 4391 :   0 - 0x0
      13'h1128: dout  = 8'b00000000; // 4392 :   0 - 0x0
      13'h1129: dout  = 8'b00000000; // 4393 :   0 - 0x0
      13'h112A: dout  = 8'b00000000; // 4394 :   0 - 0x0
      13'h112B: dout  = 8'b00000000; // 4395 :   0 - 0x0
      13'h112C: dout  = 8'b00000000; // 4396 :   0 - 0x0
      13'h112D: dout  = 8'b00000000; // 4397 :   0 - 0x0
      13'h112E: dout  = 8'b00000000; // 4398 :   0 - 0x0
      13'h112F: dout  = 8'b00000000; // 4399 :   0 - 0x0
      13'h1130: dout  = 8'b00011110; // 4400 :  30 - 0x1e -- Background 0x13
      13'h1131: dout  = 8'b00000110; // 4401 :   6 - 0x6
      13'h1132: dout  = 8'b00000110; // 4402 :   6 - 0x6
      13'h1133: dout  = 8'b00000110; // 4403 :   6 - 0x6
      13'h1134: dout  = 8'b11000110; // 4404 : 198 - 0xc6
      13'h1135: dout  = 8'b11000110; // 4405 : 198 - 0xc6
      13'h1136: dout  = 8'b01111100; // 4406 : 124 - 0x7c
      13'h1137: dout  = 8'b00000000; // 4407 :   0 - 0x0
      13'h1138: dout  = 8'b00000000; // 4408 :   0 - 0x0
      13'h1139: dout  = 8'b00000000; // 4409 :   0 - 0x0
      13'h113A: dout  = 8'b00000000; // 4410 :   0 - 0x0
      13'h113B: dout  = 8'b00000000; // 4411 :   0 - 0x0
      13'h113C: dout  = 8'b00000000; // 4412 :   0 - 0x0
      13'h113D: dout  = 8'b00000000; // 4413 :   0 - 0x0
      13'h113E: dout  = 8'b00000000; // 4414 :   0 - 0x0
      13'h113F: dout  = 8'b00000000; // 4415 :   0 - 0x0
      13'h1140: dout  = 8'b11000110; // 4416 : 198 - 0xc6 -- Background 0x14
      13'h1141: dout  = 8'b11001100; // 4417 : 204 - 0xcc
      13'h1142: dout  = 8'b11011000; // 4418 : 216 - 0xd8
      13'h1143: dout  = 8'b11110000; // 4419 : 240 - 0xf0
      13'h1144: dout  = 8'b11111000; // 4420 : 248 - 0xf8
      13'h1145: dout  = 8'b11011100; // 4421 : 220 - 0xdc
      13'h1146: dout  = 8'b11001110; // 4422 : 206 - 0xce
      13'h1147: dout  = 8'b00000000; // 4423 :   0 - 0x0
      13'h1148: dout  = 8'b00000000; // 4424 :   0 - 0x0
      13'h1149: dout  = 8'b00000000; // 4425 :   0 - 0x0
      13'h114A: dout  = 8'b00000000; // 4426 :   0 - 0x0
      13'h114B: dout  = 8'b00000000; // 4427 :   0 - 0x0
      13'h114C: dout  = 8'b00000000; // 4428 :   0 - 0x0
      13'h114D: dout  = 8'b00000000; // 4429 :   0 - 0x0
      13'h114E: dout  = 8'b00000000; // 4430 :   0 - 0x0
      13'h114F: dout  = 8'b00000000; // 4431 :   0 - 0x0
      13'h1150: dout  = 8'b01100000; // 4432 :  96 - 0x60 -- Background 0x15
      13'h1151: dout  = 8'b01100000; // 4433 :  96 - 0x60
      13'h1152: dout  = 8'b01100000; // 4434 :  96 - 0x60
      13'h1153: dout  = 8'b01100000; // 4435 :  96 - 0x60
      13'h1154: dout  = 8'b01100000; // 4436 :  96 - 0x60
      13'h1155: dout  = 8'b01100000; // 4437 :  96 - 0x60
      13'h1156: dout  = 8'b01111110; // 4438 : 126 - 0x7e
      13'h1157: dout  = 8'b00000000; // 4439 :   0 - 0x0
      13'h1158: dout  = 8'b00000000; // 4440 :   0 - 0x0
      13'h1159: dout  = 8'b00000000; // 4441 :   0 - 0x0
      13'h115A: dout  = 8'b00000000; // 4442 :   0 - 0x0
      13'h115B: dout  = 8'b00000000; // 4443 :   0 - 0x0
      13'h115C: dout  = 8'b00000000; // 4444 :   0 - 0x0
      13'h115D: dout  = 8'b00000000; // 4445 :   0 - 0x0
      13'h115E: dout  = 8'b00000000; // 4446 :   0 - 0x0
      13'h115F: dout  = 8'b00000000; // 4447 :   0 - 0x0
      13'h1160: dout  = 8'b11000110; // 4448 : 198 - 0xc6 -- Background 0x16
      13'h1161: dout  = 8'b11101110; // 4449 : 238 - 0xee
      13'h1162: dout  = 8'b11111110; // 4450 : 254 - 0xfe
      13'h1163: dout  = 8'b11111110; // 4451 : 254 - 0xfe
      13'h1164: dout  = 8'b11010110; // 4452 : 214 - 0xd6
      13'h1165: dout  = 8'b11000110; // 4453 : 198 - 0xc6
      13'h1166: dout  = 8'b11000110; // 4454 : 198 - 0xc6
      13'h1167: dout  = 8'b00000000; // 4455 :   0 - 0x0
      13'h1168: dout  = 8'b00000000; // 4456 :   0 - 0x0
      13'h1169: dout  = 8'b00000000; // 4457 :   0 - 0x0
      13'h116A: dout  = 8'b00000000; // 4458 :   0 - 0x0
      13'h116B: dout  = 8'b00000000; // 4459 :   0 - 0x0
      13'h116C: dout  = 8'b00000000; // 4460 :   0 - 0x0
      13'h116D: dout  = 8'b00000000; // 4461 :   0 - 0x0
      13'h116E: dout  = 8'b00000000; // 4462 :   0 - 0x0
      13'h116F: dout  = 8'b00000000; // 4463 :   0 - 0x0
      13'h1170: dout  = 8'b11000110; // 4464 : 198 - 0xc6 -- Background 0x17
      13'h1171: dout  = 8'b11100110; // 4465 : 230 - 0xe6
      13'h1172: dout  = 8'b11110110; // 4466 : 246 - 0xf6
      13'h1173: dout  = 8'b11111110; // 4467 : 254 - 0xfe
      13'h1174: dout  = 8'b11011110; // 4468 : 222 - 0xde
      13'h1175: dout  = 8'b11001110; // 4469 : 206 - 0xce
      13'h1176: dout  = 8'b11000110; // 4470 : 198 - 0xc6
      13'h1177: dout  = 8'b00000000; // 4471 :   0 - 0x0
      13'h1178: dout  = 8'b00000000; // 4472 :   0 - 0x0
      13'h1179: dout  = 8'b00000000; // 4473 :   0 - 0x0
      13'h117A: dout  = 8'b00000000; // 4474 :   0 - 0x0
      13'h117B: dout  = 8'b00000000; // 4475 :   0 - 0x0
      13'h117C: dout  = 8'b00000000; // 4476 :   0 - 0x0
      13'h117D: dout  = 8'b00000000; // 4477 :   0 - 0x0
      13'h117E: dout  = 8'b00000000; // 4478 :   0 - 0x0
      13'h117F: dout  = 8'b00000000; // 4479 :   0 - 0x0
      13'h1180: dout  = 8'b01111100; // 4480 : 124 - 0x7c -- Background 0x18
      13'h1181: dout  = 8'b11000110; // 4481 : 198 - 0xc6
      13'h1182: dout  = 8'b11000110; // 4482 : 198 - 0xc6
      13'h1183: dout  = 8'b11000110; // 4483 : 198 - 0xc6
      13'h1184: dout  = 8'b11000110; // 4484 : 198 - 0xc6
      13'h1185: dout  = 8'b11000110; // 4485 : 198 - 0xc6
      13'h1186: dout  = 8'b01111100; // 4486 : 124 - 0x7c
      13'h1187: dout  = 8'b00000000; // 4487 :   0 - 0x0
      13'h1188: dout  = 8'b00000000; // 4488 :   0 - 0x0
      13'h1189: dout  = 8'b00000000; // 4489 :   0 - 0x0
      13'h118A: dout  = 8'b00000000; // 4490 :   0 - 0x0
      13'h118B: dout  = 8'b00000000; // 4491 :   0 - 0x0
      13'h118C: dout  = 8'b00000000; // 4492 :   0 - 0x0
      13'h118D: dout  = 8'b00000000; // 4493 :   0 - 0x0
      13'h118E: dout  = 8'b00000000; // 4494 :   0 - 0x0
      13'h118F: dout  = 8'b00000000; // 4495 :   0 - 0x0
      13'h1190: dout  = 8'b11111100; // 4496 : 252 - 0xfc -- Background 0x19
      13'h1191: dout  = 8'b11000110; // 4497 : 198 - 0xc6
      13'h1192: dout  = 8'b11000110; // 4498 : 198 - 0xc6
      13'h1193: dout  = 8'b11000110; // 4499 : 198 - 0xc6
      13'h1194: dout  = 8'b11111100; // 4500 : 252 - 0xfc
      13'h1195: dout  = 8'b11000000; // 4501 : 192 - 0xc0
      13'h1196: dout  = 8'b11000000; // 4502 : 192 - 0xc0
      13'h1197: dout  = 8'b00000000; // 4503 :   0 - 0x0
      13'h1198: dout  = 8'b00000000; // 4504 :   0 - 0x0
      13'h1199: dout  = 8'b00000000; // 4505 :   0 - 0x0
      13'h119A: dout  = 8'b00000000; // 4506 :   0 - 0x0
      13'h119B: dout  = 8'b00000000; // 4507 :   0 - 0x0
      13'h119C: dout  = 8'b00000000; // 4508 :   0 - 0x0
      13'h119D: dout  = 8'b00000000; // 4509 :   0 - 0x0
      13'h119E: dout  = 8'b00000000; // 4510 :   0 - 0x0
      13'h119F: dout  = 8'b00000000; // 4511 :   0 - 0x0
      13'h11A0: dout  = 8'b01111100; // 4512 : 124 - 0x7c -- Background 0x1a
      13'h11A1: dout  = 8'b11000110; // 4513 : 198 - 0xc6
      13'h11A2: dout  = 8'b11000110; // 4514 : 198 - 0xc6
      13'h11A3: dout  = 8'b11000110; // 4515 : 198 - 0xc6
      13'h11A4: dout  = 8'b11011110; // 4516 : 222 - 0xde
      13'h11A5: dout  = 8'b11001100; // 4517 : 204 - 0xcc
      13'h11A6: dout  = 8'b01111010; // 4518 : 122 - 0x7a
      13'h11A7: dout  = 8'b00000000; // 4519 :   0 - 0x0
      13'h11A8: dout  = 8'b00000000; // 4520 :   0 - 0x0
      13'h11A9: dout  = 8'b00000000; // 4521 :   0 - 0x0
      13'h11AA: dout  = 8'b00000000; // 4522 :   0 - 0x0
      13'h11AB: dout  = 8'b00000000; // 4523 :   0 - 0x0
      13'h11AC: dout  = 8'b00000000; // 4524 :   0 - 0x0
      13'h11AD: dout  = 8'b00000000; // 4525 :   0 - 0x0
      13'h11AE: dout  = 8'b00000000; // 4526 :   0 - 0x0
      13'h11AF: dout  = 8'b00000000; // 4527 :   0 - 0x0
      13'h11B0: dout  = 8'b11111100; // 4528 : 252 - 0xfc -- Background 0x1b
      13'h11B1: dout  = 8'b11000110; // 4529 : 198 - 0xc6
      13'h11B2: dout  = 8'b11000110; // 4530 : 198 - 0xc6
      13'h11B3: dout  = 8'b11001110; // 4531 : 206 - 0xce
      13'h11B4: dout  = 8'b11111000; // 4532 : 248 - 0xf8
      13'h11B5: dout  = 8'b11011100; // 4533 : 220 - 0xdc
      13'h11B6: dout  = 8'b11001110; // 4534 : 206 - 0xce
      13'h11B7: dout  = 8'b00000000; // 4535 :   0 - 0x0
      13'h11B8: dout  = 8'b00000000; // 4536 :   0 - 0x0
      13'h11B9: dout  = 8'b00000000; // 4537 :   0 - 0x0
      13'h11BA: dout  = 8'b00000000; // 4538 :   0 - 0x0
      13'h11BB: dout  = 8'b00000000; // 4539 :   0 - 0x0
      13'h11BC: dout  = 8'b00000000; // 4540 :   0 - 0x0
      13'h11BD: dout  = 8'b00000000; // 4541 :   0 - 0x0
      13'h11BE: dout  = 8'b00000000; // 4542 :   0 - 0x0
      13'h11BF: dout  = 8'b00000000; // 4543 :   0 - 0x0
      13'h11C0: dout  = 8'b01111000; // 4544 : 120 - 0x78 -- Background 0x1c
      13'h11C1: dout  = 8'b11001100; // 4545 : 204 - 0xcc
      13'h11C2: dout  = 8'b11000000; // 4546 : 192 - 0xc0
      13'h11C3: dout  = 8'b01111100; // 4547 : 124 - 0x7c
      13'h11C4: dout  = 8'b00000110; // 4548 :   6 - 0x6
      13'h11C5: dout  = 8'b11000110; // 4549 : 198 - 0xc6
      13'h11C6: dout  = 8'b01111100; // 4550 : 124 - 0x7c
      13'h11C7: dout  = 8'b00000000; // 4551 :   0 - 0x0
      13'h11C8: dout  = 8'b00000000; // 4552 :   0 - 0x0
      13'h11C9: dout  = 8'b00000000; // 4553 :   0 - 0x0
      13'h11CA: dout  = 8'b00000000; // 4554 :   0 - 0x0
      13'h11CB: dout  = 8'b00000000; // 4555 :   0 - 0x0
      13'h11CC: dout  = 8'b00000000; // 4556 :   0 - 0x0
      13'h11CD: dout  = 8'b00000000; // 4557 :   0 - 0x0
      13'h11CE: dout  = 8'b00000000; // 4558 :   0 - 0x0
      13'h11CF: dout  = 8'b00000000; // 4559 :   0 - 0x0
      13'h11D0: dout  = 8'b01111110; // 4560 : 126 - 0x7e -- Background 0x1d
      13'h11D1: dout  = 8'b00011000; // 4561 :  24 - 0x18
      13'h11D2: dout  = 8'b00011000; // 4562 :  24 - 0x18
      13'h11D3: dout  = 8'b00011000; // 4563 :  24 - 0x18
      13'h11D4: dout  = 8'b00011000; // 4564 :  24 - 0x18
      13'h11D5: dout  = 8'b00011000; // 4565 :  24 - 0x18
      13'h11D6: dout  = 8'b00011000; // 4566 :  24 - 0x18
      13'h11D7: dout  = 8'b00000000; // 4567 :   0 - 0x0
      13'h11D8: dout  = 8'b00000000; // 4568 :   0 - 0x0
      13'h11D9: dout  = 8'b00000000; // 4569 :   0 - 0x0
      13'h11DA: dout  = 8'b00000000; // 4570 :   0 - 0x0
      13'h11DB: dout  = 8'b00000000; // 4571 :   0 - 0x0
      13'h11DC: dout  = 8'b00000000; // 4572 :   0 - 0x0
      13'h11DD: dout  = 8'b00000000; // 4573 :   0 - 0x0
      13'h11DE: dout  = 8'b00000000; // 4574 :   0 - 0x0
      13'h11DF: dout  = 8'b00000000; // 4575 :   0 - 0x0
      13'h11E0: dout  = 8'b11000110; // 4576 : 198 - 0xc6 -- Background 0x1e
      13'h11E1: dout  = 8'b11000110; // 4577 : 198 - 0xc6
      13'h11E2: dout  = 8'b11000110; // 4578 : 198 - 0xc6
      13'h11E3: dout  = 8'b11000110; // 4579 : 198 - 0xc6
      13'h11E4: dout  = 8'b11000110; // 4580 : 198 - 0xc6
      13'h11E5: dout  = 8'b11000110; // 4581 : 198 - 0xc6
      13'h11E6: dout  = 8'b01111100; // 4582 : 124 - 0x7c
      13'h11E7: dout  = 8'b00000000; // 4583 :   0 - 0x0
      13'h11E8: dout  = 8'b00000000; // 4584 :   0 - 0x0
      13'h11E9: dout  = 8'b00000000; // 4585 :   0 - 0x0
      13'h11EA: dout  = 8'b00000000; // 4586 :   0 - 0x0
      13'h11EB: dout  = 8'b00000000; // 4587 :   0 - 0x0
      13'h11EC: dout  = 8'b00000000; // 4588 :   0 - 0x0
      13'h11ED: dout  = 8'b00000000; // 4589 :   0 - 0x0
      13'h11EE: dout  = 8'b00000000; // 4590 :   0 - 0x0
      13'h11EF: dout  = 8'b00000000; // 4591 :   0 - 0x0
      13'h11F0: dout  = 8'b11000110; // 4592 : 198 - 0xc6 -- Background 0x1f
      13'h11F1: dout  = 8'b11000110; // 4593 : 198 - 0xc6
      13'h11F2: dout  = 8'b11000110; // 4594 : 198 - 0xc6
      13'h11F3: dout  = 8'b11101110; // 4595 : 238 - 0xee
      13'h11F4: dout  = 8'b01111100; // 4596 : 124 - 0x7c
      13'h11F5: dout  = 8'b00111000; // 4597 :  56 - 0x38
      13'h11F6: dout  = 8'b00010000; // 4598 :  16 - 0x10
      13'h11F7: dout  = 8'b00000000; // 4599 :   0 - 0x0
      13'h11F8: dout  = 8'b00000000; // 4600 :   0 - 0x0
      13'h11F9: dout  = 8'b00000000; // 4601 :   0 - 0x0
      13'h11FA: dout  = 8'b00000000; // 4602 :   0 - 0x0
      13'h11FB: dout  = 8'b00000000; // 4603 :   0 - 0x0
      13'h11FC: dout  = 8'b00000000; // 4604 :   0 - 0x0
      13'h11FD: dout  = 8'b00000000; // 4605 :   0 - 0x0
      13'h11FE: dout  = 8'b00000000; // 4606 :   0 - 0x0
      13'h11FF: dout  = 8'b00000000; // 4607 :   0 - 0x0
      13'h1200: dout  = 8'b11000110; // 4608 : 198 - 0xc6 -- Background 0x20
      13'h1201: dout  = 8'b11000110; // 4609 : 198 - 0xc6
      13'h1202: dout  = 8'b11010110; // 4610 : 214 - 0xd6
      13'h1203: dout  = 8'b11111110; // 4611 : 254 - 0xfe
      13'h1204: dout  = 8'b11111110; // 4612 : 254 - 0xfe
      13'h1205: dout  = 8'b11101110; // 4613 : 238 - 0xee
      13'h1206: dout  = 8'b11000110; // 4614 : 198 - 0xc6
      13'h1207: dout  = 8'b00000000; // 4615 :   0 - 0x0
      13'h1208: dout  = 8'b00000000; // 4616 :   0 - 0x0
      13'h1209: dout  = 8'b00000000; // 4617 :   0 - 0x0
      13'h120A: dout  = 8'b00000000; // 4618 :   0 - 0x0
      13'h120B: dout  = 8'b00000000; // 4619 :   0 - 0x0
      13'h120C: dout  = 8'b00000000; // 4620 :   0 - 0x0
      13'h120D: dout  = 8'b00000000; // 4621 :   0 - 0x0
      13'h120E: dout  = 8'b00000000; // 4622 :   0 - 0x0
      13'h120F: dout  = 8'b00000000; // 4623 :   0 - 0x0
      13'h1210: dout  = 8'b11000110; // 4624 : 198 - 0xc6 -- Background 0x21
      13'h1211: dout  = 8'b11101110; // 4625 : 238 - 0xee
      13'h1212: dout  = 8'b01111100; // 4626 : 124 - 0x7c
      13'h1213: dout  = 8'b00111000; // 4627 :  56 - 0x38
      13'h1214: dout  = 8'b01111100; // 4628 : 124 - 0x7c
      13'h1215: dout  = 8'b11101110; // 4629 : 238 - 0xee
      13'h1216: dout  = 8'b11000110; // 4630 : 198 - 0xc6
      13'h1217: dout  = 8'b00000000; // 4631 :   0 - 0x0
      13'h1218: dout  = 8'b00000000; // 4632 :   0 - 0x0
      13'h1219: dout  = 8'b00000000; // 4633 :   0 - 0x0
      13'h121A: dout  = 8'b00000000; // 4634 :   0 - 0x0
      13'h121B: dout  = 8'b00000000; // 4635 :   0 - 0x0
      13'h121C: dout  = 8'b00000000; // 4636 :   0 - 0x0
      13'h121D: dout  = 8'b00000000; // 4637 :   0 - 0x0
      13'h121E: dout  = 8'b00000000; // 4638 :   0 - 0x0
      13'h121F: dout  = 8'b00000000; // 4639 :   0 - 0x0
      13'h1220: dout  = 8'b01100110; // 4640 : 102 - 0x66 -- Background 0x22
      13'h1221: dout  = 8'b01100110; // 4641 : 102 - 0x66
      13'h1222: dout  = 8'b01100110; // 4642 : 102 - 0x66
      13'h1223: dout  = 8'b00111100; // 4643 :  60 - 0x3c
      13'h1224: dout  = 8'b00011000; // 4644 :  24 - 0x18
      13'h1225: dout  = 8'b00011000; // 4645 :  24 - 0x18
      13'h1226: dout  = 8'b00011000; // 4646 :  24 - 0x18
      13'h1227: dout  = 8'b00000000; // 4647 :   0 - 0x0
      13'h1228: dout  = 8'b00000000; // 4648 :   0 - 0x0
      13'h1229: dout  = 8'b00000000; // 4649 :   0 - 0x0
      13'h122A: dout  = 8'b00000000; // 4650 :   0 - 0x0
      13'h122B: dout  = 8'b00000000; // 4651 :   0 - 0x0
      13'h122C: dout  = 8'b00000000; // 4652 :   0 - 0x0
      13'h122D: dout  = 8'b00000000; // 4653 :   0 - 0x0
      13'h122E: dout  = 8'b00000000; // 4654 :   0 - 0x0
      13'h122F: dout  = 8'b00000000; // 4655 :   0 - 0x0
      13'h1230: dout  = 8'b11111110; // 4656 : 254 - 0xfe -- Background 0x23
      13'h1231: dout  = 8'b00001110; // 4657 :  14 - 0xe
      13'h1232: dout  = 8'b00011100; // 4658 :  28 - 0x1c
      13'h1233: dout  = 8'b00111000; // 4659 :  56 - 0x38
      13'h1234: dout  = 8'b01110000; // 4660 : 112 - 0x70
      13'h1235: dout  = 8'b11100000; // 4661 : 224 - 0xe0
      13'h1236: dout  = 8'b11111110; // 4662 : 254 - 0xfe
      13'h1237: dout  = 8'b00000000; // 4663 :   0 - 0x0
      13'h1238: dout  = 8'b00000000; // 4664 :   0 - 0x0
      13'h1239: dout  = 8'b00000000; // 4665 :   0 - 0x0
      13'h123A: dout  = 8'b00000000; // 4666 :   0 - 0x0
      13'h123B: dout  = 8'b00000000; // 4667 :   0 - 0x0
      13'h123C: dout  = 8'b00000000; // 4668 :   0 - 0x0
      13'h123D: dout  = 8'b00000000; // 4669 :   0 - 0x0
      13'h123E: dout  = 8'b00000000; // 4670 :   0 - 0x0
      13'h123F: dout  = 8'b00000000; // 4671 :   0 - 0x0
      13'h1240: dout  = 8'b00000000; // 4672 :   0 - 0x0 -- Background 0x24
      13'h1241: dout  = 8'b00000000; // 4673 :   0 - 0x0
      13'h1242: dout  = 8'b00000000; // 4674 :   0 - 0x0
      13'h1243: dout  = 8'b00000000; // 4675 :   0 - 0x0
      13'h1244: dout  = 8'b00000000; // 4676 :   0 - 0x0
      13'h1245: dout  = 8'b00000000; // 4677 :   0 - 0x0
      13'h1246: dout  = 8'b00000000; // 4678 :   0 - 0x0
      13'h1247: dout  = 8'b00000000; // 4679 :   0 - 0x0
      13'h1248: dout  = 8'b00000000; // 4680 :   0 - 0x0
      13'h1249: dout  = 8'b00000000; // 4681 :   0 - 0x0
      13'h124A: dout  = 8'b00000000; // 4682 :   0 - 0x0
      13'h124B: dout  = 8'b00000000; // 4683 :   0 - 0x0
      13'h124C: dout  = 8'b00000000; // 4684 :   0 - 0x0
      13'h124D: dout  = 8'b00000000; // 4685 :   0 - 0x0
      13'h124E: dout  = 8'b00000000; // 4686 :   0 - 0x0
      13'h124F: dout  = 8'b00000000; // 4687 :   0 - 0x0
      13'h1250: dout  = 8'b00000000; // 4688 :   0 - 0x0 -- Background 0x25
      13'h1251: dout  = 8'b00000000; // 4689 :   0 - 0x0
      13'h1252: dout  = 8'b00000110; // 4690 :   6 - 0x6
      13'h1253: dout  = 8'b00001110; // 4691 :  14 - 0xe
      13'h1254: dout  = 8'b00001000; // 4692 :   8 - 0x8
      13'h1255: dout  = 8'b00001000; // 4693 :   8 - 0x8
      13'h1256: dout  = 8'b00001000; // 4694 :   8 - 0x8
      13'h1257: dout  = 8'b00001000; // 4695 :   8 - 0x8
      13'h1258: dout  = 8'b00000000; // 4696 :   0 - 0x0
      13'h1259: dout  = 8'b00000000; // 4697 :   0 - 0x0
      13'h125A: dout  = 8'b00000000; // 4698 :   0 - 0x0
      13'h125B: dout  = 8'b00000000; // 4699 :   0 - 0x0
      13'h125C: dout  = 8'b00000000; // 4700 :   0 - 0x0
      13'h125D: dout  = 8'b00000000; // 4701 :   0 - 0x0
      13'h125E: dout  = 8'b00000000; // 4702 :   0 - 0x0
      13'h125F: dout  = 8'b00000000; // 4703 :   0 - 0x0
      13'h1260: dout  = 8'b00000000; // 4704 :   0 - 0x0 -- Background 0x26
      13'h1261: dout  = 8'b01111000; // 4705 : 120 - 0x78
      13'h1262: dout  = 8'b01100101; // 4706 : 101 - 0x65
      13'h1263: dout  = 8'b01111001; // 4707 : 121 - 0x79
      13'h1264: dout  = 8'b01100101; // 4708 : 101 - 0x65
      13'h1265: dout  = 8'b01100101; // 4709 : 101 - 0x65
      13'h1266: dout  = 8'b01111000; // 4710 : 120 - 0x78
      13'h1267: dout  = 8'b00000000; // 4711 :   0 - 0x0
      13'h1268: dout  = 8'b00000000; // 4712 :   0 - 0x0
      13'h1269: dout  = 8'b00000000; // 4713 :   0 - 0x0
      13'h126A: dout  = 8'b00000000; // 4714 :   0 - 0x0
      13'h126B: dout  = 8'b00000000; // 4715 :   0 - 0x0
      13'h126C: dout  = 8'b00000000; // 4716 :   0 - 0x0
      13'h126D: dout  = 8'b00000000; // 4717 :   0 - 0x0
      13'h126E: dout  = 8'b00000000; // 4718 :   0 - 0x0
      13'h126F: dout  = 8'b00000000; // 4719 :   0 - 0x0
      13'h1270: dout  = 8'b00000000; // 4720 :   0 - 0x0 -- Background 0x27
      13'h1271: dout  = 8'b11100100; // 4721 : 228 - 0xe4
      13'h1272: dout  = 8'b10010110; // 4722 : 150 - 0x96
      13'h1273: dout  = 8'b10010110; // 4723 : 150 - 0x96
      13'h1274: dout  = 8'b10010111; // 4724 : 151 - 0x97
      13'h1275: dout  = 8'b10010110; // 4725 : 150 - 0x96
      13'h1276: dout  = 8'b11100110; // 4726 : 230 - 0xe6
      13'h1277: dout  = 8'b00000000; // 4727 :   0 - 0x0
      13'h1278: dout  = 8'b00000000; // 4728 :   0 - 0x0
      13'h1279: dout  = 8'b00000000; // 4729 :   0 - 0x0
      13'h127A: dout  = 8'b00000000; // 4730 :   0 - 0x0
      13'h127B: dout  = 8'b00000000; // 4731 :   0 - 0x0
      13'h127C: dout  = 8'b00000000; // 4732 :   0 - 0x0
      13'h127D: dout  = 8'b00000000; // 4733 :   0 - 0x0
      13'h127E: dout  = 8'b00000000; // 4734 :   0 - 0x0
      13'h127F: dout  = 8'b00000000; // 4735 :   0 - 0x0
      13'h1280: dout  = 8'b00000000; // 4736 :   0 - 0x0 -- Background 0x28
      13'h1281: dout  = 8'b01011001; // 4737 :  89 - 0x59
      13'h1282: dout  = 8'b01011001; // 4738 :  89 - 0x59
      13'h1283: dout  = 8'b01011001; // 4739 :  89 - 0x59
      13'h1284: dout  = 8'b01011001; // 4740 :  89 - 0x59
      13'h1285: dout  = 8'b11011001; // 4741 : 217 - 0xd9
      13'h1286: dout  = 8'b01001110; // 4742 :  78 - 0x4e
      13'h1287: dout  = 8'b00000000; // 4743 :   0 - 0x0
      13'h1288: dout  = 8'b00000000; // 4744 :   0 - 0x0
      13'h1289: dout  = 8'b00000000; // 4745 :   0 - 0x0
      13'h128A: dout  = 8'b00000000; // 4746 :   0 - 0x0
      13'h128B: dout  = 8'b00000000; // 4747 :   0 - 0x0
      13'h128C: dout  = 8'b00000000; // 4748 :   0 - 0x0
      13'h128D: dout  = 8'b00000000; // 4749 :   0 - 0x0
      13'h128E: dout  = 8'b00000000; // 4750 :   0 - 0x0
      13'h128F: dout  = 8'b00000000; // 4751 :   0 - 0x0
      13'h1290: dout  = 8'b00000000; // 4752 :   0 - 0x0 -- Background 0x29
      13'h1291: dout  = 8'b00111100; // 4753 :  60 - 0x3c
      13'h1292: dout  = 8'b01110000; // 4754 : 112 - 0x70
      13'h1293: dout  = 8'b01110000; // 4755 : 112 - 0x70
      13'h1294: dout  = 8'b00111100; // 4756 :  60 - 0x3c
      13'h1295: dout  = 8'b00001100; // 4757 :  12 - 0xc
      13'h1296: dout  = 8'b01111000; // 4758 : 120 - 0x78
      13'h1297: dout  = 8'b00000000; // 4759 :   0 - 0x0
      13'h1298: dout  = 8'b00000000; // 4760 :   0 - 0x0
      13'h1299: dout  = 8'b00000000; // 4761 :   0 - 0x0
      13'h129A: dout  = 8'b00000000; // 4762 :   0 - 0x0
      13'h129B: dout  = 8'b00000000; // 4763 :   0 - 0x0
      13'h129C: dout  = 8'b00000000; // 4764 :   0 - 0x0
      13'h129D: dout  = 8'b00000000; // 4765 :   0 - 0x0
      13'h129E: dout  = 8'b00000000; // 4766 :   0 - 0x0
      13'h129F: dout  = 8'b00000000; // 4767 :   0 - 0x0
      13'h12A0: dout  = 8'b00000000; // 4768 :   0 - 0x0 -- Background 0x2a
      13'h12A1: dout  = 8'b00000000; // 4769 :   0 - 0x0
      13'h12A2: dout  = 8'b11000110; // 4770 : 198 - 0xc6
      13'h12A3: dout  = 8'b11101110; // 4771 : 238 - 0xee
      13'h12A4: dout  = 8'b00101000; // 4772 :  40 - 0x28
      13'h12A5: dout  = 8'b00101000; // 4773 :  40 - 0x28
      13'h12A6: dout  = 8'b00101000; // 4774 :  40 - 0x28
      13'h12A7: dout  = 8'b00101000; // 4775 :  40 - 0x28
      13'h12A8: dout  = 8'b00000000; // 4776 :   0 - 0x0
      13'h12A9: dout  = 8'b00000000; // 4777 :   0 - 0x0
      13'h12AA: dout  = 8'b00000000; // 4778 :   0 - 0x0
      13'h12AB: dout  = 8'b00000000; // 4779 :   0 - 0x0
      13'h12AC: dout  = 8'b00000000; // 4780 :   0 - 0x0
      13'h12AD: dout  = 8'b00000000; // 4781 :   0 - 0x0
      13'h12AE: dout  = 8'b00000000; // 4782 :   0 - 0x0
      13'h12AF: dout  = 8'b00000000; // 4783 :   0 - 0x0
      13'h12B0: dout  = 8'b00001000; // 4784 :   8 - 0x8 -- Background 0x2b
      13'h12B1: dout  = 8'b00001000; // 4785 :   8 - 0x8
      13'h12B2: dout  = 8'b00001000; // 4786 :   8 - 0x8
      13'h12B3: dout  = 8'b00001000; // 4787 :   8 - 0x8
      13'h12B4: dout  = 8'b00001110; // 4788 :  14 - 0xe
      13'h12B5: dout  = 8'b00000110; // 4789 :   6 - 0x6
      13'h12B6: dout  = 8'b00000000; // 4790 :   0 - 0x0
      13'h12B7: dout  = 8'b00000000; // 4791 :   0 - 0x0
      13'h12B8: dout  = 8'b00000000; // 4792 :   0 - 0x0
      13'h12B9: dout  = 8'b00000000; // 4793 :   0 - 0x0
      13'h12BA: dout  = 8'b00000000; // 4794 :   0 - 0x0
      13'h12BB: dout  = 8'b00000000; // 4795 :   0 - 0x0
      13'h12BC: dout  = 8'b00000000; // 4796 :   0 - 0x0
      13'h12BD: dout  = 8'b00000000; // 4797 :   0 - 0x0
      13'h12BE: dout  = 8'b00000000; // 4798 :   0 - 0x0
      13'h12BF: dout  = 8'b00000000; // 4799 :   0 - 0x0
      13'h12C0: dout  = 8'b00101000; // 4800 :  40 - 0x28 -- Background 0x2c
      13'h12C1: dout  = 8'b00101000; // 4801 :  40 - 0x28
      13'h12C2: dout  = 8'b00101000; // 4802 :  40 - 0x28
      13'h12C3: dout  = 8'b00101000; // 4803 :  40 - 0x28
      13'h12C4: dout  = 8'b11101110; // 4804 : 238 - 0xee
      13'h12C5: dout  = 8'b11000110; // 4805 : 198 - 0xc6
      13'h12C6: dout  = 8'b00000000; // 4806 :   0 - 0x0
      13'h12C7: dout  = 8'b00000000; // 4807 :   0 - 0x0
      13'h12C8: dout  = 8'b00000000; // 4808 :   0 - 0x0
      13'h12C9: dout  = 8'b00000000; // 4809 :   0 - 0x0
      13'h12CA: dout  = 8'b00000000; // 4810 :   0 - 0x0
      13'h12CB: dout  = 8'b00000000; // 4811 :   0 - 0x0
      13'h12CC: dout  = 8'b00000000; // 4812 :   0 - 0x0
      13'h12CD: dout  = 8'b00000000; // 4813 :   0 - 0x0
      13'h12CE: dout  = 8'b00000000; // 4814 :   0 - 0x0
      13'h12CF: dout  = 8'b00000000; // 4815 :   0 - 0x0
      13'h12D0: dout  = 8'b00000000; // 4816 :   0 - 0x0 -- Background 0x2d
      13'h12D1: dout  = 8'b00000000; // 4817 :   0 - 0x0
      13'h12D2: dout  = 8'b01100000; // 4818 :  96 - 0x60
      13'h12D3: dout  = 8'b01110000; // 4819 : 112 - 0x70
      13'h12D4: dout  = 8'b00010000; // 4820 :  16 - 0x10
      13'h12D5: dout  = 8'b00010000; // 4821 :  16 - 0x10
      13'h12D6: dout  = 8'b00010000; // 4822 :  16 - 0x10
      13'h12D7: dout  = 8'b00010000; // 4823 :  16 - 0x10
      13'h12D8: dout  = 8'b00000000; // 4824 :   0 - 0x0
      13'h12D9: dout  = 8'b00000000; // 4825 :   0 - 0x0
      13'h12DA: dout  = 8'b00000000; // 4826 :   0 - 0x0
      13'h12DB: dout  = 8'b00000000; // 4827 :   0 - 0x0
      13'h12DC: dout  = 8'b00000000; // 4828 :   0 - 0x0
      13'h12DD: dout  = 8'b00000000; // 4829 :   0 - 0x0
      13'h12DE: dout  = 8'b00000000; // 4830 :   0 - 0x0
      13'h12DF: dout  = 8'b00000000; // 4831 :   0 - 0x0
      13'h12E0: dout  = 8'b00011100; // 4832 :  28 - 0x1c -- Background 0x2e
      13'h12E1: dout  = 8'b00111110; // 4833 :  62 - 0x3e
      13'h12E2: dout  = 8'b00111100; // 4834 :  60 - 0x3c
      13'h12E3: dout  = 8'b00111000; // 4835 :  56 - 0x38
      13'h12E4: dout  = 8'b00110000; // 4836 :  48 - 0x30
      13'h12E5: dout  = 8'b00000000; // 4837 :   0 - 0x0
      13'h12E6: dout  = 8'b01100000; // 4838 :  96 - 0x60
      13'h12E7: dout  = 8'b00000000; // 4839 :   0 - 0x0
      13'h12E8: dout  = 8'b00000000; // 4840 :   0 - 0x0
      13'h12E9: dout  = 8'b00000000; // 4841 :   0 - 0x0
      13'h12EA: dout  = 8'b00000000; // 4842 :   0 - 0x0
      13'h12EB: dout  = 8'b00000000; // 4843 :   0 - 0x0
      13'h12EC: dout  = 8'b00000000; // 4844 :   0 - 0x0
      13'h12ED: dout  = 8'b00000000; // 4845 :   0 - 0x0
      13'h12EE: dout  = 8'b00000000; // 4846 :   0 - 0x0
      13'h12EF: dout  = 8'b00000000; // 4847 :   0 - 0x0
      13'h12F0: dout  = 8'b00010000; // 4848 :  16 - 0x10 -- Background 0x2f
      13'h12F1: dout  = 8'b00010000; // 4849 :  16 - 0x10
      13'h12F2: dout  = 8'b00010000; // 4850 :  16 - 0x10
      13'h12F3: dout  = 8'b00010000; // 4851 :  16 - 0x10
      13'h12F4: dout  = 8'b01110000; // 4852 : 112 - 0x70
      13'h12F5: dout  = 8'b01100000; // 4853 :  96 - 0x60
      13'h12F6: dout  = 8'b00000000; // 4854 :   0 - 0x0
      13'h12F7: dout  = 8'b00000000; // 4855 :   0 - 0x0
      13'h12F8: dout  = 8'b00000000; // 4856 :   0 - 0x0
      13'h12F9: dout  = 8'b00000000; // 4857 :   0 - 0x0
      13'h12FA: dout  = 8'b00000000; // 4858 :   0 - 0x0
      13'h12FB: dout  = 8'b00000000; // 4859 :   0 - 0x0
      13'h12FC: dout  = 8'b00000000; // 4860 :   0 - 0x0
      13'h12FD: dout  = 8'b00000000; // 4861 :   0 - 0x0
      13'h12FE: dout  = 8'b00000000; // 4862 :   0 - 0x0
      13'h12FF: dout  = 8'b00000000; // 4863 :   0 - 0x0
      13'h1300: dout  = 8'b11111111; // 4864 : 255 - 0xff -- Background 0x30
      13'h1301: dout  = 8'b11111111; // 4865 : 255 - 0xff
      13'h1302: dout  = 8'b00111000; // 4866 :  56 - 0x38
      13'h1303: dout  = 8'b01101100; // 4867 : 108 - 0x6c
      13'h1304: dout  = 8'b11000110; // 4868 : 198 - 0xc6
      13'h1305: dout  = 8'b10000011; // 4869 : 131 - 0x83
      13'h1306: dout  = 8'b11111111; // 4870 : 255 - 0xff
      13'h1307: dout  = 8'b11111111; // 4871 : 255 - 0xff
      13'h1308: dout  = 8'b00000000; // 4872 :   0 - 0x0
      13'h1309: dout  = 8'b00000000; // 4873 :   0 - 0x0
      13'h130A: dout  = 8'b00000000; // 4874 :   0 - 0x0
      13'h130B: dout  = 8'b00000000; // 4875 :   0 - 0x0
      13'h130C: dout  = 8'b00000000; // 4876 :   0 - 0x0
      13'h130D: dout  = 8'b00000000; // 4877 :   0 - 0x0
      13'h130E: dout  = 8'b00000000; // 4878 :   0 - 0x0
      13'h130F: dout  = 8'b00000000; // 4879 :   0 - 0x0
      13'h1310: dout  = 8'b11111111; // 4880 : 255 - 0xff -- Background 0x31
      13'h1311: dout  = 8'b00111000; // 4881 :  56 - 0x38
      13'h1312: dout  = 8'b01101100; // 4882 : 108 - 0x6c
      13'h1313: dout  = 8'b11000110; // 4883 : 198 - 0xc6
      13'h1314: dout  = 8'b10000011; // 4884 : 131 - 0x83
      13'h1315: dout  = 8'b11111111; // 4885 : 255 - 0xff
      13'h1316: dout  = 8'b11111111; // 4886 : 255 - 0xff
      13'h1317: dout  = 8'b00000000; // 4887 :   0 - 0x0
      13'h1318: dout  = 8'b00000000; // 4888 :   0 - 0x0
      13'h1319: dout  = 8'b00000000; // 4889 :   0 - 0x0
      13'h131A: dout  = 8'b00000000; // 4890 :   0 - 0x0
      13'h131B: dout  = 8'b00000000; // 4891 :   0 - 0x0
      13'h131C: dout  = 8'b00000000; // 4892 :   0 - 0x0
      13'h131D: dout  = 8'b00000000; // 4893 :   0 - 0x0
      13'h131E: dout  = 8'b00000000; // 4894 :   0 - 0x0
      13'h131F: dout  = 8'b00000000; // 4895 :   0 - 0x0
      13'h1320: dout  = 8'b00111000; // 4896 :  56 - 0x38 -- Background 0x32
      13'h1321: dout  = 8'b01101100; // 4897 : 108 - 0x6c
      13'h1322: dout  = 8'b11000110; // 4898 : 198 - 0xc6
      13'h1323: dout  = 8'b10000011; // 4899 : 131 - 0x83
      13'h1324: dout  = 8'b11111111; // 4900 : 255 - 0xff
      13'h1325: dout  = 8'b11111111; // 4901 : 255 - 0xff
      13'h1326: dout  = 8'b00000000; // 4902 :   0 - 0x0
      13'h1327: dout  = 8'b00000000; // 4903 :   0 - 0x0
      13'h1328: dout  = 8'b00000000; // 4904 :   0 - 0x0
      13'h1329: dout  = 8'b00000000; // 4905 :   0 - 0x0
      13'h132A: dout  = 8'b00000000; // 4906 :   0 - 0x0
      13'h132B: dout  = 8'b00000000; // 4907 :   0 - 0x0
      13'h132C: dout  = 8'b00000000; // 4908 :   0 - 0x0
      13'h132D: dout  = 8'b00000000; // 4909 :   0 - 0x0
      13'h132E: dout  = 8'b00000000; // 4910 :   0 - 0x0
      13'h132F: dout  = 8'b00000000; // 4911 :   0 - 0x0
      13'h1330: dout  = 8'b01101100; // 4912 : 108 - 0x6c -- Background 0x33
      13'h1331: dout  = 8'b11000110; // 4913 : 198 - 0xc6
      13'h1332: dout  = 8'b10000011; // 4914 : 131 - 0x83
      13'h1333: dout  = 8'b11111111; // 4915 : 255 - 0xff
      13'h1334: dout  = 8'b11111111; // 4916 : 255 - 0xff
      13'h1335: dout  = 8'b00000000; // 4917 :   0 - 0x0
      13'h1336: dout  = 8'b00000000; // 4918 :   0 - 0x0
      13'h1337: dout  = 8'b00000000; // 4919 :   0 - 0x0
      13'h1338: dout  = 8'b00000000; // 4920 :   0 - 0x0
      13'h1339: dout  = 8'b00000000; // 4921 :   0 - 0x0
      13'h133A: dout  = 8'b00000000; // 4922 :   0 - 0x0
      13'h133B: dout  = 8'b00000000; // 4923 :   0 - 0x0
      13'h133C: dout  = 8'b00000000; // 4924 :   0 - 0x0
      13'h133D: dout  = 8'b00000000; // 4925 :   0 - 0x0
      13'h133E: dout  = 8'b00000000; // 4926 :   0 - 0x0
      13'h133F: dout  = 8'b00000000; // 4927 :   0 - 0x0
      13'h1340: dout  = 8'b11000110; // 4928 : 198 - 0xc6 -- Background 0x34
      13'h1341: dout  = 8'b10000011; // 4929 : 131 - 0x83
      13'h1342: dout  = 8'b11111111; // 4930 : 255 - 0xff
      13'h1343: dout  = 8'b11111111; // 4931 : 255 - 0xff
      13'h1344: dout  = 8'b00000000; // 4932 :   0 - 0x0
      13'h1345: dout  = 8'b00000000; // 4933 :   0 - 0x0
      13'h1346: dout  = 8'b00000000; // 4934 :   0 - 0x0
      13'h1347: dout  = 8'b00000000; // 4935 :   0 - 0x0
      13'h1348: dout  = 8'b00000000; // 4936 :   0 - 0x0
      13'h1349: dout  = 8'b00000000; // 4937 :   0 - 0x0
      13'h134A: dout  = 8'b00000000; // 4938 :   0 - 0x0
      13'h134B: dout  = 8'b00000000; // 4939 :   0 - 0x0
      13'h134C: dout  = 8'b00000000; // 4940 :   0 - 0x0
      13'h134D: dout  = 8'b00000000; // 4941 :   0 - 0x0
      13'h134E: dout  = 8'b00000000; // 4942 :   0 - 0x0
      13'h134F: dout  = 8'b00000000; // 4943 :   0 - 0x0
      13'h1350: dout  = 8'b10000011; // 4944 : 131 - 0x83 -- Background 0x35
      13'h1351: dout  = 8'b11111111; // 4945 : 255 - 0xff
      13'h1352: dout  = 8'b11111111; // 4946 : 255 - 0xff
      13'h1353: dout  = 8'b00000000; // 4947 :   0 - 0x0
      13'h1354: dout  = 8'b00000000; // 4948 :   0 - 0x0
      13'h1355: dout  = 8'b00000000; // 4949 :   0 - 0x0
      13'h1356: dout  = 8'b00000000; // 4950 :   0 - 0x0
      13'h1357: dout  = 8'b00000000; // 4951 :   0 - 0x0
      13'h1358: dout  = 8'b00000000; // 4952 :   0 - 0x0
      13'h1359: dout  = 8'b00000000; // 4953 :   0 - 0x0
      13'h135A: dout  = 8'b00000000; // 4954 :   0 - 0x0
      13'h135B: dout  = 8'b00000000; // 4955 :   0 - 0x0
      13'h135C: dout  = 8'b00000000; // 4956 :   0 - 0x0
      13'h135D: dout  = 8'b00000000; // 4957 :   0 - 0x0
      13'h135E: dout  = 8'b00000000; // 4958 :   0 - 0x0
      13'h135F: dout  = 8'b00000000; // 4959 :   0 - 0x0
      13'h1360: dout  = 8'b11111111; // 4960 : 255 - 0xff -- Background 0x36
      13'h1361: dout  = 8'b11111111; // 4961 : 255 - 0xff
      13'h1362: dout  = 8'b00000000; // 4962 :   0 - 0x0
      13'h1363: dout  = 8'b00000000; // 4963 :   0 - 0x0
      13'h1364: dout  = 8'b00000000; // 4964 :   0 - 0x0
      13'h1365: dout  = 8'b00000000; // 4965 :   0 - 0x0
      13'h1366: dout  = 8'b00000000; // 4966 :   0 - 0x0
      13'h1367: dout  = 8'b00000000; // 4967 :   0 - 0x0
      13'h1368: dout  = 8'b00000000; // 4968 :   0 - 0x0
      13'h1369: dout  = 8'b00000000; // 4969 :   0 - 0x0
      13'h136A: dout  = 8'b00000000; // 4970 :   0 - 0x0
      13'h136B: dout  = 8'b00000000; // 4971 :   0 - 0x0
      13'h136C: dout  = 8'b00000000; // 4972 :   0 - 0x0
      13'h136D: dout  = 8'b00000000; // 4973 :   0 - 0x0
      13'h136E: dout  = 8'b00000000; // 4974 :   0 - 0x0
      13'h136F: dout  = 8'b00000000; // 4975 :   0 - 0x0
      13'h1370: dout  = 8'b11111111; // 4976 : 255 - 0xff -- Background 0x37
      13'h1371: dout  = 8'b00000000; // 4977 :   0 - 0x0
      13'h1372: dout  = 8'b00000000; // 4978 :   0 - 0x0
      13'h1373: dout  = 8'b00000000; // 4979 :   0 - 0x0
      13'h1374: dout  = 8'b00000000; // 4980 :   0 - 0x0
      13'h1375: dout  = 8'b00000000; // 4981 :   0 - 0x0
      13'h1376: dout  = 8'b00000000; // 4982 :   0 - 0x0
      13'h1377: dout  = 8'b00000000; // 4983 :   0 - 0x0
      13'h1378: dout  = 8'b00000000; // 4984 :   0 - 0x0
      13'h1379: dout  = 8'b00000000; // 4985 :   0 - 0x0
      13'h137A: dout  = 8'b00000000; // 4986 :   0 - 0x0
      13'h137B: dout  = 8'b00000000; // 4987 :   0 - 0x0
      13'h137C: dout  = 8'b00000000; // 4988 :   0 - 0x0
      13'h137D: dout  = 8'b00000000; // 4989 :   0 - 0x0
      13'h137E: dout  = 8'b00000000; // 4990 :   0 - 0x0
      13'h137F: dout  = 8'b00000000; // 4991 :   0 - 0x0
      13'h1380: dout  = 8'b00000000; // 4992 :   0 - 0x0 -- Background 0x38
      13'h1381: dout  = 8'b00000000; // 4993 :   0 - 0x0
      13'h1382: dout  = 8'b00000000; // 4994 :   0 - 0x0
      13'h1383: dout  = 8'b00000000; // 4995 :   0 - 0x0
      13'h1384: dout  = 8'b00000000; // 4996 :   0 - 0x0
      13'h1385: dout  = 8'b00000000; // 4997 :   0 - 0x0
      13'h1386: dout  = 8'b00000000; // 4998 :   0 - 0x0
      13'h1387: dout  = 8'b11111111; // 4999 : 255 - 0xff
      13'h1388: dout  = 8'b00000000; // 5000 :   0 - 0x0
      13'h1389: dout  = 8'b00000000; // 5001 :   0 - 0x0
      13'h138A: dout  = 8'b00000000; // 5002 :   0 - 0x0
      13'h138B: dout  = 8'b00000000; // 5003 :   0 - 0x0
      13'h138C: dout  = 8'b00000000; // 5004 :   0 - 0x0
      13'h138D: dout  = 8'b00000000; // 5005 :   0 - 0x0
      13'h138E: dout  = 8'b00000000; // 5006 :   0 - 0x0
      13'h138F: dout  = 8'b00000000; // 5007 :   0 - 0x0
      13'h1390: dout  = 8'b00000000; // 5008 :   0 - 0x0 -- Background 0x39
      13'h1391: dout  = 8'b00000000; // 5009 :   0 - 0x0
      13'h1392: dout  = 8'b00000000; // 5010 :   0 - 0x0
      13'h1393: dout  = 8'b00000000; // 5011 :   0 - 0x0
      13'h1394: dout  = 8'b00000000; // 5012 :   0 - 0x0
      13'h1395: dout  = 8'b00000000; // 5013 :   0 - 0x0
      13'h1396: dout  = 8'b11111111; // 5014 : 255 - 0xff
      13'h1397: dout  = 8'b11111111; // 5015 : 255 - 0xff
      13'h1398: dout  = 8'b00000000; // 5016 :   0 - 0x0
      13'h1399: dout  = 8'b00000000; // 5017 :   0 - 0x0
      13'h139A: dout  = 8'b00000000; // 5018 :   0 - 0x0
      13'h139B: dout  = 8'b00000000; // 5019 :   0 - 0x0
      13'h139C: dout  = 8'b00000000; // 5020 :   0 - 0x0
      13'h139D: dout  = 8'b00000000; // 5021 :   0 - 0x0
      13'h139E: dout  = 8'b00000000; // 5022 :   0 - 0x0
      13'h139F: dout  = 8'b00000000; // 5023 :   0 - 0x0
      13'h13A0: dout  = 8'b00000000; // 5024 :   0 - 0x0 -- Background 0x3a
      13'h13A1: dout  = 8'b00000000; // 5025 :   0 - 0x0
      13'h13A2: dout  = 8'b00000000; // 5026 :   0 - 0x0
      13'h13A3: dout  = 8'b00000000; // 5027 :   0 - 0x0
      13'h13A4: dout  = 8'b00000000; // 5028 :   0 - 0x0
      13'h13A5: dout  = 8'b11111111; // 5029 : 255 - 0xff
      13'h13A6: dout  = 8'b11111111; // 5030 : 255 - 0xff
      13'h13A7: dout  = 8'b00111000; // 5031 :  56 - 0x38
      13'h13A8: dout  = 8'b00000000; // 5032 :   0 - 0x0
      13'h13A9: dout  = 8'b00000000; // 5033 :   0 - 0x0
      13'h13AA: dout  = 8'b00000000; // 5034 :   0 - 0x0
      13'h13AB: dout  = 8'b00000000; // 5035 :   0 - 0x0
      13'h13AC: dout  = 8'b00000000; // 5036 :   0 - 0x0
      13'h13AD: dout  = 8'b00000000; // 5037 :   0 - 0x0
      13'h13AE: dout  = 8'b00000000; // 5038 :   0 - 0x0
      13'h13AF: dout  = 8'b00000000; // 5039 :   0 - 0x0
      13'h13B0: dout  = 8'b00000000; // 5040 :   0 - 0x0 -- Background 0x3b
      13'h13B1: dout  = 8'b00000000; // 5041 :   0 - 0x0
      13'h13B2: dout  = 8'b00000000; // 5042 :   0 - 0x0
      13'h13B3: dout  = 8'b00000000; // 5043 :   0 - 0x0
      13'h13B4: dout  = 8'b11111111; // 5044 : 255 - 0xff
      13'h13B5: dout  = 8'b11111111; // 5045 : 255 - 0xff
      13'h13B6: dout  = 8'b00111000; // 5046 :  56 - 0x38
      13'h13B7: dout  = 8'b01101100; // 5047 : 108 - 0x6c
      13'h13B8: dout  = 8'b00000000; // 5048 :   0 - 0x0
      13'h13B9: dout  = 8'b00000000; // 5049 :   0 - 0x0
      13'h13BA: dout  = 8'b00000000; // 5050 :   0 - 0x0
      13'h13BB: dout  = 8'b00000000; // 5051 :   0 - 0x0
      13'h13BC: dout  = 8'b00000000; // 5052 :   0 - 0x0
      13'h13BD: dout  = 8'b00000000; // 5053 :   0 - 0x0
      13'h13BE: dout  = 8'b00000000; // 5054 :   0 - 0x0
      13'h13BF: dout  = 8'b00000000; // 5055 :   0 - 0x0
      13'h13C0: dout  = 8'b00000000; // 5056 :   0 - 0x0 -- Background 0x3c
      13'h13C1: dout  = 8'b00000000; // 5057 :   0 - 0x0
      13'h13C2: dout  = 8'b00000000; // 5058 :   0 - 0x0
      13'h13C3: dout  = 8'b11111111; // 5059 : 255 - 0xff
      13'h13C4: dout  = 8'b11111111; // 5060 : 255 - 0xff
      13'h13C5: dout  = 8'b00111000; // 5061 :  56 - 0x38
      13'h13C6: dout  = 8'b01101100; // 5062 : 108 - 0x6c
      13'h13C7: dout  = 8'b11000110; // 5063 : 198 - 0xc6
      13'h13C8: dout  = 8'b00000000; // 5064 :   0 - 0x0
      13'h13C9: dout  = 8'b00000000; // 5065 :   0 - 0x0
      13'h13CA: dout  = 8'b00000000; // 5066 :   0 - 0x0
      13'h13CB: dout  = 8'b00000000; // 5067 :   0 - 0x0
      13'h13CC: dout  = 8'b00000000; // 5068 :   0 - 0x0
      13'h13CD: dout  = 8'b00000000; // 5069 :   0 - 0x0
      13'h13CE: dout  = 8'b00000000; // 5070 :   0 - 0x0
      13'h13CF: dout  = 8'b00000000; // 5071 :   0 - 0x0
      13'h13D0: dout  = 8'b00000000; // 5072 :   0 - 0x0 -- Background 0x3d
      13'h13D1: dout  = 8'b00000000; // 5073 :   0 - 0x0
      13'h13D2: dout  = 8'b11111111; // 5074 : 255 - 0xff
      13'h13D3: dout  = 8'b11111111; // 5075 : 255 - 0xff
      13'h13D4: dout  = 8'b00111000; // 5076 :  56 - 0x38
      13'h13D5: dout  = 8'b01101100; // 5077 : 108 - 0x6c
      13'h13D6: dout  = 8'b11000110; // 5078 : 198 - 0xc6
      13'h13D7: dout  = 8'b10000011; // 5079 : 131 - 0x83
      13'h13D8: dout  = 8'b00000000; // 5080 :   0 - 0x0
      13'h13D9: dout  = 8'b00000000; // 5081 :   0 - 0x0
      13'h13DA: dout  = 8'b00000000; // 5082 :   0 - 0x0
      13'h13DB: dout  = 8'b00000000; // 5083 :   0 - 0x0
      13'h13DC: dout  = 8'b00000000; // 5084 :   0 - 0x0
      13'h13DD: dout  = 8'b00000000; // 5085 :   0 - 0x0
      13'h13DE: dout  = 8'b00000000; // 5086 :   0 - 0x0
      13'h13DF: dout  = 8'b00000000; // 5087 :   0 - 0x0
      13'h13E0: dout  = 8'b00000000; // 5088 :   0 - 0x0 -- Background 0x3e
      13'h13E1: dout  = 8'b11111111; // 5089 : 255 - 0xff
      13'h13E2: dout  = 8'b11111111; // 5090 : 255 - 0xff
      13'h13E3: dout  = 8'b00111000; // 5091 :  56 - 0x38
      13'h13E4: dout  = 8'b01101100; // 5092 : 108 - 0x6c
      13'h13E5: dout  = 8'b11000110; // 5093 : 198 - 0xc6
      13'h13E6: dout  = 8'b10000011; // 5094 : 131 - 0x83
      13'h13E7: dout  = 8'b11111111; // 5095 : 255 - 0xff
      13'h13E8: dout  = 8'b00000000; // 5096 :   0 - 0x0
      13'h13E9: dout  = 8'b00000000; // 5097 :   0 - 0x0
      13'h13EA: dout  = 8'b00000000; // 5098 :   0 - 0x0
      13'h13EB: dout  = 8'b00000000; // 5099 :   0 - 0x0
      13'h13EC: dout  = 8'b00000000; // 5100 :   0 - 0x0
      13'h13ED: dout  = 8'b00000000; // 5101 :   0 - 0x0
      13'h13EE: dout  = 8'b00000000; // 5102 :   0 - 0x0
      13'h13EF: dout  = 8'b00000000; // 5103 :   0 - 0x0
      13'h13F0: dout  = 8'b00000000; // 5104 :   0 - 0x0 -- Background 0x3f
      13'h13F1: dout  = 8'b00000000; // 5105 :   0 - 0x0
      13'h13F2: dout  = 8'b00000000; // 5106 :   0 - 0x0
      13'h13F3: dout  = 8'b00000000; // 5107 :   0 - 0x0
      13'h13F4: dout  = 8'b00000000; // 5108 :   0 - 0x0
      13'h13F5: dout  = 8'b00000000; // 5109 :   0 - 0x0
      13'h13F6: dout  = 8'b00000000; // 5110 :   0 - 0x0
      13'h13F7: dout  = 8'b00000000; // 5111 :   0 - 0x0
      13'h13F8: dout  = 8'b10000001; // 5112 : 129 - 0x81
      13'h13F9: dout  = 8'b11111111; // 5113 : 255 - 0xff
      13'h13FA: dout  = 8'b10000001; // 5114 : 129 - 0x81
      13'h13FB: dout  = 8'b10000001; // 5115 : 129 - 0x81
      13'h13FC: dout  = 8'b10000001; // 5116 : 129 - 0x81
      13'h13FD: dout  = 8'b11111111; // 5117 : 255 - 0xff
      13'h13FE: dout  = 8'b10000001; // 5118 : 129 - 0x81
      13'h13FF: dout  = 8'b10000001; // 5119 : 129 - 0x81
      13'h1400: dout  = 8'b00000000; // 5120 :   0 - 0x0 -- Background 0x40
      13'h1401: dout  = 8'b00000000; // 5121 :   0 - 0x0
      13'h1402: dout  = 8'b00000000; // 5122 :   0 - 0x0
      13'h1403: dout  = 8'b00000000; // 5123 :   0 - 0x0
      13'h1404: dout  = 8'b00000000; // 5124 :   0 - 0x0
      13'h1405: dout  = 8'b00000000; // 5125 :   0 - 0x0
      13'h1406: dout  = 8'b00000000; // 5126 :   0 - 0x0
      13'h1407: dout  = 8'b11111111; // 5127 : 255 - 0xff
      13'h1408: dout  = 8'b10000001; // 5128 : 129 - 0x81
      13'h1409: dout  = 8'b11111111; // 5129 : 255 - 0xff
      13'h140A: dout  = 8'b10000001; // 5130 : 129 - 0x81
      13'h140B: dout  = 8'b10000001; // 5131 : 129 - 0x81
      13'h140C: dout  = 8'b10000001; // 5132 : 129 - 0x81
      13'h140D: dout  = 8'b11111111; // 5133 : 255 - 0xff
      13'h140E: dout  = 8'b10000001; // 5134 : 129 - 0x81
      13'h140F: dout  = 8'b00000000; // 5135 :   0 - 0x0
      13'h1410: dout  = 8'b00000000; // 5136 :   0 - 0x0 -- Background 0x41
      13'h1411: dout  = 8'b00000000; // 5137 :   0 - 0x0
      13'h1412: dout  = 8'b00000000; // 5138 :   0 - 0x0
      13'h1413: dout  = 8'b00000000; // 5139 :   0 - 0x0
      13'h1414: dout  = 8'b00000000; // 5140 :   0 - 0x0
      13'h1415: dout  = 8'b11111111; // 5141 : 255 - 0xff
      13'h1416: dout  = 8'b11111111; // 5142 : 255 - 0xff
      13'h1417: dout  = 8'b00111000; // 5143 :  56 - 0x38
      13'h1418: dout  = 8'b10000001; // 5144 : 129 - 0x81
      13'h1419: dout  = 8'b11111111; // 5145 : 255 - 0xff
      13'h141A: dout  = 8'b10000001; // 5146 : 129 - 0x81
      13'h141B: dout  = 8'b10000001; // 5147 : 129 - 0x81
      13'h141C: dout  = 8'b10000001; // 5148 : 129 - 0x81
      13'h141D: dout  = 8'b00000000; // 5149 :   0 - 0x0
      13'h141E: dout  = 8'b00000000; // 5150 :   0 - 0x0
      13'h141F: dout  = 8'b00000000; // 5151 :   0 - 0x0
      13'h1420: dout  = 8'b00000000; // 5152 :   0 - 0x0 -- Background 0x42
      13'h1421: dout  = 8'b00000000; // 5153 :   0 - 0x0
      13'h1422: dout  = 8'b00000000; // 5154 :   0 - 0x0
      13'h1423: dout  = 8'b00000000; // 5155 :   0 - 0x0
      13'h1424: dout  = 8'b11111111; // 5156 : 255 - 0xff
      13'h1425: dout  = 8'b11111111; // 5157 : 255 - 0xff
      13'h1426: dout  = 8'b00111000; // 5158 :  56 - 0x38
      13'h1427: dout  = 8'b01101100; // 5159 : 108 - 0x6c
      13'h1428: dout  = 8'b10000001; // 5160 : 129 - 0x81
      13'h1429: dout  = 8'b11111111; // 5161 : 255 - 0xff
      13'h142A: dout  = 8'b10000001; // 5162 : 129 - 0x81
      13'h142B: dout  = 8'b10000001; // 5163 : 129 - 0x81
      13'h142C: dout  = 8'b00000000; // 5164 :   0 - 0x0
      13'h142D: dout  = 8'b00000000; // 5165 :   0 - 0x0
      13'h142E: dout  = 8'b00000000; // 5166 :   0 - 0x0
      13'h142F: dout  = 8'b00000000; // 5167 :   0 - 0x0
      13'h1430: dout  = 8'b00000000; // 5168 :   0 - 0x0 -- Background 0x43
      13'h1431: dout  = 8'b00000000; // 5169 :   0 - 0x0
      13'h1432: dout  = 8'b00000000; // 5170 :   0 - 0x0
      13'h1433: dout  = 8'b11111111; // 5171 : 255 - 0xff
      13'h1434: dout  = 8'b11111111; // 5172 : 255 - 0xff
      13'h1435: dout  = 8'b00111000; // 5173 :  56 - 0x38
      13'h1436: dout  = 8'b01101100; // 5174 : 108 - 0x6c
      13'h1437: dout  = 8'b11000110; // 5175 : 198 - 0xc6
      13'h1438: dout  = 8'b10000001; // 5176 : 129 - 0x81
      13'h1439: dout  = 8'b11111111; // 5177 : 255 - 0xff
      13'h143A: dout  = 8'b10000001; // 5178 : 129 - 0x81
      13'h143B: dout  = 8'b00000000; // 5179 :   0 - 0x0
      13'h143C: dout  = 8'b00000000; // 5180 :   0 - 0x0
      13'h143D: dout  = 8'b00000000; // 5181 :   0 - 0x0
      13'h143E: dout  = 8'b00000000; // 5182 :   0 - 0x0
      13'h143F: dout  = 8'b00000000; // 5183 :   0 - 0x0
      13'h1440: dout  = 8'b00000000; // 5184 :   0 - 0x0 -- Background 0x44
      13'h1441: dout  = 8'b00000000; // 5185 :   0 - 0x0
      13'h1442: dout  = 8'b11111111; // 5186 : 255 - 0xff
      13'h1443: dout  = 8'b11111111; // 5187 : 255 - 0xff
      13'h1444: dout  = 8'b00111000; // 5188 :  56 - 0x38
      13'h1445: dout  = 8'b01101100; // 5189 : 108 - 0x6c
      13'h1446: dout  = 8'b11000110; // 5190 : 198 - 0xc6
      13'h1447: dout  = 8'b10000011; // 5191 : 131 - 0x83
      13'h1448: dout  = 8'b10000001; // 5192 : 129 - 0x81
      13'h1449: dout  = 8'b11111111; // 5193 : 255 - 0xff
      13'h144A: dout  = 8'b00000000; // 5194 :   0 - 0x0
      13'h144B: dout  = 8'b00000000; // 5195 :   0 - 0x0
      13'h144C: dout  = 8'b00000000; // 5196 :   0 - 0x0
      13'h144D: dout  = 8'b00000000; // 5197 :   0 - 0x0
      13'h144E: dout  = 8'b00000000; // 5198 :   0 - 0x0
      13'h144F: dout  = 8'b00000000; // 5199 :   0 - 0x0
      13'h1450: dout  = 8'b00000000; // 5200 :   0 - 0x0 -- Background 0x45
      13'h1451: dout  = 8'b11111111; // 5201 : 255 - 0xff
      13'h1452: dout  = 8'b11111111; // 5202 : 255 - 0xff
      13'h1453: dout  = 8'b00111000; // 5203 :  56 - 0x38
      13'h1454: dout  = 8'b01101100; // 5204 : 108 - 0x6c
      13'h1455: dout  = 8'b11000110; // 5205 : 198 - 0xc6
      13'h1456: dout  = 8'b10000011; // 5206 : 131 - 0x83
      13'h1457: dout  = 8'b11111111; // 5207 : 255 - 0xff
      13'h1458: dout  = 8'b10000001; // 5208 : 129 - 0x81
      13'h1459: dout  = 8'b00000000; // 5209 :   0 - 0x0
      13'h145A: dout  = 8'b00000000; // 5210 :   0 - 0x0
      13'h145B: dout  = 8'b00000000; // 5211 :   0 - 0x0
      13'h145C: dout  = 8'b00000000; // 5212 :   0 - 0x0
      13'h145D: dout  = 8'b00000000; // 5213 :   0 - 0x0
      13'h145E: dout  = 8'b00000000; // 5214 :   0 - 0x0
      13'h145F: dout  = 8'b00000000; // 5215 :   0 - 0x0
      13'h1460: dout  = 8'b11111111; // 5216 : 255 - 0xff -- Background 0x46
      13'h1461: dout  = 8'b00111000; // 5217 :  56 - 0x38
      13'h1462: dout  = 8'b01101100; // 5218 : 108 - 0x6c
      13'h1463: dout  = 8'b11000110; // 5219 : 198 - 0xc6
      13'h1464: dout  = 8'b10000011; // 5220 : 131 - 0x83
      13'h1465: dout  = 8'b11111111; // 5221 : 255 - 0xff
      13'h1466: dout  = 8'b11111111; // 5222 : 255 - 0xff
      13'h1467: dout  = 8'b00000000; // 5223 :   0 - 0x0
      13'h1468: dout  = 8'b00000000; // 5224 :   0 - 0x0
      13'h1469: dout  = 8'b00000000; // 5225 :   0 - 0x0
      13'h146A: dout  = 8'b00000000; // 5226 :   0 - 0x0
      13'h146B: dout  = 8'b00000000; // 5227 :   0 - 0x0
      13'h146C: dout  = 8'b00000000; // 5228 :   0 - 0x0
      13'h146D: dout  = 8'b00000000; // 5229 :   0 - 0x0
      13'h146E: dout  = 8'b00000000; // 5230 :   0 - 0x0
      13'h146F: dout  = 8'b10000001; // 5231 : 129 - 0x81
      13'h1470: dout  = 8'b00111000; // 5232 :  56 - 0x38 -- Background 0x47
      13'h1471: dout  = 8'b01101100; // 5233 : 108 - 0x6c
      13'h1472: dout  = 8'b11000110; // 5234 : 198 - 0xc6
      13'h1473: dout  = 8'b10000011; // 5235 : 131 - 0x83
      13'h1474: dout  = 8'b11111111; // 5236 : 255 - 0xff
      13'h1475: dout  = 8'b11111111; // 5237 : 255 - 0xff
      13'h1476: dout  = 8'b00000000; // 5238 :   0 - 0x0
      13'h1477: dout  = 8'b00000000; // 5239 :   0 - 0x0
      13'h1478: dout  = 8'b00000000; // 5240 :   0 - 0x0
      13'h1479: dout  = 8'b00000000; // 5241 :   0 - 0x0
      13'h147A: dout  = 8'b00000000; // 5242 :   0 - 0x0
      13'h147B: dout  = 8'b00000000; // 5243 :   0 - 0x0
      13'h147C: dout  = 8'b00000000; // 5244 :   0 - 0x0
      13'h147D: dout  = 8'b00000000; // 5245 :   0 - 0x0
      13'h147E: dout  = 8'b10000001; // 5246 : 129 - 0x81
      13'h147F: dout  = 8'b10000001; // 5247 : 129 - 0x81
      13'h1480: dout  = 8'b01101100; // 5248 : 108 - 0x6c -- Background 0x48
      13'h1481: dout  = 8'b11000110; // 5249 : 198 - 0xc6
      13'h1482: dout  = 8'b10000011; // 5250 : 131 - 0x83
      13'h1483: dout  = 8'b11111111; // 5251 : 255 - 0xff
      13'h1484: dout  = 8'b11111111; // 5252 : 255 - 0xff
      13'h1485: dout  = 8'b00000000; // 5253 :   0 - 0x0
      13'h1486: dout  = 8'b00000000; // 5254 :   0 - 0x0
      13'h1487: dout  = 8'b00000000; // 5255 :   0 - 0x0
      13'h1488: dout  = 8'b00000000; // 5256 :   0 - 0x0
      13'h1489: dout  = 8'b00000000; // 5257 :   0 - 0x0
      13'h148A: dout  = 8'b00000000; // 5258 :   0 - 0x0
      13'h148B: dout  = 8'b00000000; // 5259 :   0 - 0x0
      13'h148C: dout  = 8'b00000000; // 5260 :   0 - 0x0
      13'h148D: dout  = 8'b11111111; // 5261 : 255 - 0xff
      13'h148E: dout  = 8'b10000001; // 5262 : 129 - 0x81
      13'h148F: dout  = 8'b10000001; // 5263 : 129 - 0x81
      13'h1490: dout  = 8'b11000110; // 5264 : 198 - 0xc6 -- Background 0x49
      13'h1491: dout  = 8'b10000011; // 5265 : 131 - 0x83
      13'h1492: dout  = 8'b11111111; // 5266 : 255 - 0xff
      13'h1493: dout  = 8'b11111111; // 5267 : 255 - 0xff
      13'h1494: dout  = 8'b00000000; // 5268 :   0 - 0x0
      13'h1495: dout  = 8'b00000000; // 5269 :   0 - 0x0
      13'h1496: dout  = 8'b00000000; // 5270 :   0 - 0x0
      13'h1497: dout  = 8'b00000000; // 5271 :   0 - 0x0
      13'h1498: dout  = 8'b00000000; // 5272 :   0 - 0x0
      13'h1499: dout  = 8'b00000000; // 5273 :   0 - 0x0
      13'h149A: dout  = 8'b00000000; // 5274 :   0 - 0x0
      13'h149B: dout  = 8'b00000000; // 5275 :   0 - 0x0
      13'h149C: dout  = 8'b10000001; // 5276 : 129 - 0x81
      13'h149D: dout  = 8'b11111111; // 5277 : 255 - 0xff
      13'h149E: dout  = 8'b10000001; // 5278 : 129 - 0x81
      13'h149F: dout  = 8'b10000001; // 5279 : 129 - 0x81
      13'h14A0: dout  = 8'b10000011; // 5280 : 131 - 0x83 -- Background 0x4a
      13'h14A1: dout  = 8'b11111111; // 5281 : 255 - 0xff
      13'h14A2: dout  = 8'b11111111; // 5282 : 255 - 0xff
      13'h14A3: dout  = 8'b00000000; // 5283 :   0 - 0x0
      13'h14A4: dout  = 8'b00000000; // 5284 :   0 - 0x0
      13'h14A5: dout  = 8'b00000000; // 5285 :   0 - 0x0
      13'h14A6: dout  = 8'b00000000; // 5286 :   0 - 0x0
      13'h14A7: dout  = 8'b00000000; // 5287 :   0 - 0x0
      13'h14A8: dout  = 8'b00000000; // 5288 :   0 - 0x0
      13'h14A9: dout  = 8'b00000000; // 5289 :   0 - 0x0
      13'h14AA: dout  = 8'b00000000; // 5290 :   0 - 0x0
      13'h14AB: dout  = 8'b10000001; // 5291 : 129 - 0x81
      13'h14AC: dout  = 8'b10000001; // 5292 : 129 - 0x81
      13'h14AD: dout  = 8'b11111111; // 5293 : 255 - 0xff
      13'h14AE: dout  = 8'b10000001; // 5294 : 129 - 0x81
      13'h14AF: dout  = 8'b10000001; // 5295 : 129 - 0x81
      13'h14B0: dout  = 8'b11111111; // 5296 : 255 - 0xff -- Background 0x4b
      13'h14B1: dout  = 8'b11111111; // 5297 : 255 - 0xff
      13'h14B2: dout  = 8'b00000000; // 5298 :   0 - 0x0
      13'h14B3: dout  = 8'b00000000; // 5299 :   0 - 0x0
      13'h14B4: dout  = 8'b00000000; // 5300 :   0 - 0x0
      13'h14B5: dout  = 8'b00000000; // 5301 :   0 - 0x0
      13'h14B6: dout  = 8'b00000000; // 5302 :   0 - 0x0
      13'h14B7: dout  = 8'b00000000; // 5303 :   0 - 0x0
      13'h14B8: dout  = 8'b00000000; // 5304 :   0 - 0x0
      13'h14B9: dout  = 8'b00000000; // 5305 :   0 - 0x0
      13'h14BA: dout  = 8'b10000001; // 5306 : 129 - 0x81
      13'h14BB: dout  = 8'b10000001; // 5307 : 129 - 0x81
      13'h14BC: dout  = 8'b10000001; // 5308 : 129 - 0x81
      13'h14BD: dout  = 8'b11111111; // 5309 : 255 - 0xff
      13'h14BE: dout  = 8'b10000001; // 5310 : 129 - 0x81
      13'h14BF: dout  = 8'b10000001; // 5311 : 129 - 0x81
      13'h14C0: dout  = 8'b10111111; // 5312 : 191 - 0xbf -- Background 0x4c
      13'h14C1: dout  = 8'b01011111; // 5313 :  95 - 0x5f
      13'h14C2: dout  = 8'b01011111; // 5314 :  95 - 0x5f
      13'h14C3: dout  = 8'b01011111; // 5315 :  95 - 0x5f
      13'h14C4: dout  = 8'b00000000; // 5316 :   0 - 0x0
      13'h14C5: dout  = 8'b01011111; // 5317 :  95 - 0x5f
      13'h14C6: dout  = 8'b01010001; // 5318 :  81 - 0x51
      13'h14C7: dout  = 8'b01010101; // 5319 :  85 - 0x55
      13'h14C8: dout  = 8'b11111111; // 5320 : 255 - 0xff
      13'h14C9: dout  = 8'b01111111; // 5321 : 127 - 0x7f
      13'h14CA: dout  = 8'b01111111; // 5322 : 127 - 0x7f
      13'h14CB: dout  = 8'b01111111; // 5323 : 127 - 0x7f
      13'h14CC: dout  = 8'b01111111; // 5324 : 127 - 0x7f
      13'h14CD: dout  = 8'b01111111; // 5325 : 127 - 0x7f
      13'h14CE: dout  = 8'b01111111; // 5326 : 127 - 0x7f
      13'h14CF: dout  = 8'b01111111; // 5327 : 127 - 0x7f
      13'h14D0: dout  = 8'b01010001; // 5328 :  81 - 0x51 -- Background 0x4d
      13'h14D1: dout  = 8'b01011111; // 5329 :  95 - 0x5f
      13'h14D2: dout  = 8'b00000000; // 5330 :   0 - 0x0
      13'h14D3: dout  = 8'b01011111; // 5331 :  95 - 0x5f
      13'h14D4: dout  = 8'b01011111; // 5332 :  95 - 0x5f
      13'h14D5: dout  = 8'b01011111; // 5333 :  95 - 0x5f
      13'h14D6: dout  = 8'b01011111; // 5334 :  95 - 0x5f
      13'h14D7: dout  = 8'b10111111; // 5335 : 191 - 0xbf
      13'h14D8: dout  = 8'b01111111; // 5336 : 127 - 0x7f
      13'h14D9: dout  = 8'b01111111; // 5337 : 127 - 0x7f
      13'h14DA: dout  = 8'b01111111; // 5338 : 127 - 0x7f
      13'h14DB: dout  = 8'b01111111; // 5339 : 127 - 0x7f
      13'h14DC: dout  = 8'b01110010; // 5340 : 114 - 0x72
      13'h14DD: dout  = 8'b01111111; // 5341 : 127 - 0x7f
      13'h14DE: dout  = 8'b01111111; // 5342 : 127 - 0x7f
      13'h14DF: dout  = 8'b11111111; // 5343 : 255 - 0xff
      13'h14E0: dout  = 8'b11111111; // 5344 : 255 - 0xff -- Background 0x4e
      13'h14E1: dout  = 8'b11111110; // 5345 : 254 - 0xfe
      13'h14E2: dout  = 8'b11111110; // 5346 : 254 - 0xfe
      13'h14E3: dout  = 8'b11111110; // 5347 : 254 - 0xfe
      13'h14E4: dout  = 8'b00000000; // 5348 :   0 - 0x0
      13'h14E5: dout  = 8'b11111110; // 5349 : 254 - 0xfe
      13'h14E6: dout  = 8'b00100110; // 5350 :  38 - 0x26
      13'h14E7: dout  = 8'b00100110; // 5351 :  38 - 0x26
      13'h14E8: dout  = 8'b11111111; // 5352 : 255 - 0xff
      13'h14E9: dout  = 8'b11111110; // 5353 : 254 - 0xfe
      13'h14EA: dout  = 8'b11111110; // 5354 : 254 - 0xfe
      13'h14EB: dout  = 8'b11111110; // 5355 : 254 - 0xfe
      13'h14EC: dout  = 8'b11111110; // 5356 : 254 - 0xfe
      13'h14ED: dout  = 8'b11111110; // 5357 : 254 - 0xfe
      13'h14EE: dout  = 8'b11111110; // 5358 : 254 - 0xfe
      13'h14EF: dout  = 8'b11111110; // 5359 : 254 - 0xfe
      13'h14F0: dout  = 8'b00100010; // 5360 :  34 - 0x22 -- Background 0x4f
      13'h14F1: dout  = 8'b11111110; // 5361 : 254 - 0xfe
      13'h14F2: dout  = 8'b00000000; // 5362 :   0 - 0x0
      13'h14F3: dout  = 8'b11111110; // 5363 : 254 - 0xfe
      13'h14F4: dout  = 8'b11111110; // 5364 : 254 - 0xfe
      13'h14F5: dout  = 8'b11111110; // 5365 : 254 - 0xfe
      13'h14F6: dout  = 8'b11111110; // 5366 : 254 - 0xfe
      13'h14F7: dout  = 8'b11111111; // 5367 : 255 - 0xff
      13'h14F8: dout  = 8'b11111110; // 5368 : 254 - 0xfe
      13'h14F9: dout  = 8'b11111110; // 5369 : 254 - 0xfe
      13'h14FA: dout  = 8'b11111110; // 5370 : 254 - 0xfe
      13'h14FB: dout  = 8'b11111110; // 5371 : 254 - 0xfe
      13'h14FC: dout  = 8'b01001010; // 5372 :  74 - 0x4a
      13'h14FD: dout  = 8'b11111110; // 5373 : 254 - 0xfe
      13'h14FE: dout  = 8'b11111110; // 5374 : 254 - 0xfe
      13'h14FF: dout  = 8'b11111111; // 5375 : 255 - 0xff
      13'h1500: dout  = 8'b00000111; // 5376 :   7 - 0x7 -- Background 0x50
      13'h1501: dout  = 8'b00000000; // 5377 :   0 - 0x0
      13'h1502: dout  = 8'b00001111; // 5378 :  15 - 0xf
      13'h1503: dout  = 8'b00011111; // 5379 :  31 - 0x1f
      13'h1504: dout  = 8'b00011111; // 5380 :  31 - 0x1f
      13'h1505: dout  = 8'b00011111; // 5381 :  31 - 0x1f
      13'h1506: dout  = 8'b00011111; // 5382 :  31 - 0x1f
      13'h1507: dout  = 8'b00011111; // 5383 :  31 - 0x1f
      13'h1508: dout  = 8'b00000101; // 5384 :   5 - 0x5
      13'h1509: dout  = 8'b00001111; // 5385 :  15 - 0xf
      13'h150A: dout  = 8'b00001011; // 5386 :  11 - 0xb
      13'h150B: dout  = 8'b00011011; // 5387 :  27 - 0x1b
      13'h150C: dout  = 8'b00010011; // 5388 :  19 - 0x13
      13'h150D: dout  = 8'b00010011; // 5389 :  19 - 0x13
      13'h150E: dout  = 8'b00010011; // 5390 :  19 - 0x13
      13'h150F: dout  = 8'b00010011; // 5391 :  19 - 0x13
      13'h1510: dout  = 8'b00011111; // 5392 :  31 - 0x1f -- Background 0x51
      13'h1511: dout  = 8'b00011111; // 5393 :  31 - 0x1f
      13'h1512: dout  = 8'b00011111; // 5394 :  31 - 0x1f
      13'h1513: dout  = 8'b00011111; // 5395 :  31 - 0x1f
      13'h1514: dout  = 8'b00011111; // 5396 :  31 - 0x1f
      13'h1515: dout  = 8'b00001111; // 5397 :  15 - 0xf
      13'h1516: dout  = 8'b00000000; // 5398 :   0 - 0x0
      13'h1517: dout  = 8'b00000111; // 5399 :   7 - 0x7
      13'h1518: dout  = 8'b00010011; // 5400 :  19 - 0x13
      13'h1519: dout  = 8'b00010011; // 5401 :  19 - 0x13
      13'h151A: dout  = 8'b00010011; // 5402 :  19 - 0x13
      13'h151B: dout  = 8'b00010011; // 5403 :  19 - 0x13
      13'h151C: dout  = 8'b00011011; // 5404 :  27 - 0x1b
      13'h151D: dout  = 8'b00001011; // 5405 :  11 - 0xb
      13'h151E: dout  = 8'b00001111; // 5406 :  15 - 0xf
      13'h151F: dout  = 8'b00000101; // 5407 :   5 - 0x5
      13'h1520: dout  = 8'b00000111; // 5408 :   7 - 0x7 -- Background 0x52
      13'h1521: dout  = 8'b00000000; // 5409 :   0 - 0x0
      13'h1522: dout  = 8'b00001111; // 5410 :  15 - 0xf
      13'h1523: dout  = 8'b00011111; // 5411 :  31 - 0x1f
      13'h1524: dout  = 8'b00011111; // 5412 :  31 - 0x1f
      13'h1525: dout  = 8'b00011111; // 5413 :  31 - 0x1f
      13'h1526: dout  = 8'b00011111; // 5414 :  31 - 0x1f
      13'h1527: dout  = 8'b00011111; // 5415 :  31 - 0x1f
      13'h1528: dout  = 8'b00000101; // 5416 :   5 - 0x5
      13'h1529: dout  = 8'b00001111; // 5417 :  15 - 0xf
      13'h152A: dout  = 8'b00001011; // 5418 :  11 - 0xb
      13'h152B: dout  = 8'b00011011; // 5419 :  27 - 0x1b
      13'h152C: dout  = 8'b00010011; // 5420 :  19 - 0x13
      13'h152D: dout  = 8'b00010011; // 5421 :  19 - 0x13
      13'h152E: dout  = 8'b00010011; // 5422 :  19 - 0x13
      13'h152F: dout  = 8'b00010011; // 5423 :  19 - 0x13
      13'h1530: dout  = 8'b00011111; // 5424 :  31 - 0x1f -- Background 0x53
      13'h1531: dout  = 8'b00011111; // 5425 :  31 - 0x1f
      13'h1532: dout  = 8'b00011111; // 5426 :  31 - 0x1f
      13'h1533: dout  = 8'b00011111; // 5427 :  31 - 0x1f
      13'h1534: dout  = 8'b00011111; // 5428 :  31 - 0x1f
      13'h1535: dout  = 8'b00001111; // 5429 :  15 - 0xf
      13'h1536: dout  = 8'b00000000; // 5430 :   0 - 0x0
      13'h1537: dout  = 8'b00000111; // 5431 :   7 - 0x7
      13'h1538: dout  = 8'b00010011; // 5432 :  19 - 0x13
      13'h1539: dout  = 8'b00010011; // 5433 :  19 - 0x13
      13'h153A: dout  = 8'b00010011; // 5434 :  19 - 0x13
      13'h153B: dout  = 8'b00010011; // 5435 :  19 - 0x13
      13'h153C: dout  = 8'b00011011; // 5436 :  27 - 0x1b
      13'h153D: dout  = 8'b00001011; // 5437 :  11 - 0xb
      13'h153E: dout  = 8'b00001111; // 5438 :  15 - 0xf
      13'h153F: dout  = 8'b00000101; // 5439 :   5 - 0x5
      13'h1540: dout  = 8'b11100000; // 5440 : 224 - 0xe0 -- Background 0x54
      13'h1541: dout  = 8'b00000000; // 5441 :   0 - 0x0
      13'h1542: dout  = 8'b11110001; // 5442 : 241 - 0xf1
      13'h1543: dout  = 8'b11111011; // 5443 : 251 - 0xfb
      13'h1544: dout  = 8'b11111011; // 5444 : 251 - 0xfb
      13'h1545: dout  = 8'b11111011; // 5445 : 251 - 0xfb
      13'h1546: dout  = 8'b11111011; // 5446 : 251 - 0xfb
      13'h1547: dout  = 8'b11111011; // 5447 : 251 - 0xfb
      13'h1548: dout  = 8'b10100000; // 5448 : 160 - 0xa0
      13'h1549: dout  = 8'b11110001; // 5449 : 241 - 0xf1
      13'h154A: dout  = 8'b11010001; // 5450 : 209 - 0xd1
      13'h154B: dout  = 8'b11011011; // 5451 : 219 - 0xdb
      13'h154C: dout  = 8'b11001010; // 5452 : 202 - 0xca
      13'h154D: dout  = 8'b11001010; // 5453 : 202 - 0xca
      13'h154E: dout  = 8'b11001010; // 5454 : 202 - 0xca
      13'h154F: dout  = 8'b11001010; // 5455 : 202 - 0xca
      13'h1550: dout  = 8'b11111011; // 5456 : 251 - 0xfb -- Background 0x55
      13'h1551: dout  = 8'b11111011; // 5457 : 251 - 0xfb
      13'h1552: dout  = 8'b11111011; // 5458 : 251 - 0xfb
      13'h1553: dout  = 8'b11111011; // 5459 : 251 - 0xfb
      13'h1554: dout  = 8'b11111011; // 5460 : 251 - 0xfb
      13'h1555: dout  = 8'b11110001; // 5461 : 241 - 0xf1
      13'h1556: dout  = 8'b00000000; // 5462 :   0 - 0x0
      13'h1557: dout  = 8'b11100000; // 5463 : 224 - 0xe0
      13'h1558: dout  = 8'b11001010; // 5464 : 202 - 0xca
      13'h1559: dout  = 8'b11001010; // 5465 : 202 - 0xca
      13'h155A: dout  = 8'b11001010; // 5466 : 202 - 0xca
      13'h155B: dout  = 8'b11001010; // 5467 : 202 - 0xca
      13'h155C: dout  = 8'b11011011; // 5468 : 219 - 0xdb
      13'h155D: dout  = 8'b11010001; // 5469 : 209 - 0xd1
      13'h155E: dout  = 8'b11110001; // 5470 : 241 - 0xf1
      13'h155F: dout  = 8'b10100000; // 5471 : 160 - 0xa0
      13'h1560: dout  = 8'b11100000; // 5472 : 224 - 0xe0 -- Background 0x56
      13'h1561: dout  = 8'b00000000; // 5473 :   0 - 0x0
      13'h1562: dout  = 8'b11110001; // 5474 : 241 - 0xf1
      13'h1563: dout  = 8'b11111011; // 5475 : 251 - 0xfb
      13'h1564: dout  = 8'b11111011; // 5476 : 251 - 0xfb
      13'h1565: dout  = 8'b11111011; // 5477 : 251 - 0xfb
      13'h1566: dout  = 8'b11111011; // 5478 : 251 - 0xfb
      13'h1567: dout  = 8'b11111011; // 5479 : 251 - 0xfb
      13'h1568: dout  = 8'b10100000; // 5480 : 160 - 0xa0
      13'h1569: dout  = 8'b11110001; // 5481 : 241 - 0xf1
      13'h156A: dout  = 8'b11010001; // 5482 : 209 - 0xd1
      13'h156B: dout  = 8'b11011011; // 5483 : 219 - 0xdb
      13'h156C: dout  = 8'b11001010; // 5484 : 202 - 0xca
      13'h156D: dout  = 8'b11001010; // 5485 : 202 - 0xca
      13'h156E: dout  = 8'b11001010; // 5486 : 202 - 0xca
      13'h156F: dout  = 8'b11001010; // 5487 : 202 - 0xca
      13'h1570: dout  = 8'b11111011; // 5488 : 251 - 0xfb -- Background 0x57
      13'h1571: dout  = 8'b11111011; // 5489 : 251 - 0xfb
      13'h1572: dout  = 8'b11111011; // 5490 : 251 - 0xfb
      13'h1573: dout  = 8'b11111011; // 5491 : 251 - 0xfb
      13'h1574: dout  = 8'b11111011; // 5492 : 251 - 0xfb
      13'h1575: dout  = 8'b11110001; // 5493 : 241 - 0xf1
      13'h1576: dout  = 8'b00000000; // 5494 :   0 - 0x0
      13'h1577: dout  = 8'b11100000; // 5495 : 224 - 0xe0
      13'h1578: dout  = 8'b11001010; // 5496 : 202 - 0xca
      13'h1579: dout  = 8'b11001010; // 5497 : 202 - 0xca
      13'h157A: dout  = 8'b11001010; // 5498 : 202 - 0xca
      13'h157B: dout  = 8'b11001010; // 5499 : 202 - 0xca
      13'h157C: dout  = 8'b11011011; // 5500 : 219 - 0xdb
      13'h157D: dout  = 8'b11010001; // 5501 : 209 - 0xd1
      13'h157E: dout  = 8'b11110000; // 5502 : 240 - 0xf0
      13'h157F: dout  = 8'b10100000; // 5503 : 160 - 0xa0
      13'h1580: dout  = 8'b11111100; // 5504 : 252 - 0xfc -- Background 0x58
      13'h1581: dout  = 8'b00000000; // 5505 :   0 - 0x0
      13'h1582: dout  = 8'b11111110; // 5506 : 254 - 0xfe
      13'h1583: dout  = 8'b11111111; // 5507 : 255 - 0xff
      13'h1584: dout  = 8'b11111111; // 5508 : 255 - 0xff
      13'h1585: dout  = 8'b11111111; // 5509 : 255 - 0xff
      13'h1586: dout  = 8'b11111111; // 5510 : 255 - 0xff
      13'h1587: dout  = 8'b11111111; // 5511 : 255 - 0xff
      13'h1588: dout  = 8'b10110100; // 5512 : 180 - 0xb4
      13'h1589: dout  = 8'b11111110; // 5513 : 254 - 0xfe
      13'h158A: dout  = 8'b01111010; // 5514 : 122 - 0x7a
      13'h158B: dout  = 8'b01111011; // 5515 : 123 - 0x7b
      13'h158C: dout  = 8'b01111001; // 5516 : 121 - 0x79
      13'h158D: dout  = 8'b01111001; // 5517 : 121 - 0x79
      13'h158E: dout  = 8'b01111001; // 5518 : 121 - 0x79
      13'h158F: dout  = 8'b01111001; // 5519 : 121 - 0x79
      13'h1590: dout  = 8'b11111111; // 5520 : 255 - 0xff -- Background 0x59
      13'h1591: dout  = 8'b11111111; // 5521 : 255 - 0xff
      13'h1592: dout  = 8'b11111111; // 5522 : 255 - 0xff
      13'h1593: dout  = 8'b11111111; // 5523 : 255 - 0xff
      13'h1594: dout  = 8'b11111111; // 5524 : 255 - 0xff
      13'h1595: dout  = 8'b11111110; // 5525 : 254 - 0xfe
      13'h1596: dout  = 8'b00000000; // 5526 :   0 - 0x0
      13'h1597: dout  = 8'b11111100; // 5527 : 252 - 0xfc
      13'h1598: dout  = 8'b01111001; // 5528 : 121 - 0x79
      13'h1599: dout  = 8'b01111001; // 5529 : 121 - 0x79
      13'h159A: dout  = 8'b01111001; // 5530 : 121 - 0x79
      13'h159B: dout  = 8'b01111001; // 5531 : 121 - 0x79
      13'h159C: dout  = 8'b01111011; // 5532 : 123 - 0x7b
      13'h159D: dout  = 8'b01111010; // 5533 : 122 - 0x7a
      13'h159E: dout  = 8'b11111110; // 5534 : 254 - 0xfe
      13'h159F: dout  = 8'b10110100; // 5535 : 180 - 0xb4
      13'h15A0: dout  = 8'b11111100; // 5536 : 252 - 0xfc -- Background 0x5a
      13'h15A1: dout  = 8'b00000000; // 5537 :   0 - 0x0
      13'h15A2: dout  = 8'b11111110; // 5538 : 254 - 0xfe
      13'h15A3: dout  = 8'b11111111; // 5539 : 255 - 0xff
      13'h15A4: dout  = 8'b11111111; // 5540 : 255 - 0xff
      13'h15A5: dout  = 8'b11111111; // 5541 : 255 - 0xff
      13'h15A6: dout  = 8'b11111111; // 5542 : 255 - 0xff
      13'h15A7: dout  = 8'b11111111; // 5543 : 255 - 0xff
      13'h15A8: dout  = 8'b10110100; // 5544 : 180 - 0xb4
      13'h15A9: dout  = 8'b11111110; // 5545 : 254 - 0xfe
      13'h15AA: dout  = 8'b01111010; // 5546 : 122 - 0x7a
      13'h15AB: dout  = 8'b01111011; // 5547 : 123 - 0x7b
      13'h15AC: dout  = 8'b01111001; // 5548 : 121 - 0x79
      13'h15AD: dout  = 8'b01111001; // 5549 : 121 - 0x79
      13'h15AE: dout  = 8'b01111001; // 5550 : 121 - 0x79
      13'h15AF: dout  = 8'b01111001; // 5551 : 121 - 0x79
      13'h15B0: dout  = 8'b11111111; // 5552 : 255 - 0xff -- Background 0x5b
      13'h15B1: dout  = 8'b11111111; // 5553 : 255 - 0xff
      13'h15B2: dout  = 8'b11111111; // 5554 : 255 - 0xff
      13'h15B3: dout  = 8'b11111111; // 5555 : 255 - 0xff
      13'h15B4: dout  = 8'b11111111; // 5556 : 255 - 0xff
      13'h15B5: dout  = 8'b11111110; // 5557 : 254 - 0xfe
      13'h15B6: dout  = 8'b00000000; // 5558 :   0 - 0x0
      13'h15B7: dout  = 8'b11111100; // 5559 : 252 - 0xfc
      13'h15B8: dout  = 8'b01111001; // 5560 : 121 - 0x79
      13'h15B9: dout  = 8'b01111001; // 5561 : 121 - 0x79
      13'h15BA: dout  = 8'b01111001; // 5562 : 121 - 0x79
      13'h15BB: dout  = 8'b01111001; // 5563 : 121 - 0x79
      13'h15BC: dout  = 8'b01111011; // 5564 : 123 - 0x7b
      13'h15BD: dout  = 8'b01111010; // 5565 : 122 - 0x7a
      13'h15BE: dout  = 8'b11111110; // 5566 : 254 - 0xfe
      13'h15BF: dout  = 8'b10110100; // 5567 : 180 - 0xb4
      13'h15C0: dout  = 8'b00000000; // 5568 :   0 - 0x0 -- Background 0x5c
      13'h15C1: dout  = 8'b00000000; // 5569 :   0 - 0x0
      13'h15C2: dout  = 8'b00011111; // 5570 :  31 - 0x1f
      13'h15C3: dout  = 8'b00010000; // 5571 :  16 - 0x10
      13'h15C4: dout  = 8'b00010000; // 5572 :  16 - 0x10
      13'h15C5: dout  = 8'b00011111; // 5573 :  31 - 0x1f
      13'h15C6: dout  = 8'b00000000; // 5574 :   0 - 0x0
      13'h15C7: dout  = 8'b00000000; // 5575 :   0 - 0x0
      13'h15C8: dout  = 8'b01111111; // 5576 : 127 - 0x7f
      13'h15C9: dout  = 8'b10111111; // 5577 : 191 - 0xbf
      13'h15CA: dout  = 8'b11111111; // 5578 : 255 - 0xff
      13'h15CB: dout  = 8'b10110010; // 5579 : 178 - 0xb2
      13'h15CC: dout  = 8'b10110001; // 5580 : 177 - 0xb1
      13'h15CD: dout  = 8'b11111111; // 5581 : 255 - 0xff
      13'h15CE: dout  = 8'b10111111; // 5582 : 191 - 0xbf
      13'h15CF: dout  = 8'b01111111; // 5583 : 127 - 0x7f
      13'h15D0: dout  = 8'b00000000; // 5584 :   0 - 0x0 -- Background 0x5d
      13'h15D1: dout  = 8'b00000000; // 5585 :   0 - 0x0
      13'h15D2: dout  = 8'b11111000; // 5586 : 248 - 0xf8
      13'h15D3: dout  = 8'b00001000; // 5587 :   8 - 0x8
      13'h15D4: dout  = 8'b00001000; // 5588 :   8 - 0x8
      13'h15D5: dout  = 8'b11111000; // 5589 : 248 - 0xf8
      13'h15D6: dout  = 8'b00000000; // 5590 :   0 - 0x0
      13'h15D7: dout  = 8'b00000000; // 5591 :   0 - 0x0
      13'h15D8: dout  = 8'b11111110; // 5592 : 254 - 0xfe
      13'h15D9: dout  = 8'b11111101; // 5593 : 253 - 0xfd
      13'h15DA: dout  = 8'b11111111; // 5594 : 255 - 0xff
      13'h15DB: dout  = 8'b11001101; // 5595 : 205 - 0xcd
      13'h15DC: dout  = 8'b01101101; // 5596 : 109 - 0x6d
      13'h15DD: dout  = 8'b11111111; // 5597 : 255 - 0xff
      13'h15DE: dout  = 8'b11111101; // 5598 : 253 - 0xfd
      13'h15DF: dout  = 8'b11111110; // 5599 : 254 - 0xfe
      13'h15E0: dout  = 8'b00000000; // 5600 :   0 - 0x0 -- Background 0x5e
      13'h15E1: dout  = 8'b00000001; // 5601 :   1 - 0x1
      13'h15E2: dout  = 8'b00000010; // 5602 :   2 - 0x2
      13'h15E3: dout  = 8'b00000010; // 5603 :   2 - 0x2
      13'h15E4: dout  = 8'b11110001; // 5604 : 241 - 0xf1
      13'h15E5: dout  = 8'b00001000; // 5605 :   8 - 0x8
      13'h15E6: dout  = 8'b00000100; // 5606 :   4 - 0x4
      13'h15E7: dout  = 8'b00000011; // 5607 :   3 - 0x3
      13'h15E8: dout  = 8'b11111111; // 5608 : 255 - 0xff
      13'h15E9: dout  = 8'b11111111; // 5609 : 255 - 0xff
      13'h15EA: dout  = 8'b10101110; // 5610 : 174 - 0xae
      13'h15EB: dout  = 8'b11111110; // 5611 : 254 - 0xfe
      13'h15EC: dout  = 8'b11111111; // 5612 : 255 - 0xff
      13'h15ED: dout  = 8'b00001111; // 5613 :  15 - 0xf
      13'h15EE: dout  = 8'b00000111; // 5614 :   7 - 0x7
      13'h15EF: dout  = 8'b00000011; // 5615 :   3 - 0x3
      13'h15F0: dout  = 8'b00000000; // 5616 :   0 - 0x0 -- Background 0x5f
      13'h15F1: dout  = 8'b10000000; // 5617 : 128 - 0x80
      13'h15F2: dout  = 8'b01000000; // 5618 :  64 - 0x40
      13'h15F3: dout  = 8'b01000000; // 5619 :  64 - 0x40
      13'h15F4: dout  = 8'b10001111; // 5620 : 143 - 0x8f
      13'h15F5: dout  = 8'b00010000; // 5621 :  16 - 0x10
      13'h15F6: dout  = 8'b00100000; // 5622 :  32 - 0x20
      13'h15F7: dout  = 8'b11000000; // 5623 : 192 - 0xc0
      13'h15F8: dout  = 8'b11111111; // 5624 : 255 - 0xff
      13'h15F9: dout  = 8'b11111111; // 5625 : 255 - 0xff
      13'h15FA: dout  = 8'b01110101; // 5626 : 117 - 0x75
      13'h15FB: dout  = 8'b01111111; // 5627 : 127 - 0x7f
      13'h15FC: dout  = 8'b11111111; // 5628 : 255 - 0xff
      13'h15FD: dout  = 8'b11110000; // 5629 : 240 - 0xf0
      13'h15FE: dout  = 8'b11100000; // 5630 : 224 - 0xe0
      13'h15FF: dout  = 8'b11000000; // 5631 : 192 - 0xc0
      13'h1600: dout  = 8'b00000011; // 5632 :   3 - 0x3 -- Background 0x60
      13'h1601: dout  = 8'b00000100; // 5633 :   4 - 0x4
      13'h1602: dout  = 8'b00001000; // 5634 :   8 - 0x8
      13'h1603: dout  = 8'b11110001; // 5635 : 241 - 0xf1
      13'h1604: dout  = 8'b00000010; // 5636 :   2 - 0x2
      13'h1605: dout  = 8'b00000010; // 5637 :   2 - 0x2
      13'h1606: dout  = 8'b00000001; // 5638 :   1 - 0x1
      13'h1607: dout  = 8'b00000000; // 5639 :   0 - 0x0
      13'h1608: dout  = 8'b00000011; // 5640 :   3 - 0x3
      13'h1609: dout  = 8'b00000111; // 5641 :   7 - 0x7
      13'h160A: dout  = 8'b00001111; // 5642 :  15 - 0xf
      13'h160B: dout  = 8'b11111111; // 5643 : 255 - 0xff
      13'h160C: dout  = 8'b11111110; // 5644 : 254 - 0xfe
      13'h160D: dout  = 8'b10101110; // 5645 : 174 - 0xae
      13'h160E: dout  = 8'b11111111; // 5646 : 255 - 0xff
      13'h160F: dout  = 8'b11111111; // 5647 : 255 - 0xff
      13'h1610: dout  = 8'b11000000; // 5648 : 192 - 0xc0 -- Background 0x61
      13'h1611: dout  = 8'b00100000; // 5649 :  32 - 0x20
      13'h1612: dout  = 8'b00010000; // 5650 :  16 - 0x10
      13'h1613: dout  = 8'b10001111; // 5651 : 143 - 0x8f
      13'h1614: dout  = 8'b01000000; // 5652 :  64 - 0x40
      13'h1615: dout  = 8'b01000000; // 5653 :  64 - 0x40
      13'h1616: dout  = 8'b10000000; // 5654 : 128 - 0x80
      13'h1617: dout  = 8'b00000000; // 5655 :   0 - 0x0
      13'h1618: dout  = 8'b11000000; // 5656 : 192 - 0xc0
      13'h1619: dout  = 8'b11100000; // 5657 : 224 - 0xe0
      13'h161A: dout  = 8'b11110000; // 5658 : 240 - 0xf0
      13'h161B: dout  = 8'b11111111; // 5659 : 255 - 0xff
      13'h161C: dout  = 8'b01111111; // 5660 : 127 - 0x7f
      13'h161D: dout  = 8'b01110101; // 5661 : 117 - 0x75
      13'h161E: dout  = 8'b11111111; // 5662 : 255 - 0xff
      13'h161F: dout  = 8'b11111111; // 5663 : 255 - 0xff
      13'h1620: dout  = 8'b11111111; // 5664 : 255 - 0xff -- Background 0x62
      13'h1621: dout  = 8'b11111111; // 5665 : 255 - 0xff
      13'h1622: dout  = 8'b11000011; // 5666 : 195 - 0xc3
      13'h1623: dout  = 8'b10000001; // 5667 : 129 - 0x81
      13'h1624: dout  = 8'b10000001; // 5668 : 129 - 0x81
      13'h1625: dout  = 8'b11000011; // 5669 : 195 - 0xc3
      13'h1626: dout  = 8'b11111111; // 5670 : 255 - 0xff
      13'h1627: dout  = 8'b11111111; // 5671 : 255 - 0xff
      13'h1628: dout  = 8'b11111111; // 5672 : 255 - 0xff
      13'h1629: dout  = 8'b00000000; // 5673 :   0 - 0x0
      13'h162A: dout  = 8'b11000011; // 5674 : 195 - 0xc3
      13'h162B: dout  = 8'b10000001; // 5675 : 129 - 0x81
      13'h162C: dout  = 8'b10000001; // 5676 : 129 - 0x81
      13'h162D: dout  = 8'b11000011; // 5677 : 195 - 0xc3
      13'h162E: dout  = 8'b11111111; // 5678 : 255 - 0xff
      13'h162F: dout  = 8'b00000000; // 5679 :   0 - 0x0
      13'h1630: dout  = 8'b11111111; // 5680 : 255 - 0xff -- Background 0x63
      13'h1631: dout  = 8'b10011001; // 5681 : 153 - 0x99
      13'h1632: dout  = 8'b00000000; // 5682 :   0 - 0x0
      13'h1633: dout  = 8'b00000000; // 5683 :   0 - 0x0
      13'h1634: dout  = 8'b00000000; // 5684 :   0 - 0x0
      13'h1635: dout  = 8'b10000001; // 5685 : 129 - 0x81
      13'h1636: dout  = 8'b10000001; // 5686 : 129 - 0x81
      13'h1637: dout  = 8'b10000001; // 5687 : 129 - 0x81
      13'h1638: dout  = 8'b10000001; // 5688 : 129 - 0x81
      13'h1639: dout  = 8'b01100110; // 5689 : 102 - 0x66
      13'h163A: dout  = 8'b01111110; // 5690 : 126 - 0x7e
      13'h163B: dout  = 8'b01111110; // 5691 : 126 - 0x7e
      13'h163C: dout  = 8'b01111110; // 5692 : 126 - 0x7e
      13'h163D: dout  = 8'b11111111; // 5693 : 255 - 0xff
      13'h163E: dout  = 8'b11111111; // 5694 : 255 - 0xff
      13'h163F: dout  = 8'b01111110; // 5695 : 126 - 0x7e
      13'h1640: dout  = 8'b00000000; // 5696 :   0 - 0x0 -- Background 0x64
      13'h1641: dout  = 8'b00000000; // 5697 :   0 - 0x0
      13'h1642: dout  = 8'b00000000; // 5698 :   0 - 0x0
      13'h1643: dout  = 8'b00000000; // 5699 :   0 - 0x0
      13'h1644: dout  = 8'b01100000; // 5700 :  96 - 0x60
      13'h1645: dout  = 8'b01100000; // 5701 :  96 - 0x60
      13'h1646: dout  = 8'b00000000; // 5702 :   0 - 0x0
      13'h1647: dout  = 8'b00000000; // 5703 :   0 - 0x0
      13'h1648: dout  = 8'b00000000; // 5704 :   0 - 0x0
      13'h1649: dout  = 8'b00000000; // 5705 :   0 - 0x0
      13'h164A: dout  = 8'b00000000; // 5706 :   0 - 0x0
      13'h164B: dout  = 8'b00000000; // 5707 :   0 - 0x0
      13'h164C: dout  = 8'b00000000; // 5708 :   0 - 0x0
      13'h164D: dout  = 8'b00000000; // 5709 :   0 - 0x0
      13'h164E: dout  = 8'b00000000; // 5710 :   0 - 0x0
      13'h164F: dout  = 8'b00000000; // 5711 :   0 - 0x0
      13'h1650: dout  = 8'b00000000; // 5712 :   0 - 0x0 -- Background 0x65
      13'h1651: dout  = 8'b00000000; // 5713 :   0 - 0x0
      13'h1652: dout  = 8'b00000000; // 5714 :   0 - 0x0
      13'h1653: dout  = 8'b00000000; // 5715 :   0 - 0x0
      13'h1654: dout  = 8'b01101100; // 5716 : 108 - 0x6c
      13'h1655: dout  = 8'b01101100; // 5717 : 108 - 0x6c
      13'h1656: dout  = 8'b00001000; // 5718 :   8 - 0x8
      13'h1657: dout  = 8'b00000000; // 5719 :   0 - 0x0
      13'h1658: dout  = 8'b00000000; // 5720 :   0 - 0x0
      13'h1659: dout  = 8'b00000000; // 5721 :   0 - 0x0
      13'h165A: dout  = 8'b00000000; // 5722 :   0 - 0x0
      13'h165B: dout  = 8'b00000000; // 5723 :   0 - 0x0
      13'h165C: dout  = 8'b00000000; // 5724 :   0 - 0x0
      13'h165D: dout  = 8'b00000000; // 5725 :   0 - 0x0
      13'h165E: dout  = 8'b00000000; // 5726 :   0 - 0x0
      13'h165F: dout  = 8'b00000000; // 5727 :   0 - 0x0
      13'h1660: dout  = 8'b00111100; // 5728 :  60 - 0x3c -- Background 0x66
      13'h1661: dout  = 8'b00011000; // 5729 :  24 - 0x18
      13'h1662: dout  = 8'b00011000; // 5730 :  24 - 0x18
      13'h1663: dout  = 8'b00011000; // 5731 :  24 - 0x18
      13'h1664: dout  = 8'b00011000; // 5732 :  24 - 0x18
      13'h1665: dout  = 8'b00011000; // 5733 :  24 - 0x18
      13'h1666: dout  = 8'b00111100; // 5734 :  60 - 0x3c
      13'h1667: dout  = 8'b00000000; // 5735 :   0 - 0x0
      13'h1668: dout  = 8'b00000000; // 5736 :   0 - 0x0
      13'h1669: dout  = 8'b00000000; // 5737 :   0 - 0x0
      13'h166A: dout  = 8'b00000000; // 5738 :   0 - 0x0
      13'h166B: dout  = 8'b00000000; // 5739 :   0 - 0x0
      13'h166C: dout  = 8'b00000000; // 5740 :   0 - 0x0
      13'h166D: dout  = 8'b00000000; // 5741 :   0 - 0x0
      13'h166E: dout  = 8'b00000000; // 5742 :   0 - 0x0
      13'h166F: dout  = 8'b00000000; // 5743 :   0 - 0x0
      13'h1670: dout  = 8'b11111111; // 5744 : 255 - 0xff -- Background 0x67
      13'h1671: dout  = 8'b01100110; // 5745 : 102 - 0x66
      13'h1672: dout  = 8'b01100110; // 5746 : 102 - 0x66
      13'h1673: dout  = 8'b01100110; // 5747 : 102 - 0x66
      13'h1674: dout  = 8'b01100110; // 5748 : 102 - 0x66
      13'h1675: dout  = 8'b01100110; // 5749 : 102 - 0x66
      13'h1676: dout  = 8'b01100110; // 5750 : 102 - 0x66
      13'h1677: dout  = 8'b11111111; // 5751 : 255 - 0xff
      13'h1678: dout  = 8'b00000000; // 5752 :   0 - 0x0
      13'h1679: dout  = 8'b00000000; // 5753 :   0 - 0x0
      13'h167A: dout  = 8'b00000000; // 5754 :   0 - 0x0
      13'h167B: dout  = 8'b00000000; // 5755 :   0 - 0x0
      13'h167C: dout  = 8'b00000000; // 5756 :   0 - 0x0
      13'h167D: dout  = 8'b00000000; // 5757 :   0 - 0x0
      13'h167E: dout  = 8'b00000000; // 5758 :   0 - 0x0
      13'h167F: dout  = 8'b00000000; // 5759 :   0 - 0x0
      13'h1680: dout  = 8'b00000011; // 5760 :   3 - 0x3 -- Background 0x68
      13'h1681: dout  = 8'b00000001; // 5761 :   1 - 0x1
      13'h1682: dout  = 8'b00000000; // 5762 :   0 - 0x0
      13'h1683: dout  = 8'b00000000; // 5763 :   0 - 0x0
      13'h1684: dout  = 8'b00000000; // 5764 :   0 - 0x0
      13'h1685: dout  = 8'b00000000; // 5765 :   0 - 0x0
      13'h1686: dout  = 8'b00000000; // 5766 :   0 - 0x0
      13'h1687: dout  = 8'b00000000; // 5767 :   0 - 0x0
      13'h1688: dout  = 8'b00000011; // 5768 :   3 - 0x3
      13'h1689: dout  = 8'b00000001; // 5769 :   1 - 0x1
      13'h168A: dout  = 8'b00000000; // 5770 :   0 - 0x0
      13'h168B: dout  = 8'b00000000; // 5771 :   0 - 0x0
      13'h168C: dout  = 8'b00000000; // 5772 :   0 - 0x0
      13'h168D: dout  = 8'b00000000; // 5773 :   0 - 0x0
      13'h168E: dout  = 8'b00000000; // 5774 :   0 - 0x0
      13'h168F: dout  = 8'b00000000; // 5775 :   0 - 0x0
      13'h1690: dout  = 8'b10000011; // 5776 : 131 - 0x83 -- Background 0x69
      13'h1691: dout  = 8'b11010001; // 5777 : 209 - 0xd1
      13'h1692: dout  = 8'b11100001; // 5778 : 225 - 0xe1
      13'h1693: dout  = 8'b11010001; // 5779 : 209 - 0xd1
      13'h1694: dout  = 8'b00000010; // 5780 :   2 - 0x2
      13'h1695: dout  = 8'b10000100; // 5781 : 132 - 0x84
      13'h1696: dout  = 8'b11110000; // 5782 : 240 - 0xf0
      13'h1697: dout  = 8'b11001110; // 5783 : 206 - 0xce
      13'h1698: dout  = 8'b11111111; // 5784 : 255 - 0xff
      13'h1699: dout  = 8'b11111111; // 5785 : 255 - 0xff
      13'h169A: dout  = 8'b11111111; // 5786 : 255 - 0xff
      13'h169B: dout  = 8'b11111111; // 5787 : 255 - 0xff
      13'h169C: dout  = 8'b11111111; // 5788 : 255 - 0xff
      13'h169D: dout  = 8'b11111111; // 5789 : 255 - 0xff
      13'h169E: dout  = 8'b11111111; // 5790 : 255 - 0xff
      13'h169F: dout  = 8'b11111111; // 5791 : 255 - 0xff
      13'h16A0: dout  = 8'b11000000; // 5792 : 192 - 0xc0 -- Background 0x6a
      13'h16A1: dout  = 8'b10000000; // 5793 : 128 - 0x80
      13'h16A2: dout  = 8'b00000000; // 5794 :   0 - 0x0
      13'h16A3: dout  = 8'b00000000; // 5795 :   0 - 0x0
      13'h16A4: dout  = 8'b00000000; // 5796 :   0 - 0x0
      13'h16A5: dout  = 8'b00000000; // 5797 :   0 - 0x0
      13'h16A6: dout  = 8'b00000000; // 5798 :   0 - 0x0
      13'h16A7: dout  = 8'b00000000; // 5799 :   0 - 0x0
      13'h16A8: dout  = 8'b11000000; // 5800 : 192 - 0xc0
      13'h16A9: dout  = 8'b10000000; // 5801 : 128 - 0x80
      13'h16AA: dout  = 8'b00000000; // 5802 :   0 - 0x0
      13'h16AB: dout  = 8'b00000000; // 5803 :   0 - 0x0
      13'h16AC: dout  = 8'b00000000; // 5804 :   0 - 0x0
      13'h16AD: dout  = 8'b00000000; // 5805 :   0 - 0x0
      13'h16AE: dout  = 8'b00000000; // 5806 :   0 - 0x0
      13'h16AF: dout  = 8'b00000000; // 5807 :   0 - 0x0
      13'h16B0: dout  = 8'b11000001; // 5808 : 193 - 0xc1 -- Background 0x6b
      13'h16B1: dout  = 8'b10001011; // 5809 : 139 - 0x8b
      13'h16B2: dout  = 8'b10000111; // 5810 : 135 - 0x87
      13'h16B3: dout  = 8'b10001011; // 5811 : 139 - 0x8b
      13'h16B4: dout  = 8'b01000000; // 5812 :  64 - 0x40
      13'h16B5: dout  = 8'b00100001; // 5813 :  33 - 0x21
      13'h16B6: dout  = 8'b00001111; // 5814 :  15 - 0xf
      13'h16B7: dout  = 8'b11010011; // 5815 : 211 - 0xd3
      13'h16B8: dout  = 8'b11111111; // 5816 : 255 - 0xff
      13'h16B9: dout  = 8'b11111111; // 5817 : 255 - 0xff
      13'h16BA: dout  = 8'b11111111; // 5818 : 255 - 0xff
      13'h16BB: dout  = 8'b11111111; // 5819 : 255 - 0xff
      13'h16BC: dout  = 8'b11111111; // 5820 : 255 - 0xff
      13'h16BD: dout  = 8'b11111111; // 5821 : 255 - 0xff
      13'h16BE: dout  = 8'b11111111; // 5822 : 255 - 0xff
      13'h16BF: dout  = 8'b11111111; // 5823 : 255 - 0xff
      13'h16C0: dout  = 8'b11111111; // 5824 : 255 - 0xff -- Background 0x6c
      13'h16C1: dout  = 8'b11111111; // 5825 : 255 - 0xff
      13'h16C2: dout  = 8'b11111111; // 5826 : 255 - 0xff
      13'h16C3: dout  = 8'b00011111; // 5827 :  31 - 0x1f
      13'h16C4: dout  = 8'b00001111; // 5828 :  15 - 0xf
      13'h16C5: dout  = 8'b00011110; // 5829 :  30 - 0x1e
      13'h16C6: dout  = 8'b00111111; // 5830 :  63 - 0x3f
      13'h16C7: dout  = 8'b01111111; // 5831 : 127 - 0x7f
      13'h16C8: dout  = 8'b11111111; // 5832 : 255 - 0xff
      13'h16C9: dout  = 8'b11111111; // 5833 : 255 - 0xff
      13'h16CA: dout  = 8'b11111111; // 5834 : 255 - 0xff
      13'h16CB: dout  = 8'b00011111; // 5835 :  31 - 0x1f
      13'h16CC: dout  = 8'b00011111; // 5836 :  31 - 0x1f
      13'h16CD: dout  = 8'b00111111; // 5837 :  63 - 0x3f
      13'h16CE: dout  = 8'b01111111; // 5838 : 127 - 0x7f
      13'h16CF: dout  = 8'b11111111; // 5839 : 255 - 0xff
      13'h16D0: dout  = 8'b11111111; // 5840 : 255 - 0xff -- Background 0x6d
      13'h16D1: dout  = 8'b11111111; // 5841 : 255 - 0xff
      13'h16D2: dout  = 8'b11111111; // 5842 : 255 - 0xff
      13'h16D3: dout  = 8'b11111000; // 5843 : 248 - 0xf8
      13'h16D4: dout  = 8'b11110000; // 5844 : 240 - 0xf0
      13'h16D5: dout  = 8'b01111000; // 5845 : 120 - 0x78
      13'h16D6: dout  = 8'b11111100; // 5846 : 252 - 0xfc
      13'h16D7: dout  = 8'b11111110; // 5847 : 254 - 0xfe
      13'h16D8: dout  = 8'b11111111; // 5848 : 255 - 0xff
      13'h16D9: dout  = 8'b11111111; // 5849 : 255 - 0xff
      13'h16DA: dout  = 8'b11111111; // 5850 : 255 - 0xff
      13'h16DB: dout  = 8'b11111000; // 5851 : 248 - 0xf8
      13'h16DC: dout  = 8'b11111000; // 5852 : 248 - 0xf8
      13'h16DD: dout  = 8'b11111100; // 5853 : 252 - 0xfc
      13'h16DE: dout  = 8'b11111110; // 5854 : 254 - 0xfe
      13'h16DF: dout  = 8'b11111111; // 5855 : 255 - 0xff
      13'h16E0: dout  = 8'b00000000; // 5856 :   0 - 0x0 -- Background 0x6e
      13'h16E1: dout  = 8'b00000000; // 5857 :   0 - 0x0
      13'h16E2: dout  = 8'b00000000; // 5858 :   0 - 0x0
      13'h16E3: dout  = 8'b00000000; // 5859 :   0 - 0x0
      13'h16E4: dout  = 8'b00000000; // 5860 :   0 - 0x0
      13'h16E5: dout  = 8'b00111100; // 5861 :  60 - 0x3c
      13'h16E6: dout  = 8'b01000010; // 5862 :  66 - 0x42
      13'h16E7: dout  = 8'b10000001; // 5863 : 129 - 0x81
      13'h16E8: dout  = 8'b00000000; // 5864 :   0 - 0x0
      13'h16E9: dout  = 8'b00000000; // 5865 :   0 - 0x0
      13'h16EA: dout  = 8'b00000000; // 5866 :   0 - 0x0
      13'h16EB: dout  = 8'b00000000; // 5867 :   0 - 0x0
      13'h16EC: dout  = 8'b00000000; // 5868 :   0 - 0x0
      13'h16ED: dout  = 8'b00111100; // 5869 :  60 - 0x3c
      13'h16EE: dout  = 8'b01000010; // 5870 :  66 - 0x42
      13'h16EF: dout  = 8'b10000001; // 5871 : 129 - 0x81
      13'h16F0: dout  = 8'b10000001; // 5872 : 129 - 0x81 -- Background 0x6f
      13'h16F1: dout  = 8'b10111101; // 5873 : 189 - 0xbd
      13'h16F2: dout  = 8'b01111110; // 5874 : 126 - 0x7e
      13'h16F3: dout  = 8'b11111111; // 5875 : 255 - 0xff
      13'h16F4: dout  = 8'b11100111; // 5876 : 231 - 0xe7
      13'h16F5: dout  = 8'b11111111; // 5877 : 255 - 0xff
      13'h16F6: dout  = 8'b11111111; // 5878 : 255 - 0xff
      13'h16F7: dout  = 8'b11111111; // 5879 : 255 - 0xff
      13'h16F8: dout  = 8'b10000001; // 5880 : 129 - 0x81
      13'h16F9: dout  = 8'b10111101; // 5881 : 189 - 0xbd
      13'h16FA: dout  = 8'b01111110; // 5882 : 126 - 0x7e
      13'h16FB: dout  = 8'b10100101; // 5883 : 165 - 0xa5
      13'h16FC: dout  = 8'b11011011; // 5884 : 219 - 0xdb
      13'h16FD: dout  = 8'b11100111; // 5885 : 231 - 0xe7
      13'h16FE: dout  = 8'b11111111; // 5886 : 255 - 0xff
      13'h16FF: dout  = 8'b11111111; // 5887 : 255 - 0xff
      13'h1700: dout  = 8'b00000001; // 5888 :   1 - 0x1 -- Background 0x70
      13'h1701: dout  = 8'b00000111; // 5889 :   7 - 0x7
      13'h1702: dout  = 8'b00011111; // 5890 :  31 - 0x1f
      13'h1703: dout  = 8'b00111111; // 5891 :  63 - 0x3f
      13'h1704: dout  = 8'b01111111; // 5892 : 127 - 0x7f
      13'h1705: dout  = 8'b11111111; // 5893 : 255 - 0xff
      13'h1706: dout  = 8'b11111111; // 5894 : 255 - 0xff
      13'h1707: dout  = 8'b11011101; // 5895 : 221 - 0xdd
      13'h1708: dout  = 8'b00000000; // 5896 :   0 - 0x0
      13'h1709: dout  = 8'b00000101; // 5897 :   5 - 0x5
      13'h170A: dout  = 8'b00011001; // 5898 :  25 - 0x19
      13'h170B: dout  = 8'b00110011; // 5899 :  51 - 0x33
      13'h170C: dout  = 8'b01100011; // 5900 :  99 - 0x63
      13'h170D: dout  = 8'b11000111; // 5901 : 199 - 0xc7
      13'h170E: dout  = 8'b11000111; // 5902 : 199 - 0xc7
      13'h170F: dout  = 8'b11000100; // 5903 : 196 - 0xc4
      13'h1710: dout  = 8'b10001001; // 5904 : 137 - 0x89 -- Background 0x71
      13'h1711: dout  = 8'b00000001; // 5905 :   1 - 0x1
      13'h1712: dout  = 8'b00000001; // 5906 :   1 - 0x1
      13'h1713: dout  = 8'b00000001; // 5907 :   1 - 0x1
      13'h1714: dout  = 8'b00000001; // 5908 :   1 - 0x1
      13'h1715: dout  = 8'b00000001; // 5909 :   1 - 0x1
      13'h1716: dout  = 8'b00000000; // 5910 :   0 - 0x0
      13'h1717: dout  = 8'b00000000; // 5911 :   0 - 0x0
      13'h1718: dout  = 8'b10000000; // 5912 : 128 - 0x80
      13'h1719: dout  = 8'b00000000; // 5913 :   0 - 0x0
      13'h171A: dout  = 8'b00000000; // 5914 :   0 - 0x0
      13'h171B: dout  = 8'b00000001; // 5915 :   1 - 0x1
      13'h171C: dout  = 8'b00000001; // 5916 :   1 - 0x1
      13'h171D: dout  = 8'b00000001; // 5917 :   1 - 0x1
      13'h171E: dout  = 8'b00000000; // 5918 :   0 - 0x0
      13'h171F: dout  = 8'b00000000; // 5919 :   0 - 0x0
      13'h1720: dout  = 8'b10000000; // 5920 : 128 - 0x80 -- Background 0x72
      13'h1721: dout  = 8'b11100000; // 5921 : 224 - 0xe0
      13'h1722: dout  = 8'b11111000; // 5922 : 248 - 0xf8
      13'h1723: dout  = 8'b11111100; // 5923 : 252 - 0xfc
      13'h1724: dout  = 8'b11111110; // 5924 : 254 - 0xfe
      13'h1725: dout  = 8'b11111111; // 5925 : 255 - 0xff
      13'h1726: dout  = 8'b11111111; // 5926 : 255 - 0xff
      13'h1727: dout  = 8'b00111011; // 5927 :  59 - 0x3b
      13'h1728: dout  = 8'b00000000; // 5928 :   0 - 0x0
      13'h1729: dout  = 8'b10100000; // 5929 : 160 - 0xa0
      13'h172A: dout  = 8'b10011000; // 5930 : 152 - 0x98
      13'h172B: dout  = 8'b11001100; // 5931 : 204 - 0xcc
      13'h172C: dout  = 8'b11000110; // 5932 : 198 - 0xc6
      13'h172D: dout  = 8'b11100011; // 5933 : 227 - 0xe3
      13'h172E: dout  = 8'b11100011; // 5934 : 227 - 0xe3
      13'h172F: dout  = 8'b00100011; // 5935 :  35 - 0x23
      13'h1730: dout  = 8'b00010001; // 5936 :  17 - 0x11 -- Background 0x73
      13'h1731: dout  = 8'b00000000; // 5937 :   0 - 0x0
      13'h1732: dout  = 8'b00000000; // 5938 :   0 - 0x0
      13'h1733: dout  = 8'b00000000; // 5939 :   0 - 0x0
      13'h1734: dout  = 8'b00000000; // 5940 :   0 - 0x0
      13'h1735: dout  = 8'b01000000; // 5941 :  64 - 0x40
      13'h1736: dout  = 8'b10000000; // 5942 : 128 - 0x80
      13'h1737: dout  = 8'b00000000; // 5943 :   0 - 0x0
      13'h1738: dout  = 8'b00000001; // 5944 :   1 - 0x1
      13'h1739: dout  = 8'b00000000; // 5945 :   0 - 0x0
      13'h173A: dout  = 8'b00000000; // 5946 :   0 - 0x0
      13'h173B: dout  = 8'b00000000; // 5947 :   0 - 0x0
      13'h173C: dout  = 8'b00000000; // 5948 :   0 - 0x0
      13'h173D: dout  = 8'b01000000; // 5949 :  64 - 0x40
      13'h173E: dout  = 8'b10000000; // 5950 : 128 - 0x80
      13'h173F: dout  = 8'b00000000; // 5951 :   0 - 0x0
      13'h1740: dout  = 8'b00000001; // 5952 :   1 - 0x1 -- Background 0x74
      13'h1741: dout  = 8'b00000001; // 5953 :   1 - 0x1
      13'h1742: dout  = 8'b00000001; // 5954 :   1 - 0x1
      13'h1743: dout  = 8'b00000001; // 5955 :   1 - 0x1
      13'h1744: dout  = 8'b00000001; // 5956 :   1 - 0x1
      13'h1745: dout  = 8'b00000001; // 5957 :   1 - 0x1
      13'h1746: dout  = 8'b00000001; // 5958 :   1 - 0x1
      13'h1747: dout  = 8'b00000001; // 5959 :   1 - 0x1
      13'h1748: dout  = 8'b00000001; // 5960 :   1 - 0x1
      13'h1749: dout  = 8'b00000001; // 5961 :   1 - 0x1
      13'h174A: dout  = 8'b00000001; // 5962 :   1 - 0x1
      13'h174B: dout  = 8'b00000001; // 5963 :   1 - 0x1
      13'h174C: dout  = 8'b00000001; // 5964 :   1 - 0x1
      13'h174D: dout  = 8'b00000001; // 5965 :   1 - 0x1
      13'h174E: dout  = 8'b00000001; // 5966 :   1 - 0x1
      13'h174F: dout  = 8'b00000001; // 5967 :   1 - 0x1
      13'h1750: dout  = 8'b10000000; // 5968 : 128 - 0x80 -- Background 0x75
      13'h1751: dout  = 8'b10000000; // 5969 : 128 - 0x80
      13'h1752: dout  = 8'b10000000; // 5970 : 128 - 0x80
      13'h1753: dout  = 8'b10000000; // 5971 : 128 - 0x80
      13'h1754: dout  = 8'b10000000; // 5972 : 128 - 0x80
      13'h1755: dout  = 8'b10000000; // 5973 : 128 - 0x80
      13'h1756: dout  = 8'b10000000; // 5974 : 128 - 0x80
      13'h1757: dout  = 8'b10000000; // 5975 : 128 - 0x80
      13'h1758: dout  = 8'b10000000; // 5976 : 128 - 0x80
      13'h1759: dout  = 8'b10000000; // 5977 : 128 - 0x80
      13'h175A: dout  = 8'b10000000; // 5978 : 128 - 0x80
      13'h175B: dout  = 8'b10000000; // 5979 : 128 - 0x80
      13'h175C: dout  = 8'b10000000; // 5980 : 128 - 0x80
      13'h175D: dout  = 8'b10000000; // 5981 : 128 - 0x80
      13'h175E: dout  = 8'b10000000; // 5982 : 128 - 0x80
      13'h175F: dout  = 8'b10000000; // 5983 : 128 - 0x80
      13'h1760: dout  = 8'b00000001; // 5984 :   1 - 0x1 -- Background 0x76
      13'h1761: dout  = 8'b00000011; // 5985 :   3 - 0x3
      13'h1762: dout  = 8'b00000000; // 5986 :   0 - 0x0
      13'h1763: dout  = 8'b00000000; // 5987 :   0 - 0x0
      13'h1764: dout  = 8'b00000011; // 5988 :   3 - 0x3
      13'h1765: dout  = 8'b00011001; // 5989 :  25 - 0x19
      13'h1766: dout  = 8'b00000000; // 5990 :   0 - 0x0
      13'h1767: dout  = 8'b00000000; // 5991 :   0 - 0x0
      13'h1768: dout  = 8'b00000001; // 5992 :   1 - 0x1
      13'h1769: dout  = 8'b00000011; // 5993 :   3 - 0x3
      13'h176A: dout  = 8'b00000011; // 5994 :   3 - 0x3
      13'h176B: dout  = 8'b00000111; // 5995 :   7 - 0x7
      13'h176C: dout  = 8'b00000100; // 5996 :   4 - 0x4
      13'h176D: dout  = 8'b00011100; // 5997 :  28 - 0x1c
      13'h176E: dout  = 8'b00111111; // 5998 :  63 - 0x3f
      13'h176F: dout  = 8'b01111111; // 5999 : 127 - 0x7f
      13'h1770: dout  = 8'b00000000; // 6000 :   0 - 0x0 -- Background 0x77
      13'h1771: dout  = 8'b00000000; // 6001 :   0 - 0x0
      13'h1772: dout  = 8'b01111100; // 6002 : 124 - 0x7c
      13'h1773: dout  = 8'b00000010; // 6003 :   2 - 0x2
      13'h1774: dout  = 8'b00000001; // 6004 :   1 - 0x1
      13'h1775: dout  = 8'b00000000; // 6005 :   0 - 0x0
      13'h1776: dout  = 8'b00000000; // 6006 :   0 - 0x0
      13'h1777: dout  = 8'b00000000; // 6007 :   0 - 0x0
      13'h1778: dout  = 8'b01111111; // 6008 : 127 - 0x7f
      13'h1779: dout  = 8'b11111111; // 6009 : 255 - 0xff
      13'h177A: dout  = 8'b11111111; // 6010 : 255 - 0xff
      13'h177B: dout  = 8'b01111111; // 6011 : 127 - 0x7f
      13'h177C: dout  = 8'b01111111; // 6012 : 127 - 0x7f
      13'h177D: dout  = 8'b00011111; // 6013 :  31 - 0x1f
      13'h177E: dout  = 8'b00000011; // 6014 :   3 - 0x3
      13'h177F: dout  = 8'b00000000; // 6015 :   0 - 0x0
      13'h1780: dout  = 8'b00000000; // 6016 :   0 - 0x0 -- Background 0x78
      13'h1781: dout  = 8'b00000000; // 6017 :   0 - 0x0
      13'h1782: dout  = 8'b00000001; // 6018 :   1 - 0x1
      13'h1783: dout  = 8'b00000001; // 6019 :   1 - 0x1
      13'h1784: dout  = 8'b00000011; // 6020 :   3 - 0x3
      13'h1785: dout  = 8'b00000111; // 6021 :   7 - 0x7
      13'h1786: dout  = 8'b00000111; // 6022 :   7 - 0x7
      13'h1787: dout  = 8'b00001111; // 6023 :  15 - 0xf
      13'h1788: dout  = 8'b00000000; // 6024 :   0 - 0x0
      13'h1789: dout  = 8'b00000000; // 6025 :   0 - 0x0
      13'h178A: dout  = 8'b00000001; // 6026 :   1 - 0x1
      13'h178B: dout  = 8'b00000001; // 6027 :   1 - 0x1
      13'h178C: dout  = 8'b00000011; // 6028 :   3 - 0x3
      13'h178D: dout  = 8'b00000111; // 6029 :   7 - 0x7
      13'h178E: dout  = 8'b00000111; // 6030 :   7 - 0x7
      13'h178F: dout  = 8'b00001111; // 6031 :  15 - 0xf
      13'h1790: dout  = 8'b00001111; // 6032 :  15 - 0xf -- Background 0x79
      13'h1791: dout  = 8'b00000111; // 6033 :   7 - 0x7
      13'h1792: dout  = 8'b00001111; // 6034 :  15 - 0xf
      13'h1793: dout  = 8'b00000111; // 6035 :   7 - 0x7
      13'h1794: dout  = 8'b00000001; // 6036 :   1 - 0x1
      13'h1795: dout  = 8'b00010000; // 6037 :  16 - 0x10
      13'h1796: dout  = 8'b00100000; // 6038 :  32 - 0x20
      13'h1797: dout  = 8'b00000000; // 6039 :   0 - 0x0
      13'h1798: dout  = 8'b11111111; // 6040 : 255 - 0xff
      13'h1799: dout  = 8'b11111111; // 6041 : 255 - 0xff
      13'h179A: dout  = 8'b00111111; // 6042 :  63 - 0x3f
      13'h179B: dout  = 8'b00111111; // 6043 :  63 - 0x3f
      13'h179C: dout  = 8'b01111111; // 6044 : 127 - 0x7f
      13'h179D: dout  = 8'b11111110; // 6045 : 254 - 0xfe
      13'h179E: dout  = 8'b11111100; // 6046 : 252 - 0xfc
      13'h179F: dout  = 8'b00110000; // 6047 :  48 - 0x30
      13'h17A0: dout  = 8'b11111000; // 6048 : 248 - 0xf8 -- Background 0x7a
      13'h17A1: dout  = 8'b11111110; // 6049 : 254 - 0xfe
      13'h17A2: dout  = 8'b01111111; // 6050 : 127 - 0x7f
      13'h17A3: dout  = 8'b00011111; // 6051 :  31 - 0x1f
      13'h17A4: dout  = 8'b00001111; // 6052 :  15 - 0xf
      13'h17A5: dout  = 8'b00011001; // 6053 :  25 - 0x19
      13'h17A6: dout  = 8'b00110000; // 6054 :  48 - 0x30
      13'h17A7: dout  = 8'b01110000; // 6055 : 112 - 0x70
      13'h17A8: dout  = 8'b11111000; // 6056 : 248 - 0xf8
      13'h17A9: dout  = 8'b11111110; // 6057 : 254 - 0xfe
      13'h17AA: dout  = 8'b11111111; // 6058 : 255 - 0xff
      13'h17AB: dout  = 8'b11111111; // 6059 : 255 - 0xff
      13'h17AC: dout  = 8'b11111111; // 6060 : 255 - 0xff
      13'h17AD: dout  = 8'b11111111; // 6061 : 255 - 0xff
      13'h17AE: dout  = 8'b11111111; // 6062 : 255 - 0xff
      13'h17AF: dout  = 8'b11111111; // 6063 : 255 - 0xff
      13'h17B0: dout  = 8'b11111011; // 6064 : 251 - 0xfb -- Background 0x7b
      13'h17B1: dout  = 8'b01110011; // 6065 : 115 - 0x73
      13'h17B2: dout  = 8'b00100111; // 6066 :  39 - 0x27
      13'h17B3: dout  = 8'b00001111; // 6067 :  15 - 0xf
      13'h17B4: dout  = 8'b00011111; // 6068 :  31 - 0x1f
      13'h17B5: dout  = 8'b00011111; // 6069 :  31 - 0x1f
      13'h17B6: dout  = 8'b00111111; // 6070 :  63 - 0x3f
      13'h17B7: dout  = 8'b01111111; // 6071 : 127 - 0x7f
      13'h17B8: dout  = 8'b11111111; // 6072 : 255 - 0xff
      13'h17B9: dout  = 8'b11111111; // 6073 : 255 - 0xff
      13'h17BA: dout  = 8'b11111111; // 6074 : 255 - 0xff
      13'h17BB: dout  = 8'b11111111; // 6075 : 255 - 0xff
      13'h17BC: dout  = 8'b11111111; // 6076 : 255 - 0xff
      13'h17BD: dout  = 8'b11111111; // 6077 : 255 - 0xff
      13'h17BE: dout  = 8'b11111111; // 6078 : 255 - 0xff
      13'h17BF: dout  = 8'b01111111; // 6079 : 127 - 0x7f
      13'h17C0: dout  = 8'b11111111; // 6080 : 255 - 0xff -- Background 0x7c
      13'h17C1: dout  = 8'b11111111; // 6081 : 255 - 0xff
      13'h17C2: dout  = 8'b11111111; // 6082 : 255 - 0xff
      13'h17C3: dout  = 8'b11111111; // 6083 : 255 - 0xff
      13'h17C4: dout  = 8'b11111110; // 6084 : 254 - 0xfe
      13'h17C5: dout  = 8'b11111101; // 6085 : 253 - 0xfd
      13'h17C6: dout  = 8'b11111000; // 6086 : 248 - 0xf8
      13'h17C7: dout  = 8'b11110110; // 6087 : 246 - 0xf6
      13'h17C8: dout  = 8'b11111111; // 6088 : 255 - 0xff
      13'h17C9: dout  = 8'b11111111; // 6089 : 255 - 0xff
      13'h17CA: dout  = 8'b11111111; // 6090 : 255 - 0xff
      13'h17CB: dout  = 8'b11111111; // 6091 : 255 - 0xff
      13'h17CC: dout  = 8'b11111111; // 6092 : 255 - 0xff
      13'h17CD: dout  = 8'b11111111; // 6093 : 255 - 0xff
      13'h17CE: dout  = 8'b11111111; // 6094 : 255 - 0xff
      13'h17CF: dout  = 8'b11111111; // 6095 : 255 - 0xff
      13'h17D0: dout  = 8'b11101111; // 6096 : 239 - 0xef -- Background 0x7d
      13'h17D1: dout  = 8'b11001111; // 6097 : 207 - 0xcf
      13'h17D2: dout  = 8'b10011111; // 6098 : 159 - 0x9f
      13'h17D3: dout  = 8'b00011111; // 6099 :  31 - 0x1f
      13'h17D4: dout  = 8'b00001111; // 6100 :  15 - 0xf
      13'h17D5: dout  = 8'b00101101; // 6101 :  45 - 0x2d
      13'h17D6: dout  = 8'b01010000; // 6102 :  80 - 0x50
      13'h17D7: dout  = 8'b01000000; // 6103 :  64 - 0x40
      13'h17D8: dout  = 8'b11101111; // 6104 : 239 - 0xef
      13'h17D9: dout  = 8'b11001111; // 6105 : 207 - 0xcf
      13'h17DA: dout  = 8'b10011111; // 6106 : 159 - 0x9f
      13'h17DB: dout  = 8'b00011111; // 6107 :  31 - 0x1f
      13'h17DC: dout  = 8'b00001111; // 6108 :  15 - 0xf
      13'h17DD: dout  = 8'b01111111; // 6109 : 127 - 0x7f
      13'h17DE: dout  = 8'b11111111; // 6110 : 255 - 0xff
      13'h17DF: dout  = 8'b11111111; // 6111 : 255 - 0xff
      13'h17E0: dout  = 8'b00000000; // 6112 :   0 - 0x0 -- Background 0x7e
      13'h17E1: dout  = 8'b00000000; // 6113 :   0 - 0x0
      13'h17E2: dout  = 8'b00000000; // 6114 :   0 - 0x0
      13'h17E3: dout  = 8'b00000000; // 6115 :   0 - 0x0
      13'h17E4: dout  = 8'b11100000; // 6116 : 224 - 0xe0
      13'h17E5: dout  = 8'b11111110; // 6117 : 254 - 0xfe
      13'h17E6: dout  = 8'b11111111; // 6118 : 255 - 0xff
      13'h17E7: dout  = 8'b11110011; // 6119 : 243 - 0xf3
      13'h17E8: dout  = 8'b00000000; // 6120 :   0 - 0x0
      13'h17E9: dout  = 8'b00000000; // 6121 :   0 - 0x0
      13'h17EA: dout  = 8'b00000000; // 6122 :   0 - 0x0
      13'h17EB: dout  = 8'b11110000; // 6123 : 240 - 0xf0
      13'h17EC: dout  = 8'b11111110; // 6124 : 254 - 0xfe
      13'h17ED: dout  = 8'b11111111; // 6125 : 255 - 0xff
      13'h17EE: dout  = 8'b11111111; // 6126 : 255 - 0xff
      13'h17EF: dout  = 8'b11111111; // 6127 : 255 - 0xff
      13'h17F0: dout  = 8'b11111011; // 6128 : 251 - 0xfb -- Background 0x7f
      13'h17F1: dout  = 8'b11111011; // 6129 : 251 - 0xfb
      13'h17F2: dout  = 8'b11111011; // 6130 : 251 - 0xfb
      13'h17F3: dout  = 8'b11111011; // 6131 : 251 - 0xfb
      13'h17F4: dout  = 8'b11111011; // 6132 : 251 - 0xfb
      13'h17F5: dout  = 8'b11110011; // 6133 : 243 - 0xf3
      13'h17F6: dout  = 8'b11110111; // 6134 : 247 - 0xf7
      13'h17F7: dout  = 8'b11100111; // 6135 : 231 - 0xe7
      13'h17F8: dout  = 8'b11111111; // 6136 : 255 - 0xff
      13'h17F9: dout  = 8'b11111111; // 6137 : 255 - 0xff
      13'h17FA: dout  = 8'b11111111; // 6138 : 255 - 0xff
      13'h17FB: dout  = 8'b11111111; // 6139 : 255 - 0xff
      13'h17FC: dout  = 8'b11111111; // 6140 : 255 - 0xff
      13'h17FD: dout  = 8'b11111111; // 6141 : 255 - 0xff
      13'h17FE: dout  = 8'b11111111; // 6142 : 255 - 0xff
      13'h17FF: dout  = 8'b11111111; // 6143 : 255 - 0xff
      13'h1800: dout  = 8'b11001111; // 6144 : 207 - 0xcf -- Background 0x80
      13'h1801: dout  = 8'b10011111; // 6145 : 159 - 0x9f
      13'h1802: dout  = 8'b00111111; // 6146 :  63 - 0x3f
      13'h1803: dout  = 8'b00111111; // 6147 :  63 - 0x3f
      13'h1804: dout  = 8'b00111111; // 6148 :  63 - 0x3f
      13'h1805: dout  = 8'b00001111; // 6149 :  15 - 0xf
      13'h1806: dout  = 8'b00000011; // 6150 :   3 - 0x3
      13'h1807: dout  = 8'b00000000; // 6151 :   0 - 0x0
      13'h1808: dout  = 8'b11111111; // 6152 : 255 - 0xff
      13'h1809: dout  = 8'b11111111; // 6153 : 255 - 0xff
      13'h180A: dout  = 8'b11111111; // 6154 : 255 - 0xff
      13'h180B: dout  = 8'b11111111; // 6155 : 255 - 0xff
      13'h180C: dout  = 8'b11111111; // 6156 : 255 - 0xff
      13'h180D: dout  = 8'b11111111; // 6157 : 255 - 0xff
      13'h180E: dout  = 8'b11111111; // 6158 : 255 - 0xff
      13'h180F: dout  = 8'b11111111; // 6159 : 255 - 0xff
      13'h1810: dout  = 8'b11000000; // 6160 : 192 - 0xc0 -- Background 0x81
      13'h1811: dout  = 8'b11110000; // 6161 : 240 - 0xf0
      13'h1812: dout  = 8'b11111100; // 6162 : 252 - 0xfc
      13'h1813: dout  = 8'b11110000; // 6163 : 240 - 0xf0
      13'h1814: dout  = 8'b11110000; // 6164 : 240 - 0xf0
      13'h1815: dout  = 8'b10011000; // 6165 : 152 - 0x98
      13'h1816: dout  = 8'b00001000; // 6166 :   8 - 0x8
      13'h1817: dout  = 8'b00000000; // 6167 :   0 - 0x0
      13'h1818: dout  = 8'b11111111; // 6168 : 255 - 0xff
      13'h1819: dout  = 8'b11111111; // 6169 : 255 - 0xff
      13'h181A: dout  = 8'b11111111; // 6170 : 255 - 0xff
      13'h181B: dout  = 8'b11110000; // 6171 : 240 - 0xf0
      13'h181C: dout  = 8'b11110000; // 6172 : 240 - 0xf0
      13'h181D: dout  = 8'b11111000; // 6173 : 248 - 0xf8
      13'h181E: dout  = 8'b11111000; // 6174 : 248 - 0xf8
      13'h181F: dout  = 8'b11111000; // 6175 : 248 - 0xf8
      13'h1820: dout  = 8'b00000000; // 6176 :   0 - 0x0 -- Background 0x82
      13'h1821: dout  = 8'b00000000; // 6177 :   0 - 0x0
      13'h1822: dout  = 8'b00000000; // 6178 :   0 - 0x0
      13'h1823: dout  = 8'b00000000; // 6179 :   0 - 0x0
      13'h1824: dout  = 8'b00000000; // 6180 :   0 - 0x0
      13'h1825: dout  = 8'b00000000; // 6181 :   0 - 0x0
      13'h1826: dout  = 8'b10000000; // 6182 : 128 - 0x80
      13'h1827: dout  = 8'b11000000; // 6183 : 192 - 0xc0
      13'h1828: dout  = 8'b00000000; // 6184 :   0 - 0x0
      13'h1829: dout  = 8'b00000000; // 6185 :   0 - 0x0
      13'h182A: dout  = 8'b00000000; // 6186 :   0 - 0x0
      13'h182B: dout  = 8'b00000000; // 6187 :   0 - 0x0
      13'h182C: dout  = 8'b00000000; // 6188 :   0 - 0x0
      13'h182D: dout  = 8'b10000000; // 6189 : 128 - 0x80
      13'h182E: dout  = 8'b11000000; // 6190 : 192 - 0xc0
      13'h182F: dout  = 8'b11100000; // 6191 : 224 - 0xe0
      13'h1830: dout  = 8'b11100000; // 6192 : 224 - 0xe0 -- Background 0x83
      13'h1831: dout  = 8'b11100000; // 6193 : 224 - 0xe0
      13'h1832: dout  = 8'b11110000; // 6194 : 240 - 0xf0
      13'h1833: dout  = 8'b11110000; // 6195 : 240 - 0xf0
      13'h1834: dout  = 8'b11110000; // 6196 : 240 - 0xf0
      13'h1835: dout  = 8'b11110000; // 6197 : 240 - 0xf0
      13'h1836: dout  = 8'b11111000; // 6198 : 248 - 0xf8
      13'h1837: dout  = 8'b11111000; // 6199 : 248 - 0xf8
      13'h1838: dout  = 8'b11110000; // 6200 : 240 - 0xf0
      13'h1839: dout  = 8'b11110000; // 6201 : 240 - 0xf0
      13'h183A: dout  = 8'b11111000; // 6202 : 248 - 0xf8
      13'h183B: dout  = 8'b11111000; // 6203 : 248 - 0xf8
      13'h183C: dout  = 8'b11111000; // 6204 : 248 - 0xf8
      13'h183D: dout  = 8'b11111100; // 6205 : 252 - 0xfc
      13'h183E: dout  = 8'b11111100; // 6206 : 252 - 0xfc
      13'h183F: dout  = 8'b11111110; // 6207 : 254 - 0xfe
      13'h1840: dout  = 8'b11111110; // 6208 : 254 - 0xfe -- Background 0x84
      13'h1841: dout  = 8'b11111111; // 6209 : 255 - 0xff
      13'h1842: dout  = 8'b11111111; // 6210 : 255 - 0xff
      13'h1843: dout  = 8'b11111111; // 6211 : 255 - 0xff
      13'h1844: dout  = 8'b11111111; // 6212 : 255 - 0xff
      13'h1845: dout  = 8'b11111111; // 6213 : 255 - 0xff
      13'h1846: dout  = 8'b11111111; // 6214 : 255 - 0xff
      13'h1847: dout  = 8'b11111111; // 6215 : 255 - 0xff
      13'h1848: dout  = 8'b11111111; // 6216 : 255 - 0xff
      13'h1849: dout  = 8'b11111111; // 6217 : 255 - 0xff
      13'h184A: dout  = 8'b11111111; // 6218 : 255 - 0xff
      13'h184B: dout  = 8'b11111111; // 6219 : 255 - 0xff
      13'h184C: dout  = 8'b11111111; // 6220 : 255 - 0xff
      13'h184D: dout  = 8'b11111111; // 6221 : 255 - 0xff
      13'h184E: dout  = 8'b11111111; // 6222 : 255 - 0xff
      13'h184F: dout  = 8'b11111111; // 6223 : 255 - 0xff
      13'h1850: dout  = 8'b00111111; // 6224 :  63 - 0x3f -- Background 0x85
      13'h1851: dout  = 8'b00011111; // 6225 :  31 - 0x1f
      13'h1852: dout  = 8'b00011111; // 6226 :  31 - 0x1f
      13'h1853: dout  = 8'b00001111; // 6227 :  15 - 0xf
      13'h1854: dout  = 8'b00000111; // 6228 :   7 - 0x7
      13'h1855: dout  = 8'b00000000; // 6229 :   0 - 0x0
      13'h1856: dout  = 8'b00000000; // 6230 :   0 - 0x0
      13'h1857: dout  = 8'b00000000; // 6231 :   0 - 0x0
      13'h1858: dout  = 8'b11111111; // 6232 : 255 - 0xff
      13'h1859: dout  = 8'b11111111; // 6233 : 255 - 0xff
      13'h185A: dout  = 8'b11111111; // 6234 : 255 - 0xff
      13'h185B: dout  = 8'b00001111; // 6235 :  15 - 0xf
      13'h185C: dout  = 8'b00000111; // 6236 :   7 - 0x7
      13'h185D: dout  = 8'b00000000; // 6237 :   0 - 0x0
      13'h185E: dout  = 8'b00000000; // 6238 :   0 - 0x0
      13'h185F: dout  = 8'b00000000; // 6239 :   0 - 0x0
      13'h1860: dout  = 8'b00000000; // 6240 :   0 - 0x0 -- Background 0x86
      13'h1861: dout  = 8'b00000000; // 6241 :   0 - 0x0
      13'h1862: dout  = 8'b11000000; // 6242 : 192 - 0xc0
      13'h1863: dout  = 8'b11100000; // 6243 : 224 - 0xe0
      13'h1864: dout  = 8'b11110000; // 6244 : 240 - 0xf0
      13'h1865: dout  = 8'b11110000; // 6245 : 240 - 0xf0
      13'h1866: dout  = 8'b11110000; // 6246 : 240 - 0xf0
      13'h1867: dout  = 8'b11111000; // 6247 : 248 - 0xf8
      13'h1868: dout  = 8'b00000000; // 6248 :   0 - 0x0
      13'h1869: dout  = 8'b10000000; // 6249 : 128 - 0x80
      13'h186A: dout  = 8'b11000000; // 6250 : 192 - 0xc0
      13'h186B: dout  = 8'b11100000; // 6251 : 224 - 0xe0
      13'h186C: dout  = 8'b11110000; // 6252 : 240 - 0xf0
      13'h186D: dout  = 8'b11110000; // 6253 : 240 - 0xf0
      13'h186E: dout  = 8'b11110000; // 6254 : 240 - 0xf0
      13'h186F: dout  = 8'b11111100; // 6255 : 252 - 0xfc
      13'h1870: dout  = 8'b11111001; // 6256 : 249 - 0xf9 -- Background 0x87
      13'h1871: dout  = 8'b11111111; // 6257 : 255 - 0xff
      13'h1872: dout  = 8'b11111111; // 6258 : 255 - 0xff
      13'h1873: dout  = 8'b11111111; // 6259 : 255 - 0xff
      13'h1874: dout  = 8'b11111111; // 6260 : 255 - 0xff
      13'h1875: dout  = 8'b00001110; // 6261 :  14 - 0xe
      13'h1876: dout  = 8'b00000010; // 6262 :   2 - 0x2
      13'h1877: dout  = 8'b00010100; // 6263 :  20 - 0x14
      13'h1878: dout  = 8'b11111111; // 6264 : 255 - 0xff
      13'h1879: dout  = 8'b11111111; // 6265 : 255 - 0xff
      13'h187A: dout  = 8'b11111111; // 6266 : 255 - 0xff
      13'h187B: dout  = 8'b11111111; // 6267 : 255 - 0xff
      13'h187C: dout  = 8'b11111111; // 6268 : 255 - 0xff
      13'h187D: dout  = 8'b00001111; // 6269 :  15 - 0xf
      13'h187E: dout  = 8'b00011111; // 6270 :  31 - 0x1f
      13'h187F: dout  = 8'b00111111; // 6271 :  63 - 0x3f
      13'h1880: dout  = 8'b10000000; // 6272 : 128 - 0x80 -- Background 0x88
      13'h1881: dout  = 8'b10100000; // 6273 : 160 - 0xa0
      13'h1882: dout  = 8'b00100000; // 6274 :  32 - 0x20
      13'h1883: dout  = 8'b00100000; // 6275 :  32 - 0x20
      13'h1884: dout  = 8'b10100000; // 6276 : 160 - 0xa0
      13'h1885: dout  = 8'b10000000; // 6277 : 128 - 0x80
      13'h1886: dout  = 8'b00000000; // 6278 :   0 - 0x0
      13'h1887: dout  = 8'b00000000; // 6279 :   0 - 0x0
      13'h1888: dout  = 8'b11000000; // 6280 : 192 - 0xc0
      13'h1889: dout  = 8'b11100000; // 6281 : 224 - 0xe0
      13'h188A: dout  = 8'b11100000; // 6282 : 224 - 0xe0
      13'h188B: dout  = 8'b11100000; // 6283 : 224 - 0xe0
      13'h188C: dout  = 8'b11100000; // 6284 : 224 - 0xe0
      13'h188D: dout  = 8'b11000000; // 6285 : 192 - 0xc0
      13'h188E: dout  = 8'b11000000; // 6286 : 192 - 0xc0
      13'h188F: dout  = 8'b10000000; // 6287 : 128 - 0x80
      13'h1890: dout  = 8'b00000001; // 6288 :   1 - 0x1 -- Background 0x89
      13'h1891: dout  = 8'b00000101; // 6289 :   5 - 0x5
      13'h1892: dout  = 8'b00000100; // 6290 :   4 - 0x4
      13'h1893: dout  = 8'b00000100; // 6291 :   4 - 0x4
      13'h1894: dout  = 8'b00000101; // 6292 :   5 - 0x5
      13'h1895: dout  = 8'b00000001; // 6293 :   1 - 0x1
      13'h1896: dout  = 8'b00000000; // 6294 :   0 - 0x0
      13'h1897: dout  = 8'b00000000; // 6295 :   0 - 0x0
      13'h1898: dout  = 8'b00000011; // 6296 :   3 - 0x3
      13'h1899: dout  = 8'b00000111; // 6297 :   7 - 0x7
      13'h189A: dout  = 8'b00000111; // 6298 :   7 - 0x7
      13'h189B: dout  = 8'b00000111; // 6299 :   7 - 0x7
      13'h189C: dout  = 8'b00000111; // 6300 :   7 - 0x7
      13'h189D: dout  = 8'b00000011; // 6301 :   3 - 0x3
      13'h189E: dout  = 8'b00000011; // 6302 :   3 - 0x3
      13'h189F: dout  = 8'b00000001; // 6303 :   1 - 0x1
      13'h18A0: dout  = 8'b00000000; // 6304 :   0 - 0x0 -- Background 0x8a
      13'h18A1: dout  = 8'b00000000; // 6305 :   0 - 0x0
      13'h18A2: dout  = 8'b00000011; // 6306 :   3 - 0x3
      13'h18A3: dout  = 8'b00000111; // 6307 :   7 - 0x7
      13'h18A4: dout  = 8'b00001111; // 6308 :  15 - 0xf
      13'h18A5: dout  = 8'b00001111; // 6309 :  15 - 0xf
      13'h18A6: dout  = 8'b00001111; // 6310 :  15 - 0xf
      13'h18A7: dout  = 8'b00001111; // 6311 :  15 - 0xf
      13'h18A8: dout  = 8'b00000000; // 6312 :   0 - 0x0
      13'h18A9: dout  = 8'b00000001; // 6313 :   1 - 0x1
      13'h18AA: dout  = 8'b00000011; // 6314 :   3 - 0x3
      13'h18AB: dout  = 8'b00000111; // 6315 :   7 - 0x7
      13'h18AC: dout  = 8'b00001111; // 6316 :  15 - 0xf
      13'h18AD: dout  = 8'b00001111; // 6317 :  15 - 0xf
      13'h18AE: dout  = 8'b00001111; // 6318 :  15 - 0xf
      13'h18AF: dout  = 8'b00111111; // 6319 :  63 - 0x3f
      13'h18B0: dout  = 8'b10011111; // 6320 : 159 - 0x9f -- Background 0x8b
      13'h18B1: dout  = 8'b11111111; // 6321 : 255 - 0xff
      13'h18B2: dout  = 8'b11111111; // 6322 : 255 - 0xff
      13'h18B3: dout  = 8'b11111111; // 6323 : 255 - 0xff
      13'h18B4: dout  = 8'b11111111; // 6324 : 255 - 0xff
      13'h18B5: dout  = 8'b01110000; // 6325 : 112 - 0x70
      13'h18B6: dout  = 8'b01000000; // 6326 :  64 - 0x40
      13'h18B7: dout  = 8'b00101000; // 6327 :  40 - 0x28
      13'h18B8: dout  = 8'b11111111; // 6328 : 255 - 0xff
      13'h18B9: dout  = 8'b11111111; // 6329 : 255 - 0xff
      13'h18BA: dout  = 8'b11111111; // 6330 : 255 - 0xff
      13'h18BB: dout  = 8'b11111111; // 6331 : 255 - 0xff
      13'h18BC: dout  = 8'b11111111; // 6332 : 255 - 0xff
      13'h18BD: dout  = 8'b11110000; // 6333 : 240 - 0xf0
      13'h18BE: dout  = 8'b11111000; // 6334 : 248 - 0xf8
      13'h18BF: dout  = 8'b11111100; // 6335 : 252 - 0xfc
      13'h18C0: dout  = 8'b00000000; // 6336 :   0 - 0x0 -- Background 0x8c
      13'h18C1: dout  = 8'b00000000; // 6337 :   0 - 0x0
      13'h18C2: dout  = 8'b00000000; // 6338 :   0 - 0x0
      13'h18C3: dout  = 8'b00000000; // 6339 :   0 - 0x0
      13'h18C4: dout  = 8'b00000000; // 6340 :   0 - 0x0
      13'h18C5: dout  = 8'b00000000; // 6341 :   0 - 0x0
      13'h18C6: dout  = 8'b00000001; // 6342 :   1 - 0x1
      13'h18C7: dout  = 8'b00000011; // 6343 :   3 - 0x3
      13'h18C8: dout  = 8'b00000000; // 6344 :   0 - 0x0
      13'h18C9: dout  = 8'b00000000; // 6345 :   0 - 0x0
      13'h18CA: dout  = 8'b00000000; // 6346 :   0 - 0x0
      13'h18CB: dout  = 8'b00000000; // 6347 :   0 - 0x0
      13'h18CC: dout  = 8'b00000000; // 6348 :   0 - 0x0
      13'h18CD: dout  = 8'b00000001; // 6349 :   1 - 0x1
      13'h18CE: dout  = 8'b00000011; // 6350 :   3 - 0x3
      13'h18CF: dout  = 8'b00000111; // 6351 :   7 - 0x7
      13'h18D0: dout  = 8'b00000111; // 6352 :   7 - 0x7 -- Background 0x8d
      13'h18D1: dout  = 8'b00000111; // 6353 :   7 - 0x7
      13'h18D2: dout  = 8'b00001111; // 6354 :  15 - 0xf
      13'h18D3: dout  = 8'b00001111; // 6355 :  15 - 0xf
      13'h18D4: dout  = 8'b00001111; // 6356 :  15 - 0xf
      13'h18D5: dout  = 8'b00001111; // 6357 :  15 - 0xf
      13'h18D6: dout  = 8'b00011111; // 6358 :  31 - 0x1f
      13'h18D7: dout  = 8'b00011111; // 6359 :  31 - 0x1f
      13'h18D8: dout  = 8'b00001111; // 6360 :  15 - 0xf
      13'h18D9: dout  = 8'b00001111; // 6361 :  15 - 0xf
      13'h18DA: dout  = 8'b00011111; // 6362 :  31 - 0x1f
      13'h18DB: dout  = 8'b00011111; // 6363 :  31 - 0x1f
      13'h18DC: dout  = 8'b00011111; // 6364 :  31 - 0x1f
      13'h18DD: dout  = 8'b00111111; // 6365 :  63 - 0x3f
      13'h18DE: dout  = 8'b00111111; // 6366 :  63 - 0x3f
      13'h18DF: dout  = 8'b01111111; // 6367 : 127 - 0x7f
      13'h18E0: dout  = 8'b01111111; // 6368 : 127 - 0x7f -- Background 0x8e
      13'h18E1: dout  = 8'b11111111; // 6369 : 255 - 0xff
      13'h18E2: dout  = 8'b11111111; // 6370 : 255 - 0xff
      13'h18E3: dout  = 8'b11111111; // 6371 : 255 - 0xff
      13'h18E4: dout  = 8'b11111111; // 6372 : 255 - 0xff
      13'h18E5: dout  = 8'b11111111; // 6373 : 255 - 0xff
      13'h18E6: dout  = 8'b11111111; // 6374 : 255 - 0xff
      13'h18E7: dout  = 8'b11111111; // 6375 : 255 - 0xff
      13'h18E8: dout  = 8'b11111111; // 6376 : 255 - 0xff
      13'h18E9: dout  = 8'b11111111; // 6377 : 255 - 0xff
      13'h18EA: dout  = 8'b11111111; // 6378 : 255 - 0xff
      13'h18EB: dout  = 8'b11111111; // 6379 : 255 - 0xff
      13'h18EC: dout  = 8'b11111111; // 6380 : 255 - 0xff
      13'h18ED: dout  = 8'b11111111; // 6381 : 255 - 0xff
      13'h18EE: dout  = 8'b11111111; // 6382 : 255 - 0xff
      13'h18EF: dout  = 8'b11111111; // 6383 : 255 - 0xff
      13'h18F0: dout  = 8'b11111100; // 6384 : 252 - 0xfc -- Background 0x8f
      13'h18F1: dout  = 8'b11111000; // 6385 : 248 - 0xf8
      13'h18F2: dout  = 8'b11111000; // 6386 : 248 - 0xf8
      13'h18F3: dout  = 8'b11110000; // 6387 : 240 - 0xf0
      13'h18F4: dout  = 8'b11100000; // 6388 : 224 - 0xe0
      13'h18F5: dout  = 8'b00000000; // 6389 :   0 - 0x0
      13'h18F6: dout  = 8'b00000000; // 6390 :   0 - 0x0
      13'h18F7: dout  = 8'b00000000; // 6391 :   0 - 0x0
      13'h18F8: dout  = 8'b11111111; // 6392 : 255 - 0xff
      13'h18F9: dout  = 8'b11111111; // 6393 : 255 - 0xff
      13'h18FA: dout  = 8'b11111111; // 6394 : 255 - 0xff
      13'h18FB: dout  = 8'b11110000; // 6395 : 240 - 0xf0
      13'h18FC: dout  = 8'b11100000; // 6396 : 224 - 0xe0
      13'h18FD: dout  = 8'b00000000; // 6397 :   0 - 0x0
      13'h18FE: dout  = 8'b00000000; // 6398 :   0 - 0x0
      13'h18FF: dout  = 8'b00000000; // 6399 :   0 - 0x0
      13'h1900: dout  = 8'b00000000; // 6400 :   0 - 0x0 -- Background 0x90
      13'h1901: dout  = 8'b00000000; // 6401 :   0 - 0x0
      13'h1902: dout  = 8'b00000000; // 6402 :   0 - 0x0
      13'h1903: dout  = 8'b00000000; // 6403 :   0 - 0x0
      13'h1904: dout  = 8'b00000111; // 6404 :   7 - 0x7
      13'h1905: dout  = 8'b01111111; // 6405 : 127 - 0x7f
      13'h1906: dout  = 8'b11111111; // 6406 : 255 - 0xff
      13'h1907: dout  = 8'b11001111; // 6407 : 207 - 0xcf
      13'h1908: dout  = 8'b00000000; // 6408 :   0 - 0x0
      13'h1909: dout  = 8'b00000000; // 6409 :   0 - 0x0
      13'h190A: dout  = 8'b00000000; // 6410 :   0 - 0x0
      13'h190B: dout  = 8'b00001111; // 6411 :  15 - 0xf
      13'h190C: dout  = 8'b01111111; // 6412 : 127 - 0x7f
      13'h190D: dout  = 8'b11111111; // 6413 : 255 - 0xff
      13'h190E: dout  = 8'b11111111; // 6414 : 255 - 0xff
      13'h190F: dout  = 8'b11111111; // 6415 : 255 - 0xff
      13'h1910: dout  = 8'b11011111; // 6416 : 223 - 0xdf -- Background 0x91
      13'h1911: dout  = 8'b11011111; // 6417 : 223 - 0xdf
      13'h1912: dout  = 8'b11011111; // 6418 : 223 - 0xdf
      13'h1913: dout  = 8'b11011111; // 6419 : 223 - 0xdf
      13'h1914: dout  = 8'b11011111; // 6420 : 223 - 0xdf
      13'h1915: dout  = 8'b11001111; // 6421 : 207 - 0xcf
      13'h1916: dout  = 8'b11101111; // 6422 : 239 - 0xef
      13'h1917: dout  = 8'b11100111; // 6423 : 231 - 0xe7
      13'h1918: dout  = 8'b11111111; // 6424 : 255 - 0xff
      13'h1919: dout  = 8'b11111111; // 6425 : 255 - 0xff
      13'h191A: dout  = 8'b11111111; // 6426 : 255 - 0xff
      13'h191B: dout  = 8'b11111111; // 6427 : 255 - 0xff
      13'h191C: dout  = 8'b11111111; // 6428 : 255 - 0xff
      13'h191D: dout  = 8'b11111111; // 6429 : 255 - 0xff
      13'h191E: dout  = 8'b11111111; // 6430 : 255 - 0xff
      13'h191F: dout  = 8'b11111111; // 6431 : 255 - 0xff
      13'h1920: dout  = 8'b11110011; // 6432 : 243 - 0xf3 -- Background 0x92
      13'h1921: dout  = 8'b11111001; // 6433 : 249 - 0xf9
      13'h1922: dout  = 8'b11111100; // 6434 : 252 - 0xfc
      13'h1923: dout  = 8'b11111100; // 6435 : 252 - 0xfc
      13'h1924: dout  = 8'b11111100; // 6436 : 252 - 0xfc
      13'h1925: dout  = 8'b11110000; // 6437 : 240 - 0xf0
      13'h1926: dout  = 8'b11000000; // 6438 : 192 - 0xc0
      13'h1927: dout  = 8'b00000000; // 6439 :   0 - 0x0
      13'h1928: dout  = 8'b11111111; // 6440 : 255 - 0xff
      13'h1929: dout  = 8'b11111111; // 6441 : 255 - 0xff
      13'h192A: dout  = 8'b11111111; // 6442 : 255 - 0xff
      13'h192B: dout  = 8'b11111111; // 6443 : 255 - 0xff
      13'h192C: dout  = 8'b11111111; // 6444 : 255 - 0xff
      13'h192D: dout  = 8'b11111111; // 6445 : 255 - 0xff
      13'h192E: dout  = 8'b11111111; // 6446 : 255 - 0xff
      13'h192F: dout  = 8'b11111111; // 6447 : 255 - 0xff
      13'h1930: dout  = 8'b00000011; // 6448 :   3 - 0x3 -- Background 0x93
      13'h1931: dout  = 8'b00001111; // 6449 :  15 - 0xf
      13'h1932: dout  = 8'b00111111; // 6450 :  63 - 0x3f
      13'h1933: dout  = 8'b00001111; // 6451 :  15 - 0xf
      13'h1934: dout  = 8'b00001111; // 6452 :  15 - 0xf
      13'h1935: dout  = 8'b00011001; // 6453 :  25 - 0x19
      13'h1936: dout  = 8'b00010000; // 6454 :  16 - 0x10
      13'h1937: dout  = 8'b00000000; // 6455 :   0 - 0x0
      13'h1938: dout  = 8'b11111111; // 6456 : 255 - 0xff
      13'h1939: dout  = 8'b11111111; // 6457 : 255 - 0xff
      13'h193A: dout  = 8'b11111111; // 6458 : 255 - 0xff
      13'h193B: dout  = 8'b00001111; // 6459 :  15 - 0xf
      13'h193C: dout  = 8'b00001111; // 6460 :  15 - 0xf
      13'h193D: dout  = 8'b00011111; // 6461 :  31 - 0x1f
      13'h193E: dout  = 8'b00011111; // 6462 :  31 - 0x1f
      13'h193F: dout  = 8'b00011111; // 6463 :  31 - 0x1f
      13'h1940: dout  = 8'b00011111; // 6464 :  31 - 0x1f -- Background 0x94
      13'h1941: dout  = 8'b01111111; // 6465 : 127 - 0x7f
      13'h1942: dout  = 8'b11111110; // 6466 : 254 - 0xfe
      13'h1943: dout  = 8'b11111000; // 6467 : 248 - 0xf8
      13'h1944: dout  = 8'b11110000; // 6468 : 240 - 0xf0
      13'h1945: dout  = 8'b10011000; // 6469 : 152 - 0x98
      13'h1946: dout  = 8'b00001100; // 6470 :  12 - 0xc
      13'h1947: dout  = 8'b00001110; // 6471 :  14 - 0xe
      13'h1948: dout  = 8'b00011111; // 6472 :  31 - 0x1f
      13'h1949: dout  = 8'b01111111; // 6473 : 127 - 0x7f
      13'h194A: dout  = 8'b11111111; // 6474 : 255 - 0xff
      13'h194B: dout  = 8'b11111111; // 6475 : 255 - 0xff
      13'h194C: dout  = 8'b11111111; // 6476 : 255 - 0xff
      13'h194D: dout  = 8'b11111111; // 6477 : 255 - 0xff
      13'h194E: dout  = 8'b11111111; // 6478 : 255 - 0xff
      13'h194F: dout  = 8'b11111111; // 6479 : 255 - 0xff
      13'h1950: dout  = 8'b11011111; // 6480 : 223 - 0xdf -- Background 0x95
      13'h1951: dout  = 8'b11001110; // 6481 : 206 - 0xce
      13'h1952: dout  = 8'b11100100; // 6482 : 228 - 0xe4
      13'h1953: dout  = 8'b11110000; // 6483 : 240 - 0xf0
      13'h1954: dout  = 8'b11111000; // 6484 : 248 - 0xf8
      13'h1955: dout  = 8'b11111000; // 6485 : 248 - 0xf8
      13'h1956: dout  = 8'b11111100; // 6486 : 252 - 0xfc
      13'h1957: dout  = 8'b11111110; // 6487 : 254 - 0xfe
      13'h1958: dout  = 8'b11111111; // 6488 : 255 - 0xff
      13'h1959: dout  = 8'b11111111; // 6489 : 255 - 0xff
      13'h195A: dout  = 8'b11111111; // 6490 : 255 - 0xff
      13'h195B: dout  = 8'b11111111; // 6491 : 255 - 0xff
      13'h195C: dout  = 8'b11111111; // 6492 : 255 - 0xff
      13'h195D: dout  = 8'b11111111; // 6493 : 255 - 0xff
      13'h195E: dout  = 8'b11111111; // 6494 : 255 - 0xff
      13'h195F: dout  = 8'b11111110; // 6495 : 254 - 0xfe
      13'h1960: dout  = 8'b11111111; // 6496 : 255 - 0xff -- Background 0x96
      13'h1961: dout  = 8'b11111111; // 6497 : 255 - 0xff
      13'h1962: dout  = 8'b11111111; // 6498 : 255 - 0xff
      13'h1963: dout  = 8'b11111111; // 6499 : 255 - 0xff
      13'h1964: dout  = 8'b01111111; // 6500 : 127 - 0x7f
      13'h1965: dout  = 8'b10111111; // 6501 : 191 - 0xbf
      13'h1966: dout  = 8'b00011111; // 6502 :  31 - 0x1f
      13'h1967: dout  = 8'b01101111; // 6503 : 111 - 0x6f
      13'h1968: dout  = 8'b11111111; // 6504 : 255 - 0xff
      13'h1969: dout  = 8'b11111111; // 6505 : 255 - 0xff
      13'h196A: dout  = 8'b11111111; // 6506 : 255 - 0xff
      13'h196B: dout  = 8'b11111111; // 6507 : 255 - 0xff
      13'h196C: dout  = 8'b11111111; // 6508 : 255 - 0xff
      13'h196D: dout  = 8'b11111111; // 6509 : 255 - 0xff
      13'h196E: dout  = 8'b11111111; // 6510 : 255 - 0xff
      13'h196F: dout  = 8'b11111111; // 6511 : 255 - 0xff
      13'h1970: dout  = 8'b11110111; // 6512 : 247 - 0xf7 -- Background 0x97
      13'h1971: dout  = 8'b11110011; // 6513 : 243 - 0xf3
      13'h1972: dout  = 8'b11111001; // 6514 : 249 - 0xf9
      13'h1973: dout  = 8'b11111000; // 6515 : 248 - 0xf8
      13'h1974: dout  = 8'b11110000; // 6516 : 240 - 0xf0
      13'h1975: dout  = 8'b10110100; // 6517 : 180 - 0xb4
      13'h1976: dout  = 8'b00001010; // 6518 :  10 - 0xa
      13'h1977: dout  = 8'b00000010; // 6519 :   2 - 0x2
      13'h1978: dout  = 8'b11110111; // 6520 : 247 - 0xf7
      13'h1979: dout  = 8'b11110011; // 6521 : 243 - 0xf3
      13'h197A: dout  = 8'b11111001; // 6522 : 249 - 0xf9
      13'h197B: dout  = 8'b11111000; // 6523 : 248 - 0xf8
      13'h197C: dout  = 8'b11110000; // 6524 : 240 - 0xf0
      13'h197D: dout  = 8'b11111110; // 6525 : 254 - 0xfe
      13'h197E: dout  = 8'b11111111; // 6526 : 255 - 0xff
      13'h197F: dout  = 8'b11111111; // 6527 : 255 - 0xff
      13'h1980: dout  = 8'b10000000; // 6528 : 128 - 0x80 -- Background 0x98
      13'h1981: dout  = 8'b11000000; // 6529 : 192 - 0xc0
      13'h1982: dout  = 8'b00000000; // 6530 :   0 - 0x0
      13'h1983: dout  = 8'b00000000; // 6531 :   0 - 0x0
      13'h1984: dout  = 8'b11000000; // 6532 : 192 - 0xc0
      13'h1985: dout  = 8'b10011000; // 6533 : 152 - 0x98
      13'h1986: dout  = 8'b00000000; // 6534 :   0 - 0x0
      13'h1987: dout  = 8'b00000000; // 6535 :   0 - 0x0
      13'h1988: dout  = 8'b10000000; // 6536 : 128 - 0x80
      13'h1989: dout  = 8'b11000000; // 6537 : 192 - 0xc0
      13'h198A: dout  = 8'b11000000; // 6538 : 192 - 0xc0
      13'h198B: dout  = 8'b11100000; // 6539 : 224 - 0xe0
      13'h198C: dout  = 8'b00100000; // 6540 :  32 - 0x20
      13'h198D: dout  = 8'b00111000; // 6541 :  56 - 0x38
      13'h198E: dout  = 8'b11111100; // 6542 : 252 - 0xfc
      13'h198F: dout  = 8'b11111110; // 6543 : 254 - 0xfe
      13'h1990: dout  = 8'b00000000; // 6544 :   0 - 0x0 -- Background 0x99
      13'h1991: dout  = 8'b00000000; // 6545 :   0 - 0x0
      13'h1992: dout  = 8'b00111110; // 6546 :  62 - 0x3e
      13'h1993: dout  = 8'b01000000; // 6547 :  64 - 0x40
      13'h1994: dout  = 8'b10000000; // 6548 : 128 - 0x80
      13'h1995: dout  = 8'b00000000; // 6549 :   0 - 0x0
      13'h1996: dout  = 8'b00000000; // 6550 :   0 - 0x0
      13'h1997: dout  = 8'b00000000; // 6551 :   0 - 0x0
      13'h1998: dout  = 8'b11111110; // 6552 : 254 - 0xfe
      13'h1999: dout  = 8'b11111111; // 6553 : 255 - 0xff
      13'h199A: dout  = 8'b11111111; // 6554 : 255 - 0xff
      13'h199B: dout  = 8'b11111110; // 6555 : 254 - 0xfe
      13'h199C: dout  = 8'b11111100; // 6556 : 252 - 0xfc
      13'h199D: dout  = 8'b11111000; // 6557 : 248 - 0xf8
      13'h199E: dout  = 8'b11000000; // 6558 : 192 - 0xc0
      13'h199F: dout  = 8'b00000000; // 6559 :   0 - 0x0
      13'h19A0: dout  = 8'b00000000; // 6560 :   0 - 0x0 -- Background 0x9a
      13'h19A1: dout  = 8'b00000000; // 6561 :   0 - 0x0
      13'h19A2: dout  = 8'b10000000; // 6562 : 128 - 0x80
      13'h19A3: dout  = 8'b10000000; // 6563 : 128 - 0x80
      13'h19A4: dout  = 8'b11000000; // 6564 : 192 - 0xc0
      13'h19A5: dout  = 8'b11100000; // 6565 : 224 - 0xe0
      13'h19A6: dout  = 8'b11100000; // 6566 : 224 - 0xe0
      13'h19A7: dout  = 8'b11110000; // 6567 : 240 - 0xf0
      13'h19A8: dout  = 8'b00000000; // 6568 :   0 - 0x0
      13'h19A9: dout  = 8'b00000000; // 6569 :   0 - 0x0
      13'h19AA: dout  = 8'b10000000; // 6570 : 128 - 0x80
      13'h19AB: dout  = 8'b10000000; // 6571 : 128 - 0x80
      13'h19AC: dout  = 8'b11000000; // 6572 : 192 - 0xc0
      13'h19AD: dout  = 8'b11100000; // 6573 : 224 - 0xe0
      13'h19AE: dout  = 8'b11100000; // 6574 : 224 - 0xe0
      13'h19AF: dout  = 8'b11110000; // 6575 : 240 - 0xf0
      13'h19B0: dout  = 8'b11110000; // 6576 : 240 - 0xf0 -- Background 0x9b
      13'h19B1: dout  = 8'b11100000; // 6577 : 224 - 0xe0
      13'h19B2: dout  = 8'b11110000; // 6578 : 240 - 0xf0
      13'h19B3: dout  = 8'b11100000; // 6579 : 224 - 0xe0
      13'h19B4: dout  = 8'b10000000; // 6580 : 128 - 0x80
      13'h19B5: dout  = 8'b00001000; // 6581 :   8 - 0x8
      13'h19B6: dout  = 8'b00000100; // 6582 :   4 - 0x4
      13'h19B7: dout  = 8'b00000000; // 6583 :   0 - 0x0
      13'h19B8: dout  = 8'b11111111; // 6584 : 255 - 0xff
      13'h19B9: dout  = 8'b11111111; // 6585 : 255 - 0xff
      13'h19BA: dout  = 8'b11111100; // 6586 : 252 - 0xfc
      13'h19BB: dout  = 8'b11111100; // 6587 : 252 - 0xfc
      13'h19BC: dout  = 8'b11111110; // 6588 : 254 - 0xfe
      13'h19BD: dout  = 8'b01111110; // 6589 : 126 - 0x7e
      13'h19BE: dout  = 8'b00111111; // 6590 :  63 - 0x3f
      13'h19BF: dout  = 8'b00001100; // 6591 :  12 - 0xc
      13'h19C0: dout  = 8'b00000000; // 6592 :   0 - 0x0 -- Background 0x9c
      13'h19C1: dout  = 8'b00000000; // 6593 :   0 - 0x0
      13'h19C2: dout  = 8'b00000001; // 6594 :   1 - 0x1
      13'h19C3: dout  = 8'b00000011; // 6595 :   3 - 0x3
      13'h19C4: dout  = 8'b00000011; // 6596 :   3 - 0x3
      13'h19C5: dout  = 8'b00000011; // 6597 :   3 - 0x3
      13'h19C6: dout  = 8'b00000111; // 6598 :   7 - 0x7
      13'h19C7: dout  = 8'b00000111; // 6599 :   7 - 0x7
      13'h19C8: dout  = 8'b00000000; // 6600 :   0 - 0x0
      13'h19C9: dout  = 8'b00000001; // 6601 :   1 - 0x1
      13'h19CA: dout  = 8'b00000011; // 6602 :   3 - 0x3
      13'h19CB: dout  = 8'b00000111; // 6603 :   7 - 0x7
      13'h19CC: dout  = 8'b00000111; // 6604 :   7 - 0x7
      13'h19CD: dout  = 8'b00000111; // 6605 :   7 - 0x7
      13'h19CE: dout  = 8'b00001111; // 6606 :  15 - 0xf
      13'h19CF: dout  = 8'b00001111; // 6607 :  15 - 0xf
      13'h19D0: dout  = 8'b00000111; // 6608 :   7 - 0x7 -- Background 0x9d
      13'h19D1: dout  = 8'b00000011; // 6609 :   3 - 0x3
      13'h19D2: dout  = 8'b00000011; // 6610 :   3 - 0x3
      13'h19D3: dout  = 8'b00000011; // 6611 :   3 - 0x3
      13'h19D4: dout  = 8'b00000011; // 6612 :   3 - 0x3
      13'h19D5: dout  = 8'b00000011; // 6613 :   3 - 0x3
      13'h19D6: dout  = 8'b00000011; // 6614 :   3 - 0x3
      13'h19D7: dout  = 8'b00000001; // 6615 :   1 - 0x1
      13'h19D8: dout  = 8'b00001111; // 6616 :  15 - 0xf
      13'h19D9: dout  = 8'b00001111; // 6617 :  15 - 0xf
      13'h19DA: dout  = 8'b00000111; // 6618 :   7 - 0x7
      13'h19DB: dout  = 8'b00000111; // 6619 :   7 - 0x7
      13'h19DC: dout  = 8'b00000111; // 6620 :   7 - 0x7
      13'h19DD: dout  = 8'b00000011; // 6621 :   3 - 0x3
      13'h19DE: dout  = 8'b00000011; // 6622 :   3 - 0x3
      13'h19DF: dout  = 8'b00000001; // 6623 :   1 - 0x1
      13'h19E0: dout  = 8'b00000000; // 6624 :   0 - 0x0 -- Background 0x9e
      13'h19E1: dout  = 8'b00000000; // 6625 :   0 - 0x0
      13'h19E2: dout  = 8'b00000000; // 6626 :   0 - 0x0
      13'h19E3: dout  = 8'b00000000; // 6627 :   0 - 0x0
      13'h19E4: dout  = 8'b00000000; // 6628 :   0 - 0x0
      13'h19E5: dout  = 8'b00000001; // 6629 :   1 - 0x1
      13'h19E6: dout  = 8'b00000010; // 6630 :   2 - 0x2
      13'h19E7: dout  = 8'b00000100; // 6631 :   4 - 0x4
      13'h19E8: dout  = 8'b00000001; // 6632 :   1 - 0x1
      13'h19E9: dout  = 8'b00000001; // 6633 :   1 - 0x1
      13'h19EA: dout  = 8'b00000001; // 6634 :   1 - 0x1
      13'h19EB: dout  = 8'b00000000; // 6635 :   0 - 0x0
      13'h19EC: dout  = 8'b00000000; // 6636 :   0 - 0x0
      13'h19ED: dout  = 8'b00000011; // 6637 :   3 - 0x3
      13'h19EE: dout  = 8'b00000111; // 6638 :   7 - 0x7
      13'h19EF: dout  = 8'b00001111; // 6639 :  15 - 0xf
      13'h19F0: dout  = 8'b00000000; // 6640 :   0 - 0x0 -- Background 0x9f
      13'h19F1: dout  = 8'b00000000; // 6641 :   0 - 0x0
      13'h19F2: dout  = 8'b00000000; // 6642 :   0 - 0x0
      13'h19F3: dout  = 8'b00000000; // 6643 :   0 - 0x0
      13'h19F4: dout  = 8'b00000000; // 6644 :   0 - 0x0
      13'h19F5: dout  = 8'b00000000; // 6645 :   0 - 0x0
      13'h19F6: dout  = 8'b00011100; // 6646 :  28 - 0x1c
      13'h19F7: dout  = 8'b00111011; // 6647 :  59 - 0x3b
      13'h19F8: dout  = 8'b00000000; // 6648 :   0 - 0x0
      13'h19F9: dout  = 8'b00000000; // 6649 :   0 - 0x0
      13'h19FA: dout  = 8'b00000000; // 6650 :   0 - 0x0
      13'h19FB: dout  = 8'b00000000; // 6651 :   0 - 0x0
      13'h19FC: dout  = 8'b00000001; // 6652 :   1 - 0x1
      13'h19FD: dout  = 8'b00000011; // 6653 :   3 - 0x3
      13'h19FE: dout  = 8'b00111111; // 6654 :  63 - 0x3f
      13'h19FF: dout  = 8'b01111111; // 6655 : 127 - 0x7f
      13'h1A00: dout  = 8'b01111110; // 6656 : 126 - 0x7e -- Background 0xa0
      13'h1A01: dout  = 8'b11111110; // 6657 : 254 - 0xfe
      13'h1A02: dout  = 8'b11111111; // 6658 : 255 - 0xff
      13'h1A03: dout  = 8'b11111111; // 6659 : 255 - 0xff
      13'h1A04: dout  = 8'b11111111; // 6660 : 255 - 0xff
      13'h1A05: dout  = 8'b11111111; // 6661 : 255 - 0xff
      13'h1A06: dout  = 8'b11111101; // 6662 : 253 - 0xfd
      13'h1A07: dout  = 8'b11111001; // 6663 : 249 - 0xf9
      13'h1A08: dout  = 8'b11111111; // 6664 : 255 - 0xff
      13'h1A09: dout  = 8'b11111111; // 6665 : 255 - 0xff
      13'h1A0A: dout  = 8'b11111111; // 6666 : 255 - 0xff
      13'h1A0B: dout  = 8'b11111111; // 6667 : 255 - 0xff
      13'h1A0C: dout  = 8'b11111111; // 6668 : 255 - 0xff
      13'h1A0D: dout  = 8'b11111111; // 6669 : 255 - 0xff
      13'h1A0E: dout  = 8'b11111101; // 6670 : 253 - 0xfd
      13'h1A0F: dout  = 8'b11111001; // 6671 : 249 - 0xf9
      13'h1A10: dout  = 8'b11110011; // 6672 : 243 - 0xf3 -- Background 0xa1
      13'h1A11: dout  = 8'b11110111; // 6673 : 247 - 0xf7
      13'h1A12: dout  = 8'b11110110; // 6674 : 246 - 0xf6
      13'h1A13: dout  = 8'b11101110; // 6675 : 238 - 0xee
      13'h1A14: dout  = 8'b11111101; // 6676 : 253 - 0xfd
      13'h1A15: dout  = 8'b11111100; // 6677 : 252 - 0xfc
      13'h1A16: dout  = 8'b11111000; // 6678 : 248 - 0xf8
      13'h1A17: dout  = 8'b11100001; // 6679 : 225 - 0xe1
      13'h1A18: dout  = 8'b11110011; // 6680 : 243 - 0xf3
      13'h1A19: dout  = 8'b11111111; // 6681 : 255 - 0xff
      13'h1A1A: dout  = 8'b11111111; // 6682 : 255 - 0xff
      13'h1A1B: dout  = 8'b11111111; // 6683 : 255 - 0xff
      13'h1A1C: dout  = 8'b11111111; // 6684 : 255 - 0xff
      13'h1A1D: dout  = 8'b11111111; // 6685 : 255 - 0xff
      13'h1A1E: dout  = 8'b11111111; // 6686 : 255 - 0xff
      13'h1A1F: dout  = 8'b11111111; // 6687 : 255 - 0xff
      13'h1A20: dout  = 8'b11010011; // 6688 : 211 - 0xd3 -- Background 0xa2
      13'h1A21: dout  = 8'b11001011; // 6689 : 203 - 0xcb
      13'h1A22: dout  = 8'b11000011; // 6690 : 195 - 0xc3
      13'h1A23: dout  = 8'b11100001; // 6691 : 225 - 0xe1
      13'h1A24: dout  = 8'b11111001; // 6692 : 249 - 0xf9
      13'h1A25: dout  = 8'b00111001; // 6693 :  57 - 0x39
      13'h1A26: dout  = 8'b01000010; // 6694 :  66 - 0x42
      13'h1A27: dout  = 8'b00000000; // 6695 :   0 - 0x0
      13'h1A28: dout  = 8'b11111111; // 6696 : 255 - 0xff
      13'h1A29: dout  = 8'b11111111; // 6697 : 255 - 0xff
      13'h1A2A: dout  = 8'b11111111; // 6698 : 255 - 0xff
      13'h1A2B: dout  = 8'b11111111; // 6699 : 255 - 0xff
      13'h1A2C: dout  = 8'b11111111; // 6700 : 255 - 0xff
      13'h1A2D: dout  = 8'b11111111; // 6701 : 255 - 0xff
      13'h1A2E: dout  = 8'b11111111; // 6702 : 255 - 0xff
      13'h1A2F: dout  = 8'b11111111; // 6703 : 255 - 0xff
      13'h1A30: dout  = 8'b00000111; // 6704 :   7 - 0x7 -- Background 0xa3
      13'h1A31: dout  = 8'b00001111; // 6705 :  15 - 0xf
      13'h1A32: dout  = 8'b00011001; // 6706 :  25 - 0x19
      13'h1A33: dout  = 8'b00110000; // 6707 :  48 - 0x30
      13'h1A34: dout  = 8'b01100011; // 6708 :  99 - 0x63
      13'h1A35: dout  = 8'b01110010; // 6709 : 114 - 0x72
      13'h1A36: dout  = 8'b01110000; // 6710 : 112 - 0x70
      13'h1A37: dout  = 8'b00000001; // 6711 :   1 - 0x1
      13'h1A38: dout  = 8'b00000111; // 6712 :   7 - 0x7
      13'h1A39: dout  = 8'b00001111; // 6713 :  15 - 0xf
      13'h1A3A: dout  = 8'b00011111; // 6714 :  31 - 0x1f
      13'h1A3B: dout  = 8'b00111111; // 6715 :  63 - 0x3f
      13'h1A3C: dout  = 8'b11111100; // 6716 : 252 - 0xfc
      13'h1A3D: dout  = 8'b11111100; // 6717 : 252 - 0xfc
      13'h1A3E: dout  = 8'b11111111; // 6718 : 255 - 0xff
      13'h1A3F: dout  = 8'b11111111; // 6719 : 255 - 0xff
      13'h1A40: dout  = 8'b00000000; // 6720 :   0 - 0x0 -- Background 0xa4
      13'h1A41: dout  = 8'b00011111; // 6721 :  31 - 0x1f
      13'h1A42: dout  = 8'b00100000; // 6722 :  32 - 0x20
      13'h1A43: dout  = 8'b11000000; // 6723 : 192 - 0xc0
      13'h1A44: dout  = 8'b11000000; // 6724 : 192 - 0xc0
      13'h1A45: dout  = 8'b11110000; // 6725 : 240 - 0xf0
      13'h1A46: dout  = 8'b11111111; // 6726 : 255 - 0xff
      13'h1A47: dout  = 8'b11111111; // 6727 : 255 - 0xff
      13'h1A48: dout  = 8'b11111111; // 6728 : 255 - 0xff
      13'h1A49: dout  = 8'b11111111; // 6729 : 255 - 0xff
      13'h1A4A: dout  = 8'b11111111; // 6730 : 255 - 0xff
      13'h1A4B: dout  = 8'b11111111; // 6731 : 255 - 0xff
      13'h1A4C: dout  = 8'b11111111; // 6732 : 255 - 0xff
      13'h1A4D: dout  = 8'b11111111; // 6733 : 255 - 0xff
      13'h1A4E: dout  = 8'b11111111; // 6734 : 255 - 0xff
      13'h1A4F: dout  = 8'b11111111; // 6735 : 255 - 0xff
      13'h1A50: dout  = 8'b10101011; // 6736 : 171 - 0xab -- Background 0xa5
      13'h1A51: dout  = 8'b11000001; // 6737 : 193 - 0xc1
      13'h1A52: dout  = 8'b10000001; // 6738 : 129 - 0x81
      13'h1A53: dout  = 8'b10010001; // 6739 : 145 - 0x91
      13'h1A54: dout  = 8'b10000010; // 6740 : 130 - 0x82
      13'h1A55: dout  = 8'b11111100; // 6741 : 252 - 0xfc
      13'h1A56: dout  = 8'b11100000; // 6742 : 224 - 0xe0
      13'h1A57: dout  = 8'b11001110; // 6743 : 206 - 0xce
      13'h1A58: dout  = 8'b11111111; // 6744 : 255 - 0xff
      13'h1A59: dout  = 8'b11111111; // 6745 : 255 - 0xff
      13'h1A5A: dout  = 8'b11111111; // 6746 : 255 - 0xff
      13'h1A5B: dout  = 8'b11111111; // 6747 : 255 - 0xff
      13'h1A5C: dout  = 8'b11111111; // 6748 : 255 - 0xff
      13'h1A5D: dout  = 8'b11111111; // 6749 : 255 - 0xff
      13'h1A5E: dout  = 8'b11111111; // 6750 : 255 - 0xff
      13'h1A5F: dout  = 8'b11111111; // 6751 : 255 - 0xff
      13'h1A60: dout  = 8'b11100101; // 6752 : 229 - 0xe5 -- Background 0xa6
      13'h1A61: dout  = 8'b11011010; // 6753 : 218 - 0xda
      13'h1A62: dout  = 8'b11110000; // 6754 : 240 - 0xf0
      13'h1A63: dout  = 8'b11100000; // 6755 : 224 - 0xe0
      13'h1A64: dout  = 8'b11000000; // 6756 : 192 - 0xc0
      13'h1A65: dout  = 8'b00000000; // 6757 :   0 - 0x0
      13'h1A66: dout  = 8'b00000000; // 6758 :   0 - 0x0
      13'h1A67: dout  = 8'b00000000; // 6759 :   0 - 0x0
      13'h1A68: dout  = 8'b11111111; // 6760 : 255 - 0xff
      13'h1A69: dout  = 8'b11111111; // 6761 : 255 - 0xff
      13'h1A6A: dout  = 8'b11110000; // 6762 : 240 - 0xf0
      13'h1A6B: dout  = 8'b11100000; // 6763 : 224 - 0xe0
      13'h1A6C: dout  = 8'b11000000; // 6764 : 192 - 0xc0
      13'h1A6D: dout  = 8'b10000000; // 6765 : 128 - 0x80
      13'h1A6E: dout  = 8'b10000000; // 6766 : 128 - 0x80
      13'h1A6F: dout  = 8'b00000000; // 6767 :   0 - 0x0
      13'h1A70: dout  = 8'b11110000; // 6768 : 240 - 0xf0 -- Background 0xa7
      13'h1A71: dout  = 8'b11111000; // 6769 : 248 - 0xf8
      13'h1A72: dout  = 8'b11001100; // 6770 : 204 - 0xcc
      13'h1A73: dout  = 8'b10000110; // 6771 : 134 - 0x86
      13'h1A74: dout  = 8'b01100010; // 6772 :  98 - 0x62
      13'h1A75: dout  = 8'b00100110; // 6773 :  38 - 0x26
      13'h1A76: dout  = 8'b00000110; // 6774 :   6 - 0x6
      13'h1A77: dout  = 8'b11000000; // 6775 : 192 - 0xc0
      13'h1A78: dout  = 8'b11110000; // 6776 : 240 - 0xf0
      13'h1A79: dout  = 8'b11111000; // 6777 : 248 - 0xf8
      13'h1A7A: dout  = 8'b11111100; // 6778 : 252 - 0xfc
      13'h1A7B: dout  = 8'b11111110; // 6779 : 254 - 0xfe
      13'h1A7C: dout  = 8'b10011111; // 6780 : 159 - 0x9f
      13'h1A7D: dout  = 8'b10011111; // 6781 : 159 - 0x9f
      13'h1A7E: dout  = 8'b11111111; // 6782 : 255 - 0xff
      13'h1A7F: dout  = 8'b11111111; // 6783 : 255 - 0xff
      13'h1A80: dout  = 8'b00000000; // 6784 :   0 - 0x0 -- Background 0xa8
      13'h1A81: dout  = 8'b11111100; // 6785 : 252 - 0xfc
      13'h1A82: dout  = 8'b00000110; // 6786 :   6 - 0x6
      13'h1A83: dout  = 8'b00000011; // 6787 :   3 - 0x3
      13'h1A84: dout  = 8'b00000001; // 6788 :   1 - 0x1
      13'h1A85: dout  = 8'b00000111; // 6789 :   7 - 0x7
      13'h1A86: dout  = 8'b11111111; // 6790 : 255 - 0xff
      13'h1A87: dout  = 8'b11111111; // 6791 : 255 - 0xff
      13'h1A88: dout  = 8'b11111111; // 6792 : 255 - 0xff
      13'h1A89: dout  = 8'b11111111; // 6793 : 255 - 0xff
      13'h1A8A: dout  = 8'b11111111; // 6794 : 255 - 0xff
      13'h1A8B: dout  = 8'b11111111; // 6795 : 255 - 0xff
      13'h1A8C: dout  = 8'b11111111; // 6796 : 255 - 0xff
      13'h1A8D: dout  = 8'b11111111; // 6797 : 255 - 0xff
      13'h1A8E: dout  = 8'b11111111; // 6798 : 255 - 0xff
      13'h1A8F: dout  = 8'b11111111; // 6799 : 255 - 0xff
      13'h1A90: dout  = 8'b11010101; // 6800 : 213 - 0xd5 -- Background 0xa9
      13'h1A91: dout  = 8'b10000011; // 6801 : 131 - 0x83
      13'h1A92: dout  = 8'b10000001; // 6802 : 129 - 0x81
      13'h1A93: dout  = 8'b10001001; // 6803 : 137 - 0x89
      13'h1A94: dout  = 8'b01000001; // 6804 :  65 - 0x41
      13'h1A95: dout  = 8'b00111111; // 6805 :  63 - 0x3f
      13'h1A96: dout  = 8'b00000111; // 6806 :   7 - 0x7
      13'h1A97: dout  = 8'b11010011; // 6807 : 211 - 0xd3
      13'h1A98: dout  = 8'b11111111; // 6808 : 255 - 0xff
      13'h1A99: dout  = 8'b11111111; // 6809 : 255 - 0xff
      13'h1A9A: dout  = 8'b11111111; // 6810 : 255 - 0xff
      13'h1A9B: dout  = 8'b11111111; // 6811 : 255 - 0xff
      13'h1A9C: dout  = 8'b11111111; // 6812 : 255 - 0xff
      13'h1A9D: dout  = 8'b11111111; // 6813 : 255 - 0xff
      13'h1A9E: dout  = 8'b11111111; // 6814 : 255 - 0xff
      13'h1A9F: dout  = 8'b11111111; // 6815 : 255 - 0xff
      13'h1AA0: dout  = 8'b01101111; // 6816 : 111 - 0x6f -- Background 0xaa
      13'h1AA1: dout  = 8'b11011011; // 6817 : 219 - 0xdb
      13'h1AA2: dout  = 8'b00001111; // 6818 :  15 - 0xf
      13'h1AA3: dout  = 8'b00000111; // 6819 :   7 - 0x7
      13'h1AA4: dout  = 8'b00000011; // 6820 :   3 - 0x3
      13'h1AA5: dout  = 8'b00000000; // 6821 :   0 - 0x0
      13'h1AA6: dout  = 8'b00000000; // 6822 :   0 - 0x0
      13'h1AA7: dout  = 8'b00000000; // 6823 :   0 - 0x0
      13'h1AA8: dout  = 8'b11111111; // 6824 : 255 - 0xff
      13'h1AA9: dout  = 8'b11111111; // 6825 : 255 - 0xff
      13'h1AAA: dout  = 8'b00001111; // 6826 :  15 - 0xf
      13'h1AAB: dout  = 8'b00000111; // 6827 :   7 - 0x7
      13'h1AAC: dout  = 8'b00000011; // 6828 :   3 - 0x3
      13'h1AAD: dout  = 8'b00000001; // 6829 :   1 - 0x1
      13'h1AAE: dout  = 8'b00000001; // 6830 :   1 - 0x1
      13'h1AAF: dout  = 8'b00000000; // 6831 :   0 - 0x0
      13'h1AB0: dout  = 8'b00000000; // 6832 :   0 - 0x0 -- Background 0xab
      13'h1AB1: dout  = 8'b00000000; // 6833 :   0 - 0x0
      13'h1AB2: dout  = 8'b00000000; // 6834 :   0 - 0x0
      13'h1AB3: dout  = 8'b00000000; // 6835 :   0 - 0x0
      13'h1AB4: dout  = 8'b00000000; // 6836 :   0 - 0x0
      13'h1AB5: dout  = 8'b00000000; // 6837 :   0 - 0x0
      13'h1AB6: dout  = 8'b00111000; // 6838 :  56 - 0x38
      13'h1AB7: dout  = 8'b11011100; // 6839 : 220 - 0xdc
      13'h1AB8: dout  = 8'b00000000; // 6840 :   0 - 0x0
      13'h1AB9: dout  = 8'b00000000; // 6841 :   0 - 0x0
      13'h1ABA: dout  = 8'b00000000; // 6842 :   0 - 0x0
      13'h1ABB: dout  = 8'b00000000; // 6843 :   0 - 0x0
      13'h1ABC: dout  = 8'b10000000; // 6844 : 128 - 0x80
      13'h1ABD: dout  = 8'b11000000; // 6845 : 192 - 0xc0
      13'h1ABE: dout  = 8'b11111100; // 6846 : 252 - 0xfc
      13'h1ABF: dout  = 8'b11111110; // 6847 : 254 - 0xfe
      13'h1AC0: dout  = 8'b01111110; // 6848 : 126 - 0x7e -- Background 0xac
      13'h1AC1: dout  = 8'b01111111; // 6849 : 127 - 0x7f
      13'h1AC2: dout  = 8'b01111111; // 6850 : 127 - 0x7f
      13'h1AC3: dout  = 8'b11111111; // 6851 : 255 - 0xff
      13'h1AC4: dout  = 8'b11111111; // 6852 : 255 - 0xff
      13'h1AC5: dout  = 8'b11111111; // 6853 : 255 - 0xff
      13'h1AC6: dout  = 8'b10111111; // 6854 : 191 - 0xbf
      13'h1AC7: dout  = 8'b10011111; // 6855 : 159 - 0x9f
      13'h1AC8: dout  = 8'b11111111; // 6856 : 255 - 0xff
      13'h1AC9: dout  = 8'b11111111; // 6857 : 255 - 0xff
      13'h1ACA: dout  = 8'b11111111; // 6858 : 255 - 0xff
      13'h1ACB: dout  = 8'b11111111; // 6859 : 255 - 0xff
      13'h1ACC: dout  = 8'b11111111; // 6860 : 255 - 0xff
      13'h1ACD: dout  = 8'b11111111; // 6861 : 255 - 0xff
      13'h1ACE: dout  = 8'b10111111; // 6862 : 191 - 0xbf
      13'h1ACF: dout  = 8'b10011111; // 6863 : 159 - 0x9f
      13'h1AD0: dout  = 8'b11001111; // 6864 : 207 - 0xcf -- Background 0xad
      13'h1AD1: dout  = 8'b11101111; // 6865 : 239 - 0xef
      13'h1AD2: dout  = 8'b01101111; // 6866 : 111 - 0x6f
      13'h1AD3: dout  = 8'b01110111; // 6867 : 119 - 0x77
      13'h1AD4: dout  = 8'b10111111; // 6868 : 191 - 0xbf
      13'h1AD5: dout  = 8'b00111111; // 6869 :  63 - 0x3f
      13'h1AD6: dout  = 8'b00011111; // 6870 :  31 - 0x1f
      13'h1AD7: dout  = 8'b10000111; // 6871 : 135 - 0x87
      13'h1AD8: dout  = 8'b11001111; // 6872 : 207 - 0xcf
      13'h1AD9: dout  = 8'b11111111; // 6873 : 255 - 0xff
      13'h1ADA: dout  = 8'b11111111; // 6874 : 255 - 0xff
      13'h1ADB: dout  = 8'b11111111; // 6875 : 255 - 0xff
      13'h1ADC: dout  = 8'b11111111; // 6876 : 255 - 0xff
      13'h1ADD: dout  = 8'b11111111; // 6877 : 255 - 0xff
      13'h1ADE: dout  = 8'b11111111; // 6878 : 255 - 0xff
      13'h1ADF: dout  = 8'b11111111; // 6879 : 255 - 0xff
      13'h1AE0: dout  = 8'b11001011; // 6880 : 203 - 0xcb -- Background 0xae
      13'h1AE1: dout  = 8'b11010011; // 6881 : 211 - 0xd3
      13'h1AE2: dout  = 8'b11000011; // 6882 : 195 - 0xc3
      13'h1AE3: dout  = 8'b10000111; // 6883 : 135 - 0x87
      13'h1AE4: dout  = 8'b10011111; // 6884 : 159 - 0x9f
      13'h1AE5: dout  = 8'b10011100; // 6885 : 156 - 0x9c
      13'h1AE6: dout  = 8'b01000010; // 6886 :  66 - 0x42
      13'h1AE7: dout  = 8'b00000000; // 6887 :   0 - 0x0
      13'h1AE8: dout  = 8'b11111111; // 6888 : 255 - 0xff
      13'h1AE9: dout  = 8'b11111111; // 6889 : 255 - 0xff
      13'h1AEA: dout  = 8'b11111111; // 6890 : 255 - 0xff
      13'h1AEB: dout  = 8'b11111111; // 6891 : 255 - 0xff
      13'h1AEC: dout  = 8'b11111111; // 6892 : 255 - 0xff
      13'h1AED: dout  = 8'b11111111; // 6893 : 255 - 0xff
      13'h1AEE: dout  = 8'b11111111; // 6894 : 255 - 0xff
      13'h1AEF: dout  = 8'b11111111; // 6895 : 255 - 0xff
      13'h1AF0: dout  = 8'b00000000; // 6896 :   0 - 0x0 -- Background 0xaf
      13'h1AF1: dout  = 8'b00000000; // 6897 :   0 - 0x0
      13'h1AF2: dout  = 8'b10000000; // 6898 : 128 - 0x80
      13'h1AF3: dout  = 8'b11000000; // 6899 : 192 - 0xc0
      13'h1AF4: dout  = 8'b11000000; // 6900 : 192 - 0xc0
      13'h1AF5: dout  = 8'b11000000; // 6901 : 192 - 0xc0
      13'h1AF6: dout  = 8'b11100000; // 6902 : 224 - 0xe0
      13'h1AF7: dout  = 8'b11100000; // 6903 : 224 - 0xe0
      13'h1AF8: dout  = 8'b00000000; // 6904 :   0 - 0x0
      13'h1AF9: dout  = 8'b10000000; // 6905 : 128 - 0x80
      13'h1AFA: dout  = 8'b11000000; // 6906 : 192 - 0xc0
      13'h1AFB: dout  = 8'b11100000; // 6907 : 224 - 0xe0
      13'h1AFC: dout  = 8'b11100000; // 6908 : 224 - 0xe0
      13'h1AFD: dout  = 8'b11100000; // 6909 : 224 - 0xe0
      13'h1AFE: dout  = 8'b11110000; // 6910 : 240 - 0xf0
      13'h1AFF: dout  = 8'b11110000; // 6911 : 240 - 0xf0
      13'h1B00: dout  = 8'b11100000; // 6912 : 224 - 0xe0 -- Background 0xb0
      13'h1B01: dout  = 8'b11000000; // 6913 : 192 - 0xc0
      13'h1B02: dout  = 8'b11000000; // 6914 : 192 - 0xc0
      13'h1B03: dout  = 8'b11000000; // 6915 : 192 - 0xc0
      13'h1B04: dout  = 8'b11000000; // 6916 : 192 - 0xc0
      13'h1B05: dout  = 8'b11000000; // 6917 : 192 - 0xc0
      13'h1B06: dout  = 8'b11000000; // 6918 : 192 - 0xc0
      13'h1B07: dout  = 8'b10000000; // 6919 : 128 - 0x80
      13'h1B08: dout  = 8'b11110000; // 6920 : 240 - 0xf0
      13'h1B09: dout  = 8'b11110000; // 6921 : 240 - 0xf0
      13'h1B0A: dout  = 8'b11100000; // 6922 : 224 - 0xe0
      13'h1B0B: dout  = 8'b11100000; // 6923 : 224 - 0xe0
      13'h1B0C: dout  = 8'b11100000; // 6924 : 224 - 0xe0
      13'h1B0D: dout  = 8'b11000000; // 6925 : 192 - 0xc0
      13'h1B0E: dout  = 8'b11000000; // 6926 : 192 - 0xc0
      13'h1B0F: dout  = 8'b10000000; // 6927 : 128 - 0x80
      13'h1B10: dout  = 8'b00000000; // 6928 :   0 - 0x0 -- Background 0xb1
      13'h1B11: dout  = 8'b00000000; // 6929 :   0 - 0x0
      13'h1B12: dout  = 8'b00000000; // 6930 :   0 - 0x0
      13'h1B13: dout  = 8'b00000000; // 6931 :   0 - 0x0
      13'h1B14: dout  = 8'b00000000; // 6932 :   0 - 0x0
      13'h1B15: dout  = 8'b10000000; // 6933 : 128 - 0x80
      13'h1B16: dout  = 8'b01000000; // 6934 :  64 - 0x40
      13'h1B17: dout  = 8'b00100000; // 6935 :  32 - 0x20
      13'h1B18: dout  = 8'b10000000; // 6936 : 128 - 0x80
      13'h1B19: dout  = 8'b10000000; // 6937 : 128 - 0x80
      13'h1B1A: dout  = 8'b10000000; // 6938 : 128 - 0x80
      13'h1B1B: dout  = 8'b00000000; // 6939 :   0 - 0x0
      13'h1B1C: dout  = 8'b00000000; // 6940 :   0 - 0x0
      13'h1B1D: dout  = 8'b11000000; // 6941 : 192 - 0xc0
      13'h1B1E: dout  = 8'b11100000; // 6942 : 224 - 0xe0
      13'h1B1F: dout  = 8'b11110000; // 6943 : 240 - 0xf0
      13'h1B20: dout  = 8'b00000000; // 6944 :   0 - 0x0 -- Background 0xb2
      13'h1B21: dout  = 8'b00000000; // 6945 :   0 - 0x0
      13'h1B22: dout  = 8'b00000000; // 6946 :   0 - 0x0
      13'h1B23: dout  = 8'b00000001; // 6947 :   1 - 0x1
      13'h1B24: dout  = 8'b00000011; // 6948 :   3 - 0x3
      13'h1B25: dout  = 8'b00000111; // 6949 :   7 - 0x7
      13'h1B26: dout  = 8'b00000111; // 6950 :   7 - 0x7
      13'h1B27: dout  = 8'b00000111; // 6951 :   7 - 0x7
      13'h1B28: dout  = 8'b00000000; // 6952 :   0 - 0x0
      13'h1B29: dout  = 8'b00000000; // 6953 :   0 - 0x0
      13'h1B2A: dout  = 8'b00000001; // 6954 :   1 - 0x1
      13'h1B2B: dout  = 8'b00000011; // 6955 :   3 - 0x3
      13'h1B2C: dout  = 8'b00000111; // 6956 :   7 - 0x7
      13'h1B2D: dout  = 8'b00000111; // 6957 :   7 - 0x7
      13'h1B2E: dout  = 8'b00000111; // 6958 :   7 - 0x7
      13'h1B2F: dout  = 8'b00000111; // 6959 :   7 - 0x7
      13'h1B30: dout  = 8'b00000011; // 6960 :   3 - 0x3 -- Background 0xb3
      13'h1B31: dout  = 8'b00000001; // 6961 :   1 - 0x1
      13'h1B32: dout  = 8'b00000000; // 6962 :   0 - 0x0
      13'h1B33: dout  = 8'b00000000; // 6963 :   0 - 0x0
      13'h1B34: dout  = 8'b00000000; // 6964 :   0 - 0x0
      13'h1B35: dout  = 8'b00000000; // 6965 :   0 - 0x0
      13'h1B36: dout  = 8'b00000001; // 6966 :   1 - 0x1
      13'h1B37: dout  = 8'b00000001; // 6967 :   1 - 0x1
      13'h1B38: dout  = 8'b00000011; // 6968 :   3 - 0x3
      13'h1B39: dout  = 8'b00000001; // 6969 :   1 - 0x1
      13'h1B3A: dout  = 8'b00000000; // 6970 :   0 - 0x0
      13'h1B3B: dout  = 8'b00000000; // 6971 :   0 - 0x0
      13'h1B3C: dout  = 8'b00000000; // 6972 :   0 - 0x0
      13'h1B3D: dout  = 8'b00000001; // 6973 :   1 - 0x1
      13'h1B3E: dout  = 8'b00000011; // 6974 :   3 - 0x3
      13'h1B3F: dout  = 8'b00000011; // 6975 :   3 - 0x3
      13'h1B40: dout  = 8'b00000001; // 6976 :   1 - 0x1 -- Background 0xb4
      13'h1B41: dout  = 8'b00000001; // 6977 :   1 - 0x1
      13'h1B42: dout  = 8'b00000111; // 6978 :   7 - 0x7
      13'h1B43: dout  = 8'b00000011; // 6979 :   3 - 0x3
      13'h1B44: dout  = 8'b00000100; // 6980 :   4 - 0x4
      13'h1B45: dout  = 8'b00000000; // 6981 :   0 - 0x0
      13'h1B46: dout  = 8'b00000000; // 6982 :   0 - 0x0
      13'h1B47: dout  = 8'b00000000; // 6983 :   0 - 0x0
      13'h1B48: dout  = 8'b00000011; // 6984 :   3 - 0x3
      13'h1B49: dout  = 8'b00000011; // 6985 :   3 - 0x3
      13'h1B4A: dout  = 8'b00000111; // 6986 :   7 - 0x7
      13'h1B4B: dout  = 8'b00011111; // 6987 :  31 - 0x1f
      13'h1B4C: dout  = 8'b00111111; // 6988 :  63 - 0x3f
      13'h1B4D: dout  = 8'b00111111; // 6989 :  63 - 0x3f
      13'h1B4E: dout  = 8'b00000000; // 6990 :   0 - 0x0
      13'h1B4F: dout  = 8'b00000000; // 6991 :   0 - 0x0
      13'h1B50: dout  = 8'b00000000; // 6992 :   0 - 0x0 -- Background 0xb5
      13'h1B51: dout  = 8'b00000000; // 6993 :   0 - 0x0
      13'h1B52: dout  = 8'b00000000; // 6994 :   0 - 0x0
      13'h1B53: dout  = 8'b00000000; // 6995 :   0 - 0x0
      13'h1B54: dout  = 8'b00000000; // 6996 :   0 - 0x0
      13'h1B55: dout  = 8'b00000000; // 6997 :   0 - 0x0
      13'h1B56: dout  = 8'b00000000; // 6998 :   0 - 0x0
      13'h1B57: dout  = 8'b00000111; // 6999 :   7 - 0x7
      13'h1B58: dout  = 8'b00000000; // 7000 :   0 - 0x0
      13'h1B59: dout  = 8'b00000000; // 7001 :   0 - 0x0
      13'h1B5A: dout  = 8'b00000000; // 7002 :   0 - 0x0
      13'h1B5B: dout  = 8'b00000000; // 7003 :   0 - 0x0
      13'h1B5C: dout  = 8'b00000001; // 7004 :   1 - 0x1
      13'h1B5D: dout  = 8'b00000011; // 7005 :   3 - 0x3
      13'h1B5E: dout  = 8'b00000011; // 7006 :   3 - 0x3
      13'h1B5F: dout  = 8'b00001111; // 7007 :  15 - 0xf
      13'h1B60: dout  = 8'b00001110; // 7008 :  14 - 0xe -- Background 0xb6
      13'h1B61: dout  = 8'b00111110; // 7009 :  62 - 0x3e
      13'h1B62: dout  = 8'b01111111; // 7010 : 127 - 0x7f
      13'h1B63: dout  = 8'b11111111; // 7011 : 255 - 0xff
      13'h1B64: dout  = 8'b11111111; // 7012 : 255 - 0xff
      13'h1B65: dout  = 8'b11101111; // 7013 : 239 - 0xef
      13'h1B66: dout  = 8'b11110111; // 7014 : 247 - 0xf7
      13'h1B67: dout  = 8'b11111000; // 7015 : 248 - 0xf8
      13'h1B68: dout  = 8'b00111111; // 7016 :  63 - 0x3f
      13'h1B69: dout  = 8'b01111111; // 7017 : 127 - 0x7f
      13'h1B6A: dout  = 8'b11111111; // 7018 : 255 - 0xff
      13'h1B6B: dout  = 8'b11111111; // 7019 : 255 - 0xff
      13'h1B6C: dout  = 8'b11111111; // 7020 : 255 - 0xff
      13'h1B6D: dout  = 8'b11111111; // 7021 : 255 - 0xff
      13'h1B6E: dout  = 8'b11111111; // 7022 : 255 - 0xff
      13'h1B6F: dout  = 8'b11111111; // 7023 : 255 - 0xff
      13'h1B70: dout  = 8'b11111111; // 7024 : 255 - 0xff -- Background 0xb7
      13'h1B71: dout  = 8'b11111111; // 7025 : 255 - 0xff
      13'h1B72: dout  = 8'b11111111; // 7026 : 255 - 0xff
      13'h1B73: dout  = 8'b00011111; // 7027 :  31 - 0x1f
      13'h1B74: dout  = 8'b00011111; // 7028 :  31 - 0x1f
      13'h1B75: dout  = 8'b01111111; // 7029 : 127 - 0x7f
      13'h1B76: dout  = 8'b11111111; // 7030 : 255 - 0xff
      13'h1B77: dout  = 8'b11111110; // 7031 : 254 - 0xfe
      13'h1B78: dout  = 8'b11111111; // 7032 : 255 - 0xff
      13'h1B79: dout  = 8'b11111111; // 7033 : 255 - 0xff
      13'h1B7A: dout  = 8'b11111111; // 7034 : 255 - 0xff
      13'h1B7B: dout  = 8'b00011111; // 7035 :  31 - 0x1f
      13'h1B7C: dout  = 8'b01111111; // 7036 : 127 - 0x7f
      13'h1B7D: dout  = 8'b11111111; // 7037 : 255 - 0xff
      13'h1B7E: dout  = 8'b11111111; // 7038 : 255 - 0xff
      13'h1B7F: dout  = 8'b11111111; // 7039 : 255 - 0xff
      13'h1B80: dout  = 8'b11111111; // 7040 : 255 - 0xff -- Background 0xb8
      13'h1B81: dout  = 8'b11111111; // 7041 : 255 - 0xff
      13'h1B82: dout  = 8'b11111111; // 7042 : 255 - 0xff
      13'h1B83: dout  = 8'b11111100; // 7043 : 252 - 0xfc
      13'h1B84: dout  = 8'b11111000; // 7044 : 248 - 0xf8
      13'h1B85: dout  = 8'b10000000; // 7045 : 128 - 0x80
      13'h1B86: dout  = 8'b00000000; // 7046 :   0 - 0x0
      13'h1B87: dout  = 8'b00000000; // 7047 :   0 - 0x0
      13'h1B88: dout  = 8'b11111111; // 7048 : 255 - 0xff
      13'h1B89: dout  = 8'b11111111; // 7049 : 255 - 0xff
      13'h1B8A: dout  = 8'b11111111; // 7050 : 255 - 0xff
      13'h1B8B: dout  = 8'b11111100; // 7051 : 252 - 0xfc
      13'h1B8C: dout  = 8'b11111000; // 7052 : 248 - 0xf8
      13'h1B8D: dout  = 8'b11111000; // 7053 : 248 - 0xf8
      13'h1B8E: dout  = 8'b00000000; // 7054 :   0 - 0x0
      13'h1B8F: dout  = 8'b00000000; // 7055 :   0 - 0x0
      13'h1B90: dout  = 8'b00110000; // 7056 :  48 - 0x30 -- Background 0xb9
      13'h1B91: dout  = 8'b01111111; // 7057 : 127 - 0x7f
      13'h1B92: dout  = 8'b01111111; // 7058 : 127 - 0x7f
      13'h1B93: dout  = 8'b00111111; // 7059 :  63 - 0x3f
      13'h1B94: dout  = 8'b10000111; // 7060 : 135 - 0x87
      13'h1B95: dout  = 8'b11110000; // 7061 : 240 - 0xf0
      13'h1B96: dout  = 8'b11111111; // 7062 : 255 - 0xff
      13'h1B97: dout  = 8'b11111111; // 7063 : 255 - 0xff
      13'h1B98: dout  = 8'b11001111; // 7064 : 207 - 0xcf
      13'h1B99: dout  = 8'b10001000; // 7065 : 136 - 0x88
      13'h1B9A: dout  = 8'b11011101; // 7066 : 221 - 0xdd
      13'h1B9B: dout  = 8'b11001000; // 7067 : 200 - 0xc8
      13'h1B9C: dout  = 8'b11111000; // 7068 : 248 - 0xf8
      13'h1B9D: dout  = 8'b11111111; // 7069 : 255 - 0xff
      13'h1B9E: dout  = 8'b11111111; // 7070 : 255 - 0xff
      13'h1B9F: dout  = 8'b11111111; // 7071 : 255 - 0xff
      13'h1BA0: dout  = 8'b11100101; // 7072 : 229 - 0xe5 -- Background 0xba
      13'h1BA1: dout  = 8'b11011010; // 7073 : 218 - 0xda
      13'h1BA2: dout  = 8'b11000000; // 7074 : 192 - 0xc0
      13'h1BA3: dout  = 8'b00000000; // 7075 :   0 - 0x0
      13'h1BA4: dout  = 8'b00000000; // 7076 :   0 - 0x0
      13'h1BA5: dout  = 8'b00000000; // 7077 :   0 - 0x0
      13'h1BA6: dout  = 8'b00000000; // 7078 :   0 - 0x0
      13'h1BA7: dout  = 8'b00000000; // 7079 :   0 - 0x0
      13'h1BA8: dout  = 8'b11111111; // 7080 : 255 - 0xff
      13'h1BA9: dout  = 8'b11111111; // 7081 : 255 - 0xff
      13'h1BAA: dout  = 8'b11000000; // 7082 : 192 - 0xc0
      13'h1BAB: dout  = 8'b00000000; // 7083 :   0 - 0x0
      13'h1BAC: dout  = 8'b00000000; // 7084 :   0 - 0x0
      13'h1BAD: dout  = 8'b00000000; // 7085 :   0 - 0x0
      13'h1BAE: dout  = 8'b00000000; // 7086 :   0 - 0x0
      13'h1BAF: dout  = 8'b00000000; // 7087 :   0 - 0x0
      13'h1BB0: dout  = 8'b00000110; // 7088 :   6 - 0x6 -- Background 0xbb
      13'h1BB1: dout  = 8'b11111111; // 7089 : 255 - 0xff
      13'h1BB2: dout  = 8'b11111111; // 7090 : 255 - 0xff
      13'h1BB3: dout  = 8'b11111110; // 7091 : 254 - 0xfe
      13'h1BB4: dout  = 8'b11110001; // 7092 : 241 - 0xf1
      13'h1BB5: dout  = 8'b00000111; // 7093 :   7 - 0x7
      13'h1BB6: dout  = 8'b11111111; // 7094 : 255 - 0xff
      13'h1BB7: dout  = 8'b11111111; // 7095 : 255 - 0xff
      13'h1BB8: dout  = 8'b11111001; // 7096 : 249 - 0xf9
      13'h1BB9: dout  = 8'b10001000; // 7097 : 136 - 0x88
      13'h1BBA: dout  = 8'b11011101; // 7098 : 221 - 0xdd
      13'h1BBB: dout  = 8'b10001001; // 7099 : 137 - 0x89
      13'h1BBC: dout  = 8'b00001111; // 7100 :  15 - 0xf
      13'h1BBD: dout  = 8'b11111111; // 7101 : 255 - 0xff
      13'h1BBE: dout  = 8'b11111111; // 7102 : 255 - 0xff
      13'h1BBF: dout  = 8'b11111111; // 7103 : 255 - 0xff
      13'h1BC0: dout  = 8'b00000000; // 7104 :   0 - 0x0 -- Background 0xbc
      13'h1BC1: dout  = 8'b00000001; // 7105 :   1 - 0x1
      13'h1BC2: dout  = 8'b00000010; // 7106 :   2 - 0x2
      13'h1BC3: dout  = 8'b00000111; // 7107 :   7 - 0x7
      13'h1BC4: dout  = 8'b00000000; // 7108 :   0 - 0x0
      13'h1BC5: dout  = 8'b00000000; // 7109 :   0 - 0x0
      13'h1BC6: dout  = 8'b00100000; // 7110 :  32 - 0x20
      13'h1BC7: dout  = 8'b11111111; // 7111 : 255 - 0xff
      13'h1BC8: dout  = 8'b00000011; // 7112 :   3 - 0x3
      13'h1BC9: dout  = 8'b00000111; // 7113 :   7 - 0x7
      13'h1BCA: dout  = 8'b00001111; // 7114 :  15 - 0xf
      13'h1BCB: dout  = 8'b00000111; // 7115 :   7 - 0x7
      13'h1BCC: dout  = 8'b10000111; // 7116 : 135 - 0x87
      13'h1BCD: dout  = 8'b11000011; // 7117 : 195 - 0xc3
      13'h1BCE: dout  = 8'b11100000; // 7118 : 224 - 0xe0
      13'h1BCF: dout  = 8'b11111111; // 7119 : 255 - 0xff
      13'h1BD0: dout  = 8'b01111111; // 7120 : 127 - 0x7f -- Background 0xbd
      13'h1BD1: dout  = 8'b01111111; // 7121 : 127 - 0x7f
      13'h1BD2: dout  = 8'b01111111; // 7122 : 127 - 0x7f
      13'h1BD3: dout  = 8'b11111111; // 7123 : 255 - 0xff
      13'h1BD4: dout  = 8'b11111111; // 7124 : 255 - 0xff
      13'h1BD5: dout  = 8'b11111111; // 7125 : 255 - 0xff
      13'h1BD6: dout  = 8'b11111111; // 7126 : 255 - 0xff
      13'h1BD7: dout  = 8'b11111110; // 7127 : 254 - 0xfe
      13'h1BD8: dout  = 8'b11111111; // 7128 : 255 - 0xff
      13'h1BD9: dout  = 8'b11111111; // 7129 : 255 - 0xff
      13'h1BDA: dout  = 8'b11111111; // 7130 : 255 - 0xff
      13'h1BDB: dout  = 8'b11111111; // 7131 : 255 - 0xff
      13'h1BDC: dout  = 8'b11111111; // 7132 : 255 - 0xff
      13'h1BDD: dout  = 8'b11111111; // 7133 : 255 - 0xff
      13'h1BDE: dout  = 8'b11111111; // 7134 : 255 - 0xff
      13'h1BDF: dout  = 8'b11111110; // 7135 : 254 - 0xfe
      13'h1BE0: dout  = 8'b11111100; // 7136 : 252 - 0xfc -- Background 0xbe
      13'h1BE1: dout  = 8'b10111000; // 7137 : 184 - 0xb8
      13'h1BE2: dout  = 8'b01111000; // 7138 : 120 - 0x78
      13'h1BE3: dout  = 8'b01111000; // 7139 : 120 - 0x78
      13'h1BE4: dout  = 8'b10110000; // 7140 : 176 - 0xb0
      13'h1BE5: dout  = 8'b01111000; // 7141 : 120 - 0x78
      13'h1BE6: dout  = 8'b11111100; // 7142 : 252 - 0xfc
      13'h1BE7: dout  = 8'b11111110; // 7143 : 254 - 0xfe
      13'h1BE8: dout  = 8'b11111100; // 7144 : 252 - 0xfc
      13'h1BE9: dout  = 8'b11111000; // 7145 : 248 - 0xf8
      13'h1BEA: dout  = 8'b11111000; // 7146 : 248 - 0xf8
      13'h1BEB: dout  = 8'b11111000; // 7147 : 248 - 0xf8
      13'h1BEC: dout  = 8'b11111000; // 7148 : 248 - 0xf8
      13'h1BED: dout  = 8'b11111100; // 7149 : 252 - 0xfc
      13'h1BEE: dout  = 8'b11111110; // 7150 : 254 - 0xfe
      13'h1BEF: dout  = 8'b11111111; // 7151 : 255 - 0xff
      13'h1BF0: dout  = 8'b11111111; // 7152 : 255 - 0xff -- Background 0xbf
      13'h1BF1: dout  = 8'b11111111; // 7153 : 255 - 0xff
      13'h1BF2: dout  = 8'b11111111; // 7154 : 255 - 0xff
      13'h1BF3: dout  = 8'b11111111; // 7155 : 255 - 0xff
      13'h1BF4: dout  = 8'b11111111; // 7156 : 255 - 0xff
      13'h1BF5: dout  = 8'b10011100; // 7157 : 156 - 0x9c
      13'h1BF6: dout  = 8'b01000010; // 7158 :  66 - 0x42
      13'h1BF7: dout  = 8'b00000000; // 7159 :   0 - 0x0
      13'h1BF8: dout  = 8'b11111111; // 7160 : 255 - 0xff
      13'h1BF9: dout  = 8'b11111111; // 7161 : 255 - 0xff
      13'h1BFA: dout  = 8'b11111111; // 7162 : 255 - 0xff
      13'h1BFB: dout  = 8'b11111111; // 7163 : 255 - 0xff
      13'h1BFC: dout  = 8'b11111111; // 7164 : 255 - 0xff
      13'h1BFD: dout  = 8'b11111111; // 7165 : 255 - 0xff
      13'h1BFE: dout  = 8'b11111111; // 7166 : 255 - 0xff
      13'h1BFF: dout  = 8'b11111111; // 7167 : 255 - 0xff
      13'h1C00: dout  = 8'b00000000; // 7168 :   0 - 0x0 -- Background 0xc0
      13'h1C01: dout  = 8'b00000000; // 7169 :   0 - 0x0
      13'h1C02: dout  = 8'b00100000; // 7170 :  32 - 0x20
      13'h1C03: dout  = 8'b01000000; // 7171 :  64 - 0x40
      13'h1C04: dout  = 8'b10001010; // 7172 : 138 - 0x8a
      13'h1C05: dout  = 8'b00011110; // 7173 :  30 - 0x1e
      13'h1C06: dout  = 8'b01111110; // 7174 : 126 - 0x7e
      13'h1C07: dout  = 8'b10111110; // 7175 : 190 - 0xbe
      13'h1C08: dout  = 8'b11000000; // 7176 : 192 - 0xc0
      13'h1C09: dout  = 8'b11110000; // 7177 : 240 - 0xf0
      13'h1C0A: dout  = 8'b11111100; // 7178 : 252 - 0xfc
      13'h1C0B: dout  = 8'b11111100; // 7179 : 252 - 0xfc
      13'h1C0C: dout  = 8'b11111110; // 7180 : 254 - 0xfe
      13'h1C0D: dout  = 8'b11111110; // 7181 : 254 - 0xfe
      13'h1C0E: dout  = 8'b11111110; // 7182 : 254 - 0xfe
      13'h1C0F: dout  = 8'b11111110; // 7183 : 254 - 0xfe
      13'h1C10: dout  = 8'b11011111; // 7184 : 223 - 0xdf -- Background 0xc1
      13'h1C11: dout  = 8'b11111111; // 7185 : 255 - 0xff
      13'h1C12: dout  = 8'b11111110; // 7186 : 254 - 0xfe
      13'h1C13: dout  = 8'b11111100; // 7187 : 252 - 0xfc
      13'h1C14: dout  = 8'b11110000; // 7188 : 240 - 0xf0
      13'h1C15: dout  = 8'b11100000; // 7189 : 224 - 0xe0
      13'h1C16: dout  = 8'b10000000; // 7190 : 128 - 0x80
      13'h1C17: dout  = 8'b00000000; // 7191 :   0 - 0x0
      13'h1C18: dout  = 8'b11111111; // 7192 : 255 - 0xff
      13'h1C19: dout  = 8'b11111111; // 7193 : 255 - 0xff
      13'h1C1A: dout  = 8'b11111110; // 7194 : 254 - 0xfe
      13'h1C1B: dout  = 8'b11111100; // 7195 : 252 - 0xfc
      13'h1C1C: dout  = 8'b11110000; // 7196 : 240 - 0xf0
      13'h1C1D: dout  = 8'b11100000; // 7197 : 224 - 0xe0
      13'h1C1E: dout  = 8'b10000000; // 7198 : 128 - 0x80
      13'h1C1F: dout  = 8'b00000000; // 7199 :   0 - 0x0
      13'h1C20: dout  = 8'b00000000; // 7200 :   0 - 0x0 -- Background 0xc2
      13'h1C21: dout  = 8'b00000000; // 7201 :   0 - 0x0
      13'h1C22: dout  = 8'b00000100; // 7202 :   4 - 0x4
      13'h1C23: dout  = 8'b00000010; // 7203 :   2 - 0x2
      13'h1C24: dout  = 8'b01010001; // 7204 :  81 - 0x51
      13'h1C25: dout  = 8'b01111000; // 7205 : 120 - 0x78
      13'h1C26: dout  = 8'b01111110; // 7206 : 126 - 0x7e
      13'h1C27: dout  = 8'b11111101; // 7207 : 253 - 0xfd
      13'h1C28: dout  = 8'b00000011; // 7208 :   3 - 0x3
      13'h1C29: dout  = 8'b00001111; // 7209 :  15 - 0xf
      13'h1C2A: dout  = 8'b00111111; // 7210 :  63 - 0x3f
      13'h1C2B: dout  = 8'b00111111; // 7211 :  63 - 0x3f
      13'h1C2C: dout  = 8'b01111111; // 7212 : 127 - 0x7f
      13'h1C2D: dout  = 8'b01111111; // 7213 : 127 - 0x7f
      13'h1C2E: dout  = 8'b01111110; // 7214 : 126 - 0x7e
      13'h1C2F: dout  = 8'b11111111; // 7215 : 255 - 0xff
      13'h1C30: dout  = 8'b11111011; // 7216 : 251 - 0xfb -- Background 0xc3
      13'h1C31: dout  = 8'b11111111; // 7217 : 255 - 0xff
      13'h1C32: dout  = 8'b01111111; // 7218 : 127 - 0x7f
      13'h1C33: dout  = 8'b00111111; // 7219 :  63 - 0x3f
      13'h1C34: dout  = 8'b00001111; // 7220 :  15 - 0xf
      13'h1C35: dout  = 8'b00000111; // 7221 :   7 - 0x7
      13'h1C36: dout  = 8'b00000001; // 7222 :   1 - 0x1
      13'h1C37: dout  = 8'b00000000; // 7223 :   0 - 0x0
      13'h1C38: dout  = 8'b11111111; // 7224 : 255 - 0xff
      13'h1C39: dout  = 8'b11111111; // 7225 : 255 - 0xff
      13'h1C3A: dout  = 8'b01111111; // 7226 : 127 - 0x7f
      13'h1C3B: dout  = 8'b00111111; // 7227 :  63 - 0x3f
      13'h1C3C: dout  = 8'b00001111; // 7228 :  15 - 0xf
      13'h1C3D: dout  = 8'b00000111; // 7229 :   7 - 0x7
      13'h1C3E: dout  = 8'b00000001; // 7230 :   1 - 0x1
      13'h1C3F: dout  = 8'b00000000; // 7231 :   0 - 0x0
      13'h1C40: dout  = 8'b00000000; // 7232 :   0 - 0x0 -- Background 0xc4
      13'h1C41: dout  = 8'b10000000; // 7233 : 128 - 0x80
      13'h1C42: dout  = 8'b01000000; // 7234 :  64 - 0x40
      13'h1C43: dout  = 8'b11100000; // 7235 : 224 - 0xe0
      13'h1C44: dout  = 8'b00000000; // 7236 :   0 - 0x0
      13'h1C45: dout  = 8'b00000000; // 7237 :   0 - 0x0
      13'h1C46: dout  = 8'b00000100; // 7238 :   4 - 0x4
      13'h1C47: dout  = 8'b11111111; // 7239 : 255 - 0xff
      13'h1C48: dout  = 8'b11000000; // 7240 : 192 - 0xc0
      13'h1C49: dout  = 8'b11100000; // 7241 : 224 - 0xe0
      13'h1C4A: dout  = 8'b11110000; // 7242 : 240 - 0xf0
      13'h1C4B: dout  = 8'b11100000; // 7243 : 224 - 0xe0
      13'h1C4C: dout  = 8'b11100001; // 7244 : 225 - 0xe1
      13'h1C4D: dout  = 8'b11000011; // 7245 : 195 - 0xc3
      13'h1C4E: dout  = 8'b00000111; // 7246 :   7 - 0x7
      13'h1C4F: dout  = 8'b11111111; // 7247 : 255 - 0xff
      13'h1C50: dout  = 8'b11111110; // 7248 : 254 - 0xfe -- Background 0xc5
      13'h1C51: dout  = 8'b11111110; // 7249 : 254 - 0xfe
      13'h1C52: dout  = 8'b11111110; // 7250 : 254 - 0xfe
      13'h1C53: dout  = 8'b11111111; // 7251 : 255 - 0xff
      13'h1C54: dout  = 8'b11111111; // 7252 : 255 - 0xff
      13'h1C55: dout  = 8'b11111111; // 7253 : 255 - 0xff
      13'h1C56: dout  = 8'b11111111; // 7254 : 255 - 0xff
      13'h1C57: dout  = 8'b01111111; // 7255 : 127 - 0x7f
      13'h1C58: dout  = 8'b11111111; // 7256 : 255 - 0xff
      13'h1C59: dout  = 8'b11111111; // 7257 : 255 - 0xff
      13'h1C5A: dout  = 8'b11111111; // 7258 : 255 - 0xff
      13'h1C5B: dout  = 8'b11111111; // 7259 : 255 - 0xff
      13'h1C5C: dout  = 8'b11111111; // 7260 : 255 - 0xff
      13'h1C5D: dout  = 8'b11111111; // 7261 : 255 - 0xff
      13'h1C5E: dout  = 8'b11111111; // 7262 : 255 - 0xff
      13'h1C5F: dout  = 8'b01111111; // 7263 : 127 - 0x7f
      13'h1C60: dout  = 8'b00111111; // 7264 :  63 - 0x3f -- Background 0xc6
      13'h1C61: dout  = 8'b00011101; // 7265 :  29 - 0x1d
      13'h1C62: dout  = 8'b00011110; // 7266 :  30 - 0x1e
      13'h1C63: dout  = 8'b00011110; // 7267 :  30 - 0x1e
      13'h1C64: dout  = 8'b00001101; // 7268 :  13 - 0xd
      13'h1C65: dout  = 8'b00011110; // 7269 :  30 - 0x1e
      13'h1C66: dout  = 8'b00111111; // 7270 :  63 - 0x3f
      13'h1C67: dout  = 8'b01111111; // 7271 : 127 - 0x7f
      13'h1C68: dout  = 8'b00111111; // 7272 :  63 - 0x3f
      13'h1C69: dout  = 8'b00011111; // 7273 :  31 - 0x1f
      13'h1C6A: dout  = 8'b00011111; // 7274 :  31 - 0x1f
      13'h1C6B: dout  = 8'b00011111; // 7275 :  31 - 0x1f
      13'h1C6C: dout  = 8'b00011111; // 7276 :  31 - 0x1f
      13'h1C6D: dout  = 8'b00111111; // 7277 :  63 - 0x3f
      13'h1C6E: dout  = 8'b01111111; // 7278 : 127 - 0x7f
      13'h1C6F: dout  = 8'b11111111; // 7279 : 255 - 0xff
      13'h1C70: dout  = 8'b11111111; // 7280 : 255 - 0xff -- Background 0xc7
      13'h1C71: dout  = 8'b11111111; // 7281 : 255 - 0xff
      13'h1C72: dout  = 8'b11111111; // 7282 : 255 - 0xff
      13'h1C73: dout  = 8'b11111111; // 7283 : 255 - 0xff
      13'h1C74: dout  = 8'b11111111; // 7284 : 255 - 0xff
      13'h1C75: dout  = 8'b00111001; // 7285 :  57 - 0x39
      13'h1C76: dout  = 8'b01000010; // 7286 :  66 - 0x42
      13'h1C77: dout  = 8'b00000000; // 7287 :   0 - 0x0
      13'h1C78: dout  = 8'b11111111; // 7288 : 255 - 0xff
      13'h1C79: dout  = 8'b11111111; // 7289 : 255 - 0xff
      13'h1C7A: dout  = 8'b11111111; // 7290 : 255 - 0xff
      13'h1C7B: dout  = 8'b11111111; // 7291 : 255 - 0xff
      13'h1C7C: dout  = 8'b11111111; // 7292 : 255 - 0xff
      13'h1C7D: dout  = 8'b11111111; // 7293 : 255 - 0xff
      13'h1C7E: dout  = 8'b11111111; // 7294 : 255 - 0xff
      13'h1C7F: dout  = 8'b11111111; // 7295 : 255 - 0xff
      13'h1C80: dout  = 8'b01101111; // 7296 : 111 - 0x6f -- Background 0xc8
      13'h1C81: dout  = 8'b11011011; // 7297 : 219 - 0xdb
      13'h1C82: dout  = 8'b00000011; // 7298 :   3 - 0x3
      13'h1C83: dout  = 8'b00000000; // 7299 :   0 - 0x0
      13'h1C84: dout  = 8'b00000000; // 7300 :   0 - 0x0
      13'h1C85: dout  = 8'b00000000; // 7301 :   0 - 0x0
      13'h1C86: dout  = 8'b00000000; // 7302 :   0 - 0x0
      13'h1C87: dout  = 8'b00000000; // 7303 :   0 - 0x0
      13'h1C88: dout  = 8'b11111111; // 7304 : 255 - 0xff
      13'h1C89: dout  = 8'b11111111; // 7305 : 255 - 0xff
      13'h1C8A: dout  = 8'b00000011; // 7306 :   3 - 0x3
      13'h1C8B: dout  = 8'b00000000; // 7307 :   0 - 0x0
      13'h1C8C: dout  = 8'b00000000; // 7308 :   0 - 0x0
      13'h1C8D: dout  = 8'b00000000; // 7309 :   0 - 0x0
      13'h1C8E: dout  = 8'b00000000; // 7310 :   0 - 0x0
      13'h1C8F: dout  = 8'b00000000; // 7311 :   0 - 0x0
      13'h1C90: dout  = 8'b00000000; // 7312 :   0 - 0x0 -- Background 0xc9
      13'h1C91: dout  = 8'b00000000; // 7313 :   0 - 0x0
      13'h1C92: dout  = 8'b00000000; // 7314 :   0 - 0x0
      13'h1C93: dout  = 8'b00000000; // 7315 :   0 - 0x0
      13'h1C94: dout  = 8'b00000000; // 7316 :   0 - 0x0
      13'h1C95: dout  = 8'b00000000; // 7317 :   0 - 0x0
      13'h1C96: dout  = 8'b00000000; // 7318 :   0 - 0x0
      13'h1C97: dout  = 8'b11100000; // 7319 : 224 - 0xe0
      13'h1C98: dout  = 8'b00000000; // 7320 :   0 - 0x0
      13'h1C99: dout  = 8'b00000000; // 7321 :   0 - 0x0
      13'h1C9A: dout  = 8'b00000000; // 7322 :   0 - 0x0
      13'h1C9B: dout  = 8'b00000000; // 7323 :   0 - 0x0
      13'h1C9C: dout  = 8'b10000000; // 7324 : 128 - 0x80
      13'h1C9D: dout  = 8'b11000000; // 7325 : 192 - 0xc0
      13'h1C9E: dout  = 8'b11000000; // 7326 : 192 - 0xc0
      13'h1C9F: dout  = 8'b11110000; // 7327 : 240 - 0xf0
      13'h1CA0: dout  = 8'b01110000; // 7328 : 112 - 0x70 -- Background 0xca
      13'h1CA1: dout  = 8'b01111100; // 7329 : 124 - 0x7c
      13'h1CA2: dout  = 8'b01111110; // 7330 : 126 - 0x7e
      13'h1CA3: dout  = 8'b11111111; // 7331 : 255 - 0xff
      13'h1CA4: dout  = 8'b11111111; // 7332 : 255 - 0xff
      13'h1CA5: dout  = 8'b11110111; // 7333 : 247 - 0xf7
      13'h1CA6: dout  = 8'b11101111; // 7334 : 239 - 0xef
      13'h1CA7: dout  = 8'b00011111; // 7335 :  31 - 0x1f
      13'h1CA8: dout  = 8'b11111100; // 7336 : 252 - 0xfc
      13'h1CA9: dout  = 8'b11111110; // 7337 : 254 - 0xfe
      13'h1CAA: dout  = 8'b11111111; // 7338 : 255 - 0xff
      13'h1CAB: dout  = 8'b11111111; // 7339 : 255 - 0xff
      13'h1CAC: dout  = 8'b11111111; // 7340 : 255 - 0xff
      13'h1CAD: dout  = 8'b11111111; // 7341 : 255 - 0xff
      13'h1CAE: dout  = 8'b11111111; // 7342 : 255 - 0xff
      13'h1CAF: dout  = 8'b11111111; // 7343 : 255 - 0xff
      13'h1CB0: dout  = 8'b11111111; // 7344 : 255 - 0xff -- Background 0xcb
      13'h1CB1: dout  = 8'b11111111; // 7345 : 255 - 0xff
      13'h1CB2: dout  = 8'b11111111; // 7346 : 255 - 0xff
      13'h1CB3: dout  = 8'b11111000; // 7347 : 248 - 0xf8
      13'h1CB4: dout  = 8'b11111000; // 7348 : 248 - 0xf8
      13'h1CB5: dout  = 8'b11111110; // 7349 : 254 - 0xfe
      13'h1CB6: dout  = 8'b11111111; // 7350 : 255 - 0xff
      13'h1CB7: dout  = 8'b11111111; // 7351 : 255 - 0xff
      13'h1CB8: dout  = 8'b11111111; // 7352 : 255 - 0xff
      13'h1CB9: dout  = 8'b11111111; // 7353 : 255 - 0xff
      13'h1CBA: dout  = 8'b11111111; // 7354 : 255 - 0xff
      13'h1CBB: dout  = 8'b11111000; // 7355 : 248 - 0xf8
      13'h1CBC: dout  = 8'b11111110; // 7356 : 254 - 0xfe
      13'h1CBD: dout  = 8'b11111111; // 7357 : 255 - 0xff
      13'h1CBE: dout  = 8'b11111111; // 7358 : 255 - 0xff
      13'h1CBF: dout  = 8'b11111111; // 7359 : 255 - 0xff
      13'h1CC0: dout  = 8'b11111111; // 7360 : 255 - 0xff -- Background 0xcc
      13'h1CC1: dout  = 8'b11111111; // 7361 : 255 - 0xff
      13'h1CC2: dout  = 8'b11111111; // 7362 : 255 - 0xff
      13'h1CC3: dout  = 8'b00111111; // 7363 :  63 - 0x3f
      13'h1CC4: dout  = 8'b00011110; // 7364 :  30 - 0x1e
      13'h1CC5: dout  = 8'b00000001; // 7365 :   1 - 0x1
      13'h1CC6: dout  = 8'b00000000; // 7366 :   0 - 0x0
      13'h1CC7: dout  = 8'b00000000; // 7367 :   0 - 0x0
      13'h1CC8: dout  = 8'b11111111; // 7368 : 255 - 0xff
      13'h1CC9: dout  = 8'b11111111; // 7369 : 255 - 0xff
      13'h1CCA: dout  = 8'b11111111; // 7370 : 255 - 0xff
      13'h1CCB: dout  = 8'b00111111; // 7371 :  63 - 0x3f
      13'h1CCC: dout  = 8'b00011111; // 7372 :  31 - 0x1f
      13'h1CCD: dout  = 8'b00011111; // 7373 :  31 - 0x1f
      13'h1CCE: dout  = 8'b00000000; // 7374 :   0 - 0x0
      13'h1CCF: dout  = 8'b00000000; // 7375 :   0 - 0x0
      13'h1CD0: dout  = 8'b00000000; // 7376 :   0 - 0x0 -- Background 0xcd
      13'h1CD1: dout  = 8'b00000000; // 7377 :   0 - 0x0
      13'h1CD2: dout  = 8'b00000000; // 7378 :   0 - 0x0
      13'h1CD3: dout  = 8'b10000000; // 7379 : 128 - 0x80
      13'h1CD4: dout  = 8'b11000000; // 7380 : 192 - 0xc0
      13'h1CD5: dout  = 8'b11100000; // 7381 : 224 - 0xe0
      13'h1CD6: dout  = 8'b11100000; // 7382 : 224 - 0xe0
      13'h1CD7: dout  = 8'b11100000; // 7383 : 224 - 0xe0
      13'h1CD8: dout  = 8'b00000000; // 7384 :   0 - 0x0
      13'h1CD9: dout  = 8'b00000000; // 7385 :   0 - 0x0
      13'h1CDA: dout  = 8'b10000000; // 7386 : 128 - 0x80
      13'h1CDB: dout  = 8'b11000000; // 7387 : 192 - 0xc0
      13'h1CDC: dout  = 8'b11100000; // 7388 : 224 - 0xe0
      13'h1CDD: dout  = 8'b11100000; // 7389 : 224 - 0xe0
      13'h1CDE: dout  = 8'b11100000; // 7390 : 224 - 0xe0
      13'h1CDF: dout  = 8'b11100000; // 7391 : 224 - 0xe0
      13'h1CE0: dout  = 8'b11000000; // 7392 : 192 - 0xc0 -- Background 0xce
      13'h1CE1: dout  = 8'b10000000; // 7393 : 128 - 0x80
      13'h1CE2: dout  = 8'b00000000; // 7394 :   0 - 0x0
      13'h1CE3: dout  = 8'b00000000; // 7395 :   0 - 0x0
      13'h1CE4: dout  = 8'b00000000; // 7396 :   0 - 0x0
      13'h1CE5: dout  = 8'b00000000; // 7397 :   0 - 0x0
      13'h1CE6: dout  = 8'b10000000; // 7398 : 128 - 0x80
      13'h1CE7: dout  = 8'b10000000; // 7399 : 128 - 0x80
      13'h1CE8: dout  = 8'b11000000; // 7400 : 192 - 0xc0
      13'h1CE9: dout  = 8'b10000000; // 7401 : 128 - 0x80
      13'h1CEA: dout  = 8'b00000000; // 7402 :   0 - 0x0
      13'h1CEB: dout  = 8'b00000000; // 7403 :   0 - 0x0
      13'h1CEC: dout  = 8'b00000000; // 7404 :   0 - 0x0
      13'h1CED: dout  = 8'b10000000; // 7405 : 128 - 0x80
      13'h1CEE: dout  = 8'b11000000; // 7406 : 192 - 0xc0
      13'h1CEF: dout  = 8'b11000000; // 7407 : 192 - 0xc0
      13'h1CF0: dout  = 8'b10000000; // 7408 : 128 - 0x80 -- Background 0xcf
      13'h1CF1: dout  = 8'b10000000; // 7409 : 128 - 0x80
      13'h1CF2: dout  = 8'b11100000; // 7410 : 224 - 0xe0
      13'h1CF3: dout  = 8'b11000000; // 7411 : 192 - 0xc0
      13'h1CF4: dout  = 8'b00100000; // 7412 :  32 - 0x20
      13'h1CF5: dout  = 8'b00000000; // 7413 :   0 - 0x0
      13'h1CF6: dout  = 8'b00000000; // 7414 :   0 - 0x0
      13'h1CF7: dout  = 8'b00000000; // 7415 :   0 - 0x0
      13'h1CF8: dout  = 8'b11000000; // 7416 : 192 - 0xc0
      13'h1CF9: dout  = 8'b11000000; // 7417 : 192 - 0xc0
      13'h1CFA: dout  = 8'b11100000; // 7418 : 224 - 0xe0
      13'h1CFB: dout  = 8'b11111000; // 7419 : 248 - 0xf8
      13'h1CFC: dout  = 8'b11111100; // 7420 : 252 - 0xfc
      13'h1CFD: dout  = 8'b11111100; // 7421 : 252 - 0xfc
      13'h1CFE: dout  = 8'b00000000; // 7422 :   0 - 0x0
      13'h1CFF: dout  = 8'b00000000; // 7423 :   0 - 0x0
      13'h1D00: dout  = 8'b00011111; // 7424 :  31 - 0x1f -- Background 0xd0
      13'h1D01: dout  = 8'b00000110; // 7425 :   6 - 0x6
      13'h1D02: dout  = 8'b00000110; // 7426 :   6 - 0x6
      13'h1D03: dout  = 8'b00000110; // 7427 :   6 - 0x6
      13'h1D04: dout  = 8'b00000110; // 7428 :   6 - 0x6
      13'h1D05: dout  = 8'b00000110; // 7429 :   6 - 0x6
      13'h1D06: dout  = 8'b00000110; // 7430 :   6 - 0x6
      13'h1D07: dout  = 8'b00000000; // 7431 :   0 - 0x0
      13'h1D08: dout  = 8'b00000000; // 7432 :   0 - 0x0
      13'h1D09: dout  = 8'b00000000; // 7433 :   0 - 0x0
      13'h1D0A: dout  = 8'b00000000; // 7434 :   0 - 0x0
      13'h1D0B: dout  = 8'b00000000; // 7435 :   0 - 0x0
      13'h1D0C: dout  = 8'b00000000; // 7436 :   0 - 0x0
      13'h1D0D: dout  = 8'b00000000; // 7437 :   0 - 0x0
      13'h1D0E: dout  = 8'b00000000; // 7438 :   0 - 0x0
      13'h1D0F: dout  = 8'b00000000; // 7439 :   0 - 0x0
      13'h1D10: dout  = 8'b00111001; // 7440 :  57 - 0x39 -- Background 0xd1
      13'h1D11: dout  = 8'b01100101; // 7441 : 101 - 0x65
      13'h1D12: dout  = 8'b01100101; // 7442 : 101 - 0x65
      13'h1D13: dout  = 8'b01100101; // 7443 : 101 - 0x65
      13'h1D14: dout  = 8'b01100101; // 7444 : 101 - 0x65
      13'h1D15: dout  = 8'b01100101; // 7445 : 101 - 0x65
      13'h1D16: dout  = 8'b00111001; // 7446 :  57 - 0x39
      13'h1D17: dout  = 8'b00000000; // 7447 :   0 - 0x0
      13'h1D18: dout  = 8'b00000000; // 7448 :   0 - 0x0
      13'h1D19: dout  = 8'b00000000; // 7449 :   0 - 0x0
      13'h1D1A: dout  = 8'b00000000; // 7450 :   0 - 0x0
      13'h1D1B: dout  = 8'b00000000; // 7451 :   0 - 0x0
      13'h1D1C: dout  = 8'b00000000; // 7452 :   0 - 0x0
      13'h1D1D: dout  = 8'b00000000; // 7453 :   0 - 0x0
      13'h1D1E: dout  = 8'b00000000; // 7454 :   0 - 0x0
      13'h1D1F: dout  = 8'b00000000; // 7455 :   0 - 0x0
      13'h1D20: dout  = 8'b11100000; // 7456 : 224 - 0xe0 -- Background 0xd2
      13'h1D21: dout  = 8'b10110000; // 7457 : 176 - 0xb0
      13'h1D22: dout  = 8'b10110000; // 7458 : 176 - 0xb0
      13'h1D23: dout  = 8'b10110110; // 7459 : 182 - 0xb6
      13'h1D24: dout  = 8'b11100110; // 7460 : 230 - 0xe6
      13'h1D25: dout  = 8'b10000000; // 7461 : 128 - 0x80
      13'h1D26: dout  = 8'b10000000; // 7462 : 128 - 0x80
      13'h1D27: dout  = 8'b00000000; // 7463 :   0 - 0x0
      13'h1D28: dout  = 8'b00000000; // 7464 :   0 - 0x0
      13'h1D29: dout  = 8'b00000000; // 7465 :   0 - 0x0
      13'h1D2A: dout  = 8'b00000000; // 7466 :   0 - 0x0
      13'h1D2B: dout  = 8'b00000000; // 7467 :   0 - 0x0
      13'h1D2C: dout  = 8'b00000000; // 7468 :   0 - 0x0
      13'h1D2D: dout  = 8'b00000000; // 7469 :   0 - 0x0
      13'h1D2E: dout  = 8'b00000000; // 7470 :   0 - 0x0
      13'h1D2F: dout  = 8'b00000000; // 7471 :   0 - 0x0
      13'h1D30: dout  = 8'b00111100; // 7472 :  60 - 0x3c -- Background 0xd3
      13'h1D31: dout  = 8'b01000010; // 7473 :  66 - 0x42
      13'h1D32: dout  = 8'b10011001; // 7474 : 153 - 0x99
      13'h1D33: dout  = 8'b10100001; // 7475 : 161 - 0xa1
      13'h1D34: dout  = 8'b10100001; // 7476 : 161 - 0xa1
      13'h1D35: dout  = 8'b10011001; // 7477 : 153 - 0x99
      13'h1D36: dout  = 8'b01000010; // 7478 :  66 - 0x42
      13'h1D37: dout  = 8'b00111100; // 7479 :  60 - 0x3c
      13'h1D38: dout  = 8'b00000000; // 7480 :   0 - 0x0
      13'h1D39: dout  = 8'b00000000; // 7481 :   0 - 0x0
      13'h1D3A: dout  = 8'b00000000; // 7482 :   0 - 0x0
      13'h1D3B: dout  = 8'b00000000; // 7483 :   0 - 0x0
      13'h1D3C: dout  = 8'b00000000; // 7484 :   0 - 0x0
      13'h1D3D: dout  = 8'b00000000; // 7485 :   0 - 0x0
      13'h1D3E: dout  = 8'b00000000; // 7486 :   0 - 0x0
      13'h1D3F: dout  = 8'b00000000; // 7487 :   0 - 0x0
      13'h1D40: dout  = 8'b00000000; // 7488 :   0 - 0x0 -- Background 0xd4
      13'h1D41: dout  = 8'b00000000; // 7489 :   0 - 0x0
      13'h1D42: dout  = 8'b00000000; // 7490 :   0 - 0x0
      13'h1D43: dout  = 8'b00000011; // 7491 :   3 - 0x3
      13'h1D44: dout  = 8'b00000110; // 7492 :   6 - 0x6
      13'h1D45: dout  = 8'b00000000; // 7493 :   0 - 0x0
      13'h1D46: dout  = 8'b00000001; // 7494 :   1 - 0x1
      13'h1D47: dout  = 8'b00000111; // 7495 :   7 - 0x7
      13'h1D48: dout  = 8'b00000000; // 7496 :   0 - 0x0
      13'h1D49: dout  = 8'b00000000; // 7497 :   0 - 0x0
      13'h1D4A: dout  = 8'b00000000; // 7498 :   0 - 0x0
      13'h1D4B: dout  = 8'b00000000; // 7499 :   0 - 0x0
      13'h1D4C: dout  = 8'b00000011; // 7500 :   3 - 0x3
      13'h1D4D: dout  = 8'b00000111; // 7501 :   7 - 0x7
      13'h1D4E: dout  = 8'b00000011; // 7502 :   3 - 0x3
      13'h1D4F: dout  = 8'b00000111; // 7503 :   7 - 0x7
      13'h1D50: dout  = 8'b00001111; // 7504 :  15 - 0xf -- Background 0xd5
      13'h1D51: dout  = 8'b00011111; // 7505 :  31 - 0x1f
      13'h1D52: dout  = 8'b00111111; // 7506 :  63 - 0x3f
      13'h1D53: dout  = 8'b01111111; // 7507 : 127 - 0x7f
      13'h1D54: dout  = 8'b01111111; // 7508 : 127 - 0x7f
      13'h1D55: dout  = 8'b01111111; // 7509 : 127 - 0x7f
      13'h1D56: dout  = 8'b11111111; // 7510 : 255 - 0xff
      13'h1D57: dout  = 8'b01111111; // 7511 : 127 - 0x7f
      13'h1D58: dout  = 8'b00011111; // 7512 :  31 - 0x1f
      13'h1D59: dout  = 8'b00111111; // 7513 :  63 - 0x3f
      13'h1D5A: dout  = 8'b01111111; // 7514 : 127 - 0x7f
      13'h1D5B: dout  = 8'b11111111; // 7515 : 255 - 0xff
      13'h1D5C: dout  = 8'b11111111; // 7516 : 255 - 0xff
      13'h1D5D: dout  = 8'b11111111; // 7517 : 255 - 0xff
      13'h1D5E: dout  = 8'b11111111; // 7518 : 255 - 0xff
      13'h1D5F: dout  = 8'b01111111; // 7519 : 127 - 0x7f
      13'h1D60: dout  = 8'b00000000; // 7520 :   0 - 0x0 -- Background 0xd6
      13'h1D61: dout  = 8'b00000000; // 7521 :   0 - 0x0
      13'h1D62: dout  = 8'b00000000; // 7522 :   0 - 0x0
      13'h1D63: dout  = 8'b10000000; // 7523 : 128 - 0x80
      13'h1D64: dout  = 8'b00000000; // 7524 :   0 - 0x0
      13'h1D65: dout  = 8'b00000000; // 7525 :   0 - 0x0
      13'h1D66: dout  = 8'b00000000; // 7526 :   0 - 0x0
      13'h1D67: dout  = 8'b10100000; // 7527 : 160 - 0xa0
      13'h1D68: dout  = 8'b00000000; // 7528 :   0 - 0x0
      13'h1D69: dout  = 8'b00000000; // 7529 :   0 - 0x0
      13'h1D6A: dout  = 8'b00000000; // 7530 :   0 - 0x0
      13'h1D6B: dout  = 8'b11000000; // 7531 : 192 - 0xc0
      13'h1D6C: dout  = 8'b11100000; // 7532 : 224 - 0xe0
      13'h1D6D: dout  = 8'b11110000; // 7533 : 240 - 0xf0
      13'h1D6E: dout  = 8'b11110000; // 7534 : 240 - 0xf0
      13'h1D6F: dout  = 8'b11111000; // 7535 : 248 - 0xf8
      13'h1D70: dout  = 8'b11100000; // 7536 : 224 - 0xe0 -- Background 0xd7
      13'h1D71: dout  = 8'b11110000; // 7537 : 240 - 0xf0
      13'h1D72: dout  = 8'b11100000; // 7538 : 224 - 0xe0
      13'h1D73: dout  = 8'b11011101; // 7539 : 221 - 0xdd
      13'h1D74: dout  = 8'b11111010; // 7540 : 250 - 0xfa
      13'h1D75: dout  = 8'b11101011; // 7541 : 235 - 0xeb
      13'h1D76: dout  = 8'b10000000; // 7542 : 128 - 0x80
      13'h1D77: dout  = 8'b00000000; // 7543 :   0 - 0x0
      13'h1D78: dout  = 8'b11111100; // 7544 : 252 - 0xfc
      13'h1D79: dout  = 8'b11111000; // 7545 : 248 - 0xf8
      13'h1D7A: dout  = 8'b11110000; // 7546 : 240 - 0xf0
      13'h1D7B: dout  = 8'b11111111; // 7547 : 255 - 0xff
      13'h1D7C: dout  = 8'b11111111; // 7548 : 255 - 0xff
      13'h1D7D: dout  = 8'b11111111; // 7549 : 255 - 0xff
      13'h1D7E: dout  = 8'b11111111; // 7550 : 255 - 0xff
      13'h1D7F: dout  = 8'b11111111; // 7551 : 255 - 0xff
      13'h1D80: dout  = 8'b00000000; // 7552 :   0 - 0x0 -- Background 0xd8
      13'h1D81: dout  = 8'b00000000; // 7553 :   0 - 0x0
      13'h1D82: dout  = 8'b00000000; // 7554 :   0 - 0x0
      13'h1D83: dout  = 8'b00000011; // 7555 :   3 - 0x3
      13'h1D84: dout  = 8'b00000110; // 7556 :   6 - 0x6
      13'h1D85: dout  = 8'b00000000; // 7557 :   0 - 0x0
      13'h1D86: dout  = 8'b00000001; // 7558 :   1 - 0x1
      13'h1D87: dout  = 8'b00000001; // 7559 :   1 - 0x1
      13'h1D88: dout  = 8'b00000000; // 7560 :   0 - 0x0
      13'h1D89: dout  = 8'b00000000; // 7561 :   0 - 0x0
      13'h1D8A: dout  = 8'b00000000; // 7562 :   0 - 0x0
      13'h1D8B: dout  = 8'b00000000; // 7563 :   0 - 0x0
      13'h1D8C: dout  = 8'b00000011; // 7564 :   3 - 0x3
      13'h1D8D: dout  = 8'b00000111; // 7565 :   7 - 0x7
      13'h1D8E: dout  = 8'b00001111; // 7566 :  15 - 0xf
      13'h1D8F: dout  = 8'b00011111; // 7567 :  31 - 0x1f
      13'h1D90: dout  = 8'b00001011; // 7568 :  11 - 0xb -- Background 0xd9
      13'h1D91: dout  = 8'b00000111; // 7569 :   7 - 0x7
      13'h1D92: dout  = 8'b00000011; // 7570 :   3 - 0x3
      13'h1D93: dout  = 8'b01011101; // 7571 :  93 - 0x5d
      13'h1D94: dout  = 8'b10101111; // 7572 : 175 - 0xaf
      13'h1D95: dout  = 8'b01010011; // 7573 :  83 - 0x53
      13'h1D96: dout  = 8'b00000000; // 7574 :   0 - 0x0
      13'h1D97: dout  = 8'b00000000; // 7575 :   0 - 0x0
      13'h1D98: dout  = 8'b00111111; // 7576 :  63 - 0x3f
      13'h1D99: dout  = 8'b00011111; // 7577 :  31 - 0x1f
      13'h1D9A: dout  = 8'b00000111; // 7578 :   7 - 0x7
      13'h1D9B: dout  = 8'b11111111; // 7579 : 255 - 0xff
      13'h1D9C: dout  = 8'b11111111; // 7580 : 255 - 0xff
      13'h1D9D: dout  = 8'b11111111; // 7581 : 255 - 0xff
      13'h1D9E: dout  = 8'b11111111; // 7582 : 255 - 0xff
      13'h1D9F: dout  = 8'b11111111; // 7583 : 255 - 0xff
      13'h1DA0: dout  = 8'b00000000; // 7584 :   0 - 0x0 -- Background 0xda
      13'h1DA1: dout  = 8'b00000000; // 7585 :   0 - 0x0
      13'h1DA2: dout  = 8'b00000000; // 7586 :   0 - 0x0
      13'h1DA3: dout  = 8'b10000000; // 7587 : 128 - 0x80
      13'h1DA4: dout  = 8'b00000000; // 7588 :   0 - 0x0
      13'h1DA5: dout  = 8'b00000000; // 7589 :   0 - 0x0
      13'h1DA6: dout  = 8'b01100000; // 7590 :  96 - 0x60
      13'h1DA7: dout  = 8'b11110000; // 7591 : 240 - 0xf0
      13'h1DA8: dout  = 8'b00000000; // 7592 :   0 - 0x0
      13'h1DA9: dout  = 8'b00000000; // 7593 :   0 - 0x0
      13'h1DAA: dout  = 8'b00000000; // 7594 :   0 - 0x0
      13'h1DAB: dout  = 8'b11000000; // 7595 : 192 - 0xc0
      13'h1DAC: dout  = 8'b11000000; // 7596 : 192 - 0xc0
      13'h1DAD: dout  = 8'b11000000; // 7597 : 192 - 0xc0
      13'h1DAE: dout  = 8'b11100000; // 7598 : 224 - 0xe0
      13'h1DAF: dout  = 8'b11111000; // 7599 : 248 - 0xf8
      13'h1DB0: dout  = 8'b11111000; // 7600 : 248 - 0xf8 -- Background 0xdb
      13'h1DB1: dout  = 8'b11111100; // 7601 : 252 - 0xfc
      13'h1DB2: dout  = 8'b11111100; // 7602 : 252 - 0xfc
      13'h1DB3: dout  = 8'b11111110; // 7603 : 254 - 0xfe
      13'h1DB4: dout  = 8'b11111110; // 7604 : 254 - 0xfe
      13'h1DB5: dout  = 8'b11111111; // 7605 : 255 - 0xff
      13'h1DB6: dout  = 8'b11111111; // 7606 : 255 - 0xff
      13'h1DB7: dout  = 8'b01111110; // 7607 : 126 - 0x7e
      13'h1DB8: dout  = 8'b11111100; // 7608 : 252 - 0xfc
      13'h1DB9: dout  = 8'b11111110; // 7609 : 254 - 0xfe
      13'h1DBA: dout  = 8'b11111110; // 7610 : 254 - 0xfe
      13'h1DBB: dout  = 8'b11111111; // 7611 : 255 - 0xff
      13'h1DBC: dout  = 8'b11111111; // 7612 : 255 - 0xff
      13'h1DBD: dout  = 8'b11111111; // 7613 : 255 - 0xff
      13'h1DBE: dout  = 8'b11111111; // 7614 : 255 - 0xff
      13'h1DBF: dout  = 8'b11111110; // 7615 : 254 - 0xfe
      13'h1DC0: dout  = 8'b00000000; // 7616 :   0 - 0x0 -- Background 0xdc
      13'h1DC1: dout  = 8'b00000000; // 7617 :   0 - 0x0
      13'h1DC2: dout  = 8'b00000000; // 7618 :   0 - 0x0
      13'h1DC3: dout  = 8'b00000000; // 7619 :   0 - 0x0
      13'h1DC4: dout  = 8'b00000000; // 7620 :   0 - 0x0
      13'h1DC5: dout  = 8'b00000000; // 7621 :   0 - 0x0
      13'h1DC6: dout  = 8'b00100001; // 7622 :  33 - 0x21
      13'h1DC7: dout  = 8'b00111111; // 7623 :  63 - 0x3f
      13'h1DC8: dout  = 8'b00110110; // 7624 :  54 - 0x36
      13'h1DC9: dout  = 8'b00110110; // 7625 :  54 - 0x36
      13'h1DCA: dout  = 8'b01111110; // 7626 : 126 - 0x7e
      13'h1DCB: dout  = 8'b01111111; // 7627 : 127 - 0x7f
      13'h1DCC: dout  = 8'b01111111; // 7628 : 127 - 0x7f
      13'h1DCD: dout  = 8'b01111111; // 7629 : 127 - 0x7f
      13'h1DCE: dout  = 8'b00111111; // 7630 :  63 - 0x3f
      13'h1DCF: dout  = 8'b00111111; // 7631 :  63 - 0x3f
      13'h1DD0: dout  = 8'b00111111; // 7632 :  63 - 0x3f -- Background 0xdd
      13'h1DD1: dout  = 8'b00011111; // 7633 :  31 - 0x1f
      13'h1DD2: dout  = 8'b00011111; // 7634 :  31 - 0x1f
      13'h1DD3: dout  = 8'b00001111; // 7635 :  15 - 0xf
      13'h1DD4: dout  = 8'b00000111; // 7636 :   7 - 0x7
      13'h1DD5: dout  = 8'b00000011; // 7637 :   3 - 0x3
      13'h1DD6: dout  = 8'b00000000; // 7638 :   0 - 0x0
      13'h1DD7: dout  = 8'b00000000; // 7639 :   0 - 0x0
      13'h1DD8: dout  = 8'b00111111; // 7640 :  63 - 0x3f
      13'h1DD9: dout  = 8'b00011111; // 7641 :  31 - 0x1f
      13'h1DDA: dout  = 8'b00011111; // 7642 :  31 - 0x1f
      13'h1DDB: dout  = 8'b00001111; // 7643 :  15 - 0xf
      13'h1DDC: dout  = 8'b00000111; // 7644 :   7 - 0x7
      13'h1DDD: dout  = 8'b00000011; // 7645 :   3 - 0x3
      13'h1DDE: dout  = 8'b00000000; // 7646 :   0 - 0x0
      13'h1DDF: dout  = 8'b00000000; // 7647 :   0 - 0x0
      13'h1DE0: dout  = 8'b00111110; // 7648 :  62 - 0x3e -- Background 0xde
      13'h1DE1: dout  = 8'b00011110; // 7649 :  30 - 0x1e
      13'h1DE2: dout  = 8'b00011110; // 7650 :  30 - 0x1e
      13'h1DE3: dout  = 8'b00001110; // 7651 :  14 - 0xe
      13'h1DE4: dout  = 8'b00001111; // 7652 :  15 - 0xf
      13'h1DE5: dout  = 8'b00011111; // 7653 :  31 - 0x1f
      13'h1DE6: dout  = 8'b10011111; // 7654 : 159 - 0x9f
      13'h1DE7: dout  = 8'b10011111; // 7655 : 159 - 0x9f
      13'h1DE8: dout  = 8'b00111111; // 7656 :  63 - 0x3f
      13'h1DE9: dout  = 8'b00011111; // 7657 :  31 - 0x1f
      13'h1DEA: dout  = 8'b11011111; // 7658 : 223 - 0xdf
      13'h1DEB: dout  = 8'b11001111; // 7659 : 207 - 0xcf
      13'h1DEC: dout  = 8'b11001111; // 7660 : 207 - 0xcf
      13'h1DED: dout  = 8'b10011111; // 7661 : 159 - 0x9f
      13'h1DEE: dout  = 8'b11011111; // 7662 : 223 - 0xdf
      13'h1DEF: dout  = 8'b11111111; // 7663 : 255 - 0xff
      13'h1DF0: dout  = 8'b11011111; // 7664 : 223 - 0xdf -- Background 0xdf
      13'h1DF1: dout  = 8'b11111111; // 7665 : 255 - 0xff
      13'h1DF2: dout  = 8'b11111111; // 7666 : 255 - 0xff
      13'h1DF3: dout  = 8'b11111111; // 7667 : 255 - 0xff
      13'h1DF4: dout  = 8'b11111111; // 7668 : 255 - 0xff
      13'h1DF5: dout  = 8'b11011111; // 7669 : 223 - 0xdf
      13'h1DF6: dout  = 8'b11100111; // 7670 : 231 - 0xe7
      13'h1DF7: dout  = 8'b00000000; // 7671 :   0 - 0x0
      13'h1DF8: dout  = 8'b11111111; // 7672 : 255 - 0xff
      13'h1DF9: dout  = 8'b11111111; // 7673 : 255 - 0xff
      13'h1DFA: dout  = 8'b11111111; // 7674 : 255 - 0xff
      13'h1DFB: dout  = 8'b11111111; // 7675 : 255 - 0xff
      13'h1DFC: dout  = 8'b11111111; // 7676 : 255 - 0xff
      13'h1DFD: dout  = 8'b11111111; // 7677 : 255 - 0xff
      13'h1DFE: dout  = 8'b11111111; // 7678 : 255 - 0xff
      13'h1DFF: dout  = 8'b00001111; // 7679 :  15 - 0xf
      13'h1E00: dout  = 8'b00100000; // 7680 :  32 - 0x20 -- Background 0xe0
      13'h1E01: dout  = 8'b00001111; // 7681 :  15 - 0xf
      13'h1E02: dout  = 8'b00110000; // 7682 :  48 - 0x30
      13'h1E03: dout  = 8'b01000000; // 7683 :  64 - 0x40
      13'h1E04: dout  = 8'b10011000; // 7684 : 152 - 0x98
      13'h1E05: dout  = 8'b00111110; // 7685 :  62 - 0x3e
      13'h1E06: dout  = 8'b00011111; // 7686 :  31 - 0x1f
      13'h1E07: dout  = 8'b00000000; // 7687 :   0 - 0x0
      13'h1E08: dout  = 8'b11111111; // 7688 : 255 - 0xff
      13'h1E09: dout  = 8'b11111111; // 7689 : 255 - 0xff
      13'h1E0A: dout  = 8'b11111111; // 7690 : 255 - 0xff
      13'h1E0B: dout  = 8'b11111111; // 7691 : 255 - 0xff
      13'h1E0C: dout  = 8'b11111111; // 7692 : 255 - 0xff
      13'h1E0D: dout  = 8'b11111111; // 7693 : 255 - 0xff
      13'h1E0E: dout  = 8'b11111111; // 7694 : 255 - 0xff
      13'h1E0F: dout  = 8'b11111111; // 7695 : 255 - 0xff
      13'h1E10: dout  = 8'b10000001; // 7696 : 129 - 0x81 -- Background 0xe1
      13'h1E11: dout  = 8'b00110110; // 7697 :  54 - 0x36
      13'h1E12: dout  = 8'b00101110; // 7698 :  46 - 0x2e
      13'h1E13: dout  = 8'b10101111; // 7699 : 175 - 0xaf
      13'h1E14: dout  = 8'b10101110; // 7700 : 174 - 0xae
      13'h1E15: dout  = 8'b11010001; // 7701 : 209 - 0xd1
      13'h1E16: dout  = 8'b11101111; // 7702 : 239 - 0xef
      13'h1E17: dout  = 8'b10000111; // 7703 : 135 - 0x87
      13'h1E18: dout  = 8'b11111111; // 7704 : 255 - 0xff
      13'h1E19: dout  = 8'b11111001; // 7705 : 249 - 0xf9
      13'h1E1A: dout  = 8'b11110000; // 7706 : 240 - 0xf0
      13'h1E1B: dout  = 8'b11110000; // 7707 : 240 - 0xf0
      13'h1E1C: dout  = 8'b10110001; // 7708 : 177 - 0xb1
      13'h1E1D: dout  = 8'b11011111; // 7709 : 223 - 0xdf
      13'h1E1E: dout  = 8'b11101111; // 7710 : 239 - 0xef
      13'h1E1F: dout  = 8'b10000111; // 7711 : 135 - 0x87
      13'h1E20: dout  = 8'b00000010; // 7712 :   2 - 0x2 -- Background 0xe2
      13'h1E21: dout  = 8'b11111000; // 7713 : 248 - 0xf8
      13'h1E22: dout  = 8'b00000110; // 7714 :   6 - 0x6
      13'h1E23: dout  = 8'b00000001; // 7715 :   1 - 0x1
      13'h1E24: dout  = 8'b00001100; // 7716 :  12 - 0xc
      13'h1E25: dout  = 8'b00111110; // 7717 :  62 - 0x3e
      13'h1E26: dout  = 8'b11111100; // 7718 : 252 - 0xfc
      13'h1E27: dout  = 8'b00000000; // 7719 :   0 - 0x0
      13'h1E28: dout  = 8'b11111111; // 7720 : 255 - 0xff
      13'h1E29: dout  = 8'b11111111; // 7721 : 255 - 0xff
      13'h1E2A: dout  = 8'b11111111; // 7722 : 255 - 0xff
      13'h1E2B: dout  = 8'b11111111; // 7723 : 255 - 0xff
      13'h1E2C: dout  = 8'b11111111; // 7724 : 255 - 0xff
      13'h1E2D: dout  = 8'b11111111; // 7725 : 255 - 0xff
      13'h1E2E: dout  = 8'b11111111; // 7726 : 255 - 0xff
      13'h1E2F: dout  = 8'b11111111; // 7727 : 255 - 0xff
      13'h1E30: dout  = 8'b11000000; // 7728 : 192 - 0xc0 -- Background 0xe3
      13'h1E31: dout  = 8'b00110110; // 7729 :  54 - 0x36
      13'h1E32: dout  = 8'b00111110; // 7730 :  62 - 0x3e
      13'h1E33: dout  = 8'b01111010; // 7731 : 122 - 0x7a
      13'h1E34: dout  = 8'b10110110; // 7732 : 182 - 0xb6
      13'h1E35: dout  = 8'b11001101; // 7733 : 205 - 0xcd
      13'h1E36: dout  = 8'b11111011; // 7734 : 251 - 0xfb
      13'h1E37: dout  = 8'b11110000; // 7735 : 240 - 0xf0
      13'h1E38: dout  = 8'b11111111; // 7736 : 255 - 0xff
      13'h1E39: dout  = 8'b11001111; // 7737 : 207 - 0xcf
      13'h1E3A: dout  = 8'b10000111; // 7738 : 135 - 0x87
      13'h1E3B: dout  = 8'b10000111; // 7739 : 135 - 0x87
      13'h1E3C: dout  = 8'b11001110; // 7740 : 206 - 0xce
      13'h1E3D: dout  = 8'b11111101; // 7741 : 253 - 0xfd
      13'h1E3E: dout  = 8'b11111011; // 7742 : 251 - 0xfb
      13'h1E3F: dout  = 8'b11110000; // 7743 : 240 - 0xf0
      13'h1E40: dout  = 8'b00111110; // 7744 :  62 - 0x3e -- Background 0xe4
      13'h1E41: dout  = 8'b00111100; // 7745 :  60 - 0x3c
      13'h1E42: dout  = 8'b00111100; // 7746 :  60 - 0x3c
      13'h1E43: dout  = 8'b00111000; // 7747 :  56 - 0x38
      13'h1E44: dout  = 8'b11111000; // 7748 : 248 - 0xf8
      13'h1E45: dout  = 8'b01111100; // 7749 : 124 - 0x7c
      13'h1E46: dout  = 8'b01111110; // 7750 : 126 - 0x7e
      13'h1E47: dout  = 8'b01111000; // 7751 : 120 - 0x78
      13'h1E48: dout  = 8'b11111110; // 7752 : 254 - 0xfe
      13'h1E49: dout  = 8'b11111100; // 7753 : 252 - 0xfc
      13'h1E4A: dout  = 8'b11111100; // 7754 : 252 - 0xfc
      13'h1E4B: dout  = 8'b11111000; // 7755 : 248 - 0xf8
      13'h1E4C: dout  = 8'b11111011; // 7756 : 251 - 0xfb
      13'h1E4D: dout  = 8'b11111101; // 7757 : 253 - 0xfd
      13'h1E4E: dout  = 8'b11111110; // 7758 : 254 - 0xfe
      13'h1E4F: dout  = 8'b11111111; // 7759 : 255 - 0xff
      13'h1E50: dout  = 8'b11111000; // 7760 : 248 - 0xf8 -- Background 0xe5
      13'h1E51: dout  = 8'b01111111; // 7761 : 127 - 0x7f
      13'h1E52: dout  = 8'b01111111; // 7762 : 127 - 0x7f
      13'h1E53: dout  = 8'b11111110; // 7763 : 254 - 0xfe
      13'h1E54: dout  = 8'b11111111; // 7764 : 255 - 0xff
      13'h1E55: dout  = 8'b11111111; // 7765 : 255 - 0xff
      13'h1E56: dout  = 8'b11110011; // 7766 : 243 - 0xf3
      13'h1E57: dout  = 8'b10000001; // 7767 : 129 - 0x81
      13'h1E58: dout  = 8'b11111111; // 7768 : 255 - 0xff
      13'h1E59: dout  = 8'b11111111; // 7769 : 255 - 0xff
      13'h1E5A: dout  = 8'b11111111; // 7770 : 255 - 0xff
      13'h1E5B: dout  = 8'b11111111; // 7771 : 255 - 0xff
      13'h1E5C: dout  = 8'b11111111; // 7772 : 255 - 0xff
      13'h1E5D: dout  = 8'b11111111; // 7773 : 255 - 0xff
      13'h1E5E: dout  = 8'b11111111; // 7774 : 255 - 0xff
      13'h1E5F: dout  = 8'b11111001; // 7775 : 249 - 0xf9
      13'h1E60: dout  = 8'b00000000; // 7776 :   0 - 0x0 -- Background 0xe6
      13'h1E61: dout  = 8'b00000000; // 7777 :   0 - 0x0
      13'h1E62: dout  = 8'b00000000; // 7778 :   0 - 0x0
      13'h1E63: dout  = 8'b00010000; // 7779 :  16 - 0x10
      13'h1E64: dout  = 8'b01000000; // 7780 :  64 - 0x40
      13'h1E65: dout  = 8'b00100000; // 7781 :  32 - 0x20
      13'h1E66: dout  = 8'b00000000; // 7782 :   0 - 0x0
      13'h1E67: dout  = 8'b00000000; // 7783 :   0 - 0x0
      13'h1E68: dout  = 8'b00000000; // 7784 :   0 - 0x0
      13'h1E69: dout  = 8'b00000000; // 7785 :   0 - 0x0
      13'h1E6A: dout  = 8'b00000000; // 7786 :   0 - 0x0
      13'h1E6B: dout  = 8'b01111000; // 7787 : 120 - 0x78
      13'h1E6C: dout  = 8'b11111100; // 7788 : 252 - 0xfc
      13'h1E6D: dout  = 8'b11111100; // 7789 : 252 - 0xfc
      13'h1E6E: dout  = 8'b11111100; // 7790 : 252 - 0xfc
      13'h1E6F: dout  = 8'b11111100; // 7791 : 252 - 0xfc
      13'h1E70: dout  = 8'b00000110; // 7792 :   6 - 0x6 -- Background 0xe7
      13'h1E71: dout  = 8'b00001110; // 7793 :  14 - 0xe
      13'h1E72: dout  = 8'b01111110; // 7794 : 126 - 0x7e
      13'h1E73: dout  = 8'b11111110; // 7795 : 254 - 0xfe
      13'h1E74: dout  = 8'b11111110; // 7796 : 254 - 0xfe
      13'h1E75: dout  = 8'b11111100; // 7797 : 252 - 0xfc
      13'h1E76: dout  = 8'b11111000; // 7798 : 248 - 0xf8
      13'h1E77: dout  = 8'b11110000; // 7799 : 240 - 0xf0
      13'h1E78: dout  = 8'b11111110; // 7800 : 254 - 0xfe
      13'h1E79: dout  = 8'b11111110; // 7801 : 254 - 0xfe
      13'h1E7A: dout  = 8'b11111110; // 7802 : 254 - 0xfe
      13'h1E7B: dout  = 8'b11111110; // 7803 : 254 - 0xfe
      13'h1E7C: dout  = 8'b11111110; // 7804 : 254 - 0xfe
      13'h1E7D: dout  = 8'b11111100; // 7805 : 252 - 0xfc
      13'h1E7E: dout  = 8'b11111000; // 7806 : 248 - 0xf8
      13'h1E7F: dout  = 8'b11110000; // 7807 : 240 - 0xf0
      13'h1E80: dout  = 8'b00000000; // 7808 :   0 - 0x0 -- Background 0xe8
      13'h1E81: dout  = 8'b00000000; // 7809 :   0 - 0x0
      13'h1E82: dout  = 8'b00000000; // 7810 :   0 - 0x0
      13'h1E83: dout  = 8'b00000000; // 7811 :   0 - 0x0
      13'h1E84: dout  = 8'b00000000; // 7812 :   0 - 0x0
      13'h1E85: dout  = 8'b00000000; // 7813 :   0 - 0x0
      13'h1E86: dout  = 8'b00000000; // 7814 :   0 - 0x0
      13'h1E87: dout  = 8'b00000001; // 7815 :   1 - 0x1
      13'h1E88: dout  = 8'b00000000; // 7816 :   0 - 0x0
      13'h1E89: dout  = 8'b00000000; // 7817 :   0 - 0x0
      13'h1E8A: dout  = 8'b00000000; // 7818 :   0 - 0x0
      13'h1E8B: dout  = 8'b00000000; // 7819 :   0 - 0x0
      13'h1E8C: dout  = 8'b00000000; // 7820 :   0 - 0x0
      13'h1E8D: dout  = 8'b00000000; // 7821 :   0 - 0x0
      13'h1E8E: dout  = 8'b00000000; // 7822 :   0 - 0x0
      13'h1E8F: dout  = 8'b00000000; // 7823 :   0 - 0x0
      13'h1E90: dout  = 8'b00000010; // 7824 :   2 - 0x2 -- Background 0xe9
      13'h1E91: dout  = 8'b00000000; // 7825 :   0 - 0x0
      13'h1E92: dout  = 8'b00001000; // 7826 :   8 - 0x8
      13'h1E93: dout  = 8'b00000001; // 7827 :   1 - 0x1
      13'h1E94: dout  = 8'b00010011; // 7828 :  19 - 0x13
      13'h1E95: dout  = 8'b00000001; // 7829 :   1 - 0x1
      13'h1E96: dout  = 8'b00000000; // 7830 :   0 - 0x0
      13'h1E97: dout  = 8'b00000000; // 7831 :   0 - 0x0
      13'h1E98: dout  = 8'b00000001; // 7832 :   1 - 0x1
      13'h1E99: dout  = 8'b00001111; // 7833 :  15 - 0xf
      13'h1E9A: dout  = 8'b00011111; // 7834 :  31 - 0x1f
      13'h1E9B: dout  = 8'b00011111; // 7835 :  31 - 0x1f
      13'h1E9C: dout  = 8'b00111011; // 7836 :  59 - 0x3b
      13'h1E9D: dout  = 8'b00110011; // 7837 :  51 - 0x33
      13'h1E9E: dout  = 8'b00000001; // 7838 :   1 - 0x1
      13'h1E9F: dout  = 8'b00000001; // 7839 :   1 - 0x1
      13'h1EA0: dout  = 8'b00000000; // 7840 :   0 - 0x0 -- Background 0xea
      13'h1EA1: dout  = 8'b00000000; // 7841 :   0 - 0x0
      13'h1EA2: dout  = 8'b00000000; // 7842 :   0 - 0x0
      13'h1EA3: dout  = 8'b00000000; // 7843 :   0 - 0x0
      13'h1EA4: dout  = 8'b00000000; // 7844 :   0 - 0x0
      13'h1EA5: dout  = 8'b00000000; // 7845 :   0 - 0x0
      13'h1EA6: dout  = 8'b00000000; // 7846 :   0 - 0x0
      13'h1EA7: dout  = 8'b00000000; // 7847 :   0 - 0x0
      13'h1EA8: dout  = 8'b00000000; // 7848 :   0 - 0x0
      13'h1EA9: dout  = 8'b00000000; // 7849 :   0 - 0x0
      13'h1EAA: dout  = 8'b00000000; // 7850 :   0 - 0x0
      13'h1EAB: dout  = 8'b00110110; // 7851 :  54 - 0x36
      13'h1EAC: dout  = 8'b01101100; // 7852 : 108 - 0x6c
      13'h1EAD: dout  = 8'b11111101; // 7853 : 253 - 0xfd
      13'h1EAE: dout  = 8'b11111111; // 7854 : 255 - 0xff
      13'h1EAF: dout  = 8'b11111111; // 7855 : 255 - 0xff
      13'h1EB0: dout  = 8'b00000000; // 7856 :   0 - 0x0 -- Background 0xeb
      13'h1EB1: dout  = 8'b01000011; // 7857 :  67 - 0x43
      13'h1EB2: dout  = 8'b01111111; // 7858 : 127 - 0x7f
      13'h1EB3: dout  = 8'b01111111; // 7859 : 127 - 0x7f
      13'h1EB4: dout  = 8'b01111111; // 7860 : 127 - 0x7f
      13'h1EB5: dout  = 8'b00111111; // 7861 :  63 - 0x3f
      13'h1EB6: dout  = 8'b00011111; // 7862 :  31 - 0x1f
      13'h1EB7: dout  = 8'b00000111; // 7863 :   7 - 0x7
      13'h1EB8: dout  = 8'b11111111; // 7864 : 255 - 0xff
      13'h1EB9: dout  = 8'b01111111; // 7865 : 127 - 0x7f
      13'h1EBA: dout  = 8'b01111111; // 7866 : 127 - 0x7f
      13'h1EBB: dout  = 8'b01111111; // 7867 : 127 - 0x7f
      13'h1EBC: dout  = 8'b01111111; // 7868 : 127 - 0x7f
      13'h1EBD: dout  = 8'b00111111; // 7869 :  63 - 0x3f
      13'h1EBE: dout  = 8'b00011111; // 7870 :  31 - 0x1f
      13'h1EBF: dout  = 8'b00000111; // 7871 :   7 - 0x7
      13'h1EC0: dout  = 8'b00000000; // 7872 :   0 - 0x0 -- Background 0xec
      13'h1EC1: dout  = 8'b00000000; // 7873 :   0 - 0x0
      13'h1EC2: dout  = 8'b00000000; // 7874 :   0 - 0x0
      13'h1EC3: dout  = 8'b00000000; // 7875 :   0 - 0x0
      13'h1EC4: dout  = 8'b00000000; // 7876 :   0 - 0x0
      13'h1EC5: dout  = 8'b00000000; // 7877 :   0 - 0x0
      13'h1EC6: dout  = 8'b11000000; // 7878 : 192 - 0xc0
      13'h1EC7: dout  = 8'b00000000; // 7879 :   0 - 0x0
      13'h1EC8: dout  = 8'b00000000; // 7880 :   0 - 0x0
      13'h1EC9: dout  = 8'b00000000; // 7881 :   0 - 0x0
      13'h1ECA: dout  = 8'b00000000; // 7882 :   0 - 0x0
      13'h1ECB: dout  = 8'b00000000; // 7883 :   0 - 0x0
      13'h1ECC: dout  = 8'b00000000; // 7884 :   0 - 0x0
      13'h1ECD: dout  = 8'b00000000; // 7885 :   0 - 0x0
      13'h1ECE: dout  = 8'b00000000; // 7886 :   0 - 0x0
      13'h1ECF: dout  = 8'b11100000; // 7887 : 224 - 0xe0
      13'h1ED0: dout  = 8'b00010000; // 7888 :  16 - 0x10 -- Background 0xed
      13'h1ED1: dout  = 8'b00111000; // 7889 :  56 - 0x38
      13'h1ED2: dout  = 8'b10111111; // 7890 : 191 - 0xbf
      13'h1ED3: dout  = 8'b11111111; // 7891 : 255 - 0xff
      13'h1ED4: dout  = 8'b11111111; // 7892 : 255 - 0xff
      13'h1ED5: dout  = 8'b11111111; // 7893 : 255 - 0xff
      13'h1ED6: dout  = 8'b11111111; // 7894 : 255 - 0xff
      13'h1ED7: dout  = 8'b11111111; // 7895 : 255 - 0xff
      13'h1ED8: dout  = 8'b11111000; // 7896 : 248 - 0xf8
      13'h1ED9: dout  = 8'b11111111; // 7897 : 255 - 0xff
      13'h1EDA: dout  = 8'b11111111; // 7898 : 255 - 0xff
      13'h1EDB: dout  = 8'b11111111; // 7899 : 255 - 0xff
      13'h1EDC: dout  = 8'b11111111; // 7900 : 255 - 0xff
      13'h1EDD: dout  = 8'b11111111; // 7901 : 255 - 0xff
      13'h1EDE: dout  = 8'b11111111; // 7902 : 255 - 0xff
      13'h1EDF: dout  = 8'b11111111; // 7903 : 255 - 0xff
      13'h1EE0: dout  = 8'b01111110; // 7904 : 126 - 0x7e -- Background 0xee
      13'h1EE1: dout  = 8'b00011110; // 7905 :  30 - 0x1e
      13'h1EE2: dout  = 8'b00011110; // 7906 :  30 - 0x1e
      13'h1EE3: dout  = 8'b00001110; // 7907 :  14 - 0xe
      13'h1EE4: dout  = 8'b00001111; // 7908 :  15 - 0xf
      13'h1EE5: dout  = 8'b00011110; // 7909 :  30 - 0x1e
      13'h1EE6: dout  = 8'b00011110; // 7910 :  30 - 0x1e
      13'h1EE7: dout  = 8'b00111110; // 7911 :  62 - 0x3e
      13'h1EE8: dout  = 8'b11111111; // 7912 : 255 - 0xff
      13'h1EE9: dout  = 8'b01111111; // 7913 : 127 - 0x7f
      13'h1EEA: dout  = 8'b00011111; // 7914 :  31 - 0x1f
      13'h1EEB: dout  = 8'b00001111; // 7915 :  15 - 0xf
      13'h1EEC: dout  = 8'b00001111; // 7916 :  15 - 0xf
      13'h1EED: dout  = 8'b10011111; // 7917 : 159 - 0x9f
      13'h1EEE: dout  = 8'b10011111; // 7918 : 159 - 0x9f
      13'h1EEF: dout  = 8'b10111111; // 7919 : 191 - 0xbf
      13'h1EF0: dout  = 8'b01111111; // 7920 : 127 - 0x7f -- Background 0xef
      13'h1EF1: dout  = 8'b01111111; // 7921 : 127 - 0x7f
      13'h1EF2: dout  = 8'b10111111; // 7922 : 191 - 0xbf
      13'h1EF3: dout  = 8'b11111111; // 7923 : 255 - 0xff
      13'h1EF4: dout  = 8'b11111111; // 7924 : 255 - 0xff
      13'h1EF5: dout  = 8'b11111111; // 7925 : 255 - 0xff
      13'h1EF6: dout  = 8'b11100111; // 7926 : 231 - 0xe7
      13'h1EF7: dout  = 8'b11000000; // 7927 : 192 - 0xc0
      13'h1EF8: dout  = 8'b01111111; // 7928 : 127 - 0x7f
      13'h1EF9: dout  = 8'b11111111; // 7929 : 255 - 0xff
      13'h1EFA: dout  = 8'b11111111; // 7930 : 255 - 0xff
      13'h1EFB: dout  = 8'b11111111; // 7931 : 255 - 0xff
      13'h1EFC: dout  = 8'b11111111; // 7932 : 255 - 0xff
      13'h1EFD: dout  = 8'b11111111; // 7933 : 255 - 0xff
      13'h1EFE: dout  = 8'b11111111; // 7934 : 255 - 0xff
      13'h1EFF: dout  = 8'b11001111; // 7935 : 207 - 0xcf
      13'h1F00: dout  = 8'b00000000; // 7936 :   0 - 0x0 -- Background 0xf0
      13'h1F01: dout  = 8'b00000000; // 7937 :   0 - 0x0
      13'h1F02: dout  = 8'b00010000; // 7938 :  16 - 0x10
      13'h1F03: dout  = 8'b11111101; // 7939 : 253 - 0xfd
      13'h1F04: dout  = 8'b11111010; // 7940 : 250 - 0xfa
      13'h1F05: dout  = 8'b11101011; // 7941 : 235 - 0xeb
      13'h1F06: dout  = 8'b10000000; // 7942 : 128 - 0x80
      13'h1F07: dout  = 8'b00000000; // 7943 :   0 - 0x0
      13'h1F08: dout  = 8'b00000000; // 7944 :   0 - 0x0
      13'h1F09: dout  = 8'b00000000; // 7945 :   0 - 0x0
      13'h1F0A: dout  = 8'b11110000; // 7946 : 240 - 0xf0
      13'h1F0B: dout  = 8'b11111111; // 7947 : 255 - 0xff
      13'h1F0C: dout  = 8'b11111111; // 7948 : 255 - 0xff
      13'h1F0D: dout  = 8'b11111111; // 7949 : 255 - 0xff
      13'h1F0E: dout  = 8'b11111111; // 7950 : 255 - 0xff
      13'h1F0F: dout  = 8'b11111111; // 7951 : 255 - 0xff
      13'h1F10: dout  = 8'b00100000; // 7952 :  32 - 0x20 -- Background 0xf1
      13'h1F11: dout  = 8'b00011111; // 7953 :  31 - 0x1f
      13'h1F12: dout  = 8'b01100000; // 7954 :  96 - 0x60
      13'h1F13: dout  = 8'b10001110; // 7955 : 142 - 0x8e
      13'h1F14: dout  = 8'b00111111; // 7956 :  63 - 0x3f
      13'h1F15: dout  = 8'b01111111; // 7957 : 127 - 0x7f
      13'h1F16: dout  = 8'b01111111; // 7958 : 127 - 0x7f
      13'h1F17: dout  = 8'b01111100; // 7959 : 124 - 0x7c
      13'h1F18: dout  = 8'b11111111; // 7960 : 255 - 0xff
      13'h1F19: dout  = 8'b11111111; // 7961 : 255 - 0xff
      13'h1F1A: dout  = 8'b11111111; // 7962 : 255 - 0xff
      13'h1F1B: dout  = 8'b11110001; // 7963 : 241 - 0xf1
      13'h1F1C: dout  = 8'b11000100; // 7964 : 196 - 0xc4
      13'h1F1D: dout  = 8'b11101110; // 7965 : 238 - 0xee
      13'h1F1E: dout  = 8'b11000100; // 7966 : 196 - 0xc4
      13'h1F1F: dout  = 8'b10000011; // 7967 : 131 - 0x83
      13'h1F20: dout  = 8'b00111001; // 7968 :  57 - 0x39 -- Background 0xf2
      13'h1F21: dout  = 8'b00110110; // 7969 :  54 - 0x36
      13'h1F22: dout  = 8'b00101110; // 7970 :  46 - 0x2e
      13'h1F23: dout  = 8'b10101111; // 7971 : 175 - 0xaf
      13'h1F24: dout  = 8'b10101110; // 7972 : 174 - 0xae
      13'h1F25: dout  = 8'b11010001; // 7973 : 209 - 0xd1
      13'h1F26: dout  = 8'b11101111; // 7974 : 239 - 0xef
      13'h1F27: dout  = 8'b10000111; // 7975 : 135 - 0x87
      13'h1F28: dout  = 8'b11000111; // 7976 : 199 - 0xc7
      13'h1F29: dout  = 8'b11111001; // 7977 : 249 - 0xf9
      13'h1F2A: dout  = 8'b11110000; // 7978 : 240 - 0xf0
      13'h1F2B: dout  = 8'b11110000; // 7979 : 240 - 0xf0
      13'h1F2C: dout  = 8'b10110001; // 7980 : 177 - 0xb1
      13'h1F2D: dout  = 8'b11011111; // 7981 : 223 - 0xdf
      13'h1F2E: dout  = 8'b11101111; // 7982 : 239 - 0xef
      13'h1F2F: dout  = 8'b10000111; // 7983 : 135 - 0x87
      13'h1F30: dout  = 8'b00000000; // 7984 :   0 - 0x0 -- Background 0xf3
      13'h1F31: dout  = 8'b00000000; // 7985 :   0 - 0x0
      13'h1F32: dout  = 8'b00000100; // 7986 :   4 - 0x4
      13'h1F33: dout  = 8'b01011111; // 7987 :  95 - 0x5f
      13'h1F34: dout  = 8'b10101111; // 7988 : 175 - 0xaf
      13'h1F35: dout  = 8'b01010011; // 7989 :  83 - 0x53
      13'h1F36: dout  = 8'b00000000; // 7990 :   0 - 0x0
      13'h1F37: dout  = 8'b00000000; // 7991 :   0 - 0x0
      13'h1F38: dout  = 8'b00000000; // 7992 :   0 - 0x0
      13'h1F39: dout  = 8'b00000000; // 7993 :   0 - 0x0
      13'h1F3A: dout  = 8'b00000111; // 7994 :   7 - 0x7
      13'h1F3B: dout  = 8'b11111111; // 7995 : 255 - 0xff
      13'h1F3C: dout  = 8'b11111111; // 7996 : 255 - 0xff
      13'h1F3D: dout  = 8'b11111111; // 7997 : 255 - 0xff
      13'h1F3E: dout  = 8'b11111111; // 7998 : 255 - 0xff
      13'h1F3F: dout  = 8'b11111111; // 7999 : 255 - 0xff
      13'h1F40: dout  = 8'b00000010; // 8000 :   2 - 0x2 -- Background 0xf4
      13'h1F41: dout  = 8'b11111100; // 8001 : 252 - 0xfc
      13'h1F42: dout  = 8'b00000011; // 8002 :   3 - 0x3
      13'h1F43: dout  = 8'b00111000; // 8003 :  56 - 0x38
      13'h1F44: dout  = 8'b11111110; // 8004 : 254 - 0xfe
      13'h1F45: dout  = 8'b11111111; // 8005 : 255 - 0xff
      13'h1F46: dout  = 8'b11111111; // 8006 : 255 - 0xff
      13'h1F47: dout  = 8'b00011110; // 8007 :  30 - 0x1e
      13'h1F48: dout  = 8'b11111111; // 8008 : 255 - 0xff
      13'h1F49: dout  = 8'b11111111; // 8009 : 255 - 0xff
      13'h1F4A: dout  = 8'b11111111; // 8010 : 255 - 0xff
      13'h1F4B: dout  = 8'b11000111; // 8011 : 199 - 0xc7
      13'h1F4C: dout  = 8'b01000101; // 8012 :  69 - 0x45
      13'h1F4D: dout  = 8'b11101110; // 8013 : 238 - 0xee
      13'h1F4E: dout  = 8'b01000100; // 8014 :  68 - 0x44
      13'h1F4F: dout  = 8'b11100001; // 8015 : 225 - 0xe1
      13'h1F50: dout  = 8'b11000000; // 8016 : 192 - 0xc0 -- Background 0xf5
      13'h1F51: dout  = 8'b00110110; // 8017 :  54 - 0x36
      13'h1F52: dout  = 8'b00111110; // 8018 :  62 - 0x3e
      13'h1F53: dout  = 8'b01111010; // 8019 : 122 - 0x7a
      13'h1F54: dout  = 8'b10110110; // 8020 : 182 - 0xb6
      13'h1F55: dout  = 8'b11001101; // 8021 : 205 - 0xcd
      13'h1F56: dout  = 8'b11111011; // 8022 : 251 - 0xfb
      13'h1F57: dout  = 8'b11110000; // 8023 : 240 - 0xf0
      13'h1F58: dout  = 8'b11111111; // 8024 : 255 - 0xff
      13'h1F59: dout  = 8'b11001111; // 8025 : 207 - 0xcf
      13'h1F5A: dout  = 8'b10000111; // 8026 : 135 - 0x87
      13'h1F5B: dout  = 8'b10000111; // 8027 : 135 - 0x87
      13'h1F5C: dout  = 8'b11001110; // 8028 : 206 - 0xce
      13'h1F5D: dout  = 8'b11111101; // 8029 : 253 - 0xfd
      13'h1F5E: dout  = 8'b11111011; // 8030 : 251 - 0xfb
      13'h1F5F: dout  = 8'b11110000; // 8031 : 240 - 0xf0
      13'h1F60: dout  = 8'b00000000; // 8032 :   0 - 0x0 -- Background 0xf6
      13'h1F61: dout  = 8'b00000000; // 8033 :   0 - 0x0
      13'h1F62: dout  = 8'b00000000; // 8034 :   0 - 0x0
      13'h1F63: dout  = 8'b00000000; // 8035 :   0 - 0x0
      13'h1F64: dout  = 8'b00000000; // 8036 :   0 - 0x0
      13'h1F65: dout  = 8'b00001110; // 8037 :  14 - 0xe
      13'h1F66: dout  = 8'b00001000; // 8038 :   8 - 0x8
      13'h1F67: dout  = 8'b00001000; // 8039 :   8 - 0x8
      13'h1F68: dout  = 8'b00000000; // 8040 :   0 - 0x0
      13'h1F69: dout  = 8'b00000000; // 8041 :   0 - 0x0
      13'h1F6A: dout  = 8'b00000000; // 8042 :   0 - 0x0
      13'h1F6B: dout  = 8'b00000000; // 8043 :   0 - 0x0
      13'h1F6C: dout  = 8'b00000000; // 8044 :   0 - 0x0
      13'h1F6D: dout  = 8'b00000001; // 8045 :   1 - 0x1
      13'h1F6E: dout  = 8'b00000111; // 8046 :   7 - 0x7
      13'h1F6F: dout  = 8'b00001111; // 8047 :  15 - 0xf
      13'h1F70: dout  = 8'b00011111; // 8048 :  31 - 0x1f -- Background 0xf7
      13'h1F71: dout  = 8'b00111111; // 8049 :  63 - 0x3f
      13'h1F72: dout  = 8'b11111111; // 8050 : 255 - 0xff
      13'h1F73: dout  = 8'b11111111; // 8051 : 255 - 0xff
      13'h1F74: dout  = 8'b11111111; // 8052 : 255 - 0xff
      13'h1F75: dout  = 8'b11111111; // 8053 : 255 - 0xff
      13'h1F76: dout  = 8'b11111111; // 8054 : 255 - 0xff
      13'h1F77: dout  = 8'b01111111; // 8055 : 127 - 0x7f
      13'h1F78: dout  = 8'b00111111; // 8056 :  63 - 0x3f
      13'h1F79: dout  = 8'b11111111; // 8057 : 255 - 0xff
      13'h1F7A: dout  = 8'b11111111; // 8058 : 255 - 0xff
      13'h1F7B: dout  = 8'b11111111; // 8059 : 255 - 0xff
      13'h1F7C: dout  = 8'b11111111; // 8060 : 255 - 0xff
      13'h1F7D: dout  = 8'b11111111; // 8061 : 255 - 0xff
      13'h1F7E: dout  = 8'b11111111; // 8062 : 255 - 0xff
      13'h1F7F: dout  = 8'b11111111; // 8063 : 255 - 0xff
      13'h1F80: dout  = 8'b00111111; // 8064 :  63 - 0x3f -- Background 0xf8
      13'h1F81: dout  = 8'b00111110; // 8065 :  62 - 0x3e
      13'h1F82: dout  = 8'b00111100; // 8066 :  60 - 0x3c
      13'h1F83: dout  = 8'b10111000; // 8067 : 184 - 0xb8
      13'h1F84: dout  = 8'b01111000; // 8068 : 120 - 0x78
      13'h1F85: dout  = 8'b01111000; // 8069 : 120 - 0x78
      13'h1F86: dout  = 8'b01111110; // 8070 : 126 - 0x7e
      13'h1F87: dout  = 8'b01111110; // 8071 : 126 - 0x7e
      13'h1F88: dout  = 8'b11111111; // 8072 : 255 - 0xff
      13'h1F89: dout  = 8'b11111111; // 8073 : 255 - 0xff
      13'h1F8A: dout  = 8'b11111101; // 8074 : 253 - 0xfd
      13'h1F8B: dout  = 8'b11111000; // 8075 : 248 - 0xf8
      13'h1F8C: dout  = 8'b11111111; // 8076 : 255 - 0xff
      13'h1F8D: dout  = 8'b11111111; // 8077 : 255 - 0xff
      13'h1F8E: dout  = 8'b11111110; // 8078 : 254 - 0xfe
      13'h1F8F: dout  = 8'b11111111; // 8079 : 255 - 0xff
      13'h1F90: dout  = 8'b11111101; // 8080 : 253 - 0xfd -- Background 0xf9
      13'h1F91: dout  = 8'b01111001; // 8081 : 121 - 0x79
      13'h1F92: dout  = 8'b01111011; // 8082 : 123 - 0x7b
      13'h1F93: dout  = 8'b11111111; // 8083 : 255 - 0xff
      13'h1F94: dout  = 8'b11111111; // 8084 : 255 - 0xff
      13'h1F95: dout  = 8'b11111111; // 8085 : 255 - 0xff
      13'h1F96: dout  = 8'b11110011; // 8086 : 243 - 0xf3
      13'h1F97: dout  = 8'b10000000; // 8087 : 128 - 0x80
      13'h1F98: dout  = 8'b11111111; // 8088 : 255 - 0xff
      13'h1F99: dout  = 8'b11111111; // 8089 : 255 - 0xff
      13'h1F9A: dout  = 8'b11111111; // 8090 : 255 - 0xff
      13'h1F9B: dout  = 8'b11111111; // 8091 : 255 - 0xff
      13'h1F9C: dout  = 8'b11111111; // 8092 : 255 - 0xff
      13'h1F9D: dout  = 8'b11111111; // 8093 : 255 - 0xff
      13'h1F9E: dout  = 8'b11111111; // 8094 : 255 - 0xff
      13'h1F9F: dout  = 8'b11111000; // 8095 : 248 - 0xf8
      13'h1FA0: dout  = 8'b00000000; // 8096 :   0 - 0x0 -- Background 0xfa
      13'h1FA1: dout  = 8'b00000000; // 8097 :   0 - 0x0
      13'h1FA2: dout  = 8'b00000000; // 8098 :   0 - 0x0
      13'h1FA3: dout  = 8'b00000000; // 8099 :   0 - 0x0
      13'h1FA4: dout  = 8'b00000000; // 8100 :   0 - 0x0
      13'h1FA5: dout  = 8'b00000000; // 8101 :   0 - 0x0
      13'h1FA6: dout  = 8'b00000000; // 8102 :   0 - 0x0
      13'h1FA7: dout  = 8'b00000000; // 8103 :   0 - 0x0
      13'h1FA8: dout  = 8'b00000000; // 8104 :   0 - 0x0
      13'h1FA9: dout  = 8'b00000000; // 8105 :   0 - 0x0
      13'h1FAA: dout  = 8'b00000000; // 8106 :   0 - 0x0
      13'h1FAB: dout  = 8'b00000000; // 8107 :   0 - 0x0
      13'h1FAC: dout  = 8'b00000000; // 8108 :   0 - 0x0
      13'h1FAD: dout  = 8'b00000000; // 8109 :   0 - 0x0
      13'h1FAE: dout  = 8'b11000000; // 8110 : 192 - 0xc0
      13'h1FAF: dout  = 8'b11110000; // 8111 : 240 - 0xf0
      13'h1FB0: dout  = 8'b00010000; // 8112 :  16 - 0x10 -- Background 0xfb
      13'h1FB1: dout  = 8'b10000100; // 8113 : 132 - 0x84
      13'h1FB2: dout  = 8'b11100000; // 8114 : 224 - 0xe0
      13'h1FB3: dout  = 8'b11000000; // 8115 : 192 - 0xc0
      13'h1FB4: dout  = 8'b10000000; // 8116 : 128 - 0x80
      13'h1FB5: dout  = 8'b10000000; // 8117 : 128 - 0x80
      13'h1FB6: dout  = 8'b00000000; // 8118 :   0 - 0x0
      13'h1FB7: dout  = 8'b00000000; // 8119 :   0 - 0x0
      13'h1FB8: dout  = 8'b11111100; // 8120 : 252 - 0xfc
      13'h1FB9: dout  = 8'b11111110; // 8121 : 254 - 0xfe
      13'h1FBA: dout  = 8'b11101100; // 8122 : 236 - 0xec
      13'h1FBB: dout  = 8'b11100000; // 8123 : 224 - 0xe0
      13'h1FBC: dout  = 8'b11000000; // 8124 : 192 - 0xc0
      13'h1FBD: dout  = 8'b11000000; // 8125 : 192 - 0xc0
      13'h1FBE: dout  = 8'b10000000; // 8126 : 128 - 0x80
      13'h1FBF: dout  = 8'b10000000; // 8127 : 128 - 0x80
      13'h1FC0: dout  = 8'b00000000; // 8128 :   0 - 0x0 -- Background 0xfc
      13'h1FC1: dout  = 8'b01001000; // 8129 :  72 - 0x48
      13'h1FC2: dout  = 8'b00100000; // 8130 :  32 - 0x20
      13'h1FC3: dout  = 8'b00000000; // 8131 :   0 - 0x0
      13'h1FC4: dout  = 8'b00000000; // 8132 :   0 - 0x0
      13'h1FC5: dout  = 8'b00000100; // 8133 :   4 - 0x4
      13'h1FC6: dout  = 8'b00001110; // 8134 :  14 - 0xe
      13'h1FC7: dout  = 8'b11111110; // 8135 : 254 - 0xfe
      13'h1FC8: dout  = 8'b01110000; // 8136 : 112 - 0x70
      13'h1FC9: dout  = 8'b11111100; // 8137 : 252 - 0xfc
      13'h1FCA: dout  = 8'b11111100; // 8138 : 252 - 0xfc
      13'h1FCB: dout  = 8'b11111100; // 8139 : 252 - 0xfc
      13'h1FCC: dout  = 8'b11111100; // 8140 : 252 - 0xfc
      13'h1FCD: dout  = 8'b11111100; // 8141 : 252 - 0xfc
      13'h1FCE: dout  = 8'b11111110; // 8142 : 254 - 0xfe
      13'h1FCF: dout  = 8'b11111110; // 8143 : 254 - 0xfe
      13'h1FD0: dout  = 8'b11111110; // 8144 : 254 - 0xfe -- Background 0xfd
      13'h1FD1: dout  = 8'b11111100; // 8145 : 252 - 0xfc
      13'h1FD2: dout  = 8'b11111100; // 8146 : 252 - 0xfc
      13'h1FD3: dout  = 8'b11111000; // 8147 : 248 - 0xf8
      13'h1FD4: dout  = 8'b11110000; // 8148 : 240 - 0xf0
      13'h1FD5: dout  = 8'b11100000; // 8149 : 224 - 0xe0
      13'h1FD6: dout  = 8'b10000000; // 8150 : 128 - 0x80
      13'h1FD7: dout  = 8'b00000000; // 8151 :   0 - 0x0
      13'h1FD8: dout  = 8'b11111110; // 8152 : 254 - 0xfe
      13'h1FD9: dout  = 8'b11111100; // 8153 : 252 - 0xfc
      13'h1FDA: dout  = 8'b11111100; // 8154 : 252 - 0xfc
      13'h1FDB: dout  = 8'b11111000; // 8155 : 248 - 0xf8
      13'h1FDC: dout  = 8'b11110000; // 8156 : 240 - 0xf0
      13'h1FDD: dout  = 8'b11100000; // 8157 : 224 - 0xe0
      13'h1FDE: dout  = 8'b10000000; // 8158 : 128 - 0x80
      13'h1FDF: dout  = 8'b00000000; // 8159 :   0 - 0x0
      13'h1FE0: dout  = 8'b00001111; // 8160 :  15 - 0xf -- Background 0xfe
      13'h1FE1: dout  = 8'b00000110; // 8161 :   6 - 0x6
      13'h1FE2: dout  = 8'b00000110; // 8162 :   6 - 0x6
      13'h1FE3: dout  = 8'b00000110; // 8163 :   6 - 0x6
      13'h1FE4: dout  = 8'b00000110; // 8164 :   6 - 0x6
      13'h1FE5: dout  = 8'b00000110; // 8165 :   6 - 0x6
      13'h1FE6: dout  = 8'b00001111; // 8166 :  15 - 0xf
      13'h1FE7: dout  = 8'b00000000; // 8167 :   0 - 0x0
      13'h1FE8: dout  = 8'b00000000; // 8168 :   0 - 0x0
      13'h1FE9: dout  = 8'b00000000; // 8169 :   0 - 0x0
      13'h1FEA: dout  = 8'b00000000; // 8170 :   0 - 0x0
      13'h1FEB: dout  = 8'b00000000; // 8171 :   0 - 0x0
      13'h1FEC: dout  = 8'b00000000; // 8172 :   0 - 0x0
      13'h1FED: dout  = 8'b00000000; // 8173 :   0 - 0x0
      13'h1FEE: dout  = 8'b00000000; // 8174 :   0 - 0x0
      13'h1FEF: dout  = 8'b00000000; // 8175 :   0 - 0x0
      13'h1FF0: dout  = 8'b11110000; // 8176 : 240 - 0xf0 -- Background 0xff
      13'h1FF1: dout  = 8'b01100000; // 8177 :  96 - 0x60
      13'h1FF2: dout  = 8'b01100000; // 8178 :  96 - 0x60
      13'h1FF3: dout  = 8'b01100110; // 8179 : 102 - 0x66
      13'h1FF4: dout  = 8'b01100110; // 8180 : 102 - 0x66
      13'h1FF5: dout  = 8'b01100000; // 8181 :  96 - 0x60
      13'h1FF6: dout  = 8'b11110000; // 8182 : 240 - 0xf0
      13'h1FF7: dout  = 8'b00000000; // 8183 :   0 - 0x0
      13'h1FF8: dout  = 8'b00000000; // 8184 :   0 - 0x0
      13'h1FF9: dout  = 8'b00000000; // 8185 :   0 - 0x0
      13'h1FFA: dout  = 8'b00000000; // 8186 :   0 - 0x0
      13'h1FFB: dout  = 8'b00000000; // 8187 :   0 - 0x0
      13'h1FFC: dout  = 8'b00000000; // 8188 :   0 - 0x0
      13'h1FFD: dout  = 8'b00000000; // 8189 :   0 - 0x0
      13'h1FFE: dout  = 8'b00000000; // 8190 :   0 - 0x0
      13'h1FFF: dout  = 8'b00000000; // 8191 :   0 - 0x0
    endcase
  end

endmodule
