--- Autcmatically generated VHDL ROM from a NES memory file----
---   NAME TABLE
-- https://wiki.nesdev.com/w/index.php/PPU_nametables


---  Original memory dump file name: lawnmower_ntable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory with clock ------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_NTABLE_LAWN_00 is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(11-1 downto 0);  --2048 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_NTABLE_LAWN_00;

architecture BEHAVIORAL of ROM_NTABLE_LAWN_00 is
  signal addr_int  : natural range 0 to 2**11-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
     ------- Name Table 0---------
    "10101001", --    0 -  0x0  :  169 - 0xa9 -- line 0x0
    "10101001", --    1 -  0x1  :  169 - 0xa9
    "10101001", --    2 -  0x2  :  169 - 0xa9
    "10101001", --    3 -  0x3  :  169 - 0xa9
    "10101001", --    4 -  0x4  :  169 - 0xa9
    "10101001", --    5 -  0x5  :  169 - 0xa9
    "10101001", --    6 -  0x6  :  169 - 0xa9
    "10101001", --    7 -  0x7  :  169 - 0xa9
    "10101001", --    8 -  0x8  :  169 - 0xa9
    "10101001", --    9 -  0x9  :  169 - 0xa9
    "10101001", --   10 -  0xa  :  169 - 0xa9
    "10101001", --   11 -  0xb  :  169 - 0xa9
    "10101001", --   12 -  0xc  :  169 - 0xa9
    "10101001", --   13 -  0xd  :  169 - 0xa9
    "10101001", --   14 -  0xe  :  169 - 0xa9
    "10101001", --   15 -  0xf  :  169 - 0xa9
    "10101001", --   16 - 0x10  :  169 - 0xa9
    "10101001", --   17 - 0x11  :  169 - 0xa9
    "10101001", --   18 - 0x12  :  169 - 0xa9
    "10101001", --   19 - 0x13  :  169 - 0xa9
    "10101001", --   20 - 0x14  :  169 - 0xa9
    "10101001", --   21 - 0x15  :  169 - 0xa9
    "10101001", --   22 - 0x16  :  169 - 0xa9
    "10101001", --   23 - 0x17  :  169 - 0xa9
    "10101001", --   24 - 0x18  :  169 - 0xa9
    "10101001", --   25 - 0x19  :  169 - 0xa9
    "10101001", --   26 - 0x1a  :  169 - 0xa9
    "10101001", --   27 - 0x1b  :  169 - 0xa9
    "10101001", --   28 - 0x1c  :  169 - 0xa9
    "10101001", --   29 - 0x1d  :  169 - 0xa9
    "10101001", --   30 - 0x1e  :  169 - 0xa9
    "10101001", --   31 - 0x1f  :  169 - 0xa9
    "10101001", --   32 - 0x20  :  169 - 0xa9 -- line 0x1
    "10101001", --   33 - 0x21  :  169 - 0xa9
    "10101001", --   34 - 0x22  :  169 - 0xa9
    "10101001", --   35 - 0x23  :  169 - 0xa9
    "10101001", --   36 - 0x24  :  169 - 0xa9
    "10101001", --   37 - 0x25  :  169 - 0xa9
    "10101001", --   38 - 0x26  :  169 - 0xa9
    "10101001", --   39 - 0x27  :  169 - 0xa9
    "10101001", --   40 - 0x28  :  169 - 0xa9
    "10101001", --   41 - 0x29  :  169 - 0xa9
    "10101001", --   42 - 0x2a  :  169 - 0xa9
    "10101001", --   43 - 0x2b  :  169 - 0xa9
    "10101001", --   44 - 0x2c  :  169 - 0xa9
    "10101001", --   45 - 0x2d  :  169 - 0xa9
    "10101001", --   46 - 0x2e  :  169 - 0xa9
    "10101001", --   47 - 0x2f  :  169 - 0xa9
    "10101001", --   48 - 0x30  :  169 - 0xa9
    "10101001", --   49 - 0x31  :  169 - 0xa9
    "10101001", --   50 - 0x32  :  169 - 0xa9
    "10101001", --   51 - 0x33  :  169 - 0xa9
    "10101001", --   52 - 0x34  :  169 - 0xa9
    "10101001", --   53 - 0x35  :  169 - 0xa9
    "10101001", --   54 - 0x36  :  169 - 0xa9
    "10101001", --   55 - 0x37  :  169 - 0xa9
    "10101001", --   56 - 0x38  :  169 - 0xa9
    "10101001", --   57 - 0x39  :  169 - 0xa9
    "10101001", --   58 - 0x3a  :  169 - 0xa9
    "10101001", --   59 - 0x3b  :  169 - 0xa9
    "10101001", --   60 - 0x3c  :  169 - 0xa9
    "10101001", --   61 - 0x3d  :  169 - 0xa9
    "10101001", --   62 - 0x3e  :  169 - 0xa9
    "10101001", --   63 - 0x3f  :  169 - 0xa9
    "10101001", --   64 - 0x40  :  169 - 0xa9 -- line 0x2
    "10101001", --   65 - 0x41  :  169 - 0xa9
    "01010110", --   66 - 0x42  :   86 - 0x56
    "01010101", --   67 - 0x43  :   85 - 0x55
    "01010111", --   68 - 0x44  :   87 - 0x57
    "01011000", --   69 - 0x45  :   88 - 0x58
    "11010000", --   70 - 0x46  :  208 - 0xd0
    "11010001", --   71 - 0x47  :  209 - 0xd1
    "10101001", --   72 - 0x48  :  169 - 0xa9
    "01011101", --   73 - 0x49  :   93 - 0x5d
    "01011110", --   74 - 0x4a  :   94 - 0x5e
    "01011011", --   75 - 0x4b  :   91 - 0x5b
    "01010110", --   76 - 0x4c  :   86 - 0x56
    "11111001", --   77 - 0x4d  :  249 - 0xf9
    "11111010", --   78 - 0x4e  :  250 - 0xfa
    "11111010", --   79 - 0x4f  :  250 - 0xfa
    "11111010", --   80 - 0x50  :  250 - 0xfa
    "11111010", --   81 - 0x51  :  250 - 0xfa
    "11111010", --   82 - 0x52  :  250 - 0xfa
    "11111010", --   83 - 0x53  :  250 - 0xfa
    "11111011", --   84 - 0x54  :  251 - 0xfb
    "10101001", --   85 - 0x55  :  169 - 0xa9
    "01011001", --   86 - 0x56  :   89 - 0x59
    "01011010", --   87 - 0x57  :   90 - 0x5a
    "01011000", --   88 - 0x58  :   88 - 0x58
    "01011011", --   89 - 0x59  :   91 - 0x5b
    "11010000", --   90 - 0x5a  :  208 - 0xd0
    "11010000", --   91 - 0x5b  :  208 - 0xd0
    "11010000", --   92 - 0x5c  :  208 - 0xd0
    "01011100", --   93 - 0x5d  :   92 - 0x5c
    "10101001", --   94 - 0x5e  :  169 - 0xa9
    "10101001", --   95 - 0x5f  :  169 - 0xa9
    "10101001", --   96 - 0x60  :  169 - 0xa9 -- line 0x3
    "10101001", --   97 - 0x61  :  169 - 0xa9
    "01100110", --   98 - 0x62  :  102 - 0x66
    "01100101", --   99 - 0x63  :  101 - 0x65
    "01100111", --  100 - 0x64  :  103 - 0x67
    "01101000", --  101 - 0x65  :  104 - 0x68
    "11100000", --  102 - 0x66  :  224 - 0xe0
    "11100001", --  103 - 0x67  :  225 - 0xe1
    "10101001", --  104 - 0x68  :  169 - 0xa9
    "01101101", --  105 - 0x69  :  109 - 0x6d
    "01101110", --  106 - 0x6a  :  110 - 0x6e
    "01101011", --  107 - 0x6b  :  107 - 0x6b
    "01100110", --  108 - 0x6c  :  102 - 0x66
    "11111100", --  109 - 0x6d  :  252 - 0xfc
    "11111101", --  110 - 0x6e  :  253 - 0xfd
    "11111101", --  111 - 0x6f  :  253 - 0xfd
    "11111101", --  112 - 0x70  :  253 - 0xfd
    "11111101", --  113 - 0x71  :  253 - 0xfd
    "11111101", --  114 - 0x72  :  253 - 0xfd
    "11111101", --  115 - 0x73  :  253 - 0xfd
    "11111110", --  116 - 0x74  :  254 - 0xfe
    "10101001", --  117 - 0x75  :  169 - 0xa9
    "01101001", --  118 - 0x76  :  105 - 0x69
    "01101010", --  119 - 0x77  :  106 - 0x6a
    "01101000", --  120 - 0x78  :  104 - 0x68
    "01101011", --  121 - 0x79  :  107 - 0x6b
    "11100000", --  122 - 0x7a  :  224 - 0xe0
    "11100000", --  123 - 0x7b  :  224 - 0xe0
    "11100000", --  124 - 0x7c  :  224 - 0xe0
    "01101100", --  125 - 0x7d  :  108 - 0x6c
    "10101001", --  126 - 0x7e  :  169 - 0xa9
    "10101001", --  127 - 0x7f  :  169 - 0xa9
    "10101010", --  128 - 0x80  :  170 - 0xaa -- line 0x4
    "10101010", --  129 - 0x81  :  170 - 0xaa
    "10101010", --  130 - 0x82  :  170 - 0xaa
    "10101010", --  131 - 0x83  :  170 - 0xaa
    "10101010", --  132 - 0x84  :  170 - 0xaa
    "10101010", --  133 - 0x85  :  170 - 0xaa
    "10101010", --  134 - 0x86  :  170 - 0xaa
    "10101010", --  135 - 0x87  :  170 - 0xaa
    "10101010", --  136 - 0x88  :  170 - 0xaa
    "10101010", --  137 - 0x89  :  170 - 0xaa
    "10101010", --  138 - 0x8a  :  170 - 0xaa
    "10101010", --  139 - 0x8b  :  170 - 0xaa
    "10101010", --  140 - 0x8c  :  170 - 0xaa
    "10101010", --  141 - 0x8d  :  170 - 0xaa
    "10101010", --  142 - 0x8e  :  170 - 0xaa
    "10101010", --  143 - 0x8f  :  170 - 0xaa
    "10101010", --  144 - 0x90  :  170 - 0xaa
    "10101010", --  145 - 0x91  :  170 - 0xaa
    "10101010", --  146 - 0x92  :  170 - 0xaa
    "10101010", --  147 - 0x93  :  170 - 0xaa
    "10101010", --  148 - 0x94  :  170 - 0xaa
    "10101010", --  149 - 0x95  :  170 - 0xaa
    "10101010", --  150 - 0x96  :  170 - 0xaa
    "10101010", --  151 - 0x97  :  170 - 0xaa
    "10101010", --  152 - 0x98  :  170 - 0xaa
    "10101010", --  153 - 0x99  :  170 - 0xaa
    "10101010", --  154 - 0x9a  :  170 - 0xaa
    "10101010", --  155 - 0x9b  :  170 - 0xaa
    "10101010", --  156 - 0x9c  :  170 - 0xaa
    "10101010", --  157 - 0x9d  :  170 - 0xaa
    "10101010", --  158 - 0x9e  :  170 - 0xaa
    "10101010", --  159 - 0x9f  :  170 - 0xaa
    "10100000", --  160 - 0xa0  :  160 - 0xa0 -- line 0x5
    "10100001", --  161 - 0xa1  :  161 - 0xa1
    "10100010", --  162 - 0xa2  :  162 - 0xa2
    "10100010", --  163 - 0xa3  :  162 - 0xa2
    "10100010", --  164 - 0xa4  :  162 - 0xa2
    "10100010", --  165 - 0xa5  :  162 - 0xa2
    "10100010", --  166 - 0xa6  :  162 - 0xa2
    "10100010", --  167 - 0xa7  :  162 - 0xa2
    "10100010", --  168 - 0xa8  :  162 - 0xa2
    "10100010", --  169 - 0xa9  :  162 - 0xa2
    "10100010", --  170 - 0xaa  :  162 - 0xa2
    "10100010", --  171 - 0xab  :  162 - 0xa2
    "10100010", --  172 - 0xac  :  162 - 0xa2
    "10100010", --  173 - 0xad  :  162 - 0xa2
    "10100010", --  174 - 0xae  :  162 - 0xa2
    "10100010", --  175 - 0xaf  :  162 - 0xa2
    "10100010", --  176 - 0xb0  :  162 - 0xa2
    "10100010", --  177 - 0xb1  :  162 - 0xa2
    "10100010", --  178 - 0xb2  :  162 - 0xa2
    "10100010", --  179 - 0xb3  :  162 - 0xa2
    "10100010", --  180 - 0xb4  :  162 - 0xa2
    "10100010", --  181 - 0xb5  :  162 - 0xa2
    "10100010", --  182 - 0xb6  :  162 - 0xa2
    "10100010", --  183 - 0xb7  :  162 - 0xa2
    "10100010", --  184 - 0xb8  :  162 - 0xa2
    "10100010", --  185 - 0xb9  :  162 - 0xa2
    "10100010", --  186 - 0xba  :  162 - 0xa2
    "10100010", --  187 - 0xbb  :  162 - 0xa2
    "10100010", --  188 - 0xbc  :  162 - 0xa2
    "10100010", --  189 - 0xbd  :  162 - 0xa2
    "10100110", --  190 - 0xbe  :  166 - 0xa6
    "10100000", --  191 - 0xbf  :  160 - 0xa0
    "10100000", --  192 - 0xc0  :  160 - 0xa0 -- line 0x6
    "10100011", --  193 - 0xc1  :  163 - 0xa3
    "10000000", --  194 - 0xc2  :  128 - 0x80
    "10000001", --  195 - 0xc3  :  129 - 0x81
    "10000000", --  196 - 0xc4  :  128 - 0x80
    "10000001", --  197 - 0xc5  :  129 - 0x81
    "10000000", --  198 - 0xc6  :  128 - 0x80
    "10000010", --  199 - 0xc7  :  130 - 0x82
    "10000000", --  200 - 0xc8  :  128 - 0x80
    "10000001", --  201 - 0xc9  :  129 - 0x81
    "10000001", --  202 - 0xca  :  129 - 0x81
    "10000000", --  203 - 0xcb  :  128 - 0x80
    "10000000", --  204 - 0xcc  :  128 - 0x80
    "10000001", --  205 - 0xcd  :  129 - 0x81
    "10000010", --  206 - 0xce  :  130 - 0x82
    "10000011", --  207 - 0xcf  :  131 - 0x83
    "10000010", --  208 - 0xd0  :  130 - 0x82
    "10000011", --  209 - 0xd1  :  131 - 0x83
    "10000000", --  210 - 0xd2  :  128 - 0x80
    "10000010", --  211 - 0xd3  :  130 - 0x82
    "10000000", --  212 - 0xd4  :  128 - 0x80
    "10000010", --  213 - 0xd5  :  130 - 0x82
    "10000010", --  214 - 0xd6  :  130 - 0x82
    "10000011", --  215 - 0xd7  :  131 - 0x83
    "10000010", --  216 - 0xd8  :  130 - 0x82
    "10000011", --  217 - 0xd9  :  131 - 0x83
    "10000001", --  218 - 0xda  :  129 - 0x81
    "10000000", --  219 - 0xdb  :  128 - 0x80
    "10000000", --  220 - 0xdc  :  128 - 0x80
    "10000001", --  221 - 0xdd  :  129 - 0x81
    "10100111", --  222 - 0xde  :  167 - 0xa7
    "10100000", --  223 - 0xdf  :  160 - 0xa0
    "10100000", --  224 - 0xe0  :  160 - 0xa0 -- line 0x7
    "10100011", --  225 - 0xe1  :  163 - 0xa3
    "10010000", --  226 - 0xe2  :  144 - 0x90
    "10010001", --  227 - 0xe3  :  145 - 0x91
    "10010000", --  228 - 0xe4  :  144 - 0x90
    "10010001", --  229 - 0xe5  :  145 - 0x91
    "10010010", --  230 - 0xe6  :  146 - 0x92
    "10010001", --  231 - 0xe7  :  145 - 0x91
    "10010000", --  232 - 0xe8  :  144 - 0x90
    "10010001", --  233 - 0xe9  :  145 - 0x91
    "10010011", --  234 - 0xea  :  147 - 0x93
    "10010010", --  235 - 0xeb  :  146 - 0x92
    "10010000", --  236 - 0xec  :  144 - 0x90
    "10010001", --  237 - 0xed  :  145 - 0x91
    "10010010", --  238 - 0xee  :  146 - 0x92
    "10010011", --  239 - 0xef  :  147 - 0x93
    "10010010", --  240 - 0xf0  :  146 - 0x92
    "10010011", --  241 - 0xf1  :  147 - 0x93
    "10010010", --  242 - 0xf2  :  146 - 0x92
    "10010001", --  243 - 0xf3  :  145 - 0x91
    "10010010", --  244 - 0xf4  :  146 - 0x92
    "10010001", --  245 - 0xf5  :  145 - 0x91
    "10010010", --  246 - 0xf6  :  146 - 0x92
    "10010011", --  247 - 0xf7  :  147 - 0x93
    "10010010", --  248 - 0xf8  :  146 - 0x92
    "10010011", --  249 - 0xf9  :  147 - 0x93
    "10010011", --  250 - 0xfa  :  147 - 0x93
    "10010010", --  251 - 0xfb  :  146 - 0x92
    "10010000", --  252 - 0xfc  :  144 - 0x90
    "10010001", --  253 - 0xfd  :  145 - 0x91
    "10100111", --  254 - 0xfe  :  167 - 0xa7
    "10100000", --  255 - 0xff  :  160 - 0xa0
    "10100000", --  256 - 0x100  :  160 - 0xa0 -- line 0x8
    "10100011", --  257 - 0x101  :  163 - 0xa3
    "10000010", --  258 - 0x102  :  130 - 0x82
    "10000011", --  259 - 0x103  :  131 - 0x83
    "10000101", --  260 - 0x104  :  133 - 0x85
    "10000110", --  261 - 0x105  :  134 - 0x86
    "10000101", --  262 - 0x106  :  133 - 0x85
    "10000110", --  263 - 0x107  :  134 - 0x86
    "10000101", --  264 - 0x108  :  133 - 0x85
    "10000110", --  265 - 0x109  :  134 - 0x86
    "10000101", --  266 - 0x10a  :  133 - 0x85
    "10000110", --  267 - 0x10b  :  134 - 0x86
    "10000100", --  268 - 0x10c  :  132 - 0x84
    "10000111", --  269 - 0x10d  :  135 - 0x87
    "10000110", --  270 - 0x10e  :  134 - 0x86
    "10000111", --  271 - 0x10f  :  135 - 0x87
    "10000100", --  272 - 0x110  :  132 - 0x84
    "10000101", --  273 - 0x111  :  133 - 0x85
    "10000101", --  274 - 0x112  :  133 - 0x85
    "10000110", --  275 - 0x113  :  134 - 0x86
    "10000101", --  276 - 0x114  :  133 - 0x85
    "10000110", --  277 - 0x115  :  134 - 0x86
    "10000110", --  278 - 0x116  :  134 - 0x86
    "10000111", --  279 - 0x117  :  135 - 0x87
    "10000110", --  280 - 0x118  :  134 - 0x86
    "10000111", --  281 - 0x119  :  135 - 0x87
    "10000100", --  282 - 0x11a  :  132 - 0x84
    "10000101", --  283 - 0x11b  :  133 - 0x85
    "10000010", --  284 - 0x11c  :  130 - 0x82
    "10000011", --  285 - 0x11d  :  131 - 0x83
    "10100111", --  286 - 0x11e  :  167 - 0xa7
    "10100000", --  287 - 0x11f  :  160 - 0xa0
    "10100000", --  288 - 0x120  :  160 - 0xa0 -- line 0x9
    "10100011", --  289 - 0x121  :  163 - 0xa3
    "10010010", --  290 - 0x122  :  146 - 0x92
    "10010011", --  291 - 0x123  :  147 - 0x93
    "10010111", --  292 - 0x124  :  151 - 0x97
    "10010100", --  293 - 0x125  :  148 - 0x94
    "10010111", --  294 - 0x126  :  151 - 0x97
    "10010100", --  295 - 0x127  :  148 - 0x94
    "10010111", --  296 - 0x128  :  151 - 0x97
    "10010100", --  297 - 0x129  :  148 - 0x94
    "10010111", --  298 - 0x12a  :  151 - 0x97
    "10010100", --  299 - 0x12b  :  148 - 0x94
    "10010110", --  300 - 0x12c  :  150 - 0x96
    "10010101", --  301 - 0x12d  :  149 - 0x95
    "10010110", --  302 - 0x12e  :  150 - 0x96
    "10010111", --  303 - 0x12f  :  151 - 0x97
    "10010100", --  304 - 0x130  :  148 - 0x94
    "10010101", --  305 - 0x131  :  149 - 0x95
    "10010111", --  306 - 0x132  :  151 - 0x97
    "10010100", --  307 - 0x133  :  148 - 0x94
    "10010111", --  308 - 0x134  :  151 - 0x97
    "10010100", --  309 - 0x135  :  148 - 0x94
    "10010110", --  310 - 0x136  :  150 - 0x96
    "10010111", --  311 - 0x137  :  151 - 0x97
    "10010110", --  312 - 0x138  :  150 - 0x96
    "10010111", --  313 - 0x139  :  151 - 0x97
    "10010100", --  314 - 0x13a  :  148 - 0x94
    "10010101", --  315 - 0x13b  :  149 - 0x95
    "10010010", --  316 - 0x13c  :  146 - 0x92
    "10010011", --  317 - 0x13d  :  147 - 0x93
    "10100111", --  318 - 0x13e  :  167 - 0xa7
    "10100000", --  319 - 0x13f  :  160 - 0xa0
    "10100000", --  320 - 0x140  :  160 - 0xa0 -- line 0xa
    "10100011", --  321 - 0x141  :  163 - 0xa3
    "10000000", --  322 - 0x142  :  128 - 0x80
    "10000010", --  323 - 0x143  :  130 - 0x82
    "10000100", --  324 - 0x144  :  132 - 0x84
    "10000111", --  325 - 0x145  :  135 - 0x87
    "10000101", --  326 - 0x146  :  133 - 0x85
    "10000110", --  327 - 0x147  :  134 - 0x86
    "10000100", --  328 - 0x148  :  132 - 0x84
    "10000111", --  329 - 0x149  :  135 - 0x87
    "10000100", --  330 - 0x14a  :  132 - 0x84
    "10000111", --  331 - 0x14b  :  135 - 0x87
    "10000110", --  332 - 0x14c  :  134 - 0x86
    "10000111", --  333 - 0x14d  :  135 - 0x87
    "10000100", --  334 - 0x14e  :  132 - 0x84
    "10000101", --  335 - 0x14f  :  133 - 0x85
    "10000100", --  336 - 0x150  :  132 - 0x84
    "10000101", --  337 - 0x151  :  133 - 0x85
    "10000110", --  338 - 0x152  :  134 - 0x86
    "10000111", --  339 - 0x153  :  135 - 0x87
    "10000100", --  340 - 0x154  :  132 - 0x84
    "10000101", --  341 - 0x155  :  133 - 0x85
    "10000101", --  342 - 0x156  :  133 - 0x85
    "10000110", --  343 - 0x157  :  134 - 0x86
    "10000100", --  344 - 0x158  :  132 - 0x84
    "10000111", --  345 - 0x159  :  135 - 0x87
    "10000100", --  346 - 0x15a  :  132 - 0x84
    "10000111", --  347 - 0x15b  :  135 - 0x87
    "10000000", --  348 - 0x15c  :  128 - 0x80
    "10000001", --  349 - 0x15d  :  129 - 0x81
    "10100111", --  350 - 0x15e  :  167 - 0xa7
    "10100000", --  351 - 0x15f  :  160 - 0xa0
    "10100000", --  352 - 0x160  :  160 - 0xa0 -- line 0xb
    "10100011", --  353 - 0x161  :  163 - 0xa3
    "10010010", --  354 - 0x162  :  146 - 0x92
    "10010001", --  355 - 0x163  :  145 - 0x91
    "10010110", --  356 - 0x164  :  150 - 0x96
    "10010101", --  357 - 0x165  :  149 - 0x95
    "10010111", --  358 - 0x166  :  151 - 0x97
    "10010100", --  359 - 0x167  :  148 - 0x94
    "10010110", --  360 - 0x168  :  150 - 0x96
    "10010101", --  361 - 0x169  :  149 - 0x95
    "10010110", --  362 - 0x16a  :  150 - 0x96
    "10010101", --  363 - 0x16b  :  149 - 0x95
    "10010110", --  364 - 0x16c  :  150 - 0x96
    "10010111", --  365 - 0x16d  :  151 - 0x97
    "10010100", --  366 - 0x16e  :  148 - 0x94
    "10010101", --  367 - 0x16f  :  149 - 0x95
    "10010100", --  368 - 0x170  :  148 - 0x94
    "10010101", --  369 - 0x171  :  149 - 0x95
    "10010110", --  370 - 0x172  :  150 - 0x96
    "10010111", --  371 - 0x173  :  151 - 0x97
    "10010100", --  372 - 0x174  :  148 - 0x94
    "10010101", --  373 - 0x175  :  149 - 0x95
    "10010111", --  374 - 0x176  :  151 - 0x97
    "10010100", --  375 - 0x177  :  148 - 0x94
    "10010110", --  376 - 0x178  :  150 - 0x96
    "10010101", --  377 - 0x179  :  149 - 0x95
    "10010110", --  378 - 0x17a  :  150 - 0x96
    "10010101", --  379 - 0x17b  :  149 - 0x95
    "10010000", --  380 - 0x17c  :  144 - 0x90
    "10010001", --  381 - 0x17d  :  145 - 0x91
    "10100111", --  382 - 0x17e  :  167 - 0xa7
    "10100000", --  383 - 0x17f  :  160 - 0xa0
    "10100000", --  384 - 0x180  :  160 - 0xa0 -- line 0xc
    "10100011", --  385 - 0x181  :  163 - 0xa3
    "10000010", --  386 - 0x182  :  130 - 0x82
    "10000011", --  387 - 0x183  :  131 - 0x83
    "10000110", --  388 - 0x184  :  134 - 0x86
    "10000111", --  389 - 0x185  :  135 - 0x87
    "10000100", --  390 - 0x186  :  132 - 0x84
    "10000101", --  391 - 0x187  :  133 - 0x85
    "10000100", --  392 - 0x188  :  132 - 0x84
    "10000111", --  393 - 0x189  :  135 - 0x87
    "10000100", --  394 - 0x18a  :  132 - 0x84
    "10000111", --  395 - 0x18b  :  135 - 0x87
    "10000110", --  396 - 0x18c  :  134 - 0x86
    "10000111", --  397 - 0x18d  :  135 - 0x87
    "10000100", --  398 - 0x18e  :  132 - 0x84
    "10000111", --  399 - 0x18f  :  135 - 0x87
    "10000110", --  400 - 0x190  :  134 - 0x86
    "10000111", --  401 - 0x191  :  135 - 0x87
    "10000110", --  402 - 0x192  :  134 - 0x86
    "10000111", --  403 - 0x193  :  135 - 0x87
    "10000110", --  404 - 0x194  :  134 - 0x86
    "10000111", --  405 - 0x195  :  135 - 0x87
    "10000110", --  406 - 0x196  :  134 - 0x86
    "10000111", --  407 - 0x197  :  135 - 0x87
    "10000101", --  408 - 0x198  :  133 - 0x85
    "10000110", --  409 - 0x199  :  134 - 0x86
    "10000100", --  410 - 0x19a  :  132 - 0x84
    "10000111", --  411 - 0x19b  :  135 - 0x87
    "10000000", --  412 - 0x19c  :  128 - 0x80
    "10000010", --  413 - 0x19d  :  130 - 0x82
    "10100111", --  414 - 0x19e  :  167 - 0xa7
    "10100000", --  415 - 0x19f  :  160 - 0xa0
    "10100000", --  416 - 0x1a0  :  160 - 0xa0 -- line 0xd
    "10100011", --  417 - 0x1a1  :  163 - 0xa3
    "10010010", --  418 - 0x1a2  :  146 - 0x92
    "10010011", --  419 - 0x1a3  :  147 - 0x93
    "10010110", --  420 - 0x1a4  :  150 - 0x96
    "10010111", --  421 - 0x1a5  :  151 - 0x97
    "10010100", --  422 - 0x1a6  :  148 - 0x94
    "10010101", --  423 - 0x1a7  :  149 - 0x95
    "10010110", --  424 - 0x1a8  :  150 - 0x96
    "10010101", --  425 - 0x1a9  :  149 - 0x95
    "10010110", --  426 - 0x1aa  :  150 - 0x96
    "10010101", --  427 - 0x1ab  :  149 - 0x95
    "10010110", --  428 - 0x1ac  :  150 - 0x96
    "10010111", --  429 - 0x1ad  :  151 - 0x97
    "10010110", --  430 - 0x1ae  :  150 - 0x96
    "10010101", --  431 - 0x1af  :  149 - 0x95
    "10010110", --  432 - 0x1b0  :  150 - 0x96
    "10010111", --  433 - 0x1b1  :  151 - 0x97
    "10010110", --  434 - 0x1b2  :  150 - 0x96
    "10010111", --  435 - 0x1b3  :  151 - 0x97
    "10010110", --  436 - 0x1b4  :  150 - 0x96
    "10010111", --  437 - 0x1b5  :  151 - 0x97
    "10010110", --  438 - 0x1b6  :  150 - 0x96
    "10010111", --  439 - 0x1b7  :  151 - 0x97
    "10010111", --  440 - 0x1b8  :  151 - 0x97
    "10010100", --  441 - 0x1b9  :  148 - 0x94
    "10010110", --  442 - 0x1ba  :  150 - 0x96
    "10010101", --  443 - 0x1bb  :  149 - 0x95
    "10010010", --  444 - 0x1bc  :  146 - 0x92
    "10010001", --  445 - 0x1bd  :  145 - 0x91
    "10100111", --  446 - 0x1be  :  167 - 0xa7
    "10100000", --  447 - 0x1bf  :  160 - 0xa0
    "10100000", --  448 - 0x1c0  :  160 - 0xa0 -- line 0xe
    "10100011", --  449 - 0x1c1  :  163 - 0xa3
    "10000000", --  450 - 0x1c2  :  128 - 0x80
    "10000001", --  451 - 0x1c3  :  129 - 0x81
    "10000101", --  452 - 0x1c4  :  133 - 0x85
    "10000110", --  453 - 0x1c5  :  134 - 0x86
    "10000100", --  454 - 0x1c6  :  132 - 0x84
    "10000101", --  455 - 0x1c7  :  133 - 0x85
    "10000100", --  456 - 0x1c8  :  132 - 0x84
    "10000101", --  457 - 0x1c9  :  133 - 0x85
    "10000100", --  458 - 0x1ca  :  132 - 0x84
    "10000111", --  459 - 0x1cb  :  135 - 0x87
    "10000001", --  460 - 0x1cc  :  129 - 0x81
    "10000000", --  461 - 0x1cd  :  128 - 0x80
    "10000010", --  462 - 0x1ce  :  130 - 0x82
    "10000011", --  463 - 0x1cf  :  131 - 0x83
    "10000010", --  464 - 0x1d0  :  130 - 0x82
    "10000011", --  465 - 0x1d1  :  131 - 0x83
    "10000001", --  466 - 0x1d2  :  129 - 0x81
    "10000000", --  467 - 0x1d3  :  128 - 0x80
    "10000101", --  468 - 0x1d4  :  133 - 0x85
    "10000110", --  469 - 0x1d5  :  134 - 0x86
    "10000110", --  470 - 0x1d6  :  134 - 0x86
    "10000111", --  471 - 0x1d7  :  135 - 0x87
    "10000100", --  472 - 0x1d8  :  132 - 0x84
    "10000111", --  473 - 0x1d9  :  135 - 0x87
    "10000100", --  474 - 0x1da  :  132 - 0x84
    "10000111", --  475 - 0x1db  :  135 - 0x87
    "10000000", --  476 - 0x1dc  :  128 - 0x80
    "10000001", --  477 - 0x1dd  :  129 - 0x81
    "10100111", --  478 - 0x1de  :  167 - 0xa7
    "10100000", --  479 - 0x1df  :  160 - 0xa0
    "10100000", --  480 - 0x1e0  :  160 - 0xa0 -- line 0xf
    "10100011", --  481 - 0x1e1  :  163 - 0xa3
    "10010000", --  482 - 0x1e2  :  144 - 0x90
    "10010001", --  483 - 0x1e3  :  145 - 0x91
    "10010111", --  484 - 0x1e4  :  151 - 0x97
    "10010100", --  485 - 0x1e5  :  148 - 0x94
    "10010100", --  486 - 0x1e6  :  148 - 0x94
    "10010101", --  487 - 0x1e7  :  149 - 0x95
    "10010100", --  488 - 0x1e8  :  148 - 0x94
    "10010101", --  489 - 0x1e9  :  149 - 0x95
    "10010110", --  490 - 0x1ea  :  150 - 0x96
    "10010101", --  491 - 0x1eb  :  149 - 0x95
    "10010011", --  492 - 0x1ec  :  147 - 0x93
    "10010010", --  493 - 0x1ed  :  146 - 0x92
    "10010010", --  494 - 0x1ee  :  146 - 0x92
    "10010011", --  495 - 0x1ef  :  147 - 0x93
    "10010010", --  496 - 0x1f0  :  146 - 0x92
    "10010011", --  497 - 0x1f1  :  147 - 0x93
    "10010011", --  498 - 0x1f2  :  147 - 0x93
    "10010010", --  499 - 0x1f3  :  146 - 0x92
    "10010111", --  500 - 0x1f4  :  151 - 0x97
    "10010100", --  501 - 0x1f5  :  148 - 0x94
    "10010110", --  502 - 0x1f6  :  150 - 0x96
    "10010111", --  503 - 0x1f7  :  151 - 0x97
    "10010110", --  504 - 0x1f8  :  150 - 0x96
    "10010101", --  505 - 0x1f9  :  149 - 0x95
    "10010110", --  506 - 0x1fa  :  150 - 0x96
    "10010101", --  507 - 0x1fb  :  149 - 0x95
    "10010000", --  508 - 0x1fc  :  144 - 0x90
    "10010001", --  509 - 0x1fd  :  145 - 0x91
    "10100111", --  510 - 0x1fe  :  167 - 0xa7
    "10100000", --  511 - 0x1ff  :  160 - 0xa0
    "10100000", --  512 - 0x200  :  160 - 0xa0 -- line 0x10
    "10100011", --  513 - 0x201  :  163 - 0xa3
    "10000010", --  514 - 0x202  :  130 - 0x82
    "10000011", --  515 - 0x203  :  131 - 0x83
    "10000101", --  516 - 0x204  :  133 - 0x85
    "10000110", --  517 - 0x205  :  134 - 0x86
    "10000101", --  518 - 0x206  :  133 - 0x85
    "10000110", --  519 - 0x207  :  134 - 0x86
    "10000101", --  520 - 0x208  :  133 - 0x85
    "10000110", --  521 - 0x209  :  134 - 0x86
    "10000101", --  522 - 0x20a  :  133 - 0x85
    "10000110", --  523 - 0x20b  :  134 - 0x86
    "10000000", --  524 - 0x20c  :  128 - 0x80
    "10000010", --  525 - 0x20d  :  130 - 0x82
    "10000010", --  526 - 0x20e  :  130 - 0x82
    "10000011", --  527 - 0x20f  :  131 - 0x83
    "10000000", --  528 - 0x210  :  128 - 0x80
    "10000001", --  529 - 0x211  :  129 - 0x81
    "10000001", --  530 - 0x212  :  129 - 0x81
    "10000000", --  531 - 0x213  :  128 - 0x80
    "10000101", --  532 - 0x214  :  133 - 0x85
    "10000110", --  533 - 0x215  :  134 - 0x86
    "10000110", --  534 - 0x216  :  134 - 0x86
    "10000111", --  535 - 0x217  :  135 - 0x87
    "10000110", --  536 - 0x218  :  134 - 0x86
    "10000111", --  537 - 0x219  :  135 - 0x87
    "10000100", --  538 - 0x21a  :  132 - 0x84
    "10000101", --  539 - 0x21b  :  133 - 0x85
    "10000010", --  540 - 0x21c  :  130 - 0x82
    "10000011", --  541 - 0x21d  :  131 - 0x83
    "10100111", --  542 - 0x21e  :  167 - 0xa7
    "10100000", --  543 - 0x21f  :  160 - 0xa0
    "10100000", --  544 - 0x220  :  160 - 0xa0 -- line 0x11
    "10100011", --  545 - 0x221  :  163 - 0xa3
    "10010010", --  546 - 0x222  :  146 - 0x92
    "10010011", --  547 - 0x223  :  147 - 0x93
    "10010111", --  548 - 0x224  :  151 - 0x97
    "10010100", --  549 - 0x225  :  148 - 0x94
    "10010111", --  550 - 0x226  :  151 - 0x97
    "10010100", --  551 - 0x227  :  148 - 0x94
    "10010111", --  552 - 0x228  :  151 - 0x97
    "10010100", --  553 - 0x229  :  148 - 0x94
    "10010111", --  554 - 0x22a  :  151 - 0x97
    "10010100", --  555 - 0x22b  :  148 - 0x94
    "10010010", --  556 - 0x22c  :  146 - 0x92
    "10010001", --  557 - 0x22d  :  145 - 0x91
    "10010010", --  558 - 0x22e  :  146 - 0x92
    "10010011", --  559 - 0x22f  :  147 - 0x93
    "10010000", --  560 - 0x230  :  144 - 0x90
    "10010001", --  561 - 0x231  :  145 - 0x91
    "10010011", --  562 - 0x232  :  147 - 0x93
    "10010010", --  563 - 0x233  :  146 - 0x92
    "10010111", --  564 - 0x234  :  151 - 0x97
    "10010100", --  565 - 0x235  :  148 - 0x94
    "10010110", --  566 - 0x236  :  150 - 0x96
    "10010111", --  567 - 0x237  :  151 - 0x97
    "10010110", --  568 - 0x238  :  150 - 0x96
    "10010111", --  569 - 0x239  :  151 - 0x97
    "10010100", --  570 - 0x23a  :  148 - 0x94
    "10010101", --  571 - 0x23b  :  149 - 0x95
    "10010010", --  572 - 0x23c  :  146 - 0x92
    "10010011", --  573 - 0x23d  :  147 - 0x93
    "10100111", --  574 - 0x23e  :  167 - 0xa7
    "10100000", --  575 - 0x23f  :  160 - 0xa0
    "10100000", --  576 - 0x240  :  160 - 0xa0 -- line 0x12
    "10100011", --  577 - 0x241  :  163 - 0xa3
    "10000000", --  578 - 0x242  :  128 - 0x80
    "10000010", --  579 - 0x243  :  130 - 0x82
    "10000100", --  580 - 0x244  :  132 - 0x84
    "10000111", --  581 - 0x245  :  135 - 0x87
    "10000101", --  582 - 0x246  :  133 - 0x85
    "10000110", --  583 - 0x247  :  134 - 0x86
    "10000100", --  584 - 0x248  :  132 - 0x84
    "10000111", --  585 - 0x249  :  135 - 0x87
    "10000100", --  586 - 0x24a  :  132 - 0x84
    "10000111", --  587 - 0x24b  :  135 - 0x87
    "10000010", --  588 - 0x24c  :  130 - 0x82
    "10000011", --  589 - 0x24d  :  131 - 0x83
    "10000000", --  590 - 0x24e  :  128 - 0x80
    "10000001", --  591 - 0x24f  :  129 - 0x81
    "10000000", --  592 - 0x250  :  128 - 0x80
    "10000001", --  593 - 0x251  :  129 - 0x81
    "10000010", --  594 - 0x252  :  130 - 0x82
    "10000011", --  595 - 0x253  :  131 - 0x83
    "10000100", --  596 - 0x254  :  132 - 0x84
    "10000101", --  597 - 0x255  :  133 - 0x85
    "10000101", --  598 - 0x256  :  133 - 0x85
    "10000110", --  599 - 0x257  :  134 - 0x86
    "10000100", --  600 - 0x258  :  132 - 0x84
    "10000111", --  601 - 0x259  :  135 - 0x87
    "10000100", --  602 - 0x25a  :  132 - 0x84
    "10000111", --  603 - 0x25b  :  135 - 0x87
    "10000000", --  604 - 0x25c  :  128 - 0x80
    "10000001", --  605 - 0x25d  :  129 - 0x81
    "10100111", --  606 - 0x25e  :  167 - 0xa7
    "10100000", --  607 - 0x25f  :  160 - 0xa0
    "10100000", --  608 - 0x260  :  160 - 0xa0 -- line 0x13
    "10100011", --  609 - 0x261  :  163 - 0xa3
    "10010010", --  610 - 0x262  :  146 - 0x92
    "10010001", --  611 - 0x263  :  145 - 0x91
    "10010110", --  612 - 0x264  :  150 - 0x96
    "10010101", --  613 - 0x265  :  149 - 0x95
    "10010111", --  614 - 0x266  :  151 - 0x97
    "10010100", --  615 - 0x267  :  148 - 0x94
    "10010110", --  616 - 0x268  :  150 - 0x96
    "10010101", --  617 - 0x269  :  149 - 0x95
    "10010110", --  618 - 0x26a  :  150 - 0x96
    "10010101", --  619 - 0x26b  :  149 - 0x95
    "10010010", --  620 - 0x26c  :  146 - 0x92
    "10010011", --  621 - 0x26d  :  147 - 0x93
    "10010000", --  622 - 0x26e  :  144 - 0x90
    "10010001", --  623 - 0x26f  :  145 - 0x91
    "10010000", --  624 - 0x270  :  144 - 0x90
    "10010001", --  625 - 0x271  :  145 - 0x91
    "10010010", --  626 - 0x272  :  146 - 0x92
    "10010011", --  627 - 0x273  :  147 - 0x93
    "10010100", --  628 - 0x274  :  148 - 0x94
    "10010101", --  629 - 0x275  :  149 - 0x95
    "10010111", --  630 - 0x276  :  151 - 0x97
    "10010100", --  631 - 0x277  :  148 - 0x94
    "10010110", --  632 - 0x278  :  150 - 0x96
    "10010101", --  633 - 0x279  :  149 - 0x95
    "10010110", --  634 - 0x27a  :  150 - 0x96
    "10010101", --  635 - 0x27b  :  149 - 0x95
    "10010000", --  636 - 0x27c  :  144 - 0x90
    "10010001", --  637 - 0x27d  :  145 - 0x91
    "10100111", --  638 - 0x27e  :  167 - 0xa7
    "10100000", --  639 - 0x27f  :  160 - 0xa0
    "10100000", --  640 - 0x280  :  160 - 0xa0 -- line 0x14
    "10100011", --  641 - 0x281  :  163 - 0xa3
    "10000010", --  642 - 0x282  :  130 - 0x82
    "10000011", --  643 - 0x283  :  131 - 0x83
    "10000110", --  644 - 0x284  :  134 - 0x86
    "10000111", --  645 - 0x285  :  135 - 0x87
    "10000100", --  646 - 0x286  :  132 - 0x84
    "10000101", --  647 - 0x287  :  133 - 0x85
    "10000100", --  648 - 0x288  :  132 - 0x84
    "10000111", --  649 - 0x289  :  135 - 0x87
    "10000100", --  650 - 0x28a  :  132 - 0x84
    "10000111", --  651 - 0x28b  :  135 - 0x87
    "10000110", --  652 - 0x28c  :  134 - 0x86
    "10000111", --  653 - 0x28d  :  135 - 0x87
    "10000100", --  654 - 0x28e  :  132 - 0x84
    "10000111", --  655 - 0x28f  :  135 - 0x87
    "10000110", --  656 - 0x290  :  134 - 0x86
    "10000111", --  657 - 0x291  :  135 - 0x87
    "10000110", --  658 - 0x292  :  134 - 0x86
    "10000111", --  659 - 0x293  :  135 - 0x87
    "10000110", --  660 - 0x294  :  134 - 0x86
    "10000111", --  661 - 0x295  :  135 - 0x87
    "10000110", --  662 - 0x296  :  134 - 0x86
    "10000111", --  663 - 0x297  :  135 - 0x87
    "10000101", --  664 - 0x298  :  133 - 0x85
    "10000110", --  665 - 0x299  :  134 - 0x86
    "10000100", --  666 - 0x29a  :  132 - 0x84
    "10000111", --  667 - 0x29b  :  135 - 0x87
    "10000000", --  668 - 0x29c  :  128 - 0x80
    "10000010", --  669 - 0x29d  :  130 - 0x82
    "10100111", --  670 - 0x29e  :  167 - 0xa7
    "10100000", --  671 - 0x29f  :  160 - 0xa0
    "10100000", --  672 - 0x2a0  :  160 - 0xa0 -- line 0x15
    "10100011", --  673 - 0x2a1  :  163 - 0xa3
    "10010010", --  674 - 0x2a2  :  146 - 0x92
    "10010011", --  675 - 0x2a3  :  147 - 0x93
    "10010110", --  676 - 0x2a4  :  150 - 0x96
    "10010111", --  677 - 0x2a5  :  151 - 0x97
    "10010100", --  678 - 0x2a6  :  148 - 0x94
    "10010101", --  679 - 0x2a7  :  149 - 0x95
    "10010110", --  680 - 0x2a8  :  150 - 0x96
    "10010101", --  681 - 0x2a9  :  149 - 0x95
    "10010110", --  682 - 0x2aa  :  150 - 0x96
    "10010101", --  683 - 0x2ab  :  149 - 0x95
    "10010110", --  684 - 0x2ac  :  150 - 0x96
    "10010111", --  685 - 0x2ad  :  151 - 0x97
    "10010110", --  686 - 0x2ae  :  150 - 0x96
    "10010101", --  687 - 0x2af  :  149 - 0x95
    "10010110", --  688 - 0x2b0  :  150 - 0x96
    "10010111", --  689 - 0x2b1  :  151 - 0x97
    "10010110", --  690 - 0x2b2  :  150 - 0x96
    "10010111", --  691 - 0x2b3  :  151 - 0x97
    "10010110", --  692 - 0x2b4  :  150 - 0x96
    "10010111", --  693 - 0x2b5  :  151 - 0x97
    "10010110", --  694 - 0x2b6  :  150 - 0x96
    "10010111", --  695 - 0x2b7  :  151 - 0x97
    "10010111", --  696 - 0x2b8  :  151 - 0x97
    "10010100", --  697 - 0x2b9  :  148 - 0x94
    "10010110", --  698 - 0x2ba  :  150 - 0x96
    "10010101", --  699 - 0x2bb  :  149 - 0x95
    "10010010", --  700 - 0x2bc  :  146 - 0x92
    "10010001", --  701 - 0x2bd  :  145 - 0x91
    "10100111", --  702 - 0x2be  :  167 - 0xa7
    "10100000", --  703 - 0x2bf  :  160 - 0xa0
    "10100000", --  704 - 0x2c0  :  160 - 0xa0 -- line 0x16
    "10100011", --  705 - 0x2c1  :  163 - 0xa3
    "10000000", --  706 - 0x2c2  :  128 - 0x80
    "10000001", --  707 - 0x2c3  :  129 - 0x81
    "10000101", --  708 - 0x2c4  :  133 - 0x85
    "10000110", --  709 - 0x2c5  :  134 - 0x86
    "10000100", --  710 - 0x2c6  :  132 - 0x84
    "10000101", --  711 - 0x2c7  :  133 - 0x85
    "10000100", --  712 - 0x2c8  :  132 - 0x84
    "10000101", --  713 - 0x2c9  :  133 - 0x85
    "10000100", --  714 - 0x2ca  :  132 - 0x84
    "10000111", --  715 - 0x2cb  :  135 - 0x87
    "10000101", --  716 - 0x2cc  :  133 - 0x85
    "10000110", --  717 - 0x2cd  :  134 - 0x86
    "10000110", --  718 - 0x2ce  :  134 - 0x86
    "10000111", --  719 - 0x2cf  :  135 - 0x87
    "10000110", --  720 - 0x2d0  :  134 - 0x86
    "10000111", --  721 - 0x2d1  :  135 - 0x87
    "10000101", --  722 - 0x2d2  :  133 - 0x85
    "10000110", --  723 - 0x2d3  :  134 - 0x86
    "10000101", --  724 - 0x2d4  :  133 - 0x85
    "10000110", --  725 - 0x2d5  :  134 - 0x86
    "10000110", --  726 - 0x2d6  :  134 - 0x86
    "10000111", --  727 - 0x2d7  :  135 - 0x87
    "10000100", --  728 - 0x2d8  :  132 - 0x84
    "10000111", --  729 - 0x2d9  :  135 - 0x87
    "10000100", --  730 - 0x2da  :  132 - 0x84
    "10000111", --  731 - 0x2db  :  135 - 0x87
    "10000000", --  732 - 0x2dc  :  128 - 0x80
    "10000001", --  733 - 0x2dd  :  129 - 0x81
    "10100111", --  734 - 0x2de  :  167 - 0xa7
    "10100000", --  735 - 0x2df  :  160 - 0xa0
    "10100000", --  736 - 0x2e0  :  160 - 0xa0 -- line 0x17
    "10100011", --  737 - 0x2e1  :  163 - 0xa3
    "10010000", --  738 - 0x2e2  :  144 - 0x90
    "10010001", --  739 - 0x2e3  :  145 - 0x91
    "10010111", --  740 - 0x2e4  :  151 - 0x97
    "10010100", --  741 - 0x2e5  :  148 - 0x94
    "10010100", --  742 - 0x2e6  :  148 - 0x94
    "10010101", --  743 - 0x2e7  :  149 - 0x95
    "10010100", --  744 - 0x2e8  :  148 - 0x94
    "10010101", --  745 - 0x2e9  :  149 - 0x95
    "10010110", --  746 - 0x2ea  :  150 - 0x96
    "10010101", --  747 - 0x2eb  :  149 - 0x95
    "10010111", --  748 - 0x2ec  :  151 - 0x97
    "10010100", --  749 - 0x2ed  :  148 - 0x94
    "10010110", --  750 - 0x2ee  :  150 - 0x96
    "10010111", --  751 - 0x2ef  :  151 - 0x97
    "10010110", --  752 - 0x2f0  :  150 - 0x96
    "10010111", --  753 - 0x2f1  :  151 - 0x97
    "10010111", --  754 - 0x2f2  :  151 - 0x97
    "10010100", --  755 - 0x2f3  :  148 - 0x94
    "10010111", --  756 - 0x2f4  :  151 - 0x97
    "10010100", --  757 - 0x2f5  :  148 - 0x94
    "10010110", --  758 - 0x2f6  :  150 - 0x96
    "10010111", --  759 - 0x2f7  :  151 - 0x97
    "10010110", --  760 - 0x2f8  :  150 - 0x96
    "10010101", --  761 - 0x2f9  :  149 - 0x95
    "10010110", --  762 - 0x2fa  :  150 - 0x96
    "10010101", --  763 - 0x2fb  :  149 - 0x95
    "10010000", --  764 - 0x2fc  :  144 - 0x90
    "10010001", --  765 - 0x2fd  :  145 - 0x91
    "10100111", --  766 - 0x2fe  :  167 - 0xa7
    "10100000", --  767 - 0x2ff  :  160 - 0xa0
    "10100000", --  768 - 0x300  :  160 - 0xa0 -- line 0x18
    "10100011", --  769 - 0x301  :  163 - 0xa3
    "10000000", --  770 - 0x302  :  128 - 0x80
    "10000010", --  771 - 0x303  :  130 - 0x82
    "10000100", --  772 - 0x304  :  132 - 0x84
    "10000111", --  773 - 0x305  :  135 - 0x87
    "10000100", --  774 - 0x306  :  132 - 0x84
    "10000111", --  775 - 0x307  :  135 - 0x87
    "10000100", --  776 - 0x308  :  132 - 0x84
    "10000111", --  777 - 0x309  :  135 - 0x87
    "10000110", --  778 - 0x30a  :  134 - 0x86
    "10000111", --  779 - 0x30b  :  135 - 0x87
    "10000101", --  780 - 0x30c  :  133 - 0x85
    "10000110", --  781 - 0x30d  :  134 - 0x86
    "10000100", --  782 - 0x30e  :  132 - 0x84
    "10000111", --  783 - 0x30f  :  135 - 0x87
    "10000100", --  784 - 0x310  :  132 - 0x84
    "10000101", --  785 - 0x311  :  133 - 0x85
    "10000100", --  786 - 0x312  :  132 - 0x84
    "10000111", --  787 - 0x313  :  135 - 0x87
    "10000110", --  788 - 0x314  :  134 - 0x86
    "10000111", --  789 - 0x315  :  135 - 0x87
    "10000110", --  790 - 0x316  :  134 - 0x86
    "10000111", --  791 - 0x317  :  135 - 0x87
    "10000100", --  792 - 0x318  :  132 - 0x84
    "10000111", --  793 - 0x319  :  135 - 0x87
    "10000101", --  794 - 0x31a  :  133 - 0x85
    "10000110", --  795 - 0x31b  :  134 - 0x86
    "10000000", --  796 - 0x31c  :  128 - 0x80
    "10000010", --  797 - 0x31d  :  130 - 0x82
    "10100111", --  798 - 0x31e  :  167 - 0xa7
    "10100000", --  799 - 0x31f  :  160 - 0xa0
    "10100000", --  800 - 0x320  :  160 - 0xa0 -- line 0x19
    "10100011", --  801 - 0x321  :  163 - 0xa3
    "10010010", --  802 - 0x322  :  146 - 0x92
    "10010001", --  803 - 0x323  :  145 - 0x91
    "10010110", --  804 - 0x324  :  150 - 0x96
    "10010101", --  805 - 0x325  :  149 - 0x95
    "10010110", --  806 - 0x326  :  150 - 0x96
    "10010101", --  807 - 0x327  :  149 - 0x95
    "10010110", --  808 - 0x328  :  150 - 0x96
    "10010101", --  809 - 0x329  :  149 - 0x95
    "10010110", --  810 - 0x32a  :  150 - 0x96
    "10010111", --  811 - 0x32b  :  151 - 0x97
    "10010111", --  812 - 0x32c  :  151 - 0x97
    "10010100", --  813 - 0x32d  :  148 - 0x94
    "10010110", --  814 - 0x32e  :  150 - 0x96
    "10010101", --  815 - 0x32f  :  149 - 0x95
    "10010100", --  816 - 0x330  :  148 - 0x94
    "10010101", --  817 - 0x331  :  149 - 0x95
    "10010110", --  818 - 0x332  :  150 - 0x96
    "10010101", --  819 - 0x333  :  149 - 0x95
    "10010110", --  820 - 0x334  :  150 - 0x96
    "10010111", --  821 - 0x335  :  151 - 0x97
    "10010110", --  822 - 0x336  :  150 - 0x96
    "10010111", --  823 - 0x337  :  151 - 0x97
    "10010110", --  824 - 0x338  :  150 - 0x96
    "10010101", --  825 - 0x339  :  149 - 0x95
    "10010111", --  826 - 0x33a  :  151 - 0x97
    "10010100", --  827 - 0x33b  :  148 - 0x94
    "10010010", --  828 - 0x33c  :  146 - 0x92
    "10010001", --  829 - 0x33d  :  145 - 0x91
    "10100111", --  830 - 0x33e  :  167 - 0xa7
    "10100000", --  831 - 0x33f  :  160 - 0xa0
    "10100000", --  832 - 0x340  :  160 - 0xa0 -- line 0x1a
    "10100011", --  833 - 0x341  :  163 - 0xa3
    "10000001", --  834 - 0x342  :  129 - 0x81
    "10000000", --  835 - 0x343  :  128 - 0x80
    "10000000", --  836 - 0x344  :  128 - 0x80
    "10000001", --  837 - 0x345  :  129 - 0x81
    "10000010", --  838 - 0x346  :  130 - 0x82
    "10000011", --  839 - 0x347  :  131 - 0x83
    "10000001", --  840 - 0x348  :  129 - 0x81
    "10000000", --  841 - 0x349  :  128 - 0x80
    "10000001", --  842 - 0x34a  :  129 - 0x81
    "10000000", --  843 - 0x34b  :  128 - 0x80
    "10000000", --  844 - 0x34c  :  128 - 0x80
    "10000010", --  845 - 0x34d  :  130 - 0x82
    "10000000", --  846 - 0x34e  :  128 - 0x80
    "10000001", --  847 - 0x34f  :  129 - 0x81
    "10000001", --  848 - 0x350  :  129 - 0x81
    "10000000", --  849 - 0x351  :  128 - 0x80
    "10000000", --  850 - 0x352  :  128 - 0x80
    "10000010", --  851 - 0x353  :  130 - 0x82
    "10000000", --  852 - 0x354  :  128 - 0x80
    "10000001", --  853 - 0x355  :  129 - 0x81
    "10000010", --  854 - 0x356  :  130 - 0x82
    "10000011", --  855 - 0x357  :  131 - 0x83
    "10000001", --  856 - 0x358  :  129 - 0x81
    "10000000", --  857 - 0x359  :  128 - 0x80
    "10000000", --  858 - 0x35a  :  128 - 0x80
    "10000001", --  859 - 0x35b  :  129 - 0x81
    "10000000", --  860 - 0x35c  :  128 - 0x80
    "10000001", --  861 - 0x35d  :  129 - 0x81
    "10100111", --  862 - 0x35e  :  167 - 0xa7
    "10100000", --  863 - 0x35f  :  160 - 0xa0
    "10100000", --  864 - 0x360  :  160 - 0xa0 -- line 0x1b
    "10100011", --  865 - 0x361  :  163 - 0xa3
    "10010011", --  866 - 0x362  :  147 - 0x93
    "10010010", --  867 - 0x363  :  146 - 0x92
    "10010000", --  868 - 0x364  :  144 - 0x90
    "10010001", --  869 - 0x365  :  145 - 0x91
    "10010010", --  870 - 0x366  :  146 - 0x92
    "10010011", --  871 - 0x367  :  147 - 0x93
    "10010011", --  872 - 0x368  :  147 - 0x93
    "10010010", --  873 - 0x369  :  146 - 0x92
    "10010011", --  874 - 0x36a  :  147 - 0x93
    "10010010", --  875 - 0x36b  :  146 - 0x92
    "10010010", --  876 - 0x36c  :  146 - 0x92
    "10010001", --  877 - 0x36d  :  145 - 0x91
    "10010000", --  878 - 0x36e  :  144 - 0x90
    "10010001", --  879 - 0x36f  :  145 - 0x91
    "10010011", --  880 - 0x370  :  147 - 0x93
    "10010010", --  881 - 0x371  :  146 - 0x92
    "10010010", --  882 - 0x372  :  146 - 0x92
    "10010001", --  883 - 0x373  :  145 - 0x91
    "10010000", --  884 - 0x374  :  144 - 0x90
    "10010001", --  885 - 0x375  :  145 - 0x91
    "10010010", --  886 - 0x376  :  146 - 0x92
    "10010011", --  887 - 0x377  :  147 - 0x93
    "10010011", --  888 - 0x378  :  147 - 0x93
    "10010010", --  889 - 0x379  :  146 - 0x92
    "10010000", --  890 - 0x37a  :  144 - 0x90
    "10010001", --  891 - 0x37b  :  145 - 0x91
    "10010000", --  892 - 0x37c  :  144 - 0x90
    "10010001", --  893 - 0x37d  :  145 - 0x91
    "10100111", --  894 - 0x37e  :  167 - 0xa7
    "10100000", --  895 - 0x37f  :  160 - 0xa0
    "10100000", --  896 - 0x380  :  160 - 0xa0 -- line 0x1c
    "10100100", --  897 - 0x381  :  164 - 0xa4
    "10100101", --  898 - 0x382  :  165 - 0xa5
    "10100101", --  899 - 0x383  :  165 - 0xa5
    "10100101", --  900 - 0x384  :  165 - 0xa5
    "10100101", --  901 - 0x385  :  165 - 0xa5
    "10100101", --  902 - 0x386  :  165 - 0xa5
    "10100101", --  903 - 0x387  :  165 - 0xa5
    "10100101", --  904 - 0x388  :  165 - 0xa5
    "10100101", --  905 - 0x389  :  165 - 0xa5
    "10100101", --  906 - 0x38a  :  165 - 0xa5
    "10100101", --  907 - 0x38b  :  165 - 0xa5
    "10100101", --  908 - 0x38c  :  165 - 0xa5
    "10100101", --  909 - 0x38d  :  165 - 0xa5
    "10100101", --  910 - 0x38e  :  165 - 0xa5
    "10100101", --  911 - 0x38f  :  165 - 0xa5
    "10100101", --  912 - 0x390  :  165 - 0xa5
    "10100101", --  913 - 0x391  :  165 - 0xa5
    "10100101", --  914 - 0x392  :  165 - 0xa5
    "10100101", --  915 - 0x393  :  165 - 0xa5
    "10100101", --  916 - 0x394  :  165 - 0xa5
    "10100101", --  917 - 0x395  :  165 - 0xa5
    "10100101", --  918 - 0x396  :  165 - 0xa5
    "10100101", --  919 - 0x397  :  165 - 0xa5
    "10100101", --  920 - 0x398  :  165 - 0xa5
    "10100101", --  921 - 0x399  :  165 - 0xa5
    "10100101", --  922 - 0x39a  :  165 - 0xa5
    "10100101", --  923 - 0x39b  :  165 - 0xa5
    "10100101", --  924 - 0x39c  :  165 - 0xa5
    "10100101", --  925 - 0x39d  :  165 - 0xa5
    "10101000", --  926 - 0x39e  :  168 - 0xa8
    "10100000", --  927 - 0x39f  :  160 - 0xa0
    "10100000", --  928 - 0x3a0  :  160 - 0xa0 -- line 0x1d
    "10100000", --  929 - 0x3a1  :  160 - 0xa0
    "10100000", --  930 - 0x3a2  :  160 - 0xa0
    "10100000", --  931 - 0x3a3  :  160 - 0xa0
    "10100000", --  932 - 0x3a4  :  160 - 0xa0
    "10100000", --  933 - 0x3a5  :  160 - 0xa0
    "10100000", --  934 - 0x3a6  :  160 - 0xa0
    "10100000", --  935 - 0x3a7  :  160 - 0xa0
    "10100000", --  936 - 0x3a8  :  160 - 0xa0
    "10100000", --  937 - 0x3a9  :  160 - 0xa0
    "10100000", --  938 - 0x3aa  :  160 - 0xa0
    "10100000", --  939 - 0x3ab  :  160 - 0xa0
    "10100000", --  940 - 0x3ac  :  160 - 0xa0
    "10100000", --  941 - 0x3ad  :  160 - 0xa0
    "10100000", --  942 - 0x3ae  :  160 - 0xa0
    "10100000", --  943 - 0x3af  :  160 - 0xa0
    "10100000", --  944 - 0x3b0  :  160 - 0xa0
    "10100000", --  945 - 0x3b1  :  160 - 0xa0
    "10100000", --  946 - 0x3b2  :  160 - 0xa0
    "10100000", --  947 - 0x3b3  :  160 - 0xa0
    "10100000", --  948 - 0x3b4  :  160 - 0xa0
    "10100000", --  949 - 0x3b5  :  160 - 0xa0
    "10100000", --  950 - 0x3b6  :  160 - 0xa0
    "10100000", --  951 - 0x3b7  :  160 - 0xa0
    "10100000", --  952 - 0x3b8  :  160 - 0xa0
    "10100000", --  953 - 0x3b9  :  160 - 0xa0
    "10100000", --  954 - 0x3ba  :  160 - 0xa0
    "10100000", --  955 - 0x3bb  :  160 - 0xa0
    "10100000", --  956 - 0x3bc  :  160 - 0xa0
    "10100000", --  957 - 0x3bd  :  160 - 0xa0
    "10100000", --  958 - 0x3be  :  160 - 0xa0
    "10100000", --  959 - 0x3bf  :  160 - 0xa0
        ---- Attribute Table 0----
    "00000000", --  960 - 0x3c0  :    0 - 0x0
    "00000000", --  961 - 0x3c1  :    0 - 0x0
    "00000000", --  962 - 0x3c2  :    0 - 0x0
    "00000000", --  963 - 0x3c3  :    0 - 0x0
    "00000000", --  964 - 0x3c4  :    0 - 0x0
    "00000000", --  965 - 0x3c5  :    0 - 0x0
    "00000000", --  966 - 0x3c6  :    0 - 0x0
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "10000000", --  968 - 0x3c8  :  128 - 0x80
    "10100000", --  969 - 0x3c9  :  160 - 0xa0
    "10100000", --  970 - 0x3ca  :  160 - 0xa0
    "10100000", --  971 - 0x3cb  :  160 - 0xa0
    "10100000", --  972 - 0x3cc  :  160 - 0xa0
    "10100000", --  973 - 0x3cd  :  160 - 0xa0
    "10100000", --  974 - 0x3ce  :  160 - 0xa0
    "00100000", --  975 - 0x3cf  :   32 - 0x20
    "10001000", --  976 - 0x3d0  :  136 - 0x88
    "10101010", --  977 - 0x3d1  :  170 - 0xaa
    "10101010", --  978 - 0x3d2  :  170 - 0xaa
    "10101010", --  979 - 0x3d3  :  170 - 0xaa
    "10101010", --  980 - 0x3d4  :  170 - 0xaa
    "10101010", --  981 - 0x3d5  :  170 - 0xaa
    "10101010", --  982 - 0x3d6  :  170 - 0xaa
    "00100010", --  983 - 0x3d7  :   34 - 0x22
    "10001000", --  984 - 0x3d8  :  136 - 0x88
    "10101010", --  985 - 0x3d9  :  170 - 0xaa
    "10101010", --  986 - 0x3da  :  170 - 0xaa
    "10101010", --  987 - 0x3db  :  170 - 0xaa
    "10101010", --  988 - 0x3dc  :  170 - 0xaa
    "10101010", --  989 - 0x3dd  :  170 - 0xaa
    "10101010", --  990 - 0x3de  :  170 - 0xaa
    "00100010", --  991 - 0x3df  :   34 - 0x22
    "10001000", --  992 - 0x3e0  :  136 - 0x88
    "10101010", --  993 - 0x3e1  :  170 - 0xaa
    "10101010", --  994 - 0x3e2  :  170 - 0xaa
    "10101010", --  995 - 0x3e3  :  170 - 0xaa
    "10101010", --  996 - 0x3e4  :  170 - 0xaa
    "10101010", --  997 - 0x3e5  :  170 - 0xaa
    "10101010", --  998 - 0x3e6  :  170 - 0xaa
    "00100010", --  999 - 0x3e7  :   34 - 0x22
    "10001000", -- 1000 - 0x3e8  :  136 - 0x88
    "10101010", -- 1001 - 0x3e9  :  170 - 0xaa
    "10101010", -- 1002 - 0x3ea  :  170 - 0xaa
    "10101010", -- 1003 - 0x3eb  :  170 - 0xaa
    "10101010", -- 1004 - 0x3ec  :  170 - 0xaa
    "10101010", -- 1005 - 0x3ed  :  170 - 0xaa
    "10101010", -- 1006 - 0x3ee  :  170 - 0xaa
    "00100010", -- 1007 - 0x3ef  :   34 - 0x22
    "10001000", -- 1008 - 0x3f0  :  136 - 0x88
    "10101010", -- 1009 - 0x3f1  :  170 - 0xaa
    "10101010", -- 1010 - 0x3f2  :  170 - 0xaa
    "10101010", -- 1011 - 0x3f3  :  170 - 0xaa
    "10101010", -- 1012 - 0x3f4  :  170 - 0xaa
    "10101010", -- 1013 - 0x3f5  :  170 - 0xaa
    "10101010", -- 1014 - 0x3f6  :  170 - 0xaa
    "00100010", -- 1015 - 0x3f7  :   34 - 0x22
    "00000000", -- 1016 - 0x3f8  :    0 - 0x0
    "00000000", -- 1017 - 0x3f9  :    0 - 0x0
    "00000000", -- 1018 - 0x3fa  :    0 - 0x0
    "00000000", -- 1019 - 0x3fb  :    0 - 0x0
    "00000000", -- 1020 - 0x3fc  :    0 - 0x0
    "00000000", -- 1021 - 0x3fd  :    0 - 0x0
    "00000000", -- 1022 - 0x3fe  :    0 - 0x0
    "00000000", -- 1023 - 0x3ff  :    0 - 0x0
     ------- Name Table 1---------
    "00000000", -- 1024 - 0x400  :    0 - 0x0 -- line 0x0
    "00000000", -- 1025 - 0x401  :    0 - 0x0
    "00000000", -- 1026 - 0x402  :    0 - 0x0
    "00000000", -- 1027 - 0x403  :    0 - 0x0
    "00000000", -- 1028 - 0x404  :    0 - 0x0
    "00000000", -- 1029 - 0x405  :    0 - 0x0
    "00000000", -- 1030 - 0x406  :    0 - 0x0
    "00000000", -- 1031 - 0x407  :    0 - 0x0
    "00000000", -- 1032 - 0x408  :    0 - 0x0
    "00000000", -- 1033 - 0x409  :    0 - 0x0
    "00000000", -- 1034 - 0x40a  :    0 - 0x0
    "00000000", -- 1035 - 0x40b  :    0 - 0x0
    "00000000", -- 1036 - 0x40c  :    0 - 0x0
    "00000000", -- 1037 - 0x40d  :    0 - 0x0
    "00000000", -- 1038 - 0x40e  :    0 - 0x0
    "00000000", -- 1039 - 0x40f  :    0 - 0x0
    "00000000", -- 1040 - 0x410  :    0 - 0x0
    "00000000", -- 1041 - 0x411  :    0 - 0x0
    "00000000", -- 1042 - 0x412  :    0 - 0x0
    "00000000", -- 1043 - 0x413  :    0 - 0x0
    "00000000", -- 1044 - 0x414  :    0 - 0x0
    "00000000", -- 1045 - 0x415  :    0 - 0x0
    "00000000", -- 1046 - 0x416  :    0 - 0x0
    "00000000", -- 1047 - 0x417  :    0 - 0x0
    "00000000", -- 1048 - 0x418  :    0 - 0x0
    "00000000", -- 1049 - 0x419  :    0 - 0x0
    "00000000", -- 1050 - 0x41a  :    0 - 0x0
    "00000000", -- 1051 - 0x41b  :    0 - 0x0
    "00000000", -- 1052 - 0x41c  :    0 - 0x0
    "00000000", -- 1053 - 0x41d  :    0 - 0x0
    "00000000", -- 1054 - 0x41e  :    0 - 0x0
    "00000000", -- 1055 - 0x41f  :    0 - 0x0
    "00000000", -- 1056 - 0x420  :    0 - 0x0 -- line 0x1
    "00000000", -- 1057 - 0x421  :    0 - 0x0
    "00000000", -- 1058 - 0x422  :    0 - 0x0
    "00000000", -- 1059 - 0x423  :    0 - 0x0
    "00000000", -- 1060 - 0x424  :    0 - 0x0
    "00000000", -- 1061 - 0x425  :    0 - 0x0
    "00000000", -- 1062 - 0x426  :    0 - 0x0
    "00000000", -- 1063 - 0x427  :    0 - 0x0
    "00000000", -- 1064 - 0x428  :    0 - 0x0
    "00000000", -- 1065 - 0x429  :    0 - 0x0
    "00000000", -- 1066 - 0x42a  :    0 - 0x0
    "00000000", -- 1067 - 0x42b  :    0 - 0x0
    "00000000", -- 1068 - 0x42c  :    0 - 0x0
    "00000000", -- 1069 - 0x42d  :    0 - 0x0
    "00000000", -- 1070 - 0x42e  :    0 - 0x0
    "00000000", -- 1071 - 0x42f  :    0 - 0x0
    "00000000", -- 1072 - 0x430  :    0 - 0x0
    "00000000", -- 1073 - 0x431  :    0 - 0x0
    "00000000", -- 1074 - 0x432  :    0 - 0x0
    "00000000", -- 1075 - 0x433  :    0 - 0x0
    "00000000", -- 1076 - 0x434  :    0 - 0x0
    "00000000", -- 1077 - 0x435  :    0 - 0x0
    "00000000", -- 1078 - 0x436  :    0 - 0x0
    "00000000", -- 1079 - 0x437  :    0 - 0x0
    "00000000", -- 1080 - 0x438  :    0 - 0x0
    "00000000", -- 1081 - 0x439  :    0 - 0x0
    "00000000", -- 1082 - 0x43a  :    0 - 0x0
    "00000000", -- 1083 - 0x43b  :    0 - 0x0
    "00000000", -- 1084 - 0x43c  :    0 - 0x0
    "00000000", -- 1085 - 0x43d  :    0 - 0x0
    "00000000", -- 1086 - 0x43e  :    0 - 0x0
    "00000000", -- 1087 - 0x43f  :    0 - 0x0
    "00000000", -- 1088 - 0x440  :    0 - 0x0 -- line 0x2
    "00000000", -- 1089 - 0x441  :    0 - 0x0
    "00000000", -- 1090 - 0x442  :    0 - 0x0
    "00000000", -- 1091 - 0x443  :    0 - 0x0
    "00000000", -- 1092 - 0x444  :    0 - 0x0
    "00000000", -- 1093 - 0x445  :    0 - 0x0
    "00000000", -- 1094 - 0x446  :    0 - 0x0
    "00000000", -- 1095 - 0x447  :    0 - 0x0
    "00000000", -- 1096 - 0x448  :    0 - 0x0
    "00000000", -- 1097 - 0x449  :    0 - 0x0
    "00000000", -- 1098 - 0x44a  :    0 - 0x0
    "00000000", -- 1099 - 0x44b  :    0 - 0x0
    "00000000", -- 1100 - 0x44c  :    0 - 0x0
    "00000000", -- 1101 - 0x44d  :    0 - 0x0
    "00000000", -- 1102 - 0x44e  :    0 - 0x0
    "00000000", -- 1103 - 0x44f  :    0 - 0x0
    "00000000", -- 1104 - 0x450  :    0 - 0x0
    "00000000", -- 1105 - 0x451  :    0 - 0x0
    "00000000", -- 1106 - 0x452  :    0 - 0x0
    "00000000", -- 1107 - 0x453  :    0 - 0x0
    "00000000", -- 1108 - 0x454  :    0 - 0x0
    "00000000", -- 1109 - 0x455  :    0 - 0x0
    "00000000", -- 1110 - 0x456  :    0 - 0x0
    "00000000", -- 1111 - 0x457  :    0 - 0x0
    "00000000", -- 1112 - 0x458  :    0 - 0x0
    "00000000", -- 1113 - 0x459  :    0 - 0x0
    "00000000", -- 1114 - 0x45a  :    0 - 0x0
    "00000000", -- 1115 - 0x45b  :    0 - 0x0
    "00000000", -- 1116 - 0x45c  :    0 - 0x0
    "00000000", -- 1117 - 0x45d  :    0 - 0x0
    "00000000", -- 1118 - 0x45e  :    0 - 0x0
    "00000000", -- 1119 - 0x45f  :    0 - 0x0
    "00000000", -- 1120 - 0x460  :    0 - 0x0 -- line 0x3
    "00000000", -- 1121 - 0x461  :    0 - 0x0
    "00000000", -- 1122 - 0x462  :    0 - 0x0
    "00000000", -- 1123 - 0x463  :    0 - 0x0
    "00000000", -- 1124 - 0x464  :    0 - 0x0
    "00000000", -- 1125 - 0x465  :    0 - 0x0
    "00000000", -- 1126 - 0x466  :    0 - 0x0
    "00000000", -- 1127 - 0x467  :    0 - 0x0
    "00000000", -- 1128 - 0x468  :    0 - 0x0
    "00000000", -- 1129 - 0x469  :    0 - 0x0
    "00000000", -- 1130 - 0x46a  :    0 - 0x0
    "00000000", -- 1131 - 0x46b  :    0 - 0x0
    "00000000", -- 1132 - 0x46c  :    0 - 0x0
    "00000000", -- 1133 - 0x46d  :    0 - 0x0
    "00000000", -- 1134 - 0x46e  :    0 - 0x0
    "00000000", -- 1135 - 0x46f  :    0 - 0x0
    "00000000", -- 1136 - 0x470  :    0 - 0x0
    "00000000", -- 1137 - 0x471  :    0 - 0x0
    "00000000", -- 1138 - 0x472  :    0 - 0x0
    "00000000", -- 1139 - 0x473  :    0 - 0x0
    "00000000", -- 1140 - 0x474  :    0 - 0x0
    "00000000", -- 1141 - 0x475  :    0 - 0x0
    "00000000", -- 1142 - 0x476  :    0 - 0x0
    "00000000", -- 1143 - 0x477  :    0 - 0x0
    "00000000", -- 1144 - 0x478  :    0 - 0x0
    "00000000", -- 1145 - 0x479  :    0 - 0x0
    "00000000", -- 1146 - 0x47a  :    0 - 0x0
    "00000000", -- 1147 - 0x47b  :    0 - 0x0
    "00000000", -- 1148 - 0x47c  :    0 - 0x0
    "00000000", -- 1149 - 0x47d  :    0 - 0x0
    "00000000", -- 1150 - 0x47e  :    0 - 0x0
    "00000000", -- 1151 - 0x47f  :    0 - 0x0
    "00000000", -- 1152 - 0x480  :    0 - 0x0 -- line 0x4
    "00000000", -- 1153 - 0x481  :    0 - 0x0
    "00000000", -- 1154 - 0x482  :    0 - 0x0
    "00000000", -- 1155 - 0x483  :    0 - 0x0
    "00000000", -- 1156 - 0x484  :    0 - 0x0
    "00000000", -- 1157 - 0x485  :    0 - 0x0
    "00000000", -- 1158 - 0x486  :    0 - 0x0
    "00000000", -- 1159 - 0x487  :    0 - 0x0
    "00000000", -- 1160 - 0x488  :    0 - 0x0
    "00000000", -- 1161 - 0x489  :    0 - 0x0
    "00000000", -- 1162 - 0x48a  :    0 - 0x0
    "00000000", -- 1163 - 0x48b  :    0 - 0x0
    "00000000", -- 1164 - 0x48c  :    0 - 0x0
    "00000000", -- 1165 - 0x48d  :    0 - 0x0
    "00000000", -- 1166 - 0x48e  :    0 - 0x0
    "00000000", -- 1167 - 0x48f  :    0 - 0x0
    "00000000", -- 1168 - 0x490  :    0 - 0x0
    "00000000", -- 1169 - 0x491  :    0 - 0x0
    "00000000", -- 1170 - 0x492  :    0 - 0x0
    "00000000", -- 1171 - 0x493  :    0 - 0x0
    "00000000", -- 1172 - 0x494  :    0 - 0x0
    "00000000", -- 1173 - 0x495  :    0 - 0x0
    "00000000", -- 1174 - 0x496  :    0 - 0x0
    "00000000", -- 1175 - 0x497  :    0 - 0x0
    "00000000", -- 1176 - 0x498  :    0 - 0x0
    "00000000", -- 1177 - 0x499  :    0 - 0x0
    "00000000", -- 1178 - 0x49a  :    0 - 0x0
    "00000000", -- 1179 - 0x49b  :    0 - 0x0
    "00000000", -- 1180 - 0x49c  :    0 - 0x0
    "00000000", -- 1181 - 0x49d  :    0 - 0x0
    "00000000", -- 1182 - 0x49e  :    0 - 0x0
    "00000000", -- 1183 - 0x49f  :    0 - 0x0
    "00000000", -- 1184 - 0x4a0  :    0 - 0x0 -- line 0x5
    "00000000", -- 1185 - 0x4a1  :    0 - 0x0
    "00000000", -- 1186 - 0x4a2  :    0 - 0x0
    "00000000", -- 1187 - 0x4a3  :    0 - 0x0
    "00000000", -- 1188 - 0x4a4  :    0 - 0x0
    "00000000", -- 1189 - 0x4a5  :    0 - 0x0
    "00000000", -- 1190 - 0x4a6  :    0 - 0x0
    "00000000", -- 1191 - 0x4a7  :    0 - 0x0
    "00000000", -- 1192 - 0x4a8  :    0 - 0x0
    "00000000", -- 1193 - 0x4a9  :    0 - 0x0
    "00000000", -- 1194 - 0x4aa  :    0 - 0x0
    "00000000", -- 1195 - 0x4ab  :    0 - 0x0
    "00000000", -- 1196 - 0x4ac  :    0 - 0x0
    "00000000", -- 1197 - 0x4ad  :    0 - 0x0
    "00000000", -- 1198 - 0x4ae  :    0 - 0x0
    "00000000", -- 1199 - 0x4af  :    0 - 0x0
    "00000000", -- 1200 - 0x4b0  :    0 - 0x0
    "00000000", -- 1201 - 0x4b1  :    0 - 0x0
    "00000000", -- 1202 - 0x4b2  :    0 - 0x0
    "00000000", -- 1203 - 0x4b3  :    0 - 0x0
    "00000000", -- 1204 - 0x4b4  :    0 - 0x0
    "00000000", -- 1205 - 0x4b5  :    0 - 0x0
    "00000000", -- 1206 - 0x4b6  :    0 - 0x0
    "00000000", -- 1207 - 0x4b7  :    0 - 0x0
    "00000000", -- 1208 - 0x4b8  :    0 - 0x0
    "00000000", -- 1209 - 0x4b9  :    0 - 0x0
    "00000000", -- 1210 - 0x4ba  :    0 - 0x0
    "00000000", -- 1211 - 0x4bb  :    0 - 0x0
    "00000000", -- 1212 - 0x4bc  :    0 - 0x0
    "00000000", -- 1213 - 0x4bd  :    0 - 0x0
    "00000000", -- 1214 - 0x4be  :    0 - 0x0
    "00000000", -- 1215 - 0x4bf  :    0 - 0x0
    "00000000", -- 1216 - 0x4c0  :    0 - 0x0 -- line 0x6
    "00000000", -- 1217 - 0x4c1  :    0 - 0x0
    "00000000", -- 1218 - 0x4c2  :    0 - 0x0
    "00000000", -- 1219 - 0x4c3  :    0 - 0x0
    "00000000", -- 1220 - 0x4c4  :    0 - 0x0
    "00000000", -- 1221 - 0x4c5  :    0 - 0x0
    "00000000", -- 1222 - 0x4c6  :    0 - 0x0
    "00000000", -- 1223 - 0x4c7  :    0 - 0x0
    "00000000", -- 1224 - 0x4c8  :    0 - 0x0
    "00000000", -- 1225 - 0x4c9  :    0 - 0x0
    "00000000", -- 1226 - 0x4ca  :    0 - 0x0
    "00000000", -- 1227 - 0x4cb  :    0 - 0x0
    "00000000", -- 1228 - 0x4cc  :    0 - 0x0
    "00000000", -- 1229 - 0x4cd  :    0 - 0x0
    "00000000", -- 1230 - 0x4ce  :    0 - 0x0
    "00000000", -- 1231 - 0x4cf  :    0 - 0x0
    "00000000", -- 1232 - 0x4d0  :    0 - 0x0
    "00000000", -- 1233 - 0x4d1  :    0 - 0x0
    "00000000", -- 1234 - 0x4d2  :    0 - 0x0
    "00000000", -- 1235 - 0x4d3  :    0 - 0x0
    "00000000", -- 1236 - 0x4d4  :    0 - 0x0
    "00000000", -- 1237 - 0x4d5  :    0 - 0x0
    "00000000", -- 1238 - 0x4d6  :    0 - 0x0
    "00000000", -- 1239 - 0x4d7  :    0 - 0x0
    "00000000", -- 1240 - 0x4d8  :    0 - 0x0
    "00000000", -- 1241 - 0x4d9  :    0 - 0x0
    "00000000", -- 1242 - 0x4da  :    0 - 0x0
    "00000000", -- 1243 - 0x4db  :    0 - 0x0
    "00000000", -- 1244 - 0x4dc  :    0 - 0x0
    "00000000", -- 1245 - 0x4dd  :    0 - 0x0
    "00000000", -- 1246 - 0x4de  :    0 - 0x0
    "00000000", -- 1247 - 0x4df  :    0 - 0x0
    "00000000", -- 1248 - 0x4e0  :    0 - 0x0 -- line 0x7
    "00000000", -- 1249 - 0x4e1  :    0 - 0x0
    "00000000", -- 1250 - 0x4e2  :    0 - 0x0
    "00000000", -- 1251 - 0x4e3  :    0 - 0x0
    "00000000", -- 1252 - 0x4e4  :    0 - 0x0
    "00000000", -- 1253 - 0x4e5  :    0 - 0x0
    "00000000", -- 1254 - 0x4e6  :    0 - 0x0
    "00000000", -- 1255 - 0x4e7  :    0 - 0x0
    "00000000", -- 1256 - 0x4e8  :    0 - 0x0
    "00000000", -- 1257 - 0x4e9  :    0 - 0x0
    "00000000", -- 1258 - 0x4ea  :    0 - 0x0
    "00000000", -- 1259 - 0x4eb  :    0 - 0x0
    "00000000", -- 1260 - 0x4ec  :    0 - 0x0
    "00000000", -- 1261 - 0x4ed  :    0 - 0x0
    "00000000", -- 1262 - 0x4ee  :    0 - 0x0
    "00000000", -- 1263 - 0x4ef  :    0 - 0x0
    "00000000", -- 1264 - 0x4f0  :    0 - 0x0
    "00000000", -- 1265 - 0x4f1  :    0 - 0x0
    "00000000", -- 1266 - 0x4f2  :    0 - 0x0
    "00000000", -- 1267 - 0x4f3  :    0 - 0x0
    "00000000", -- 1268 - 0x4f4  :    0 - 0x0
    "00000000", -- 1269 - 0x4f5  :    0 - 0x0
    "00000000", -- 1270 - 0x4f6  :    0 - 0x0
    "00000000", -- 1271 - 0x4f7  :    0 - 0x0
    "00000000", -- 1272 - 0x4f8  :    0 - 0x0
    "00000000", -- 1273 - 0x4f9  :    0 - 0x0
    "00000000", -- 1274 - 0x4fa  :    0 - 0x0
    "00000000", -- 1275 - 0x4fb  :    0 - 0x0
    "00000000", -- 1276 - 0x4fc  :    0 - 0x0
    "00000000", -- 1277 - 0x4fd  :    0 - 0x0
    "00000000", -- 1278 - 0x4fe  :    0 - 0x0
    "00000000", -- 1279 - 0x4ff  :    0 - 0x0
    "00000000", -- 1280 - 0x500  :    0 - 0x0 -- line 0x8
    "00000000", -- 1281 - 0x501  :    0 - 0x0
    "00000000", -- 1282 - 0x502  :    0 - 0x0
    "00000000", -- 1283 - 0x503  :    0 - 0x0
    "00000000", -- 1284 - 0x504  :    0 - 0x0
    "00000000", -- 1285 - 0x505  :    0 - 0x0
    "00000000", -- 1286 - 0x506  :    0 - 0x0
    "00000000", -- 1287 - 0x507  :    0 - 0x0
    "00000000", -- 1288 - 0x508  :    0 - 0x0
    "00000000", -- 1289 - 0x509  :    0 - 0x0
    "00000000", -- 1290 - 0x50a  :    0 - 0x0
    "00000000", -- 1291 - 0x50b  :    0 - 0x0
    "00000000", -- 1292 - 0x50c  :    0 - 0x0
    "00000000", -- 1293 - 0x50d  :    0 - 0x0
    "00000000", -- 1294 - 0x50e  :    0 - 0x0
    "00000000", -- 1295 - 0x50f  :    0 - 0x0
    "00000000", -- 1296 - 0x510  :    0 - 0x0
    "00000000", -- 1297 - 0x511  :    0 - 0x0
    "00000000", -- 1298 - 0x512  :    0 - 0x0
    "00000000", -- 1299 - 0x513  :    0 - 0x0
    "00000000", -- 1300 - 0x514  :    0 - 0x0
    "00000000", -- 1301 - 0x515  :    0 - 0x0
    "00000000", -- 1302 - 0x516  :    0 - 0x0
    "00000000", -- 1303 - 0x517  :    0 - 0x0
    "00000000", -- 1304 - 0x518  :    0 - 0x0
    "00000000", -- 1305 - 0x519  :    0 - 0x0
    "00000000", -- 1306 - 0x51a  :    0 - 0x0
    "00000000", -- 1307 - 0x51b  :    0 - 0x0
    "00000000", -- 1308 - 0x51c  :    0 - 0x0
    "00000000", -- 1309 - 0x51d  :    0 - 0x0
    "00000000", -- 1310 - 0x51e  :    0 - 0x0
    "00000000", -- 1311 - 0x51f  :    0 - 0x0
    "00000000", -- 1312 - 0x520  :    0 - 0x0 -- line 0x9
    "00000000", -- 1313 - 0x521  :    0 - 0x0
    "00000000", -- 1314 - 0x522  :    0 - 0x0
    "00000000", -- 1315 - 0x523  :    0 - 0x0
    "00000000", -- 1316 - 0x524  :    0 - 0x0
    "00000000", -- 1317 - 0x525  :    0 - 0x0
    "00000000", -- 1318 - 0x526  :    0 - 0x0
    "00000000", -- 1319 - 0x527  :    0 - 0x0
    "00000000", -- 1320 - 0x528  :    0 - 0x0
    "00000000", -- 1321 - 0x529  :    0 - 0x0
    "00000000", -- 1322 - 0x52a  :    0 - 0x0
    "00000000", -- 1323 - 0x52b  :    0 - 0x0
    "00000000", -- 1324 - 0x52c  :    0 - 0x0
    "00000000", -- 1325 - 0x52d  :    0 - 0x0
    "00000000", -- 1326 - 0x52e  :    0 - 0x0
    "00000000", -- 1327 - 0x52f  :    0 - 0x0
    "00000000", -- 1328 - 0x530  :    0 - 0x0
    "00000000", -- 1329 - 0x531  :    0 - 0x0
    "00000000", -- 1330 - 0x532  :    0 - 0x0
    "00000000", -- 1331 - 0x533  :    0 - 0x0
    "00000000", -- 1332 - 0x534  :    0 - 0x0
    "00000000", -- 1333 - 0x535  :    0 - 0x0
    "00000000", -- 1334 - 0x536  :    0 - 0x0
    "00000000", -- 1335 - 0x537  :    0 - 0x0
    "00000000", -- 1336 - 0x538  :    0 - 0x0
    "00000000", -- 1337 - 0x539  :    0 - 0x0
    "00000000", -- 1338 - 0x53a  :    0 - 0x0
    "00000000", -- 1339 - 0x53b  :    0 - 0x0
    "00000000", -- 1340 - 0x53c  :    0 - 0x0
    "00000000", -- 1341 - 0x53d  :    0 - 0x0
    "00000000", -- 1342 - 0x53e  :    0 - 0x0
    "00000000", -- 1343 - 0x53f  :    0 - 0x0
    "00000000", -- 1344 - 0x540  :    0 - 0x0 -- line 0xa
    "00000000", -- 1345 - 0x541  :    0 - 0x0
    "00000000", -- 1346 - 0x542  :    0 - 0x0
    "00000000", -- 1347 - 0x543  :    0 - 0x0
    "00000000", -- 1348 - 0x544  :    0 - 0x0
    "00000000", -- 1349 - 0x545  :    0 - 0x0
    "00000000", -- 1350 - 0x546  :    0 - 0x0
    "00000000", -- 1351 - 0x547  :    0 - 0x0
    "00000000", -- 1352 - 0x548  :    0 - 0x0
    "00000000", -- 1353 - 0x549  :    0 - 0x0
    "00000000", -- 1354 - 0x54a  :    0 - 0x0
    "00000000", -- 1355 - 0x54b  :    0 - 0x0
    "00000000", -- 1356 - 0x54c  :    0 - 0x0
    "00000000", -- 1357 - 0x54d  :    0 - 0x0
    "00000000", -- 1358 - 0x54e  :    0 - 0x0
    "00000000", -- 1359 - 0x54f  :    0 - 0x0
    "00000000", -- 1360 - 0x550  :    0 - 0x0
    "00000000", -- 1361 - 0x551  :    0 - 0x0
    "00000000", -- 1362 - 0x552  :    0 - 0x0
    "00000000", -- 1363 - 0x553  :    0 - 0x0
    "00000000", -- 1364 - 0x554  :    0 - 0x0
    "00000000", -- 1365 - 0x555  :    0 - 0x0
    "00000000", -- 1366 - 0x556  :    0 - 0x0
    "00000000", -- 1367 - 0x557  :    0 - 0x0
    "00000000", -- 1368 - 0x558  :    0 - 0x0
    "00000000", -- 1369 - 0x559  :    0 - 0x0
    "00000000", -- 1370 - 0x55a  :    0 - 0x0
    "00000000", -- 1371 - 0x55b  :    0 - 0x0
    "00000000", -- 1372 - 0x55c  :    0 - 0x0
    "00000000", -- 1373 - 0x55d  :    0 - 0x0
    "00000000", -- 1374 - 0x55e  :    0 - 0x0
    "00000000", -- 1375 - 0x55f  :    0 - 0x0
    "00000000", -- 1376 - 0x560  :    0 - 0x0 -- line 0xb
    "00000000", -- 1377 - 0x561  :    0 - 0x0
    "00000000", -- 1378 - 0x562  :    0 - 0x0
    "00000000", -- 1379 - 0x563  :    0 - 0x0
    "00000000", -- 1380 - 0x564  :    0 - 0x0
    "00000000", -- 1381 - 0x565  :    0 - 0x0
    "00000000", -- 1382 - 0x566  :    0 - 0x0
    "00000000", -- 1383 - 0x567  :    0 - 0x0
    "00000000", -- 1384 - 0x568  :    0 - 0x0
    "00000000", -- 1385 - 0x569  :    0 - 0x0
    "00000000", -- 1386 - 0x56a  :    0 - 0x0
    "00000000", -- 1387 - 0x56b  :    0 - 0x0
    "00000000", -- 1388 - 0x56c  :    0 - 0x0
    "00000000", -- 1389 - 0x56d  :    0 - 0x0
    "00000000", -- 1390 - 0x56e  :    0 - 0x0
    "00000000", -- 1391 - 0x56f  :    0 - 0x0
    "00000000", -- 1392 - 0x570  :    0 - 0x0
    "00000000", -- 1393 - 0x571  :    0 - 0x0
    "00000000", -- 1394 - 0x572  :    0 - 0x0
    "00000000", -- 1395 - 0x573  :    0 - 0x0
    "00000000", -- 1396 - 0x574  :    0 - 0x0
    "00000000", -- 1397 - 0x575  :    0 - 0x0
    "00000000", -- 1398 - 0x576  :    0 - 0x0
    "00000000", -- 1399 - 0x577  :    0 - 0x0
    "00000000", -- 1400 - 0x578  :    0 - 0x0
    "00000000", -- 1401 - 0x579  :    0 - 0x0
    "00000000", -- 1402 - 0x57a  :    0 - 0x0
    "00000000", -- 1403 - 0x57b  :    0 - 0x0
    "00000000", -- 1404 - 0x57c  :    0 - 0x0
    "00000000", -- 1405 - 0x57d  :    0 - 0x0
    "00000000", -- 1406 - 0x57e  :    0 - 0x0
    "00000000", -- 1407 - 0x57f  :    0 - 0x0
    "00000000", -- 1408 - 0x580  :    0 - 0x0 -- line 0xc
    "00000000", -- 1409 - 0x581  :    0 - 0x0
    "00000000", -- 1410 - 0x582  :    0 - 0x0
    "00000000", -- 1411 - 0x583  :    0 - 0x0
    "00000000", -- 1412 - 0x584  :    0 - 0x0
    "00000000", -- 1413 - 0x585  :    0 - 0x0
    "00000000", -- 1414 - 0x586  :    0 - 0x0
    "00000000", -- 1415 - 0x587  :    0 - 0x0
    "00000000", -- 1416 - 0x588  :    0 - 0x0
    "00000000", -- 1417 - 0x589  :    0 - 0x0
    "00000000", -- 1418 - 0x58a  :    0 - 0x0
    "00000000", -- 1419 - 0x58b  :    0 - 0x0
    "00000000", -- 1420 - 0x58c  :    0 - 0x0
    "00000000", -- 1421 - 0x58d  :    0 - 0x0
    "00000000", -- 1422 - 0x58e  :    0 - 0x0
    "00000000", -- 1423 - 0x58f  :    0 - 0x0
    "00000000", -- 1424 - 0x590  :    0 - 0x0
    "00000000", -- 1425 - 0x591  :    0 - 0x0
    "00000000", -- 1426 - 0x592  :    0 - 0x0
    "00000000", -- 1427 - 0x593  :    0 - 0x0
    "00000000", -- 1428 - 0x594  :    0 - 0x0
    "00000000", -- 1429 - 0x595  :    0 - 0x0
    "00000000", -- 1430 - 0x596  :    0 - 0x0
    "00000000", -- 1431 - 0x597  :    0 - 0x0
    "00000000", -- 1432 - 0x598  :    0 - 0x0
    "00000000", -- 1433 - 0x599  :    0 - 0x0
    "00000000", -- 1434 - 0x59a  :    0 - 0x0
    "00000000", -- 1435 - 0x59b  :    0 - 0x0
    "00000000", -- 1436 - 0x59c  :    0 - 0x0
    "00000000", -- 1437 - 0x59d  :    0 - 0x0
    "00000000", -- 1438 - 0x59e  :    0 - 0x0
    "00000000", -- 1439 - 0x59f  :    0 - 0x0
    "00000000", -- 1440 - 0x5a0  :    0 - 0x0 -- line 0xd
    "00000000", -- 1441 - 0x5a1  :    0 - 0x0
    "00000000", -- 1442 - 0x5a2  :    0 - 0x0
    "00000000", -- 1443 - 0x5a3  :    0 - 0x0
    "00000000", -- 1444 - 0x5a4  :    0 - 0x0
    "00000000", -- 1445 - 0x5a5  :    0 - 0x0
    "00000000", -- 1446 - 0x5a6  :    0 - 0x0
    "00000000", -- 1447 - 0x5a7  :    0 - 0x0
    "00000000", -- 1448 - 0x5a8  :    0 - 0x0
    "00000000", -- 1449 - 0x5a9  :    0 - 0x0
    "00000000", -- 1450 - 0x5aa  :    0 - 0x0
    "00000000", -- 1451 - 0x5ab  :    0 - 0x0
    "00000000", -- 1452 - 0x5ac  :    0 - 0x0
    "00000000", -- 1453 - 0x5ad  :    0 - 0x0
    "00000000", -- 1454 - 0x5ae  :    0 - 0x0
    "00000000", -- 1455 - 0x5af  :    0 - 0x0
    "00000000", -- 1456 - 0x5b0  :    0 - 0x0
    "00000000", -- 1457 - 0x5b1  :    0 - 0x0
    "00000000", -- 1458 - 0x5b2  :    0 - 0x0
    "00000000", -- 1459 - 0x5b3  :    0 - 0x0
    "00000000", -- 1460 - 0x5b4  :    0 - 0x0
    "00000000", -- 1461 - 0x5b5  :    0 - 0x0
    "00000000", -- 1462 - 0x5b6  :    0 - 0x0
    "00000000", -- 1463 - 0x5b7  :    0 - 0x0
    "00000000", -- 1464 - 0x5b8  :    0 - 0x0
    "00000000", -- 1465 - 0x5b9  :    0 - 0x0
    "00000000", -- 1466 - 0x5ba  :    0 - 0x0
    "00000000", -- 1467 - 0x5bb  :    0 - 0x0
    "00000000", -- 1468 - 0x5bc  :    0 - 0x0
    "00000000", -- 1469 - 0x5bd  :    0 - 0x0
    "00000000", -- 1470 - 0x5be  :    0 - 0x0
    "00000000", -- 1471 - 0x5bf  :    0 - 0x0
    "00000000", -- 1472 - 0x5c0  :    0 - 0x0 -- line 0xe
    "00000000", -- 1473 - 0x5c1  :    0 - 0x0
    "00000000", -- 1474 - 0x5c2  :    0 - 0x0
    "00000000", -- 1475 - 0x5c3  :    0 - 0x0
    "00000000", -- 1476 - 0x5c4  :    0 - 0x0
    "00000000", -- 1477 - 0x5c5  :    0 - 0x0
    "00000000", -- 1478 - 0x5c6  :    0 - 0x0
    "00000000", -- 1479 - 0x5c7  :    0 - 0x0
    "00000000", -- 1480 - 0x5c8  :    0 - 0x0
    "00000000", -- 1481 - 0x5c9  :    0 - 0x0
    "00000000", -- 1482 - 0x5ca  :    0 - 0x0
    "00000000", -- 1483 - 0x5cb  :    0 - 0x0
    "00000000", -- 1484 - 0x5cc  :    0 - 0x0
    "00000000", -- 1485 - 0x5cd  :    0 - 0x0
    "00000000", -- 1486 - 0x5ce  :    0 - 0x0
    "00000000", -- 1487 - 0x5cf  :    0 - 0x0
    "00000000", -- 1488 - 0x5d0  :    0 - 0x0
    "00000000", -- 1489 - 0x5d1  :    0 - 0x0
    "00000000", -- 1490 - 0x5d2  :    0 - 0x0
    "00000000", -- 1491 - 0x5d3  :    0 - 0x0
    "00000000", -- 1492 - 0x5d4  :    0 - 0x0
    "00000000", -- 1493 - 0x5d5  :    0 - 0x0
    "00000000", -- 1494 - 0x5d6  :    0 - 0x0
    "00000000", -- 1495 - 0x5d7  :    0 - 0x0
    "00000000", -- 1496 - 0x5d8  :    0 - 0x0
    "00000000", -- 1497 - 0x5d9  :    0 - 0x0
    "00000000", -- 1498 - 0x5da  :    0 - 0x0
    "00000000", -- 1499 - 0x5db  :    0 - 0x0
    "00000000", -- 1500 - 0x5dc  :    0 - 0x0
    "00000000", -- 1501 - 0x5dd  :    0 - 0x0
    "00000000", -- 1502 - 0x5de  :    0 - 0x0
    "00000000", -- 1503 - 0x5df  :    0 - 0x0
    "00000000", -- 1504 - 0x5e0  :    0 - 0x0 -- line 0xf
    "00000000", -- 1505 - 0x5e1  :    0 - 0x0
    "00000000", -- 1506 - 0x5e2  :    0 - 0x0
    "00000000", -- 1507 - 0x5e3  :    0 - 0x0
    "00000000", -- 1508 - 0x5e4  :    0 - 0x0
    "00000000", -- 1509 - 0x5e5  :    0 - 0x0
    "00000000", -- 1510 - 0x5e6  :    0 - 0x0
    "00000000", -- 1511 - 0x5e7  :    0 - 0x0
    "00000000", -- 1512 - 0x5e8  :    0 - 0x0
    "00000000", -- 1513 - 0x5e9  :    0 - 0x0
    "00000000", -- 1514 - 0x5ea  :    0 - 0x0
    "00000000", -- 1515 - 0x5eb  :    0 - 0x0
    "00000000", -- 1516 - 0x5ec  :    0 - 0x0
    "00000000", -- 1517 - 0x5ed  :    0 - 0x0
    "00000000", -- 1518 - 0x5ee  :    0 - 0x0
    "00000000", -- 1519 - 0x5ef  :    0 - 0x0
    "00000000", -- 1520 - 0x5f0  :    0 - 0x0
    "00000000", -- 1521 - 0x5f1  :    0 - 0x0
    "00000000", -- 1522 - 0x5f2  :    0 - 0x0
    "00000000", -- 1523 - 0x5f3  :    0 - 0x0
    "00000000", -- 1524 - 0x5f4  :    0 - 0x0
    "00000000", -- 1525 - 0x5f5  :    0 - 0x0
    "00000000", -- 1526 - 0x5f6  :    0 - 0x0
    "00000000", -- 1527 - 0x5f7  :    0 - 0x0
    "00000000", -- 1528 - 0x5f8  :    0 - 0x0
    "00000000", -- 1529 - 0x5f9  :    0 - 0x0
    "00000000", -- 1530 - 0x5fa  :    0 - 0x0
    "00000000", -- 1531 - 0x5fb  :    0 - 0x0
    "00000000", -- 1532 - 0x5fc  :    0 - 0x0
    "00000000", -- 1533 - 0x5fd  :    0 - 0x0
    "00000000", -- 1534 - 0x5fe  :    0 - 0x0
    "00000000", -- 1535 - 0x5ff  :    0 - 0x0
    "00000000", -- 1536 - 0x600  :    0 - 0x0 -- line 0x10
    "00000000", -- 1537 - 0x601  :    0 - 0x0
    "00000000", -- 1538 - 0x602  :    0 - 0x0
    "00000000", -- 1539 - 0x603  :    0 - 0x0
    "00000000", -- 1540 - 0x604  :    0 - 0x0
    "00000000", -- 1541 - 0x605  :    0 - 0x0
    "00000000", -- 1542 - 0x606  :    0 - 0x0
    "00000000", -- 1543 - 0x607  :    0 - 0x0
    "00000000", -- 1544 - 0x608  :    0 - 0x0
    "00000000", -- 1545 - 0x609  :    0 - 0x0
    "00000000", -- 1546 - 0x60a  :    0 - 0x0
    "00000000", -- 1547 - 0x60b  :    0 - 0x0
    "00000000", -- 1548 - 0x60c  :    0 - 0x0
    "00000000", -- 1549 - 0x60d  :    0 - 0x0
    "00000000", -- 1550 - 0x60e  :    0 - 0x0
    "00000000", -- 1551 - 0x60f  :    0 - 0x0
    "00000000", -- 1552 - 0x610  :    0 - 0x0
    "00000000", -- 1553 - 0x611  :    0 - 0x0
    "00000000", -- 1554 - 0x612  :    0 - 0x0
    "00000000", -- 1555 - 0x613  :    0 - 0x0
    "00000000", -- 1556 - 0x614  :    0 - 0x0
    "00000000", -- 1557 - 0x615  :    0 - 0x0
    "00000000", -- 1558 - 0x616  :    0 - 0x0
    "00000000", -- 1559 - 0x617  :    0 - 0x0
    "00000000", -- 1560 - 0x618  :    0 - 0x0
    "00000000", -- 1561 - 0x619  :    0 - 0x0
    "00000000", -- 1562 - 0x61a  :    0 - 0x0
    "00000000", -- 1563 - 0x61b  :    0 - 0x0
    "00000000", -- 1564 - 0x61c  :    0 - 0x0
    "00000000", -- 1565 - 0x61d  :    0 - 0x0
    "00000000", -- 1566 - 0x61e  :    0 - 0x0
    "00000000", -- 1567 - 0x61f  :    0 - 0x0
    "00000000", -- 1568 - 0x620  :    0 - 0x0 -- line 0x11
    "00000000", -- 1569 - 0x621  :    0 - 0x0
    "00000000", -- 1570 - 0x622  :    0 - 0x0
    "00000000", -- 1571 - 0x623  :    0 - 0x0
    "00000000", -- 1572 - 0x624  :    0 - 0x0
    "00000000", -- 1573 - 0x625  :    0 - 0x0
    "00000000", -- 1574 - 0x626  :    0 - 0x0
    "00000000", -- 1575 - 0x627  :    0 - 0x0
    "00000000", -- 1576 - 0x628  :    0 - 0x0
    "00000000", -- 1577 - 0x629  :    0 - 0x0
    "00000000", -- 1578 - 0x62a  :    0 - 0x0
    "00000000", -- 1579 - 0x62b  :    0 - 0x0
    "00000000", -- 1580 - 0x62c  :    0 - 0x0
    "00000000", -- 1581 - 0x62d  :    0 - 0x0
    "00000000", -- 1582 - 0x62e  :    0 - 0x0
    "00000000", -- 1583 - 0x62f  :    0 - 0x0
    "00000000", -- 1584 - 0x630  :    0 - 0x0
    "00000000", -- 1585 - 0x631  :    0 - 0x0
    "00000000", -- 1586 - 0x632  :    0 - 0x0
    "00000000", -- 1587 - 0x633  :    0 - 0x0
    "00000000", -- 1588 - 0x634  :    0 - 0x0
    "00000000", -- 1589 - 0x635  :    0 - 0x0
    "00000000", -- 1590 - 0x636  :    0 - 0x0
    "00000000", -- 1591 - 0x637  :    0 - 0x0
    "00000000", -- 1592 - 0x638  :    0 - 0x0
    "00000000", -- 1593 - 0x639  :    0 - 0x0
    "00000000", -- 1594 - 0x63a  :    0 - 0x0
    "00000000", -- 1595 - 0x63b  :    0 - 0x0
    "00000000", -- 1596 - 0x63c  :    0 - 0x0
    "00000000", -- 1597 - 0x63d  :    0 - 0x0
    "00000000", -- 1598 - 0x63e  :    0 - 0x0
    "00000000", -- 1599 - 0x63f  :    0 - 0x0
    "00000000", -- 1600 - 0x640  :    0 - 0x0 -- line 0x12
    "00000000", -- 1601 - 0x641  :    0 - 0x0
    "00000000", -- 1602 - 0x642  :    0 - 0x0
    "00000000", -- 1603 - 0x643  :    0 - 0x0
    "00000000", -- 1604 - 0x644  :    0 - 0x0
    "00000000", -- 1605 - 0x645  :    0 - 0x0
    "00000000", -- 1606 - 0x646  :    0 - 0x0
    "00000000", -- 1607 - 0x647  :    0 - 0x0
    "00000000", -- 1608 - 0x648  :    0 - 0x0
    "00000000", -- 1609 - 0x649  :    0 - 0x0
    "00000000", -- 1610 - 0x64a  :    0 - 0x0
    "00000000", -- 1611 - 0x64b  :    0 - 0x0
    "00000000", -- 1612 - 0x64c  :    0 - 0x0
    "00000000", -- 1613 - 0x64d  :    0 - 0x0
    "00000000", -- 1614 - 0x64e  :    0 - 0x0
    "00000000", -- 1615 - 0x64f  :    0 - 0x0
    "00000000", -- 1616 - 0x650  :    0 - 0x0
    "00000000", -- 1617 - 0x651  :    0 - 0x0
    "00000000", -- 1618 - 0x652  :    0 - 0x0
    "00000000", -- 1619 - 0x653  :    0 - 0x0
    "00000000", -- 1620 - 0x654  :    0 - 0x0
    "00000000", -- 1621 - 0x655  :    0 - 0x0
    "00000000", -- 1622 - 0x656  :    0 - 0x0
    "00000000", -- 1623 - 0x657  :    0 - 0x0
    "00000000", -- 1624 - 0x658  :    0 - 0x0
    "00000000", -- 1625 - 0x659  :    0 - 0x0
    "00000000", -- 1626 - 0x65a  :    0 - 0x0
    "00000000", -- 1627 - 0x65b  :    0 - 0x0
    "00000000", -- 1628 - 0x65c  :    0 - 0x0
    "00000000", -- 1629 - 0x65d  :    0 - 0x0
    "00000000", -- 1630 - 0x65e  :    0 - 0x0
    "00000000", -- 1631 - 0x65f  :    0 - 0x0
    "00000000", -- 1632 - 0x660  :    0 - 0x0 -- line 0x13
    "00000000", -- 1633 - 0x661  :    0 - 0x0
    "00000000", -- 1634 - 0x662  :    0 - 0x0
    "00000000", -- 1635 - 0x663  :    0 - 0x0
    "00000000", -- 1636 - 0x664  :    0 - 0x0
    "00000000", -- 1637 - 0x665  :    0 - 0x0
    "00000000", -- 1638 - 0x666  :    0 - 0x0
    "00000000", -- 1639 - 0x667  :    0 - 0x0
    "00000000", -- 1640 - 0x668  :    0 - 0x0
    "00000000", -- 1641 - 0x669  :    0 - 0x0
    "00000000", -- 1642 - 0x66a  :    0 - 0x0
    "00000000", -- 1643 - 0x66b  :    0 - 0x0
    "00000000", -- 1644 - 0x66c  :    0 - 0x0
    "00000000", -- 1645 - 0x66d  :    0 - 0x0
    "00000000", -- 1646 - 0x66e  :    0 - 0x0
    "00000000", -- 1647 - 0x66f  :    0 - 0x0
    "00000000", -- 1648 - 0x670  :    0 - 0x0
    "00000000", -- 1649 - 0x671  :    0 - 0x0
    "00000000", -- 1650 - 0x672  :    0 - 0x0
    "00000000", -- 1651 - 0x673  :    0 - 0x0
    "00000000", -- 1652 - 0x674  :    0 - 0x0
    "00000000", -- 1653 - 0x675  :    0 - 0x0
    "00000000", -- 1654 - 0x676  :    0 - 0x0
    "00000000", -- 1655 - 0x677  :    0 - 0x0
    "00000000", -- 1656 - 0x678  :    0 - 0x0
    "00000000", -- 1657 - 0x679  :    0 - 0x0
    "00000000", -- 1658 - 0x67a  :    0 - 0x0
    "00000000", -- 1659 - 0x67b  :    0 - 0x0
    "00000000", -- 1660 - 0x67c  :    0 - 0x0
    "00000000", -- 1661 - 0x67d  :    0 - 0x0
    "00000000", -- 1662 - 0x67e  :    0 - 0x0
    "00000000", -- 1663 - 0x67f  :    0 - 0x0
    "00000000", -- 1664 - 0x680  :    0 - 0x0 -- line 0x14
    "00000000", -- 1665 - 0x681  :    0 - 0x0
    "00000000", -- 1666 - 0x682  :    0 - 0x0
    "00000000", -- 1667 - 0x683  :    0 - 0x0
    "00000000", -- 1668 - 0x684  :    0 - 0x0
    "00000000", -- 1669 - 0x685  :    0 - 0x0
    "00000000", -- 1670 - 0x686  :    0 - 0x0
    "00000000", -- 1671 - 0x687  :    0 - 0x0
    "00000000", -- 1672 - 0x688  :    0 - 0x0
    "00000000", -- 1673 - 0x689  :    0 - 0x0
    "00000000", -- 1674 - 0x68a  :    0 - 0x0
    "00000000", -- 1675 - 0x68b  :    0 - 0x0
    "00000000", -- 1676 - 0x68c  :    0 - 0x0
    "00000000", -- 1677 - 0x68d  :    0 - 0x0
    "00000000", -- 1678 - 0x68e  :    0 - 0x0
    "00000000", -- 1679 - 0x68f  :    0 - 0x0
    "00000000", -- 1680 - 0x690  :    0 - 0x0
    "00000000", -- 1681 - 0x691  :    0 - 0x0
    "00000000", -- 1682 - 0x692  :    0 - 0x0
    "00000000", -- 1683 - 0x693  :    0 - 0x0
    "00000000", -- 1684 - 0x694  :    0 - 0x0
    "00000000", -- 1685 - 0x695  :    0 - 0x0
    "00000000", -- 1686 - 0x696  :    0 - 0x0
    "00000000", -- 1687 - 0x697  :    0 - 0x0
    "00000000", -- 1688 - 0x698  :    0 - 0x0
    "00000000", -- 1689 - 0x699  :    0 - 0x0
    "00000000", -- 1690 - 0x69a  :    0 - 0x0
    "00000000", -- 1691 - 0x69b  :    0 - 0x0
    "00000000", -- 1692 - 0x69c  :    0 - 0x0
    "00000000", -- 1693 - 0x69d  :    0 - 0x0
    "00000000", -- 1694 - 0x69e  :    0 - 0x0
    "00000000", -- 1695 - 0x69f  :    0 - 0x0
    "00000000", -- 1696 - 0x6a0  :    0 - 0x0 -- line 0x15
    "00000000", -- 1697 - 0x6a1  :    0 - 0x0
    "00000000", -- 1698 - 0x6a2  :    0 - 0x0
    "00000000", -- 1699 - 0x6a3  :    0 - 0x0
    "00000000", -- 1700 - 0x6a4  :    0 - 0x0
    "00000000", -- 1701 - 0x6a5  :    0 - 0x0
    "00000000", -- 1702 - 0x6a6  :    0 - 0x0
    "00000000", -- 1703 - 0x6a7  :    0 - 0x0
    "00000000", -- 1704 - 0x6a8  :    0 - 0x0
    "00000000", -- 1705 - 0x6a9  :    0 - 0x0
    "00000000", -- 1706 - 0x6aa  :    0 - 0x0
    "00000000", -- 1707 - 0x6ab  :    0 - 0x0
    "00000000", -- 1708 - 0x6ac  :    0 - 0x0
    "00000000", -- 1709 - 0x6ad  :    0 - 0x0
    "00000000", -- 1710 - 0x6ae  :    0 - 0x0
    "00000000", -- 1711 - 0x6af  :    0 - 0x0
    "00000000", -- 1712 - 0x6b0  :    0 - 0x0
    "00000000", -- 1713 - 0x6b1  :    0 - 0x0
    "00000000", -- 1714 - 0x6b2  :    0 - 0x0
    "00000000", -- 1715 - 0x6b3  :    0 - 0x0
    "00000000", -- 1716 - 0x6b4  :    0 - 0x0
    "00000000", -- 1717 - 0x6b5  :    0 - 0x0
    "00000000", -- 1718 - 0x6b6  :    0 - 0x0
    "00000000", -- 1719 - 0x6b7  :    0 - 0x0
    "00000000", -- 1720 - 0x6b8  :    0 - 0x0
    "00000000", -- 1721 - 0x6b9  :    0 - 0x0
    "00000000", -- 1722 - 0x6ba  :    0 - 0x0
    "00000000", -- 1723 - 0x6bb  :    0 - 0x0
    "00000000", -- 1724 - 0x6bc  :    0 - 0x0
    "00000000", -- 1725 - 0x6bd  :    0 - 0x0
    "00000000", -- 1726 - 0x6be  :    0 - 0x0
    "00000000", -- 1727 - 0x6bf  :    0 - 0x0
    "00000000", -- 1728 - 0x6c0  :    0 - 0x0 -- line 0x16
    "00000000", -- 1729 - 0x6c1  :    0 - 0x0
    "00000000", -- 1730 - 0x6c2  :    0 - 0x0
    "00000000", -- 1731 - 0x6c3  :    0 - 0x0
    "00000000", -- 1732 - 0x6c4  :    0 - 0x0
    "00000000", -- 1733 - 0x6c5  :    0 - 0x0
    "00000000", -- 1734 - 0x6c6  :    0 - 0x0
    "00000000", -- 1735 - 0x6c7  :    0 - 0x0
    "00000000", -- 1736 - 0x6c8  :    0 - 0x0
    "00000000", -- 1737 - 0x6c9  :    0 - 0x0
    "00000000", -- 1738 - 0x6ca  :    0 - 0x0
    "00000000", -- 1739 - 0x6cb  :    0 - 0x0
    "00000000", -- 1740 - 0x6cc  :    0 - 0x0
    "00000000", -- 1741 - 0x6cd  :    0 - 0x0
    "00000000", -- 1742 - 0x6ce  :    0 - 0x0
    "00000000", -- 1743 - 0x6cf  :    0 - 0x0
    "00000000", -- 1744 - 0x6d0  :    0 - 0x0
    "00000000", -- 1745 - 0x6d1  :    0 - 0x0
    "00000000", -- 1746 - 0x6d2  :    0 - 0x0
    "00000000", -- 1747 - 0x6d3  :    0 - 0x0
    "00000000", -- 1748 - 0x6d4  :    0 - 0x0
    "00000000", -- 1749 - 0x6d5  :    0 - 0x0
    "00000000", -- 1750 - 0x6d6  :    0 - 0x0
    "00000000", -- 1751 - 0x6d7  :    0 - 0x0
    "00000000", -- 1752 - 0x6d8  :    0 - 0x0
    "00000000", -- 1753 - 0x6d9  :    0 - 0x0
    "00000000", -- 1754 - 0x6da  :    0 - 0x0
    "00000000", -- 1755 - 0x6db  :    0 - 0x0
    "00000000", -- 1756 - 0x6dc  :    0 - 0x0
    "00000000", -- 1757 - 0x6dd  :    0 - 0x0
    "00000000", -- 1758 - 0x6de  :    0 - 0x0
    "00000000", -- 1759 - 0x6df  :    0 - 0x0
    "00000000", -- 1760 - 0x6e0  :    0 - 0x0 -- line 0x17
    "00000000", -- 1761 - 0x6e1  :    0 - 0x0
    "00000000", -- 1762 - 0x6e2  :    0 - 0x0
    "00000000", -- 1763 - 0x6e3  :    0 - 0x0
    "00000000", -- 1764 - 0x6e4  :    0 - 0x0
    "00000000", -- 1765 - 0x6e5  :    0 - 0x0
    "00000000", -- 1766 - 0x6e6  :    0 - 0x0
    "00000000", -- 1767 - 0x6e7  :    0 - 0x0
    "00000000", -- 1768 - 0x6e8  :    0 - 0x0
    "00000000", -- 1769 - 0x6e9  :    0 - 0x0
    "00000000", -- 1770 - 0x6ea  :    0 - 0x0
    "00000000", -- 1771 - 0x6eb  :    0 - 0x0
    "00000000", -- 1772 - 0x6ec  :    0 - 0x0
    "00000000", -- 1773 - 0x6ed  :    0 - 0x0
    "00000000", -- 1774 - 0x6ee  :    0 - 0x0
    "00000000", -- 1775 - 0x6ef  :    0 - 0x0
    "00000000", -- 1776 - 0x6f0  :    0 - 0x0
    "00000000", -- 1777 - 0x6f1  :    0 - 0x0
    "00000000", -- 1778 - 0x6f2  :    0 - 0x0
    "00000000", -- 1779 - 0x6f3  :    0 - 0x0
    "00000000", -- 1780 - 0x6f4  :    0 - 0x0
    "00000000", -- 1781 - 0x6f5  :    0 - 0x0
    "00000000", -- 1782 - 0x6f6  :    0 - 0x0
    "00000000", -- 1783 - 0x6f7  :    0 - 0x0
    "00000000", -- 1784 - 0x6f8  :    0 - 0x0
    "00000000", -- 1785 - 0x6f9  :    0 - 0x0
    "00000000", -- 1786 - 0x6fa  :    0 - 0x0
    "00000000", -- 1787 - 0x6fb  :    0 - 0x0
    "00000000", -- 1788 - 0x6fc  :    0 - 0x0
    "00000000", -- 1789 - 0x6fd  :    0 - 0x0
    "00000000", -- 1790 - 0x6fe  :    0 - 0x0
    "00000000", -- 1791 - 0x6ff  :    0 - 0x0
    "00000000", -- 1792 - 0x700  :    0 - 0x0 -- line 0x18
    "00000000", -- 1793 - 0x701  :    0 - 0x0
    "00000000", -- 1794 - 0x702  :    0 - 0x0
    "00000000", -- 1795 - 0x703  :    0 - 0x0
    "00000000", -- 1796 - 0x704  :    0 - 0x0
    "00000000", -- 1797 - 0x705  :    0 - 0x0
    "00000000", -- 1798 - 0x706  :    0 - 0x0
    "00000000", -- 1799 - 0x707  :    0 - 0x0
    "00000000", -- 1800 - 0x708  :    0 - 0x0
    "00000000", -- 1801 - 0x709  :    0 - 0x0
    "00000000", -- 1802 - 0x70a  :    0 - 0x0
    "00000000", -- 1803 - 0x70b  :    0 - 0x0
    "00000000", -- 1804 - 0x70c  :    0 - 0x0
    "00000000", -- 1805 - 0x70d  :    0 - 0x0
    "00000000", -- 1806 - 0x70e  :    0 - 0x0
    "00000000", -- 1807 - 0x70f  :    0 - 0x0
    "00000000", -- 1808 - 0x710  :    0 - 0x0
    "00000000", -- 1809 - 0x711  :    0 - 0x0
    "00000000", -- 1810 - 0x712  :    0 - 0x0
    "00000000", -- 1811 - 0x713  :    0 - 0x0
    "00000000", -- 1812 - 0x714  :    0 - 0x0
    "00000000", -- 1813 - 0x715  :    0 - 0x0
    "00000000", -- 1814 - 0x716  :    0 - 0x0
    "00000000", -- 1815 - 0x717  :    0 - 0x0
    "00000000", -- 1816 - 0x718  :    0 - 0x0
    "00000000", -- 1817 - 0x719  :    0 - 0x0
    "00000000", -- 1818 - 0x71a  :    0 - 0x0
    "00000000", -- 1819 - 0x71b  :    0 - 0x0
    "00000000", -- 1820 - 0x71c  :    0 - 0x0
    "00000000", -- 1821 - 0x71d  :    0 - 0x0
    "00000000", -- 1822 - 0x71e  :    0 - 0x0
    "00000000", -- 1823 - 0x71f  :    0 - 0x0
    "00000000", -- 1824 - 0x720  :    0 - 0x0 -- line 0x19
    "00000000", -- 1825 - 0x721  :    0 - 0x0
    "00000000", -- 1826 - 0x722  :    0 - 0x0
    "00000000", -- 1827 - 0x723  :    0 - 0x0
    "00000000", -- 1828 - 0x724  :    0 - 0x0
    "00000000", -- 1829 - 0x725  :    0 - 0x0
    "00000000", -- 1830 - 0x726  :    0 - 0x0
    "00000000", -- 1831 - 0x727  :    0 - 0x0
    "00000000", -- 1832 - 0x728  :    0 - 0x0
    "00000000", -- 1833 - 0x729  :    0 - 0x0
    "00000000", -- 1834 - 0x72a  :    0 - 0x0
    "00000000", -- 1835 - 0x72b  :    0 - 0x0
    "00000000", -- 1836 - 0x72c  :    0 - 0x0
    "00000000", -- 1837 - 0x72d  :    0 - 0x0
    "00000000", -- 1838 - 0x72e  :    0 - 0x0
    "00000000", -- 1839 - 0x72f  :    0 - 0x0
    "00000000", -- 1840 - 0x730  :    0 - 0x0
    "00000000", -- 1841 - 0x731  :    0 - 0x0
    "00000000", -- 1842 - 0x732  :    0 - 0x0
    "00000000", -- 1843 - 0x733  :    0 - 0x0
    "00000000", -- 1844 - 0x734  :    0 - 0x0
    "00000000", -- 1845 - 0x735  :    0 - 0x0
    "00000000", -- 1846 - 0x736  :    0 - 0x0
    "00000000", -- 1847 - 0x737  :    0 - 0x0
    "00000000", -- 1848 - 0x738  :    0 - 0x0
    "00000000", -- 1849 - 0x739  :    0 - 0x0
    "00000000", -- 1850 - 0x73a  :    0 - 0x0
    "00000000", -- 1851 - 0x73b  :    0 - 0x0
    "00000000", -- 1852 - 0x73c  :    0 - 0x0
    "00000000", -- 1853 - 0x73d  :    0 - 0x0
    "00000000", -- 1854 - 0x73e  :    0 - 0x0
    "00000000", -- 1855 - 0x73f  :    0 - 0x0
    "00000000", -- 1856 - 0x740  :    0 - 0x0 -- line 0x1a
    "00000000", -- 1857 - 0x741  :    0 - 0x0
    "00000000", -- 1858 - 0x742  :    0 - 0x0
    "00000000", -- 1859 - 0x743  :    0 - 0x0
    "00000000", -- 1860 - 0x744  :    0 - 0x0
    "00000000", -- 1861 - 0x745  :    0 - 0x0
    "00000000", -- 1862 - 0x746  :    0 - 0x0
    "00000000", -- 1863 - 0x747  :    0 - 0x0
    "00000000", -- 1864 - 0x748  :    0 - 0x0
    "00000000", -- 1865 - 0x749  :    0 - 0x0
    "00000000", -- 1866 - 0x74a  :    0 - 0x0
    "00000000", -- 1867 - 0x74b  :    0 - 0x0
    "00000000", -- 1868 - 0x74c  :    0 - 0x0
    "00000000", -- 1869 - 0x74d  :    0 - 0x0
    "00000000", -- 1870 - 0x74e  :    0 - 0x0
    "00000000", -- 1871 - 0x74f  :    0 - 0x0
    "00000000", -- 1872 - 0x750  :    0 - 0x0
    "00000000", -- 1873 - 0x751  :    0 - 0x0
    "00000000", -- 1874 - 0x752  :    0 - 0x0
    "00000000", -- 1875 - 0x753  :    0 - 0x0
    "00000000", -- 1876 - 0x754  :    0 - 0x0
    "00000000", -- 1877 - 0x755  :    0 - 0x0
    "00000000", -- 1878 - 0x756  :    0 - 0x0
    "00000000", -- 1879 - 0x757  :    0 - 0x0
    "00000000", -- 1880 - 0x758  :    0 - 0x0
    "00000000", -- 1881 - 0x759  :    0 - 0x0
    "00000000", -- 1882 - 0x75a  :    0 - 0x0
    "00000000", -- 1883 - 0x75b  :    0 - 0x0
    "00000000", -- 1884 - 0x75c  :    0 - 0x0
    "00000000", -- 1885 - 0x75d  :    0 - 0x0
    "00000000", -- 1886 - 0x75e  :    0 - 0x0
    "00000000", -- 1887 - 0x75f  :    0 - 0x0
    "00000000", -- 1888 - 0x760  :    0 - 0x0 -- line 0x1b
    "00000000", -- 1889 - 0x761  :    0 - 0x0
    "00000000", -- 1890 - 0x762  :    0 - 0x0
    "00000000", -- 1891 - 0x763  :    0 - 0x0
    "00000000", -- 1892 - 0x764  :    0 - 0x0
    "00000000", -- 1893 - 0x765  :    0 - 0x0
    "00000000", -- 1894 - 0x766  :    0 - 0x0
    "00000000", -- 1895 - 0x767  :    0 - 0x0
    "00000000", -- 1896 - 0x768  :    0 - 0x0
    "00000000", -- 1897 - 0x769  :    0 - 0x0
    "00000000", -- 1898 - 0x76a  :    0 - 0x0
    "00000000", -- 1899 - 0x76b  :    0 - 0x0
    "00000000", -- 1900 - 0x76c  :    0 - 0x0
    "00000000", -- 1901 - 0x76d  :    0 - 0x0
    "00000000", -- 1902 - 0x76e  :    0 - 0x0
    "00000000", -- 1903 - 0x76f  :    0 - 0x0
    "00000000", -- 1904 - 0x770  :    0 - 0x0
    "00000000", -- 1905 - 0x771  :    0 - 0x0
    "00000000", -- 1906 - 0x772  :    0 - 0x0
    "00000000", -- 1907 - 0x773  :    0 - 0x0
    "00000000", -- 1908 - 0x774  :    0 - 0x0
    "00000000", -- 1909 - 0x775  :    0 - 0x0
    "00000000", -- 1910 - 0x776  :    0 - 0x0
    "00000000", -- 1911 - 0x777  :    0 - 0x0
    "00000000", -- 1912 - 0x778  :    0 - 0x0
    "00000000", -- 1913 - 0x779  :    0 - 0x0
    "00000000", -- 1914 - 0x77a  :    0 - 0x0
    "00000000", -- 1915 - 0x77b  :    0 - 0x0
    "00000000", -- 1916 - 0x77c  :    0 - 0x0
    "00000000", -- 1917 - 0x77d  :    0 - 0x0
    "00000000", -- 1918 - 0x77e  :    0 - 0x0
    "00000000", -- 1919 - 0x77f  :    0 - 0x0
    "10100101", -- 1920 - 0x780  :  165 - 0xa5 -- line 0x1c
    "10100101", -- 1921 - 0x781  :  165 - 0xa5
    "10100101", -- 1922 - 0x782  :  165 - 0xa5
    "10100101", -- 1923 - 0x783  :  165 - 0xa5
    "10100101", -- 1924 - 0x784  :  165 - 0xa5
    "10100101", -- 1925 - 0x785  :  165 - 0xa5
    "10100101", -- 1926 - 0x786  :  165 - 0xa5
    "10100101", -- 1927 - 0x787  :  165 - 0xa5
    "10100101", -- 1928 - 0x788  :  165 - 0xa5
    "10100101", -- 1929 - 0x789  :  165 - 0xa5
    "10100101", -- 1930 - 0x78a  :  165 - 0xa5
    "10100101", -- 1931 - 0x78b  :  165 - 0xa5
    "10100101", -- 1932 - 0x78c  :  165 - 0xa5
    "10100101", -- 1933 - 0x78d  :  165 - 0xa5
    "10100101", -- 1934 - 0x78e  :  165 - 0xa5
    "10100101", -- 1935 - 0x78f  :  165 - 0xa5
    "10100101", -- 1936 - 0x790  :  165 - 0xa5
    "10100101", -- 1937 - 0x791  :  165 - 0xa5
    "10100101", -- 1938 - 0x792  :  165 - 0xa5
    "10100101", -- 1939 - 0x793  :  165 - 0xa5
    "10100101", -- 1940 - 0x794  :  165 - 0xa5
    "10100101", -- 1941 - 0x795  :  165 - 0xa5
    "10100101", -- 1942 - 0x796  :  165 - 0xa5
    "10100101", -- 1943 - 0x797  :  165 - 0xa5
    "10100101", -- 1944 - 0x798  :  165 - 0xa5
    "10100101", -- 1945 - 0x799  :  165 - 0xa5
    "10100101", -- 1946 - 0x79a  :  165 - 0xa5
    "10100101", -- 1947 - 0x79b  :  165 - 0xa5
    "10100101", -- 1948 - 0x79c  :  165 - 0xa5
    "10100101", -- 1949 - 0x79d  :  165 - 0xa5
    "10100101", -- 1950 - 0x79e  :  165 - 0xa5
    "10100101", -- 1951 - 0x79f  :  165 - 0xa5
    "10100000", -- 1952 - 0x7a0  :  160 - 0xa0 -- line 0x1d
    "10100000", -- 1953 - 0x7a1  :  160 - 0xa0
    "10100000", -- 1954 - 0x7a2  :  160 - 0xa0
    "10100000", -- 1955 - 0x7a3  :  160 - 0xa0
    "10100000", -- 1956 - 0x7a4  :  160 - 0xa0
    "10100000", -- 1957 - 0x7a5  :  160 - 0xa0
    "10100000", -- 1958 - 0x7a6  :  160 - 0xa0
    "10100000", -- 1959 - 0x7a7  :  160 - 0xa0
    "10100000", -- 1960 - 0x7a8  :  160 - 0xa0
    "10100000", -- 1961 - 0x7a9  :  160 - 0xa0
    "10100000", -- 1962 - 0x7aa  :  160 - 0xa0
    "10100000", -- 1963 - 0x7ab  :  160 - 0xa0
    "10100000", -- 1964 - 0x7ac  :  160 - 0xa0
    "10100000", -- 1965 - 0x7ad  :  160 - 0xa0
    "10100000", -- 1966 - 0x7ae  :  160 - 0xa0
    "10100000", -- 1967 - 0x7af  :  160 - 0xa0
    "10100000", -- 1968 - 0x7b0  :  160 - 0xa0
    "10100000", -- 1969 - 0x7b1  :  160 - 0xa0
    "10100000", -- 1970 - 0x7b2  :  160 - 0xa0
    "10100000", -- 1971 - 0x7b3  :  160 - 0xa0
    "10100000", -- 1972 - 0x7b4  :  160 - 0xa0
    "10100000", -- 1973 - 0x7b5  :  160 - 0xa0
    "10100000", -- 1974 - 0x7b6  :  160 - 0xa0
    "10100000", -- 1975 - 0x7b7  :  160 - 0xa0
    "10100000", -- 1976 - 0x7b8  :  160 - 0xa0
    "10100000", -- 1977 - 0x7b9  :  160 - 0xa0
    "10100000", -- 1978 - 0x7ba  :  160 - 0xa0
    "10100000", -- 1979 - 0x7bb  :  160 - 0xa0
    "10100000", -- 1980 - 0x7bc  :  160 - 0xa0
    "10100000", -- 1981 - 0x7bd  :  160 - 0xa0
    "10100000", -- 1982 - 0x7be  :  160 - 0xa0
    "10100000", -- 1983 - 0x7bf  :  160 - 0xa0
        ---- Attribute Table 1----
    "00000000", -- 1984 - 0x7c0  :    0 - 0x0
    "00000000", -- 1985 - 0x7c1  :    0 - 0x0
    "00000000", -- 1986 - 0x7c2  :    0 - 0x0
    "00000000", -- 1987 - 0x7c3  :    0 - 0x0
    "00000000", -- 1988 - 0x7c4  :    0 - 0x0
    "00000000", -- 1989 - 0x7c5  :    0 - 0x0
    "00000000", -- 1990 - 0x7c6  :    0 - 0x0
    "00000000", -- 1991 - 0x7c7  :    0 - 0x0
    "00000000", -- 1992 - 0x7c8  :    0 - 0x0
    "00000000", -- 1993 - 0x7c9  :    0 - 0x0
    "00000000", -- 1994 - 0x7ca  :    0 - 0x0
    "00000000", -- 1995 - 0x7cb  :    0 - 0x0
    "00000000", -- 1996 - 0x7cc  :    0 - 0x0
    "00000000", -- 1997 - 0x7cd  :    0 - 0x0
    "00000000", -- 1998 - 0x7ce  :    0 - 0x0
    "00000000", -- 1999 - 0x7cf  :    0 - 0x0
    "00000000", -- 2000 - 0x7d0  :    0 - 0x0
    "00000000", -- 2001 - 0x7d1  :    0 - 0x0
    "00000000", -- 2002 - 0x7d2  :    0 - 0x0
    "00000000", -- 2003 - 0x7d3  :    0 - 0x0
    "00000000", -- 2004 - 0x7d4  :    0 - 0x0
    "00000000", -- 2005 - 0x7d5  :    0 - 0x0
    "00000000", -- 2006 - 0x7d6  :    0 - 0x0
    "00000000", -- 2007 - 0x7d7  :    0 - 0x0
    "00000000", -- 2008 - 0x7d8  :    0 - 0x0
    "00000000", -- 2009 - 0x7d9  :    0 - 0x0
    "00000000", -- 2010 - 0x7da  :    0 - 0x0
    "00000000", -- 2011 - 0x7db  :    0 - 0x0
    "00000000", -- 2012 - 0x7dc  :    0 - 0x0
    "00000000", -- 2013 - 0x7dd  :    0 - 0x0
    "00000000", -- 2014 - 0x7de  :    0 - 0x0
    "00000000", -- 2015 - 0x7df  :    0 - 0x0
    "00000000", -- 2016 - 0x7e0  :    0 - 0x0
    "00000000", -- 2017 - 0x7e1  :    0 - 0x0
    "00000000", -- 2018 - 0x7e2  :    0 - 0x0
    "00000000", -- 2019 - 0x7e3  :    0 - 0x0
    "00000000", -- 2020 - 0x7e4  :    0 - 0x0
    "00000000", -- 2021 - 0x7e5  :    0 - 0x0
    "00000000", -- 2022 - 0x7e6  :    0 - 0x0
    "00000000", -- 2023 - 0x7e7  :    0 - 0x0
    "00000000", -- 2024 - 0x7e8  :    0 - 0x0
    "00000000", -- 2025 - 0x7e9  :    0 - 0x0
    "00000000", -- 2026 - 0x7ea  :    0 - 0x0
    "00000000", -- 2027 - 0x7eb  :    0 - 0x0
    "00000000", -- 2028 - 0x7ec  :    0 - 0x0
    "00000000", -- 2029 - 0x7ed  :    0 - 0x0
    "00000000", -- 2030 - 0x7ee  :    0 - 0x0
    "00000000", -- 2031 - 0x7ef  :    0 - 0x0
    "00000000", -- 2032 - 0x7f0  :    0 - 0x0
    "00000000", -- 2033 - 0x7f1  :    0 - 0x0
    "00000000", -- 2034 - 0x7f2  :    0 - 0x0
    "00000000", -- 2035 - 0x7f3  :    0 - 0x0
    "00000000", -- 2036 - 0x7f4  :    0 - 0x0
    "00000000", -- 2037 - 0x7f5  :    0 - 0x0
    "00000000", -- 2038 - 0x7f6  :    0 - 0x0
    "00000000", -- 2039 - 0x7f7  :    0 - 0x0
    "00000000", -- 2040 - 0x7f8  :    0 - 0x0
    "00000000", -- 2041 - 0x7f9  :    0 - 0x0
    "00000000", -- 2042 - 0x7fa  :    0 - 0x0
    "00000000", -- 2043 - 0x7fb  :    0 - 0x0
    "00000000", -- 2044 - 0x7fc  :    0 - 0x0
    "00000000", -- 2045 - 0x7fd  :    0 - 0x0
    "00000000", -- 2046 - 0x7fe  :    0 - 0x0
    "00000000"  -- 2047 - 0x7ff  :    0 - 0x0
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
