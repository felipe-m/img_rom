//- Autcmatically generated verilog ROM from a NES memory file----
//-   PATTERN TABLE WITH ONLY ONE COLOR PLANE
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


//-  Original memory dump file name: nova_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_PTABLE_NOVA_color0
  (
     input     clk,   // clock
     input      [12-1:0] addr,  //4096 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                              //  address:   value 
                              //    dec  : dec - hex
          // Sprite pattern Table
      12'h0: dout <= 8'b11111111; //    0 : 255 - 0xff -- Sprite 0x0
      12'h1: dout <= 8'b11111111; //    1 : 255 - 0xff
      12'h2: dout <= 8'b11000000; //    2 : 192 - 0xc0
      12'h3: dout <= 8'b11000000; //    3 : 192 - 0xc0
      12'h4: dout <= 8'b11000000; //    4 : 192 - 0xc0
      12'h5: dout <= 8'b11000000; //    5 : 192 - 0xc0
      12'h6: dout <= 8'b11010101; //    6 : 213 - 0xd5
      12'h7: dout <= 8'b11111111; //    7 : 255 - 0xff
      12'h8: dout <= 8'b11111111; //    8 : 255 - 0xff -- Sprite 0x1
      12'h9: dout <= 8'b11111111; //    9 : 255 - 0xff
      12'hA: dout <= 8'b11001110; //   10 : 206 - 0xce
      12'hB: dout <= 8'b11000110; //   11 : 198 - 0xc6
      12'hC: dout <= 8'b11001110; //   12 : 206 - 0xce
      12'hD: dout <= 8'b11000110; //   13 : 198 - 0xc6
      12'hE: dout <= 8'b11101110; //   14 : 238 - 0xee
      12'hF: dout <= 8'b11111111; //   15 : 255 - 0xff
      12'h10: dout <= 8'b11111111; //   16 : 255 - 0xff -- Sprite 0x2
      12'h11: dout <= 8'b11111111; //   17 : 255 - 0xff
      12'h12: dout <= 8'b01110001; //   18 : 113 - 0x71
      12'h13: dout <= 8'b00110011; //   19 :  51 - 0x33
      12'h14: dout <= 8'b01110001; //   20 : 113 - 0x71
      12'h15: dout <= 8'b00110011; //   21 :  51 - 0x33
      12'h16: dout <= 8'b01110101; //   22 : 117 - 0x75
      12'h17: dout <= 8'b11111111; //   23 : 255 - 0xff
      12'h18: dout <= 8'b11111111; //   24 : 255 - 0xff -- Sprite 0x3
      12'h19: dout <= 8'b11111111; //   25 : 255 - 0xff
      12'h1A: dout <= 8'b00000011; //   26 :   3 - 0x3
      12'h1B: dout <= 8'b00000001; //   27 :   1 - 0x1
      12'h1C: dout <= 8'b00000011; //   28 :   3 - 0x3
      12'h1D: dout <= 8'b00000001; //   29 :   1 - 0x1
      12'h1E: dout <= 8'b10101011; //   30 : 171 - 0xab
      12'h1F: dout <= 8'b11111111; //   31 : 255 - 0xff
      12'h20: dout <= 8'b11111111; //   32 : 255 - 0xff -- Sprite 0x4
      12'h21: dout <= 8'b11111111; //   33 : 255 - 0xff
      12'h22: dout <= 8'b11100000; //   34 : 224 - 0xe0
      12'h23: dout <= 8'b11000110; //   35 : 198 - 0xc6
      12'h24: dout <= 8'b11000110; //   36 : 198 - 0xc6
      12'h25: dout <= 8'b11110110; //   37 : 246 - 0xf6
      12'h26: dout <= 8'b11110000; //   38 : 240 - 0xf0
      12'h27: dout <= 8'b11110001; //   39 : 241 - 0xf1
      12'h28: dout <= 8'b11000111; //   40 : 199 - 0xc7 -- Sprite 0x5
      12'h29: dout <= 8'b11001111; //   41 : 207 - 0xcf
      12'h2A: dout <= 8'b11011111; //   42 : 223 - 0xdf
      12'h2B: dout <= 8'b11011111; //   43 : 223 - 0xdf
      12'h2C: dout <= 8'b11001110; //   44 : 206 - 0xce
      12'h2D: dout <= 8'b11100000; //   45 : 224 - 0xe0
      12'h2E: dout <= 8'b11111111; //   46 : 255 - 0xff
      12'h2F: dout <= 8'b11111111; //   47 : 255 - 0xff
      12'h30: dout <= 8'b11111111; //   48 : 255 - 0xff -- Sprite 0x6
      12'h31: dout <= 8'b11111111; //   49 : 255 - 0xff
      12'h32: dout <= 8'b00000111; //   50 :   7 - 0x7
      12'h33: dout <= 8'b01100011; //   51 :  99 - 0x63
      12'h34: dout <= 8'b01100011; //   52 :  99 - 0x63
      12'h35: dout <= 8'b01101111; //   53 : 111 - 0x6f
      12'h36: dout <= 8'b00001111; //   54 :  15 - 0xf
      12'h37: dout <= 8'b10001111; //   55 : 143 - 0x8f
      12'h38: dout <= 8'b11100011; //   56 : 227 - 0xe3 -- Sprite 0x7
      12'h39: dout <= 8'b11110011; //   57 : 243 - 0xf3
      12'h3A: dout <= 8'b11111011; //   58 : 251 - 0xfb
      12'h3B: dout <= 8'b11111011; //   59 : 251 - 0xfb
      12'h3C: dout <= 8'b01110011; //   60 : 115 - 0x73
      12'h3D: dout <= 8'b00000111; //   61 :   7 - 0x7
      12'h3E: dout <= 8'b11111111; //   62 : 255 - 0xff
      12'h3F: dout <= 8'b11111111; //   63 : 255 - 0xff
      12'h40: dout <= 8'b11111111; //   64 : 255 - 0xff -- Sprite 0x8
      12'h41: dout <= 8'b11010101; //   65 : 213 - 0xd5
      12'h42: dout <= 8'b10101010; //   66 : 170 - 0xaa
      12'h43: dout <= 8'b11010101; //   67 : 213 - 0xd5
      12'h44: dout <= 8'b10101010; //   68 : 170 - 0xaa
      12'h45: dout <= 8'b11010101; //   69 : 213 - 0xd5
      12'h46: dout <= 8'b10101010; //   70 : 170 - 0xaa
      12'h47: dout <= 8'b11010101; //   71 : 213 - 0xd5
      12'h48: dout <= 8'b10101010; //   72 : 170 - 0xaa -- Sprite 0x9
      12'h49: dout <= 8'b11010101; //   73 : 213 - 0xd5
      12'h4A: dout <= 8'b10101010; //   74 : 170 - 0xaa
      12'h4B: dout <= 8'b11010101; //   75 : 213 - 0xd5
      12'h4C: dout <= 8'b10101010; //   76 : 170 - 0xaa
      12'h4D: dout <= 8'b11110101; //   77 : 245 - 0xf5
      12'h4E: dout <= 8'b10101010; //   78 : 170 - 0xaa
      12'h4F: dout <= 8'b11111111; //   79 : 255 - 0xff
      12'h50: dout <= 8'b11111111; //   80 : 255 - 0xff -- Sprite 0xa
      12'h51: dout <= 8'b01010101; //   81 :  85 - 0x55
      12'h52: dout <= 8'b10101111; //   82 : 175 - 0xaf
      12'h53: dout <= 8'b01010101; //   83 :  85 - 0x55
      12'h54: dout <= 8'b10101011; //   84 : 171 - 0xab
      12'h55: dout <= 8'b01010101; //   85 :  85 - 0x55
      12'h56: dout <= 8'b10101011; //   86 : 171 - 0xab
      12'h57: dout <= 8'b01010101; //   87 :  85 - 0x55
      12'h58: dout <= 8'b10101011; //   88 : 171 - 0xab -- Sprite 0xb
      12'h59: dout <= 8'b01010101; //   89 :  85 - 0x55
      12'h5A: dout <= 8'b10101011; //   90 : 171 - 0xab
      12'h5B: dout <= 8'b01010101; //   91 :  85 - 0x55
      12'h5C: dout <= 8'b10101011; //   92 : 171 - 0xab
      12'h5D: dout <= 8'b01010101; //   93 :  85 - 0x55
      12'h5E: dout <= 8'b10101011; //   94 : 171 - 0xab
      12'h5F: dout <= 8'b11111111; //   95 : 255 - 0xff
      12'h60: dout <= 8'b11111111; //   96 : 255 - 0xff -- Sprite 0xc
      12'h61: dout <= 8'b11010101; //   97 : 213 - 0xd5
      12'h62: dout <= 8'b10100000; //   98 : 160 - 0xa0
      12'h63: dout <= 8'b11010000; //   99 : 208 - 0xd0
      12'h64: dout <= 8'b10001111; //  100 : 143 - 0x8f
      12'h65: dout <= 8'b11001000; //  101 : 200 - 0xc8
      12'h66: dout <= 8'b10001000; //  102 : 136 - 0x88
      12'h67: dout <= 8'b11001000; //  103 : 200 - 0xc8
      12'h68: dout <= 8'b10001000; //  104 : 136 - 0x88 -- Sprite 0xd
      12'h69: dout <= 8'b11001000; //  105 : 200 - 0xc8
      12'h6A: dout <= 8'b10001000; //  106 : 136 - 0x88
      12'h6B: dout <= 8'b11001111; //  107 : 207 - 0xcf
      12'h6C: dout <= 8'b10010000; //  108 : 144 - 0x90
      12'h6D: dout <= 8'b11100000; //  109 : 224 - 0xe0
      12'h6E: dout <= 8'b11101010; //  110 : 234 - 0xea
      12'h6F: dout <= 8'b11111111; //  111 : 255 - 0xff
      12'h70: dout <= 8'b11111111; //  112 : 255 - 0xff -- Sprite 0xe
      12'h71: dout <= 8'b01011011; //  113 :  91 - 0x5b
      12'h72: dout <= 8'b00000111; //  114 :   7 - 0x7
      12'h73: dout <= 8'b00001001; //  115 :   9 - 0x9
      12'h74: dout <= 8'b11110011; //  116 : 243 - 0xf3
      12'h75: dout <= 8'b00010001; //  117 :  17 - 0x11
      12'h76: dout <= 8'b00010011; //  118 :  19 - 0x13
      12'h77: dout <= 8'b00010001; //  119 :  17 - 0x11
      12'h78: dout <= 8'b00010011; //  120 :  19 - 0x13 -- Sprite 0xf
      12'h79: dout <= 8'b00010001; //  121 :  17 - 0x11
      12'h7A: dout <= 8'b00010011; //  122 :  19 - 0x13
      12'h7B: dout <= 8'b11110001; //  123 : 241 - 0xf1
      12'h7C: dout <= 8'b00001011; //  124 :  11 - 0xb
      12'h7D: dout <= 8'b00000101; //  125 :   5 - 0x5
      12'h7E: dout <= 8'b10101011; //  126 : 171 - 0xab
      12'h7F: dout <= 8'b11111111; //  127 : 255 - 0xff
      12'h80: dout <= 8'b11010000; //  128 : 208 - 0xd0 -- Sprite 0x10
      12'h81: dout <= 8'b10010000; //  129 : 144 - 0x90
      12'h82: dout <= 8'b11011111; //  130 : 223 - 0xdf
      12'h83: dout <= 8'b10011010; //  131 : 154 - 0x9a
      12'h84: dout <= 8'b11010101; //  132 : 213 - 0xd5
      12'h85: dout <= 8'b10011111; //  133 : 159 - 0x9f
      12'h86: dout <= 8'b11010000; //  134 : 208 - 0xd0
      12'h87: dout <= 8'b10010000; //  135 : 144 - 0x90
      12'h88: dout <= 8'b00001001; //  136 :   9 - 0x9 -- Sprite 0x11
      12'h89: dout <= 8'b00001011; //  137 :  11 - 0xb
      12'h8A: dout <= 8'b11111001; //  138 : 249 - 0xf9
      12'h8B: dout <= 8'b10101011; //  139 : 171 - 0xab
      12'h8C: dout <= 8'b01011001; //  140 :  89 - 0x59
      12'h8D: dout <= 8'b11111011; //  141 : 251 - 0xfb
      12'h8E: dout <= 8'b00001001; //  142 :   9 - 0x9
      12'h8F: dout <= 8'b00001011; //  143 :  11 - 0xb
      12'h90: dout <= 8'b00011000; //  144 :  24 - 0x18 -- Sprite 0x12
      12'h91: dout <= 8'b00010100; //  145 :  20 - 0x14
      12'h92: dout <= 8'b00010100; //  146 :  20 - 0x14
      12'h93: dout <= 8'b00111010; //  147 :  58 - 0x3a
      12'h94: dout <= 8'b00111010; //  148 :  58 - 0x3a
      12'h95: dout <= 8'b01111010; //  149 : 122 - 0x7a
      12'h96: dout <= 8'b01111010; //  150 : 122 - 0x7a
      12'h97: dout <= 8'b01111010; //  151 : 122 - 0x7a
      12'h98: dout <= 8'b11111011; //  152 : 251 - 0xfb -- Sprite 0x13
      12'h99: dout <= 8'b11111101; //  153 : 253 - 0xfd
      12'h9A: dout <= 8'b11111101; //  154 : 253 - 0xfd
      12'h9B: dout <= 8'b11111101; //  155 : 253 - 0xfd
      12'h9C: dout <= 8'b11111101; //  156 : 253 - 0xfd
      12'h9D: dout <= 8'b11111101; //  157 : 253 - 0xfd
      12'h9E: dout <= 8'b10000001; //  158 : 129 - 0x81
      12'h9F: dout <= 8'b11111111; //  159 : 255 - 0xff
      12'hA0: dout <= 8'b00000000; //  160 :   0 - 0x0 -- Sprite 0x14
      12'hA1: dout <= 8'b00000111; //  161 :   7 - 0x7
      12'hA2: dout <= 8'b00000010; //  162 :   2 - 0x2
      12'hA3: dout <= 8'b00000100; //  163 :   4 - 0x4
      12'hA4: dout <= 8'b00000011; //  164 :   3 - 0x3
      12'hA5: dout <= 8'b00000011; //  165 :   3 - 0x3
      12'hA6: dout <= 8'b00001101; //  166 :  13 - 0xd
      12'hA7: dout <= 8'b00010111; //  167 :  23 - 0x17
      12'hA8: dout <= 8'b00101111; //  168 :  47 - 0x2f -- Sprite 0x15
      12'hA9: dout <= 8'b01001111; //  169 :  79 - 0x4f
      12'hAA: dout <= 8'b01001111; //  170 :  79 - 0x4f
      12'hAB: dout <= 8'b01001111; //  171 :  79 - 0x4f
      12'hAC: dout <= 8'b01001111; //  172 :  79 - 0x4f
      12'hAD: dout <= 8'b00100111; //  173 :  39 - 0x27
      12'hAE: dout <= 8'b00010000; //  174 :  16 - 0x10
      12'hAF: dout <= 8'b00001111; //  175 :  15 - 0xf
      12'hB0: dout <= 8'b00000000; //  176 :   0 - 0x0 -- Sprite 0x16
      12'hB1: dout <= 8'b11100000; //  177 : 224 - 0xe0
      12'hB2: dout <= 8'b10100000; //  178 : 160 - 0xa0
      12'hB3: dout <= 8'b00100000; //  179 :  32 - 0x20
      12'hB4: dout <= 8'b11000000; //  180 : 192 - 0xc0
      12'hB5: dout <= 8'b01000000; //  181 :  64 - 0x40
      12'hB6: dout <= 8'b00110000; //  182 :  48 - 0x30
      12'hB7: dout <= 8'b11101000; //  183 : 232 - 0xe8
      12'hB8: dout <= 8'b11110100; //  184 : 244 - 0xf4 -- Sprite 0x17
      12'hB9: dout <= 8'b11110010; //  185 : 242 - 0xf2
      12'hBA: dout <= 8'b11110010; //  186 : 242 - 0xf2
      12'hBB: dout <= 8'b11110010; //  187 : 242 - 0xf2
      12'hBC: dout <= 8'b11110010; //  188 : 242 - 0xf2
      12'hBD: dout <= 8'b11100100; //  189 : 228 - 0xe4
      12'hBE: dout <= 8'b00001000; //  190 :   8 - 0x8
      12'hBF: dout <= 8'b11110000; //  191 : 240 - 0xf0
      12'hC0: dout <= 8'b00111111; //  192 :  63 - 0x3f -- Sprite 0x18
      12'hC1: dout <= 8'b01000000; //  193 :  64 - 0x40
      12'hC2: dout <= 8'b01000000; //  194 :  64 - 0x40
      12'hC3: dout <= 8'b10000000; //  195 : 128 - 0x80
      12'hC4: dout <= 8'b10000000; //  196 : 128 - 0x80
      12'hC5: dout <= 8'b01111111; //  197 : 127 - 0x7f
      12'hC6: dout <= 8'b00000001; //  198 :   1 - 0x1
      12'hC7: dout <= 8'b01111111; //  199 : 127 - 0x7f
      12'hC8: dout <= 8'b11111100; //  200 : 252 - 0xfc -- Sprite 0x19
      12'hC9: dout <= 8'b00000010; //  201 :   2 - 0x2
      12'hCA: dout <= 8'b00000010; //  202 :   2 - 0x2
      12'hCB: dout <= 8'b00000001; //  203 :   1 - 0x1
      12'hCC: dout <= 8'b00000001; //  204 :   1 - 0x1
      12'hCD: dout <= 8'b11111110; //  205 : 254 - 0xfe
      12'hCE: dout <= 8'b10000000; //  206 : 128 - 0x80
      12'hCF: dout <= 8'b11111110; //  207 : 254 - 0xfe
      12'hD0: dout <= 8'b00000000; //  208 :   0 - 0x0 -- Sprite 0x1a
      12'hD1: dout <= 8'b00000000; //  209 :   0 - 0x0
      12'hD2: dout <= 8'b00111111; //  210 :  63 - 0x3f
      12'hD3: dout <= 8'b01000000; //  211 :  64 - 0x40
      12'hD4: dout <= 8'b01000000; //  212 :  64 - 0x40
      12'hD5: dout <= 8'b10000000; //  213 : 128 - 0x80
      12'hD6: dout <= 8'b10000000; //  214 : 128 - 0x80
      12'hD7: dout <= 8'b01111111; //  215 : 127 - 0x7f
      12'hD8: dout <= 8'b00000000; //  216 :   0 - 0x0 -- Sprite 0x1b
      12'hD9: dout <= 8'b00000000; //  217 :   0 - 0x0
      12'hDA: dout <= 8'b11111100; //  218 : 252 - 0xfc
      12'hDB: dout <= 8'b00000010; //  219 :   2 - 0x2
      12'hDC: dout <= 8'b00000010; //  220 :   2 - 0x2
      12'hDD: dout <= 8'b00000001; //  221 :   1 - 0x1
      12'hDE: dout <= 8'b00000001; //  222 :   1 - 0x1
      12'hDF: dout <= 8'b11111110; //  223 : 254 - 0xfe
      12'hE0: dout <= 8'b01111111; //  224 : 127 - 0x7f -- Sprite 0x1c
      12'hE1: dout <= 8'b10000000; //  225 : 128 - 0x80
      12'hE2: dout <= 8'b10000000; //  226 : 128 - 0x80
      12'hE3: dout <= 8'b10000000; //  227 : 128 - 0x80
      12'hE4: dout <= 8'b10011011; //  228 : 155 - 0x9b
      12'hE5: dout <= 8'b10100100; //  229 : 164 - 0xa4
      12'hE6: dout <= 8'b10100110; //  230 : 166 - 0xa6
      12'hE7: dout <= 8'b10000000; //  231 : 128 - 0x80
      12'hE8: dout <= 8'b10000000; //  232 : 128 - 0x80 -- Sprite 0x1d
      12'hE9: dout <= 8'b01111111; //  233 : 127 - 0x7f
      12'hEA: dout <= 8'b00000010; //  234 :   2 - 0x2
      12'hEB: dout <= 8'b00000010; //  235 :   2 - 0x2
      12'hEC: dout <= 8'b00000010; //  236 :   2 - 0x2
      12'hED: dout <= 8'b00000010; //  237 :   2 - 0x2
      12'hEE: dout <= 8'b00000010; //  238 :   2 - 0x2
      12'hEF: dout <= 8'b00001111; //  239 :  15 - 0xf
      12'hF0: dout <= 8'b11111110; //  240 : 254 - 0xfe -- Sprite 0x1e
      12'hF1: dout <= 8'b00000001; //  241 :   1 - 0x1
      12'hF2: dout <= 8'b00000001; //  242 :   1 - 0x1
      12'hF3: dout <= 8'b00000001; //  243 :   1 - 0x1
      12'hF4: dout <= 8'b01000001; //  244 :  65 - 0x41
      12'hF5: dout <= 8'b11110101; //  245 : 245 - 0xf5
      12'hF6: dout <= 8'b00011101; //  246 :  29 - 0x1d
      12'hF7: dout <= 8'b00000001; //  247 :   1 - 0x1
      12'hF8: dout <= 8'b00000001; //  248 :   1 - 0x1 -- Sprite 0x1f
      12'hF9: dout <= 8'b11111110; //  249 : 254 - 0xfe
      12'hFA: dout <= 8'b01000000; //  250 :  64 - 0x40
      12'hFB: dout <= 8'b01000000; //  251 :  64 - 0x40
      12'hFC: dout <= 8'b01000000; //  252 :  64 - 0x40
      12'hFD: dout <= 8'b01000000; //  253 :  64 - 0x40
      12'hFE: dout <= 8'b01000000; //  254 :  64 - 0x40
      12'hFF: dout <= 8'b11110000; //  255 : 240 - 0xf0
      12'h100: dout <= 8'b00000111; //  256 :   7 - 0x7 -- Sprite 0x20
      12'h101: dout <= 8'b00011111; //  257 :  31 - 0x1f
      12'h102: dout <= 8'b00111111; //  258 :  63 - 0x3f
      12'h103: dout <= 8'b01111111; //  259 : 127 - 0x7f
      12'h104: dout <= 8'b01111111; //  260 : 127 - 0x7f
      12'h105: dout <= 8'b11111111; //  261 : 255 - 0xff
      12'h106: dout <= 8'b11111111; //  262 : 255 - 0xff
      12'h107: dout <= 8'b11111111; //  263 : 255 - 0xff
      12'h108: dout <= 8'b11100000; //  264 : 224 - 0xe0 -- Sprite 0x21
      12'h109: dout <= 8'b11111000; //  265 : 248 - 0xf8
      12'h10A: dout <= 8'b11111100; //  266 : 252 - 0xfc
      12'h10B: dout <= 8'b11111110; //  267 : 254 - 0xfe
      12'h10C: dout <= 8'b11111110; //  268 : 254 - 0xfe
      12'h10D: dout <= 8'b11111111; //  269 : 255 - 0xff
      12'h10E: dout <= 8'b11111111; //  270 : 255 - 0xff
      12'h10F: dout <= 8'b11111111; //  271 : 255 - 0xff
      12'h110: dout <= 8'b00000111; //  272 :   7 - 0x7 -- Sprite 0x22
      12'h111: dout <= 8'b00011111; //  273 :  31 - 0x1f
      12'h112: dout <= 8'b00111111; //  274 :  63 - 0x3f
      12'h113: dout <= 8'b01111111; //  275 : 127 - 0x7f
      12'h114: dout <= 8'b01111111; //  276 : 127 - 0x7f
      12'h115: dout <= 8'b11111111; //  277 : 255 - 0xff
      12'h116: dout <= 8'b11111111; //  278 : 255 - 0xff
      12'h117: dout <= 8'b11111111; //  279 : 255 - 0xff
      12'h118: dout <= 8'b11100000; //  280 : 224 - 0xe0 -- Sprite 0x23
      12'h119: dout <= 8'b11111000; //  281 : 248 - 0xf8
      12'h11A: dout <= 8'b11111100; //  282 : 252 - 0xfc
      12'h11B: dout <= 8'b11111110; //  283 : 254 - 0xfe
      12'h11C: dout <= 8'b11111110; //  284 : 254 - 0xfe
      12'h11D: dout <= 8'b11111111; //  285 : 255 - 0xff
      12'h11E: dout <= 8'b11111111; //  286 : 255 - 0xff
      12'h11F: dout <= 8'b11111111; //  287 : 255 - 0xff
      12'h120: dout <= 8'b00000000; //  288 :   0 - 0x0 -- Sprite 0x24
      12'h121: dout <= 8'b00000000; //  289 :   0 - 0x0
      12'h122: dout <= 8'b00000000; //  290 :   0 - 0x0
      12'h123: dout <= 8'b00000000; //  291 :   0 - 0x0
      12'h124: dout <= 8'b00000000; //  292 :   0 - 0x0
      12'h125: dout <= 8'b00000000; //  293 :   0 - 0x0
      12'h126: dout <= 8'b00000000; //  294 :   0 - 0x0
      12'h127: dout <= 8'b00000000; //  295 :   0 - 0x0
      12'h128: dout <= 8'b00101111; //  296 :  47 - 0x2f -- Sprite 0x25
      12'h129: dout <= 8'b01001111; //  297 :  79 - 0x4f
      12'h12A: dout <= 8'b01001111; //  298 :  79 - 0x4f
      12'h12B: dout <= 8'b01001111; //  299 :  79 - 0x4f
      12'h12C: dout <= 8'b01001111; //  300 :  79 - 0x4f
      12'h12D: dout <= 8'b00100111; //  301 :  39 - 0x27
      12'h12E: dout <= 8'b00010000; //  302 :  16 - 0x10
      12'h12F: dout <= 8'b00001111; //  303 :  15 - 0xf
      12'h130: dout <= 8'b00000000; //  304 :   0 - 0x0 -- Sprite 0x26
      12'h131: dout <= 8'b11100000; //  305 : 224 - 0xe0
      12'h132: dout <= 8'b10100000; //  306 : 160 - 0xa0
      12'h133: dout <= 8'b00100000; //  307 :  32 - 0x20
      12'h134: dout <= 8'b11000000; //  308 : 192 - 0xc0
      12'h135: dout <= 8'b01000000; //  309 :  64 - 0x40
      12'h136: dout <= 8'b00110000; //  310 :  48 - 0x30
      12'h137: dout <= 8'b11101000; //  311 : 232 - 0xe8
      12'h138: dout <= 8'b11110100; //  312 : 244 - 0xf4 -- Sprite 0x27
      12'h139: dout <= 8'b11110010; //  313 : 242 - 0xf2
      12'h13A: dout <= 8'b11110010; //  314 : 242 - 0xf2
      12'h13B: dout <= 8'b11110010; //  315 : 242 - 0xf2
      12'h13C: dout <= 8'b11110010; //  316 : 242 - 0xf2
      12'h13D: dout <= 8'b11100100; //  317 : 228 - 0xe4
      12'h13E: dout <= 8'b00001000; //  318 :   8 - 0x8
      12'h13F: dout <= 8'b11110000; //  319 : 240 - 0xf0
      12'h140: dout <= 8'b11111111; //  320 : 255 - 0xff -- Sprite 0x28
      12'h141: dout <= 8'b11010101; //  321 : 213 - 0xd5
      12'h142: dout <= 8'b10100011; //  322 : 163 - 0xa3
      12'h143: dout <= 8'b11010111; //  323 : 215 - 0xd7
      12'h144: dout <= 8'b10001111; //  324 : 143 - 0x8f
      12'h145: dout <= 8'b11001111; //  325 : 207 - 0xcf
      12'h146: dout <= 8'b10001011; //  326 : 139 - 0x8b
      12'h147: dout <= 8'b11001011; //  327 : 203 - 0xcb
      12'h148: dout <= 8'b10001111; //  328 : 143 - 0x8f -- Sprite 0x29
      12'h149: dout <= 8'b11001111; //  329 : 207 - 0xcf
      12'h14A: dout <= 8'b10001111; //  330 : 143 - 0x8f
      12'h14B: dout <= 8'b11001111; //  331 : 207 - 0xcf
      12'h14C: dout <= 8'b10010000; //  332 : 144 - 0x90
      12'h14D: dout <= 8'b11100000; //  333 : 224 - 0xe0
      12'h14E: dout <= 8'b11101010; //  334 : 234 - 0xea
      12'h14F: dout <= 8'b11111111; //  335 : 255 - 0xff
      12'h150: dout <= 8'b11111111; //  336 : 255 - 0xff -- Sprite 0x2a
      12'h151: dout <= 8'b11011011; //  337 : 219 - 0xdb
      12'h152: dout <= 8'b11000111; //  338 : 199 - 0xc7
      12'h153: dout <= 8'b11101001; //  339 : 233 - 0xe9
      12'h154: dout <= 8'b11110011; //  340 : 243 - 0xf3
      12'h155: dout <= 8'b11110001; //  341 : 241 - 0xf1
      12'h156: dout <= 8'b11010011; //  342 : 211 - 0xd3
      12'h157: dout <= 8'b11010001; //  343 : 209 - 0xd1
      12'h158: dout <= 8'b11110011; //  344 : 243 - 0xf3 -- Sprite 0x2b
      12'h159: dout <= 8'b11110001; //  345 : 241 - 0xf1
      12'h15A: dout <= 8'b11110011; //  346 : 243 - 0xf3
      12'h15B: dout <= 8'b11110001; //  347 : 241 - 0xf1
      12'h15C: dout <= 8'b00001011; //  348 :  11 - 0xb
      12'h15D: dout <= 8'b00000101; //  349 :   5 - 0x5
      12'h15E: dout <= 8'b10101011; //  350 : 171 - 0xab
      12'h15F: dout <= 8'b11111111; //  351 : 255 - 0xff
      12'h160: dout <= 8'b00000000; //  352 :   0 - 0x0 -- Sprite 0x2c
      12'h161: dout <= 8'b00000000; //  353 :   0 - 0x0
      12'h162: dout <= 8'b00000000; //  354 :   0 - 0x0
      12'h163: dout <= 8'b00000000; //  355 :   0 - 0x0
      12'h164: dout <= 8'b00000000; //  356 :   0 - 0x0
      12'h165: dout <= 8'b00000000; //  357 :   0 - 0x0
      12'h166: dout <= 8'b00000000; //  358 :   0 - 0x0
      12'h167: dout <= 8'b00000000; //  359 :   0 - 0x0
      12'h168: dout <= 8'b00101111; //  360 :  47 - 0x2f -- Sprite 0x2d
      12'h169: dout <= 8'b01001111; //  361 :  79 - 0x4f
      12'h16A: dout <= 8'b01001111; //  362 :  79 - 0x4f
      12'h16B: dout <= 8'b01001111; //  363 :  79 - 0x4f
      12'h16C: dout <= 8'b01001111; //  364 :  79 - 0x4f
      12'h16D: dout <= 8'b00100111; //  365 :  39 - 0x27
      12'h16E: dout <= 8'b00010000; //  366 :  16 - 0x10
      12'h16F: dout <= 8'b00001111; //  367 :  15 - 0xf
      12'h170: dout <= 8'b00000000; //  368 :   0 - 0x0 -- Sprite 0x2e
      12'h171: dout <= 8'b00000000; //  369 :   0 - 0x0
      12'h172: dout <= 8'b00000000; //  370 :   0 - 0x0
      12'h173: dout <= 8'b00000000; //  371 :   0 - 0x0
      12'h174: dout <= 8'b00000000; //  372 :   0 - 0x0
      12'h175: dout <= 8'b00000000; //  373 :   0 - 0x0
      12'h176: dout <= 8'b00000000; //  374 :   0 - 0x0
      12'h177: dout <= 8'b00000000; //  375 :   0 - 0x0
      12'h178: dout <= 8'b11110100; //  376 : 244 - 0xf4 -- Sprite 0x2f
      12'h179: dout <= 8'b11110010; //  377 : 242 - 0xf2
      12'h17A: dout <= 8'b11110010; //  378 : 242 - 0xf2
      12'h17B: dout <= 8'b11110010; //  379 : 242 - 0xf2
      12'h17C: dout <= 8'b11110010; //  380 : 242 - 0xf2
      12'h17D: dout <= 8'b11100100; //  381 : 228 - 0xe4
      12'h17E: dout <= 8'b00001000; //  382 :   8 - 0x8
      12'h17F: dout <= 8'b11110000; //  383 : 240 - 0xf0
      12'h180: dout <= 8'b00011000; //  384 :  24 - 0x18 -- Sprite 0x30
      12'h181: dout <= 8'b00100100; //  385 :  36 - 0x24
      12'h182: dout <= 8'b01000010; //  386 :  66 - 0x42
      12'h183: dout <= 8'b10100101; //  387 : 165 - 0xa5
      12'h184: dout <= 8'b11100111; //  388 : 231 - 0xe7
      12'h185: dout <= 8'b00100100; //  389 :  36 - 0x24
      12'h186: dout <= 8'b00100100; //  390 :  36 - 0x24
      12'h187: dout <= 8'b00111100; //  391 :  60 - 0x3c
      12'h188: dout <= 8'b00111100; //  392 :  60 - 0x3c -- Sprite 0x31
      12'h189: dout <= 8'b00100100; //  393 :  36 - 0x24
      12'h18A: dout <= 8'b00100100; //  394 :  36 - 0x24
      12'h18B: dout <= 8'b01100110; //  395 : 102 - 0x66
      12'h18C: dout <= 8'b10100101; //  396 : 165 - 0xa5
      12'h18D: dout <= 8'b01000010; //  397 :  66 - 0x42
      12'h18E: dout <= 8'b00100100; //  398 :  36 - 0x24
      12'h18F: dout <= 8'b00011000; //  399 :  24 - 0x18
      12'h190: dout <= 8'b00000010; //  400 :   2 - 0x2 -- Sprite 0x32
      12'h191: dout <= 8'b00000010; //  401 :   2 - 0x2
      12'h192: dout <= 8'b00000011; //  402 :   3 - 0x3
      12'h193: dout <= 8'b00000010; //  403 :   2 - 0x2
      12'h194: dout <= 8'b00000010; //  404 :   2 - 0x2
      12'h195: dout <= 8'b00000010; //  405 :   2 - 0x2
      12'h196: dout <= 8'b00000011; //  406 :   3 - 0x3
      12'h197: dout <= 8'b00000010; //  407 :   2 - 0x2
      12'h198: dout <= 8'b01000000; //  408 :  64 - 0x40 -- Sprite 0x33
      12'h199: dout <= 8'b11000000; //  409 : 192 - 0xc0
      12'h19A: dout <= 8'b01000000; //  410 :  64 - 0x40
      12'h19B: dout <= 8'b01000000; //  411 :  64 - 0x40
      12'h19C: dout <= 8'b01000000; //  412 :  64 - 0x40
      12'h19D: dout <= 8'b11000000; //  413 : 192 - 0xc0
      12'h19E: dout <= 8'b01000000; //  414 :  64 - 0x40
      12'h19F: dout <= 8'b01000000; //  415 :  64 - 0x40
      12'h1A0: dout <= 8'b00000000; //  416 :   0 - 0x0 -- Sprite 0x34
      12'h1A1: dout <= 8'b00011000; //  417 :  24 - 0x18
      12'h1A2: dout <= 8'b00111100; //  418 :  60 - 0x3c
      12'h1A3: dout <= 8'b01100010; //  419 :  98 - 0x62
      12'h1A4: dout <= 8'b01100001; //  420 :  97 - 0x61
      12'h1A5: dout <= 8'b11000000; //  421 : 192 - 0xc0
      12'h1A6: dout <= 8'b11000000; //  422 : 192 - 0xc0
      12'h1A7: dout <= 8'b11000000; //  423 : 192 - 0xc0
      12'h1A8: dout <= 8'b01100000; //  424 :  96 - 0x60 -- Sprite 0x35
      12'h1A9: dout <= 8'b01100000; //  425 :  96 - 0x60
      12'h1AA: dout <= 8'b00110000; //  426 :  48 - 0x30
      12'h1AB: dout <= 8'b00011000; //  427 :  24 - 0x18
      12'h1AC: dout <= 8'b00001100; //  428 :  12 - 0xc
      12'h1AD: dout <= 8'b00000110; //  429 :   6 - 0x6
      12'h1AE: dout <= 8'b00000010; //  430 :   2 - 0x2
      12'h1AF: dout <= 8'b00000001; //  431 :   1 - 0x1
      12'h1B0: dout <= 8'b00000000; //  432 :   0 - 0x0 -- Sprite 0x36
      12'h1B1: dout <= 8'b00011000; //  433 :  24 - 0x18
      12'h1B2: dout <= 8'b00100100; //  434 :  36 - 0x24
      12'h1B3: dout <= 8'b01000010; //  435 :  66 - 0x42
      12'h1B4: dout <= 8'b10000010; //  436 : 130 - 0x82
      12'h1B5: dout <= 8'b00000001; //  437 :   1 - 0x1
      12'h1B6: dout <= 8'b00000001; //  438 :   1 - 0x1
      12'h1B7: dout <= 8'b00000001; //  439 :   1 - 0x1
      12'h1B8: dout <= 8'b00000010; //  440 :   2 - 0x2 -- Sprite 0x37
      12'h1B9: dout <= 8'b00000010; //  441 :   2 - 0x2
      12'h1BA: dout <= 8'b00000100; //  442 :   4 - 0x4
      12'h1BB: dout <= 8'b00001000; //  443 :   8 - 0x8
      12'h1BC: dout <= 8'b00010000; //  444 :  16 - 0x10
      12'h1BD: dout <= 8'b00100000; //  445 :  32 - 0x20
      12'h1BE: dout <= 8'b01000000; //  446 :  64 - 0x40
      12'h1BF: dout <= 8'b10000000; //  447 : 128 - 0x80
      12'h1C0: dout <= 8'b00000000; //  448 :   0 - 0x0 -- Sprite 0x38
      12'h1C1: dout <= 8'b00000110; //  449 :   6 - 0x6
      12'h1C2: dout <= 8'b00001101; //  450 :  13 - 0xd
      12'h1C3: dout <= 8'b00001100; //  451 :  12 - 0xc
      12'h1C4: dout <= 8'b00001100; //  452 :  12 - 0xc
      12'h1C5: dout <= 8'b00000110; //  453 :   6 - 0x6
      12'h1C6: dout <= 8'b00000010; //  454 :   2 - 0x2
      12'h1C7: dout <= 8'b00000001; //  455 :   1 - 0x1
      12'h1C8: dout <= 8'b11111111; //  456 : 255 - 0xff -- Sprite 0x39
      12'h1C9: dout <= 8'b00000000; //  457 :   0 - 0x0
      12'h1CA: dout <= 8'b00000000; //  458 :   0 - 0x0
      12'h1CB: dout <= 8'b00000000; //  459 :   0 - 0x0
      12'h1CC: dout <= 8'b00000000; //  460 :   0 - 0x0
      12'h1CD: dout <= 8'b00000000; //  461 :   0 - 0x0
      12'h1CE: dout <= 8'b00000000; //  462 :   0 - 0x0
      12'h1CF: dout <= 8'b00000000; //  463 :   0 - 0x0
      12'h1D0: dout <= 8'b00000000; //  464 :   0 - 0x0 -- Sprite 0x3a
      12'h1D1: dout <= 8'b01100000; //  465 :  96 - 0x60
      12'h1D2: dout <= 8'b10010000; //  466 : 144 - 0x90
      12'h1D3: dout <= 8'b00010000; //  467 :  16 - 0x10
      12'h1D4: dout <= 8'b00010000; //  468 :  16 - 0x10
      12'h1D5: dout <= 8'b00100000; //  469 :  32 - 0x20
      12'h1D6: dout <= 8'b01000000; //  470 :  64 - 0x40
      12'h1D7: dout <= 8'b10000000; //  471 : 128 - 0x80
      12'h1D8: dout <= 8'b00000000; //  472 :   0 - 0x0 -- Sprite 0x3b
      12'h1D9: dout <= 8'b01010100; //  473 :  84 - 0x54
      12'h1DA: dout <= 8'b00000010; //  474 :   2 - 0x2
      12'h1DB: dout <= 8'b01000000; //  475 :  64 - 0x40
      12'h1DC: dout <= 8'b00000010; //  476 :   2 - 0x2
      12'h1DD: dout <= 8'b01000000; //  477 :  64 - 0x40
      12'h1DE: dout <= 8'b00101010; //  478 :  42 - 0x2a
      12'h1DF: dout <= 8'b00000000; //  479 :   0 - 0x0
      12'h1E0: dout <= 8'b11111111; //  480 : 255 - 0xff -- Sprite 0x3c
      12'h1E1: dout <= 8'b11111111; //  481 : 255 - 0xff
      12'h1E2: dout <= 8'b11111111; //  482 : 255 - 0xff
      12'h1E3: dout <= 8'b11111111; //  483 : 255 - 0xff
      12'h1E4: dout <= 8'b11111111; //  484 : 255 - 0xff
      12'h1E5: dout <= 8'b11111111; //  485 : 255 - 0xff
      12'h1E6: dout <= 8'b11111111; //  486 : 255 - 0xff
      12'h1E7: dout <= 8'b11111111; //  487 : 255 - 0xff
      12'h1E8: dout <= 8'b00000000; //  488 :   0 - 0x0 -- Sprite 0x3d
      12'h1E9: dout <= 8'b00000000; //  489 :   0 - 0x0
      12'h1EA: dout <= 8'b00000000; //  490 :   0 - 0x0
      12'h1EB: dout <= 8'b00000000; //  491 :   0 - 0x0
      12'h1EC: dout <= 8'b00000000; //  492 :   0 - 0x0
      12'h1ED: dout <= 8'b00000000; //  493 :   0 - 0x0
      12'h1EE: dout <= 8'b00000000; //  494 :   0 - 0x0
      12'h1EF: dout <= 8'b00000000; //  495 :   0 - 0x0
      12'h1F0: dout <= 8'b11111111; //  496 : 255 - 0xff -- Sprite 0x3e
      12'h1F1: dout <= 8'b11111111; //  497 : 255 - 0xff
      12'h1F2: dout <= 8'b11111111; //  498 : 255 - 0xff
      12'h1F3: dout <= 8'b11111111; //  499 : 255 - 0xff
      12'h1F4: dout <= 8'b11111111; //  500 : 255 - 0xff
      12'h1F5: dout <= 8'b11111111; //  501 : 255 - 0xff
      12'h1F6: dout <= 8'b11111111; //  502 : 255 - 0xff
      12'h1F7: dout <= 8'b11111111; //  503 : 255 - 0xff
      12'h1F8: dout <= 8'b00000000; //  504 :   0 - 0x0 -- Sprite 0x3f
      12'h1F9: dout <= 8'b00000000; //  505 :   0 - 0x0
      12'h1FA: dout <= 8'b00000000; //  506 :   0 - 0x0
      12'h1FB: dout <= 8'b00000000; //  507 :   0 - 0x0
      12'h1FC: dout <= 8'b00000000; //  508 :   0 - 0x0
      12'h1FD: dout <= 8'b00000000; //  509 :   0 - 0x0
      12'h1FE: dout <= 8'b00000000; //  510 :   0 - 0x0
      12'h1FF: dout <= 8'b00000000; //  511 :   0 - 0x0
      12'h200: dout <= 8'b00111100; //  512 :  60 - 0x3c -- Sprite 0x40
      12'h201: dout <= 8'b01000010; //  513 :  66 - 0x42
      12'h202: dout <= 8'b10011001; //  514 : 153 - 0x99
      12'h203: dout <= 8'b10100101; //  515 : 165 - 0xa5
      12'h204: dout <= 8'b10100101; //  516 : 165 - 0xa5
      12'h205: dout <= 8'b10011010; //  517 : 154 - 0x9a
      12'h206: dout <= 8'b01000000; //  518 :  64 - 0x40
      12'h207: dout <= 8'b00111100; //  519 :  60 - 0x3c
      12'h208: dout <= 8'b00001100; //  520 :  12 - 0xc -- Sprite 0x41
      12'h209: dout <= 8'b00010010; //  521 :  18 - 0x12
      12'h20A: dout <= 8'b00100010; //  522 :  34 - 0x22
      12'h20B: dout <= 8'b00100010; //  523 :  34 - 0x22
      12'h20C: dout <= 8'b01111110; //  524 : 126 - 0x7e
      12'h20D: dout <= 8'b00100010; //  525 :  34 - 0x22
      12'h20E: dout <= 8'b00100100; //  526 :  36 - 0x24
      12'h20F: dout <= 8'b00000000; //  527 :   0 - 0x0
      12'h210: dout <= 8'b00111100; //  528 :  60 - 0x3c -- Sprite 0x42
      12'h211: dout <= 8'b01000010; //  529 :  66 - 0x42
      12'h212: dout <= 8'b01010010; //  530 :  82 - 0x52
      12'h213: dout <= 8'b00011100; //  531 :  28 - 0x1c
      12'h214: dout <= 8'b00010010; //  532 :  18 - 0x12
      12'h215: dout <= 8'b00110010; //  533 :  50 - 0x32
      12'h216: dout <= 8'b00011100; //  534 :  28 - 0x1c
      12'h217: dout <= 8'b00000000; //  535 :   0 - 0x0
      12'h218: dout <= 8'b00011000; //  536 :  24 - 0x18 -- Sprite 0x43
      12'h219: dout <= 8'b00100100; //  537 :  36 - 0x24
      12'h21A: dout <= 8'b01010100; //  538 :  84 - 0x54
      12'h21B: dout <= 8'b01001000; //  539 :  72 - 0x48
      12'h21C: dout <= 8'b01000010; //  540 :  66 - 0x42
      12'h21D: dout <= 8'b00100100; //  541 :  36 - 0x24
      12'h21E: dout <= 8'b00011000; //  542 :  24 - 0x18
      12'h21F: dout <= 8'b00000000; //  543 :   0 - 0x0
      12'h220: dout <= 8'b01011000; //  544 :  88 - 0x58 -- Sprite 0x44
      12'h221: dout <= 8'b11100100; //  545 : 228 - 0xe4
      12'h222: dout <= 8'b01000010; //  546 :  66 - 0x42
      12'h223: dout <= 8'b01000010; //  547 :  66 - 0x42
      12'h224: dout <= 8'b00100010; //  548 :  34 - 0x22
      12'h225: dout <= 8'b01100100; //  549 : 100 - 0x64
      12'h226: dout <= 8'b00111000; //  550 :  56 - 0x38
      12'h227: dout <= 8'b00000000; //  551 :   0 - 0x0
      12'h228: dout <= 8'b00011100; //  552 :  28 - 0x1c -- Sprite 0x45
      12'h229: dout <= 8'b00100000; //  553 :  32 - 0x20
      12'h22A: dout <= 8'b00100000; //  554 :  32 - 0x20
      12'h22B: dout <= 8'b00101100; //  555 :  44 - 0x2c
      12'h22C: dout <= 8'b01110000; //  556 : 112 - 0x70
      12'h22D: dout <= 8'b00100010; //  557 :  34 - 0x22
      12'h22E: dout <= 8'b00011100; //  558 :  28 - 0x1c
      12'h22F: dout <= 8'b00000000; //  559 :   0 - 0x0
      12'h230: dout <= 8'b00011100; //  560 :  28 - 0x1c -- Sprite 0x46
      12'h231: dout <= 8'b00100000; //  561 :  32 - 0x20
      12'h232: dout <= 8'b00100000; //  562 :  32 - 0x20
      12'h233: dout <= 8'b00101100; //  563 :  44 - 0x2c
      12'h234: dout <= 8'b01110000; //  564 : 112 - 0x70
      12'h235: dout <= 8'b00010000; //  565 :  16 - 0x10
      12'h236: dout <= 8'b00010000; //  566 :  16 - 0x10
      12'h237: dout <= 8'b00000000; //  567 :   0 - 0x0
      12'h238: dout <= 8'b00011000; //  568 :  24 - 0x18 -- Sprite 0x47
      12'h239: dout <= 8'b00100100; //  569 :  36 - 0x24
      12'h23A: dout <= 8'b01000000; //  570 :  64 - 0x40
      12'h23B: dout <= 8'b01001110; //  571 :  78 - 0x4e
      12'h23C: dout <= 8'b01000010; //  572 :  66 - 0x42
      12'h23D: dout <= 8'b00100100; //  573 :  36 - 0x24
      12'h23E: dout <= 8'b00011000; //  574 :  24 - 0x18
      12'h23F: dout <= 8'b00000000; //  575 :   0 - 0x0
      12'h240: dout <= 8'b00100000; //  576 :  32 - 0x20 -- Sprite 0x48
      12'h241: dout <= 8'b01000100; //  577 :  68 - 0x44
      12'h242: dout <= 8'b01000100; //  578 :  68 - 0x44
      12'h243: dout <= 8'b01000100; //  579 :  68 - 0x44
      12'h244: dout <= 8'b11111100; //  580 : 252 - 0xfc
      12'h245: dout <= 8'b01000100; //  581 :  68 - 0x44
      12'h246: dout <= 8'b01001000; //  582 :  72 - 0x48
      12'h247: dout <= 8'b00000000; //  583 :   0 - 0x0
      12'h248: dout <= 8'b00010000; //  584 :  16 - 0x10 -- Sprite 0x49
      12'h249: dout <= 8'b00010000; //  585 :  16 - 0x10
      12'h24A: dout <= 8'b00010000; //  586 :  16 - 0x10
      12'h24B: dout <= 8'b00010000; //  587 :  16 - 0x10
      12'h24C: dout <= 8'b00010000; //  588 :  16 - 0x10
      12'h24D: dout <= 8'b00001000; //  589 :   8 - 0x8
      12'h24E: dout <= 8'b00001000; //  590 :   8 - 0x8
      12'h24F: dout <= 8'b00000000; //  591 :   0 - 0x0
      12'h250: dout <= 8'b00001000; //  592 :   8 - 0x8 -- Sprite 0x4a
      12'h251: dout <= 8'b00001000; //  593 :   8 - 0x8
      12'h252: dout <= 8'b00000100; //  594 :   4 - 0x4
      12'h253: dout <= 8'b00000100; //  595 :   4 - 0x4
      12'h254: dout <= 8'b01000100; //  596 :  68 - 0x44
      12'h255: dout <= 8'b01001000; //  597 :  72 - 0x48
      12'h256: dout <= 8'b00110000; //  598 :  48 - 0x30
      12'h257: dout <= 8'b00000000; //  599 :   0 - 0x0
      12'h258: dout <= 8'b01000100; //  600 :  68 - 0x44 -- Sprite 0x4b
      12'h259: dout <= 8'b01000100; //  601 :  68 - 0x44
      12'h25A: dout <= 8'b01001000; //  602 :  72 - 0x48
      12'h25B: dout <= 8'b01110000; //  603 : 112 - 0x70
      12'h25C: dout <= 8'b01001000; //  604 :  72 - 0x48
      12'h25D: dout <= 8'b00100100; //  605 :  36 - 0x24
      12'h25E: dout <= 8'b00100010; //  606 :  34 - 0x22
      12'h25F: dout <= 8'b00000000; //  607 :   0 - 0x0
      12'h260: dout <= 8'b00010000; //  608 :  16 - 0x10 -- Sprite 0x4c
      12'h261: dout <= 8'b00100000; //  609 :  32 - 0x20
      12'h262: dout <= 8'b00100000; //  610 :  32 - 0x20
      12'h263: dout <= 8'b00100000; //  611 :  32 - 0x20
      12'h264: dout <= 8'b01000000; //  612 :  64 - 0x40
      12'h265: dout <= 8'b01000000; //  613 :  64 - 0x40
      12'h266: dout <= 8'b01000110; //  614 :  70 - 0x46
      12'h267: dout <= 8'b00111000; //  615 :  56 - 0x38
      12'h268: dout <= 8'b00100100; //  616 :  36 - 0x24 -- Sprite 0x4d
      12'h269: dout <= 8'b01011010; //  617 :  90 - 0x5a
      12'h26A: dout <= 8'b01011010; //  618 :  90 - 0x5a
      12'h26B: dout <= 8'b01011010; //  619 :  90 - 0x5a
      12'h26C: dout <= 8'b01000010; //  620 :  66 - 0x42
      12'h26D: dout <= 8'b01000010; //  621 :  66 - 0x42
      12'h26E: dout <= 8'b00100010; //  622 :  34 - 0x22
      12'h26F: dout <= 8'b00000000; //  623 :   0 - 0x0
      12'h270: dout <= 8'b00100100; //  624 :  36 - 0x24 -- Sprite 0x4e
      12'h271: dout <= 8'b01010010; //  625 :  82 - 0x52
      12'h272: dout <= 8'b01010010; //  626 :  82 - 0x52
      12'h273: dout <= 8'b01010010; //  627 :  82 - 0x52
      12'h274: dout <= 8'b01010010; //  628 :  82 - 0x52
      12'h275: dout <= 8'b01010010; //  629 :  82 - 0x52
      12'h276: dout <= 8'b01001100; //  630 :  76 - 0x4c
      12'h277: dout <= 8'b00000000; //  631 :   0 - 0x0
      12'h278: dout <= 8'b00111000; //  632 :  56 - 0x38 -- Sprite 0x4f
      12'h279: dout <= 8'b01000100; //  633 :  68 - 0x44
      12'h27A: dout <= 8'b10000010; //  634 : 130 - 0x82
      12'h27B: dout <= 8'b10000010; //  635 : 130 - 0x82
      12'h27C: dout <= 8'b10000010; //  636 : 130 - 0x82
      12'h27D: dout <= 8'b01000100; //  637 :  68 - 0x44
      12'h27E: dout <= 8'b00111000; //  638 :  56 - 0x38
      12'h27F: dout <= 8'b00000000; //  639 :   0 - 0x0
      12'h280: dout <= 8'b01111111; //  640 : 127 - 0x7f -- Sprite 0x50
      12'h281: dout <= 8'b11000000; //  641 : 192 - 0xc0
      12'h282: dout <= 8'b10000000; //  642 : 128 - 0x80
      12'h283: dout <= 8'b10000000; //  643 : 128 - 0x80
      12'h284: dout <= 8'b10000000; //  644 : 128 - 0x80
      12'h285: dout <= 8'b11000011; //  645 : 195 - 0xc3
      12'h286: dout <= 8'b11111111; //  646 : 255 - 0xff
      12'h287: dout <= 8'b11111111; //  647 : 255 - 0xff
      12'h288: dout <= 8'b11111110; //  648 : 254 - 0xfe -- Sprite 0x51
      12'h289: dout <= 8'b00000011; //  649 :   3 - 0x3
      12'h28A: dout <= 8'b00000001; //  650 :   1 - 0x1
      12'h28B: dout <= 8'b00000001; //  651 :   1 - 0x1
      12'h28C: dout <= 8'b00000001; //  652 :   1 - 0x1
      12'h28D: dout <= 8'b11000011; //  653 : 195 - 0xc3
      12'h28E: dout <= 8'b11111111; //  654 : 255 - 0xff
      12'h28F: dout <= 8'b11111111; //  655 : 255 - 0xff
      12'h290: dout <= 8'b00000000; //  656 :   0 - 0x0 -- Sprite 0x52
      12'h291: dout <= 8'b00000111; //  657 :   7 - 0x7
      12'h292: dout <= 8'b00001100; //  658 :  12 - 0xc
      12'h293: dout <= 8'b00011000; //  659 :  24 - 0x18
      12'h294: dout <= 8'b00110000; //  660 :  48 - 0x30
      12'h295: dout <= 8'b01100000; //  661 :  96 - 0x60
      12'h296: dout <= 8'b01000000; //  662 :  64 - 0x40
      12'h297: dout <= 8'b01001111; //  663 :  79 - 0x4f
      12'h298: dout <= 8'b00000000; //  664 :   0 - 0x0 -- Sprite 0x53
      12'h299: dout <= 8'b11110000; //  665 : 240 - 0xf0
      12'h29A: dout <= 8'b01010000; //  666 :  80 - 0x50
      12'h29B: dout <= 8'b01001000; //  667 :  72 - 0x48
      12'h29C: dout <= 8'b01001100; //  668 :  76 - 0x4c
      12'h29D: dout <= 8'b01000100; //  669 :  68 - 0x44
      12'h29E: dout <= 8'b10000010; //  670 : 130 - 0x82
      12'h29F: dout <= 8'b10000011; //  671 : 131 - 0x83
      12'h2A0: dout <= 8'b01111111; //  672 : 127 - 0x7f -- Sprite 0x54
      12'h2A1: dout <= 8'b11011110; //  673 : 222 - 0xde
      12'h2A2: dout <= 8'b10001110; //  674 : 142 - 0x8e
      12'h2A3: dout <= 8'b11000101; //  675 : 197 - 0xc5
      12'h2A4: dout <= 8'b10010010; //  676 : 146 - 0x92
      12'h2A5: dout <= 8'b11000111; //  677 : 199 - 0xc7
      12'h2A6: dout <= 8'b11100010; //  678 : 226 - 0xe2
      12'h2A7: dout <= 8'b11010000; //  679 : 208 - 0xd0
      12'h2A8: dout <= 8'b11111111; //  680 : 255 - 0xff -- Sprite 0x55
      12'h2A9: dout <= 8'b11011110; //  681 : 222 - 0xde
      12'h2AA: dout <= 8'b10001110; //  682 : 142 - 0x8e
      12'h2AB: dout <= 8'b11000101; //  683 : 197 - 0xc5
      12'h2AC: dout <= 8'b10010010; //  684 : 146 - 0x92
      12'h2AD: dout <= 8'b01000111; //  685 :  71 - 0x47
      12'h2AE: dout <= 8'b11100010; //  686 : 226 - 0xe2
      12'h2AF: dout <= 8'b01010000; //  687 :  80 - 0x50
      12'h2B0: dout <= 8'b11111110; //  688 : 254 - 0xfe -- Sprite 0x56
      12'h2B1: dout <= 8'b11011111; //  689 : 223 - 0xdf
      12'h2B2: dout <= 8'b10001111; //  690 : 143 - 0x8f
      12'h2B3: dout <= 8'b11000101; //  691 : 197 - 0xc5
      12'h2B4: dout <= 8'b10010011; //  692 : 147 - 0x93
      12'h2B5: dout <= 8'b01000111; //  693 :  71 - 0x47
      12'h2B6: dout <= 8'b11100011; //  694 : 227 - 0xe3
      12'h2B7: dout <= 8'b01010001; //  695 :  81 - 0x51
      12'h2B8: dout <= 8'b01111111; //  696 : 127 - 0x7f -- Sprite 0x57
      12'h2B9: dout <= 8'b10000000; //  697 : 128 - 0x80
      12'h2BA: dout <= 8'b10110011; //  698 : 179 - 0xb3
      12'h2BB: dout <= 8'b01001100; //  699 :  76 - 0x4c
      12'h2BC: dout <= 8'b00111111; //  700 :  63 - 0x3f
      12'h2BD: dout <= 8'b00000011; //  701 :   3 - 0x3
      12'h2BE: dout <= 8'b00000000; //  702 :   0 - 0x0
      12'h2BF: dout <= 8'b00000000; //  703 :   0 - 0x0
      12'h2C0: dout <= 8'b11111111; //  704 : 255 - 0xff -- Sprite 0x58
      12'h2C1: dout <= 8'b00000000; //  705 :   0 - 0x0
      12'h2C2: dout <= 8'b00110011; //  706 :  51 - 0x33
      12'h2C3: dout <= 8'b11001100; //  707 : 204 - 0xcc
      12'h2C4: dout <= 8'b00110011; //  708 :  51 - 0x33
      12'h2C5: dout <= 8'b11111111; //  709 : 255 - 0xff
      12'h2C6: dout <= 8'b00000000; //  710 :   0 - 0x0
      12'h2C7: dout <= 8'b00000000; //  711 :   0 - 0x0
      12'h2C8: dout <= 8'b11111110; //  712 : 254 - 0xfe -- Sprite 0x59
      12'h2C9: dout <= 8'b00000001; //  713 :   1 - 0x1
      12'h2CA: dout <= 8'b00110011; //  714 :  51 - 0x33
      12'h2CB: dout <= 8'b11001110; //  715 : 206 - 0xce
      12'h2CC: dout <= 8'b00111100; //  716 :  60 - 0x3c
      12'h2CD: dout <= 8'b11000000; //  717 : 192 - 0xc0
      12'h2CE: dout <= 8'b00000000; //  718 :   0 - 0x0
      12'h2CF: dout <= 8'b00000000; //  719 :   0 - 0x0
      12'h2D0: dout <= 8'b00000000; //  720 :   0 - 0x0 -- Sprite 0x5a
      12'h2D1: dout <= 8'b00000000; //  721 :   0 - 0x0
      12'h2D2: dout <= 8'b00000000; //  722 :   0 - 0x0
      12'h2D3: dout <= 8'b00000000; //  723 :   0 - 0x0
      12'h2D4: dout <= 8'b00000000; //  724 :   0 - 0x0
      12'h2D5: dout <= 8'b00000000; //  725 :   0 - 0x0
      12'h2D6: dout <= 8'b00000000; //  726 :   0 - 0x0
      12'h2D7: dout <= 8'b00000000; //  727 :   0 - 0x0
      12'h2D8: dout <= 8'b00000000; //  728 :   0 - 0x0 -- Sprite 0x5b
      12'h2D9: dout <= 8'b00000000; //  729 :   0 - 0x0
      12'h2DA: dout <= 8'b00000000; //  730 :   0 - 0x0
      12'h2DB: dout <= 8'b00000001; //  731 :   1 - 0x1
      12'h2DC: dout <= 8'b00000011; //  732 :   3 - 0x3
      12'h2DD: dout <= 8'b00000011; //  733 :   3 - 0x3
      12'h2DE: dout <= 8'b00000111; //  734 :   7 - 0x7
      12'h2DF: dout <= 8'b00111111; //  735 :  63 - 0x3f
      12'h2E0: dout <= 8'b00000000; //  736 :   0 - 0x0 -- Sprite 0x5c
      12'h2E1: dout <= 8'b00000001; //  737 :   1 - 0x1
      12'h2E2: dout <= 8'b01111111; //  738 : 127 - 0x7f
      12'h2E3: dout <= 8'b11111111; //  739 : 255 - 0xff
      12'h2E4: dout <= 8'b11111111; //  740 : 255 - 0xff
      12'h2E5: dout <= 8'b11111111; //  741 : 255 - 0xff
      12'h2E6: dout <= 8'b11111111; //  742 : 255 - 0xff
      12'h2E7: dout <= 8'b11111111; //  743 : 255 - 0xff
      12'h2E8: dout <= 8'b11111111; //  744 : 255 - 0xff -- Sprite 0x5d
      12'h2E9: dout <= 8'b11111111; //  745 : 255 - 0xff
      12'h2EA: dout <= 8'b11111111; //  746 : 255 - 0xff
      12'h2EB: dout <= 8'b11111111; //  747 : 255 - 0xff
      12'h2EC: dout <= 8'b11111111; //  748 : 255 - 0xff
      12'h2ED: dout <= 8'b11111111; //  749 : 255 - 0xff
      12'h2EE: dout <= 8'b11111111; //  750 : 255 - 0xff
      12'h2EF: dout <= 8'b11111111; //  751 : 255 - 0xff
      12'h2F0: dout <= 8'b00000000; //  752 :   0 - 0x0 -- Sprite 0x5e
      12'h2F1: dout <= 8'b10000000; //  753 : 128 - 0x80
      12'h2F2: dout <= 8'b11111110; //  754 : 254 - 0xfe
      12'h2F3: dout <= 8'b11111111; //  755 : 255 - 0xff
      12'h2F4: dout <= 8'b11111111; //  756 : 255 - 0xff
      12'h2F5: dout <= 8'b11111111; //  757 : 255 - 0xff
      12'h2F6: dout <= 8'b11111111; //  758 : 255 - 0xff
      12'h2F7: dout <= 8'b11111111; //  759 : 255 - 0xff
      12'h2F8: dout <= 8'b00000000; //  760 :   0 - 0x0 -- Sprite 0x5f
      12'h2F9: dout <= 8'b00000000; //  761 :   0 - 0x0
      12'h2FA: dout <= 8'b00000000; //  762 :   0 - 0x0
      12'h2FB: dout <= 8'b10000000; //  763 : 128 - 0x80
      12'h2FC: dout <= 8'b11000000; //  764 : 192 - 0xc0
      12'h2FD: dout <= 8'b11000000; //  765 : 192 - 0xc0
      12'h2FE: dout <= 8'b11100000; //  766 : 224 - 0xe0
      12'h2FF: dout <= 8'b11111000; //  767 : 248 - 0xf8
      12'h300: dout <= 8'b11111111; //  768 : 255 - 0xff -- Sprite 0x60
      12'h301: dout <= 8'b11111111; //  769 : 255 - 0xff
      12'h302: dout <= 8'b11111111; //  770 : 255 - 0xff
      12'h303: dout <= 8'b11111111; //  771 : 255 - 0xff
      12'h304: dout <= 8'b11111111; //  772 : 255 - 0xff
      12'h305: dout <= 8'b11111111; //  773 : 255 - 0xff
      12'h306: dout <= 8'b11111111; //  774 : 255 - 0xff
      12'h307: dout <= 8'b11111111; //  775 : 255 - 0xff
      12'h308: dout <= 8'b11111111; //  776 : 255 - 0xff -- Sprite 0x61
      12'h309: dout <= 8'b11111111; //  777 : 255 - 0xff
      12'h30A: dout <= 8'b11111111; //  778 : 255 - 0xff
      12'h30B: dout <= 8'b11111111; //  779 : 255 - 0xff
      12'h30C: dout <= 8'b11111111; //  780 : 255 - 0xff
      12'h30D: dout <= 8'b11111111; //  781 : 255 - 0xff
      12'h30E: dout <= 8'b11111111; //  782 : 255 - 0xff
      12'h30F: dout <= 8'b11111111; //  783 : 255 - 0xff
      12'h310: dout <= 8'b01111000; //  784 : 120 - 0x78 -- Sprite 0x62
      12'h311: dout <= 8'b01100000; //  785 :  96 - 0x60
      12'h312: dout <= 8'b01000000; //  786 :  64 - 0x40
      12'h313: dout <= 8'b01000000; //  787 :  64 - 0x40
      12'h314: dout <= 8'b01000000; //  788 :  64 - 0x40
      12'h315: dout <= 8'b01100000; //  789 :  96 - 0x60
      12'h316: dout <= 8'b00110000; //  790 :  48 - 0x30
      12'h317: dout <= 8'b00011111; //  791 :  31 - 0x1f
      12'h318: dout <= 8'b10000001; //  792 : 129 - 0x81 -- Sprite 0x63
      12'h319: dout <= 8'b10000011; //  793 : 131 - 0x83
      12'h31A: dout <= 8'b11000001; //  794 : 193 - 0xc1
      12'h31B: dout <= 8'b01000011; //  795 :  67 - 0x43
      12'h31C: dout <= 8'b01000001; //  796 :  65 - 0x41
      12'h31D: dout <= 8'b01100011; //  797 :  99 - 0x63
      12'h31E: dout <= 8'b00100110; //  798 :  38 - 0x26
      12'h31F: dout <= 8'b11111000; //  799 : 248 - 0xf8
      12'h320: dout <= 8'b10111001; //  800 : 185 - 0xb9 -- Sprite 0x64
      12'h321: dout <= 8'b10010100; //  801 : 148 - 0x94
      12'h322: dout <= 8'b10001110; //  802 : 142 - 0x8e
      12'h323: dout <= 8'b11000101; //  803 : 197 - 0xc5
      12'h324: dout <= 8'b10010010; //  804 : 146 - 0x92
      12'h325: dout <= 8'b11000111; //  805 : 199 - 0xc7
      12'h326: dout <= 8'b11100010; //  806 : 226 - 0xe2
      12'h327: dout <= 8'b11010000; //  807 : 208 - 0xd0
      12'h328: dout <= 8'b10111001; //  808 : 185 - 0xb9 -- Sprite 0x65
      12'h329: dout <= 8'b00010100; //  809 :  20 - 0x14
      12'h32A: dout <= 8'b10001110; //  810 : 142 - 0x8e
      12'h32B: dout <= 8'b11000101; //  811 : 197 - 0xc5
      12'h32C: dout <= 8'b10010010; //  812 : 146 - 0x92
      12'h32D: dout <= 8'b01000111; //  813 :  71 - 0x47
      12'h32E: dout <= 8'b11100010; //  814 : 226 - 0xe2
      12'h32F: dout <= 8'b01010000; //  815 :  80 - 0x50
      12'h330: dout <= 8'b10111001; //  816 : 185 - 0xb9 -- Sprite 0x66
      12'h331: dout <= 8'b00010101; //  817 :  21 - 0x15
      12'h332: dout <= 8'b10001111; //  818 : 143 - 0x8f
      12'h333: dout <= 8'b11000101; //  819 : 197 - 0xc5
      12'h334: dout <= 8'b10010011; //  820 : 147 - 0x93
      12'h335: dout <= 8'b01000111; //  821 :  71 - 0x47
      12'h336: dout <= 8'b11100011; //  822 : 227 - 0xe3
      12'h337: dout <= 8'b01010001; //  823 :  81 - 0x51
      12'h338: dout <= 8'b01111111; //  824 : 127 - 0x7f -- Sprite 0x67
      12'h339: dout <= 8'b10000000; //  825 : 128 - 0x80
      12'h33A: dout <= 8'b11001100; //  826 : 204 - 0xcc
      12'h33B: dout <= 8'b01111111; //  827 : 127 - 0x7f
      12'h33C: dout <= 8'b00111111; //  828 :  63 - 0x3f
      12'h33D: dout <= 8'b00000011; //  829 :   3 - 0x3
      12'h33E: dout <= 8'b00000000; //  830 :   0 - 0x0
      12'h33F: dout <= 8'b00000000; //  831 :   0 - 0x0
      12'h340: dout <= 8'b11111111; //  832 : 255 - 0xff -- Sprite 0x68
      12'h341: dout <= 8'b00000000; //  833 :   0 - 0x0
      12'h342: dout <= 8'b11001100; //  834 : 204 - 0xcc
      12'h343: dout <= 8'b00110011; //  835 :  51 - 0x33
      12'h344: dout <= 8'b11111111; //  836 : 255 - 0xff
      12'h345: dout <= 8'b11111111; //  837 : 255 - 0xff
      12'h346: dout <= 8'b00000000; //  838 :   0 - 0x0
      12'h347: dout <= 8'b00000000; //  839 :   0 - 0x0
      12'h348: dout <= 8'b11111110; //  840 : 254 - 0xfe -- Sprite 0x69
      12'h349: dout <= 8'b00000001; //  841 :   1 - 0x1
      12'h34A: dout <= 8'b11001101; //  842 : 205 - 0xcd
      12'h34B: dout <= 8'b00111110; //  843 :  62 - 0x3e
      12'h34C: dout <= 8'b11111100; //  844 : 252 - 0xfc
      12'h34D: dout <= 8'b11000000; //  845 : 192 - 0xc0
      12'h34E: dout <= 8'b00000000; //  846 :   0 - 0x0
      12'h34F: dout <= 8'b00000000; //  847 :   0 - 0x0
      12'h350: dout <= 8'b00000000; //  848 :   0 - 0x0 -- Sprite 0x6a
      12'h351: dout <= 8'b00000000; //  849 :   0 - 0x0
      12'h352: dout <= 8'b00000000; //  850 :   0 - 0x0
      12'h353: dout <= 8'b00000000; //  851 :   0 - 0x0
      12'h354: dout <= 8'b00000000; //  852 :   0 - 0x0
      12'h355: dout <= 8'b00000000; //  853 :   0 - 0x0
      12'h356: dout <= 8'b00000000; //  854 :   0 - 0x0
      12'h357: dout <= 8'b00000000; //  855 :   0 - 0x0
      12'h358: dout <= 8'b01111111; //  856 : 127 - 0x7f -- Sprite 0x6b
      12'h359: dout <= 8'b11111111; //  857 : 255 - 0xff
      12'h35A: dout <= 8'b11111111; //  858 : 255 - 0xff
      12'h35B: dout <= 8'b11111111; //  859 : 255 - 0xff
      12'h35C: dout <= 8'b01111111; //  860 : 127 - 0x7f
      12'h35D: dout <= 8'b00110000; //  861 :  48 - 0x30
      12'h35E: dout <= 8'b00001111; //  862 :  15 - 0xf
      12'h35F: dout <= 8'b00000000; //  863 :   0 - 0x0
      12'h360: dout <= 8'b11111111; //  864 : 255 - 0xff -- Sprite 0x6c
      12'h361: dout <= 8'b11111111; //  865 : 255 - 0xff
      12'h362: dout <= 8'b11111111; //  866 : 255 - 0xff
      12'h363: dout <= 8'b11111111; //  867 : 255 - 0xff
      12'h364: dout <= 8'b11111111; //  868 : 255 - 0xff
      12'h365: dout <= 8'b11111110; //  869 : 254 - 0xfe
      12'h366: dout <= 8'b00000001; //  870 :   1 - 0x1
      12'h367: dout <= 8'b11111110; //  871 : 254 - 0xfe
      12'h368: dout <= 8'b00000000; //  872 :   0 - 0x0 -- Sprite 0x6d
      12'h369: dout <= 8'b00000000; //  873 :   0 - 0x0
      12'h36A: dout <= 8'b00000000; //  874 :   0 - 0x0
      12'h36B: dout <= 8'b00000000; //  875 :   0 - 0x0
      12'h36C: dout <= 8'b00000000; //  876 :   0 - 0x0
      12'h36D: dout <= 8'b00000000; //  877 :   0 - 0x0
      12'h36E: dout <= 8'b00000000; //  878 :   0 - 0x0
      12'h36F: dout <= 8'b00000000; //  879 :   0 - 0x0
      12'h370: dout <= 8'b00000000; //  880 :   0 - 0x0 -- Sprite 0x6e
      12'h371: dout <= 8'b00000000; //  881 :   0 - 0x0
      12'h372: dout <= 8'b00000000; //  882 :   0 - 0x0
      12'h373: dout <= 8'b00000000; //  883 :   0 - 0x0
      12'h374: dout <= 8'b00000000; //  884 :   0 - 0x0
      12'h375: dout <= 8'b00000000; //  885 :   0 - 0x0
      12'h376: dout <= 8'b00000000; //  886 :   0 - 0x0
      12'h377: dout <= 8'b00000000; //  887 :   0 - 0x0
      12'h378: dout <= 8'b11111100; //  888 : 252 - 0xfc -- Sprite 0x6f
      12'h379: dout <= 8'b11111110; //  889 : 254 - 0xfe
      12'h37A: dout <= 8'b11111111; //  890 : 255 - 0xff
      12'h37B: dout <= 8'b11111111; //  891 : 255 - 0xff
      12'h37C: dout <= 8'b11110010; //  892 : 242 - 0xf2
      12'h37D: dout <= 8'b00001100; //  893 :  12 - 0xc
      12'h37E: dout <= 8'b11110000; //  894 : 240 - 0xf0
      12'h37F: dout <= 8'b00000000; //  895 :   0 - 0x0
      12'h380: dout <= 8'b01111111; //  896 : 127 - 0x7f -- Sprite 0x70
      12'h381: dout <= 8'b11000000; //  897 : 192 - 0xc0
      12'h382: dout <= 8'b10000000; //  898 : 128 - 0x80
      12'h383: dout <= 8'b10000000; //  899 : 128 - 0x80
      12'h384: dout <= 8'b11100011; //  900 : 227 - 0xe3
      12'h385: dout <= 8'b11111111; //  901 : 255 - 0xff
      12'h386: dout <= 8'b11111111; //  902 : 255 - 0xff
      12'h387: dout <= 8'b11111111; //  903 : 255 - 0xff
      12'h388: dout <= 8'b11111111; //  904 : 255 - 0xff -- Sprite 0x71
      12'h389: dout <= 8'b00000000; //  905 :   0 - 0x0
      12'h38A: dout <= 8'b00000000; //  906 :   0 - 0x0
      12'h38B: dout <= 8'b00000000; //  907 :   0 - 0x0
      12'h38C: dout <= 8'b00000000; //  908 :   0 - 0x0
      12'h38D: dout <= 8'b11000011; //  909 : 195 - 0xc3
      12'h38E: dout <= 8'b11111111; //  910 : 255 - 0xff
      12'h38F: dout <= 8'b11111111; //  911 : 255 - 0xff
      12'h390: dout <= 8'b11111110; //  912 : 254 - 0xfe -- Sprite 0x72
      12'h391: dout <= 8'b00000011; //  913 :   3 - 0x3
      12'h392: dout <= 8'b00000001; //  914 :   1 - 0x1
      12'h393: dout <= 8'b00000001; //  915 :   1 - 0x1
      12'h394: dout <= 8'b11000111; //  916 : 199 - 0xc7
      12'h395: dout <= 8'b11111111; //  917 : 255 - 0xff
      12'h396: dout <= 8'b11111111; //  918 : 255 - 0xff
      12'h397: dout <= 8'b11111111; //  919 : 255 - 0xff
      12'h398: dout <= 8'b11111111; //  920 : 255 - 0xff -- Sprite 0x73
      12'h399: dout <= 8'b11111111; //  921 : 255 - 0xff
      12'h39A: dout <= 8'b11111111; //  922 : 255 - 0xff
      12'h39B: dout <= 8'b11111111; //  923 : 255 - 0xff
      12'h39C: dout <= 8'b11111111; //  924 : 255 - 0xff
      12'h39D: dout <= 8'b11111111; //  925 : 255 - 0xff
      12'h39E: dout <= 8'b11111111; //  926 : 255 - 0xff
      12'h39F: dout <= 8'b11111111; //  927 : 255 - 0xff
      12'h3A0: dout <= 8'b10111001; //  928 : 185 - 0xb9 -- Sprite 0x74
      12'h3A1: dout <= 8'b10010100; //  929 : 148 - 0x94
      12'h3A2: dout <= 8'b10001110; //  930 : 142 - 0x8e
      12'h3A3: dout <= 8'b11000101; //  931 : 197 - 0xc5
      12'h3A4: dout <= 8'b10010010; //  932 : 146 - 0x92
      12'h3A5: dout <= 8'b11000111; //  933 : 199 - 0xc7
      12'h3A6: dout <= 8'b11100010; //  934 : 226 - 0xe2
      12'h3A7: dout <= 8'b01111111; //  935 : 127 - 0x7f
      12'h3A8: dout <= 8'b10111001; //  936 : 185 - 0xb9 -- Sprite 0x75
      12'h3A9: dout <= 8'b00010100; //  937 :  20 - 0x14
      12'h3AA: dout <= 8'b10001110; //  938 : 142 - 0x8e
      12'h3AB: dout <= 8'b11000101; //  939 : 197 - 0xc5
      12'h3AC: dout <= 8'b10010010; //  940 : 146 - 0x92
      12'h3AD: dout <= 8'b01000111; //  941 :  71 - 0x47
      12'h3AE: dout <= 8'b11100010; //  942 : 226 - 0xe2
      12'h3AF: dout <= 8'b11111111; //  943 : 255 - 0xff
      12'h3B0: dout <= 8'b10111001; //  944 : 185 - 0xb9 -- Sprite 0x76
      12'h3B1: dout <= 8'b00010101; //  945 :  21 - 0x15
      12'h3B2: dout <= 8'b10001111; //  946 : 143 - 0x8f
      12'h3B3: dout <= 8'b11000101; //  947 : 197 - 0xc5
      12'h3B4: dout <= 8'b10010011; //  948 : 147 - 0x93
      12'h3B5: dout <= 8'b01000111; //  949 :  71 - 0x47
      12'h3B6: dout <= 8'b11100011; //  950 : 227 - 0xe3
      12'h3B7: dout <= 8'b11111110; //  951 : 254 - 0xfe
      12'h3B8: dout <= 8'b11111111; //  952 : 255 - 0xff -- Sprite 0x77
      12'h3B9: dout <= 8'b11111111; //  953 : 255 - 0xff
      12'h3BA: dout <= 8'b11111111; //  954 : 255 - 0xff
      12'h3BB: dout <= 8'b11111111; //  955 : 255 - 0xff
      12'h3BC: dout <= 8'b11111111; //  956 : 255 - 0xff
      12'h3BD: dout <= 8'b11111111; //  957 : 255 - 0xff
      12'h3BE: dout <= 8'b11111111; //  958 : 255 - 0xff
      12'h3BF: dout <= 8'b11111111; //  959 : 255 - 0xff
      12'h3C0: dout <= 8'b00000000; //  960 :   0 - 0x0 -- Sprite 0x78
      12'h3C1: dout <= 8'b00000000; //  961 :   0 - 0x0
      12'h3C2: dout <= 8'b00000000; //  962 :   0 - 0x0
      12'h3C3: dout <= 8'b00000000; //  963 :   0 - 0x0
      12'h3C4: dout <= 8'b00000000; //  964 :   0 - 0x0
      12'h3C5: dout <= 8'b00000000; //  965 :   0 - 0x0
      12'h3C6: dout <= 8'b00000000; //  966 :   0 - 0x0
      12'h3C7: dout <= 8'b00000000; //  967 :   0 - 0x0
      12'h3C8: dout <= 8'b00000000; //  968 :   0 - 0x0 -- Sprite 0x79
      12'h3C9: dout <= 8'b00000000; //  969 :   0 - 0x0
      12'h3CA: dout <= 8'b00000000; //  970 :   0 - 0x0
      12'h3CB: dout <= 8'b00000000; //  971 :   0 - 0x0
      12'h3CC: dout <= 8'b00000000; //  972 :   0 - 0x0
      12'h3CD: dout <= 8'b00000000; //  973 :   0 - 0x0
      12'h3CE: dout <= 8'b00000000; //  974 :   0 - 0x0
      12'h3CF: dout <= 8'b00000000; //  975 :   0 - 0x0
      12'h3D0: dout <= 8'b00000000; //  976 :   0 - 0x0 -- Sprite 0x7a
      12'h3D1: dout <= 8'b00000000; //  977 :   0 - 0x0
      12'h3D2: dout <= 8'b00000000; //  978 :   0 - 0x0
      12'h3D3: dout <= 8'b00000000; //  979 :   0 - 0x0
      12'h3D4: dout <= 8'b00000000; //  980 :   0 - 0x0
      12'h3D5: dout <= 8'b00000000; //  981 :   0 - 0x0
      12'h3D6: dout <= 8'b00000000; //  982 :   0 - 0x0
      12'h3D7: dout <= 8'b00000000; //  983 :   0 - 0x0
      12'h3D8: dout <= 8'b00000000; //  984 :   0 - 0x0 -- Sprite 0x7b
      12'h3D9: dout <= 8'b00000000; //  985 :   0 - 0x0
      12'h3DA: dout <= 8'b00000000; //  986 :   0 - 0x0
      12'h3DB: dout <= 8'b00000000; //  987 :   0 - 0x0
      12'h3DC: dout <= 8'b00000000; //  988 :   0 - 0x0
      12'h3DD: dout <= 8'b00000000; //  989 :   0 - 0x0
      12'h3DE: dout <= 8'b00000000; //  990 :   0 - 0x0
      12'h3DF: dout <= 8'b00000000; //  991 :   0 - 0x0
      12'h3E0: dout <= 8'b00100010; //  992 :  34 - 0x22 -- Sprite 0x7c
      12'h3E1: dout <= 8'b01010101; //  993 :  85 - 0x55
      12'h3E2: dout <= 8'b10101010; //  994 : 170 - 0xaa
      12'h3E3: dout <= 8'b00000101; //  995 :   5 - 0x5
      12'h3E4: dout <= 8'b00000100; //  996 :   4 - 0x4
      12'h3E5: dout <= 8'b00001010; //  997 :  10 - 0xa
      12'h3E6: dout <= 8'b01010000; //  998 :  80 - 0x50
      12'h3E7: dout <= 8'b00000010; //  999 :   2 - 0x2
      12'h3E8: dout <= 8'b01110011; // 1000 : 115 - 0x73 -- Sprite 0x7d
      12'h3E9: dout <= 8'b11111111; // 1001 : 255 - 0xff
      12'h3EA: dout <= 8'b11111111; // 1002 : 255 - 0xff
      12'h3EB: dout <= 8'b10111101; // 1003 : 189 - 0xbd
      12'h3EC: dout <= 8'b01101110; // 1004 : 110 - 0x6e
      12'h3ED: dout <= 8'b00001010; // 1005 :  10 - 0xa
      12'h3EE: dout <= 8'b01010000; // 1006 :  80 - 0x50
      12'h3EF: dout <= 8'b00000010; // 1007 :   2 - 0x2
      12'h3F0: dout <= 8'b00100000; // 1008 :  32 - 0x20 -- Sprite 0x7e
      12'h3F1: dout <= 8'b01010000; // 1009 :  80 - 0x50
      12'h3F2: dout <= 8'b10000100; // 1010 : 132 - 0x84
      12'h3F3: dout <= 8'b00000000; // 1011 :   0 - 0x0
      12'h3F4: dout <= 8'b00100100; // 1012 :  36 - 0x24
      12'h3F5: dout <= 8'b01011010; // 1013 :  90 - 0x5a
      12'h3F6: dout <= 8'b00010000; // 1014 :  16 - 0x10
      12'h3F7: dout <= 8'b00000000; // 1015 :   0 - 0x0
      12'h3F8: dout <= 8'b11111111; // 1016 : 255 - 0xff -- Sprite 0x7f
      12'h3F9: dout <= 8'b01010000; // 1017 :  80 - 0x50
      12'h3FA: dout <= 8'b10000100; // 1018 : 132 - 0x84
      12'h3FB: dout <= 8'b00000000; // 1019 :   0 - 0x0
      12'h3FC: dout <= 8'b00100100; // 1020 :  36 - 0x24
      12'h3FD: dout <= 8'b01011010; // 1021 :  90 - 0x5a
      12'h3FE: dout <= 8'b00010000; // 1022 :  16 - 0x10
      12'h3FF: dout <= 8'b00000000; // 1023 :   0 - 0x0
      12'h400: dout <= 8'b11111111; // 1024 : 255 - 0xff -- Sprite 0x80
      12'h401: dout <= 8'b10000000; // 1025 : 128 - 0x80
      12'h402: dout <= 8'b11001111; // 1026 : 207 - 0xcf
      12'h403: dout <= 8'b01001000; // 1027 :  72 - 0x48
      12'h404: dout <= 8'b11001111; // 1028 : 207 - 0xcf
      12'h405: dout <= 8'b10000000; // 1029 : 128 - 0x80
      12'h406: dout <= 8'b11001111; // 1030 : 207 - 0xcf
      12'h407: dout <= 8'b01001000; // 1031 :  72 - 0x48
      12'h408: dout <= 8'b11111111; // 1032 : 255 - 0xff -- Sprite 0x81
      12'h409: dout <= 8'b10000000; // 1033 : 128 - 0x80
      12'h40A: dout <= 8'b11111111; // 1034 : 255 - 0xff
      12'h40B: dout <= 8'b10000000; // 1035 : 128 - 0x80
      12'h40C: dout <= 8'b10000000; // 1036 : 128 - 0x80
      12'h40D: dout <= 8'b11011111; // 1037 : 223 - 0xdf
      12'h40E: dout <= 8'b10110000; // 1038 : 176 - 0xb0
      12'h40F: dout <= 8'b11000000; // 1039 : 192 - 0xc0
      12'h410: dout <= 8'b11111111; // 1040 : 255 - 0xff -- Sprite 0x82
      12'h411: dout <= 8'b00000001; // 1041 :   1 - 0x1
      12'h412: dout <= 8'b11110011; // 1042 : 243 - 0xf3
      12'h413: dout <= 8'b00010010; // 1043 :  18 - 0x12
      12'h414: dout <= 8'b11110011; // 1044 : 243 - 0xf3
      12'h415: dout <= 8'b00000001; // 1045 :   1 - 0x1
      12'h416: dout <= 8'b11110011; // 1046 : 243 - 0xf3
      12'h417: dout <= 8'b00010010; // 1047 :  18 - 0x12
      12'h418: dout <= 8'b11111111; // 1048 : 255 - 0xff -- Sprite 0x83
      12'h419: dout <= 8'b00000000; // 1049 :   0 - 0x0
      12'h41A: dout <= 8'b11111111; // 1050 : 255 - 0xff
      12'h41B: dout <= 8'b00000000; // 1051 :   0 - 0x0
      12'h41C: dout <= 8'b00000000; // 1052 :   0 - 0x0
      12'h41D: dout <= 8'b11111111; // 1053 : 255 - 0xff
      12'h41E: dout <= 8'b00000000; // 1054 :   0 - 0x0
      12'h41F: dout <= 8'b00000000; // 1055 :   0 - 0x0
      12'h420: dout <= 8'b11111111; // 1056 : 255 - 0xff -- Sprite 0x84
      12'h421: dout <= 8'b10000010; // 1057 : 130 - 0x82
      12'h422: dout <= 8'b00010000; // 1058 :  16 - 0x10
      12'h423: dout <= 8'b00000000; // 1059 :   0 - 0x0
      12'h424: dout <= 8'b00000000; // 1060 :   0 - 0x0
      12'h425: dout <= 8'b00010000; // 1061 :  16 - 0x10
      12'h426: dout <= 8'b01000100; // 1062 :  68 - 0x44
      12'h427: dout <= 8'b11111111; // 1063 : 255 - 0xff
      12'h428: dout <= 8'b11111111; // 1064 : 255 - 0xff -- Sprite 0x85
      12'h429: dout <= 8'b00000001; // 1065 :   1 - 0x1
      12'h42A: dout <= 8'b11111111; // 1066 : 255 - 0xff
      12'h42B: dout <= 8'b00000001; // 1067 :   1 - 0x1
      12'h42C: dout <= 8'b00000001; // 1068 :   1 - 0x1
      12'h42D: dout <= 8'b11110011; // 1069 : 243 - 0xf3
      12'h42E: dout <= 8'b00001101; // 1070 :  13 - 0xd
      12'h42F: dout <= 8'b00000011; // 1071 :   3 - 0x3
      12'h430: dout <= 8'b00000000; // 1072 :   0 - 0x0 -- Sprite 0x86
      12'h431: dout <= 8'b00000000; // 1073 :   0 - 0x0
      12'h432: dout <= 8'b00000000; // 1074 :   0 - 0x0
      12'h433: dout <= 8'b00000000; // 1075 :   0 - 0x0
      12'h434: dout <= 8'b00000000; // 1076 :   0 - 0x0
      12'h435: dout <= 8'b00000000; // 1077 :   0 - 0x0
      12'h436: dout <= 8'b00000000; // 1078 :   0 - 0x0
      12'h437: dout <= 8'b00000000; // 1079 :   0 - 0x0
      12'h438: dout <= 8'b00000000; // 1080 :   0 - 0x0 -- Sprite 0x87
      12'h439: dout <= 8'b00000000; // 1081 :   0 - 0x0
      12'h43A: dout <= 8'b00000000; // 1082 :   0 - 0x0
      12'h43B: dout <= 8'b00000000; // 1083 :   0 - 0x0
      12'h43C: dout <= 8'b00000000; // 1084 :   0 - 0x0
      12'h43D: dout <= 8'b00000000; // 1085 :   0 - 0x0
      12'h43E: dout <= 8'b00000000; // 1086 :   0 - 0x0
      12'h43F: dout <= 8'b00000000; // 1087 :   0 - 0x0
      12'h440: dout <= 8'b00000111; // 1088 :   7 - 0x7 -- Sprite 0x88
      12'h441: dout <= 8'b00011110; // 1089 :  30 - 0x1e
      12'h442: dout <= 8'b00101111; // 1090 :  47 - 0x2f
      12'h443: dout <= 8'b01010011; // 1091 :  83 - 0x53
      12'h444: dout <= 8'b01101110; // 1092 : 110 - 0x6e
      12'h445: dout <= 8'b11011011; // 1093 : 219 - 0xdb
      12'h446: dout <= 8'b11111010; // 1094 : 250 - 0xfa
      12'h447: dout <= 8'b11010101; // 1095 : 213 - 0xd5
      12'h448: dout <= 8'b10111011; // 1096 : 187 - 0xbb -- Sprite 0x89
      12'h449: dout <= 8'b11110010; // 1097 : 242 - 0xf2
      12'h44A: dout <= 8'b11011101; // 1098 : 221 - 0xdd
      12'h44B: dout <= 8'b01001111; // 1099 :  79 - 0x4f
      12'h44C: dout <= 8'b01111011; // 1100 : 123 - 0x7b
      12'h44D: dout <= 8'b00110010; // 1101 :  50 - 0x32
      12'h44E: dout <= 8'b00011111; // 1102 :  31 - 0x1f
      12'h44F: dout <= 8'b00000111; // 1103 :   7 - 0x7
      12'h450: dout <= 8'b11100000; // 1104 : 224 - 0xe0 -- Sprite 0x8a
      12'h451: dout <= 8'b11011000; // 1105 : 216 - 0xd8
      12'h452: dout <= 8'b01010100; // 1106 :  84 - 0x54
      12'h453: dout <= 8'b11101010; // 1107 : 234 - 0xea
      12'h454: dout <= 8'b10111010; // 1108 : 186 - 0xba
      12'h455: dout <= 8'b10010011; // 1109 : 147 - 0x93
      12'h456: dout <= 8'b11011111; // 1110 : 223 - 0xdf
      12'h457: dout <= 8'b10111101; // 1111 : 189 - 0xbd
      12'h458: dout <= 8'b01101011; // 1112 : 107 - 0x6b -- Sprite 0x8b
      12'h459: dout <= 8'b10011111; // 1113 : 159 - 0x9f
      12'h45A: dout <= 8'b01011101; // 1114 :  93 - 0x5d
      12'h45B: dout <= 8'b10110110; // 1115 : 182 - 0xb6
      12'h45C: dout <= 8'b11101010; // 1116 : 234 - 0xea
      12'h45D: dout <= 8'b11001100; // 1117 : 204 - 0xcc
      12'h45E: dout <= 8'b01111000; // 1118 : 120 - 0x78
      12'h45F: dout <= 8'b11100000; // 1119 : 224 - 0xe0
      12'h460: dout <= 8'b00000111; // 1120 :   7 - 0x7 -- Sprite 0x8c
      12'h461: dout <= 8'b00011000; // 1121 :  24 - 0x18
      12'h462: dout <= 8'b00100011; // 1122 :  35 - 0x23
      12'h463: dout <= 8'b01001100; // 1123 :  76 - 0x4c
      12'h464: dout <= 8'b01110000; // 1124 : 112 - 0x70
      12'h465: dout <= 8'b10100001; // 1125 : 161 - 0xa1
      12'h466: dout <= 8'b10100110; // 1126 : 166 - 0xa6
      12'h467: dout <= 8'b10101000; // 1127 : 168 - 0xa8
      12'h468: dout <= 8'b10100101; // 1128 : 165 - 0xa5 -- Sprite 0x8d
      12'h469: dout <= 8'b10100010; // 1129 : 162 - 0xa2
      12'h46A: dout <= 8'b10010000; // 1130 : 144 - 0x90
      12'h46B: dout <= 8'b01001000; // 1131 :  72 - 0x48
      12'h46C: dout <= 8'b01000111; // 1132 :  71 - 0x47
      12'h46D: dout <= 8'b00100000; // 1133 :  32 - 0x20
      12'h46E: dout <= 8'b00011001; // 1134 :  25 - 0x19
      12'h46F: dout <= 8'b00000111; // 1135 :   7 - 0x7
      12'h470: dout <= 8'b11100000; // 1136 : 224 - 0xe0 -- Sprite 0x8e
      12'h471: dout <= 8'b00011000; // 1137 :  24 - 0x18
      12'h472: dout <= 8'b00000100; // 1138 :   4 - 0x4
      12'h473: dout <= 8'b11000010; // 1139 : 194 - 0xc2
      12'h474: dout <= 8'b00110010; // 1140 :  50 - 0x32
      12'h475: dout <= 8'b00001001; // 1141 :   9 - 0x9
      12'h476: dout <= 8'b11000101; // 1142 : 197 - 0xc5
      12'h477: dout <= 8'b00100101; // 1143 :  37 - 0x25
      12'h478: dout <= 8'b10100101; // 1144 : 165 - 0xa5 -- Sprite 0x8f
      12'h479: dout <= 8'b01100101; // 1145 : 101 - 0x65
      12'h47A: dout <= 8'b01000101; // 1146 :  69 - 0x45
      12'h47B: dout <= 8'b10001010; // 1147 : 138 - 0x8a
      12'h47C: dout <= 8'b10010010; // 1148 : 146 - 0x92
      12'h47D: dout <= 8'b00100100; // 1149 :  36 - 0x24
      12'h47E: dout <= 8'b11011000; // 1150 : 216 - 0xd8
      12'h47F: dout <= 8'b11100000; // 1151 : 224 - 0xe0
      12'h480: dout <= 8'b00000000; // 1152 :   0 - 0x0 -- Sprite 0x90
      12'h481: dout <= 8'b00000000; // 1153 :   0 - 0x0
      12'h482: dout <= 8'b00100000; // 1154 :  32 - 0x20
      12'h483: dout <= 8'b00110000; // 1155 :  48 - 0x30
      12'h484: dout <= 8'b00101100; // 1156 :  44 - 0x2c
      12'h485: dout <= 8'b00100010; // 1157 :  34 - 0x22
      12'h486: dout <= 8'b00010001; // 1158 :  17 - 0x11
      12'h487: dout <= 8'b00001000; // 1159 :   8 - 0x8
      12'h488: dout <= 8'b00000100; // 1160 :   4 - 0x4 -- Sprite 0x91
      12'h489: dout <= 8'b11110010; // 1161 : 242 - 0xf2
      12'h48A: dout <= 8'b11001111; // 1162 : 207 - 0xcf
      12'h48B: dout <= 8'b00110000; // 1163 :  48 - 0x30
      12'h48C: dout <= 8'b00001100; // 1164 :  12 - 0xc
      12'h48D: dout <= 8'b11111111; // 1165 : 255 - 0xff
      12'h48E: dout <= 8'b10000000; // 1166 : 128 - 0x80
      12'h48F: dout <= 8'b11111111; // 1167 : 255 - 0xff
      12'h490: dout <= 8'b01000010; // 1168 :  66 - 0x42 -- Sprite 0x92
      12'h491: dout <= 8'b10100101; // 1169 : 165 - 0xa5
      12'h492: dout <= 8'b10100101; // 1170 : 165 - 0xa5
      12'h493: dout <= 8'b10011001; // 1171 : 153 - 0x99
      12'h494: dout <= 8'b10011001; // 1172 : 153 - 0x99
      12'h495: dout <= 8'b10011001; // 1173 : 153 - 0x99
      12'h496: dout <= 8'b00000001; // 1174 :   1 - 0x1
      12'h497: dout <= 8'b00000000; // 1175 :   0 - 0x0
      12'h498: dout <= 8'b11111111; // 1176 : 255 - 0xff -- Sprite 0x93
      12'h499: dout <= 8'b11111111; // 1177 : 255 - 0xff
      12'h49A: dout <= 8'b11111111; // 1178 : 255 - 0xff
      12'h49B: dout <= 8'b10000001; // 1179 : 129 - 0x81
      12'h49C: dout <= 8'b11111111; // 1180 : 255 - 0xff
      12'h49D: dout <= 8'b11111111; // 1181 : 255 - 0xff
      12'h49E: dout <= 8'b11111111; // 1182 : 255 - 0xff
      12'h49F: dout <= 8'b10000001; // 1183 : 129 - 0x81
      12'h4A0: dout <= 8'b00000000; // 1184 :   0 - 0x0 -- Sprite 0x94
      12'h4A1: dout <= 8'b00000000; // 1185 :   0 - 0x0
      12'h4A2: dout <= 8'b00000100; // 1186 :   4 - 0x4
      12'h4A3: dout <= 8'b00001100; // 1187 :  12 - 0xc
      12'h4A4: dout <= 8'b00110100; // 1188 :  52 - 0x34
      12'h4A5: dout <= 8'b01000100; // 1189 :  68 - 0x44
      12'h4A6: dout <= 8'b10001000; // 1190 : 136 - 0x88
      12'h4A7: dout <= 8'b00010000; // 1191 :  16 - 0x10
      12'h4A8: dout <= 8'b00100000; // 1192 :  32 - 0x20 -- Sprite 0x95
      12'h4A9: dout <= 8'b01001111; // 1193 :  79 - 0x4f
      12'h4AA: dout <= 8'b11110011; // 1194 : 243 - 0xf3
      12'h4AB: dout <= 8'b00001100; // 1195 :  12 - 0xc
      12'h4AC: dout <= 8'b00110000; // 1196 :  48 - 0x30
      12'h4AD: dout <= 8'b11111111; // 1197 : 255 - 0xff
      12'h4AE: dout <= 8'b00000001; // 1198 :   1 - 0x1
      12'h4AF: dout <= 8'b11111111; // 1199 : 255 - 0xff
      12'h4B0: dout <= 8'b01111111; // 1200 : 127 - 0x7f -- Sprite 0x96
      12'h4B1: dout <= 8'b11111111; // 1201 : 255 - 0xff
      12'h4B2: dout <= 8'b11111111; // 1202 : 255 - 0xff
      12'h4B3: dout <= 8'b11111111; // 1203 : 255 - 0xff
      12'h4B4: dout <= 8'b11111011; // 1204 : 251 - 0xfb
      12'h4B5: dout <= 8'b11111111; // 1205 : 255 - 0xff
      12'h4B6: dout <= 8'b11111111; // 1206 : 255 - 0xff
      12'h4B7: dout <= 8'b11111111; // 1207 : 255 - 0xff
      12'h4B8: dout <= 8'b11111111; // 1208 : 255 - 0xff -- Sprite 0x97
      12'h4B9: dout <= 8'b11111111; // 1209 : 255 - 0xff
      12'h4BA: dout <= 8'b11111111; // 1210 : 255 - 0xff
      12'h4BB: dout <= 8'b11111111; // 1211 : 255 - 0xff
      12'h4BC: dout <= 8'b11111111; // 1212 : 255 - 0xff
      12'h4BD: dout <= 8'b11111111; // 1213 : 255 - 0xff
      12'h4BE: dout <= 8'b11111110; // 1214 : 254 - 0xfe
      12'h4BF: dout <= 8'b11111111; // 1215 : 255 - 0xff
      12'h4C0: dout <= 8'b11111111; // 1216 : 255 - 0xff -- Sprite 0x98
      12'h4C1: dout <= 8'b10111111; // 1217 : 191 - 0xbf
      12'h4C2: dout <= 8'b11111111; // 1218 : 255 - 0xff
      12'h4C3: dout <= 8'b11111111; // 1219 : 255 - 0xff
      12'h4C4: dout <= 8'b11111011; // 1220 : 251 - 0xfb
      12'h4C5: dout <= 8'b11111111; // 1221 : 255 - 0xff
      12'h4C6: dout <= 8'b11111111; // 1222 : 255 - 0xff
      12'h4C7: dout <= 8'b11111111; // 1223 : 255 - 0xff
      12'h4C8: dout <= 8'b11111111; // 1224 : 255 - 0xff -- Sprite 0x99
      12'h4C9: dout <= 8'b11111111; // 1225 : 255 - 0xff
      12'h4CA: dout <= 8'b11111111; // 1226 : 255 - 0xff
      12'h4CB: dout <= 8'b11111111; // 1227 : 255 - 0xff
      12'h4CC: dout <= 8'b11111111; // 1228 : 255 - 0xff
      12'h4CD: dout <= 8'b11111111; // 1229 : 255 - 0xff
      12'h4CE: dout <= 8'b11111110; // 1230 : 254 - 0xfe
      12'h4CF: dout <= 8'b11111111; // 1231 : 255 - 0xff
      12'h4D0: dout <= 8'b11111110; // 1232 : 254 - 0xfe -- Sprite 0x9a
      12'h4D1: dout <= 8'b11111111; // 1233 : 255 - 0xff
      12'h4D2: dout <= 8'b11111111; // 1234 : 255 - 0xff
      12'h4D3: dout <= 8'b11111111; // 1235 : 255 - 0xff
      12'h4D4: dout <= 8'b11111011; // 1236 : 251 - 0xfb
      12'h4D5: dout <= 8'b11111111; // 1237 : 255 - 0xff
      12'h4D6: dout <= 8'b11111111; // 1238 : 255 - 0xff
      12'h4D7: dout <= 8'b11111111; // 1239 : 255 - 0xff
      12'h4D8: dout <= 8'b11111111; // 1240 : 255 - 0xff -- Sprite 0x9b
      12'h4D9: dout <= 8'b11111111; // 1241 : 255 - 0xff
      12'h4DA: dout <= 8'b11111111; // 1242 : 255 - 0xff
      12'h4DB: dout <= 8'b11111111; // 1243 : 255 - 0xff
      12'h4DC: dout <= 8'b11111111; // 1244 : 255 - 0xff
      12'h4DD: dout <= 8'b11111111; // 1245 : 255 - 0xff
      12'h4DE: dout <= 8'b11111111; // 1246 : 255 - 0xff
      12'h4DF: dout <= 8'b11111111; // 1247 : 255 - 0xff
      12'h4E0: dout <= 8'b11111111; // 1248 : 255 - 0xff -- Sprite 0x9c
      12'h4E1: dout <= 8'b11111111; // 1249 : 255 - 0xff
      12'h4E2: dout <= 8'b10100000; // 1250 : 160 - 0xa0
      12'h4E3: dout <= 8'b10010000; // 1251 : 144 - 0x90
      12'h4E4: dout <= 8'b10001000; // 1252 : 136 - 0x88
      12'h4E5: dout <= 8'b10000100; // 1253 : 132 - 0x84
      12'h4E6: dout <= 8'b01101010; // 1254 : 106 - 0x6a
      12'h4E7: dout <= 8'b00111111; // 1255 :  63 - 0x3f
      12'h4E8: dout <= 8'b11111111; // 1256 : 255 - 0xff -- Sprite 0x9d
      12'h4E9: dout <= 8'b11111111; // 1257 : 255 - 0xff
      12'h4EA: dout <= 8'b00100001; // 1258 :  33 - 0x21
      12'h4EB: dout <= 8'b00010001; // 1259 :  17 - 0x11
      12'h4EC: dout <= 8'b00001001; // 1260 :   9 - 0x9
      12'h4ED: dout <= 8'b00000101; // 1261 :   5 - 0x5
      12'h4EE: dout <= 8'b10101010; // 1262 : 170 - 0xaa
      12'h4EF: dout <= 8'b11111100; // 1263 : 252 - 0xfc
      12'h4F0: dout <= 8'b11111111; // 1264 : 255 - 0xff -- Sprite 0x9e
      12'h4F1: dout <= 8'b11111111; // 1265 : 255 - 0xff
      12'h4F2: dout <= 8'b00100000; // 1266 :  32 - 0x20
      12'h4F3: dout <= 8'b00010000; // 1267 :  16 - 0x10
      12'h4F4: dout <= 8'b00001000; // 1268 :   8 - 0x8
      12'h4F5: dout <= 8'b00000100; // 1269 :   4 - 0x4
      12'h4F6: dout <= 8'b10101010; // 1270 : 170 - 0xaa
      12'h4F7: dout <= 8'b11111111; // 1271 : 255 - 0xff
      12'h4F8: dout <= 8'b00000000; // 1272 :   0 - 0x0 -- Sprite 0x9f
      12'h4F9: dout <= 8'b00000000; // 1273 :   0 - 0x0
      12'h4FA: dout <= 8'b00000000; // 1274 :   0 - 0x0
      12'h4FB: dout <= 8'b00000000; // 1275 :   0 - 0x0
      12'h4FC: dout <= 8'b00000000; // 1276 :   0 - 0x0
      12'h4FD: dout <= 8'b00000000; // 1277 :   0 - 0x0
      12'h4FE: dout <= 8'b00000000; // 1278 :   0 - 0x0
      12'h4FF: dout <= 8'b00000000; // 1279 :   0 - 0x0
      12'h500: dout <= 8'b11111111; // 1280 : 255 - 0xff -- Sprite 0xa0
      12'h501: dout <= 8'b11010101; // 1281 : 213 - 0xd5
      12'h502: dout <= 8'b11111111; // 1282 : 255 - 0xff
      12'h503: dout <= 8'b00000010; // 1283 :   2 - 0x2
      12'h504: dout <= 8'b00000010; // 1284 :   2 - 0x2
      12'h505: dout <= 8'b00000010; // 1285 :   2 - 0x2
      12'h506: dout <= 8'b00000010; // 1286 :   2 - 0x2
      12'h507: dout <= 8'b00000010; // 1287 :   2 - 0x2
      12'h508: dout <= 8'b00000010; // 1288 :   2 - 0x2 -- Sprite 0xa1
      12'h509: dout <= 8'b00000010; // 1289 :   2 - 0x2
      12'h50A: dout <= 8'b00000010; // 1290 :   2 - 0x2
      12'h50B: dout <= 8'b00000010; // 1291 :   2 - 0x2
      12'h50C: dout <= 8'b00000010; // 1292 :   2 - 0x2
      12'h50D: dout <= 8'b00000010; // 1293 :   2 - 0x2
      12'h50E: dout <= 8'b00000010; // 1294 :   2 - 0x2
      12'h50F: dout <= 8'b00000010; // 1295 :   2 - 0x2
      12'h510: dout <= 8'b11111111; // 1296 : 255 - 0xff -- Sprite 0xa2
      12'h511: dout <= 8'b01010101; // 1297 :  85 - 0x55
      12'h512: dout <= 8'b11111111; // 1298 : 255 - 0xff
      12'h513: dout <= 8'b01000000; // 1299 :  64 - 0x40
      12'h514: dout <= 8'b01000000; // 1300 :  64 - 0x40
      12'h515: dout <= 8'b01000000; // 1301 :  64 - 0x40
      12'h516: dout <= 8'b01000000; // 1302 :  64 - 0x40
      12'h517: dout <= 8'b01000000; // 1303 :  64 - 0x40
      12'h518: dout <= 8'b01000000; // 1304 :  64 - 0x40 -- Sprite 0xa3
      12'h519: dout <= 8'b01000000; // 1305 :  64 - 0x40
      12'h51A: dout <= 8'b01000000; // 1306 :  64 - 0x40
      12'h51B: dout <= 8'b01000000; // 1307 :  64 - 0x40
      12'h51C: dout <= 8'b01000000; // 1308 :  64 - 0x40
      12'h51D: dout <= 8'b01000000; // 1309 :  64 - 0x40
      12'h51E: dout <= 8'b01000000; // 1310 :  64 - 0x40
      12'h51F: dout <= 8'b01000000; // 1311 :  64 - 0x40
      12'h520: dout <= 8'b00110001; // 1312 :  49 - 0x31 -- Sprite 0xa4
      12'h521: dout <= 8'b01001000; // 1313 :  72 - 0x48
      12'h522: dout <= 8'b01000101; // 1314 :  69 - 0x45
      12'h523: dout <= 8'b10000101; // 1315 : 133 - 0x85
      12'h524: dout <= 8'b10000011; // 1316 : 131 - 0x83
      12'h525: dout <= 8'b10000010; // 1317 : 130 - 0x82
      12'h526: dout <= 8'b01100010; // 1318 :  98 - 0x62
      12'h527: dout <= 8'b00010010; // 1319 :  18 - 0x12
      12'h528: dout <= 8'b00110010; // 1320 :  50 - 0x32 -- Sprite 0xa5
      12'h529: dout <= 8'b00100010; // 1321 :  34 - 0x22
      12'h52A: dout <= 8'b01000010; // 1322 :  66 - 0x42
      12'h52B: dout <= 8'b01000000; // 1323 :  64 - 0x40
      12'h52C: dout <= 8'b01000000; // 1324 :  64 - 0x40
      12'h52D: dout <= 8'b00100000; // 1325 :  32 - 0x20
      12'h52E: dout <= 8'b00011110; // 1326 :  30 - 0x1e
      12'h52F: dout <= 8'b00000111; // 1327 :   7 - 0x7
      12'h530: dout <= 8'b10000000; // 1328 : 128 - 0x80 -- Sprite 0xa6
      12'h531: dout <= 8'b11100000; // 1329 : 224 - 0xe0
      12'h532: dout <= 8'b00111000; // 1330 :  56 - 0x38
      12'h533: dout <= 8'b00100100; // 1331 :  36 - 0x24
      12'h534: dout <= 8'b00000100; // 1332 :   4 - 0x4
      12'h535: dout <= 8'b00001000; // 1333 :   8 - 0x8
      12'h536: dout <= 8'b00110000; // 1334 :  48 - 0x30
      12'h537: dout <= 8'b00100000; // 1335 :  32 - 0x20
      12'h538: dout <= 8'b00110000; // 1336 :  48 - 0x30 -- Sprite 0xa7
      12'h539: dout <= 8'b00001000; // 1337 :   8 - 0x8
      12'h53A: dout <= 8'b00001000; // 1338 :   8 - 0x8
      12'h53B: dout <= 8'b00110000; // 1339 :  48 - 0x30
      12'h53C: dout <= 8'b00100000; // 1340 :  32 - 0x20
      12'h53D: dout <= 8'b00100000; // 1341 :  32 - 0x20
      12'h53E: dout <= 8'b00110000; // 1342 :  48 - 0x30
      12'h53F: dout <= 8'b11110000; // 1343 : 240 - 0xf0
      12'h540: dout <= 8'b11111111; // 1344 : 255 - 0xff -- Sprite 0xa8
      12'h541: dout <= 8'b11010010; // 1345 : 210 - 0xd2
      12'h542: dout <= 8'b11110100; // 1346 : 244 - 0xf4
      12'h543: dout <= 8'b11011000; // 1347 : 216 - 0xd8
      12'h544: dout <= 8'b11111000; // 1348 : 248 - 0xf8
      12'h545: dout <= 8'b11010100; // 1349 : 212 - 0xd4
      12'h546: dout <= 8'b11110010; // 1350 : 242 - 0xf2
      12'h547: dout <= 8'b11010001; // 1351 : 209 - 0xd1
      12'h548: dout <= 8'b11110001; // 1352 : 241 - 0xf1 -- Sprite 0xa9
      12'h549: dout <= 8'b11010010; // 1353 : 210 - 0xd2
      12'h54A: dout <= 8'b11110100; // 1354 : 244 - 0xf4
      12'h54B: dout <= 8'b11011000; // 1355 : 216 - 0xd8
      12'h54C: dout <= 8'b11111000; // 1356 : 248 - 0xf8
      12'h54D: dout <= 8'b11010100; // 1357 : 212 - 0xd4
      12'h54E: dout <= 8'b11110010; // 1358 : 242 - 0xf2
      12'h54F: dout <= 8'b11111111; // 1359 : 255 - 0xff
      12'h550: dout <= 8'b11111111; // 1360 : 255 - 0xff -- Sprite 0xaa
      12'h551: dout <= 8'b01000010; // 1361 :  66 - 0x42
      12'h552: dout <= 8'b00100100; // 1362 :  36 - 0x24
      12'h553: dout <= 8'b00011000; // 1363 :  24 - 0x18
      12'h554: dout <= 8'b00011000; // 1364 :  24 - 0x18
      12'h555: dout <= 8'b00100100; // 1365 :  36 - 0x24
      12'h556: dout <= 8'b01000010; // 1366 :  66 - 0x42
      12'h557: dout <= 8'b10000001; // 1367 : 129 - 0x81
      12'h558: dout <= 8'b10000001; // 1368 : 129 - 0x81 -- Sprite 0xab
      12'h559: dout <= 8'b01000010; // 1369 :  66 - 0x42
      12'h55A: dout <= 8'b00100100; // 1370 :  36 - 0x24
      12'h55B: dout <= 8'b00011000; // 1371 :  24 - 0x18
      12'h55C: dout <= 8'b00011000; // 1372 :  24 - 0x18
      12'h55D: dout <= 8'b00100100; // 1373 :  36 - 0x24
      12'h55E: dout <= 8'b01000010; // 1374 :  66 - 0x42
      12'h55F: dout <= 8'b11111111; // 1375 : 255 - 0xff
      12'h560: dout <= 8'b11111111; // 1376 : 255 - 0xff -- Sprite 0xac
      12'h561: dout <= 8'b01001101; // 1377 :  77 - 0x4d
      12'h562: dout <= 8'b00101111; // 1378 :  47 - 0x2f
      12'h563: dout <= 8'b00011101; // 1379 :  29 - 0x1d
      12'h564: dout <= 8'b00011111; // 1380 :  31 - 0x1f
      12'h565: dout <= 8'b00101101; // 1381 :  45 - 0x2d
      12'h566: dout <= 8'b01001111; // 1382 :  79 - 0x4f
      12'h567: dout <= 8'b10001101; // 1383 : 141 - 0x8d
      12'h568: dout <= 8'b10001111; // 1384 : 143 - 0x8f -- Sprite 0xad
      12'h569: dout <= 8'b01001101; // 1385 :  77 - 0x4d
      12'h56A: dout <= 8'b00101111; // 1386 :  47 - 0x2f
      12'h56B: dout <= 8'b00011101; // 1387 :  29 - 0x1d
      12'h56C: dout <= 8'b00011111; // 1388 :  31 - 0x1f
      12'h56D: dout <= 8'b00101101; // 1389 :  45 - 0x2d
      12'h56E: dout <= 8'b01001111; // 1390 :  79 - 0x4f
      12'h56F: dout <= 8'b11111111; // 1391 : 255 - 0xff
      12'h570: dout <= 8'b00000001; // 1392 :   1 - 0x1 -- Sprite 0xae
      12'h571: dout <= 8'b00000011; // 1393 :   3 - 0x3
      12'h572: dout <= 8'b00000110; // 1394 :   6 - 0x6
      12'h573: dout <= 8'b00000111; // 1395 :   7 - 0x7
      12'h574: dout <= 8'b00000111; // 1396 :   7 - 0x7
      12'h575: dout <= 8'b00000111; // 1397 :   7 - 0x7
      12'h576: dout <= 8'b00000110; // 1398 :   6 - 0x6
      12'h577: dout <= 8'b00000111; // 1399 :   7 - 0x7
      12'h578: dout <= 8'b00000110; // 1400 :   6 - 0x6 -- Sprite 0xaf
      12'h579: dout <= 8'b00000110; // 1401 :   6 - 0x6
      12'h57A: dout <= 8'b00001110; // 1402 :  14 - 0xe
      12'h57B: dout <= 8'b00001111; // 1403 :  15 - 0xf
      12'h57C: dout <= 8'b00001110; // 1404 :  14 - 0xe
      12'h57D: dout <= 8'b00011010; // 1405 :  26 - 0x1a
      12'h57E: dout <= 8'b00011011; // 1406 :  27 - 0x1b
      12'h57F: dout <= 8'b00001111; // 1407 :  15 - 0xf
      12'h580: dout <= 8'b00000000; // 1408 :   0 - 0x0 -- Sprite 0xb0
      12'h581: dout <= 8'b11000000; // 1409 : 192 - 0xc0
      12'h582: dout <= 8'b11110000; // 1410 : 240 - 0xf0
      12'h583: dout <= 8'b10001000; // 1411 : 136 - 0x88
      12'h584: dout <= 8'b00010100; // 1412 :  20 - 0x14
      12'h585: dout <= 8'b01101000; // 1413 : 104 - 0x68
      12'h586: dout <= 8'b10101000; // 1414 : 168 - 0xa8
      12'h587: dout <= 8'b00101100; // 1415 :  44 - 0x2c
      12'h588: dout <= 8'b00000100; // 1416 :   4 - 0x4 -- Sprite 0xb1
      12'h589: dout <= 8'b00111000; // 1417 :  56 - 0x38
      12'h58A: dout <= 8'b00010000; // 1418 :  16 - 0x10
      12'h58B: dout <= 8'b10100000; // 1419 : 160 - 0xa0
      12'h58C: dout <= 8'b01100000; // 1420 :  96 - 0x60
      12'h58D: dout <= 8'b00100000; // 1421 :  32 - 0x20
      12'h58E: dout <= 8'b00010000; // 1422 :  16 - 0x10
      12'h58F: dout <= 8'b10001000; // 1423 : 136 - 0x88
      12'h590: dout <= 8'b00001111; // 1424 :  15 - 0xf -- Sprite 0xb2
      12'h591: dout <= 8'b00011011; // 1425 :  27 - 0x1b
      12'h592: dout <= 8'b00011011; // 1426 :  27 - 0x1b
      12'h593: dout <= 8'b00001110; // 1427 :  14 - 0xe
      12'h594: dout <= 8'b00000110; // 1428 :   6 - 0x6
      12'h595: dout <= 8'b00001100; // 1429 :  12 - 0xc
      12'h596: dout <= 8'b00001100; // 1430 :  12 - 0xc
      12'h597: dout <= 8'b00111111; // 1431 :  63 - 0x3f
      12'h598: dout <= 8'b01111111; // 1432 : 127 - 0x7f -- Sprite 0xb3
      12'h599: dout <= 8'b01100000; // 1433 :  96 - 0x60
      12'h59A: dout <= 8'b01100000; // 1434 :  96 - 0x60
      12'h59B: dout <= 8'b01100000; // 1435 :  96 - 0x60
      12'h59C: dout <= 8'b01100000; // 1436 :  96 - 0x60
      12'h59D: dout <= 8'b01100000; // 1437 :  96 - 0x60
      12'h59E: dout <= 8'b01101010; // 1438 : 106 - 0x6a
      12'h59F: dout <= 8'b01111111; // 1439 : 127 - 0x7f
      12'h5A0: dout <= 8'b01001000; // 1440 :  72 - 0x48 -- Sprite 0xb4
      12'h5A1: dout <= 8'b00110000; // 1441 :  48 - 0x30
      12'h5A2: dout <= 8'b00010000; // 1442 :  16 - 0x10
      12'h5A3: dout <= 8'b00010000; // 1443 :  16 - 0x10
      12'h5A4: dout <= 8'b00001000; // 1444 :   8 - 0x8
      12'h5A5: dout <= 8'b00001000; // 1445 :   8 - 0x8
      12'h5A6: dout <= 8'b00001000; // 1446 :   8 - 0x8
      12'h5A7: dout <= 8'b11111100; // 1447 : 252 - 0xfc
      12'h5A8: dout <= 8'b11111110; // 1448 : 254 - 0xfe -- Sprite 0xb5
      12'h5A9: dout <= 8'b00000110; // 1449 :   6 - 0x6
      12'h5AA: dout <= 8'b00000010; // 1450 :   2 - 0x2
      12'h5AB: dout <= 8'b00000110; // 1451 :   6 - 0x6
      12'h5AC: dout <= 8'b00000010; // 1452 :   2 - 0x2
      12'h5AD: dout <= 8'b00000110; // 1453 :   6 - 0x6
      12'h5AE: dout <= 8'b10101010; // 1454 : 170 - 0xaa
      12'h5AF: dout <= 8'b11111110; // 1455 : 254 - 0xfe
      12'h5B0: dout <= 8'b11111111; // 1456 : 255 - 0xff -- Sprite 0xb6
      12'h5B1: dout <= 8'b10000000; // 1457 : 128 - 0x80
      12'h5B2: dout <= 8'b10000000; // 1458 : 128 - 0x80
      12'h5B3: dout <= 8'b10000000; // 1459 : 128 - 0x80
      12'h5B4: dout <= 8'b10000000; // 1460 : 128 - 0x80
      12'h5B5: dout <= 8'b10000000; // 1461 : 128 - 0x80
      12'h5B6: dout <= 8'b10010101; // 1462 : 149 - 0x95
      12'h5B7: dout <= 8'b11111111; // 1463 : 255 - 0xff
      12'h5B8: dout <= 8'b11111111; // 1464 : 255 - 0xff -- Sprite 0xb7
      12'h5B9: dout <= 8'b10000100; // 1465 : 132 - 0x84
      12'h5BA: dout <= 8'b10001100; // 1466 : 140 - 0x8c
      12'h5BB: dout <= 8'b10000100; // 1467 : 132 - 0x84
      12'h5BC: dout <= 8'b10001100; // 1468 : 140 - 0x8c
      12'h5BD: dout <= 8'b10000100; // 1469 : 132 - 0x84
      12'h5BE: dout <= 8'b10101100; // 1470 : 172 - 0xac
      12'h5BF: dout <= 8'b11111111; // 1471 : 255 - 0xff
      12'h5C0: dout <= 8'b11111111; // 1472 : 255 - 0xff -- Sprite 0xb8
      12'h5C1: dout <= 8'b00100001; // 1473 :  33 - 0x21
      12'h5C2: dout <= 8'b01100001; // 1474 :  97 - 0x61
      12'h5C3: dout <= 8'b00100011; // 1475 :  35 - 0x23
      12'h5C4: dout <= 8'b01100001; // 1476 :  97 - 0x61
      12'h5C5: dout <= 8'b00100011; // 1477 :  35 - 0x23
      12'h5C6: dout <= 8'b01100101; // 1478 : 101 - 0x65
      12'h5C7: dout <= 8'b11111111; // 1479 : 255 - 0xff
      12'h5C8: dout <= 8'b11111111; // 1480 : 255 - 0xff -- Sprite 0xb9
      12'h5C9: dout <= 8'b00000001; // 1481 :   1 - 0x1
      12'h5CA: dout <= 8'b00000011; // 1482 :   3 - 0x3
      12'h5CB: dout <= 8'b00000001; // 1483 :   1 - 0x1
      12'h5CC: dout <= 8'b00000011; // 1484 :   3 - 0x3
      12'h5CD: dout <= 8'b00000001; // 1485 :   1 - 0x1
      12'h5CE: dout <= 8'b10101011; // 1486 : 171 - 0xab
      12'h5CF: dout <= 8'b11111111; // 1487 : 255 - 0xff
      12'h5D0: dout <= 8'b11111111; // 1488 : 255 - 0xff -- Sprite 0xba
      12'h5D1: dout <= 8'b11010101; // 1489 : 213 - 0xd5
      12'h5D2: dout <= 8'b10101010; // 1490 : 170 - 0xaa
      12'h5D3: dout <= 8'b11111111; // 1491 : 255 - 0xff
      12'h5D4: dout <= 8'b10000000; // 1492 : 128 - 0x80
      12'h5D5: dout <= 8'b10000000; // 1493 : 128 - 0x80
      12'h5D6: dout <= 8'b10010101; // 1494 : 149 - 0x95
      12'h5D7: dout <= 8'b11111111; // 1495 : 255 - 0xff
      12'h5D8: dout <= 8'b00000000; // 1496 :   0 - 0x0 -- Sprite 0xbb
      12'h5D9: dout <= 8'b00000000; // 1497 :   0 - 0x0
      12'h5DA: dout <= 8'b00000000; // 1498 :   0 - 0x0
      12'h5DB: dout <= 8'b00000000; // 1499 :   0 - 0x0
      12'h5DC: dout <= 8'b00000000; // 1500 :   0 - 0x0
      12'h5DD: dout <= 8'b00000000; // 1501 :   0 - 0x0
      12'h5DE: dout <= 8'b00000000; // 1502 :   0 - 0x0
      12'h5DF: dout <= 8'b00000000; // 1503 :   0 - 0x0
      12'h5E0: dout <= 8'b11111111; // 1504 : 255 - 0xff -- Sprite 0xbc
      12'h5E1: dout <= 8'b01010101; // 1505 :  85 - 0x55
      12'h5E2: dout <= 8'b10101011; // 1506 : 171 - 0xab
      12'h5E3: dout <= 8'b11111111; // 1507 : 255 - 0xff
      12'h5E4: dout <= 8'b01100001; // 1508 :  97 - 0x61
      12'h5E5: dout <= 8'b00100011; // 1509 :  35 - 0x23
      12'h5E6: dout <= 8'b01100101; // 1510 : 101 - 0x65
      12'h5E7: dout <= 8'b11111111; // 1511 : 255 - 0xff
      12'h5E8: dout <= 8'b00000000; // 1512 :   0 - 0x0 -- Sprite 0xbd
      12'h5E9: dout <= 8'b00000000; // 1513 :   0 - 0x0
      12'h5EA: dout <= 8'b00000000; // 1514 :   0 - 0x0
      12'h5EB: dout <= 8'b00000000; // 1515 :   0 - 0x0
      12'h5EC: dout <= 8'b00000000; // 1516 :   0 - 0x0
      12'h5ED: dout <= 8'b00000000; // 1517 :   0 - 0x0
      12'h5EE: dout <= 8'b00000000; // 1518 :   0 - 0x0
      12'h5EF: dout <= 8'b00000000; // 1519 :   0 - 0x0
      12'h5F0: dout <= 8'b00000000; // 1520 :   0 - 0x0 -- Sprite 0xbe
      12'h5F1: dout <= 8'b00000000; // 1521 :   0 - 0x0
      12'h5F2: dout <= 8'b00000000; // 1522 :   0 - 0x0
      12'h5F3: dout <= 8'b00000000; // 1523 :   0 - 0x0
      12'h5F4: dout <= 8'b00000000; // 1524 :   0 - 0x0
      12'h5F5: dout <= 8'b00000000; // 1525 :   0 - 0x0
      12'h5F6: dout <= 8'b00000000; // 1526 :   0 - 0x0
      12'h5F7: dout <= 8'b00000000; // 1527 :   0 - 0x0
      12'h5F8: dout <= 8'b00000000; // 1528 :   0 - 0x0 -- Sprite 0xbf
      12'h5F9: dout <= 8'b00000000; // 1529 :   0 - 0x0
      12'h5FA: dout <= 8'b00000000; // 1530 :   0 - 0x0
      12'h5FB: dout <= 8'b00000000; // 1531 :   0 - 0x0
      12'h5FC: dout <= 8'b00000000; // 1532 :   0 - 0x0
      12'h5FD: dout <= 8'b00000000; // 1533 :   0 - 0x0
      12'h5FE: dout <= 8'b00000000; // 1534 :   0 - 0x0
      12'h5FF: dout <= 8'b00000000; // 1535 :   0 - 0x0
      12'h600: dout <= 8'b00000000; // 1536 :   0 - 0x0 -- Sprite 0xc0
      12'h601: dout <= 8'b00000000; // 1537 :   0 - 0x0
      12'h602: dout <= 8'b00000000; // 1538 :   0 - 0x0
      12'h603: dout <= 8'b00000000; // 1539 :   0 - 0x0
      12'h604: dout <= 8'b00000000; // 1540 :   0 - 0x0
      12'h605: dout <= 8'b00000000; // 1541 :   0 - 0x0
      12'h606: dout <= 8'b00000000; // 1542 :   0 - 0x0
      12'h607: dout <= 8'b00000000; // 1543 :   0 - 0x0
      12'h608: dout <= 8'b00000000; // 1544 :   0 - 0x0 -- Sprite 0xc1
      12'h609: dout <= 8'b00000000; // 1545 :   0 - 0x0
      12'h60A: dout <= 8'b00000000; // 1546 :   0 - 0x0
      12'h60B: dout <= 8'b00000000; // 1547 :   0 - 0x0
      12'h60C: dout <= 8'b00000000; // 1548 :   0 - 0x0
      12'h60D: dout <= 8'b00000000; // 1549 :   0 - 0x0
      12'h60E: dout <= 8'b00000000; // 1550 :   0 - 0x0
      12'h60F: dout <= 8'b00000000; // 1551 :   0 - 0x0
      12'h610: dout <= 8'b00000000; // 1552 :   0 - 0x0 -- Sprite 0xc2
      12'h611: dout <= 8'b00000000; // 1553 :   0 - 0x0
      12'h612: dout <= 8'b00000000; // 1554 :   0 - 0x0
      12'h613: dout <= 8'b00000000; // 1555 :   0 - 0x0
      12'h614: dout <= 8'b00000000; // 1556 :   0 - 0x0
      12'h615: dout <= 8'b00000000; // 1557 :   0 - 0x0
      12'h616: dout <= 8'b00000000; // 1558 :   0 - 0x0
      12'h617: dout <= 8'b00000000; // 1559 :   0 - 0x0
      12'h618: dout <= 8'b00000000; // 1560 :   0 - 0x0 -- Sprite 0xc3
      12'h619: dout <= 8'b00000000; // 1561 :   0 - 0x0
      12'h61A: dout <= 8'b00000000; // 1562 :   0 - 0x0
      12'h61B: dout <= 8'b00000000; // 1563 :   0 - 0x0
      12'h61C: dout <= 8'b00000000; // 1564 :   0 - 0x0
      12'h61D: dout <= 8'b00000000; // 1565 :   0 - 0x0
      12'h61E: dout <= 8'b00000000; // 1566 :   0 - 0x0
      12'h61F: dout <= 8'b00000000; // 1567 :   0 - 0x0
      12'h620: dout <= 8'b00000000; // 1568 :   0 - 0x0 -- Sprite 0xc4
      12'h621: dout <= 8'b00000000; // 1569 :   0 - 0x0
      12'h622: dout <= 8'b00000000; // 1570 :   0 - 0x0
      12'h623: dout <= 8'b00000000; // 1571 :   0 - 0x0
      12'h624: dout <= 8'b00000000; // 1572 :   0 - 0x0
      12'h625: dout <= 8'b00000000; // 1573 :   0 - 0x0
      12'h626: dout <= 8'b00000000; // 1574 :   0 - 0x0
      12'h627: dout <= 8'b00000000; // 1575 :   0 - 0x0
      12'h628: dout <= 8'b00000000; // 1576 :   0 - 0x0 -- Sprite 0xc5
      12'h629: dout <= 8'b00000000; // 1577 :   0 - 0x0
      12'h62A: dout <= 8'b00000001; // 1578 :   1 - 0x1
      12'h62B: dout <= 8'b00000110; // 1579 :   6 - 0x6
      12'h62C: dout <= 8'b00001010; // 1580 :  10 - 0xa
      12'h62D: dout <= 8'b00010100; // 1581 :  20 - 0x14
      12'h62E: dout <= 8'b00010000; // 1582 :  16 - 0x10
      12'h62F: dout <= 8'b00101000; // 1583 :  40 - 0x28
      12'h630: dout <= 8'b00011111; // 1584 :  31 - 0x1f -- Sprite 0xc6
      12'h631: dout <= 8'b01100000; // 1585 :  96 - 0x60
      12'h632: dout <= 8'b10100000; // 1586 : 160 - 0xa0
      12'h633: dout <= 8'b01000000; // 1587 :  64 - 0x40
      12'h634: dout <= 8'b00000000; // 1588 :   0 - 0x0
      12'h635: dout <= 8'b00000000; // 1589 :   0 - 0x0
      12'h636: dout <= 8'b00000000; // 1590 :   0 - 0x0
      12'h637: dout <= 8'b00000000; // 1591 :   0 - 0x0
      12'h638: dout <= 8'b00110000; // 1592 :  48 - 0x30 -- Sprite 0xc7
      12'h639: dout <= 8'b01000000; // 1593 :  64 - 0x40
      12'h63A: dout <= 8'b01100000; // 1594 :  96 - 0x60
      12'h63B: dout <= 8'b11000000; // 1595 : 192 - 0xc0
      12'h63C: dout <= 8'b10000000; // 1596 : 128 - 0x80
      12'h63D: dout <= 8'b10100000; // 1597 : 160 - 0xa0
      12'h63E: dout <= 8'b11000000; // 1598 : 192 - 0xc0
      12'h63F: dout <= 8'b10000000; // 1599 : 128 - 0x80
      12'h640: dout <= 8'b11111111; // 1600 : 255 - 0xff -- Sprite 0xc8
      12'h641: dout <= 8'b00000000; // 1601 :   0 - 0x0
      12'h642: dout <= 8'b00000000; // 1602 :   0 - 0x0
      12'h643: dout <= 8'b00000000; // 1603 :   0 - 0x0
      12'h644: dout <= 8'b00000000; // 1604 :   0 - 0x0
      12'h645: dout <= 8'b00000000; // 1605 :   0 - 0x0
      12'h646: dout <= 8'b00000000; // 1606 :   0 - 0x0
      12'h647: dout <= 8'b00000000; // 1607 :   0 - 0x0
      12'h648: dout <= 8'b00010100; // 1608 :  20 - 0x14 -- Sprite 0xc9
      12'h649: dout <= 8'b00101010; // 1609 :  42 - 0x2a
      12'h64A: dout <= 8'b00010110; // 1610 :  22 - 0x16
      12'h64B: dout <= 8'b00101011; // 1611 :  43 - 0x2b
      12'h64C: dout <= 8'b00010101; // 1612 :  21 - 0x15
      12'h64D: dout <= 8'b00101011; // 1613 :  43 - 0x2b
      12'h64E: dout <= 8'b00010101; // 1614 :  21 - 0x15
      12'h64F: dout <= 8'b00101011; // 1615 :  43 - 0x2b
      12'h650: dout <= 8'b00000000; // 1616 :   0 - 0x0 -- Sprite 0xca
      12'h651: dout <= 8'b00000100; // 1617 :   4 - 0x4
      12'h652: dout <= 8'b00000100; // 1618 :   4 - 0x4
      12'h653: dout <= 8'b00000101; // 1619 :   5 - 0x5
      12'h654: dout <= 8'b00010101; // 1620 :  21 - 0x15
      12'h655: dout <= 8'b00010101; // 1621 :  21 - 0x15
      12'h656: dout <= 8'b01010101; // 1622 :  85 - 0x55
      12'h657: dout <= 8'b01010101; // 1623 :  85 - 0x55
      12'h658: dout <= 8'b00000000; // 1624 :   0 - 0x0 -- Sprite 0xcb
      12'h659: dout <= 8'b00000000; // 1625 :   0 - 0x0
      12'h65A: dout <= 8'b00010000; // 1626 :  16 - 0x10
      12'h65B: dout <= 8'b00010000; // 1627 :  16 - 0x10
      12'h65C: dout <= 8'b01010001; // 1628 :  81 - 0x51
      12'h65D: dout <= 8'b01010101; // 1629 :  85 - 0x55
      12'h65E: dout <= 8'b01010101; // 1630 :  85 - 0x55
      12'h65F: dout <= 8'b01010101; // 1631 :  85 - 0x55
      12'h660: dout <= 8'b00000000; // 1632 :   0 - 0x0 -- Sprite 0xcc
      12'h661: dout <= 8'b00000000; // 1633 :   0 - 0x0
      12'h662: dout <= 8'b00000000; // 1634 :   0 - 0x0
      12'h663: dout <= 8'b00000101; // 1635 :   5 - 0x5
      12'h664: dout <= 8'b00001111; // 1636 :  15 - 0xf
      12'h665: dout <= 8'b00000111; // 1637 :   7 - 0x7
      12'h666: dout <= 8'b00000011; // 1638 :   3 - 0x3
      12'h667: dout <= 8'b00000001; // 1639 :   1 - 0x1
      12'h668: dout <= 8'b00000000; // 1640 :   0 - 0x0 -- Sprite 0xcd
      12'h669: dout <= 8'b00000000; // 1641 :   0 - 0x0
      12'h66A: dout <= 8'b10000000; // 1642 : 128 - 0x80
      12'h66B: dout <= 8'b11010000; // 1643 : 208 - 0xd0
      12'h66C: dout <= 8'b11111000; // 1644 : 248 - 0xf8
      12'h66D: dout <= 8'b11110000; // 1645 : 240 - 0xf0
      12'h66E: dout <= 8'b11100000; // 1646 : 224 - 0xe0
      12'h66F: dout <= 8'b11000000; // 1647 : 192 - 0xc0
      12'h670: dout <= 8'b00000000; // 1648 :   0 - 0x0 -- Sprite 0xce
      12'h671: dout <= 8'b00000000; // 1649 :   0 - 0x0
      12'h672: dout <= 8'b00000000; // 1650 :   0 - 0x0
      12'h673: dout <= 8'b01111000; // 1651 : 120 - 0x78
      12'h674: dout <= 8'b11001111; // 1652 : 207 - 0xcf
      12'h675: dout <= 8'b10000000; // 1653 : 128 - 0x80
      12'h676: dout <= 8'b11001111; // 1654 : 207 - 0xcf
      12'h677: dout <= 8'b01001000; // 1655 :  72 - 0x48
      12'h678: dout <= 8'b00000000; // 1656 :   0 - 0x0 -- Sprite 0xcf
      12'h679: dout <= 8'b00000000; // 1657 :   0 - 0x0
      12'h67A: dout <= 8'b00000000; // 1658 :   0 - 0x0
      12'h67B: dout <= 8'b00011110; // 1659 :  30 - 0x1e
      12'h67C: dout <= 8'b11110011; // 1660 : 243 - 0xf3
      12'h67D: dout <= 8'b00000001; // 1661 :   1 - 0x1
      12'h67E: dout <= 8'b11110011; // 1662 : 243 - 0xf3
      12'h67F: dout <= 8'b00010010; // 1663 :  18 - 0x12
      12'h680: dout <= 8'b00000000; // 1664 :   0 - 0x0 -- Sprite 0xd0
      12'h681: dout <= 8'b00000000; // 1665 :   0 - 0x0
      12'h682: dout <= 8'b00000000; // 1666 :   0 - 0x0
      12'h683: dout <= 8'b00000000; // 1667 :   0 - 0x0
      12'h684: dout <= 8'b00000000; // 1668 :   0 - 0x0
      12'h685: dout <= 8'b00000000; // 1669 :   0 - 0x0
      12'h686: dout <= 8'b00000000; // 1670 :   0 - 0x0
      12'h687: dout <= 8'b00000000; // 1671 :   0 - 0x0
      12'h688: dout <= 8'b00000000; // 1672 :   0 - 0x0 -- Sprite 0xd1
      12'h689: dout <= 8'b00000000; // 1673 :   0 - 0x0
      12'h68A: dout <= 8'b00000000; // 1674 :   0 - 0x0
      12'h68B: dout <= 8'b00000000; // 1675 :   0 - 0x0
      12'h68C: dout <= 8'b00000000; // 1676 :   0 - 0x0
      12'h68D: dout <= 8'b00000000; // 1677 :   0 - 0x0
      12'h68E: dout <= 8'b00000000; // 1678 :   0 - 0x0
      12'h68F: dout <= 8'b00000000; // 1679 :   0 - 0x0
      12'h690: dout <= 8'b00001000; // 1680 :   8 - 0x8 -- Sprite 0xd2
      12'h691: dout <= 8'b00001100; // 1681 :  12 - 0xc
      12'h692: dout <= 8'b00001000; // 1682 :   8 - 0x8
      12'h693: dout <= 8'b00001000; // 1683 :   8 - 0x8
      12'h694: dout <= 8'b00001010; // 1684 :  10 - 0xa
      12'h695: dout <= 8'b00001000; // 1685 :   8 - 0x8
      12'h696: dout <= 8'b00001000; // 1686 :   8 - 0x8
      12'h697: dout <= 8'b00001100; // 1687 :  12 - 0xc
      12'h698: dout <= 8'b00010000; // 1688 :  16 - 0x10 -- Sprite 0xd3
      12'h699: dout <= 8'b00010000; // 1689 :  16 - 0x10
      12'h69A: dout <= 8'b00110000; // 1690 :  48 - 0x30
      12'h69B: dout <= 8'b00010000; // 1691 :  16 - 0x10
      12'h69C: dout <= 8'b01010000; // 1692 :  80 - 0x50
      12'h69D: dout <= 8'b00010000; // 1693 :  16 - 0x10
      12'h69E: dout <= 8'b00110000; // 1694 :  48 - 0x30
      12'h69F: dout <= 8'b00010000; // 1695 :  16 - 0x10
      12'h6A0: dout <= 8'b00000000; // 1696 :   0 - 0x0 -- Sprite 0xd4
      12'h6A1: dout <= 8'b00000000; // 1697 :   0 - 0x0
      12'h6A2: dout <= 8'b00000000; // 1698 :   0 - 0x0
      12'h6A3: dout <= 8'b00000000; // 1699 :   0 - 0x0
      12'h6A4: dout <= 8'b00000000; // 1700 :   0 - 0x0
      12'h6A5: dout <= 8'b00000000; // 1701 :   0 - 0x0
      12'h6A6: dout <= 8'b00000000; // 1702 :   0 - 0x0
      12'h6A7: dout <= 8'b00000000; // 1703 :   0 - 0x0
      12'h6A8: dout <= 8'b11111000; // 1704 : 248 - 0xf8 -- Sprite 0xd5
      12'h6A9: dout <= 8'b00000110; // 1705 :   6 - 0x6
      12'h6AA: dout <= 8'b00000001; // 1706 :   1 - 0x1
      12'h6AB: dout <= 8'b00000000; // 1707 :   0 - 0x0
      12'h6AC: dout <= 8'b00000000; // 1708 :   0 - 0x0
      12'h6AD: dout <= 8'b00000000; // 1709 :   0 - 0x0
      12'h6AE: dout <= 8'b00000000; // 1710 :   0 - 0x0
      12'h6AF: dout <= 8'b00000000; // 1711 :   0 - 0x0
      12'h6B0: dout <= 8'b00000000; // 1712 :   0 - 0x0 -- Sprite 0xd6
      12'h6B1: dout <= 8'b00000000; // 1713 :   0 - 0x0
      12'h6B2: dout <= 8'b10000000; // 1714 : 128 - 0x80
      12'h6B3: dout <= 8'b01100000; // 1715 :  96 - 0x60
      12'h6B4: dout <= 8'b01010000; // 1716 :  80 - 0x50
      12'h6B5: dout <= 8'b10101000; // 1717 : 168 - 0xa8
      12'h6B6: dout <= 8'b01011000; // 1718 :  88 - 0x58
      12'h6B7: dout <= 8'b00101100; // 1719 :  44 - 0x2c
      12'h6B8: dout <= 8'b10100000; // 1720 : 160 - 0xa0 -- Sprite 0xd7
      12'h6B9: dout <= 8'b11000000; // 1721 : 192 - 0xc0
      12'h6BA: dout <= 8'b10000000; // 1722 : 128 - 0x80
      12'h6BB: dout <= 8'b01010000; // 1723 :  80 - 0x50
      12'h6BC: dout <= 8'b01100000; // 1724 :  96 - 0x60
      12'h6BD: dout <= 8'b00111000; // 1725 :  56 - 0x38
      12'h6BE: dout <= 8'b00001000; // 1726 :   8 - 0x8
      12'h6BF: dout <= 8'b00000111; // 1727 :   7 - 0x7
      12'h6C0: dout <= 8'b00000000; // 1728 :   0 - 0x0 -- Sprite 0xd8
      12'h6C1: dout <= 8'b00000000; // 1729 :   0 - 0x0
      12'h6C2: dout <= 8'b00000000; // 1730 :   0 - 0x0
      12'h6C3: dout <= 8'b00000000; // 1731 :   0 - 0x0
      12'h6C4: dout <= 8'b00000000; // 1732 :   0 - 0x0
      12'h6C5: dout <= 8'b00000000; // 1733 :   0 - 0x0
      12'h6C6: dout <= 8'b00000000; // 1734 :   0 - 0x0
      12'h6C7: dout <= 8'b11111111; // 1735 : 255 - 0xff
      12'h6C8: dout <= 8'b00010101; // 1736 :  21 - 0x15 -- Sprite 0xd9
      12'h6C9: dout <= 8'b00101011; // 1737 :  43 - 0x2b
      12'h6CA: dout <= 8'b00010101; // 1738 :  21 - 0x15
      12'h6CB: dout <= 8'b00101010; // 1739 :  42 - 0x2a
      12'h6CC: dout <= 8'b01010110; // 1740 :  86 - 0x56
      12'h6CD: dout <= 8'b10101100; // 1741 : 172 - 0xac
      12'h6CE: dout <= 8'b01010000; // 1742 :  80 - 0x50
      12'h6CF: dout <= 8'b11100000; // 1743 : 224 - 0xe0
      12'h6D0: dout <= 8'b00000001; // 1744 :   1 - 0x1 -- Sprite 0xda
      12'h6D1: dout <= 8'b00001101; // 1745 :  13 - 0xd
      12'h6D2: dout <= 8'b00010011; // 1746 :  19 - 0x13
      12'h6D3: dout <= 8'b00001101; // 1747 :  13 - 0xd
      12'h6D4: dout <= 8'b00000001; // 1748 :   1 - 0x1
      12'h6D5: dout <= 8'b00000001; // 1749 :   1 - 0x1
      12'h6D6: dout <= 8'b00000001; // 1750 :   1 - 0x1
      12'h6D7: dout <= 8'b00000001; // 1751 :   1 - 0x1
      12'h6D8: dout <= 8'b11000000; // 1752 : 192 - 0xc0 -- Sprite 0xdb
      12'h6D9: dout <= 8'b01000000; // 1753 :  64 - 0x40
      12'h6DA: dout <= 8'b01000000; // 1754 :  64 - 0x40
      12'h6DB: dout <= 8'b01011000; // 1755 :  88 - 0x58
      12'h6DC: dout <= 8'b01100100; // 1756 : 100 - 0x64
      12'h6DD: dout <= 8'b01011000; // 1757 :  88 - 0x58
      12'h6DE: dout <= 8'b01000000; // 1758 :  64 - 0x40
      12'h6DF: dout <= 8'b01000000; // 1759 :  64 - 0x40
      12'h6E0: dout <= 8'b00000000; // 1760 :   0 - 0x0 -- Sprite 0xdc
      12'h6E1: dout <= 8'b00000000; // 1761 :   0 - 0x0
      12'h6E2: dout <= 8'b00000000; // 1762 :   0 - 0x0
      12'h6E3: dout <= 8'b00000110; // 1763 :   6 - 0x6
      12'h6E4: dout <= 8'b00000111; // 1764 :   7 - 0x7
      12'h6E5: dout <= 8'b00000111; // 1765 :   7 - 0x7
      12'h6E6: dout <= 8'b00000111; // 1766 :   7 - 0x7
      12'h6E7: dout <= 8'b00000011; // 1767 :   3 - 0x3
      12'h6E8: dout <= 8'b00000000; // 1768 :   0 - 0x0 -- Sprite 0xdd
      12'h6E9: dout <= 8'b00000000; // 1769 :   0 - 0x0
      12'h6EA: dout <= 8'b00000000; // 1770 :   0 - 0x0
      12'h6EB: dout <= 8'b10110000; // 1771 : 176 - 0xb0
      12'h6EC: dout <= 8'b11110000; // 1772 : 240 - 0xf0
      12'h6ED: dout <= 8'b11110000; // 1773 : 240 - 0xf0
      12'h6EE: dout <= 8'b11110000; // 1774 : 240 - 0xf0
      12'h6EF: dout <= 8'b11100000; // 1775 : 224 - 0xe0
      12'h6F0: dout <= 8'b11001111; // 1776 : 207 - 0xcf -- Sprite 0xde
      12'h6F1: dout <= 8'b10000000; // 1777 : 128 - 0x80
      12'h6F2: dout <= 8'b11001111; // 1778 : 207 - 0xcf
      12'h6F3: dout <= 8'b01001000; // 1779 :  72 - 0x48
      12'h6F4: dout <= 8'b01001000; // 1780 :  72 - 0x48
      12'h6F5: dout <= 8'b01001000; // 1781 :  72 - 0x48
      12'h6F6: dout <= 8'b01001000; // 1782 :  72 - 0x48
      12'h6F7: dout <= 8'b01001000; // 1783 :  72 - 0x48
      12'h6F8: dout <= 8'b11110011; // 1784 : 243 - 0xf3 -- Sprite 0xdf
      12'h6F9: dout <= 8'b00000001; // 1785 :   1 - 0x1
      12'h6FA: dout <= 8'b11110011; // 1786 : 243 - 0xf3
      12'h6FB: dout <= 8'b00010010; // 1787 :  18 - 0x12
      12'h6FC: dout <= 8'b00010010; // 1788 :  18 - 0x12
      12'h6FD: dout <= 8'b00010010; // 1789 :  18 - 0x12
      12'h6FE: dout <= 8'b00010010; // 1790 :  18 - 0x12
      12'h6FF: dout <= 8'b00010010; // 1791 :  18 - 0x12
      12'h700: dout <= 8'b00000000; // 1792 :   0 - 0x0 -- Sprite 0xe0
      12'h701: dout <= 8'b00000000; // 1793 :   0 - 0x0
      12'h702: dout <= 8'b00000000; // 1794 :   0 - 0x0
      12'h703: dout <= 8'b00000000; // 1795 :   0 - 0x0
      12'h704: dout <= 8'b00000000; // 1796 :   0 - 0x0
      12'h705: dout <= 8'b00000000; // 1797 :   0 - 0x0
      12'h706: dout <= 8'b00000000; // 1798 :   0 - 0x0
      12'h707: dout <= 8'b00000000; // 1799 :   0 - 0x0
      12'h708: dout <= 8'b00000000; // 1800 :   0 - 0x0 -- Sprite 0xe1
      12'h709: dout <= 8'b00000000; // 1801 :   0 - 0x0
      12'h70A: dout <= 8'b00000000; // 1802 :   0 - 0x0
      12'h70B: dout <= 8'b00000000; // 1803 :   0 - 0x0
      12'h70C: dout <= 8'b00000000; // 1804 :   0 - 0x0
      12'h70D: dout <= 8'b00000000; // 1805 :   0 - 0x0
      12'h70E: dout <= 8'b00000000; // 1806 :   0 - 0x0
      12'h70F: dout <= 8'b00000000; // 1807 :   0 - 0x0
      12'h710: dout <= 8'b00000000; // 1808 :   0 - 0x0 -- Sprite 0xe2
      12'h711: dout <= 8'b00000000; // 1809 :   0 - 0x0
      12'h712: dout <= 8'b00000000; // 1810 :   0 - 0x0
      12'h713: dout <= 8'b00000000; // 1811 :   0 - 0x0
      12'h714: dout <= 8'b00000000; // 1812 :   0 - 0x0
      12'h715: dout <= 8'b00000000; // 1813 :   0 - 0x0
      12'h716: dout <= 8'b00000000; // 1814 :   0 - 0x0
      12'h717: dout <= 8'b00000000; // 1815 :   0 - 0x0
      12'h718: dout <= 8'b00000000; // 1816 :   0 - 0x0 -- Sprite 0xe3
      12'h719: dout <= 8'b00000000; // 1817 :   0 - 0x0
      12'h71A: dout <= 8'b00000000; // 1818 :   0 - 0x0
      12'h71B: dout <= 8'b00000000; // 1819 :   0 - 0x0
      12'h71C: dout <= 8'b00000000; // 1820 :   0 - 0x0
      12'h71D: dout <= 8'b00000000; // 1821 :   0 - 0x0
      12'h71E: dout <= 8'b00000000; // 1822 :   0 - 0x0
      12'h71F: dout <= 8'b00000000; // 1823 :   0 - 0x0
      12'h720: dout <= 8'b00000000; // 1824 :   0 - 0x0 -- Sprite 0xe4
      12'h721: dout <= 8'b00000000; // 1825 :   0 - 0x0
      12'h722: dout <= 8'b00000000; // 1826 :   0 - 0x0
      12'h723: dout <= 8'b00000000; // 1827 :   0 - 0x0
      12'h724: dout <= 8'b00000000; // 1828 :   0 - 0x0
      12'h725: dout <= 8'b00000000; // 1829 :   0 - 0x0
      12'h726: dout <= 8'b00000000; // 1830 :   0 - 0x0
      12'h727: dout <= 8'b00000000; // 1831 :   0 - 0x0
      12'h728: dout <= 8'b00000000; // 1832 :   0 - 0x0 -- Sprite 0xe5
      12'h729: dout <= 8'b00000000; // 1833 :   0 - 0x0
      12'h72A: dout <= 8'b00000000; // 1834 :   0 - 0x0
      12'h72B: dout <= 8'b00000000; // 1835 :   0 - 0x0
      12'h72C: dout <= 8'b00000000; // 1836 :   0 - 0x0
      12'h72D: dout <= 8'b00000000; // 1837 :   0 - 0x0
      12'h72E: dout <= 8'b00000000; // 1838 :   0 - 0x0
      12'h72F: dout <= 8'b00000000; // 1839 :   0 - 0x0
      12'h730: dout <= 8'b00000000; // 1840 :   0 - 0x0 -- Sprite 0xe6
      12'h731: dout <= 8'b00000000; // 1841 :   0 - 0x0
      12'h732: dout <= 8'b00000000; // 1842 :   0 - 0x0
      12'h733: dout <= 8'b00000000; // 1843 :   0 - 0x0
      12'h734: dout <= 8'b00000000; // 1844 :   0 - 0x0
      12'h735: dout <= 8'b00000000; // 1845 :   0 - 0x0
      12'h736: dout <= 8'b00000000; // 1846 :   0 - 0x0
      12'h737: dout <= 8'b00000000; // 1847 :   0 - 0x0
      12'h738: dout <= 8'b00000000; // 1848 :   0 - 0x0 -- Sprite 0xe7
      12'h739: dout <= 8'b00000000; // 1849 :   0 - 0x0
      12'h73A: dout <= 8'b00000000; // 1850 :   0 - 0x0
      12'h73B: dout <= 8'b00000000; // 1851 :   0 - 0x0
      12'h73C: dout <= 8'b00000000; // 1852 :   0 - 0x0
      12'h73D: dout <= 8'b00000000; // 1853 :   0 - 0x0
      12'h73E: dout <= 8'b00000000; // 1854 :   0 - 0x0
      12'h73F: dout <= 8'b00000000; // 1855 :   0 - 0x0
      12'h740: dout <= 8'b00000000; // 1856 :   0 - 0x0 -- Sprite 0xe8
      12'h741: dout <= 8'b00000000; // 1857 :   0 - 0x0
      12'h742: dout <= 8'b00000000; // 1858 :   0 - 0x0
      12'h743: dout <= 8'b00000000; // 1859 :   0 - 0x0
      12'h744: dout <= 8'b00000000; // 1860 :   0 - 0x0
      12'h745: dout <= 8'b00000000; // 1861 :   0 - 0x0
      12'h746: dout <= 8'b00000000; // 1862 :   0 - 0x0
      12'h747: dout <= 8'b00000000; // 1863 :   0 - 0x0
      12'h748: dout <= 8'b00000000; // 1864 :   0 - 0x0 -- Sprite 0xe9
      12'h749: dout <= 8'b00000000; // 1865 :   0 - 0x0
      12'h74A: dout <= 8'b00000000; // 1866 :   0 - 0x0
      12'h74B: dout <= 8'b00000000; // 1867 :   0 - 0x0
      12'h74C: dout <= 8'b00000000; // 1868 :   0 - 0x0
      12'h74D: dout <= 8'b00000000; // 1869 :   0 - 0x0
      12'h74E: dout <= 8'b00000000; // 1870 :   0 - 0x0
      12'h74F: dout <= 8'b00000000; // 1871 :   0 - 0x0
      12'h750: dout <= 8'b00000000; // 1872 :   0 - 0x0 -- Sprite 0xea
      12'h751: dout <= 8'b00000000; // 1873 :   0 - 0x0
      12'h752: dout <= 8'b00000000; // 1874 :   0 - 0x0
      12'h753: dout <= 8'b00000000; // 1875 :   0 - 0x0
      12'h754: dout <= 8'b00000000; // 1876 :   0 - 0x0
      12'h755: dout <= 8'b00000000; // 1877 :   0 - 0x0
      12'h756: dout <= 8'b00000000; // 1878 :   0 - 0x0
      12'h757: dout <= 8'b00000000; // 1879 :   0 - 0x0
      12'h758: dout <= 8'b00000000; // 1880 :   0 - 0x0 -- Sprite 0xeb
      12'h759: dout <= 8'b00000000; // 1881 :   0 - 0x0
      12'h75A: dout <= 8'b00000000; // 1882 :   0 - 0x0
      12'h75B: dout <= 8'b00000000; // 1883 :   0 - 0x0
      12'h75C: dout <= 8'b00000000; // 1884 :   0 - 0x0
      12'h75D: dout <= 8'b00000000; // 1885 :   0 - 0x0
      12'h75E: dout <= 8'b00000000; // 1886 :   0 - 0x0
      12'h75F: dout <= 8'b00000000; // 1887 :   0 - 0x0
      12'h760: dout <= 8'b00000000; // 1888 :   0 - 0x0 -- Sprite 0xec
      12'h761: dout <= 8'b00000000; // 1889 :   0 - 0x0
      12'h762: dout <= 8'b00000000; // 1890 :   0 - 0x0
      12'h763: dout <= 8'b00000000; // 1891 :   0 - 0x0
      12'h764: dout <= 8'b00000000; // 1892 :   0 - 0x0
      12'h765: dout <= 8'b00000000; // 1893 :   0 - 0x0
      12'h766: dout <= 8'b00000000; // 1894 :   0 - 0x0
      12'h767: dout <= 8'b00000000; // 1895 :   0 - 0x0
      12'h768: dout <= 8'b00000000; // 1896 :   0 - 0x0 -- Sprite 0xed
      12'h769: dout <= 8'b00000000; // 1897 :   0 - 0x0
      12'h76A: dout <= 8'b00000000; // 1898 :   0 - 0x0
      12'h76B: dout <= 8'b00000000; // 1899 :   0 - 0x0
      12'h76C: dout <= 8'b00000000; // 1900 :   0 - 0x0
      12'h76D: dout <= 8'b00000000; // 1901 :   0 - 0x0
      12'h76E: dout <= 8'b00000000; // 1902 :   0 - 0x0
      12'h76F: dout <= 8'b00000000; // 1903 :   0 - 0x0
      12'h770: dout <= 8'b00000000; // 1904 :   0 - 0x0 -- Sprite 0xee
      12'h771: dout <= 8'b00000000; // 1905 :   0 - 0x0
      12'h772: dout <= 8'b00000000; // 1906 :   0 - 0x0
      12'h773: dout <= 8'b00000000; // 1907 :   0 - 0x0
      12'h774: dout <= 8'b00000000; // 1908 :   0 - 0x0
      12'h775: dout <= 8'b00000000; // 1909 :   0 - 0x0
      12'h776: dout <= 8'b00000000; // 1910 :   0 - 0x0
      12'h777: dout <= 8'b00000000; // 1911 :   0 - 0x0
      12'h778: dout <= 8'b00000000; // 1912 :   0 - 0x0 -- Sprite 0xef
      12'h779: dout <= 8'b00000000; // 1913 :   0 - 0x0
      12'h77A: dout <= 8'b00000000; // 1914 :   0 - 0x0
      12'h77B: dout <= 8'b00000000; // 1915 :   0 - 0x0
      12'h77C: dout <= 8'b00000000; // 1916 :   0 - 0x0
      12'h77D: dout <= 8'b00000000; // 1917 :   0 - 0x0
      12'h77E: dout <= 8'b00000000; // 1918 :   0 - 0x0
      12'h77F: dout <= 8'b00000000; // 1919 :   0 - 0x0
      12'h780: dout <= 8'b00000000; // 1920 :   0 - 0x0 -- Sprite 0xf0
      12'h781: dout <= 8'b00000000; // 1921 :   0 - 0x0
      12'h782: dout <= 8'b00000000; // 1922 :   0 - 0x0
      12'h783: dout <= 8'b00000000; // 1923 :   0 - 0x0
      12'h784: dout <= 8'b00000000; // 1924 :   0 - 0x0
      12'h785: dout <= 8'b00000000; // 1925 :   0 - 0x0
      12'h786: dout <= 8'b00000000; // 1926 :   0 - 0x0
      12'h787: dout <= 8'b00000000; // 1927 :   0 - 0x0
      12'h788: dout <= 8'b00000000; // 1928 :   0 - 0x0 -- Sprite 0xf1
      12'h789: dout <= 8'b00000000; // 1929 :   0 - 0x0
      12'h78A: dout <= 8'b00000000; // 1930 :   0 - 0x0
      12'h78B: dout <= 8'b00000000; // 1931 :   0 - 0x0
      12'h78C: dout <= 8'b00000000; // 1932 :   0 - 0x0
      12'h78D: dout <= 8'b00000000; // 1933 :   0 - 0x0
      12'h78E: dout <= 8'b00000000; // 1934 :   0 - 0x0
      12'h78F: dout <= 8'b00000000; // 1935 :   0 - 0x0
      12'h790: dout <= 8'b00000000; // 1936 :   0 - 0x0 -- Sprite 0xf2
      12'h791: dout <= 8'b00000000; // 1937 :   0 - 0x0
      12'h792: dout <= 8'b00000000; // 1938 :   0 - 0x0
      12'h793: dout <= 8'b00000000; // 1939 :   0 - 0x0
      12'h794: dout <= 8'b00000000; // 1940 :   0 - 0x0
      12'h795: dout <= 8'b00000000; // 1941 :   0 - 0x0
      12'h796: dout <= 8'b00000000; // 1942 :   0 - 0x0
      12'h797: dout <= 8'b00000000; // 1943 :   0 - 0x0
      12'h798: dout <= 8'b00000000; // 1944 :   0 - 0x0 -- Sprite 0xf3
      12'h799: dout <= 8'b00000000; // 1945 :   0 - 0x0
      12'h79A: dout <= 8'b00000000; // 1946 :   0 - 0x0
      12'h79B: dout <= 8'b00000000; // 1947 :   0 - 0x0
      12'h79C: dout <= 8'b00000000; // 1948 :   0 - 0x0
      12'h79D: dout <= 8'b00000000; // 1949 :   0 - 0x0
      12'h79E: dout <= 8'b00000000; // 1950 :   0 - 0x0
      12'h79F: dout <= 8'b00000000; // 1951 :   0 - 0x0
      12'h7A0: dout <= 8'b00000000; // 1952 :   0 - 0x0 -- Sprite 0xf4
      12'h7A1: dout <= 8'b00000000; // 1953 :   0 - 0x0
      12'h7A2: dout <= 8'b00000000; // 1954 :   0 - 0x0
      12'h7A3: dout <= 8'b00000000; // 1955 :   0 - 0x0
      12'h7A4: dout <= 8'b00000000; // 1956 :   0 - 0x0
      12'h7A5: dout <= 8'b00000000; // 1957 :   0 - 0x0
      12'h7A6: dout <= 8'b00000000; // 1958 :   0 - 0x0
      12'h7A7: dout <= 8'b00000000; // 1959 :   0 - 0x0
      12'h7A8: dout <= 8'b00000000; // 1960 :   0 - 0x0 -- Sprite 0xf5
      12'h7A9: dout <= 8'b00000000; // 1961 :   0 - 0x0
      12'h7AA: dout <= 8'b00000000; // 1962 :   0 - 0x0
      12'h7AB: dout <= 8'b00000000; // 1963 :   0 - 0x0
      12'h7AC: dout <= 8'b00000000; // 1964 :   0 - 0x0
      12'h7AD: dout <= 8'b00000000; // 1965 :   0 - 0x0
      12'h7AE: dout <= 8'b00000000; // 1966 :   0 - 0x0
      12'h7AF: dout <= 8'b00000000; // 1967 :   0 - 0x0
      12'h7B0: dout <= 8'b00000000; // 1968 :   0 - 0x0 -- Sprite 0xf6
      12'h7B1: dout <= 8'b00000000; // 1969 :   0 - 0x0
      12'h7B2: dout <= 8'b00000000; // 1970 :   0 - 0x0
      12'h7B3: dout <= 8'b00000000; // 1971 :   0 - 0x0
      12'h7B4: dout <= 8'b00000000; // 1972 :   0 - 0x0
      12'h7B5: dout <= 8'b00000000; // 1973 :   0 - 0x0
      12'h7B6: dout <= 8'b00000000; // 1974 :   0 - 0x0
      12'h7B7: dout <= 8'b00000000; // 1975 :   0 - 0x0
      12'h7B8: dout <= 8'b00000000; // 1976 :   0 - 0x0 -- Sprite 0xf7
      12'h7B9: dout <= 8'b00000000; // 1977 :   0 - 0x0
      12'h7BA: dout <= 8'b00000000; // 1978 :   0 - 0x0
      12'h7BB: dout <= 8'b00000000; // 1979 :   0 - 0x0
      12'h7BC: dout <= 8'b00000000; // 1980 :   0 - 0x0
      12'h7BD: dout <= 8'b00000000; // 1981 :   0 - 0x0
      12'h7BE: dout <= 8'b00000000; // 1982 :   0 - 0x0
      12'h7BF: dout <= 8'b00000000; // 1983 :   0 - 0x0
      12'h7C0: dout <= 8'b00000000; // 1984 :   0 - 0x0 -- Sprite 0xf8
      12'h7C1: dout <= 8'b00000000; // 1985 :   0 - 0x0
      12'h7C2: dout <= 8'b00000000; // 1986 :   0 - 0x0
      12'h7C3: dout <= 8'b00000000; // 1987 :   0 - 0x0
      12'h7C4: dout <= 8'b00000000; // 1988 :   0 - 0x0
      12'h7C5: dout <= 8'b00000000; // 1989 :   0 - 0x0
      12'h7C6: dout <= 8'b00000000; // 1990 :   0 - 0x0
      12'h7C7: dout <= 8'b00000000; // 1991 :   0 - 0x0
      12'h7C8: dout <= 8'b00000000; // 1992 :   0 - 0x0 -- Sprite 0xf9
      12'h7C9: dout <= 8'b00000000; // 1993 :   0 - 0x0
      12'h7CA: dout <= 8'b00000000; // 1994 :   0 - 0x0
      12'h7CB: dout <= 8'b00000000; // 1995 :   0 - 0x0
      12'h7CC: dout <= 8'b00000000; // 1996 :   0 - 0x0
      12'h7CD: dout <= 8'b00000000; // 1997 :   0 - 0x0
      12'h7CE: dout <= 8'b00000000; // 1998 :   0 - 0x0
      12'h7CF: dout <= 8'b00000000; // 1999 :   0 - 0x0
      12'h7D0: dout <= 8'b00000000; // 2000 :   0 - 0x0 -- Sprite 0xfa
      12'h7D1: dout <= 8'b00000000; // 2001 :   0 - 0x0
      12'h7D2: dout <= 8'b00000000; // 2002 :   0 - 0x0
      12'h7D3: dout <= 8'b00000000; // 2003 :   0 - 0x0
      12'h7D4: dout <= 8'b00000000; // 2004 :   0 - 0x0
      12'h7D5: dout <= 8'b00000000; // 2005 :   0 - 0x0
      12'h7D6: dout <= 8'b00000000; // 2006 :   0 - 0x0
      12'h7D7: dout <= 8'b00000000; // 2007 :   0 - 0x0
      12'h7D8: dout <= 8'b00000000; // 2008 :   0 - 0x0 -- Sprite 0xfb
      12'h7D9: dout <= 8'b00000000; // 2009 :   0 - 0x0
      12'h7DA: dout <= 8'b00000000; // 2010 :   0 - 0x0
      12'h7DB: dout <= 8'b00000000; // 2011 :   0 - 0x0
      12'h7DC: dout <= 8'b00000000; // 2012 :   0 - 0x0
      12'h7DD: dout <= 8'b00000000; // 2013 :   0 - 0x0
      12'h7DE: dout <= 8'b00000000; // 2014 :   0 - 0x0
      12'h7DF: dout <= 8'b00000000; // 2015 :   0 - 0x0
      12'h7E0: dout <= 8'b00000000; // 2016 :   0 - 0x0 -- Sprite 0xfc
      12'h7E1: dout <= 8'b00000000; // 2017 :   0 - 0x0
      12'h7E2: dout <= 8'b10001110; // 2018 : 142 - 0x8e
      12'h7E3: dout <= 8'b10001010; // 2019 : 138 - 0x8a
      12'h7E4: dout <= 8'b10001010; // 2020 : 138 - 0x8a
      12'h7E5: dout <= 8'b10001010; // 2021 : 138 - 0x8a
      12'h7E6: dout <= 8'b10001010; // 2022 : 138 - 0x8a
      12'h7E7: dout <= 8'b11101110; // 2023 : 238 - 0xee
      12'h7E8: dout <= 8'b00000000; // 2024 :   0 - 0x0 -- Sprite 0xfd
      12'h7E9: dout <= 8'b00000000; // 2025 :   0 - 0x0
      12'h7EA: dout <= 8'b01001100; // 2026 :  76 - 0x4c
      12'h7EB: dout <= 8'b10101010; // 2027 : 170 - 0xaa
      12'h7EC: dout <= 8'b10101010; // 2028 : 170 - 0xaa
      12'h7ED: dout <= 8'b11101010; // 2029 : 234 - 0xea
      12'h7EE: dout <= 8'b10101010; // 2030 : 170 - 0xaa
      12'h7EF: dout <= 8'b10101100; // 2031 : 172 - 0xac
      12'h7F0: dout <= 8'b00000000; // 2032 :   0 - 0x0 -- Sprite 0xfe
      12'h7F1: dout <= 8'b00000000; // 2033 :   0 - 0x0
      12'h7F2: dout <= 8'b11101100; // 2034 : 236 - 0xec
      12'h7F3: dout <= 8'b01001010; // 2035 :  74 - 0x4a
      12'h7F4: dout <= 8'b01001010; // 2036 :  74 - 0x4a
      12'h7F5: dout <= 8'b01001010; // 2037 :  74 - 0x4a
      12'h7F6: dout <= 8'b01001010; // 2038 :  74 - 0x4a
      12'h7F7: dout <= 8'b11101010; // 2039 : 234 - 0xea
      12'h7F8: dout <= 8'b00000000; // 2040 :   0 - 0x0 -- Sprite 0xff
      12'h7F9: dout <= 8'b00000000; // 2041 :   0 - 0x0
      12'h7FA: dout <= 8'b01100000; // 2042 :  96 - 0x60
      12'h7FB: dout <= 8'b10001000; // 2043 : 136 - 0x88
      12'h7FC: dout <= 8'b10100000; // 2044 : 160 - 0xa0
      12'h7FD: dout <= 8'b10100000; // 2045 : 160 - 0xa0
      12'h7FE: dout <= 8'b10101000; // 2046 : 168 - 0xa8
      12'h7FF: dout <= 8'b01000000; // 2047 :  64 - 0x40
          // Background pattern Table
      12'h800: dout <= 8'b00000000; // 2048 :   0 - 0x0 -- Background 0x0
      12'h801: dout <= 8'b00001111; // 2049 :  15 - 0xf
      12'h802: dout <= 8'b00000100; // 2050 :   4 - 0x4
      12'h803: dout <= 8'b00000011; // 2051 :   3 - 0x3
      12'h804: dout <= 8'b00000011; // 2052 :   3 - 0x3
      12'h805: dout <= 8'b00000011; // 2053 :   3 - 0x3
      12'h806: dout <= 8'b00000100; // 2054 :   4 - 0x4
      12'h807: dout <= 8'b00111010; // 2055 :  58 - 0x3a
      12'h808: dout <= 8'b00000000; // 2056 :   0 - 0x0 -- Background 0x1
      12'h809: dout <= 8'b00111000; // 2057 :  56 - 0x38
      12'h80A: dout <= 8'b11000110; // 2058 : 198 - 0xc6
      12'h80B: dout <= 8'b11001011; // 2059 : 203 - 0xcb
      12'h80C: dout <= 8'b11011100; // 2060 : 220 - 0xdc
      12'h80D: dout <= 8'b00111010; // 2061 :  58 - 0x3a
      12'h80E: dout <= 8'b10011010; // 2062 : 154 - 0x9a
      12'h80F: dout <= 8'b10000001; // 2063 : 129 - 0x81
      12'h810: dout <= 8'b01000101; // 2064 :  69 - 0x45 -- Background 0x2
      12'h811: dout <= 8'b10000111; // 2065 : 135 - 0x87
      12'h812: dout <= 8'b10000011; // 2066 : 131 - 0x83
      12'h813: dout <= 8'b10000001; // 2067 : 129 - 0x81
      12'h814: dout <= 8'b10000001; // 2068 : 129 - 0x81
      12'h815: dout <= 8'b10000001; // 2069 : 129 - 0x81
      12'h816: dout <= 8'b01000001; // 2070 :  65 - 0x41
      12'h817: dout <= 8'b00100001; // 2071 :  33 - 0x21
      12'h818: dout <= 8'b01111111; // 2072 : 127 - 0x7f -- Background 0x3
      12'h819: dout <= 8'b01111110; // 2073 : 126 - 0x7e
      12'h81A: dout <= 8'b11111100; // 2074 : 252 - 0xfc
      12'h81B: dout <= 8'b00111000; // 2075 :  56 - 0x38
      12'h81C: dout <= 8'b00011000; // 2076 :  24 - 0x18
      12'h81D: dout <= 8'b10001100; // 2077 : 140 - 0x8c
      12'h81E: dout <= 8'b11000100; // 2078 : 196 - 0xc4
      12'h81F: dout <= 8'b11111100; // 2079 : 252 - 0xfc
      12'h820: dout <= 8'b00100011; // 2080 :  35 - 0x23 -- Background 0x4
      12'h821: dout <= 8'b00100011; // 2081 :  35 - 0x23
      12'h822: dout <= 8'b00100001; // 2082 :  33 - 0x21
      12'h823: dout <= 8'b00100000; // 2083 :  32 - 0x20
      12'h824: dout <= 8'b00010011; // 2084 :  19 - 0x13
      12'h825: dout <= 8'b00001100; // 2085 :  12 - 0xc
      12'h826: dout <= 8'b00000000; // 2086 :   0 - 0x0
      12'h827: dout <= 8'b00000000; // 2087 :   0 - 0x0
      12'h828: dout <= 8'b11111100; // 2088 : 252 - 0xfc -- Background 0x5
      12'h829: dout <= 8'b11111100; // 2089 : 252 - 0xfc
      12'h82A: dout <= 8'b11111100; // 2090 : 252 - 0xfc
      12'h82B: dout <= 8'b11111100; // 2091 : 252 - 0xfc
      12'h82C: dout <= 8'b10010000; // 2092 : 144 - 0x90
      12'h82D: dout <= 8'b10010000; // 2093 : 144 - 0x90
      12'h82E: dout <= 8'b10001000; // 2094 : 136 - 0x88
      12'h82F: dout <= 8'b11111000; // 2095 : 248 - 0xf8
      12'h830: dout <= 8'b00100011; // 2096 :  35 - 0x23 -- Background 0x6
      12'h831: dout <= 8'b00100011; // 2097 :  35 - 0x23
      12'h832: dout <= 8'b00100001; // 2098 :  33 - 0x21
      12'h833: dout <= 8'b00100000; // 2099 :  32 - 0x20
      12'h834: dout <= 8'b00010011; // 2100 :  19 - 0x13
      12'h835: dout <= 8'b00001101; // 2101 :  13 - 0xd
      12'h836: dout <= 8'b00000010; // 2102 :   2 - 0x2
      12'h837: dout <= 8'b00000001; // 2103 :   1 - 0x1
      12'h838: dout <= 8'b11111100; // 2104 : 252 - 0xfc -- Background 0x7
      12'h839: dout <= 8'b11111100; // 2105 : 252 - 0xfc
      12'h83A: dout <= 8'b11111100; // 2106 : 252 - 0xfc
      12'h83B: dout <= 8'b11111100; // 2107 : 252 - 0xfc
      12'h83C: dout <= 8'b10100100; // 2108 : 164 - 0xa4
      12'h83D: dout <= 8'b00100100; // 2109 :  36 - 0x24
      12'h83E: dout <= 8'b01010010; // 2110 :  82 - 0x52
      12'h83F: dout <= 8'b11101110; // 2111 : 238 - 0xee
      12'h840: dout <= 8'b00100011; // 2112 :  35 - 0x23 -- Background 0x8
      12'h841: dout <= 8'b00100011; // 2113 :  35 - 0x23
      12'h842: dout <= 8'b00100001; // 2114 :  33 - 0x21
      12'h843: dout <= 8'b00100000; // 2115 :  32 - 0x20
      12'h844: dout <= 8'b00010011; // 2116 :  19 - 0x13
      12'h845: dout <= 8'b00001101; // 2117 :  13 - 0xd
      12'h846: dout <= 8'b00000001; // 2118 :   1 - 0x1
      12'h847: dout <= 8'b00000001; // 2119 :   1 - 0x1
      12'h848: dout <= 8'b11111110; // 2120 : 254 - 0xfe -- Background 0x9
      12'h849: dout <= 8'b11111110; // 2121 : 254 - 0xfe
      12'h84A: dout <= 8'b11111110; // 2122 : 254 - 0xfe
      12'h84B: dout <= 8'b11111111; // 2123 : 255 - 0xff
      12'h84C: dout <= 8'b10010001; // 2124 : 145 - 0x91
      12'h84D: dout <= 8'b00101111; // 2125 :  47 - 0x2f
      12'h84E: dout <= 8'b01000000; // 2126 :  64 - 0x40
      12'h84F: dout <= 8'b11100000; // 2127 : 224 - 0xe0
      12'h850: dout <= 8'b00100011; // 2128 :  35 - 0x23 -- Background 0xa
      12'h851: dout <= 8'b00100011; // 2129 :  35 - 0x23
      12'h852: dout <= 8'b00100001; // 2130 :  33 - 0x21
      12'h853: dout <= 8'b00100000; // 2131 :  32 - 0x20
      12'h854: dout <= 8'b00010011; // 2132 :  19 - 0x13
      12'h855: dout <= 8'b00001110; // 2133 :  14 - 0xe
      12'h856: dout <= 8'b00000001; // 2134 :   1 - 0x1
      12'h857: dout <= 8'b00000000; // 2135 :   0 - 0x0
      12'h858: dout <= 8'b11111110; // 2136 : 254 - 0xfe -- Background 0xb
      12'h859: dout <= 8'b11111110; // 2137 : 254 - 0xfe
      12'h85A: dout <= 8'b11111110; // 2138 : 254 - 0xfe
      12'h85B: dout <= 8'b11111100; // 2139 : 252 - 0xfc
      12'h85C: dout <= 8'b00100100; // 2140 :  36 - 0x24
      12'h85D: dout <= 8'b00100010; // 2141 :  34 - 0x22
      12'h85E: dout <= 8'b11010010; // 2142 : 210 - 0xd2
      12'h85F: dout <= 8'b00001111; // 2143 :  15 - 0xf
      12'h860: dout <= 8'b01111111; // 2144 : 127 - 0x7f -- Background 0xc
      12'h861: dout <= 8'b01111110; // 2145 : 126 - 0x7e
      12'h862: dout <= 8'b11111100; // 2146 : 252 - 0xfc
      12'h863: dout <= 8'b00000010; // 2147 :   2 - 0x2
      12'h864: dout <= 8'b00000100; // 2148 :   4 - 0x4
      12'h865: dout <= 8'b11111100; // 2149 : 252 - 0xfc
      12'h866: dout <= 8'b11111100; // 2150 : 252 - 0xfc
      12'h867: dout <= 8'b11111110; // 2151 : 254 - 0xfe
      12'h868: dout <= 8'b01000101; // 2152 :  69 - 0x45 -- Background 0xd
      12'h869: dout <= 8'b10000111; // 2153 : 135 - 0x87
      12'h86A: dout <= 8'b10000011; // 2154 : 131 - 0x83
      12'h86B: dout <= 8'b10000010; // 2155 : 130 - 0x82
      12'h86C: dout <= 8'b10000010; // 2156 : 130 - 0x82
      12'h86D: dout <= 8'b10000100; // 2157 : 132 - 0x84
      12'h86E: dout <= 8'b01000100; // 2158 :  68 - 0x44
      12'h86F: dout <= 8'b00100100; // 2159 :  36 - 0x24
      12'h870: dout <= 8'b01111111; // 2160 : 127 - 0x7f -- Background 0xe
      12'h871: dout <= 8'b01111110; // 2161 : 126 - 0x7e
      12'h872: dout <= 8'b11111100; // 2162 : 252 - 0xfc
      12'h873: dout <= 8'b11111000; // 2163 : 248 - 0xf8
      12'h874: dout <= 8'b01111000; // 2164 : 120 - 0x78
      12'h875: dout <= 8'b01111100; // 2165 : 124 - 0x7c
      12'h876: dout <= 8'b11111100; // 2166 : 252 - 0xfc
      12'h877: dout <= 8'b11111110; // 2167 : 254 - 0xfe
      12'h878: dout <= 8'b00000000; // 2168 :   0 - 0x0 -- Background 0xf
      12'h879: dout <= 8'b00001111; // 2169 :  15 - 0xf
      12'h87A: dout <= 8'b00000100; // 2170 :   4 - 0x4
      12'h87B: dout <= 8'b00000011; // 2171 :   3 - 0x3
      12'h87C: dout <= 8'b00000011; // 2172 :   3 - 0x3
      12'h87D: dout <= 8'b00000011; // 2173 :   3 - 0x3
      12'h87E: dout <= 8'b00000100; // 2174 :   4 - 0x4
      12'h87F: dout <= 8'b00000010; // 2175 :   2 - 0x2
      12'h880: dout <= 8'b00000111; // 2176 :   7 - 0x7 -- Background 0x10
      12'h881: dout <= 8'b00001100; // 2177 :  12 - 0xc
      12'h882: dout <= 8'b00010000; // 2178 :  16 - 0x10
      12'h883: dout <= 8'b00010000; // 2179 :  16 - 0x10
      12'h884: dout <= 8'b00010000; // 2180 :  16 - 0x10
      12'h885: dout <= 8'b00100000; // 2181 :  32 - 0x20
      12'h886: dout <= 8'b00100000; // 2182 :  32 - 0x20
      12'h887: dout <= 8'b00100001; // 2183 :  33 - 0x21
      12'h888: dout <= 8'b11111111; // 2184 : 255 - 0xff -- Background 0x11
      12'h889: dout <= 8'b01111110; // 2185 : 126 - 0x7e
      12'h88A: dout <= 8'b01111100; // 2186 : 124 - 0x7c
      12'h88B: dout <= 8'b01111000; // 2187 : 120 - 0x78
      12'h88C: dout <= 8'b01011000; // 2188 :  88 - 0x58
      12'h88D: dout <= 8'b10001100; // 2189 : 140 - 0x8c
      12'h88E: dout <= 8'b11000100; // 2190 : 196 - 0xc4
      12'h88F: dout <= 8'b11111100; // 2191 : 252 - 0xfc
      12'h890: dout <= 8'b00100011; // 2192 :  35 - 0x23 -- Background 0x12
      12'h891: dout <= 8'b00100011; // 2193 :  35 - 0x23
      12'h892: dout <= 8'b00100001; // 2194 :  33 - 0x21
      12'h893: dout <= 8'b00100000; // 2195 :  32 - 0x20
      12'h894: dout <= 8'b00010011; // 2196 :  19 - 0x13
      12'h895: dout <= 8'b00001100; // 2197 :  12 - 0xc
      12'h896: dout <= 8'b00000000; // 2198 :   0 - 0x0
      12'h897: dout <= 8'b00000000; // 2199 :   0 - 0x0
      12'h898: dout <= 8'b00000001; // 2200 :   1 - 0x1 -- Background 0x13
      12'h899: dout <= 8'b00000001; // 2201 :   1 - 0x1
      12'h89A: dout <= 8'b00000011; // 2202 :   3 - 0x3
      12'h89B: dout <= 8'b00000100; // 2203 :   4 - 0x4
      12'h89C: dout <= 8'b00001000; // 2204 :   8 - 0x8
      12'h89D: dout <= 8'b00010000; // 2205 :  16 - 0x10
      12'h89E: dout <= 8'b00010000; // 2206 :  16 - 0x10
      12'h89F: dout <= 8'b00100000; // 2207 :  32 - 0x20
      12'h8A0: dout <= 8'b01111111; // 2208 : 127 - 0x7f -- Background 0x14
      12'h8A1: dout <= 8'b11111110; // 2209 : 254 - 0xfe
      12'h8A2: dout <= 8'b00000110; // 2210 :   6 - 0x6
      12'h8A3: dout <= 8'b00000001; // 2211 :   1 - 0x1
      12'h8A4: dout <= 8'b00000001; // 2212 :   1 - 0x1
      12'h8A5: dout <= 8'b00000001; // 2213 :   1 - 0x1
      12'h8A6: dout <= 8'b00000111; // 2214 :   7 - 0x7
      12'h8A7: dout <= 8'b11111110; // 2215 : 254 - 0xfe
      12'h8A8: dout <= 8'b00000101; // 2216 :   5 - 0x5 -- Background 0x15
      12'h8A9: dout <= 8'b00000101; // 2217 :   5 - 0x5
      12'h8AA: dout <= 8'b00000111; // 2218 :   7 - 0x7
      12'h8AB: dout <= 8'b00000100; // 2219 :   4 - 0x4
      12'h8AC: dout <= 8'b00000100; // 2220 :   4 - 0x4
      12'h8AD: dout <= 8'b00001111; // 2221 :  15 - 0xf
      12'h8AE: dout <= 8'b00110000; // 2222 :  48 - 0x30
      12'h8AF: dout <= 8'b01000000; // 2223 :  64 - 0x40
      12'h8B0: dout <= 8'b11111100; // 2224 : 252 - 0xfc -- Background 0x16
      12'h8B1: dout <= 8'b11111000; // 2225 : 248 - 0xf8
      12'h8B2: dout <= 8'b11110000; // 2226 : 240 - 0xf0
      12'h8B3: dout <= 8'b11100000; // 2227 : 224 - 0xe0
      12'h8B4: dout <= 8'b01100000; // 2228 :  96 - 0x60
      12'h8B5: dout <= 8'b11110000; // 2229 : 240 - 0xf0
      12'h8B6: dout <= 8'b00011100; // 2230 :  28 - 0x1c
      12'h8B7: dout <= 8'b00000010; // 2231 :   2 - 0x2
      12'h8B8: dout <= 8'b10000000; // 2232 : 128 - 0x80 -- Background 0x17
      12'h8B9: dout <= 8'b10000000; // 2233 : 128 - 0x80
      12'h8BA: dout <= 8'b10000000; // 2234 : 128 - 0x80
      12'h8BB: dout <= 8'b10000011; // 2235 : 131 - 0x83
      12'h8BC: dout <= 8'b01001111; // 2236 :  79 - 0x4f
      12'h8BD: dout <= 8'b00110010; // 2237 :  50 - 0x32
      12'h8BE: dout <= 8'b00000010; // 2238 :   2 - 0x2
      12'h8BF: dout <= 8'b00000011; // 2239 :   3 - 0x3
      12'h8C0: dout <= 8'b00000010; // 2240 :   2 - 0x2 -- Background 0x18
      12'h8C1: dout <= 8'b00000001; // 2241 :   1 - 0x1
      12'h8C2: dout <= 8'b00000010; // 2242 :   2 - 0x2
      12'h8C3: dout <= 8'b11111100; // 2243 : 252 - 0xfc
      12'h8C4: dout <= 8'b11000000; // 2244 : 192 - 0xc0
      12'h8C5: dout <= 8'b01000000; // 2245 :  64 - 0x40
      12'h8C6: dout <= 8'b00100000; // 2246 :  32 - 0x20
      12'h8C7: dout <= 8'b11100000; // 2247 : 224 - 0xe0
      12'h8C8: dout <= 8'b00001011; // 2248 :  11 - 0xb -- Background 0x19
      12'h8C9: dout <= 8'b00001011; // 2249 :  11 - 0xb
      12'h8CA: dout <= 8'b00001111; // 2250 :  15 - 0xf
      12'h8CB: dout <= 8'b00001001; // 2251 :   9 - 0x9
      12'h8CC: dout <= 8'b00001000; // 2252 :   8 - 0x8
      12'h8CD: dout <= 8'b00001001; // 2253 :   9 - 0x9
      12'h8CE: dout <= 8'b00001111; // 2254 :  15 - 0xf
      12'h8CF: dout <= 8'b00110000; // 2255 :  48 - 0x30
      12'h8D0: dout <= 8'b11111000; // 2256 : 248 - 0xf8 -- Background 0x1a
      12'h8D1: dout <= 8'b11110000; // 2257 : 240 - 0xf0
      12'h8D2: dout <= 8'b11100000; // 2258 : 224 - 0xe0
      12'h8D3: dout <= 8'b11000000; // 2259 : 192 - 0xc0
      12'h8D4: dout <= 8'b11000000; // 2260 : 192 - 0xc0
      12'h8D5: dout <= 8'b11000000; // 2261 : 192 - 0xc0
      12'h8D6: dout <= 8'b11111000; // 2262 : 248 - 0xf8
      12'h8D7: dout <= 8'b00011111; // 2263 :  31 - 0x1f
      12'h8D8: dout <= 8'b01000000; // 2264 :  64 - 0x40 -- Background 0x1b
      12'h8D9: dout <= 8'b01000000; // 2265 :  64 - 0x40
      12'h8DA: dout <= 8'b10000000; // 2266 : 128 - 0x80
      12'h8DB: dout <= 8'b10000000; // 2267 : 128 - 0x80
      12'h8DC: dout <= 8'b01000000; // 2268 :  64 - 0x40
      12'h8DD: dout <= 8'b00111111; // 2269 :  63 - 0x3f
      12'h8DE: dout <= 8'b00000100; // 2270 :   4 - 0x4
      12'h8DF: dout <= 8'b00000111; // 2271 :   7 - 0x7
      12'h8E0: dout <= 8'b00000000; // 2272 :   0 - 0x0 -- Background 0x1c
      12'h8E1: dout <= 8'b00000000; // 2273 :   0 - 0x0
      12'h8E2: dout <= 8'b00000000; // 2274 :   0 - 0x0
      12'h8E3: dout <= 8'b00000000; // 2275 :   0 - 0x0
      12'h8E4: dout <= 8'b00000000; // 2276 :   0 - 0x0
      12'h8E5: dout <= 8'b11111111; // 2277 : 255 - 0xff
      12'h8E6: dout <= 8'b01000000; // 2278 :  64 - 0x40
      12'h8E7: dout <= 8'b11000000; // 2279 : 192 - 0xc0
      12'h8E8: dout <= 8'b11000000; // 2280 : 192 - 0xc0 -- Background 0x1d
      12'h8E9: dout <= 8'b00100000; // 2281 :  32 - 0x20
      12'h8EA: dout <= 8'b00100000; // 2282 :  32 - 0x20
      12'h8EB: dout <= 8'b00100000; // 2283 :  32 - 0x20
      12'h8EC: dout <= 8'b01000000; // 2284 :  64 - 0x40
      12'h8ED: dout <= 8'b10000000; // 2285 : 128 - 0x80
      12'h8EE: dout <= 8'b00000000; // 2286 :   0 - 0x0
      12'h8EF: dout <= 8'b00000000; // 2287 :   0 - 0x0
      12'h8F0: dout <= 8'b01111111; // 2288 : 127 - 0x7f -- Background 0x1e
      12'h8F1: dout <= 8'b01100010; // 2289 :  98 - 0x62
      12'h8F2: dout <= 8'b11000100; // 2290 : 196 - 0xc4
      12'h8F3: dout <= 8'b00011000; // 2291 :  24 - 0x18
      12'h8F4: dout <= 8'b00111100; // 2292 :  60 - 0x3c
      12'h8F5: dout <= 8'b11111110; // 2293 : 254 - 0xfe
      12'h8F6: dout <= 8'b11111110; // 2294 : 254 - 0xfe
      12'h8F7: dout <= 8'b11111110; // 2295 : 254 - 0xfe
      12'h8F8: dout <= 8'b00000000; // 2296 :   0 - 0x0 -- Background 0x1f
      12'h8F9: dout <= 8'b00111000; // 2297 :  56 - 0x38
      12'h8FA: dout <= 8'b11000110; // 2298 : 198 - 0xc6
      12'h8FB: dout <= 8'b11001011; // 2299 : 203 - 0xcb
      12'h8FC: dout <= 8'b11011100; // 2300 : 220 - 0xdc
      12'h8FD: dout <= 8'b00111010; // 2301 :  58 - 0x3a
      12'h8FE: dout <= 8'b10011010; // 2302 : 154 - 0x9a
      12'h8FF: dout <= 8'b11100001; // 2303 : 225 - 0xe1
      12'h900: dout <= 8'b00000000; // 2304 :   0 - 0x0 -- Background 0x20
      12'h901: dout <= 8'b00011100; // 2305 :  28 - 0x1c
      12'h902: dout <= 8'b00010011; // 2306 :  19 - 0x13
      12'h903: dout <= 8'b00001000; // 2307 :   8 - 0x8
      12'h904: dout <= 8'b00010000; // 2308 :  16 - 0x10
      12'h905: dout <= 8'b00001000; // 2309 :   8 - 0x8
      12'h906: dout <= 8'b00010000; // 2310 :  16 - 0x10
      12'h907: dout <= 8'b00010000; // 2311 :  16 - 0x10
      12'h908: dout <= 8'b00000000; // 2312 :   0 - 0x0 -- Background 0x21
      12'h909: dout <= 8'b00111000; // 2313 :  56 - 0x38
      12'h90A: dout <= 8'b11001000; // 2314 : 200 - 0xc8
      12'h90B: dout <= 8'b00010000; // 2315 :  16 - 0x10
      12'h90C: dout <= 8'b00001000; // 2316 :   8 - 0x8
      12'h90D: dout <= 8'b00010000; // 2317 :  16 - 0x10
      12'h90E: dout <= 8'b00001000; // 2318 :   8 - 0x8
      12'h90F: dout <= 8'b00001000; // 2319 :   8 - 0x8
      12'h910: dout <= 8'b00001000; // 2320 :   8 - 0x8 -- Background 0x22
      12'h911: dout <= 8'b00011100; // 2321 :  28 - 0x1c
      12'h912: dout <= 8'b00100111; // 2322 :  39 - 0x27
      12'h913: dout <= 8'b00101111; // 2323 :  47 - 0x2f
      12'h914: dout <= 8'b00011111; // 2324 :  31 - 0x1f
      12'h915: dout <= 8'b00001111; // 2325 :  15 - 0xf
      12'h916: dout <= 8'b00001111; // 2326 :  15 - 0xf
      12'h917: dout <= 8'b00001111; // 2327 :  15 - 0xf
      12'h918: dout <= 8'b00010000; // 2328 :  16 - 0x10 -- Background 0x23
      12'h919: dout <= 8'b00111100; // 2329 :  60 - 0x3c
      12'h91A: dout <= 8'b11000010; // 2330 : 194 - 0xc2
      12'h91B: dout <= 8'b10000010; // 2331 : 130 - 0x82
      12'h91C: dout <= 8'b10000010; // 2332 : 130 - 0x82
      12'h91D: dout <= 8'b10000010; // 2333 : 130 - 0x82
      12'h91E: dout <= 8'b00010010; // 2334 :  18 - 0x12
      12'h91F: dout <= 8'b00011100; // 2335 :  28 - 0x1c
      12'h920: dout <= 8'b00001111; // 2336 :  15 - 0xf -- Background 0x24
      12'h921: dout <= 8'b00001110; // 2337 :  14 - 0xe
      12'h922: dout <= 8'b00010100; // 2338 :  20 - 0x14
      12'h923: dout <= 8'b00010100; // 2339 :  20 - 0x14
      12'h924: dout <= 8'b00010010; // 2340 :  18 - 0x12
      12'h925: dout <= 8'b00100101; // 2341 :  37 - 0x25
      12'h926: dout <= 8'b01000100; // 2342 :  68 - 0x44
      12'h927: dout <= 8'b00111000; // 2343 :  56 - 0x38
      12'h928: dout <= 8'b00010000; // 2344 :  16 - 0x10 -- Background 0x25
      12'h929: dout <= 8'b00010000; // 2345 :  16 - 0x10
      12'h92A: dout <= 8'b00010000; // 2346 :  16 - 0x10
      12'h92B: dout <= 8'b00101100; // 2347 :  44 - 0x2c
      12'h92C: dout <= 8'b01000100; // 2348 :  68 - 0x44
      12'h92D: dout <= 8'b11000100; // 2349 : 196 - 0xc4
      12'h92E: dout <= 8'b00111000; // 2350 :  56 - 0x38
      12'h92F: dout <= 8'b00000000; // 2351 :   0 - 0x0
      12'h930: dout <= 8'b00000000; // 2352 :   0 - 0x0 -- Background 0x26
      12'h931: dout <= 8'b00000000; // 2353 :   0 - 0x0
      12'h932: dout <= 8'b00000000; // 2354 :   0 - 0x0
      12'h933: dout <= 8'b00000000; // 2355 :   0 - 0x0
      12'h934: dout <= 8'b00000000; // 2356 :   0 - 0x0
      12'h935: dout <= 8'b00000000; // 2357 :   0 - 0x0
      12'h936: dout <= 8'b00000000; // 2358 :   0 - 0x0
      12'h937: dout <= 8'b00000000; // 2359 :   0 - 0x0
      12'h938: dout <= 8'b00000000; // 2360 :   0 - 0x0 -- Background 0x27
      12'h939: dout <= 8'b00000000; // 2361 :   0 - 0x0
      12'h93A: dout <= 8'b00000000; // 2362 :   0 - 0x0
      12'h93B: dout <= 8'b00000000; // 2363 :   0 - 0x0
      12'h93C: dout <= 8'b00000000; // 2364 :   0 - 0x0
      12'h93D: dout <= 8'b00000000; // 2365 :   0 - 0x0
      12'h93E: dout <= 8'b00000000; // 2366 :   0 - 0x0
      12'h93F: dout <= 8'b00000000; // 2367 :   0 - 0x0
      12'h940: dout <= 8'b00000000; // 2368 :   0 - 0x0 -- Background 0x28
      12'h941: dout <= 8'b00000000; // 2369 :   0 - 0x0
      12'h942: dout <= 8'b00000000; // 2370 :   0 - 0x0
      12'h943: dout <= 8'b00000000; // 2371 :   0 - 0x0
      12'h944: dout <= 8'b00000000; // 2372 :   0 - 0x0
      12'h945: dout <= 8'b00000000; // 2373 :   0 - 0x0
      12'h946: dout <= 8'b00000000; // 2374 :   0 - 0x0
      12'h947: dout <= 8'b00000000; // 2375 :   0 - 0x0
      12'h948: dout <= 8'b00100000; // 2376 :  32 - 0x20 -- Background 0x29
      12'h949: dout <= 8'b00100000; // 2377 :  32 - 0x20
      12'h94A: dout <= 8'b00100000; // 2378 :  32 - 0x20
      12'h94B: dout <= 8'b00100000; // 2379 :  32 - 0x20
      12'h94C: dout <= 8'b00010011; // 2380 :  19 - 0x13
      12'h94D: dout <= 8'b00001101; // 2381 :  13 - 0xd
      12'h94E: dout <= 8'b00000010; // 2382 :   2 - 0x2
      12'h94F: dout <= 8'b00000001; // 2383 :   1 - 0x1
      12'h950: dout <= 8'b00100000; // 2384 :  32 - 0x20 -- Background 0x2a
      12'h951: dout <= 8'b00100000; // 2385 :  32 - 0x20
      12'h952: dout <= 8'b00100000; // 2386 :  32 - 0x20
      12'h953: dout <= 8'b00100000; // 2387 :  32 - 0x20
      12'h954: dout <= 8'b00010011; // 2388 :  19 - 0x13
      12'h955: dout <= 8'b00001101; // 2389 :  13 - 0xd
      12'h956: dout <= 8'b00000001; // 2390 :   1 - 0x1
      12'h957: dout <= 8'b00000001; // 2391 :   1 - 0x1
      12'h958: dout <= 8'b00000000; // 2392 :   0 - 0x0 -- Background 0x2b
      12'h959: dout <= 8'b00000000; // 2393 :   0 - 0x0
      12'h95A: dout <= 8'b00000000; // 2394 :   0 - 0x0
      12'h95B: dout <= 8'b00000000; // 2395 :   0 - 0x0
      12'h95C: dout <= 8'b00000000; // 2396 :   0 - 0x0
      12'h95D: dout <= 8'b00000000; // 2397 :   0 - 0x0
      12'h95E: dout <= 8'b00000000; // 2398 :   0 - 0x0
      12'h95F: dout <= 8'b00000000; // 2399 :   0 - 0x0
      12'h960: dout <= 8'b00000000; // 2400 :   0 - 0x0 -- Background 0x2c
      12'h961: dout <= 8'b00000000; // 2401 :   0 - 0x0
      12'h962: dout <= 8'b00000000; // 2402 :   0 - 0x0
      12'h963: dout <= 8'b00000000; // 2403 :   0 - 0x0
      12'h964: dout <= 8'b00000000; // 2404 :   0 - 0x0
      12'h965: dout <= 8'b00000000; // 2405 :   0 - 0x0
      12'h966: dout <= 8'b00000000; // 2406 :   0 - 0x0
      12'h967: dout <= 8'b00000000; // 2407 :   0 - 0x0
      12'h968: dout <= 8'b00111100; // 2408 :  60 - 0x3c -- Background 0x2d
      12'h969: dout <= 8'b00000000; // 2409 :   0 - 0x0
      12'h96A: dout <= 8'b10000001; // 2410 : 129 - 0x81
      12'h96B: dout <= 8'b10011001; // 2411 : 153 - 0x99
      12'h96C: dout <= 8'b10011001; // 2412 : 153 - 0x99
      12'h96D: dout <= 8'b10000001; // 2413 : 129 - 0x81
      12'h96E: dout <= 8'b00000000; // 2414 :   0 - 0x0
      12'h96F: dout <= 8'b00111100; // 2415 :  60 - 0x3c
      12'h970: dout <= 8'b00000000; // 2416 :   0 - 0x0 -- Background 0x2e
      12'h971: dout <= 8'b00000000; // 2417 :   0 - 0x0
      12'h972: dout <= 8'b00000000; // 2418 :   0 - 0x0
      12'h973: dout <= 8'b00000000; // 2419 :   0 - 0x0
      12'h974: dout <= 8'b00000000; // 2420 :   0 - 0x0
      12'h975: dout <= 8'b00000000; // 2421 :   0 - 0x0
      12'h976: dout <= 8'b00000000; // 2422 :   0 - 0x0
      12'h977: dout <= 8'b00000000; // 2423 :   0 - 0x0
      12'h978: dout <= 8'b10011111; // 2424 : 159 - 0x9f -- Background 0x2f
      12'h979: dout <= 8'b10011110; // 2425 : 158 - 0x9e
      12'h97A: dout <= 8'b10011100; // 2426 : 156 - 0x9c
      12'h97B: dout <= 8'b00011000; // 2427 :  24 - 0x18
      12'h97C: dout <= 8'b00111000; // 2428 :  56 - 0x38
      12'h97D: dout <= 8'b11111100; // 2429 : 252 - 0xfc
      12'h97E: dout <= 8'b11111100; // 2430 : 252 - 0xfc
      12'h97F: dout <= 8'b11111100; // 2431 : 252 - 0xfc
      12'h980: dout <= 8'b01111111; // 2432 : 127 - 0x7f -- Background 0x30
      12'h981: dout <= 8'b01111110; // 2433 : 126 - 0x7e
      12'h982: dout <= 8'b11111100; // 2434 : 252 - 0xfc
      12'h983: dout <= 8'b00111000; // 2435 :  56 - 0x38
      12'h984: dout <= 8'b00111000; // 2436 :  56 - 0x38
      12'h985: dout <= 8'b00000100; // 2437 :   4 - 0x4
      12'h986: dout <= 8'b10000100; // 2438 : 132 - 0x84
      12'h987: dout <= 8'b11111100; // 2439 : 252 - 0xfc
      12'h988: dout <= 8'b01111111; // 2440 : 127 - 0x7f -- Background 0x31
      12'h989: dout <= 8'b01111110; // 2441 : 126 - 0x7e
      12'h98A: dout <= 8'b11111100; // 2442 : 252 - 0xfc
      12'h98B: dout <= 8'b00111000; // 2443 :  56 - 0x38
      12'h98C: dout <= 8'b00111000; // 2444 :  56 - 0x38
      12'h98D: dout <= 8'b00011100; // 2445 :  28 - 0x1c
      12'h98E: dout <= 8'b10000100; // 2446 : 132 - 0x84
      12'h98F: dout <= 8'b11000100; // 2447 : 196 - 0xc4
      12'h990: dout <= 8'b01111111; // 2448 : 127 - 0x7f -- Background 0x32
      12'h991: dout <= 8'b01111110; // 2449 : 126 - 0x7e
      12'h992: dout <= 8'b11111100; // 2450 : 252 - 0xfc
      12'h993: dout <= 8'b00111000; // 2451 :  56 - 0x38
      12'h994: dout <= 8'b00100100; // 2452 :  36 - 0x24
      12'h995: dout <= 8'b00000100; // 2453 :   4 - 0x4
      12'h996: dout <= 8'b10011100; // 2454 : 156 - 0x9c
      12'h997: dout <= 8'b11111100; // 2455 : 252 - 0xfc
      12'h998: dout <= 8'b00100011; // 2456 :  35 - 0x23 -- Background 0x33
      12'h999: dout <= 8'b00100011; // 2457 :  35 - 0x23
      12'h99A: dout <= 8'b00100001; // 2458 :  33 - 0x21
      12'h99B: dout <= 8'b00100000; // 2459 :  32 - 0x20
      12'h99C: dout <= 8'b00010011; // 2460 :  19 - 0x13
      12'h99D: dout <= 8'b00001101; // 2461 :  13 - 0xd
      12'h99E: dout <= 8'b00000001; // 2462 :   1 - 0x1
      12'h99F: dout <= 8'b00000001; // 2463 :   1 - 0x1
      12'h9A0: dout <= 8'b11111100; // 2464 : 252 - 0xfc -- Background 0x34
      12'h9A1: dout <= 8'b11111100; // 2465 : 252 - 0xfc
      12'h9A2: dout <= 8'b11111100; // 2466 : 252 - 0xfc
      12'h9A3: dout <= 8'b11111100; // 2467 : 252 - 0xfc
      12'h9A4: dout <= 8'b10100100; // 2468 : 164 - 0xa4
      12'h9A5: dout <= 8'b00100100; // 2469 :  36 - 0x24
      12'h9A6: dout <= 8'b00010010; // 2470 :  18 - 0x12
      12'h9A7: dout <= 8'b11101110; // 2471 : 238 - 0xee
      12'h9A8: dout <= 8'b00100011; // 2472 :  35 - 0x23 -- Background 0x35
      12'h9A9: dout <= 8'b00100011; // 2473 :  35 - 0x23
      12'h9AA: dout <= 8'b00100001; // 2474 :  33 - 0x21
      12'h9AB: dout <= 8'b00100000; // 2475 :  32 - 0x20
      12'h9AC: dout <= 8'b00010011; // 2476 :  19 - 0x13
      12'h9AD: dout <= 8'b00001110; // 2477 :  14 - 0xe
      12'h9AE: dout <= 8'b00000010; // 2478 :   2 - 0x2
      12'h9AF: dout <= 8'b00000001; // 2479 :   1 - 0x1
      12'h9B0: dout <= 8'b11111100; // 2480 : 252 - 0xfc -- Background 0x36
      12'h9B1: dout <= 8'b11111100; // 2481 : 252 - 0xfc
      12'h9B2: dout <= 8'b11111100; // 2482 : 252 - 0xfc
      12'h9B3: dout <= 8'b11111100; // 2483 : 252 - 0xfc
      12'h9B4: dout <= 8'b10100110; // 2484 : 166 - 0xa6
      12'h9B5: dout <= 8'b00110001; // 2485 :  49 - 0x31
      12'h9B6: dout <= 8'b01001001; // 2486 :  73 - 0x49
      12'h9B7: dout <= 8'b11000110; // 2487 : 198 - 0xc6
      12'h9B8: dout <= 8'b11111100; // 2488 : 252 - 0xfc -- Background 0x37
      12'h9B9: dout <= 8'b11111100; // 2489 : 252 - 0xfc
      12'h9BA: dout <= 8'b11111100; // 2490 : 252 - 0xfc
      12'h9BB: dout <= 8'b11111100; // 2491 : 252 - 0xfc
      12'h9BC: dout <= 8'b10100100; // 2492 : 164 - 0xa4
      12'h9BD: dout <= 8'b00100100; // 2493 :  36 - 0x24
      12'h9BE: dout <= 8'b00010010; // 2494 :  18 - 0x12
      12'h9BF: dout <= 8'b11101110; // 2495 : 238 - 0xee
      12'h9C0: dout <= 8'b00000000; // 2496 :   0 - 0x0 -- Background 0x38
      12'h9C1: dout <= 8'b00000000; // 2497 :   0 - 0x0
      12'h9C2: dout <= 8'b00000000; // 2498 :   0 - 0x0
      12'h9C3: dout <= 8'b00000000; // 2499 :   0 - 0x0
      12'h9C4: dout <= 8'b00000000; // 2500 :   0 - 0x0
      12'h9C5: dout <= 8'b00000000; // 2501 :   0 - 0x0
      12'h9C6: dout <= 8'b00000000; // 2502 :   0 - 0x0
      12'h9C7: dout <= 8'b00000000; // 2503 :   0 - 0x0
      12'h9C8: dout <= 8'b00000000; // 2504 :   0 - 0x0 -- Background 0x39
      12'h9C9: dout <= 8'b00000000; // 2505 :   0 - 0x0
      12'h9CA: dout <= 8'b00000000; // 2506 :   0 - 0x0
      12'h9CB: dout <= 8'b00000000; // 2507 :   0 - 0x0
      12'h9CC: dout <= 8'b00000000; // 2508 :   0 - 0x0
      12'h9CD: dout <= 8'b00000000; // 2509 :   0 - 0x0
      12'h9CE: dout <= 8'b00000000; // 2510 :   0 - 0x0
      12'h9CF: dout <= 8'b00000000; // 2511 :   0 - 0x0
      12'h9D0: dout <= 8'b00000000; // 2512 :   0 - 0x0 -- Background 0x3a
      12'h9D1: dout <= 8'b00000000; // 2513 :   0 - 0x0
      12'h9D2: dout <= 8'b00000000; // 2514 :   0 - 0x0
      12'h9D3: dout <= 8'b00000000; // 2515 :   0 - 0x0
      12'h9D4: dout <= 8'b00000000; // 2516 :   0 - 0x0
      12'h9D5: dout <= 8'b00000000; // 2517 :   0 - 0x0
      12'h9D6: dout <= 8'b00000000; // 2518 :   0 - 0x0
      12'h9D7: dout <= 8'b00000000; // 2519 :   0 - 0x0
      12'h9D8: dout <= 8'b00000000; // 2520 :   0 - 0x0 -- Background 0x3b
      12'h9D9: dout <= 8'b00000000; // 2521 :   0 - 0x0
      12'h9DA: dout <= 8'b00000000; // 2522 :   0 - 0x0
      12'h9DB: dout <= 8'b00000000; // 2523 :   0 - 0x0
      12'h9DC: dout <= 8'b00000000; // 2524 :   0 - 0x0
      12'h9DD: dout <= 8'b00000000; // 2525 :   0 - 0x0
      12'h9DE: dout <= 8'b00000000; // 2526 :   0 - 0x0
      12'h9DF: dout <= 8'b00000000; // 2527 :   0 - 0x0
      12'h9E0: dout <= 8'b00000000; // 2528 :   0 - 0x0 -- Background 0x3c
      12'h9E1: dout <= 8'b00000000; // 2529 :   0 - 0x0
      12'h9E2: dout <= 8'b00000000; // 2530 :   0 - 0x0
      12'h9E3: dout <= 8'b00000000; // 2531 :   0 - 0x0
      12'h9E4: dout <= 8'b00000000; // 2532 :   0 - 0x0
      12'h9E5: dout <= 8'b00000000; // 2533 :   0 - 0x0
      12'h9E6: dout <= 8'b00000000; // 2534 :   0 - 0x0
      12'h9E7: dout <= 8'b00000000; // 2535 :   0 - 0x0
      12'h9E8: dout <= 8'b00000000; // 2536 :   0 - 0x0 -- Background 0x3d
      12'h9E9: dout <= 8'b00000000; // 2537 :   0 - 0x0
      12'h9EA: dout <= 8'b00000000; // 2538 :   0 - 0x0
      12'h9EB: dout <= 8'b00000000; // 2539 :   0 - 0x0
      12'h9EC: dout <= 8'b00000000; // 2540 :   0 - 0x0
      12'h9ED: dout <= 8'b00000000; // 2541 :   0 - 0x0
      12'h9EE: dout <= 8'b00000000; // 2542 :   0 - 0x0
      12'h9EF: dout <= 8'b00000000; // 2543 :   0 - 0x0
      12'h9F0: dout <= 8'b00000000; // 2544 :   0 - 0x0 -- Background 0x3e
      12'h9F1: dout <= 8'b00000000; // 2545 :   0 - 0x0
      12'h9F2: dout <= 8'b00000000; // 2546 :   0 - 0x0
      12'h9F3: dout <= 8'b00000000; // 2547 :   0 - 0x0
      12'h9F4: dout <= 8'b00000000; // 2548 :   0 - 0x0
      12'h9F5: dout <= 8'b00000000; // 2549 :   0 - 0x0
      12'h9F6: dout <= 8'b00000000; // 2550 :   0 - 0x0
      12'h9F7: dout <= 8'b00000000; // 2551 :   0 - 0x0
      12'h9F8: dout <= 8'b00000000; // 2552 :   0 - 0x0 -- Background 0x3f
      12'h9F9: dout <= 8'b00000000; // 2553 :   0 - 0x0
      12'h9FA: dout <= 8'b00000000; // 2554 :   0 - 0x0
      12'h9FB: dout <= 8'b00000000; // 2555 :   0 - 0x0
      12'h9FC: dout <= 8'b00000000; // 2556 :   0 - 0x0
      12'h9FD: dout <= 8'b00000000; // 2557 :   0 - 0x0
      12'h9FE: dout <= 8'b00000000; // 2558 :   0 - 0x0
      12'h9FF: dout <= 8'b00000000; // 2559 :   0 - 0x0
      12'hA00: dout <= 8'b00000000; // 2560 :   0 - 0x0 -- Background 0x40
      12'hA01: dout <= 8'b00111110; // 2561 :  62 - 0x3e
      12'hA02: dout <= 8'b01111111; // 2562 : 127 - 0x7f
      12'hA03: dout <= 8'b01111111; // 2563 : 127 - 0x7f
      12'hA04: dout <= 8'b01111111; // 2564 : 127 - 0x7f
      12'hA05: dout <= 8'b01111111; // 2565 : 127 - 0x7f
      12'hA06: dout <= 8'b01111111; // 2566 : 127 - 0x7f
      12'hA07: dout <= 8'b00111110; // 2567 :  62 - 0x3e
      12'hA08: dout <= 8'b00000000; // 2568 :   0 - 0x0 -- Background 0x41
      12'hA09: dout <= 8'b00111100; // 2569 :  60 - 0x3c
      12'hA0A: dout <= 8'b00011100; // 2570 :  28 - 0x1c
      12'hA0B: dout <= 8'b00011100; // 2571 :  28 - 0x1c
      12'hA0C: dout <= 8'b00011100; // 2572 :  28 - 0x1c
      12'hA0D: dout <= 8'b00011100; // 2573 :  28 - 0x1c
      12'hA0E: dout <= 8'b00011100; // 2574 :  28 - 0x1c
      12'hA0F: dout <= 8'b00011100; // 2575 :  28 - 0x1c
      12'hA10: dout <= 8'b00000000; // 2576 :   0 - 0x0 -- Background 0x42
      12'hA11: dout <= 8'b01111100; // 2577 : 124 - 0x7c
      12'hA12: dout <= 8'b01111111; // 2578 : 127 - 0x7f
      12'hA13: dout <= 8'b01100111; // 2579 : 103 - 0x67
      12'hA14: dout <= 8'b00111111; // 2580 :  63 - 0x3f
      12'hA15: dout <= 8'b01111110; // 2581 : 126 - 0x7e
      12'hA16: dout <= 8'b01111111; // 2582 : 127 - 0x7f
      12'hA17: dout <= 8'b01111111; // 2583 : 127 - 0x7f
      12'hA18: dout <= 8'b00000000; // 2584 :   0 - 0x0 -- Background 0x43
      12'hA19: dout <= 8'b01111110; // 2585 : 126 - 0x7e
      12'hA1A: dout <= 8'b01111111; // 2586 : 127 - 0x7f
      12'hA1B: dout <= 8'b01111111; // 2587 : 127 - 0x7f
      12'hA1C: dout <= 8'b00011111; // 2588 :  31 - 0x1f
      12'hA1D: dout <= 8'b01110111; // 2589 : 119 - 0x77
      12'hA1E: dout <= 8'b01111111; // 2590 : 127 - 0x7f
      12'hA1F: dout <= 8'b01111110; // 2591 : 126 - 0x7e
      12'hA20: dout <= 8'b00000000; // 2592 :   0 - 0x0 -- Background 0x44
      12'hA21: dout <= 8'b00001110; // 2593 :  14 - 0xe
      12'hA22: dout <= 8'b00011110; // 2594 :  30 - 0x1e
      12'hA23: dout <= 8'b00111110; // 2595 :  62 - 0x3e
      12'hA24: dout <= 8'b01111110; // 2596 : 126 - 0x7e
      12'hA25: dout <= 8'b01111111; // 2597 : 127 - 0x7f
      12'hA26: dout <= 8'b01111110; // 2598 : 126 - 0x7e
      12'hA27: dout <= 8'b00001100; // 2599 :  12 - 0xc
      12'hA28: dout <= 8'b00000000; // 2600 :   0 - 0x0 -- Background 0x45
      12'hA29: dout <= 8'b01111111; // 2601 : 127 - 0x7f
      12'hA2A: dout <= 8'b01111111; // 2602 : 127 - 0x7f
      12'hA2B: dout <= 8'b01111111; // 2603 : 127 - 0x7f
      12'hA2C: dout <= 8'b01111111; // 2604 : 127 - 0x7f
      12'hA2D: dout <= 8'b01110111; // 2605 : 119 - 0x77
      12'hA2E: dout <= 8'b01111111; // 2606 : 127 - 0x7f
      12'hA2F: dout <= 8'b01111110; // 2607 : 126 - 0x7e
      12'hA30: dout <= 8'b00000000; // 2608 :   0 - 0x0 -- Background 0x46
      12'hA31: dout <= 8'b00111110; // 2609 :  62 - 0x3e
      12'hA32: dout <= 8'b01111110; // 2610 : 126 - 0x7e
      12'hA33: dout <= 8'b01111111; // 2611 : 127 - 0x7f
      12'hA34: dout <= 8'b01111111; // 2612 : 127 - 0x7f
      12'hA35: dout <= 8'b01110111; // 2613 : 119 - 0x77
      12'hA36: dout <= 8'b01111111; // 2614 : 127 - 0x7f
      12'hA37: dout <= 8'b00111110; // 2615 :  62 - 0x3e
      12'hA38: dout <= 8'b00000000; // 2616 :   0 - 0x0 -- Background 0x47
      12'hA39: dout <= 8'b01111110; // 2617 : 126 - 0x7e
      12'hA3A: dout <= 8'b01111110; // 2618 : 126 - 0x7e
      12'hA3B: dout <= 8'b00011110; // 2619 :  30 - 0x1e
      12'hA3C: dout <= 8'b00011100; // 2620 :  28 - 0x1c
      12'hA3D: dout <= 8'b00111100; // 2621 :  60 - 0x3c
      12'hA3E: dout <= 8'b00111000; // 2622 :  56 - 0x38
      12'hA3F: dout <= 8'b00111000; // 2623 :  56 - 0x38
      12'hA40: dout <= 8'b00000000; // 2624 :   0 - 0x0 -- Background 0x48
      12'hA41: dout <= 8'b00111110; // 2625 :  62 - 0x3e
      12'hA42: dout <= 8'b01111111; // 2626 : 127 - 0x7f
      12'hA43: dout <= 8'b01111111; // 2627 : 127 - 0x7f
      12'hA44: dout <= 8'b01111111; // 2628 : 127 - 0x7f
      12'hA45: dout <= 8'b01111111; // 2629 : 127 - 0x7f
      12'hA46: dout <= 8'b01111111; // 2630 : 127 - 0x7f
      12'hA47: dout <= 8'b00111110; // 2631 :  62 - 0x3e
      12'hA48: dout <= 8'b00000000; // 2632 :   0 - 0x0 -- Background 0x49
      12'hA49: dout <= 8'b00111110; // 2633 :  62 - 0x3e
      12'hA4A: dout <= 8'b01111111; // 2634 : 127 - 0x7f
      12'hA4B: dout <= 8'b01110111; // 2635 : 119 - 0x77
      12'hA4C: dout <= 8'b01111111; // 2636 : 127 - 0x7f
      12'hA4D: dout <= 8'b01111111; // 2637 : 127 - 0x7f
      12'hA4E: dout <= 8'b00111111; // 2638 :  63 - 0x3f
      12'hA4F: dout <= 8'b00111110; // 2639 :  62 - 0x3e
      12'hA50: dout <= 8'b11111111; // 2640 : 255 - 0xff -- Background 0x4a
      12'hA51: dout <= 8'b10011001; // 2641 : 153 - 0x99
      12'hA52: dout <= 8'b10011001; // 2642 : 153 - 0x99
      12'hA53: dout <= 8'b10011001; // 2643 : 153 - 0x99
      12'hA54: dout <= 8'b10011001; // 2644 : 153 - 0x99
      12'hA55: dout <= 8'b10011001; // 2645 : 153 - 0x99
      12'hA56: dout <= 8'b10011001; // 2646 : 153 - 0x99
      12'hA57: dout <= 8'b11111111; // 2647 : 255 - 0xff
      12'hA58: dout <= 8'b11110000; // 2648 : 240 - 0xf0 -- Background 0x4b
      12'hA59: dout <= 8'b10010000; // 2649 : 144 - 0x90
      12'hA5A: dout <= 8'b10010000; // 2650 : 144 - 0x90
      12'hA5B: dout <= 8'b10010000; // 2651 : 144 - 0x90
      12'hA5C: dout <= 8'b10010000; // 2652 : 144 - 0x90
      12'hA5D: dout <= 8'b10010000; // 2653 : 144 - 0x90
      12'hA5E: dout <= 8'b10010000; // 2654 : 144 - 0x90
      12'hA5F: dout <= 8'b11110000; // 2655 : 240 - 0xf0
      12'hA60: dout <= 8'b11111111; // 2656 : 255 - 0xff -- Background 0x4c
      12'hA61: dout <= 8'b11111111; // 2657 : 255 - 0xff
      12'hA62: dout <= 8'b11111111; // 2658 : 255 - 0xff
      12'hA63: dout <= 8'b11111111; // 2659 : 255 - 0xff
      12'hA64: dout <= 8'b11111111; // 2660 : 255 - 0xff
      12'hA65: dout <= 8'b11111111; // 2661 : 255 - 0xff
      12'hA66: dout <= 8'b11111111; // 2662 : 255 - 0xff
      12'hA67: dout <= 8'b11111111; // 2663 : 255 - 0xff
      12'hA68: dout <= 8'b11111111; // 2664 : 255 - 0xff -- Background 0x4d
      12'hA69: dout <= 8'b11111111; // 2665 : 255 - 0xff
      12'hA6A: dout <= 8'b11111111; // 2666 : 255 - 0xff
      12'hA6B: dout <= 8'b11111111; // 2667 : 255 - 0xff
      12'hA6C: dout <= 8'b11111111; // 2668 : 255 - 0xff
      12'hA6D: dout <= 8'b11111111; // 2669 : 255 - 0xff
      12'hA6E: dout <= 8'b11111111; // 2670 : 255 - 0xff
      12'hA6F: dout <= 8'b11111111; // 2671 : 255 - 0xff
      12'hA70: dout <= 8'b11111111; // 2672 : 255 - 0xff -- Background 0x4e
      12'hA71: dout <= 8'b11111111; // 2673 : 255 - 0xff
      12'hA72: dout <= 8'b11111111; // 2674 : 255 - 0xff
      12'hA73: dout <= 8'b11111111; // 2675 : 255 - 0xff
      12'hA74: dout <= 8'b11111111; // 2676 : 255 - 0xff
      12'hA75: dout <= 8'b11111111; // 2677 : 255 - 0xff
      12'hA76: dout <= 8'b11111111; // 2678 : 255 - 0xff
      12'hA77: dout <= 8'b11111111; // 2679 : 255 - 0xff
      12'hA78: dout <= 8'b11111111; // 2680 : 255 - 0xff -- Background 0x4f
      12'hA79: dout <= 8'b11111111; // 2681 : 255 - 0xff
      12'hA7A: dout <= 8'b11111111; // 2682 : 255 - 0xff
      12'hA7B: dout <= 8'b11111111; // 2683 : 255 - 0xff
      12'hA7C: dout <= 8'b11111111; // 2684 : 255 - 0xff
      12'hA7D: dout <= 8'b11111111; // 2685 : 255 - 0xff
      12'hA7E: dout <= 8'b11111111; // 2686 : 255 - 0xff
      12'hA7F: dout <= 8'b11111111; // 2687 : 255 - 0xff
      12'hA80: dout <= 8'b00010000; // 2688 :  16 - 0x10 -- Background 0x50
      12'hA81: dout <= 8'b00101000; // 2689 :  40 - 0x28
      12'hA82: dout <= 8'b11101110; // 2690 : 238 - 0xee
      12'hA83: dout <= 8'b10000010; // 2691 : 130 - 0x82
      12'hA84: dout <= 8'b01000100; // 2692 :  68 - 0x44
      12'hA85: dout <= 8'b01000100; // 2693 :  68 - 0x44
      12'hA86: dout <= 8'b10010010; // 2694 : 146 - 0x92
      12'hA87: dout <= 8'b11101110; // 2695 : 238 - 0xee
      12'hA88: dout <= 8'b00010000; // 2696 :  16 - 0x10 -- Background 0x51
      12'hA89: dout <= 8'b00101000; // 2697 :  40 - 0x28
      12'hA8A: dout <= 8'b11101110; // 2698 : 238 - 0xee
      12'hA8B: dout <= 8'b10000010; // 2699 : 130 - 0x82
      12'hA8C: dout <= 8'b01000100; // 2700 :  68 - 0x44
      12'hA8D: dout <= 8'b01000100; // 2701 :  68 - 0x44
      12'hA8E: dout <= 8'b10010010; // 2702 : 146 - 0x92
      12'hA8F: dout <= 8'b11101110; // 2703 : 238 - 0xee
      12'hA90: dout <= 8'b00010000; // 2704 :  16 - 0x10 -- Background 0x52
      12'hA91: dout <= 8'b00111000; // 2705 :  56 - 0x38
      12'hA92: dout <= 8'b11111110; // 2706 : 254 - 0xfe
      12'hA93: dout <= 8'b11111110; // 2707 : 254 - 0xfe
      12'hA94: dout <= 8'b01111100; // 2708 : 124 - 0x7c
      12'hA95: dout <= 8'b01111100; // 2709 : 124 - 0x7c
      12'hA96: dout <= 8'b11111110; // 2710 : 254 - 0xfe
      12'hA97: dout <= 8'b11101110; // 2711 : 238 - 0xee
      12'hA98: dout <= 8'b11111111; // 2712 : 255 - 0xff -- Background 0x53
      12'hA99: dout <= 8'b11111111; // 2713 : 255 - 0xff
      12'hA9A: dout <= 8'b11111111; // 2714 : 255 - 0xff
      12'hA9B: dout <= 8'b11111111; // 2715 : 255 - 0xff
      12'hA9C: dout <= 8'b11111111; // 2716 : 255 - 0xff
      12'hA9D: dout <= 8'b11111111; // 2717 : 255 - 0xff
      12'hA9E: dout <= 8'b11111111; // 2718 : 255 - 0xff
      12'hA9F: dout <= 8'b11111111; // 2719 : 255 - 0xff
      12'hAA0: dout <= 8'b00000000; // 2720 :   0 - 0x0 -- Background 0x54
      12'hAA1: dout <= 8'b00000000; // 2721 :   0 - 0x0
      12'hAA2: dout <= 8'b00000000; // 2722 :   0 - 0x0
      12'hAA3: dout <= 8'b00000000; // 2723 :   0 - 0x0
      12'hAA4: dout <= 8'b00000000; // 2724 :   0 - 0x0
      12'hAA5: dout <= 8'b00000000; // 2725 :   0 - 0x0
      12'hAA6: dout <= 8'b00000000; // 2726 :   0 - 0x0
      12'hAA7: dout <= 8'b00000000; // 2727 :   0 - 0x0
      12'hAA8: dout <= 8'b11111111; // 2728 : 255 - 0xff -- Background 0x55
      12'hAA9: dout <= 8'b11111111; // 2729 : 255 - 0xff
      12'hAAA: dout <= 8'b11111111; // 2730 : 255 - 0xff
      12'hAAB: dout <= 8'b11111111; // 2731 : 255 - 0xff
      12'hAAC: dout <= 8'b11111111; // 2732 : 255 - 0xff
      12'hAAD: dout <= 8'b11111111; // 2733 : 255 - 0xff
      12'hAAE: dout <= 8'b11111111; // 2734 : 255 - 0xff
      12'hAAF: dout <= 8'b11111111; // 2735 : 255 - 0xff
      12'hAB0: dout <= 8'b00101010; // 2736 :  42 - 0x2a -- Background 0x56
      12'hAB1: dout <= 8'b01000101; // 2737 :  69 - 0x45
      12'hAB2: dout <= 8'b00001000; // 2738 :   8 - 0x8
      12'hAB3: dout <= 8'b00010101; // 2739 :  21 - 0x15
      12'hAB4: dout <= 8'b00100000; // 2740 :  32 - 0x20
      12'hAB5: dout <= 8'b01000101; // 2741 :  69 - 0x45
      12'hAB6: dout <= 8'b10101000; // 2742 : 168 - 0xa8
      12'hAB7: dout <= 8'b00000000; // 2743 :   0 - 0x0
      12'hAB8: dout <= 8'b00001000; // 2744 :   8 - 0x8 -- Background 0x57
      12'hAB9: dout <= 8'b01010101; // 2745 :  85 - 0x55
      12'hABA: dout <= 8'b10100000; // 2746 : 160 - 0xa0
      12'hABB: dout <= 8'b00010000; // 2747 :  16 - 0x10
      12'hABC: dout <= 8'b10000000; // 2748 : 128 - 0x80
      12'hABD: dout <= 8'b00010100; // 2749 :  20 - 0x14
      12'hABE: dout <= 8'b00100010; // 2750 :  34 - 0x22
      12'hABF: dout <= 8'b00000000; // 2751 :   0 - 0x0
      12'hAC0: dout <= 8'b11111111; // 2752 : 255 - 0xff -- Background 0x58
      12'hAC1: dout <= 8'b11010101; // 2753 : 213 - 0xd5
      12'hAC2: dout <= 8'b10100000; // 2754 : 160 - 0xa0
      12'hAC3: dout <= 8'b11010000; // 2755 : 208 - 0xd0
      12'hAC4: dout <= 8'b10001111; // 2756 : 143 - 0x8f
      12'hAC5: dout <= 8'b11001000; // 2757 : 200 - 0xc8
      12'hAC6: dout <= 8'b10001000; // 2758 : 136 - 0x88
      12'hAC7: dout <= 8'b11001000; // 2759 : 200 - 0xc8
      12'hAC8: dout <= 8'b10001000; // 2760 : 136 - 0x88 -- Background 0x59
      12'hAC9: dout <= 8'b11001000; // 2761 : 200 - 0xc8
      12'hACA: dout <= 8'b10001000; // 2762 : 136 - 0x88
      12'hACB: dout <= 8'b11001111; // 2763 : 207 - 0xcf
      12'hACC: dout <= 8'b10010000; // 2764 : 144 - 0x90
      12'hACD: dout <= 8'b11100000; // 2765 : 224 - 0xe0
      12'hACE: dout <= 8'b11101010; // 2766 : 234 - 0xea
      12'hACF: dout <= 8'b11111111; // 2767 : 255 - 0xff
      12'hAD0: dout <= 8'b11111111; // 2768 : 255 - 0xff -- Background 0x5a
      12'hAD1: dout <= 8'b01011011; // 2769 :  91 - 0x5b
      12'hAD2: dout <= 8'b00000111; // 2770 :   7 - 0x7
      12'hAD3: dout <= 8'b00001001; // 2771 :   9 - 0x9
      12'hAD4: dout <= 8'b11110011; // 2772 : 243 - 0xf3
      12'hAD5: dout <= 8'b00010001; // 2773 :  17 - 0x11
      12'hAD6: dout <= 8'b00010011; // 2774 :  19 - 0x13
      12'hAD7: dout <= 8'b00010001; // 2775 :  17 - 0x11
      12'hAD8: dout <= 8'b00010011; // 2776 :  19 - 0x13 -- Background 0x5b
      12'hAD9: dout <= 8'b00010001; // 2777 :  17 - 0x11
      12'hADA: dout <= 8'b00010011; // 2778 :  19 - 0x13
      12'hADB: dout <= 8'b11110001; // 2779 : 241 - 0xf1
      12'hADC: dout <= 8'b00001011; // 2780 :  11 - 0xb
      12'hADD: dout <= 8'b00000101; // 2781 :   5 - 0x5
      12'hADE: dout <= 8'b10101011; // 2782 : 171 - 0xab
      12'hADF: dout <= 8'b11111111; // 2783 : 255 - 0xff
      12'hAE0: dout <= 8'b00011100; // 2784 :  28 - 0x1c -- Background 0x5c
      12'hAE1: dout <= 8'b00100010; // 2785 :  34 - 0x22
      12'hAE2: dout <= 8'b01000001; // 2786 :  65 - 0x41
      12'hAE3: dout <= 8'b01000001; // 2787 :  65 - 0x41
      12'hAE4: dout <= 8'b01000001; // 2788 :  65 - 0x41
      12'hAE5: dout <= 8'b00100010; // 2789 :  34 - 0x22
      12'hAE6: dout <= 8'b00100010; // 2790 :  34 - 0x22
      12'hAE7: dout <= 8'b00011100; // 2791 :  28 - 0x1c
      12'hAE8: dout <= 8'b00001000; // 2792 :   8 - 0x8 -- Background 0x5d
      12'hAE9: dout <= 8'b00010000; // 2793 :  16 - 0x10
      12'hAEA: dout <= 8'b00010000; // 2794 :  16 - 0x10
      12'hAEB: dout <= 8'b00001000; // 2795 :   8 - 0x8
      12'hAEC: dout <= 8'b00000100; // 2796 :   4 - 0x4
      12'hAED: dout <= 8'b00000100; // 2797 :   4 - 0x4
      12'hAEE: dout <= 8'b00001000; // 2798 :   8 - 0x8
      12'hAEF: dout <= 8'b00010000; // 2799 :  16 - 0x10
      12'hAF0: dout <= 8'b00110110; // 2800 :  54 - 0x36 -- Background 0x5e
      12'hAF1: dout <= 8'b01101011; // 2801 : 107 - 0x6b
      12'hAF2: dout <= 8'b01001001; // 2802 :  73 - 0x49
      12'hAF3: dout <= 8'b01000001; // 2803 :  65 - 0x41
      12'hAF4: dout <= 8'b01000001; // 2804 :  65 - 0x41
      12'hAF5: dout <= 8'b00100010; // 2805 :  34 - 0x22
      12'hAF6: dout <= 8'b00010100; // 2806 :  20 - 0x14
      12'hAF7: dout <= 8'b00001000; // 2807 :   8 - 0x8
      12'hAF8: dout <= 8'b00111110; // 2808 :  62 - 0x3e -- Background 0x5f
      12'hAF9: dout <= 8'b01101011; // 2809 : 107 - 0x6b
      12'hAFA: dout <= 8'b00100010; // 2810 :  34 - 0x22
      12'hAFB: dout <= 8'b01100011; // 2811 :  99 - 0x63
      12'hAFC: dout <= 8'b00100010; // 2812 :  34 - 0x22
      12'hAFD: dout <= 8'b01100011; // 2813 :  99 - 0x63
      12'hAFE: dout <= 8'b00100010; // 2814 :  34 - 0x22
      12'hAFF: dout <= 8'b01111111; // 2815 : 127 - 0x7f
      12'hB00: dout <= 8'b11111111; // 2816 : 255 - 0xff -- Background 0x60
      12'hB01: dout <= 8'b11111111; // 2817 : 255 - 0xff
      12'hB02: dout <= 8'b11111111; // 2818 : 255 - 0xff
      12'hB03: dout <= 8'b11111111; // 2819 : 255 - 0xff
      12'hB04: dout <= 8'b11010101; // 2820 : 213 - 0xd5
      12'hB05: dout <= 8'b10101010; // 2821 : 170 - 0xaa
      12'hB06: dout <= 8'b11010101; // 2822 : 213 - 0xd5
      12'hB07: dout <= 8'b11111111; // 2823 : 255 - 0xff
      12'hB08: dout <= 8'b11111111; // 2824 : 255 - 0xff -- Background 0x61
      12'hB09: dout <= 8'b11111111; // 2825 : 255 - 0xff
      12'hB0A: dout <= 8'b11111111; // 2826 : 255 - 0xff
      12'hB0B: dout <= 8'b11111111; // 2827 : 255 - 0xff
      12'hB0C: dout <= 8'b01010101; // 2828 :  85 - 0x55
      12'hB0D: dout <= 8'b10101010; // 2829 : 170 - 0xaa
      12'hB0E: dout <= 8'b01010101; // 2830 :  85 - 0x55
      12'hB0F: dout <= 8'b11111111; // 2831 : 255 - 0xff
      12'hB10: dout <= 8'b11111111; // 2832 : 255 - 0xff -- Background 0x62
      12'hB11: dout <= 8'b11111111; // 2833 : 255 - 0xff
      12'hB12: dout <= 8'b11111111; // 2834 : 255 - 0xff
      12'hB13: dout <= 8'b11111111; // 2835 : 255 - 0xff
      12'hB14: dout <= 8'b01010101; // 2836 :  85 - 0x55
      12'hB15: dout <= 8'b10101011; // 2837 : 171 - 0xab
      12'hB16: dout <= 8'b01010101; // 2838 :  85 - 0x55
      12'hB17: dout <= 8'b11111111; // 2839 : 255 - 0xff
      12'hB18: dout <= 8'b00000000; // 2840 :   0 - 0x0 -- Background 0x63
      12'hB19: dout <= 8'b00000000; // 2841 :   0 - 0x0
      12'hB1A: dout <= 8'b00000000; // 2842 :   0 - 0x0
      12'hB1B: dout <= 8'b00000000; // 2843 :   0 - 0x0
      12'hB1C: dout <= 8'b00000000; // 2844 :   0 - 0x0
      12'hB1D: dout <= 8'b00000000; // 2845 :   0 - 0x0
      12'hB1E: dout <= 8'b00000000; // 2846 :   0 - 0x0
      12'hB1F: dout <= 8'b00000000; // 2847 :   0 - 0x0
      12'hB20: dout <= 8'b00000001; // 2848 :   1 - 0x1 -- Background 0x64
      12'hB21: dout <= 8'b00000001; // 2849 :   1 - 0x1
      12'hB22: dout <= 8'b00000011; // 2850 :   3 - 0x3
      12'hB23: dout <= 8'b00000011; // 2851 :   3 - 0x3
      12'hB24: dout <= 8'b00000110; // 2852 :   6 - 0x6
      12'hB25: dout <= 8'b00000110; // 2853 :   6 - 0x6
      12'hB26: dout <= 8'b00001100; // 2854 :  12 - 0xc
      12'hB27: dout <= 8'b00001100; // 2855 :  12 - 0xc
      12'hB28: dout <= 8'b00011000; // 2856 :  24 - 0x18 -- Background 0x65
      12'hB29: dout <= 8'b00011000; // 2857 :  24 - 0x18
      12'hB2A: dout <= 8'b00110000; // 2858 :  48 - 0x30
      12'hB2B: dout <= 8'b00110000; // 2859 :  48 - 0x30
      12'hB2C: dout <= 8'b01100000; // 2860 :  96 - 0x60
      12'hB2D: dout <= 8'b01100000; // 2861 :  96 - 0x60
      12'hB2E: dout <= 8'b11101010; // 2862 : 234 - 0xea
      12'hB2F: dout <= 8'b11111111; // 2863 : 255 - 0xff
      12'hB30: dout <= 8'b10000000; // 2864 : 128 - 0x80 -- Background 0x66
      12'hB31: dout <= 8'b10000000; // 2865 : 128 - 0x80
      12'hB32: dout <= 8'b11000000; // 2866 : 192 - 0xc0
      12'hB33: dout <= 8'b01000000; // 2867 :  64 - 0x40
      12'hB34: dout <= 8'b10100000; // 2868 : 160 - 0xa0
      12'hB35: dout <= 8'b01100000; // 2869 :  96 - 0x60
      12'hB36: dout <= 8'b00110000; // 2870 :  48 - 0x30
      12'hB37: dout <= 8'b00010000; // 2871 :  16 - 0x10
      12'hB38: dout <= 8'b00101000; // 2872 :  40 - 0x28 -- Background 0x67
      12'hB39: dout <= 8'b00011000; // 2873 :  24 - 0x18
      12'hB3A: dout <= 8'b00001100; // 2874 :  12 - 0xc
      12'hB3B: dout <= 8'b00010100; // 2875 :  20 - 0x14
      12'hB3C: dout <= 8'b00001010; // 2876 :  10 - 0xa
      12'hB3D: dout <= 8'b00000110; // 2877 :   6 - 0x6
      12'hB3E: dout <= 8'b10101011; // 2878 : 171 - 0xab
      12'hB3F: dout <= 8'b11111111; // 2879 : 255 - 0xff
      12'hB40: dout <= 8'b00000000; // 2880 :   0 - 0x0 -- Background 0x68
      12'hB41: dout <= 8'b00000000; // 2881 :   0 - 0x0
      12'hB42: dout <= 8'b00000000; // 2882 :   0 - 0x0
      12'hB43: dout <= 8'b00000000; // 2883 :   0 - 0x0
      12'hB44: dout <= 8'b00000000; // 2884 :   0 - 0x0
      12'hB45: dout <= 8'b00000000; // 2885 :   0 - 0x0
      12'hB46: dout <= 8'b00000000; // 2886 :   0 - 0x0
      12'hB47: dout <= 8'b00000000; // 2887 :   0 - 0x0
      12'hB48: dout <= 8'b00000000; // 2888 :   0 - 0x0 -- Background 0x69
      12'hB49: dout <= 8'b00000000; // 2889 :   0 - 0x0
      12'hB4A: dout <= 8'b00000000; // 2890 :   0 - 0x0
      12'hB4B: dout <= 8'b00000000; // 2891 :   0 - 0x0
      12'hB4C: dout <= 8'b00000000; // 2892 :   0 - 0x0
      12'hB4D: dout <= 8'b00000000; // 2893 :   0 - 0x0
      12'hB4E: dout <= 8'b00000000; // 2894 :   0 - 0x0
      12'hB4F: dout <= 8'b00000000; // 2895 :   0 - 0x0
      12'hB50: dout <= 8'b00000000; // 2896 :   0 - 0x0 -- Background 0x6a
      12'hB51: dout <= 8'b00000000; // 2897 :   0 - 0x0
      12'hB52: dout <= 8'b00000000; // 2898 :   0 - 0x0
      12'hB53: dout <= 8'b00000000; // 2899 :   0 - 0x0
      12'hB54: dout <= 8'b00000000; // 2900 :   0 - 0x0
      12'hB55: dout <= 8'b00000000; // 2901 :   0 - 0x0
      12'hB56: dout <= 8'b00000000; // 2902 :   0 - 0x0
      12'hB57: dout <= 8'b00000000; // 2903 :   0 - 0x0
      12'hB58: dout <= 8'b00000000; // 2904 :   0 - 0x0 -- Background 0x6b
      12'hB59: dout <= 8'b00000000; // 2905 :   0 - 0x0
      12'hB5A: dout <= 8'b00000000; // 2906 :   0 - 0x0
      12'hB5B: dout <= 8'b00000000; // 2907 :   0 - 0x0
      12'hB5C: dout <= 8'b00000000; // 2908 :   0 - 0x0
      12'hB5D: dout <= 8'b00000000; // 2909 :   0 - 0x0
      12'hB5E: dout <= 8'b00000000; // 2910 :   0 - 0x0
      12'hB5F: dout <= 8'b00000000; // 2911 :   0 - 0x0
      12'hB60: dout <= 8'b00000000; // 2912 :   0 - 0x0 -- Background 0x6c
      12'hB61: dout <= 8'b00000000; // 2913 :   0 - 0x0
      12'hB62: dout <= 8'b00000000; // 2914 :   0 - 0x0
      12'hB63: dout <= 8'b00000000; // 2915 :   0 - 0x0
      12'hB64: dout <= 8'b00000000; // 2916 :   0 - 0x0
      12'hB65: dout <= 8'b00000000; // 2917 :   0 - 0x0
      12'hB66: dout <= 8'b00000000; // 2918 :   0 - 0x0
      12'hB67: dout <= 8'b00000000; // 2919 :   0 - 0x0
      12'hB68: dout <= 8'b00000000; // 2920 :   0 - 0x0 -- Background 0x6d
      12'hB69: dout <= 8'b00000000; // 2921 :   0 - 0x0
      12'hB6A: dout <= 8'b00000000; // 2922 :   0 - 0x0
      12'hB6B: dout <= 8'b00000000; // 2923 :   0 - 0x0
      12'hB6C: dout <= 8'b00000000; // 2924 :   0 - 0x0
      12'hB6D: dout <= 8'b00000000; // 2925 :   0 - 0x0
      12'hB6E: dout <= 8'b00000000; // 2926 :   0 - 0x0
      12'hB6F: dout <= 8'b00000000; // 2927 :   0 - 0x0
      12'hB70: dout <= 8'b00000000; // 2928 :   0 - 0x0 -- Background 0x6e
      12'hB71: dout <= 8'b00000000; // 2929 :   0 - 0x0
      12'hB72: dout <= 8'b00000000; // 2930 :   0 - 0x0
      12'hB73: dout <= 8'b00000000; // 2931 :   0 - 0x0
      12'hB74: dout <= 8'b00000000; // 2932 :   0 - 0x0
      12'hB75: dout <= 8'b00000000; // 2933 :   0 - 0x0
      12'hB76: dout <= 8'b00000000; // 2934 :   0 - 0x0
      12'hB77: dout <= 8'b00000000; // 2935 :   0 - 0x0
      12'hB78: dout <= 8'b00000000; // 2936 :   0 - 0x0 -- Background 0x6f
      12'hB79: dout <= 8'b00000000; // 2937 :   0 - 0x0
      12'hB7A: dout <= 8'b00000000; // 2938 :   0 - 0x0
      12'hB7B: dout <= 8'b00000000; // 2939 :   0 - 0x0
      12'hB7C: dout <= 8'b00000000; // 2940 :   0 - 0x0
      12'hB7D: dout <= 8'b00000000; // 2941 :   0 - 0x0
      12'hB7E: dout <= 8'b00000000; // 2942 :   0 - 0x0
      12'hB7F: dout <= 8'b00000000; // 2943 :   0 - 0x0
      12'hB80: dout <= 8'b00000000; // 2944 :   0 - 0x0 -- Background 0x70
      12'hB81: dout <= 8'b00000000; // 2945 :   0 - 0x0
      12'hB82: dout <= 8'b00000000; // 2946 :   0 - 0x0
      12'hB83: dout <= 8'b00000000; // 2947 :   0 - 0x0
      12'hB84: dout <= 8'b00000000; // 2948 :   0 - 0x0
      12'hB85: dout <= 8'b00000000; // 2949 :   0 - 0x0
      12'hB86: dout <= 8'b00000000; // 2950 :   0 - 0x0
      12'hB87: dout <= 8'b00000000; // 2951 :   0 - 0x0
      12'hB88: dout <= 8'b00000000; // 2952 :   0 - 0x0 -- Background 0x71
      12'hB89: dout <= 8'b00000000; // 2953 :   0 - 0x0
      12'hB8A: dout <= 8'b00000000; // 2954 :   0 - 0x0
      12'hB8B: dout <= 8'b00000000; // 2955 :   0 - 0x0
      12'hB8C: dout <= 8'b00000000; // 2956 :   0 - 0x0
      12'hB8D: dout <= 8'b00000000; // 2957 :   0 - 0x0
      12'hB8E: dout <= 8'b00000000; // 2958 :   0 - 0x0
      12'hB8F: dout <= 8'b00000000; // 2959 :   0 - 0x0
      12'hB90: dout <= 8'b00000000; // 2960 :   0 - 0x0 -- Background 0x72
      12'hB91: dout <= 8'b00000000; // 2961 :   0 - 0x0
      12'hB92: dout <= 8'b00000000; // 2962 :   0 - 0x0
      12'hB93: dout <= 8'b00000000; // 2963 :   0 - 0x0
      12'hB94: dout <= 8'b00000000; // 2964 :   0 - 0x0
      12'hB95: dout <= 8'b00000000; // 2965 :   0 - 0x0
      12'hB96: dout <= 8'b00000000; // 2966 :   0 - 0x0
      12'hB97: dout <= 8'b00000000; // 2967 :   0 - 0x0
      12'hB98: dout <= 8'b00000000; // 2968 :   0 - 0x0 -- Background 0x73
      12'hB99: dout <= 8'b00000000; // 2969 :   0 - 0x0
      12'hB9A: dout <= 8'b00000000; // 2970 :   0 - 0x0
      12'hB9B: dout <= 8'b00000000; // 2971 :   0 - 0x0
      12'hB9C: dout <= 8'b00000000; // 2972 :   0 - 0x0
      12'hB9D: dout <= 8'b00000000; // 2973 :   0 - 0x0
      12'hB9E: dout <= 8'b00000000; // 2974 :   0 - 0x0
      12'hB9F: dout <= 8'b00000000; // 2975 :   0 - 0x0
      12'hBA0: dout <= 8'b00000000; // 2976 :   0 - 0x0 -- Background 0x74
      12'hBA1: dout <= 8'b00000000; // 2977 :   0 - 0x0
      12'hBA2: dout <= 8'b00000000; // 2978 :   0 - 0x0
      12'hBA3: dout <= 8'b00000000; // 2979 :   0 - 0x0
      12'hBA4: dout <= 8'b00000000; // 2980 :   0 - 0x0
      12'hBA5: dout <= 8'b00000000; // 2981 :   0 - 0x0
      12'hBA6: dout <= 8'b00000000; // 2982 :   0 - 0x0
      12'hBA7: dout <= 8'b00000000; // 2983 :   0 - 0x0
      12'hBA8: dout <= 8'b00000000; // 2984 :   0 - 0x0 -- Background 0x75
      12'hBA9: dout <= 8'b00000000; // 2985 :   0 - 0x0
      12'hBAA: dout <= 8'b00000000; // 2986 :   0 - 0x0
      12'hBAB: dout <= 8'b00000000; // 2987 :   0 - 0x0
      12'hBAC: dout <= 8'b00000000; // 2988 :   0 - 0x0
      12'hBAD: dout <= 8'b00000000; // 2989 :   0 - 0x0
      12'hBAE: dout <= 8'b00000000; // 2990 :   0 - 0x0
      12'hBAF: dout <= 8'b00000000; // 2991 :   0 - 0x0
      12'hBB0: dout <= 8'b00000000; // 2992 :   0 - 0x0 -- Background 0x76
      12'hBB1: dout <= 8'b00000000; // 2993 :   0 - 0x0
      12'hBB2: dout <= 8'b00000000; // 2994 :   0 - 0x0
      12'hBB3: dout <= 8'b00000000; // 2995 :   0 - 0x0
      12'hBB4: dout <= 8'b00000000; // 2996 :   0 - 0x0
      12'hBB5: dout <= 8'b00000000; // 2997 :   0 - 0x0
      12'hBB6: dout <= 8'b00000000; // 2998 :   0 - 0x0
      12'hBB7: dout <= 8'b00000000; // 2999 :   0 - 0x0
      12'hBB8: dout <= 8'b00000000; // 3000 :   0 - 0x0 -- Background 0x77
      12'hBB9: dout <= 8'b00000000; // 3001 :   0 - 0x0
      12'hBBA: dout <= 8'b00000000; // 3002 :   0 - 0x0
      12'hBBB: dout <= 8'b00000000; // 3003 :   0 - 0x0
      12'hBBC: dout <= 8'b00000000; // 3004 :   0 - 0x0
      12'hBBD: dout <= 8'b00000000; // 3005 :   0 - 0x0
      12'hBBE: dout <= 8'b00000000; // 3006 :   0 - 0x0
      12'hBBF: dout <= 8'b00000000; // 3007 :   0 - 0x0
      12'hBC0: dout <= 8'b00000000; // 3008 :   0 - 0x0 -- Background 0x78
      12'hBC1: dout <= 8'b00000000; // 3009 :   0 - 0x0
      12'hBC2: dout <= 8'b00000000; // 3010 :   0 - 0x0
      12'hBC3: dout <= 8'b00000000; // 3011 :   0 - 0x0
      12'hBC4: dout <= 8'b00000000; // 3012 :   0 - 0x0
      12'hBC5: dout <= 8'b00000000; // 3013 :   0 - 0x0
      12'hBC6: dout <= 8'b00000000; // 3014 :   0 - 0x0
      12'hBC7: dout <= 8'b00000000; // 3015 :   0 - 0x0
      12'hBC8: dout <= 8'b00000000; // 3016 :   0 - 0x0 -- Background 0x79
      12'hBC9: dout <= 8'b00000000; // 3017 :   0 - 0x0
      12'hBCA: dout <= 8'b00000000; // 3018 :   0 - 0x0
      12'hBCB: dout <= 8'b00000000; // 3019 :   0 - 0x0
      12'hBCC: dout <= 8'b00000000; // 3020 :   0 - 0x0
      12'hBCD: dout <= 8'b00000000; // 3021 :   0 - 0x0
      12'hBCE: dout <= 8'b00000000; // 3022 :   0 - 0x0
      12'hBCF: dout <= 8'b00000000; // 3023 :   0 - 0x0
      12'hBD0: dout <= 8'b00000000; // 3024 :   0 - 0x0 -- Background 0x7a
      12'hBD1: dout <= 8'b00000000; // 3025 :   0 - 0x0
      12'hBD2: dout <= 8'b00000000; // 3026 :   0 - 0x0
      12'hBD3: dout <= 8'b00000000; // 3027 :   0 - 0x0
      12'hBD4: dout <= 8'b00000000; // 3028 :   0 - 0x0
      12'hBD5: dout <= 8'b00000000; // 3029 :   0 - 0x0
      12'hBD6: dout <= 8'b00000000; // 3030 :   0 - 0x0
      12'hBD7: dout <= 8'b00000000; // 3031 :   0 - 0x0
      12'hBD8: dout <= 8'b00000000; // 3032 :   0 - 0x0 -- Background 0x7b
      12'hBD9: dout <= 8'b00000000; // 3033 :   0 - 0x0
      12'hBDA: dout <= 8'b00000000; // 3034 :   0 - 0x0
      12'hBDB: dout <= 8'b00000000; // 3035 :   0 - 0x0
      12'hBDC: dout <= 8'b00000000; // 3036 :   0 - 0x0
      12'hBDD: dout <= 8'b00000000; // 3037 :   0 - 0x0
      12'hBDE: dout <= 8'b00000000; // 3038 :   0 - 0x0
      12'hBDF: dout <= 8'b00000000; // 3039 :   0 - 0x0
      12'hBE0: dout <= 8'b00000000; // 3040 :   0 - 0x0 -- Background 0x7c
      12'hBE1: dout <= 8'b00000000; // 3041 :   0 - 0x0
      12'hBE2: dout <= 8'b00000000; // 3042 :   0 - 0x0
      12'hBE3: dout <= 8'b00000000; // 3043 :   0 - 0x0
      12'hBE4: dout <= 8'b00000000; // 3044 :   0 - 0x0
      12'hBE5: dout <= 8'b00000000; // 3045 :   0 - 0x0
      12'hBE6: dout <= 8'b00000000; // 3046 :   0 - 0x0
      12'hBE7: dout <= 8'b00000000; // 3047 :   0 - 0x0
      12'hBE8: dout <= 8'b00000000; // 3048 :   0 - 0x0 -- Background 0x7d
      12'hBE9: dout <= 8'b00000000; // 3049 :   0 - 0x0
      12'hBEA: dout <= 8'b00000000; // 3050 :   0 - 0x0
      12'hBEB: dout <= 8'b00000000; // 3051 :   0 - 0x0
      12'hBEC: dout <= 8'b00000000; // 3052 :   0 - 0x0
      12'hBED: dout <= 8'b00000000; // 3053 :   0 - 0x0
      12'hBEE: dout <= 8'b00000000; // 3054 :   0 - 0x0
      12'hBEF: dout <= 8'b00000000; // 3055 :   0 - 0x0
      12'hBF0: dout <= 8'b00000000; // 3056 :   0 - 0x0 -- Background 0x7e
      12'hBF1: dout <= 8'b00000000; // 3057 :   0 - 0x0
      12'hBF2: dout <= 8'b00000000; // 3058 :   0 - 0x0
      12'hBF3: dout <= 8'b00000000; // 3059 :   0 - 0x0
      12'hBF4: dout <= 8'b00000000; // 3060 :   0 - 0x0
      12'hBF5: dout <= 8'b00000000; // 3061 :   0 - 0x0
      12'hBF6: dout <= 8'b00000000; // 3062 :   0 - 0x0
      12'hBF7: dout <= 8'b00000000; // 3063 :   0 - 0x0
      12'hBF8: dout <= 8'b00000000; // 3064 :   0 - 0x0 -- Background 0x7f
      12'hBF9: dout <= 8'b00000000; // 3065 :   0 - 0x0
      12'hBFA: dout <= 8'b00000000; // 3066 :   0 - 0x0
      12'hBFB: dout <= 8'b00000000; // 3067 :   0 - 0x0
      12'hBFC: dout <= 8'b00000000; // 3068 :   0 - 0x0
      12'hBFD: dout <= 8'b00000000; // 3069 :   0 - 0x0
      12'hBFE: dout <= 8'b00000000; // 3070 :   0 - 0x0
      12'hBFF: dout <= 8'b00000000; // 3071 :   0 - 0x0
      12'hC00: dout <= 8'b00000011; // 3072 :   3 - 0x3 -- Background 0x80
      12'hC01: dout <= 8'b00001111; // 3073 :  15 - 0xf
      12'hC02: dout <= 8'b00011100; // 3074 :  28 - 0x1c
      12'hC03: dout <= 8'b00110000; // 3075 :  48 - 0x30
      12'hC04: dout <= 8'b00100000; // 3076 :  32 - 0x20
      12'hC05: dout <= 8'b01000000; // 3077 :  64 - 0x40
      12'hC06: dout <= 8'b01000000; // 3078 :  64 - 0x40
      12'hC07: dout <= 8'b01111111; // 3079 : 127 - 0x7f
      12'hC08: dout <= 8'b00000001; // 3080 :   1 - 0x1 -- Background 0x81
      12'hC09: dout <= 8'b00000001; // 3081 :   1 - 0x1
      12'hC0A: dout <= 8'b00000001; // 3082 :   1 - 0x1
      12'hC0B: dout <= 8'b00000001; // 3083 :   1 - 0x1
      12'hC0C: dout <= 8'b00000001; // 3084 :   1 - 0x1
      12'hC0D: dout <= 8'b00000001; // 3085 :   1 - 0x1
      12'hC0E: dout <= 8'b00000011; // 3086 :   3 - 0x3
      12'hC0F: dout <= 8'b00000011; // 3087 :   3 - 0x3
      12'hC10: dout <= 8'b11000000; // 3088 : 192 - 0xc0 -- Background 0x82
      12'hC11: dout <= 8'b11110000; // 3089 : 240 - 0xf0
      12'hC12: dout <= 8'b00111000; // 3090 :  56 - 0x38
      12'hC13: dout <= 8'b00001110; // 3091 :  14 - 0xe
      12'hC14: dout <= 8'b00011110; // 3092 :  30 - 0x1e
      12'hC15: dout <= 8'b00011110; // 3093 :  30 - 0x1e
      12'hC16: dout <= 8'b00000010; // 3094 :   2 - 0x2
      12'hC17: dout <= 8'b11111110; // 3095 : 254 - 0xfe
      12'hC18: dout <= 8'b10000000; // 3096 : 128 - 0x80 -- Background 0x83
      12'hC19: dout <= 8'b10000000; // 3097 : 128 - 0x80
      12'hC1A: dout <= 8'b10000000; // 3098 : 128 - 0x80
      12'hC1B: dout <= 8'b10000000; // 3099 : 128 - 0x80
      12'hC1C: dout <= 8'b10000000; // 3100 : 128 - 0x80
      12'hC1D: dout <= 8'b11100000; // 3101 : 224 - 0xe0
      12'hC1E: dout <= 8'b00010000; // 3102 :  16 - 0x10
      12'hC1F: dout <= 8'b11110000; // 3103 : 240 - 0xf0
      12'hC20: dout <= 8'b00000011; // 3104 :   3 - 0x3 -- Background 0x84
      12'hC21: dout <= 8'b00001111; // 3105 :  15 - 0xf
      12'hC22: dout <= 8'b00011100; // 3106 :  28 - 0x1c
      12'hC23: dout <= 8'b00110000; // 3107 :  48 - 0x30
      12'hC24: dout <= 8'b00100000; // 3108 :  32 - 0x20
      12'hC25: dout <= 8'b01000000; // 3109 :  64 - 0x40
      12'hC26: dout <= 8'b01000000; // 3110 :  64 - 0x40
      12'hC27: dout <= 8'b01111111; // 3111 : 127 - 0x7f
      12'hC28: dout <= 8'b00000011; // 3112 :   3 - 0x3 -- Background 0x85
      12'hC29: dout <= 8'b00000110; // 3113 :   6 - 0x6
      12'hC2A: dout <= 8'b00000110; // 3114 :   6 - 0x6
      12'hC2B: dout <= 8'b00011100; // 3115 :  28 - 0x1c
      12'hC2C: dout <= 8'b00011000; // 3116 :  24 - 0x18
      12'hC2D: dout <= 8'b00110110; // 3117 :  54 - 0x36
      12'hC2E: dout <= 8'b00110001; // 3118 :  49 - 0x31
      12'hC2F: dout <= 8'b00001111; // 3119 :  15 - 0xf
      12'hC30: dout <= 8'b11000000; // 3120 : 192 - 0xc0 -- Background 0x86
      12'hC31: dout <= 8'b11110000; // 3121 : 240 - 0xf0
      12'hC32: dout <= 8'b00111000; // 3122 :  56 - 0x38
      12'hC33: dout <= 8'b00001110; // 3123 :  14 - 0xe
      12'hC34: dout <= 8'b00011110; // 3124 :  30 - 0x1e
      12'hC35: dout <= 8'b00011110; // 3125 :  30 - 0x1e
      12'hC36: dout <= 8'b00000010; // 3126 :   2 - 0x2
      12'hC37: dout <= 8'b11111110; // 3127 : 254 - 0xfe
      12'hC38: dout <= 8'b11000000; // 3128 : 192 - 0xc0 -- Background 0x87
      12'hC39: dout <= 8'b01100000; // 3129 :  96 - 0x60
      12'hC3A: dout <= 8'b01100000; // 3130 :  96 - 0x60
      12'hC3B: dout <= 8'b00110000; // 3131 :  48 - 0x30
      12'hC3C: dout <= 8'b00111110; // 3132 :  62 - 0x3e
      12'hC3D: dout <= 8'b00011001; // 3133 :  25 - 0x19
      12'hC3E: dout <= 8'b00110011; // 3134 :  51 - 0x33
      12'hC3F: dout <= 8'b00111100; // 3135 :  60 - 0x3c
      12'hC40: dout <= 8'b00000011; // 3136 :   3 - 0x3 -- Background 0x88
      12'hC41: dout <= 8'b00000111; // 3137 :   7 - 0x7
      12'hC42: dout <= 8'b00000111; // 3138 :   7 - 0x7
      12'hC43: dout <= 8'b00001011; // 3139 :  11 - 0xb
      12'hC44: dout <= 8'b00010000; // 3140 :  16 - 0x10
      12'hC45: dout <= 8'b01100000; // 3141 :  96 - 0x60
      12'hC46: dout <= 8'b11110000; // 3142 : 240 - 0xf0
      12'hC47: dout <= 8'b11110000; // 3143 : 240 - 0xf0
      12'hC48: dout <= 8'b11110000; // 3144 : 240 - 0xf0 -- Background 0x89
      12'hC49: dout <= 8'b11110000; // 3145 : 240 - 0xf0
      12'hC4A: dout <= 8'b01100000; // 3146 :  96 - 0x60
      12'hC4B: dout <= 8'b00010000; // 3147 :  16 - 0x10
      12'hC4C: dout <= 8'b00001011; // 3148 :  11 - 0xb
      12'hC4D: dout <= 8'b00000111; // 3149 :   7 - 0x7
      12'hC4E: dout <= 8'b00000111; // 3150 :   7 - 0x7
      12'hC4F: dout <= 8'b00000011; // 3151 :   3 - 0x3
      12'hC50: dout <= 8'b00000000; // 3152 :   0 - 0x0 -- Background 0x8a
      12'hC51: dout <= 8'b00011100; // 3153 :  28 - 0x1c
      12'hC52: dout <= 8'b00111111; // 3154 :  63 - 0x3f
      12'hC53: dout <= 8'b01111000; // 3155 : 120 - 0x78
      12'hC54: dout <= 8'b01110000; // 3156 : 112 - 0x70
      12'hC55: dout <= 8'b01100000; // 3157 :  96 - 0x60
      12'hC56: dout <= 8'b00100000; // 3158 :  32 - 0x20
      12'hC57: dout <= 8'b00100000; // 3159 :  32 - 0x20
      12'hC58: dout <= 8'b00100000; // 3160 :  32 - 0x20 -- Background 0x8b
      12'hC59: dout <= 8'b00100000; // 3161 :  32 - 0x20
      12'hC5A: dout <= 8'b01100000; // 3162 :  96 - 0x60
      12'hC5B: dout <= 8'b01110000; // 3163 : 112 - 0x70
      12'hC5C: dout <= 8'b01111000; // 3164 : 120 - 0x78
      12'hC5D: dout <= 8'b00111111; // 3165 :  63 - 0x3f
      12'hC5E: dout <= 8'b00011100; // 3166 :  28 - 0x1c
      12'hC5F: dout <= 8'b00000000; // 3167 :   0 - 0x0
      12'hC60: dout <= 8'b00000011; // 3168 :   3 - 0x3 -- Background 0x8c
      12'hC61: dout <= 8'b00001100; // 3169 :  12 - 0xc
      12'hC62: dout <= 8'b00011110; // 3170 :  30 - 0x1e
      12'hC63: dout <= 8'b00100110; // 3171 :  38 - 0x26
      12'hC64: dout <= 8'b01000110; // 3172 :  70 - 0x46
      12'hC65: dout <= 8'b01100100; // 3173 : 100 - 0x64
      12'hC66: dout <= 8'b01110000; // 3174 : 112 - 0x70
      12'hC67: dout <= 8'b11110000; // 3175 : 240 - 0xf0
      12'hC68: dout <= 8'b10101010; // 3176 : 170 - 0xaa -- Background 0x8d
      12'hC69: dout <= 8'b11111111; // 3177 : 255 - 0xff
      12'hC6A: dout <= 8'b01111111; // 3178 : 127 - 0x7f
      12'hC6B: dout <= 8'b00111001; // 3179 :  57 - 0x39
      12'hC6C: dout <= 8'b00011001; // 3180 :  25 - 0x19
      12'hC6D: dout <= 8'b00001011; // 3181 :  11 - 0xb
      12'hC6E: dout <= 8'b00001000; // 3182 :   8 - 0x8
      12'hC6F: dout <= 8'b00000111; // 3183 :   7 - 0x7
      12'hC70: dout <= 8'b11000000; // 3184 : 192 - 0xc0 -- Background 0x8e
      12'hC71: dout <= 8'b00110000; // 3185 :  48 - 0x30
      12'hC72: dout <= 8'b00001000; // 3186 :   8 - 0x8
      12'hC73: dout <= 8'b01000100; // 3187 :  68 - 0x44
      12'hC74: dout <= 8'b01100010; // 3188 :  98 - 0x62
      12'hC75: dout <= 8'b01100010; // 3189 :  98 - 0x62
      12'hC76: dout <= 8'b00000001; // 3190 :   1 - 0x1
      12'hC77: dout <= 8'b00111111; // 3191 :  63 - 0x3f
      12'hC78: dout <= 8'b10001011; // 3192 : 139 - 0x8b -- Background 0x8f
      12'hC79: dout <= 8'b11000001; // 3193 : 193 - 0xc1
      12'hC7A: dout <= 8'b11111110; // 3194 : 254 - 0xfe
      12'hC7B: dout <= 8'b11111100; // 3195 : 252 - 0xfc
      12'hC7C: dout <= 8'b11110000; // 3196 : 240 - 0xf0
      12'hC7D: dout <= 8'b11110000; // 3197 : 240 - 0xf0
      12'hC7E: dout <= 8'b11111000; // 3198 : 248 - 0xf8
      12'hC7F: dout <= 8'b11110000; // 3199 : 240 - 0xf0
      12'hC80: dout <= 8'b00000011; // 3200 :   3 - 0x3 -- Background 0x90
      12'hC81: dout <= 8'b00001110; // 3201 :  14 - 0xe
      12'hC82: dout <= 8'b00010110; // 3202 :  22 - 0x16
      12'hC83: dout <= 8'b00100110; // 3203 :  38 - 0x26
      12'hC84: dout <= 8'b01100011; // 3204 :  99 - 0x63
      12'hC85: dout <= 8'b01110010; // 3205 : 114 - 0x72
      12'hC86: dout <= 8'b01110000; // 3206 : 112 - 0x70
      12'hC87: dout <= 8'b11010000; // 3207 : 208 - 0xd0
      12'hC88: dout <= 8'b10101010; // 3208 : 170 - 0xaa -- Background 0x91
      12'hC89: dout <= 8'b11111111; // 3209 : 255 - 0xff
      12'hC8A: dout <= 8'b01111111; // 3210 : 127 - 0x7f
      12'hC8B: dout <= 8'b00111100; // 3211 :  60 - 0x3c
      12'hC8C: dout <= 8'b00011100; // 3212 :  28 - 0x1c
      12'hC8D: dout <= 8'b00000100; // 3213 :   4 - 0x4
      12'hC8E: dout <= 8'b00000010; // 3214 :   2 - 0x2
      12'hC8F: dout <= 8'b00000001; // 3215 :   1 - 0x1
      12'hC90: dout <= 8'b11000000; // 3216 : 192 - 0xc0 -- Background 0x92
      12'hC91: dout <= 8'b00110000; // 3217 :  48 - 0x30
      12'hC92: dout <= 8'b00001000; // 3218 :   8 - 0x8
      12'hC93: dout <= 8'b00100100; // 3219 :  36 - 0x24
      12'hC94: dout <= 8'b00110010; // 3220 :  50 - 0x32
      12'hC95: dout <= 8'b00110010; // 3221 :  50 - 0x32
      12'hC96: dout <= 8'b00000001; // 3222 :   1 - 0x1
      12'hC97: dout <= 8'b00011111; // 3223 :  31 - 0x1f
      12'hC98: dout <= 8'b10001011; // 3224 : 139 - 0x8b -- Background 0x93
      12'hC99: dout <= 8'b11000001; // 3225 : 193 - 0xc1
      12'hC9A: dout <= 8'b11111110; // 3226 : 254 - 0xfe
      12'hC9B: dout <= 8'b11111100; // 3227 : 252 - 0xfc
      12'hC9C: dout <= 8'b11110000; // 3228 : 240 - 0xf0
      12'hC9D: dout <= 8'b11000000; // 3229 : 192 - 0xc0
      12'hC9E: dout <= 8'b00100000; // 3230 :  32 - 0x20
      12'hC9F: dout <= 8'b11100000; // 3231 : 224 - 0xe0
      12'hCA0: dout <= 8'b00000011; // 3232 :   3 - 0x3 -- Background 0x94
      12'hCA1: dout <= 8'b00001111; // 3233 :  15 - 0xf
      12'hCA2: dout <= 8'b00010011; // 3234 :  19 - 0x13
      12'hCA3: dout <= 8'b00110001; // 3235 :  49 - 0x31
      12'hCA4: dout <= 8'b01111001; // 3236 : 121 - 0x79
      12'hCA5: dout <= 8'b01011001; // 3237 :  89 - 0x59
      12'hCA6: dout <= 8'b01001000; // 3238 :  72 - 0x48
      12'hCA7: dout <= 8'b11001100; // 3239 : 204 - 0xcc
      12'hCA8: dout <= 8'b10010101; // 3240 : 149 - 0x95 -- Background 0x95
      12'hCA9: dout <= 8'b11111111; // 3241 : 255 - 0xff
      12'hCAA: dout <= 8'b01111111; // 3242 : 127 - 0x7f
      12'hCAB: dout <= 8'b00111110; // 3243 :  62 - 0x3e
      12'hCAC: dout <= 8'b00011111; // 3244 :  31 - 0x1f
      12'hCAD: dout <= 8'b00001111; // 3245 :  15 - 0xf
      12'hCAE: dout <= 8'b00001111; // 3246 :  15 - 0xf
      12'hCAF: dout <= 8'b00000111; // 3247 :   7 - 0x7
      12'hCB0: dout <= 8'b11000000; // 3248 : 192 - 0xc0 -- Background 0x96
      12'hCB1: dout <= 8'b00110000; // 3249 :  48 - 0x30
      12'hCB2: dout <= 8'b00001000; // 3250 :   8 - 0x8
      12'hCB3: dout <= 8'b10010100; // 3251 : 148 - 0x94
      12'hCB4: dout <= 8'b10011010; // 3252 : 154 - 0x9a
      12'hCB5: dout <= 8'b00011010; // 3253 :  26 - 0x1a
      12'hCB6: dout <= 8'b00000001; // 3254 :   1 - 0x1
      12'hCB7: dout <= 8'b00001111; // 3255 :  15 - 0xf
      12'hCB8: dout <= 8'b01000101; // 3256 :  69 - 0x45 -- Background 0x97
      12'hCB9: dout <= 8'b11100001; // 3257 : 225 - 0xe1
      12'hCBA: dout <= 8'b11111110; // 3258 : 254 - 0xfe
      12'hCBB: dout <= 8'b01111100; // 3259 : 124 - 0x7c
      12'hCBC: dout <= 8'b00110000; // 3260 :  48 - 0x30
      12'hCBD: dout <= 8'b00110000; // 3261 :  48 - 0x30
      12'hCBE: dout <= 8'b10001000; // 3262 : 136 - 0x88
      12'hCBF: dout <= 8'b01111000; // 3263 : 120 - 0x78
      12'hCC0: dout <= 8'b00000001; // 3264 :   1 - 0x1 -- Background 0x98
      12'hCC1: dout <= 8'b00000000; // 3265 :   0 - 0x0
      12'hCC2: dout <= 8'b00000000; // 3266 :   0 - 0x0
      12'hCC3: dout <= 8'b00000000; // 3267 :   0 - 0x0
      12'hCC4: dout <= 8'b00000001; // 3268 :   1 - 0x1
      12'hCC5: dout <= 8'b00000001; // 3269 :   1 - 0x1
      12'hCC6: dout <= 8'b00000010; // 3270 :   2 - 0x2
      12'hCC7: dout <= 8'b00000110; // 3271 :   6 - 0x6
      12'hCC8: dout <= 8'b01111000; // 3272 : 120 - 0x78 -- Background 0x99
      12'hCC9: dout <= 8'b00101010; // 3273 :  42 - 0x2a
      12'hCCA: dout <= 8'b01010100; // 3274 :  84 - 0x54
      12'hCCB: dout <= 8'b00101001; // 3275 :  41 - 0x29
      12'hCCC: dout <= 8'b00101111; // 3276 :  47 - 0x2f
      12'hCCD: dout <= 8'b00110111; // 3277 :  55 - 0x37
      12'hCCE: dout <= 8'b00000011; // 3278 :   3 - 0x3
      12'hCCF: dout <= 8'b00000111; // 3279 :   7 - 0x7
      12'hCD0: dout <= 8'b10110000; // 3280 : 176 - 0xb0 -- Background 0x9a
      12'hCD1: dout <= 8'b11101000; // 3281 : 232 - 0xe8
      12'hCD2: dout <= 8'b10001100; // 3282 : 140 - 0x8c
      12'hCD3: dout <= 8'b10011110; // 3283 : 158 - 0x9e
      12'hCD4: dout <= 8'b00011111; // 3284 :  31 - 0x1f
      12'hCD5: dout <= 8'b00001111; // 3285 :  15 - 0xf
      12'hCD6: dout <= 8'b10010110; // 3286 : 150 - 0x96
      12'hCD7: dout <= 8'b00011100; // 3287 :  28 - 0x1c
      12'hCD8: dout <= 8'b00001100; // 3288 :  12 - 0xc -- Background 0x9b
      12'hCD9: dout <= 8'b00111000; // 3289 :  56 - 0x38
      12'hCDA: dout <= 8'b11101000; // 3290 : 232 - 0xe8
      12'hCDB: dout <= 8'b11010000; // 3291 : 208 - 0xd0
      12'hCDC: dout <= 8'b11100000; // 3292 : 224 - 0xe0
      12'hCDD: dout <= 8'b10000000; // 3293 : 128 - 0x80
      12'hCDE: dout <= 8'b00000000; // 3294 :   0 - 0x0
      12'hCDF: dout <= 8'b10000000; // 3295 : 128 - 0x80
      12'hCE0: dout <= 8'b00000001; // 3296 :   1 - 0x1 -- Background 0x9c
      12'hCE1: dout <= 8'b00000000; // 3297 :   0 - 0x0
      12'hCE2: dout <= 8'b00000000; // 3298 :   0 - 0x0
      12'hCE3: dout <= 8'b00000000; // 3299 :   0 - 0x0
      12'hCE4: dout <= 8'b00000001; // 3300 :   1 - 0x1
      12'hCE5: dout <= 8'b00000001; // 3301 :   1 - 0x1
      12'hCE6: dout <= 8'b00000010; // 3302 :   2 - 0x2
      12'hCE7: dout <= 8'b00000110; // 3303 :   6 - 0x6
      12'hCE8: dout <= 8'b01111000; // 3304 : 120 - 0x78 -- Background 0x9d
      12'hCE9: dout <= 8'b00101010; // 3305 :  42 - 0x2a
      12'hCEA: dout <= 8'b01010100; // 3306 :  84 - 0x54
      12'hCEB: dout <= 8'b00101001; // 3307 :  41 - 0x29
      12'hCEC: dout <= 8'b00101111; // 3308 :  47 - 0x2f
      12'hCED: dout <= 8'b00111100; // 3309 :  60 - 0x3c
      12'hCEE: dout <= 8'b00011110; // 3310 :  30 - 0x1e
      12'hCEF: dout <= 8'b00000000; // 3311 :   0 - 0x0
      12'hCF0: dout <= 8'b10110000; // 3312 : 176 - 0xb0 -- Background 0x9e
      12'hCF1: dout <= 8'b11101000; // 3313 : 232 - 0xe8
      12'hCF2: dout <= 8'b10001100; // 3314 : 140 - 0x8c
      12'hCF3: dout <= 8'b10011110; // 3315 : 158 - 0x9e
      12'hCF4: dout <= 8'b00011111; // 3316 :  31 - 0x1f
      12'hCF5: dout <= 8'b00001111; // 3317 :  15 - 0xf
      12'hCF6: dout <= 8'b10010110; // 3318 : 150 - 0x96
      12'hCF7: dout <= 8'b00011100; // 3319 :  28 - 0x1c
      12'hCF8: dout <= 8'b00001100; // 3320 :  12 - 0xc -- Background 0x9f
      12'hCF9: dout <= 8'b00111000; // 3321 :  56 - 0x38
      12'hCFA: dout <= 8'b11101000; // 3322 : 232 - 0xe8
      12'hCFB: dout <= 8'b11110000; // 3323 : 240 - 0xf0
      12'hCFC: dout <= 8'b11000000; // 3324 : 192 - 0xc0
      12'hCFD: dout <= 8'b01110000; // 3325 : 112 - 0x70
      12'hCFE: dout <= 8'b11000000; // 3326 : 192 - 0xc0
      12'hCFF: dout <= 8'b00000000; // 3327 :   0 - 0x0
      12'hD00: dout <= 8'b00000011; // 3328 :   3 - 0x3 -- Background 0xa0
      12'hD01: dout <= 8'b00001111; // 3329 :  15 - 0xf
      12'hD02: dout <= 8'b00011100; // 3330 :  28 - 0x1c
      12'hD03: dout <= 8'b00110000; // 3331 :  48 - 0x30
      12'hD04: dout <= 8'b01100000; // 3332 :  96 - 0x60
      12'hD05: dout <= 8'b01100000; // 3333 :  96 - 0x60
      12'hD06: dout <= 8'b11000000; // 3334 : 192 - 0xc0
      12'hD07: dout <= 8'b11000000; // 3335 : 192 - 0xc0
      12'hD08: dout <= 8'b11000000; // 3336 : 192 - 0xc0 -- Background 0xa1
      12'hD09: dout <= 8'b11000000; // 3337 : 192 - 0xc0
      12'hD0A: dout <= 8'b01100000; // 3338 :  96 - 0x60
      12'hD0B: dout <= 8'b01100000; // 3339 :  96 - 0x60
      12'hD0C: dout <= 8'b00110000; // 3340 :  48 - 0x30
      12'hD0D: dout <= 8'b00011010; // 3341 :  26 - 0x1a
      12'hD0E: dout <= 8'b00001101; // 3342 :  13 - 0xd
      12'hD0F: dout <= 8'b00000011; // 3343 :   3 - 0x3
      12'hD10: dout <= 8'b11000000; // 3344 : 192 - 0xc0 -- Background 0xa2
      12'hD11: dout <= 8'b11110000; // 3345 : 240 - 0xf0
      12'hD12: dout <= 8'b00111000; // 3346 :  56 - 0x38
      12'hD13: dout <= 8'b00001100; // 3347 :  12 - 0xc
      12'hD14: dout <= 8'b00000110; // 3348 :   6 - 0x6
      12'hD15: dout <= 8'b00000010; // 3349 :   2 - 0x2
      12'hD16: dout <= 8'b00000101; // 3350 :   5 - 0x5
      12'hD17: dout <= 8'b00000011; // 3351 :   3 - 0x3
      12'hD18: dout <= 8'b00000101; // 3352 :   5 - 0x5 -- Background 0xa3
      12'hD19: dout <= 8'b00001011; // 3353 :  11 - 0xb
      12'hD1A: dout <= 8'b00010110; // 3354 :  22 - 0x16
      12'hD1B: dout <= 8'b00101010; // 3355 :  42 - 0x2a
      12'hD1C: dout <= 8'b01010100; // 3356 :  84 - 0x54
      12'hD1D: dout <= 8'b10101000; // 3357 : 168 - 0xa8
      12'hD1E: dout <= 8'b01110000; // 3358 : 112 - 0x70
      12'hD1F: dout <= 8'b11000000; // 3359 : 192 - 0xc0
      12'hD20: dout <= 8'b00000000; // 3360 :   0 - 0x0 -- Background 0xa4
      12'hD21: dout <= 8'b00001111; // 3361 :  15 - 0xf
      12'hD22: dout <= 8'b00011111; // 3362 :  31 - 0x1f
      12'hD23: dout <= 8'b00110001; // 3363 :  49 - 0x31
      12'hD24: dout <= 8'b00111111; // 3364 :  63 - 0x3f
      12'hD25: dout <= 8'b01111111; // 3365 : 127 - 0x7f
      12'hD26: dout <= 8'b11111111; // 3366 : 255 - 0xff
      12'hD27: dout <= 8'b11011111; // 3367 : 223 - 0xdf
      12'hD28: dout <= 8'b11000000; // 3368 : 192 - 0xc0 -- Background 0xa5
      12'hD29: dout <= 8'b11000111; // 3369 : 199 - 0xc7
      12'hD2A: dout <= 8'b01101111; // 3370 : 111 - 0x6f
      12'hD2B: dout <= 8'b01100111; // 3371 : 103 - 0x67
      12'hD2C: dout <= 8'b01100011; // 3372 :  99 - 0x63
      12'hD2D: dout <= 8'b00110000; // 3373 :  48 - 0x30
      12'hD2E: dout <= 8'b00011000; // 3374 :  24 - 0x18
      12'hD2F: dout <= 8'b00000111; // 3375 :   7 - 0x7
      12'hD30: dout <= 8'b00000000; // 3376 :   0 - 0x0 -- Background 0xa6
      12'hD31: dout <= 8'b11110000; // 3377 : 240 - 0xf0
      12'hD32: dout <= 8'b11111000; // 3378 : 248 - 0xf8
      12'hD33: dout <= 8'b10001100; // 3379 : 140 - 0x8c
      12'hD34: dout <= 8'b11111100; // 3380 : 252 - 0xfc
      12'hD35: dout <= 8'b11111110; // 3381 : 254 - 0xfe
      12'hD36: dout <= 8'b11111101; // 3382 : 253 - 0xfd
      12'hD37: dout <= 8'b11111001; // 3383 : 249 - 0xf9
      12'hD38: dout <= 8'b00000011; // 3384 :   3 - 0x3 -- Background 0xa7
      12'hD39: dout <= 8'b11100101; // 3385 : 229 - 0xe5
      12'hD3A: dout <= 8'b11110010; // 3386 : 242 - 0xf2
      12'hD3B: dout <= 8'b11100110; // 3387 : 230 - 0xe6
      12'hD3C: dout <= 8'b11001010; // 3388 : 202 - 0xca
      12'hD3D: dout <= 8'b00010100; // 3389 :  20 - 0x14
      12'hD3E: dout <= 8'b00111000; // 3390 :  56 - 0x38
      12'hD3F: dout <= 8'b11100000; // 3391 : 224 - 0xe0
      12'hD40: dout <= 8'b00000000; // 3392 :   0 - 0x0 -- Background 0xa8
      12'hD41: dout <= 8'b00001111; // 3393 :  15 - 0xf
      12'hD42: dout <= 8'b00011111; // 3394 :  31 - 0x1f
      12'hD43: dout <= 8'b00110001; // 3395 :  49 - 0x31
      12'hD44: dout <= 8'b00111111; // 3396 :  63 - 0x3f
      12'hD45: dout <= 8'b01111111; // 3397 : 127 - 0x7f
      12'hD46: dout <= 8'b11111111; // 3398 : 255 - 0xff
      12'hD47: dout <= 8'b11011111; // 3399 : 223 - 0xdf
      12'hD48: dout <= 8'b11000000; // 3400 : 192 - 0xc0 -- Background 0xa9
      12'hD49: dout <= 8'b11000011; // 3401 : 195 - 0xc3
      12'hD4A: dout <= 8'b11000111; // 3402 : 199 - 0xc7
      12'hD4B: dout <= 8'b11001111; // 3403 : 207 - 0xcf
      12'hD4C: dout <= 8'b11000111; // 3404 : 199 - 0xc7
      12'hD4D: dout <= 8'b11000000; // 3405 : 192 - 0xc0
      12'hD4E: dout <= 8'b11100000; // 3406 : 224 - 0xe0
      12'hD4F: dout <= 8'b11111111; // 3407 : 255 - 0xff
      12'hD50: dout <= 8'b00000000; // 3408 :   0 - 0x0 -- Background 0xaa
      12'hD51: dout <= 8'b11110000; // 3409 : 240 - 0xf0
      12'hD52: dout <= 8'b11111000; // 3410 : 248 - 0xf8
      12'hD53: dout <= 8'b10001100; // 3411 : 140 - 0x8c
      12'hD54: dout <= 8'b11111100; // 3412 : 252 - 0xfc
      12'hD55: dout <= 8'b11111110; // 3413 : 254 - 0xfe
      12'hD56: dout <= 8'b11111101; // 3414 : 253 - 0xfd
      12'hD57: dout <= 8'b11111001; // 3415 : 249 - 0xf9
      12'hD58: dout <= 8'b00000011; // 3416 :   3 - 0x3 -- Background 0xab
      12'hD59: dout <= 8'b11000101; // 3417 : 197 - 0xc5
      12'hD5A: dout <= 8'b11100011; // 3418 : 227 - 0xe3
      12'hD5B: dout <= 8'b11110101; // 3419 : 245 - 0xf5
      12'hD5C: dout <= 8'b11100011; // 3420 : 227 - 0xe3
      12'hD5D: dout <= 8'b00000101; // 3421 :   5 - 0x5
      12'hD5E: dout <= 8'b00001011; // 3422 :  11 - 0xb
      12'hD5F: dout <= 8'b11111111; // 3423 : 255 - 0xff
      12'hD60: dout <= 8'b10000011; // 3424 : 131 - 0x83 -- Background 0xac
      12'hD61: dout <= 8'b10001100; // 3425 : 140 - 0x8c
      12'hD62: dout <= 8'b10010000; // 3426 : 144 - 0x90
      12'hD63: dout <= 8'b10010000; // 3427 : 144 - 0x90
      12'hD64: dout <= 8'b11100000; // 3428 : 224 - 0xe0
      12'hD65: dout <= 8'b10100000; // 3429 : 160 - 0xa0
      12'hD66: dout <= 8'b10101111; // 3430 : 175 - 0xaf
      12'hD67: dout <= 8'b01101111; // 3431 : 111 - 0x6f
      12'hD68: dout <= 8'b11111011; // 3432 : 251 - 0xfb -- Background 0xad
      12'hD69: dout <= 8'b00000101; // 3433 :   5 - 0x5
      12'hD6A: dout <= 8'b00000101; // 3434 :   5 - 0x5
      12'hD6B: dout <= 8'b00000101; // 3435 :   5 - 0x5
      12'hD6C: dout <= 8'b01000101; // 3436 :  69 - 0x45
      12'hD6D: dout <= 8'b01100101; // 3437 : 101 - 0x65
      12'hD6E: dout <= 8'b11110101; // 3438 : 245 - 0xf5
      12'hD6F: dout <= 8'b11111101; // 3439 : 253 - 0xfd
      12'hD70: dout <= 8'b10000011; // 3440 : 131 - 0x83 -- Background 0xae
      12'hD71: dout <= 8'b10001100; // 3441 : 140 - 0x8c
      12'hD72: dout <= 8'b10010000; // 3442 : 144 - 0x90
      12'hD73: dout <= 8'b10010000; // 3443 : 144 - 0x90
      12'hD74: dout <= 8'b11100000; // 3444 : 224 - 0xe0
      12'hD75: dout <= 8'b10100000; // 3445 : 160 - 0xa0
      12'hD76: dout <= 8'b10101111; // 3446 : 175 - 0xaf
      12'hD77: dout <= 8'b01101111; // 3447 : 111 - 0x6f
      12'hD78: dout <= 8'b11111011; // 3448 : 251 - 0xfb -- Background 0xaf
      12'hD79: dout <= 8'b00000101; // 3449 :   5 - 0x5
      12'hD7A: dout <= 8'b00000101; // 3450 :   5 - 0x5
      12'hD7B: dout <= 8'b00000101; // 3451 :   5 - 0x5
      12'hD7C: dout <= 8'b11000101; // 3452 : 197 - 0xc5
      12'hD7D: dout <= 8'b11100101; // 3453 : 229 - 0xe5
      12'hD7E: dout <= 8'b11110101; // 3454 : 245 - 0xf5
      12'hD7F: dout <= 8'b11111101; // 3455 : 253 - 0xfd
      12'hD80: dout <= 8'b00000000; // 3456 :   0 - 0x0 -- Background 0xb0
      12'hD81: dout <= 8'b00000011; // 3457 :   3 - 0x3
      12'hD82: dout <= 8'b00001111; // 3458 :  15 - 0xf
      12'hD83: dout <= 8'b00111111; // 3459 :  63 - 0x3f
      12'hD84: dout <= 8'b01111111; // 3460 : 127 - 0x7f
      12'hD85: dout <= 8'b01111111; // 3461 : 127 - 0x7f
      12'hD86: dout <= 8'b11111111; // 3462 : 255 - 0xff
      12'hD87: dout <= 8'b11111111; // 3463 : 255 - 0xff
      12'hD88: dout <= 8'b11111111; // 3464 : 255 - 0xff -- Background 0xb1
      12'hD89: dout <= 8'b10001111; // 3465 : 143 - 0x8f
      12'hD8A: dout <= 8'b10000000; // 3466 : 128 - 0x80
      12'hD8B: dout <= 8'b11110000; // 3467 : 240 - 0xf0
      12'hD8C: dout <= 8'b11111111; // 3468 : 255 - 0xff
      12'hD8D: dout <= 8'b11111111; // 3469 : 255 - 0xff
      12'hD8E: dout <= 8'b01111111; // 3470 : 127 - 0x7f
      12'hD8F: dout <= 8'b00001111; // 3471 :  15 - 0xf
      12'hD90: dout <= 8'b00000000; // 3472 :   0 - 0x0 -- Background 0xb2
      12'hD91: dout <= 8'b11000000; // 3473 : 192 - 0xc0
      12'hD92: dout <= 8'b11110000; // 3474 : 240 - 0xf0
      12'hD93: dout <= 8'b11111100; // 3475 : 252 - 0xfc
      12'hD94: dout <= 8'b11111110; // 3476 : 254 - 0xfe
      12'hD95: dout <= 8'b11111110; // 3477 : 254 - 0xfe
      12'hD96: dout <= 8'b11111111; // 3478 : 255 - 0xff
      12'hD97: dout <= 8'b11111111; // 3479 : 255 - 0xff
      12'hD98: dout <= 8'b11111111; // 3480 : 255 - 0xff -- Background 0xb3
      12'hD99: dout <= 8'b11110001; // 3481 : 241 - 0xf1
      12'hD9A: dout <= 8'b00000001; // 3482 :   1 - 0x1
      12'hD9B: dout <= 8'b00001111; // 3483 :  15 - 0xf
      12'hD9C: dout <= 8'b11111111; // 3484 : 255 - 0xff
      12'hD9D: dout <= 8'b11111111; // 3485 : 255 - 0xff
      12'hD9E: dout <= 8'b11111110; // 3486 : 254 - 0xfe
      12'hD9F: dout <= 8'b11110000; // 3487 : 240 - 0xf0
      12'hDA0: dout <= 8'b00000000; // 3488 :   0 - 0x0 -- Background 0xb4
      12'hDA1: dout <= 8'b00000011; // 3489 :   3 - 0x3
      12'hDA2: dout <= 8'b00001110; // 3490 :  14 - 0xe
      12'hDA3: dout <= 8'b00110101; // 3491 :  53 - 0x35
      12'hDA4: dout <= 8'b01101110; // 3492 : 110 - 0x6e
      12'hDA5: dout <= 8'b01010101; // 3493 :  85 - 0x55
      12'hDA6: dout <= 8'b10111010; // 3494 : 186 - 0xba
      12'hDA7: dout <= 8'b11010111; // 3495 : 215 - 0xd7
      12'hDA8: dout <= 8'b11111010; // 3496 : 250 - 0xfa -- Background 0xb5
      12'hDA9: dout <= 8'b10001111; // 3497 : 143 - 0x8f
      12'hDAA: dout <= 8'b10000000; // 3498 : 128 - 0x80
      12'hDAB: dout <= 8'b11110000; // 3499 : 240 - 0xf0
      12'hDAC: dout <= 8'b10101111; // 3500 : 175 - 0xaf
      12'hDAD: dout <= 8'b11010101; // 3501 : 213 - 0xd5
      12'hDAE: dout <= 8'b01111010; // 3502 : 122 - 0x7a
      12'hDAF: dout <= 8'b00001111; // 3503 :  15 - 0xf
      12'hDB0: dout <= 8'b00000000; // 3504 :   0 - 0x0 -- Background 0xb6
      12'hDB1: dout <= 8'b11000000; // 3505 : 192 - 0xc0
      12'hDB2: dout <= 8'b10110000; // 3506 : 176 - 0xb0
      12'hDB3: dout <= 8'b01011100; // 3507 :  92 - 0x5c
      12'hDB4: dout <= 8'b11101010; // 3508 : 234 - 0xea
      12'hDB5: dout <= 8'b01011110; // 3509 :  94 - 0x5e
      12'hDB6: dout <= 8'b10101011; // 3510 : 171 - 0xab
      12'hDB7: dout <= 8'b01110101; // 3511 : 117 - 0x75
      12'hDB8: dout <= 8'b10101111; // 3512 : 175 - 0xaf -- Background 0xb7
      12'hDB9: dout <= 8'b11110001; // 3513 : 241 - 0xf1
      12'hDBA: dout <= 8'b00000001; // 3514 :   1 - 0x1
      12'hDBB: dout <= 8'b00001111; // 3515 :  15 - 0xf
      12'hDBC: dout <= 8'b11111011; // 3516 : 251 - 0xfb
      12'hDBD: dout <= 8'b01010101; // 3517 :  85 - 0x55
      12'hDBE: dout <= 8'b10101110; // 3518 : 174 - 0xae
      12'hDBF: dout <= 8'b11110000; // 3519 : 240 - 0xf0
      12'hDC0: dout <= 8'b00000000; // 3520 :   0 - 0x0 -- Background 0xb8
      12'hDC1: dout <= 8'b00000011; // 3521 :   3 - 0x3
      12'hDC2: dout <= 8'b00001100; // 3522 :  12 - 0xc
      12'hDC3: dout <= 8'b00110000; // 3523 :  48 - 0x30
      12'hDC4: dout <= 8'b01000100; // 3524 :  68 - 0x44
      12'hDC5: dout <= 8'b01000000; // 3525 :  64 - 0x40
      12'hDC6: dout <= 8'b10010000; // 3526 : 144 - 0x90
      12'hDC7: dout <= 8'b10000010; // 3527 : 130 - 0x82
      12'hDC8: dout <= 8'b11110000; // 3528 : 240 - 0xf0 -- Background 0xb9
      12'hDC9: dout <= 8'b11111111; // 3529 : 255 - 0xff
      12'hDCA: dout <= 8'b11111111; // 3530 : 255 - 0xff
      12'hDCB: dout <= 8'b11111111; // 3531 : 255 - 0xff
      12'hDCC: dout <= 8'b10001111; // 3532 : 143 - 0x8f
      12'hDCD: dout <= 8'b10000000; // 3533 : 128 - 0x80
      12'hDCE: dout <= 8'b01110000; // 3534 : 112 - 0x70
      12'hDCF: dout <= 8'b00001111; // 3535 :  15 - 0xf
      12'hDD0: dout <= 8'b00000000; // 3536 :   0 - 0x0 -- Background 0xba
      12'hDD1: dout <= 8'b11000000; // 3537 : 192 - 0xc0
      12'hDD2: dout <= 8'b00110000; // 3538 :  48 - 0x30
      12'hDD3: dout <= 8'b00001100; // 3539 :  12 - 0xc
      12'hDD4: dout <= 8'b01000010; // 3540 :  66 - 0x42
      12'hDD5: dout <= 8'b00001010; // 3541 :  10 - 0xa
      12'hDD6: dout <= 8'b00000001; // 3542 :   1 - 0x1
      12'hDD7: dout <= 8'b00100001; // 3543 :  33 - 0x21
      12'hDD8: dout <= 8'b00001111; // 3544 :  15 - 0xf -- Background 0xbb
      12'hDD9: dout <= 8'b11111111; // 3545 : 255 - 0xff
      12'hDDA: dout <= 8'b11111111; // 3546 : 255 - 0xff
      12'hDDB: dout <= 8'b11111111; // 3547 : 255 - 0xff
      12'hDDC: dout <= 8'b11110001; // 3548 : 241 - 0xf1
      12'hDDD: dout <= 8'b00000001; // 3549 :   1 - 0x1
      12'hDDE: dout <= 8'b00001110; // 3550 :  14 - 0xe
      12'hDDF: dout <= 8'b11110000; // 3551 : 240 - 0xf0
      12'hDE0: dout <= 8'b11110011; // 3552 : 243 - 0xf3 -- Background 0xbc
      12'hDE1: dout <= 8'b11111111; // 3553 : 255 - 0xff
      12'hDE2: dout <= 8'b11000100; // 3554 : 196 - 0xc4
      12'hDE3: dout <= 8'b11000000; // 3555 : 192 - 0xc0
      12'hDE4: dout <= 8'b01000000; // 3556 :  64 - 0x40
      12'hDE5: dout <= 8'b01100011; // 3557 :  99 - 0x63
      12'hDE6: dout <= 8'b11000111; // 3558 : 199 - 0xc7
      12'hDE7: dout <= 8'b11000110; // 3559 : 198 - 0xc6
      12'hDE8: dout <= 8'b11000110; // 3560 : 198 - 0xc6 -- Background 0xbd
      12'hDE9: dout <= 8'b11000110; // 3561 : 198 - 0xc6
      12'hDEA: dout <= 8'b01100011; // 3562 :  99 - 0x63
      12'hDEB: dout <= 8'b01000000; // 3563 :  64 - 0x40
      12'hDEC: dout <= 8'b11000000; // 3564 : 192 - 0xc0
      12'hDED: dout <= 8'b11000100; // 3565 : 196 - 0xc4
      12'hDEE: dout <= 8'b11001100; // 3566 : 204 - 0xcc
      12'hDEF: dout <= 8'b11110011; // 3567 : 243 - 0xf3
      12'hDF0: dout <= 8'b11001111; // 3568 : 207 - 0xcf -- Background 0xbe
      12'hDF1: dout <= 8'b11111111; // 3569 : 255 - 0xff
      12'hDF2: dout <= 8'b00100001; // 3570 :  33 - 0x21
      12'hDF3: dout <= 8'b00000001; // 3571 :   1 - 0x1
      12'hDF4: dout <= 8'b00000010; // 3572 :   2 - 0x2
      12'hDF5: dout <= 8'b11000110; // 3573 : 198 - 0xc6
      12'hDF6: dout <= 8'b11100001; // 3574 : 225 - 0xe1
      12'hDF7: dout <= 8'b00100001; // 3575 :  33 - 0x21
      12'hDF8: dout <= 8'b00100001; // 3576 :  33 - 0x21 -- Background 0xbf
      12'hDF9: dout <= 8'b00100001; // 3577 :  33 - 0x21
      12'hDFA: dout <= 8'b11000110; // 3578 : 198 - 0xc6
      12'hDFB: dout <= 8'b00000010; // 3579 :   2 - 0x2
      12'hDFC: dout <= 8'b00000001; // 3580 :   1 - 0x1
      12'hDFD: dout <= 8'b00100001; // 3581 :  33 - 0x21
      12'hDFE: dout <= 8'b00110001; // 3582 :  49 - 0x31
      12'hDFF: dout <= 8'b11001111; // 3583 : 207 - 0xcf
      12'hE00: dout <= 8'b00000000; // 3584 :   0 - 0x0 -- Background 0xc0
      12'hE01: dout <= 8'b01010000; // 3585 :  80 - 0x50
      12'hE02: dout <= 8'b10110011; // 3586 : 179 - 0xb3
      12'hE03: dout <= 8'b10010111; // 3587 : 151 - 0x97
      12'hE04: dout <= 8'b10011111; // 3588 : 159 - 0x9f
      12'hE05: dout <= 8'b01101111; // 3589 : 111 - 0x6f
      12'hE06: dout <= 8'b00011111; // 3590 :  31 - 0x1f
      12'hE07: dout <= 8'b00011111; // 3591 :  31 - 0x1f
      12'hE08: dout <= 8'b00011111; // 3592 :  31 - 0x1f -- Background 0xc1
      12'hE09: dout <= 8'b00011111; // 3593 :  31 - 0x1f
      12'hE0A: dout <= 8'b00001111; // 3594 :  15 - 0xf
      12'hE0B: dout <= 8'b00000111; // 3595 :   7 - 0x7
      12'hE0C: dout <= 8'b00011101; // 3596 :  29 - 0x1d
      12'hE0D: dout <= 8'b00101100; // 3597 :  44 - 0x2c
      12'hE0E: dout <= 8'b01010100; // 3598 :  84 - 0x54
      12'hE0F: dout <= 8'b01111100; // 3599 : 124 - 0x7c
      12'hE10: dout <= 8'b00000000; // 3600 :   0 - 0x0 -- Background 0xc2
      12'hE11: dout <= 8'b00001010; // 3601 :  10 - 0xa
      12'hE12: dout <= 8'b11001101; // 3602 : 205 - 0xcd
      12'hE13: dout <= 8'b11101001; // 3603 : 233 - 0xe9
      12'hE14: dout <= 8'b11111001; // 3604 : 249 - 0xf9
      12'hE15: dout <= 8'b11110110; // 3605 : 246 - 0xf6
      12'hE16: dout <= 8'b11110000; // 3606 : 240 - 0xf0
      12'hE17: dout <= 8'b11111000; // 3607 : 248 - 0xf8
      12'hE18: dout <= 8'b11111000; // 3608 : 248 - 0xf8 -- Background 0xc3
      12'hE19: dout <= 8'b11111000; // 3609 : 248 - 0xf8
      12'hE1A: dout <= 8'b11110000; // 3610 : 240 - 0xf0
      12'hE1B: dout <= 8'b11000000; // 3611 : 192 - 0xc0
      12'hE1C: dout <= 8'b10111000; // 3612 : 184 - 0xb8
      12'hE1D: dout <= 8'b00110100; // 3613 :  52 - 0x34
      12'hE1E: dout <= 8'b00101010; // 3614 :  42 - 0x2a
      12'hE1F: dout <= 8'b00111110; // 3615 :  62 - 0x3e
      12'hE20: dout <= 8'b00000101; // 3616 :   5 - 0x5 -- Background 0xc4
      12'hE21: dout <= 8'b00001010; // 3617 :  10 - 0xa
      12'hE22: dout <= 8'b00001000; // 3618 :   8 - 0x8
      12'hE23: dout <= 8'b00001111; // 3619 :  15 - 0xf
      12'hE24: dout <= 8'b00000001; // 3620 :   1 - 0x1
      12'hE25: dout <= 8'b00000011; // 3621 :   3 - 0x3
      12'hE26: dout <= 8'b00000111; // 3622 :   7 - 0x7
      12'hE27: dout <= 8'b00001111; // 3623 :  15 - 0xf
      12'hE28: dout <= 8'b00001111; // 3624 :  15 - 0xf -- Background 0xc5
      12'hE29: dout <= 8'b11101111; // 3625 : 239 - 0xef
      12'hE2A: dout <= 8'b11011111; // 3626 : 223 - 0xdf
      12'hE2B: dout <= 8'b10101111; // 3627 : 175 - 0xaf
      12'hE2C: dout <= 8'b01100111; // 3628 : 103 - 0x67
      12'hE2D: dout <= 8'b00001101; // 3629 :  13 - 0xd
      12'hE2E: dout <= 8'b00001010; // 3630 :  10 - 0xa
      12'hE2F: dout <= 8'b00000111; // 3631 :   7 - 0x7
      12'hE30: dout <= 8'b00000000; // 3632 :   0 - 0x0 -- Background 0xc6
      12'hE31: dout <= 8'b10000000; // 3633 : 128 - 0x80
      12'hE32: dout <= 8'b10000000; // 3634 : 128 - 0x80
      12'hE33: dout <= 8'b11110000; // 3635 : 240 - 0xf0
      12'hE34: dout <= 8'b11111000; // 3636 : 248 - 0xf8
      12'hE35: dout <= 8'b11111100; // 3637 : 252 - 0xfc
      12'hE36: dout <= 8'b11111100; // 3638 : 252 - 0xfc
      12'hE37: dout <= 8'b11111100; // 3639 : 252 - 0xfc
      12'hE38: dout <= 8'b11111100; // 3640 : 252 - 0xfc -- Background 0xc7
      12'hE39: dout <= 8'b11111110; // 3641 : 254 - 0xfe
      12'hE3A: dout <= 8'b11111001; // 3642 : 249 - 0xf9
      12'hE3B: dout <= 8'b11111010; // 3643 : 250 - 0xfa
      12'hE3C: dout <= 8'b11101001; // 3644 : 233 - 0xe9
      12'hE3D: dout <= 8'b00001110; // 3645 :  14 - 0xe
      12'hE3E: dout <= 8'b10000000; // 3646 : 128 - 0x80
      12'hE3F: dout <= 8'b00000000; // 3647 :   0 - 0x0
      12'hE40: dout <= 8'b00000000; // 3648 :   0 - 0x0 -- Background 0xc8
      12'hE41: dout <= 8'b11000000; // 3649 : 192 - 0xc0
      12'hE42: dout <= 8'b10100000; // 3650 : 160 - 0xa0
      12'hE43: dout <= 8'b11010011; // 3651 : 211 - 0xd3
      12'hE44: dout <= 8'b10110111; // 3652 : 183 - 0xb7
      12'hE45: dout <= 8'b11111111; // 3653 : 255 - 0xff
      12'hE46: dout <= 8'b00001111; // 3654 :  15 - 0xf
      12'hE47: dout <= 8'b00011111; // 3655 :  31 - 0x1f
      12'hE48: dout <= 8'b00011111; // 3656 :  31 - 0x1f -- Background 0xc9
      12'hE49: dout <= 8'b00001111; // 3657 :  15 - 0xf
      12'hE4A: dout <= 8'b11110111; // 3658 : 247 - 0xf7
      12'hE4B: dout <= 8'b10110111; // 3659 : 183 - 0xb7
      12'hE4C: dout <= 8'b11010011; // 3660 : 211 - 0xd3
      12'hE4D: dout <= 8'b10100000; // 3661 : 160 - 0xa0
      12'hE4E: dout <= 8'b11000000; // 3662 : 192 - 0xc0
      12'hE4F: dout <= 8'b00000000; // 3663 :   0 - 0x0
      12'hE50: dout <= 8'b00011100; // 3664 :  28 - 0x1c -- Background 0xca
      12'hE51: dout <= 8'b00100010; // 3665 :  34 - 0x22
      12'hE52: dout <= 8'b00100100; // 3666 :  36 - 0x24
      12'hE53: dout <= 8'b11011110; // 3667 : 222 - 0xde
      12'hE54: dout <= 8'b11110000; // 3668 : 240 - 0xf0
      12'hE55: dout <= 8'b11111000; // 3669 : 248 - 0xf8
      12'hE56: dout <= 8'b11111100; // 3670 : 252 - 0xfc
      12'hE57: dout <= 8'b11111100; // 3671 : 252 - 0xfc
      12'hE58: dout <= 8'b11111100; // 3672 : 252 - 0xfc -- Background 0xcb
      12'hE59: dout <= 8'b11111100; // 3673 : 252 - 0xfc
      12'hE5A: dout <= 8'b11111000; // 3674 : 248 - 0xf8
      12'hE5B: dout <= 8'b11110000; // 3675 : 240 - 0xf0
      12'hE5C: dout <= 8'b10011110; // 3676 : 158 - 0x9e
      12'hE5D: dout <= 8'b00100100; // 3677 :  36 - 0x24
      12'hE5E: dout <= 8'b00100010; // 3678 :  34 - 0x22
      12'hE5F: dout <= 8'b00011100; // 3679 :  28 - 0x1c
      12'hE60: dout <= 8'b00001110; // 3680 :  14 - 0xe -- Background 0xcc
      12'hE61: dout <= 8'b00010110; // 3681 :  22 - 0x16
      12'hE62: dout <= 8'b00011010; // 3682 :  26 - 0x1a
      12'hE63: dout <= 8'b00000100; // 3683 :   4 - 0x4
      12'hE64: dout <= 8'b01101111; // 3684 : 111 - 0x6f
      12'hE65: dout <= 8'b10111111; // 3685 : 191 - 0xbf
      12'hE66: dout <= 8'b11011111; // 3686 : 223 - 0xdf
      12'hE67: dout <= 8'b10111111; // 3687 : 191 - 0xbf
      12'hE68: dout <= 8'b01011111; // 3688 :  95 - 0x5f -- Background 0xcd
      12'hE69: dout <= 8'b00011111; // 3689 :  31 - 0x1f
      12'hE6A: dout <= 8'b00011111; // 3690 :  31 - 0x1f
      12'hE6B: dout <= 8'b00001111; // 3691 :  15 - 0xf
      12'hE6C: dout <= 8'b00111111; // 3692 :  63 - 0x3f
      12'hE6D: dout <= 8'b00100011; // 3693 :  35 - 0x23
      12'hE6E: dout <= 8'b00101010; // 3694 :  42 - 0x2a
      12'hE6F: dout <= 8'b00010100; // 3695 :  20 - 0x14
      12'hE70: dout <= 8'b00000000; // 3696 :   0 - 0x0 -- Background 0xce
      12'hE71: dout <= 8'b00000000; // 3697 :   0 - 0x0
      12'hE72: dout <= 8'b00000000; // 3698 :   0 - 0x0
      12'hE73: dout <= 8'b00000000; // 3699 :   0 - 0x0
      12'hE74: dout <= 8'b10001110; // 3700 : 142 - 0x8e
      12'hE75: dout <= 8'b11001001; // 3701 : 201 - 0xc9
      12'hE76: dout <= 8'b11101010; // 3702 : 234 - 0xea
      12'hE77: dout <= 8'b11111001; // 3703 : 249 - 0xf9
      12'hE78: dout <= 8'b11111110; // 3704 : 254 - 0xfe -- Background 0xcf
      12'hE79: dout <= 8'b11111000; // 3705 : 248 - 0xf8
      12'hE7A: dout <= 8'b11111000; // 3706 : 248 - 0xf8
      12'hE7B: dout <= 8'b11111000; // 3707 : 248 - 0xf8
      12'hE7C: dout <= 8'b11110000; // 3708 : 240 - 0xf0
      12'hE7D: dout <= 8'b11100000; // 3709 : 224 - 0xe0
      12'hE7E: dout <= 8'b00000000; // 3710 :   0 - 0x0
      12'hE7F: dout <= 8'b00000000; // 3711 :   0 - 0x0
      12'hE80: dout <= 8'b00000000; // 3712 :   0 - 0x0 -- Background 0xd0
      12'hE81: dout <= 8'b00000000; // 3713 :   0 - 0x0
      12'hE82: dout <= 8'b00000100; // 3714 :   4 - 0x4
      12'hE83: dout <= 8'b00100110; // 3715 :  38 - 0x26
      12'hE84: dout <= 8'b00101011; // 3716 :  43 - 0x2b
      12'hE85: dout <= 8'b01110001; // 3717 : 113 - 0x71
      12'hE86: dout <= 8'b01000000; // 3718 :  64 - 0x40
      12'hE87: dout <= 8'b01000111; // 3719 :  71 - 0x47
      12'hE88: dout <= 8'b10001111; // 3720 : 143 - 0x8f -- Background 0xd1
      12'hE89: dout <= 8'b10001111; // 3721 : 143 - 0x8f
      12'hE8A: dout <= 8'b01001111; // 3722 :  79 - 0x4f
      12'hE8B: dout <= 8'b01001111; // 3723 :  79 - 0x4f
      12'hE8C: dout <= 8'b00111111; // 3724 :  63 - 0x3f
      12'hE8D: dout <= 8'b00010011; // 3725 :  19 - 0x13
      12'hE8E: dout <= 8'b00010001; // 3726 :  17 - 0x11
      12'hE8F: dout <= 8'b00011111; // 3727 :  31 - 0x1f
      12'hE90: dout <= 8'b00000000; // 3728 :   0 - 0x0 -- Background 0xd2
      12'hE91: dout <= 8'b10000000; // 3729 : 128 - 0x80
      12'hE92: dout <= 8'b11001000; // 3730 : 200 - 0xc8
      12'hE93: dout <= 8'b11010100; // 3731 : 212 - 0xd4
      12'hE94: dout <= 8'b00100100; // 3732 :  36 - 0x24
      12'hE95: dout <= 8'b00000010; // 3733 :   2 - 0x2
      12'hE96: dout <= 8'b00000010; // 3734 :   2 - 0x2
      12'hE97: dout <= 8'b11110010; // 3735 : 242 - 0xf2
      12'hE98: dout <= 8'b11110010; // 3736 : 242 - 0xf2 -- Background 0xd3
      12'hE99: dout <= 8'b11110010; // 3737 : 242 - 0xf2
      12'hE9A: dout <= 8'b11110100; // 3738 : 244 - 0xf4
      12'hE9B: dout <= 8'b11110100; // 3739 : 244 - 0xf4
      12'hE9C: dout <= 8'b11110100; // 3740 : 244 - 0xf4
      12'hE9D: dout <= 8'b11001000; // 3741 : 200 - 0xc8
      12'hE9E: dout <= 8'b01000100; // 3742 :  68 - 0x44
      12'hE9F: dout <= 8'b01111100; // 3743 : 124 - 0x7c
      12'hEA0: dout <= 8'b00000000; // 3744 :   0 - 0x0 -- Background 0xd4
      12'hEA1: dout <= 8'b00000000; // 3745 :   0 - 0x0
      12'hEA2: dout <= 8'b00000000; // 3746 :   0 - 0x0
      12'hEA3: dout <= 8'b00001001; // 3747 :   9 - 0x9
      12'hEA4: dout <= 8'b00011010; // 3748 :  26 - 0x1a
      12'hEA5: dout <= 8'b00010100; // 3749 :  20 - 0x14
      12'hEA6: dout <= 8'b00100000; // 3750 :  32 - 0x20
      12'hEA7: dout <= 8'b01000111; // 3751 :  71 - 0x47
      12'hEA8: dout <= 8'b10001111; // 3752 : 143 - 0x8f -- Background 0xd5
      12'hEA9: dout <= 8'b10001111; // 3753 : 143 - 0x8f
      12'hEAA: dout <= 8'b01001111; // 3754 :  79 - 0x4f
      12'hEAB: dout <= 8'b01001111; // 3755 :  79 - 0x4f
      12'hEAC: dout <= 8'b00111111; // 3756 :  63 - 0x3f
      12'hEAD: dout <= 8'b01000111; // 3757 :  71 - 0x47
      12'hEAE: dout <= 8'b00100010; // 3758 :  34 - 0x22
      12'hEAF: dout <= 8'b00011100; // 3759 :  28 - 0x1c
      12'hEB0: dout <= 8'b00000000; // 3760 :   0 - 0x0 -- Background 0xd6
      12'hEB1: dout <= 8'b01000000; // 3761 :  64 - 0x40
      12'hEB2: dout <= 8'b11000000; // 3762 : 192 - 0xc0
      12'hEB3: dout <= 8'b00101100; // 3763 :  44 - 0x2c
      12'hEB4: dout <= 8'b00110100; // 3764 :  52 - 0x34
      12'hEB5: dout <= 8'b00000100; // 3765 :   4 - 0x4
      12'hEB6: dout <= 8'b00000010; // 3766 :   2 - 0x2
      12'hEB7: dout <= 8'b11110010; // 3767 : 242 - 0xf2
      12'hEB8: dout <= 8'b11110010; // 3768 : 242 - 0xf2 -- Background 0xd7
      12'hEB9: dout <= 8'b11110010; // 3769 : 242 - 0xf2
      12'hEBA: dout <= 8'b11110100; // 3770 : 244 - 0xf4
      12'hEBB: dout <= 8'b11110111; // 3771 : 247 - 0xf7
      12'hEBC: dout <= 8'b11111101; // 3772 : 253 - 0xfd
      12'hEBD: dout <= 8'b11100001; // 3773 : 225 - 0xe1
      12'hEBE: dout <= 8'b00010010; // 3774 :  18 - 0x12
      12'hEBF: dout <= 8'b00001100; // 3775 :  12 - 0xc
      12'hEC0: dout <= 8'b01111000; // 3776 : 120 - 0x78 -- Background 0xd8
      12'hEC1: dout <= 8'b01001110; // 3777 :  78 - 0x4e
      12'hEC2: dout <= 8'b11000010; // 3778 : 194 - 0xc2
      12'hEC3: dout <= 8'b10011010; // 3779 : 154 - 0x9a
      12'hEC4: dout <= 8'b10011011; // 3780 : 155 - 0x9b
      12'hEC5: dout <= 8'b11011001; // 3781 : 217 - 0xd9
      12'hEC6: dout <= 8'b01100011; // 3782 :  99 - 0x63
      12'hEC7: dout <= 8'b00111110; // 3783 :  62 - 0x3e
      12'hEC8: dout <= 8'b00011110; // 3784 :  30 - 0x1e -- Background 0xd9
      12'hEC9: dout <= 8'b01110001; // 3785 : 113 - 0x71
      12'hECA: dout <= 8'b01001001; // 3786 :  73 - 0x49
      12'hECB: dout <= 8'b10111001; // 3787 : 185 - 0xb9
      12'hECC: dout <= 8'b10011101; // 3788 : 157 - 0x9d
      12'hECD: dout <= 8'b01010010; // 3789 :  82 - 0x52
      12'hECE: dout <= 8'b01110010; // 3790 : 114 - 0x72
      12'hECF: dout <= 8'b00011110; // 3791 :  30 - 0x1e
      12'hED0: dout <= 8'b01100000; // 3792 :  96 - 0x60 -- Background 0xda
      12'hED1: dout <= 8'b01011110; // 3793 :  94 - 0x5e
      12'hED2: dout <= 8'b10001001; // 3794 : 137 - 0x89
      12'hED3: dout <= 8'b10111101; // 3795 : 189 - 0xbd
      12'hED4: dout <= 8'b10011101; // 3796 : 157 - 0x9d
      12'hED5: dout <= 8'b11010011; // 3797 : 211 - 0xd3
      12'hED6: dout <= 8'b01000110; // 3798 :  70 - 0x46
      12'hED7: dout <= 8'b01111100; // 3799 : 124 - 0x7c
      12'hED8: dout <= 8'b00011110; // 3800 :  30 - 0x1e -- Background 0xdb
      12'hED9: dout <= 8'b00100011; // 3801 :  35 - 0x23
      12'hEDA: dout <= 8'b01001001; // 3802 :  73 - 0x49
      12'hEDB: dout <= 8'b10111101; // 3803 : 189 - 0xbd
      12'hEDC: dout <= 8'b10011001; // 3804 : 153 - 0x99
      12'hEDD: dout <= 8'b01000011; // 3805 :  67 - 0x43
      12'hEDE: dout <= 8'b01101110; // 3806 : 110 - 0x6e
      12'hEDF: dout <= 8'b00011000; // 3807 :  24 - 0x18
      12'hEE0: dout <= 8'b00000000; // 3808 :   0 - 0x0 -- Background 0xdc
      12'hEE1: dout <= 8'b00000000; // 3809 :   0 - 0x0
      12'hEE2: dout <= 8'b00000001; // 3810 :   1 - 0x1
      12'hEE3: dout <= 8'b00000010; // 3811 :   2 - 0x2
      12'hEE4: dout <= 8'b00000100; // 3812 :   4 - 0x4
      12'hEE5: dout <= 8'b00000010; // 3813 :   2 - 0x2
      12'hEE6: dout <= 8'b00011110; // 3814 :  30 - 0x1e
      12'hEE7: dout <= 8'b00010000; // 3815 :  16 - 0x10
      12'hEE8: dout <= 8'b00001000; // 3816 :   8 - 0x8 -- Background 0xdd
      12'hEE9: dout <= 8'b00001101; // 3817 :  13 - 0xd
      12'hEEA: dout <= 8'b00111010; // 3818 :  58 - 0x3a
      12'hEEB: dout <= 8'b00100101; // 3819 :  37 - 0x25
      12'hEEC: dout <= 8'b00011011; // 3820 :  27 - 0x1b
      12'hEED: dout <= 8'b00001111; // 3821 :  15 - 0xf
      12'hEEE: dout <= 8'b00000111; // 3822 :   7 - 0x7
      12'hEEF: dout <= 8'b00000011; // 3823 :   3 - 0x3
      12'hEF0: dout <= 8'b00000000; // 3824 :   0 - 0x0 -- Background 0xde
      12'hEF1: dout <= 8'b00000000; // 3825 :   0 - 0x0
      12'hEF2: dout <= 8'b00000000; // 3826 :   0 - 0x0
      12'hEF3: dout <= 8'b11000000; // 3827 : 192 - 0xc0
      12'hEF4: dout <= 8'b01000000; // 3828 :  64 - 0x40
      12'hEF5: dout <= 8'b01011000; // 3829 :  88 - 0x58
      12'hEF6: dout <= 8'b01101000; // 3830 : 104 - 0x68
      12'hEF7: dout <= 8'b00001000; // 3831 :   8 - 0x8
      12'hEF8: dout <= 8'b00010000; // 3832 :  16 - 0x10 -- Background 0xdf
      12'hEF9: dout <= 8'b01011100; // 3833 :  92 - 0x5c
      12'hEFA: dout <= 8'b10101000; // 3834 : 168 - 0xa8
      12'hEFB: dout <= 8'b11011000; // 3835 : 216 - 0xd8
      12'hEFC: dout <= 8'b10111000; // 3836 : 184 - 0xb8
      12'hEFD: dout <= 8'b11110000; // 3837 : 240 - 0xf0
      12'hEFE: dout <= 8'b11100000; // 3838 : 224 - 0xe0
      12'hEFF: dout <= 8'b11000000; // 3839 : 192 - 0xc0
      12'hF00: dout <= 8'b00000000; // 3840 :   0 - 0x0 -- Background 0xe0
      12'hF01: dout <= 8'b00000000; // 3841 :   0 - 0x0
      12'hF02: dout <= 8'b00000000; // 3842 :   0 - 0x0
      12'hF03: dout <= 8'b00010011; // 3843 :  19 - 0x13
      12'hF04: dout <= 8'b00010011; // 3844 :  19 - 0x13
      12'hF05: dout <= 8'b00110111; // 3845 :  55 - 0x37
      12'hF06: dout <= 8'b00110111; // 3846 :  55 - 0x37
      12'hF07: dout <= 8'b00000111; // 3847 :   7 - 0x7
      12'hF08: dout <= 8'b00000111; // 3848 :   7 - 0x7 -- Background 0xe1
      12'hF09: dout <= 8'b00000100; // 3849 :   4 - 0x4
      12'hF0A: dout <= 8'b00000000; // 3850 :   0 - 0x0
      12'hF0B: dout <= 8'b00000000; // 3851 :   0 - 0x0
      12'hF0C: dout <= 8'b00000000; // 3852 :   0 - 0x0
      12'hF0D: dout <= 8'b00100000; // 3853 :  32 - 0x20
      12'hF0E: dout <= 8'b01110000; // 3854 : 112 - 0x70
      12'hF0F: dout <= 8'b11111000; // 3855 : 248 - 0xf8
      12'hF10: dout <= 8'b00000000; // 3856 :   0 - 0x0 -- Background 0xe2
      12'hF11: dout <= 8'b00000000; // 3857 :   0 - 0x0
      12'hF12: dout <= 8'b00000000; // 3858 :   0 - 0x0
      12'hF13: dout <= 8'b11111000; // 3859 : 248 - 0xf8
      12'hF14: dout <= 8'b11111100; // 3860 : 252 - 0xfc
      12'hF15: dout <= 8'b11111100; // 3861 : 252 - 0xfc
      12'hF16: dout <= 8'b11111100; // 3862 : 252 - 0xfc
      12'hF17: dout <= 8'b11111101; // 3863 : 253 - 0xfd
      12'hF18: dout <= 8'b11111100; // 3864 : 252 - 0xfc -- Background 0xe3
      12'hF19: dout <= 8'b00011100; // 3865 :  28 - 0x1c
      12'hF1A: dout <= 8'b11000000; // 3866 : 192 - 0xc0
      12'hF1B: dout <= 8'b11100000; // 3867 : 224 - 0xe0
      12'hF1C: dout <= 8'b00000000; // 3868 :   0 - 0x0
      12'hF1D: dout <= 8'b00000000; // 3869 :   0 - 0x0
      12'hF1E: dout <= 8'b00000110; // 3870 :   6 - 0x6
      12'hF1F: dout <= 8'b00001111; // 3871 :  15 - 0xf
      12'hF20: dout <= 8'b00000000; // 3872 :   0 - 0x0 -- Background 0xe4
      12'hF21: dout <= 8'b00000000; // 3873 :   0 - 0x0
      12'hF22: dout <= 8'b00000000; // 3874 :   0 - 0x0
      12'hF23: dout <= 8'b00010011; // 3875 :  19 - 0x13
      12'hF24: dout <= 8'b00010011; // 3876 :  19 - 0x13
      12'hF25: dout <= 8'b00110111; // 3877 :  55 - 0x37
      12'hF26: dout <= 8'b00110111; // 3878 :  55 - 0x37
      12'hF27: dout <= 8'b00000111; // 3879 :   7 - 0x7
      12'hF28: dout <= 8'b00000111; // 3880 :   7 - 0x7 -- Background 0xe5
      12'hF29: dout <= 8'b00000100; // 3881 :   4 - 0x4
      12'hF2A: dout <= 8'b00000001; // 3882 :   1 - 0x1
      12'hF2B: dout <= 8'b00000000; // 3883 :   0 - 0x0
      12'hF2C: dout <= 8'b00000000; // 3884 :   0 - 0x0
      12'hF2D: dout <= 8'b00100000; // 3885 :  32 - 0x20
      12'hF2E: dout <= 8'b01110000; // 3886 : 112 - 0x70
      12'hF2F: dout <= 8'b11111000; // 3887 : 248 - 0xf8
      12'hF30: dout <= 8'b00000000; // 3888 :   0 - 0x0 -- Background 0xe6
      12'hF31: dout <= 8'b00000000; // 3889 :   0 - 0x0
      12'hF32: dout <= 8'b00000000; // 3890 :   0 - 0x0
      12'hF33: dout <= 8'b11111100; // 3891 : 252 - 0xfc
      12'hF34: dout <= 8'b11111100; // 3892 : 252 - 0xfc
      12'hF35: dout <= 8'b11111100; // 3893 : 252 - 0xfc
      12'hF36: dout <= 8'b11111100; // 3894 : 252 - 0xfc
      12'hF37: dout <= 8'b11111101; // 3895 : 253 - 0xfd
      12'hF38: dout <= 8'b11111100; // 3896 : 252 - 0xfc -- Background 0xe7
      12'hF39: dout <= 8'b00001100; // 3897 :  12 - 0xc
      12'hF3A: dout <= 8'b11000000; // 3898 : 192 - 0xc0
      12'hF3B: dout <= 8'b11110000; // 3899 : 240 - 0xf0
      12'hF3C: dout <= 8'b11110000; // 3900 : 240 - 0xf0
      12'hF3D: dout <= 8'b00000000; // 3901 :   0 - 0x0
      12'hF3E: dout <= 8'b00000110; // 3902 :   6 - 0x6
      12'hF3F: dout <= 8'b00001111; // 3903 :  15 - 0xf
      12'hF40: dout <= 8'b11111111; // 3904 : 255 - 0xff -- Background 0xe8
      12'hF41: dout <= 8'b11111111; // 3905 : 255 - 0xff
      12'hF42: dout <= 8'b01111111; // 3906 : 127 - 0x7f
      12'hF43: dout <= 8'b01111111; // 3907 : 127 - 0x7f
      12'hF44: dout <= 8'b01111111; // 3908 : 127 - 0x7f
      12'hF45: dout <= 8'b00111111; // 3909 :  63 - 0x3f
      12'hF46: dout <= 8'b00111111; // 3910 :  63 - 0x3f
      12'hF47: dout <= 8'b00111111; // 3911 :  63 - 0x3f
      12'hF48: dout <= 8'b00111100; // 3912 :  60 - 0x3c -- Background 0xe9
      12'hF49: dout <= 8'b00111110; // 3913 :  62 - 0x3e
      12'hF4A: dout <= 8'b00011111; // 3914 :  31 - 0x1f
      12'hF4B: dout <= 8'b00001111; // 3915 :  15 - 0xf
      12'hF4C: dout <= 8'b00000111; // 3916 :   7 - 0x7
      12'hF4D: dout <= 8'b00000000; // 3917 :   0 - 0x0
      12'hF4E: dout <= 8'b00000000; // 3918 :   0 - 0x0
      12'hF4F: dout <= 8'b00000000; // 3919 :   0 - 0x0
      12'hF50: dout <= 8'b11111111; // 3920 : 255 - 0xff -- Background 0xea
      12'hF51: dout <= 8'b11111110; // 3921 : 254 - 0xfe
      12'hF52: dout <= 8'b11111110; // 3922 : 254 - 0xfe
      12'hF53: dout <= 8'b11111100; // 3923 : 252 - 0xfc
      12'hF54: dout <= 8'b11111000; // 3924 : 248 - 0xf8
      12'hF55: dout <= 8'b11110000; // 3925 : 240 - 0xf0
      12'hF56: dout <= 8'b10110000; // 3926 : 176 - 0xb0
      12'hF57: dout <= 8'b00111001; // 3927 :  57 - 0x39
      12'hF58: dout <= 8'b00011111; // 3928 :  31 - 0x1f -- Background 0xeb
      12'hF59: dout <= 8'b11001111; // 3929 : 207 - 0xcf
      12'hF5A: dout <= 8'b11000110; // 3930 : 198 - 0xc6
      12'hF5B: dout <= 8'b10000000; // 3931 : 128 - 0x80
      12'hF5C: dout <= 8'b00000000; // 3932 :   0 - 0x0
      12'hF5D: dout <= 8'b00000000; // 3933 :   0 - 0x0
      12'hF5E: dout <= 8'b00000000; // 3934 :   0 - 0x0
      12'hF5F: dout <= 8'b00000000; // 3935 :   0 - 0x0
      12'hF60: dout <= 8'b00000000; // 3936 :   0 - 0x0 -- Background 0xec
      12'hF61: dout <= 8'b00000000; // 3937 :   0 - 0x0
      12'hF62: dout <= 8'b00000000; // 3938 :   0 - 0x0
      12'hF63: dout <= 8'b00000000; // 3939 :   0 - 0x0
      12'hF64: dout <= 8'b00000000; // 3940 :   0 - 0x0
      12'hF65: dout <= 8'b00000000; // 3941 :   0 - 0x0
      12'hF66: dout <= 8'b00001100; // 3942 :  12 - 0xc
      12'hF67: dout <= 8'b00001100; // 3943 :  12 - 0xc
      12'hF68: dout <= 8'b00110000; // 3944 :  48 - 0x30 -- Background 0xed
      12'hF69: dout <= 8'b01000011; // 3945 :  67 - 0x43
      12'hF6A: dout <= 8'b01000000; // 3946 :  64 - 0x40
      12'hF6B: dout <= 8'b01100000; // 3947 :  96 - 0x60
      12'hF6C: dout <= 8'b00000011; // 3948 :   3 - 0x3
      12'hF6D: dout <= 8'b00000000; // 3949 :   0 - 0x0
      12'hF6E: dout <= 8'b01111111; // 3950 : 127 - 0x7f
      12'hF6F: dout <= 8'b00000000; // 3951 :   0 - 0x0
      12'hF70: dout <= 8'b00000000; // 3952 :   0 - 0x0 -- Background 0xee
      12'hF71: dout <= 8'b00000000; // 3953 :   0 - 0x0
      12'hF72: dout <= 8'b00000000; // 3954 :   0 - 0x0
      12'hF73: dout <= 8'b00000000; // 3955 :   0 - 0x0
      12'hF74: dout <= 8'b00000000; // 3956 :   0 - 0x0
      12'hF75: dout <= 8'b00000000; // 3957 :   0 - 0x0
      12'hF76: dout <= 8'b00110000; // 3958 :  48 - 0x30
      12'hF77: dout <= 8'b00110000; // 3959 :  48 - 0x30
      12'hF78: dout <= 8'b00001110; // 3960 :  14 - 0xe -- Background 0xef
      12'hF79: dout <= 8'b11001011; // 3961 : 203 - 0xcb
      12'hF7A: dout <= 8'b00000000; // 3962 :   0 - 0x0
      12'hF7B: dout <= 8'b00000000; // 3963 :   0 - 0x0
      12'hF7C: dout <= 8'b11000000; // 3964 : 192 - 0xc0
      12'hF7D: dout <= 8'b00000000; // 3965 :   0 - 0x0
      12'hF7E: dout <= 8'b11111110; // 3966 : 254 - 0xfe
      12'hF7F: dout <= 8'b00000000; // 3967 :   0 - 0x0
      12'hF80: dout <= 8'b00000000; // 3968 :   0 - 0x0 -- Background 0xf0
      12'hF81: dout <= 8'b00000000; // 3969 :   0 - 0x0
      12'hF82: dout <= 8'b00000000; // 3970 :   0 - 0x0
      12'hF83: dout <= 8'b00000000; // 3971 :   0 - 0x0
      12'hF84: dout <= 8'b00000000; // 3972 :   0 - 0x0
      12'hF85: dout <= 8'b00000000; // 3973 :   0 - 0x0
      12'hF86: dout <= 8'b00001100; // 3974 :  12 - 0xc
      12'hF87: dout <= 8'b00001100; // 3975 :  12 - 0xc
      12'hF88: dout <= 8'b00110000; // 3976 :  48 - 0x30 -- Background 0xf1
      12'hF89: dout <= 8'b00100011; // 3977 :  35 - 0x23
      12'hF8A: dout <= 8'b00100000; // 3978 :  32 - 0x20
      12'hF8B: dout <= 8'b01100000; // 3979 :  96 - 0x60
      12'hF8C: dout <= 8'b00000011; // 3980 :   3 - 0x3
      12'hF8D: dout <= 8'b00000000; // 3981 :   0 - 0x0
      12'hF8E: dout <= 8'b01111111; // 3982 : 127 - 0x7f
      12'hF8F: dout <= 8'b00000000; // 3983 :   0 - 0x0
      12'hF90: dout <= 8'b00000000; // 3984 :   0 - 0x0 -- Background 0xf2
      12'hF91: dout <= 8'b00000000; // 3985 :   0 - 0x0
      12'hF92: dout <= 8'b00000000; // 3986 :   0 - 0x0
      12'hF93: dout <= 8'b00000000; // 3987 :   0 - 0x0
      12'hF94: dout <= 8'b00000000; // 3988 :   0 - 0x0
      12'hF95: dout <= 8'b00000000; // 3989 :   0 - 0x0
      12'hF96: dout <= 8'b00110000; // 3990 :  48 - 0x30
      12'hF97: dout <= 8'b00110000; // 3991 :  48 - 0x30
      12'hF98: dout <= 8'b00001001; // 3992 :   9 - 0x9 -- Background 0xf3
      12'hF99: dout <= 8'b11001111; // 3993 : 207 - 0xcf
      12'hF9A: dout <= 8'b00000000; // 3994 :   0 - 0x0
      12'hF9B: dout <= 8'b00000000; // 3995 :   0 - 0x0
      12'hF9C: dout <= 8'b11000000; // 3996 : 192 - 0xc0
      12'hF9D: dout <= 8'b00000000; // 3997 :   0 - 0x0
      12'hF9E: dout <= 8'b11111110; // 3998 : 254 - 0xfe
      12'hF9F: dout <= 8'b00000000; // 3999 :   0 - 0x0
      12'hFA0: dout <= 8'b00111111; // 4000 :  63 - 0x3f -- Background 0xf4
      12'hFA1: dout <= 8'b00110101; // 4001 :  53 - 0x35
      12'hFA2: dout <= 8'b00011010; // 4002 :  26 - 0x1a
      12'hFA3: dout <= 8'b00001101; // 4003 :  13 - 0xd
      12'hFA4: dout <= 8'b00001010; // 4004 :  10 - 0xa
      12'hFA5: dout <= 8'b00001101; // 4005 :  13 - 0xd
      12'hFA6: dout <= 8'b00001000; // 4006 :   8 - 0x8
      12'hFA7: dout <= 8'b00111000; // 4007 :  56 - 0x38
      12'hFA8: dout <= 8'b01110011; // 4008 : 115 - 0x73 -- Background 0xf5
      12'hFA9: dout <= 8'b11000100; // 4009 : 196 - 0xc4
      12'hFAA: dout <= 8'b11000100; // 4010 : 196 - 0xc4
      12'hFAB: dout <= 8'b11000000; // 4011 : 192 - 0xc0
      12'hFAC: dout <= 8'b11000001; // 4012 : 193 - 0xc1
      12'hFAD: dout <= 8'b11000000; // 4013 : 192 - 0xc0
      12'hFAE: dout <= 8'b01100001; // 4014 :  97 - 0x61
      12'hFAF: dout <= 8'b00111111; // 4015 :  63 - 0x3f
      12'hFB0: dout <= 8'b11111100; // 4016 : 252 - 0xfc -- Background 0xf6
      12'hFB1: dout <= 8'b01010100; // 4017 :  84 - 0x54
      12'hFB2: dout <= 8'b10101000; // 4018 : 168 - 0xa8
      12'hFB3: dout <= 8'b01010000; // 4019 :  80 - 0x50
      12'hFB4: dout <= 8'b10110000; // 4020 : 176 - 0xb0
      12'hFB5: dout <= 8'b01010000; // 4021 :  80 - 0x50
      12'hFB6: dout <= 8'b10010000; // 4022 : 144 - 0x90
      12'hFB7: dout <= 8'b00011100; // 4023 :  28 - 0x1c
      12'hFB8: dout <= 8'b10000110; // 4024 : 134 - 0x86 -- Background 0xf7
      12'hFB9: dout <= 8'b01000010; // 4025 :  66 - 0x42
      12'hFBA: dout <= 8'b01000111; // 4026 :  71 - 0x47
      12'hFBB: dout <= 8'b01000001; // 4027 :  65 - 0x41
      12'hFBC: dout <= 8'b10000011; // 4028 : 131 - 0x83
      12'hFBD: dout <= 8'b00000001; // 4029 :   1 - 0x1
      12'hFBE: dout <= 8'b10000110; // 4030 : 134 - 0x86
      12'hFBF: dout <= 8'b11111100; // 4031 : 252 - 0xfc
      12'hFC0: dout <= 8'b11100100; // 4032 : 228 - 0xe4 -- Background 0xf8
      12'hFC1: dout <= 8'b11100100; // 4033 : 228 - 0xe4
      12'hFC2: dout <= 8'b11101111; // 4034 : 239 - 0xef
      12'hFC3: dout <= 8'b11101111; // 4035 : 239 - 0xef
      12'hFC4: dout <= 8'b11111111; // 4036 : 255 - 0xff
      12'hFC5: dout <= 8'b11111111; // 4037 : 255 - 0xff
      12'hFC6: dout <= 8'b01111111; // 4038 : 127 - 0x7f
      12'hFC7: dout <= 8'b01111111; // 4039 : 127 - 0x7f
      12'hFC8: dout <= 8'b00111111; // 4040 :  63 - 0x3f -- Background 0xf9
      12'hFC9: dout <= 8'b01111111; // 4041 : 127 - 0x7f
      12'hFCA: dout <= 8'b01111111; // 4042 : 127 - 0x7f
      12'hFCB: dout <= 8'b11111111; // 4043 : 255 - 0xff
      12'hFCC: dout <= 8'b11111111; // 4044 : 255 - 0xff
      12'hFCD: dout <= 8'b11111111; // 4045 : 255 - 0xff
      12'hFCE: dout <= 8'b11111111; // 4046 : 255 - 0xff
      12'hFCF: dout <= 8'b11111111; // 4047 : 255 - 0xff
      12'hFD0: dout <= 8'b00010011; // 4048 :  19 - 0x13 -- Background 0xfa
      12'hFD1: dout <= 8'b00010011; // 4049 :  19 - 0x13
      12'hFD2: dout <= 8'b11111011; // 4050 : 251 - 0xfb
      12'hFD3: dout <= 8'b11111011; // 4051 : 251 - 0xfb
      12'hFD4: dout <= 8'b11111111; // 4052 : 255 - 0xff
      12'hFD5: dout <= 8'b11111111; // 4053 : 255 - 0xff
      12'hFD6: dout <= 8'b11111110; // 4054 : 254 - 0xfe
      12'hFD7: dout <= 8'b11111110; // 4055 : 254 - 0xfe
      12'hFD8: dout <= 8'b11111110; // 4056 : 254 - 0xfe -- Background 0xfb
      12'hFD9: dout <= 8'b11111111; // 4057 : 255 - 0xff
      12'hFDA: dout <= 8'b11111111; // 4058 : 255 - 0xff
      12'hFDB: dout <= 8'b11111111; // 4059 : 255 - 0xff
      12'hFDC: dout <= 8'b11111111; // 4060 : 255 - 0xff
      12'hFDD: dout <= 8'b11111111; // 4061 : 255 - 0xff
      12'hFDE: dout <= 8'b11111111; // 4062 : 255 - 0xff
      12'hFDF: dout <= 8'b11111111; // 4063 : 255 - 0xff
      12'hFE0: dout <= 8'b00000000; // 4064 :   0 - 0x0 -- Background 0xfc
      12'hFE1: dout <= 8'b00000000; // 4065 :   0 - 0x0
      12'hFE2: dout <= 8'b01111100; // 4066 : 124 - 0x7c
      12'hFE3: dout <= 8'b11111110; // 4067 : 254 - 0xfe
      12'hFE4: dout <= 8'b11111110; // 4068 : 254 - 0xfe
      12'hFE5: dout <= 8'b01111100; // 4069 : 124 - 0x7c
      12'hFE6: dout <= 8'b01000100; // 4070 :  68 - 0x44
      12'hFE7: dout <= 8'b10000010; // 4071 : 130 - 0x82
      12'hFE8: dout <= 8'b10000010; // 4072 : 130 - 0x82 -- Background 0xfd
      12'hFE9: dout <= 8'b10000010; // 4073 : 130 - 0x82
      12'hFEA: dout <= 8'b10000010; // 4074 : 130 - 0x82
      12'hFEB: dout <= 8'b11000110; // 4075 : 198 - 0xc6
      12'hFEC: dout <= 8'b11111110; // 4076 : 254 - 0xfe
      12'hFED: dout <= 8'b11111110; // 4077 : 254 - 0xfe
      12'hFEE: dout <= 8'b10111010; // 4078 : 186 - 0xba
      12'hFEF: dout <= 8'b01111100; // 4079 : 124 - 0x7c
      12'hFF0: dout <= 8'b00000000; // 4080 :   0 - 0x0 -- Background 0xfe
      12'hFF1: dout <= 8'b00011001; // 4081 :  25 - 0x19
      12'hFF2: dout <= 8'b00111110; // 4082 :  62 - 0x3e
      12'hFF3: dout <= 8'b00111100; // 4083 :  60 - 0x3c
      12'hFF4: dout <= 8'b00111100; // 4084 :  60 - 0x3c
      12'hFF5: dout <= 8'b00111100; // 4085 :  60 - 0x3c
      12'hFF6: dout <= 8'b00111110; // 4086 :  62 - 0x3e
      12'hFF7: dout <= 8'b00011001; // 4087 :  25 - 0x19
      12'hFF8: dout <= 8'b00000000; // 4088 :   0 - 0x0 -- Background 0xff
      12'hFF9: dout <= 8'b11111110; // 4089 : 254 - 0xfe
      12'hFFA: dout <= 8'b00011101; // 4090 :  29 - 0x1d
      12'hFFB: dout <= 8'b00001111; // 4091 :  15 - 0xf
      12'hFFC: dout <= 8'b00001111; // 4092 :  15 - 0xf
      12'hFFD: dout <= 8'b00001111; // 4093 :  15 - 0xf
      12'hFFE: dout <= 8'b00011101; // 4094 :  29 - 0x1d
      12'hFFF: dout <= 8'b11111110; // 4095 : 254 - 0xfe
    endcase
  end

endmodule
