//-   Background Pattern table COLOR PLANE 1
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
//- Autcmatically generated verilog ROM from a NES memory file----


//-  Original memory dump file name: nova_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_PTABLE_NOVA_BG_PLN1
  (
     //input     clk,   // clock
     input      [11-1:0] addr,  //2048 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Background pattern Table COLOR PLANE 1
      11'h0: dout  = 8'b00000000; //    0 :   0 - 0x0 -- Background 0x0
      11'h1: dout  = 8'b01111111; //    1 : 127 - 0x7f
      11'h2: dout  = 8'b01111111; //    2 : 127 - 0x7f
      11'h3: dout  = 8'b01111111; //    3 : 127 - 0x7f
      11'h4: dout  = 8'b01111111; //    4 : 127 - 0x7f
      11'h5: dout  = 8'b01111111; //    5 : 127 - 0x7f
      11'h6: dout  = 8'b01101010; //    6 : 106 - 0x6a
      11'h7: dout  = 8'b00000000; //    7 :   0 - 0x0
      11'h8: dout  = 8'b00000000; //    8 :   0 - 0x0 -- Background 0x1
      11'h9: dout  = 8'b01111011; //    9 : 123 - 0x7b
      11'hA: dout  = 8'b01110011; //   10 : 115 - 0x73
      11'hB: dout  = 8'b01111011; //   11 : 123 - 0x7b
      11'hC: dout  = 8'b01110011; //   12 : 115 - 0x73
      11'hD: dout  = 8'b01111011; //   13 : 123 - 0x7b
      11'hE: dout  = 8'b01010011; //   14 :  83 - 0x53
      11'hF: dout  = 8'b00000000; //   15 :   0 - 0x0
      11'h10: dout  = 8'b00000000; //   16 :   0 - 0x0 -- Background 0x2
      11'h11: dout  = 8'b11011110; //   17 : 222 - 0xde
      11'h12: dout  = 8'b10011110; //   18 : 158 - 0x9e
      11'h13: dout  = 8'b11011100; //   19 : 220 - 0xdc
      11'h14: dout  = 8'b10011110; //   20 : 158 - 0x9e
      11'h15: dout  = 8'b11011100; //   21 : 220 - 0xdc
      11'h16: dout  = 8'b10011010; //   22 : 154 - 0x9a
      11'h17: dout  = 8'b00000000; //   23 :   0 - 0x0
      11'h18: dout  = 8'b00000000; //   24 :   0 - 0x0 -- Background 0x3
      11'h19: dout  = 8'b11111110; //   25 : 254 - 0xfe
      11'h1A: dout  = 8'b11111100; //   26 : 252 - 0xfc
      11'h1B: dout  = 8'b11111110; //   27 : 254 - 0xfe
      11'h1C: dout  = 8'b11111100; //   28 : 252 - 0xfc
      11'h1D: dout  = 8'b11111110; //   29 : 254 - 0xfe
      11'h1E: dout  = 8'b01010100; //   30 :  84 - 0x54
      11'h1F: dout  = 8'b00000000; //   31 :   0 - 0x0
      11'h20: dout  = 8'b00000000; //   32 :   0 - 0x0 -- Background 0x4
      11'h21: dout  = 8'b01111111; //   33 : 127 - 0x7f
      11'h22: dout  = 8'b01011111; //   34 :  95 - 0x5f
      11'h23: dout  = 8'b01111001; //   35 : 121 - 0x79
      11'h24: dout  = 8'b01111001; //   36 : 121 - 0x79
      11'h25: dout  = 8'b01001001; //   37 :  73 - 0x49
      11'h26: dout  = 8'b01001111; //   38 :  79 - 0x4f
      11'h27: dout  = 8'b01001110; //   39 :  78 - 0x4e
      11'h28: dout  = 8'b01111000; //   40 : 120 - 0x78 -- Background 0x5
      11'h29: dout  = 8'b01110000; //   41 : 112 - 0x70
      11'h2A: dout  = 8'b01100000; //   42 :  96 - 0x60
      11'h2B: dout  = 8'b01100000; //   43 :  96 - 0x60
      11'h2C: dout  = 8'b01110001; //   44 : 113 - 0x71
      11'h2D: dout  = 8'b01011111; //   45 :  95 - 0x5f
      11'h2E: dout  = 8'b01111111; //   46 : 127 - 0x7f
      11'h2F: dout  = 8'b00000000; //   47 :   0 - 0x0
      11'h30: dout  = 8'b00000000; //   48 :   0 - 0x0 -- Background 0x6
      11'h31: dout  = 8'b11111110; //   49 : 254 - 0xfe
      11'h32: dout  = 8'b11111010; //   50 : 250 - 0xfa
      11'h33: dout  = 8'b10011110; //   51 : 158 - 0x9e
      11'h34: dout  = 8'b10011110; //   52 : 158 - 0x9e
      11'h35: dout  = 8'b10010010; //   53 : 146 - 0x92
      11'h36: dout  = 8'b11110010; //   54 : 242 - 0xf2
      11'h37: dout  = 8'b01110010; //   55 : 114 - 0x72
      11'h38: dout  = 8'b00011110; //   56 :  30 - 0x1e -- Background 0x7
      11'h39: dout  = 8'b00001110; //   57 :  14 - 0xe
      11'h3A: dout  = 8'b00000110; //   58 :   6 - 0x6
      11'h3B: dout  = 8'b00000110; //   59 :   6 - 0x6
      11'h3C: dout  = 8'b10001110; //   60 : 142 - 0x8e
      11'h3D: dout  = 8'b11111010; //   61 : 250 - 0xfa
      11'h3E: dout  = 8'b11111110; //   62 : 254 - 0xfe
      11'h3F: dout  = 8'b00000000; //   63 :   0 - 0x0
      11'h40: dout  = 8'b00000000; //   64 :   0 - 0x0 -- Background 0x8
      11'h41: dout  = 8'b01111111; //   65 : 127 - 0x7f
      11'h42: dout  = 8'b01011111; //   66 :  95 - 0x5f
      11'h43: dout  = 8'b01111111; //   67 : 127 - 0x7f
      11'h44: dout  = 8'b01111111; //   68 : 127 - 0x7f
      11'h45: dout  = 8'b01111111; //   69 : 127 - 0x7f
      11'h46: dout  = 8'b01111111; //   70 : 127 - 0x7f
      11'h47: dout  = 8'b01111111; //   71 : 127 - 0x7f
      11'h48: dout  = 8'b01111111; //   72 : 127 - 0x7f -- Background 0x9
      11'h49: dout  = 8'b01111111; //   73 : 127 - 0x7f
      11'h4A: dout  = 8'b01111111; //   74 : 127 - 0x7f
      11'h4B: dout  = 8'b01111111; //   75 : 127 - 0x7f
      11'h4C: dout  = 8'b01111111; //   76 : 127 - 0x7f
      11'h4D: dout  = 8'b01011111; //   77 :  95 - 0x5f
      11'h4E: dout  = 8'b01111111; //   78 : 127 - 0x7f
      11'h4F: dout  = 8'b00000000; //   79 :   0 - 0x0
      11'h50: dout  = 8'b00000000; //   80 :   0 - 0x0 -- Background 0xa
      11'h51: dout  = 8'b11111110; //   81 : 254 - 0xfe
      11'h52: dout  = 8'b11111010; //   82 : 250 - 0xfa
      11'h53: dout  = 8'b11111110; //   83 : 254 - 0xfe
      11'h54: dout  = 8'b11111110; //   84 : 254 - 0xfe
      11'h55: dout  = 8'b11111110; //   85 : 254 - 0xfe
      11'h56: dout  = 8'b11111110; //   86 : 254 - 0xfe
      11'h57: dout  = 8'b11111110; //   87 : 254 - 0xfe
      11'h58: dout  = 8'b11111110; //   88 : 254 - 0xfe -- Background 0xb
      11'h59: dout  = 8'b11111110; //   89 : 254 - 0xfe
      11'h5A: dout  = 8'b11111110; //   90 : 254 - 0xfe
      11'h5B: dout  = 8'b11111110; //   91 : 254 - 0xfe
      11'h5C: dout  = 8'b11111110; //   92 : 254 - 0xfe
      11'h5D: dout  = 8'b11111010; //   93 : 250 - 0xfa
      11'h5E: dout  = 8'b11111110; //   94 : 254 - 0xfe
      11'h5F: dout  = 8'b00000000; //   95 :   0 - 0x0
      11'h60: dout  = 8'b00000000; //   96 :   0 - 0x0 -- Background 0xc
      11'h61: dout  = 8'b00111111; //   97 :  63 - 0x3f
      11'h62: dout  = 8'b01011111; //   98 :  95 - 0x5f
      11'h63: dout  = 8'b01101111; //   99 : 111 - 0x6f
      11'h64: dout  = 8'b01110000; //  100 : 112 - 0x70
      11'h65: dout  = 8'b01110111; //  101 : 119 - 0x77
      11'h66: dout  = 8'b01110111; //  102 : 119 - 0x77
      11'h67: dout  = 8'b01110111; //  103 : 119 - 0x77
      11'h68: dout  = 8'b01110111; //  104 : 119 - 0x77 -- Background 0xd
      11'h69: dout  = 8'b01110111; //  105 : 119 - 0x77
      11'h6A: dout  = 8'b01110111; //  106 : 119 - 0x77
      11'h6B: dout  = 8'b01110000; //  107 : 112 - 0x70
      11'h6C: dout  = 8'b01101111; //  108 : 111 - 0x6f
      11'h6D: dout  = 8'b01011111; //  109 :  95 - 0x5f
      11'h6E: dout  = 8'b00010101; //  110 :  21 - 0x15
      11'h6F: dout  = 8'b00000000; //  111 :   0 - 0x0
      11'h70: dout  = 8'b00000000; //  112 :   0 - 0x0 -- Background 0xe
      11'h71: dout  = 8'b11111100; //  113 : 252 - 0xfc
      11'h72: dout  = 8'b11111000; //  114 : 248 - 0xf8
      11'h73: dout  = 8'b11110110; //  115 : 246 - 0xf6
      11'h74: dout  = 8'b00001100; //  116 :  12 - 0xc
      11'h75: dout  = 8'b11101110; //  117 : 238 - 0xee
      11'h76: dout  = 8'b11101100; //  118 : 236 - 0xec
      11'h77: dout  = 8'b11101110; //  119 : 238 - 0xee
      11'h78: dout  = 8'b11101100; //  120 : 236 - 0xec -- Background 0xf
      11'h79: dout  = 8'b11101110; //  121 : 238 - 0xee
      11'h7A: dout  = 8'b11101100; //  122 : 236 - 0xec
      11'h7B: dout  = 8'b00001110; //  123 :  14 - 0xe
      11'h7C: dout  = 8'b11110100; //  124 : 244 - 0xf4
      11'h7D: dout  = 8'b11111010; //  125 : 250 - 0xfa
      11'h7E: dout  = 8'b01010100; //  126 :  84 - 0x54
      11'h7F: dout  = 8'b00000000; //  127 :   0 - 0x0
      11'h80: dout  = 8'b01100000; //  128 :  96 - 0x60 -- Background 0x10
      11'h81: dout  = 8'b01100000; //  129 :  96 - 0x60
      11'h82: dout  = 8'b01100000; //  130 :  96 - 0x60
      11'h83: dout  = 8'b01101111; //  131 : 111 - 0x6f
      11'h84: dout  = 8'b01101010; //  132 : 106 - 0x6a
      11'h85: dout  = 8'b01100000; //  133 :  96 - 0x60
      11'h86: dout  = 8'b01100000; //  134 :  96 - 0x60
      11'h87: dout  = 8'b01100000; //  135 :  96 - 0x60
      11'h88: dout  = 8'b00000110; //  136 :   6 - 0x6 -- Background 0x11
      11'h89: dout  = 8'b00000100; //  137 :   4 - 0x4
      11'h8A: dout  = 8'b00000110; //  138 :   6 - 0x6
      11'h8B: dout  = 8'b11110100; //  139 : 244 - 0xf4
      11'h8C: dout  = 8'b10100110; //  140 : 166 - 0xa6
      11'h8D: dout  = 8'b00000100; //  141 :   4 - 0x4
      11'h8E: dout  = 8'b00000110; //  142 :   6 - 0x6
      11'h8F: dout  = 8'b00000100; //  143 :   4 - 0x4
      11'h90: dout  = 8'b00000000; //  144 :   0 - 0x0 -- Background 0x12
      11'h91: dout  = 8'b00001000; //  145 :   8 - 0x8
      11'h92: dout  = 8'b00001000; //  146 :   8 - 0x8
      11'h93: dout  = 8'b00011100; //  147 :  28 - 0x1c
      11'h94: dout  = 8'b00011100; //  148 :  28 - 0x1c
      11'h95: dout  = 8'b00111100; //  149 :  60 - 0x3c
      11'h96: dout  = 8'b00111100; //  150 :  60 - 0x3c
      11'h97: dout  = 8'b00111100; //  151 :  60 - 0x3c
      11'h98: dout  = 8'b00111100; //  152 :  60 - 0x3c -- Background 0x13
      11'h99: dout  = 8'b01111110; //  153 : 126 - 0x7e
      11'h9A: dout  = 8'b01111110; //  154 : 126 - 0x7e
      11'h9B: dout  = 8'b01111110; //  155 : 126 - 0x7e
      11'h9C: dout  = 8'b01111110; //  156 : 126 - 0x7e
      11'h9D: dout  = 8'b01111110; //  157 : 126 - 0x7e
      11'h9E: dout  = 8'b01111110; //  158 : 126 - 0x7e
      11'h9F: dout  = 8'b00000000; //  159 :   0 - 0x0
      11'hA0: dout  = 8'b00000000; //  160 :   0 - 0x0 -- Background 0x14
      11'hA1: dout  = 8'b00000000; //  161 :   0 - 0x0
      11'hA2: dout  = 8'b00000101; //  162 :   5 - 0x5
      11'hA3: dout  = 8'b00000011; //  163 :   3 - 0x3
      11'hA4: dout  = 8'b00000000; //  164 :   0 - 0x0
      11'hA5: dout  = 8'b00000000; //  165 :   0 - 0x0
      11'hA6: dout  = 8'b00000010; //  166 :   2 - 0x2
      11'hA7: dout  = 8'b00001111; //  167 :  15 - 0xf
      11'hA8: dout  = 8'b00011100; //  168 :  28 - 0x1c -- Background 0x15
      11'hA9: dout  = 8'b00111010; //  169 :  58 - 0x3a
      11'hAA: dout  = 8'b00111100; //  170 :  60 - 0x3c
      11'hAB: dout  = 8'b00111111; //  171 :  63 - 0x3f
      11'hAC: dout  = 8'b00111000; //  172 :  56 - 0x38
      11'hAD: dout  = 8'b00011110; //  173 :  30 - 0x1e
      11'hAE: dout  = 8'b00001111; //  174 :  15 - 0xf
      11'hAF: dout  = 8'b00000000; //  175 :   0 - 0x0
      11'hB0: dout  = 8'b00000000; //  176 :   0 - 0x0 -- Background 0x16
      11'hB1: dout  = 8'b00000000; //  177 :   0 - 0x0
      11'hB2: dout  = 8'b01000000; //  178 :  64 - 0x40
      11'hB3: dout  = 8'b11000000; //  179 : 192 - 0xc0
      11'hB4: dout  = 8'b00000000; //  180 :   0 - 0x0
      11'hB5: dout  = 8'b10000000; //  181 : 128 - 0x80
      11'hB6: dout  = 8'b11000000; //  182 : 192 - 0xc0
      11'hB7: dout  = 8'b01110000; //  183 : 112 - 0x70
      11'hB8: dout  = 8'b00011000; //  184 :  24 - 0x18 -- Background 0x17
      11'hB9: dout  = 8'b11111100; //  185 : 252 - 0xfc
      11'hBA: dout  = 8'b00111100; //  186 :  60 - 0x3c
      11'hBB: dout  = 8'b01011100; //  187 :  92 - 0x5c
      11'hBC: dout  = 8'b00111100; //  188 :  60 - 0x3c
      11'hBD: dout  = 8'b11111000; //  189 : 248 - 0xf8
      11'hBE: dout  = 8'b11110000; //  190 : 240 - 0xf0
      11'hBF: dout  = 8'b00000000; //  191 :   0 - 0x0
      11'hC0: dout  = 8'b00000000; //  192 :   0 - 0x0 -- Background 0x18
      11'hC1: dout  = 8'b00111111; //  193 :  63 - 0x3f
      11'hC2: dout  = 8'b00111111; //  194 :  63 - 0x3f
      11'hC3: dout  = 8'b01111111; //  195 : 127 - 0x7f
      11'hC4: dout  = 8'b01111111; //  196 : 127 - 0x7f
      11'hC5: dout  = 8'b00000000; //  197 :   0 - 0x0
      11'hC6: dout  = 8'b00000000; //  198 :   0 - 0x0
      11'hC7: dout  = 8'b00000000; //  199 :   0 - 0x0
      11'hC8: dout  = 8'b00000000; //  200 :   0 - 0x0 -- Background 0x19
      11'hC9: dout  = 8'b11111100; //  201 : 252 - 0xfc
      11'hCA: dout  = 8'b11111100; //  202 : 252 - 0xfc
      11'hCB: dout  = 8'b11111110; //  203 : 254 - 0xfe
      11'hCC: dout  = 8'b11111110; //  204 : 254 - 0xfe
      11'hCD: dout  = 8'b00000000; //  205 :   0 - 0x0
      11'hCE: dout  = 8'b00000000; //  206 :   0 - 0x0
      11'hCF: dout  = 8'b00000000; //  207 :   0 - 0x0
      11'hD0: dout  = 8'b00000000; //  208 :   0 - 0x0 -- Background 0x1a
      11'hD1: dout  = 8'b00000000; //  209 :   0 - 0x0
      11'hD2: dout  = 8'b00000000; //  210 :   0 - 0x0
      11'hD3: dout  = 8'b00111111; //  211 :  63 - 0x3f
      11'hD4: dout  = 8'b00111111; //  212 :  63 - 0x3f
      11'hD5: dout  = 8'b01111111; //  213 : 127 - 0x7f
      11'hD6: dout  = 8'b01111111; //  214 : 127 - 0x7f
      11'hD7: dout  = 8'b00000000; //  215 :   0 - 0x0
      11'hD8: dout  = 8'b00000000; //  216 :   0 - 0x0 -- Background 0x1b
      11'hD9: dout  = 8'b00000000; //  217 :   0 - 0x0
      11'hDA: dout  = 8'b00000000; //  218 :   0 - 0x0
      11'hDB: dout  = 8'b11111100; //  219 : 252 - 0xfc
      11'hDC: dout  = 8'b11111100; //  220 : 252 - 0xfc
      11'hDD: dout  = 8'b11111110; //  221 : 254 - 0xfe
      11'hDE: dout  = 8'b11111110; //  222 : 254 - 0xfe
      11'hDF: dout  = 8'b00000000; //  223 :   0 - 0x0
      11'hE0: dout  = 8'b00000000; //  224 :   0 - 0x0 -- Background 0x1c
      11'hE1: dout  = 8'b01111111; //  225 : 127 - 0x7f
      11'hE2: dout  = 8'b01111111; //  226 : 127 - 0x7f
      11'hE3: dout  = 8'b01111111; //  227 : 127 - 0x7f
      11'hE4: dout  = 8'b01100100; //  228 : 100 - 0x64
      11'hE5: dout  = 8'b01011011; //  229 :  91 - 0x5b
      11'hE6: dout  = 8'b01011001; //  230 :  89 - 0x59
      11'hE7: dout  = 8'b01111111; //  231 : 127 - 0x7f
      11'hE8: dout  = 8'b01111111; //  232 : 127 - 0x7f -- Background 0x1d
      11'hE9: dout  = 8'b00000000; //  233 :   0 - 0x0
      11'hEA: dout  = 8'b00000001; //  234 :   1 - 0x1
      11'hEB: dout  = 8'b00000001; //  235 :   1 - 0x1
      11'hEC: dout  = 8'b00000001; //  236 :   1 - 0x1
      11'hED: dout  = 8'b00000001; //  237 :   1 - 0x1
      11'hEE: dout  = 8'b00000001; //  238 :   1 - 0x1
      11'hEF: dout  = 8'b00000000; //  239 :   0 - 0x0
      11'hF0: dout  = 8'b00000000; //  240 :   0 - 0x0 -- Background 0x1e
      11'hF1: dout  = 8'b11111110; //  241 : 254 - 0xfe
      11'hF2: dout  = 8'b11111110; //  242 : 254 - 0xfe
      11'hF3: dout  = 8'b11111110; //  243 : 254 - 0xfe
      11'hF4: dout  = 8'b10111110; //  244 : 190 - 0xbe
      11'hF5: dout  = 8'b00001010; //  245 :  10 - 0xa
      11'hF6: dout  = 8'b11100010; //  246 : 226 - 0xe2
      11'hF7: dout  = 8'b11111110; //  247 : 254 - 0xfe
      11'hF8: dout  = 8'b11111110; //  248 : 254 - 0xfe -- Background 0x1f
      11'hF9: dout  = 8'b00000000; //  249 :   0 - 0x0
      11'hFA: dout  = 8'b10000000; //  250 : 128 - 0x80
      11'hFB: dout  = 8'b10000000; //  251 : 128 - 0x80
      11'hFC: dout  = 8'b10000000; //  252 : 128 - 0x80
      11'hFD: dout  = 8'b10000000; //  253 : 128 - 0x80
      11'hFE: dout  = 8'b10000000; //  254 : 128 - 0x80
      11'hFF: dout  = 8'b00000000; //  255 :   0 - 0x0
      11'h100: dout  = 8'b00000000; //  256 :   0 - 0x0 -- Background 0x20
      11'h101: dout  = 8'b00000000; //  257 :   0 - 0x0
      11'h102: dout  = 8'b00000000; //  258 :   0 - 0x0
      11'h103: dout  = 8'b00000000; //  259 :   0 - 0x0
      11'h104: dout  = 8'b00000000; //  260 :   0 - 0x0
      11'h105: dout  = 8'b00000000; //  261 :   0 - 0x0
      11'h106: dout  = 8'b00000000; //  262 :   0 - 0x0
      11'h107: dout  = 8'b00000000; //  263 :   0 - 0x0
      11'h108: dout  = 8'b00000000; //  264 :   0 - 0x0 -- Background 0x21
      11'h109: dout  = 8'b00000000; //  265 :   0 - 0x0
      11'h10A: dout  = 8'b00000000; //  266 :   0 - 0x0
      11'h10B: dout  = 8'b00000000; //  267 :   0 - 0x0
      11'h10C: dout  = 8'b00000000; //  268 :   0 - 0x0
      11'h10D: dout  = 8'b00000000; //  269 :   0 - 0x0
      11'h10E: dout  = 8'b00000000; //  270 :   0 - 0x0
      11'h10F: dout  = 8'b00000000; //  271 :   0 - 0x0
      11'h110: dout  = 8'b00000000; //  272 :   0 - 0x0 -- Background 0x22
      11'h111: dout  = 8'b00000000; //  273 :   0 - 0x0
      11'h112: dout  = 8'b00011000; //  274 :  24 - 0x18
      11'h113: dout  = 8'b00010000; //  275 :  16 - 0x10
      11'h114: dout  = 8'b00011010; //  276 :  26 - 0x1a
      11'h115: dout  = 8'b00010001; //  277 :  17 - 0x11
      11'h116: dout  = 8'b00011010; //  278 :  26 - 0x1a
      11'h117: dout  = 8'b00000000; //  279 :   0 - 0x0
      11'h118: dout  = 8'b00000000; //  280 :   0 - 0x0 -- Background 0x23
      11'h119: dout  = 8'b00000000; //  281 :   0 - 0x0
      11'h11A: dout  = 8'b00000000; //  282 :   0 - 0x0
      11'h11B: dout  = 8'b00101000; //  283 :  40 - 0x28
      11'h11C: dout  = 8'b10001100; //  284 : 140 - 0x8c
      11'h11D: dout  = 8'b00101000; //  285 :  40 - 0x28
      11'h11E: dout  = 8'b10101100; //  286 : 172 - 0xac
      11'h11F: dout  = 8'b00000000; //  287 :   0 - 0x0
      11'h120: dout  = 8'b00000000; //  288 :   0 - 0x0 -- Background 0x24
      11'h121: dout  = 8'b00000000; //  289 :   0 - 0x0
      11'h122: dout  = 8'b00000000; //  290 :   0 - 0x0
      11'h123: dout  = 8'b00000000; //  291 :   0 - 0x0
      11'h124: dout  = 8'b00000000; //  292 :   0 - 0x0
      11'h125: dout  = 8'b00000000; //  293 :   0 - 0x0
      11'h126: dout  = 8'b00000000; //  294 :   0 - 0x0
      11'h127: dout  = 8'b00000000; //  295 :   0 - 0x0
      11'h128: dout  = 8'b00011100; //  296 :  28 - 0x1c -- Background 0x25
      11'h129: dout  = 8'b00111001; //  297 :  57 - 0x39
      11'h12A: dout  = 8'b00111111; //  298 :  63 - 0x3f
      11'h12B: dout  = 8'b00111110; //  299 :  62 - 0x3e
      11'h12C: dout  = 8'b00111111; //  300 :  63 - 0x3f
      11'h12D: dout  = 8'b00011110; //  301 :  30 - 0x1e
      11'h12E: dout  = 8'b00001111; //  302 :  15 - 0xf
      11'h12F: dout  = 8'b00000000; //  303 :   0 - 0x0
      11'h130: dout  = 8'b00000000; //  304 :   0 - 0x0 -- Background 0x26
      11'h131: dout  = 8'b00000000; //  305 :   0 - 0x0
      11'h132: dout  = 8'b01000000; //  306 :  64 - 0x40
      11'h133: dout  = 8'b11000000; //  307 : 192 - 0xc0
      11'h134: dout  = 8'b00000000; //  308 :   0 - 0x0
      11'h135: dout  = 8'b10000000; //  309 : 128 - 0x80
      11'h136: dout  = 8'b11000000; //  310 : 192 - 0xc0
      11'h137: dout  = 8'b11110000; //  311 : 240 - 0xf0
      11'h138: dout  = 8'b00111000; //  312 :  56 - 0x38 -- Background 0x27
      11'h139: dout  = 8'b10011100; //  313 : 156 - 0x9c
      11'h13A: dout  = 8'b10011100; //  314 : 156 - 0x9c
      11'h13B: dout  = 8'b00111100; //  315 :  60 - 0x3c
      11'h13C: dout  = 8'b11111100; //  316 : 252 - 0xfc
      11'h13D: dout  = 8'b01111000; //  317 : 120 - 0x78
      11'h13E: dout  = 8'b11110000; //  318 : 240 - 0xf0
      11'h13F: dout  = 8'b00000000; //  319 :   0 - 0x0
      11'h140: dout  = 8'b00000000; //  320 :   0 - 0x0 -- Background 0x28
      11'h141: dout  = 8'b00111110; //  321 :  62 - 0x3e
      11'h142: dout  = 8'b01011101; //  322 :  93 - 0x5d
      11'h143: dout  = 8'b01101011; //  323 : 107 - 0x6b
      11'h144: dout  = 8'b01110101; //  324 : 117 - 0x75
      11'h145: dout  = 8'b01110001; //  325 : 113 - 0x71
      11'h146: dout  = 8'b01110101; //  326 : 117 - 0x75
      11'h147: dout  = 8'b01110100; //  327 : 116 - 0x74
      11'h148: dout  = 8'b01110000; //  328 : 112 - 0x70 -- Background 0x29
      11'h149: dout  = 8'b01110111; //  329 : 119 - 0x77
      11'h14A: dout  = 8'b01110111; //  330 : 119 - 0x77
      11'h14B: dout  = 8'b01110000; //  331 : 112 - 0x70
      11'h14C: dout  = 8'b01101111; //  332 : 111 - 0x6f
      11'h14D: dout  = 8'b01011111; //  333 :  95 - 0x5f
      11'h14E: dout  = 8'b00010101; //  334 :  21 - 0x15
      11'h14F: dout  = 8'b00000000; //  335 :   0 - 0x0
      11'h150: dout  = 8'b00000000; //  336 :   0 - 0x0 -- Background 0x2a
      11'h151: dout  = 8'b01111100; //  337 : 124 - 0x7c
      11'h152: dout  = 8'b10111000; //  338 : 184 - 0xb8
      11'h153: dout  = 8'b11010110; //  339 : 214 - 0xd6
      11'h154: dout  = 8'b10101100; //  340 : 172 - 0xac
      11'h155: dout  = 8'b10001110; //  341 : 142 - 0x8e
      11'h156: dout  = 8'b10101100; //  342 : 172 - 0xac
      11'h157: dout  = 8'b00101110; //  343 :  46 - 0x2e
      11'h158: dout  = 8'b00001100; //  344 :  12 - 0xc -- Background 0x2b
      11'h159: dout  = 8'b11101110; //  345 : 238 - 0xee
      11'h15A: dout  = 8'b11101100; //  346 : 236 - 0xec
      11'h15B: dout  = 8'b00001110; //  347 :  14 - 0xe
      11'h15C: dout  = 8'b11110100; //  348 : 244 - 0xf4
      11'h15D: dout  = 8'b11111010; //  349 : 250 - 0xfa
      11'h15E: dout  = 8'b01010100; //  350 :  84 - 0x54
      11'h15F: dout  = 8'b00000000; //  351 :   0 - 0x0
      11'h160: dout  = 8'b00000000; //  352 :   0 - 0x0 -- Background 0x2c
      11'h161: dout  = 8'b00000000; //  353 :   0 - 0x0
      11'h162: dout  = 8'b00000000; //  354 :   0 - 0x0
      11'h163: dout  = 8'b00000000; //  355 :   0 - 0x0
      11'h164: dout  = 8'b00000000; //  356 :   0 - 0x0
      11'h165: dout  = 8'b00000000; //  357 :   0 - 0x0
      11'h166: dout  = 8'b00000000; //  358 :   0 - 0x0
      11'h167: dout  = 8'b00000000; //  359 :   0 - 0x0
      11'h168: dout  = 8'b00011110; //  360 :  30 - 0x1e -- Background 0x2d
      11'h169: dout  = 8'b00111110; //  361 :  62 - 0x3e
      11'h16A: dout  = 8'b00111110; //  362 :  62 - 0x3e
      11'h16B: dout  = 8'b00111110; //  363 :  62 - 0x3e
      11'h16C: dout  = 8'b00111111; //  364 :  63 - 0x3f
      11'h16D: dout  = 8'b00011110; //  365 :  30 - 0x1e
      11'h16E: dout  = 8'b00001111; //  366 :  15 - 0xf
      11'h16F: dout  = 8'b00000000; //  367 :   0 - 0x0
      11'h170: dout  = 8'b00000000; //  368 :   0 - 0x0 -- Background 0x2e
      11'h171: dout  = 8'b00000000; //  369 :   0 - 0x0
      11'h172: dout  = 8'b00000000; //  370 :   0 - 0x0
      11'h173: dout  = 8'b00000000; //  371 :   0 - 0x0
      11'h174: dout  = 8'b00000000; //  372 :   0 - 0x0
      11'h175: dout  = 8'b00000000; //  373 :   0 - 0x0
      11'h176: dout  = 8'b00000000; //  374 :   0 - 0x0
      11'h177: dout  = 8'b00000000; //  375 :   0 - 0x0
      11'h178: dout  = 8'b01111000; //  376 : 120 - 0x78 -- Background 0x2f
      11'h179: dout  = 8'b01111100; //  377 : 124 - 0x7c
      11'h17A: dout  = 8'b01111100; //  378 : 124 - 0x7c
      11'h17B: dout  = 8'b01111100; //  379 : 124 - 0x7c
      11'h17C: dout  = 8'b11111100; //  380 : 252 - 0xfc
      11'h17D: dout  = 8'b01111000; //  381 : 120 - 0x78
      11'h17E: dout  = 8'b11110000; //  382 : 240 - 0xf0
      11'h17F: dout  = 8'b00000000; //  383 :   0 - 0x0
      11'h180: dout  = 8'b00000000; //  384 :   0 - 0x0 -- Background 0x30
      11'h181: dout  = 8'b00011000; //  385 :  24 - 0x18
      11'h182: dout  = 8'b00111100; //  386 :  60 - 0x3c
      11'h183: dout  = 8'b01011010; //  387 :  90 - 0x5a
      11'h184: dout  = 8'b00011000; //  388 :  24 - 0x18
      11'h185: dout  = 8'b00011000; //  389 :  24 - 0x18
      11'h186: dout  = 8'b00011000; //  390 :  24 - 0x18
      11'h187: dout  = 8'b00000000; //  391 :   0 - 0x0
      11'h188: dout  = 8'b00000000; //  392 :   0 - 0x0 -- Background 0x31
      11'h189: dout  = 8'b00011000; //  393 :  24 - 0x18
      11'h18A: dout  = 8'b00011000; //  394 :  24 - 0x18
      11'h18B: dout  = 8'b00011000; //  395 :  24 - 0x18
      11'h18C: dout  = 8'b01011010; //  396 :  90 - 0x5a
      11'h18D: dout  = 8'b00111100; //  397 :  60 - 0x3c
      11'h18E: dout  = 8'b00011000; //  398 :  24 - 0x18
      11'h18F: dout  = 8'b00000000; //  399 :   0 - 0x0
      11'h190: dout  = 8'b00000001; //  400 :   1 - 0x1 -- Background 0x32
      11'h191: dout  = 8'b00000001; //  401 :   1 - 0x1
      11'h192: dout  = 8'b00000000; //  402 :   0 - 0x0
      11'h193: dout  = 8'b00000001; //  403 :   1 - 0x1
      11'h194: dout  = 8'b00000001; //  404 :   1 - 0x1
      11'h195: dout  = 8'b00000001; //  405 :   1 - 0x1
      11'h196: dout  = 8'b00000000; //  406 :   0 - 0x0
      11'h197: dout  = 8'b00000001; //  407 :   1 - 0x1
      11'h198: dout  = 8'b10000000; //  408 : 128 - 0x80 -- Background 0x33
      11'h199: dout  = 8'b00000000; //  409 :   0 - 0x0
      11'h19A: dout  = 8'b10000000; //  410 : 128 - 0x80
      11'h19B: dout  = 8'b10000000; //  411 : 128 - 0x80
      11'h19C: dout  = 8'b10000000; //  412 : 128 - 0x80
      11'h19D: dout  = 8'b00000000; //  413 :   0 - 0x0
      11'h19E: dout  = 8'b10000000; //  414 : 128 - 0x80
      11'h19F: dout  = 8'b10000000; //  415 : 128 - 0x80
      11'h1A0: dout  = 8'b00000000; //  416 :   0 - 0x0 -- Background 0x34
      11'h1A1: dout  = 8'b00000000; //  417 :   0 - 0x0
      11'h1A2: dout  = 8'b00011000; //  418 :  24 - 0x18
      11'h1A3: dout  = 8'b00111100; //  419 :  60 - 0x3c
      11'h1A4: dout  = 8'b00111110; //  420 :  62 - 0x3e
      11'h1A5: dout  = 8'b01111111; //  421 : 127 - 0x7f
      11'h1A6: dout  = 8'b01111111; //  422 : 127 - 0x7f
      11'h1A7: dout  = 8'b01111111; //  423 : 127 - 0x7f
      11'h1A8: dout  = 8'b00111111; //  424 :  63 - 0x3f -- Background 0x35
      11'h1A9: dout  = 8'b00111111; //  425 :  63 - 0x3f
      11'h1AA: dout  = 8'b00011111; //  426 :  31 - 0x1f
      11'h1AB: dout  = 8'b00001111; //  427 :  15 - 0xf
      11'h1AC: dout  = 8'b00000111; //  428 :   7 - 0x7
      11'h1AD: dout  = 8'b00000011; //  429 :   3 - 0x3
      11'h1AE: dout  = 8'b00000001; //  430 :   1 - 0x1
      11'h1AF: dout  = 8'b00000000; //  431 :   0 - 0x0
      11'h1B0: dout  = 8'b00000000; //  432 :   0 - 0x0 -- Background 0x36
      11'h1B1: dout  = 8'b00000000; //  433 :   0 - 0x0
      11'h1B2: dout  = 8'b00011000; //  434 :  24 - 0x18
      11'h1B3: dout  = 8'b00111100; //  435 :  60 - 0x3c
      11'h1B4: dout  = 8'b01111100; //  436 : 124 - 0x7c
      11'h1B5: dout  = 8'b11111110; //  437 : 254 - 0xfe
      11'h1B6: dout  = 8'b11111110; //  438 : 254 - 0xfe
      11'h1B7: dout  = 8'b11111110; //  439 : 254 - 0xfe
      11'h1B8: dout  = 8'b11111100; //  440 : 252 - 0xfc -- Background 0x37
      11'h1B9: dout  = 8'b11111100; //  441 : 252 - 0xfc
      11'h1BA: dout  = 8'b11111000; //  442 : 248 - 0xf8
      11'h1BB: dout  = 8'b11110000; //  443 : 240 - 0xf0
      11'h1BC: dout  = 8'b11100000; //  444 : 224 - 0xe0
      11'h1BD: dout  = 8'b11000000; //  445 : 192 - 0xc0
      11'h1BE: dout  = 8'b10000000; //  446 : 128 - 0x80
      11'h1BF: dout  = 8'b00000000; //  447 :   0 - 0x0
      11'h1C0: dout  = 8'b00000000; //  448 :   0 - 0x0 -- Background 0x38
      11'h1C1: dout  = 8'b00000000; //  449 :   0 - 0x0
      11'h1C2: dout  = 8'b00000110; //  450 :   6 - 0x6
      11'h1C3: dout  = 8'b00000111; //  451 :   7 - 0x7
      11'h1C4: dout  = 8'b00000111; //  452 :   7 - 0x7
      11'h1C5: dout  = 8'b00000011; //  453 :   3 - 0x3
      11'h1C6: dout  = 8'b00000001; //  454 :   1 - 0x1
      11'h1C7: dout  = 8'b00000000; //  455 :   0 - 0x0
      11'h1C8: dout  = 8'b00000000; //  456 :   0 - 0x0 -- Background 0x39
      11'h1C9: dout  = 8'b00000000; //  457 :   0 - 0x0
      11'h1CA: dout  = 8'b00000000; //  458 :   0 - 0x0
      11'h1CB: dout  = 8'b00000000; //  459 :   0 - 0x0
      11'h1CC: dout  = 8'b00000000; //  460 :   0 - 0x0
      11'h1CD: dout  = 8'b00000000; //  461 :   0 - 0x0
      11'h1CE: dout  = 8'b00000000; //  462 :   0 - 0x0
      11'h1CF: dout  = 8'b00000000; //  463 :   0 - 0x0
      11'h1D0: dout  = 8'b00000000; //  464 :   0 - 0x0 -- Background 0x3a
      11'h1D1: dout  = 8'b00000000; //  465 :   0 - 0x0
      11'h1D2: dout  = 8'b01100000; //  466 :  96 - 0x60
      11'h1D3: dout  = 8'b11100000; //  467 : 224 - 0xe0
      11'h1D4: dout  = 8'b11100000; //  468 : 224 - 0xe0
      11'h1D5: dout  = 8'b11000000; //  469 : 192 - 0xc0
      11'h1D6: dout  = 8'b10000000; //  470 : 128 - 0x80
      11'h1D7: dout  = 8'b00000000; //  471 :   0 - 0x0
      11'h1D8: dout  = 8'b00000000; //  472 :   0 - 0x0 -- Background 0x3b
      11'h1D9: dout  = 8'b00101010; //  473 :  42 - 0x2a
      11'h1DA: dout  = 8'b01000000; //  474 :  64 - 0x40
      11'h1DB: dout  = 8'b00000010; //  475 :   2 - 0x2
      11'h1DC: dout  = 8'b01000000; //  476 :  64 - 0x40
      11'h1DD: dout  = 8'b00000010; //  477 :   2 - 0x2
      11'h1DE: dout  = 8'b01010100; //  478 :  84 - 0x54
      11'h1DF: dout  = 8'b00000000; //  479 :   0 - 0x0
      11'h1E0: dout  = 8'b00000000; //  480 :   0 - 0x0 -- Background 0x3c
      11'h1E1: dout  = 8'b00000000; //  481 :   0 - 0x0
      11'h1E2: dout  = 8'b00000000; //  482 :   0 - 0x0
      11'h1E3: dout  = 8'b00000000; //  483 :   0 - 0x0
      11'h1E4: dout  = 8'b00000000; //  484 :   0 - 0x0
      11'h1E5: dout  = 8'b00000000; //  485 :   0 - 0x0
      11'h1E6: dout  = 8'b00000000; //  486 :   0 - 0x0
      11'h1E7: dout  = 8'b00000000; //  487 :   0 - 0x0
      11'h1E8: dout  = 8'b11111111; //  488 : 255 - 0xff -- Background 0x3d
      11'h1E9: dout  = 8'b11111111; //  489 : 255 - 0xff
      11'h1EA: dout  = 8'b11111111; //  490 : 255 - 0xff
      11'h1EB: dout  = 8'b11111111; //  491 : 255 - 0xff
      11'h1EC: dout  = 8'b11111111; //  492 : 255 - 0xff
      11'h1ED: dout  = 8'b11111111; //  493 : 255 - 0xff
      11'h1EE: dout  = 8'b11111111; //  494 : 255 - 0xff
      11'h1EF: dout  = 8'b11111111; //  495 : 255 - 0xff
      11'h1F0: dout  = 8'b11111111; //  496 : 255 - 0xff -- Background 0x3e
      11'h1F1: dout  = 8'b11111111; //  497 : 255 - 0xff
      11'h1F2: dout  = 8'b11111111; //  498 : 255 - 0xff
      11'h1F3: dout  = 8'b11111111; //  499 : 255 - 0xff
      11'h1F4: dout  = 8'b11111111; //  500 : 255 - 0xff
      11'h1F5: dout  = 8'b11111111; //  501 : 255 - 0xff
      11'h1F6: dout  = 8'b11111111; //  502 : 255 - 0xff
      11'h1F7: dout  = 8'b11111111; //  503 : 255 - 0xff
      11'h1F8: dout  = 8'b00000000; //  504 :   0 - 0x0 -- Background 0x3f
      11'h1F9: dout  = 8'b00000000; //  505 :   0 - 0x0
      11'h1FA: dout  = 8'b00000000; //  506 :   0 - 0x0
      11'h1FB: dout  = 8'b00000000; //  507 :   0 - 0x0
      11'h1FC: dout  = 8'b00000000; //  508 :   0 - 0x0
      11'h1FD: dout  = 8'b00000000; //  509 :   0 - 0x0
      11'h1FE: dout  = 8'b00000000; //  510 :   0 - 0x0
      11'h1FF: dout  = 8'b00000000; //  511 :   0 - 0x0
      11'h200: dout  = 8'b00000000; //  512 :   0 - 0x0 -- Background 0x40
      11'h201: dout  = 8'b00000000; //  513 :   0 - 0x0
      11'h202: dout  = 8'b00000000; //  514 :   0 - 0x0
      11'h203: dout  = 8'b00000000; //  515 :   0 - 0x0
      11'h204: dout  = 8'b00000000; //  516 :   0 - 0x0
      11'h205: dout  = 8'b00000000; //  517 :   0 - 0x0
      11'h206: dout  = 8'b00000000; //  518 :   0 - 0x0
      11'h207: dout  = 8'b00000000; //  519 :   0 - 0x0
      11'h208: dout  = 8'b00000000; //  520 :   0 - 0x0 -- Background 0x41
      11'h209: dout  = 8'b00000000; //  521 :   0 - 0x0
      11'h20A: dout  = 8'b00000000; //  522 :   0 - 0x0
      11'h20B: dout  = 8'b00000000; //  523 :   0 - 0x0
      11'h20C: dout  = 8'b00000000; //  524 :   0 - 0x0
      11'h20D: dout  = 8'b00000000; //  525 :   0 - 0x0
      11'h20E: dout  = 8'b00000000; //  526 :   0 - 0x0
      11'h20F: dout  = 8'b00000000; //  527 :   0 - 0x0
      11'h210: dout  = 8'b00000000; //  528 :   0 - 0x0 -- Background 0x42
      11'h211: dout  = 8'b00000000; //  529 :   0 - 0x0
      11'h212: dout  = 8'b00000000; //  530 :   0 - 0x0
      11'h213: dout  = 8'b00000000; //  531 :   0 - 0x0
      11'h214: dout  = 8'b00000000; //  532 :   0 - 0x0
      11'h215: dout  = 8'b00000000; //  533 :   0 - 0x0
      11'h216: dout  = 8'b00000000; //  534 :   0 - 0x0
      11'h217: dout  = 8'b00000000; //  535 :   0 - 0x0
      11'h218: dout  = 8'b00000000; //  536 :   0 - 0x0 -- Background 0x43
      11'h219: dout  = 8'b00000000; //  537 :   0 - 0x0
      11'h21A: dout  = 8'b00000000; //  538 :   0 - 0x0
      11'h21B: dout  = 8'b00000000; //  539 :   0 - 0x0
      11'h21C: dout  = 8'b00000000; //  540 :   0 - 0x0
      11'h21D: dout  = 8'b00000000; //  541 :   0 - 0x0
      11'h21E: dout  = 8'b00000000; //  542 :   0 - 0x0
      11'h21F: dout  = 8'b00000000; //  543 :   0 - 0x0
      11'h220: dout  = 8'b00000000; //  544 :   0 - 0x0 -- Background 0x44
      11'h221: dout  = 8'b00000000; //  545 :   0 - 0x0
      11'h222: dout  = 8'b00000000; //  546 :   0 - 0x0
      11'h223: dout  = 8'b00000000; //  547 :   0 - 0x0
      11'h224: dout  = 8'b00000000; //  548 :   0 - 0x0
      11'h225: dout  = 8'b00000000; //  549 :   0 - 0x0
      11'h226: dout  = 8'b00000000; //  550 :   0 - 0x0
      11'h227: dout  = 8'b00000000; //  551 :   0 - 0x0
      11'h228: dout  = 8'b00000000; //  552 :   0 - 0x0 -- Background 0x45
      11'h229: dout  = 8'b00000000; //  553 :   0 - 0x0
      11'h22A: dout  = 8'b00000000; //  554 :   0 - 0x0
      11'h22B: dout  = 8'b00000000; //  555 :   0 - 0x0
      11'h22C: dout  = 8'b00000000; //  556 :   0 - 0x0
      11'h22D: dout  = 8'b00000000; //  557 :   0 - 0x0
      11'h22E: dout  = 8'b00000000; //  558 :   0 - 0x0
      11'h22F: dout  = 8'b00000000; //  559 :   0 - 0x0
      11'h230: dout  = 8'b00000000; //  560 :   0 - 0x0 -- Background 0x46
      11'h231: dout  = 8'b00000000; //  561 :   0 - 0x0
      11'h232: dout  = 8'b00000000; //  562 :   0 - 0x0
      11'h233: dout  = 8'b00000000; //  563 :   0 - 0x0
      11'h234: dout  = 8'b00000000; //  564 :   0 - 0x0
      11'h235: dout  = 8'b00000000; //  565 :   0 - 0x0
      11'h236: dout  = 8'b00000000; //  566 :   0 - 0x0
      11'h237: dout  = 8'b00000000; //  567 :   0 - 0x0
      11'h238: dout  = 8'b00000000; //  568 :   0 - 0x0 -- Background 0x47
      11'h239: dout  = 8'b00000000; //  569 :   0 - 0x0
      11'h23A: dout  = 8'b00000000; //  570 :   0 - 0x0
      11'h23B: dout  = 8'b00000000; //  571 :   0 - 0x0
      11'h23C: dout  = 8'b00000000; //  572 :   0 - 0x0
      11'h23D: dout  = 8'b00000000; //  573 :   0 - 0x0
      11'h23E: dout  = 8'b00000000; //  574 :   0 - 0x0
      11'h23F: dout  = 8'b00000000; //  575 :   0 - 0x0
      11'h240: dout  = 8'b00000000; //  576 :   0 - 0x0 -- Background 0x48
      11'h241: dout  = 8'b00000000; //  577 :   0 - 0x0
      11'h242: dout  = 8'b00000000; //  578 :   0 - 0x0
      11'h243: dout  = 8'b00000000; //  579 :   0 - 0x0
      11'h244: dout  = 8'b00000000; //  580 :   0 - 0x0
      11'h245: dout  = 8'b00000000; //  581 :   0 - 0x0
      11'h246: dout  = 8'b00000000; //  582 :   0 - 0x0
      11'h247: dout  = 8'b00000000; //  583 :   0 - 0x0
      11'h248: dout  = 8'b00000000; //  584 :   0 - 0x0 -- Background 0x49
      11'h249: dout  = 8'b00000000; //  585 :   0 - 0x0
      11'h24A: dout  = 8'b00000000; //  586 :   0 - 0x0
      11'h24B: dout  = 8'b00000000; //  587 :   0 - 0x0
      11'h24C: dout  = 8'b00000000; //  588 :   0 - 0x0
      11'h24D: dout  = 8'b00000000; //  589 :   0 - 0x0
      11'h24E: dout  = 8'b00000000; //  590 :   0 - 0x0
      11'h24F: dout  = 8'b00000000; //  591 :   0 - 0x0
      11'h250: dout  = 8'b00000000; //  592 :   0 - 0x0 -- Background 0x4a
      11'h251: dout  = 8'b00000000; //  593 :   0 - 0x0
      11'h252: dout  = 8'b00000000; //  594 :   0 - 0x0
      11'h253: dout  = 8'b00000000; //  595 :   0 - 0x0
      11'h254: dout  = 8'b00000000; //  596 :   0 - 0x0
      11'h255: dout  = 8'b00000000; //  597 :   0 - 0x0
      11'h256: dout  = 8'b00000000; //  598 :   0 - 0x0
      11'h257: dout  = 8'b00000000; //  599 :   0 - 0x0
      11'h258: dout  = 8'b00000000; //  600 :   0 - 0x0 -- Background 0x4b
      11'h259: dout  = 8'b00000000; //  601 :   0 - 0x0
      11'h25A: dout  = 8'b00000000; //  602 :   0 - 0x0
      11'h25B: dout  = 8'b00000000; //  603 :   0 - 0x0
      11'h25C: dout  = 8'b00000000; //  604 :   0 - 0x0
      11'h25D: dout  = 8'b00000000; //  605 :   0 - 0x0
      11'h25E: dout  = 8'b00000000; //  606 :   0 - 0x0
      11'h25F: dout  = 8'b00000000; //  607 :   0 - 0x0
      11'h260: dout  = 8'b00000000; //  608 :   0 - 0x0 -- Background 0x4c
      11'h261: dout  = 8'b00000000; //  609 :   0 - 0x0
      11'h262: dout  = 8'b00000000; //  610 :   0 - 0x0
      11'h263: dout  = 8'b00000000; //  611 :   0 - 0x0
      11'h264: dout  = 8'b00000000; //  612 :   0 - 0x0
      11'h265: dout  = 8'b00000000; //  613 :   0 - 0x0
      11'h266: dout  = 8'b00000000; //  614 :   0 - 0x0
      11'h267: dout  = 8'b00000000; //  615 :   0 - 0x0
      11'h268: dout  = 8'b00000000; //  616 :   0 - 0x0 -- Background 0x4d
      11'h269: dout  = 8'b00000000; //  617 :   0 - 0x0
      11'h26A: dout  = 8'b00000000; //  618 :   0 - 0x0
      11'h26B: dout  = 8'b00000000; //  619 :   0 - 0x0
      11'h26C: dout  = 8'b00000000; //  620 :   0 - 0x0
      11'h26D: dout  = 8'b00000000; //  621 :   0 - 0x0
      11'h26E: dout  = 8'b00000000; //  622 :   0 - 0x0
      11'h26F: dout  = 8'b00000000; //  623 :   0 - 0x0
      11'h270: dout  = 8'b00000000; //  624 :   0 - 0x0 -- Background 0x4e
      11'h271: dout  = 8'b00000000; //  625 :   0 - 0x0
      11'h272: dout  = 8'b00000000; //  626 :   0 - 0x0
      11'h273: dout  = 8'b00000000; //  627 :   0 - 0x0
      11'h274: dout  = 8'b00000000; //  628 :   0 - 0x0
      11'h275: dout  = 8'b00000000; //  629 :   0 - 0x0
      11'h276: dout  = 8'b00000000; //  630 :   0 - 0x0
      11'h277: dout  = 8'b00000000; //  631 :   0 - 0x0
      11'h278: dout  = 8'b00000000; //  632 :   0 - 0x0 -- Background 0x4f
      11'h279: dout  = 8'b00000000; //  633 :   0 - 0x0
      11'h27A: dout  = 8'b00000000; //  634 :   0 - 0x0
      11'h27B: dout  = 8'b00000000; //  635 :   0 - 0x0
      11'h27C: dout  = 8'b00000000; //  636 :   0 - 0x0
      11'h27D: dout  = 8'b00000000; //  637 :   0 - 0x0
      11'h27E: dout  = 8'b00000000; //  638 :   0 - 0x0
      11'h27F: dout  = 8'b00000000; //  639 :   0 - 0x0
      11'h280: dout  = 8'b00000000; //  640 :   0 - 0x0 -- Background 0x50
      11'h281: dout  = 8'b00111111; //  641 :  63 - 0x3f
      11'h282: dout  = 8'b01111111; //  642 : 127 - 0x7f
      11'h283: dout  = 8'b01111111; //  643 : 127 - 0x7f
      11'h284: dout  = 8'b01111111; //  644 : 127 - 0x7f
      11'h285: dout  = 8'b00111100; //  645 :  60 - 0x3c
      11'h286: dout  = 8'b00000000; //  646 :   0 - 0x0
      11'h287: dout  = 8'b01000000; //  647 :  64 - 0x40
      11'h288: dout  = 8'b00000000; //  648 :   0 - 0x0 -- Background 0x51
      11'h289: dout  = 8'b11111100; //  649 : 252 - 0xfc
      11'h28A: dout  = 8'b11111110; //  650 : 254 - 0xfe
      11'h28B: dout  = 8'b11111110; //  651 : 254 - 0xfe
      11'h28C: dout  = 8'b11111110; //  652 : 254 - 0xfe
      11'h28D: dout  = 8'b00111100; //  653 :  60 - 0x3c
      11'h28E: dout  = 8'b00000000; //  654 :   0 - 0x0
      11'h28F: dout  = 8'b00000010; //  655 :   2 - 0x2
      11'h290: dout  = 8'b00000000; //  656 :   0 - 0x0 -- Background 0x52
      11'h291: dout  = 8'b00000000; //  657 :   0 - 0x0
      11'h292: dout  = 8'b00000011; //  658 :   3 - 0x3
      11'h293: dout  = 8'b00000111; //  659 :   7 - 0x7
      11'h294: dout  = 8'b00001111; //  660 :  15 - 0xf
      11'h295: dout  = 8'b00011111; //  661 :  31 - 0x1f
      11'h296: dout  = 8'b00111111; //  662 :  63 - 0x3f
      11'h297: dout  = 8'b00110000; //  663 :  48 - 0x30
      11'h298: dout  = 8'b00000000; //  664 :   0 - 0x0 -- Background 0x53
      11'h299: dout  = 8'b00000000; //  665 :   0 - 0x0
      11'h29A: dout  = 8'b10100000; //  666 : 160 - 0xa0
      11'h29B: dout  = 8'b10110000; //  667 : 176 - 0xb0
      11'h29C: dout  = 8'b10110000; //  668 : 176 - 0xb0
      11'h29D: dout  = 8'b10111000; //  669 : 184 - 0xb8
      11'h29E: dout  = 8'b01111100; //  670 : 124 - 0x7c
      11'h29F: dout  = 8'b01111100; //  671 : 124 - 0x7c
      11'h2A0: dout  = 8'b00000000; //  672 :   0 - 0x0 -- Background 0x54
      11'h2A1: dout  = 8'b00100001; //  673 :  33 - 0x21
      11'h2A2: dout  = 8'b01110001; //  674 : 113 - 0x71
      11'h2A3: dout  = 8'b00111010; //  675 :  58 - 0x3a
      11'h2A4: dout  = 8'b01101101; //  676 : 109 - 0x6d
      11'h2A5: dout  = 8'b00111000; //  677 :  56 - 0x38
      11'h2A6: dout  = 8'b00011101; //  678 :  29 - 0x1d
      11'h2A7: dout  = 8'b00101111; //  679 :  47 - 0x2f
      11'h2A8: dout  = 8'b00000000; //  680 :   0 - 0x0 -- Background 0x55
      11'h2A9: dout  = 8'b00100001; //  681 :  33 - 0x21
      11'h2AA: dout  = 8'b01110001; //  682 : 113 - 0x71
      11'h2AB: dout  = 8'b00111010; //  683 :  58 - 0x3a
      11'h2AC: dout  = 8'b01101101; //  684 : 109 - 0x6d
      11'h2AD: dout  = 8'b10111000; //  685 : 184 - 0xb8
      11'h2AE: dout  = 8'b00011101; //  686 :  29 - 0x1d
      11'h2AF: dout  = 8'b10101111; //  687 : 175 - 0xaf
      11'h2B0: dout  = 8'b00000000; //  688 :   0 - 0x0 -- Background 0x56
      11'h2B1: dout  = 8'b00100000; //  689 :  32 - 0x20
      11'h2B2: dout  = 8'b01110000; //  690 : 112 - 0x70
      11'h2B3: dout  = 8'b00111010; //  691 :  58 - 0x3a
      11'h2B4: dout  = 8'b01101100; //  692 : 108 - 0x6c
      11'h2B5: dout  = 8'b10111000; //  693 : 184 - 0xb8
      11'h2B6: dout  = 8'b00011100; //  694 :  28 - 0x1c
      11'h2B7: dout  = 8'b10101110; //  695 : 174 - 0xae
      11'h2B8: dout  = 8'b00000000; //  696 :   0 - 0x0 -- Background 0x57
      11'h2B9: dout  = 8'b01111111; //  697 : 127 - 0x7f
      11'h2BA: dout  = 8'b01001100; //  698 :  76 - 0x4c
      11'h2BB: dout  = 8'b00110011; //  699 :  51 - 0x33
      11'h2BC: dout  = 8'b00000000; //  700 :   0 - 0x0
      11'h2BD: dout  = 8'b00000000; //  701 :   0 - 0x0
      11'h2BE: dout  = 8'b00000000; //  702 :   0 - 0x0
      11'h2BF: dout  = 8'b00000000; //  703 :   0 - 0x0
      11'h2C0: dout  = 8'b00000000; //  704 :   0 - 0x0 -- Background 0x58
      11'h2C1: dout  = 8'b11111111; //  705 : 255 - 0xff
      11'h2C2: dout  = 8'b11001100; //  706 : 204 - 0xcc
      11'h2C3: dout  = 8'b00110011; //  707 :  51 - 0x33
      11'h2C4: dout  = 8'b11001100; //  708 : 204 - 0xcc
      11'h2C5: dout  = 8'b00000000; //  709 :   0 - 0x0
      11'h2C6: dout  = 8'b00000000; //  710 :   0 - 0x0
      11'h2C7: dout  = 8'b00000000; //  711 :   0 - 0x0
      11'h2C8: dout  = 8'b00000000; //  712 :   0 - 0x0 -- Background 0x59
      11'h2C9: dout  = 8'b11111110; //  713 : 254 - 0xfe
      11'h2CA: dout  = 8'b11001100; //  714 : 204 - 0xcc
      11'h2CB: dout  = 8'b00110000; //  715 :  48 - 0x30
      11'h2CC: dout  = 8'b11000000; //  716 : 192 - 0xc0
      11'h2CD: dout  = 8'b00000000; //  717 :   0 - 0x0
      11'h2CE: dout  = 8'b00000000; //  718 :   0 - 0x0
      11'h2CF: dout  = 8'b00000000; //  719 :   0 - 0x0
      11'h2D0: dout  = 8'b00000000; //  720 :   0 - 0x0 -- Background 0x5a
      11'h2D1: dout  = 8'b00000000; //  721 :   0 - 0x0
      11'h2D2: dout  = 8'b00000000; //  722 :   0 - 0x0
      11'h2D3: dout  = 8'b00000000; //  723 :   0 - 0x0
      11'h2D4: dout  = 8'b00000000; //  724 :   0 - 0x0
      11'h2D5: dout  = 8'b00000000; //  725 :   0 - 0x0
      11'h2D6: dout  = 8'b00000000; //  726 :   0 - 0x0
      11'h2D7: dout  = 8'b00000000; //  727 :   0 - 0x0
      11'h2D8: dout  = 8'b00000000; //  728 :   0 - 0x0 -- Background 0x5b
      11'h2D9: dout  = 8'b00000000; //  729 :   0 - 0x0
      11'h2DA: dout  = 8'b00000000; //  730 :   0 - 0x0
      11'h2DB: dout  = 8'b00000000; //  731 :   0 - 0x0
      11'h2DC: dout  = 8'b00000001; //  732 :   1 - 0x1
      11'h2DD: dout  = 8'b00000001; //  733 :   1 - 0x1
      11'h2DE: dout  = 8'b00000011; //  734 :   3 - 0x3
      11'h2DF: dout  = 8'b00000011; //  735 :   3 - 0x3
      11'h2E0: dout  = 8'b00000000; //  736 :   0 - 0x0 -- Background 0x5c
      11'h2E1: dout  = 8'b00000000; //  737 :   0 - 0x0
      11'h2E2: dout  = 8'b00000001; //  738 :   1 - 0x1
      11'h2E3: dout  = 8'b01111110; //  739 : 126 - 0x7e
      11'h2E4: dout  = 8'b11111111; //  740 : 255 - 0xff
      11'h2E5: dout  = 8'b11111111; //  741 : 255 - 0xff
      11'h2E6: dout  = 8'b11111111; //  742 : 255 - 0xff
      11'h2E7: dout  = 8'b11111111; //  743 : 255 - 0xff
      11'h2E8: dout  = 8'b00000000; //  744 :   0 - 0x0 -- Background 0x5d
      11'h2E9: dout  = 8'b11111111; //  745 : 255 - 0xff
      11'h2EA: dout  = 8'b11111111; //  746 : 255 - 0xff
      11'h2EB: dout  = 8'b11111111; //  747 : 255 - 0xff
      11'h2EC: dout  = 8'b01111111; //  748 : 127 - 0x7f
      11'h2ED: dout  = 8'b11111111; //  749 : 255 - 0xff
      11'h2EE: dout  = 8'b11111111; //  750 : 255 - 0xff
      11'h2EF: dout  = 8'b11111111; //  751 : 255 - 0xff
      11'h2F0: dout  = 8'b00000000; //  752 :   0 - 0x0 -- Background 0x5e
      11'h2F1: dout  = 8'b00000000; //  753 :   0 - 0x0
      11'h2F2: dout  = 8'b10000000; //  754 : 128 - 0x80
      11'h2F3: dout  = 8'b01111110; //  755 : 126 - 0x7e
      11'h2F4: dout  = 8'b10111111; //  756 : 191 - 0xbf
      11'h2F5: dout  = 8'b11111111; //  757 : 255 - 0xff
      11'h2F6: dout  = 8'b11111111; //  758 : 255 - 0xff
      11'h2F7: dout  = 8'b11111111; //  759 : 255 - 0xff
      11'h2F8: dout  = 8'b00000000; //  760 :   0 - 0x0 -- Background 0x5f
      11'h2F9: dout  = 8'b00000000; //  761 :   0 - 0x0
      11'h2FA: dout  = 8'b00000000; //  762 :   0 - 0x0
      11'h2FB: dout  = 8'b00000000; //  763 :   0 - 0x0
      11'h2FC: dout  = 8'b10000000; //  764 : 128 - 0x80
      11'h2FD: dout  = 8'b10000000; //  765 : 128 - 0x80
      11'h2FE: dout  = 8'b11000000; //  766 : 192 - 0xc0
      11'h2FF: dout  = 8'b11000000; //  767 : 192 - 0xc0
      11'h300: dout  = 8'b01111111; //  768 : 127 - 0x7f -- Background 0x60
      11'h301: dout  = 8'b01111111; //  769 : 127 - 0x7f
      11'h302: dout  = 8'b01111101; //  770 : 125 - 0x7d
      11'h303: dout  = 8'b01111111; //  771 : 127 - 0x7f
      11'h304: dout  = 8'b00111111; //  772 :  63 - 0x3f
      11'h305: dout  = 8'b01111111; //  773 : 127 - 0x7f
      11'h306: dout  = 8'b01111111; //  774 : 127 - 0x7f
      11'h307: dout  = 8'b01110111; //  775 : 119 - 0x77
      11'h308: dout  = 8'b11111110; //  776 : 254 - 0xfe -- Background 0x61
      11'h309: dout  = 8'b11111110; //  777 : 254 - 0xfe
      11'h30A: dout  = 8'b11111100; //  778 : 252 - 0xfc
      11'h30B: dout  = 8'b11111110; //  779 : 254 - 0xfe
      11'h30C: dout  = 8'b10111110; //  780 : 190 - 0xbe
      11'h30D: dout  = 8'b11111110; //  781 : 254 - 0xfe
      11'h30E: dout  = 8'b11111110; //  782 : 254 - 0xfe
      11'h30F: dout  = 8'b11110110; //  783 : 246 - 0xf6
      11'h310: dout  = 8'b00000111; //  784 :   7 - 0x7 -- Background 0x62
      11'h311: dout  = 8'b00011111; //  785 :  31 - 0x1f
      11'h312: dout  = 8'b00111111; //  786 :  63 - 0x3f
      11'h313: dout  = 8'b00111111; //  787 :  63 - 0x3f
      11'h314: dout  = 8'b00111111; //  788 :  63 - 0x3f
      11'h315: dout  = 8'b00011111; //  789 :  31 - 0x1f
      11'h316: dout  = 8'b00001111; //  790 :  15 - 0xf
      11'h317: dout  = 8'b00000000; //  791 :   0 - 0x0
      11'h318: dout  = 8'b01111110; //  792 : 126 - 0x7e -- Background 0x63
      11'h319: dout  = 8'b01111100; //  793 : 124 - 0x7c
      11'h31A: dout  = 8'b00111110; //  794 :  62 - 0x3e
      11'h31B: dout  = 8'b10111100; //  795 : 188 - 0xbc
      11'h31C: dout  = 8'b10111110; //  796 : 190 - 0xbe
      11'h31D: dout  = 8'b10011100; //  797 : 156 - 0x9c
      11'h31E: dout  = 8'b11011000; //  798 : 216 - 0xd8
      11'h31F: dout  = 8'b00000000; //  799 :   0 - 0x0
      11'h320: dout  = 8'b01000110; //  800 :  70 - 0x46 -- Background 0x64
      11'h321: dout  = 8'b01101011; //  801 : 107 - 0x6b
      11'h322: dout  = 8'b01110001; //  802 : 113 - 0x71
      11'h323: dout  = 8'b00111010; //  803 :  58 - 0x3a
      11'h324: dout  = 8'b01101101; //  804 : 109 - 0x6d
      11'h325: dout  = 8'b00111000; //  805 :  56 - 0x38
      11'h326: dout  = 8'b00011101; //  806 :  29 - 0x1d
      11'h327: dout  = 8'b00101111; //  807 :  47 - 0x2f
      11'h328: dout  = 8'b01000110; //  808 :  70 - 0x46 -- Background 0x65
      11'h329: dout  = 8'b11101011; //  809 : 235 - 0xeb
      11'h32A: dout  = 8'b01110001; //  810 : 113 - 0x71
      11'h32B: dout  = 8'b00111010; //  811 :  58 - 0x3a
      11'h32C: dout  = 8'b01101101; //  812 : 109 - 0x6d
      11'h32D: dout  = 8'b10111000; //  813 : 184 - 0xb8
      11'h32E: dout  = 8'b00011101; //  814 :  29 - 0x1d
      11'h32F: dout  = 8'b10101111; //  815 : 175 - 0xaf
      11'h330: dout  = 8'b01000110; //  816 :  70 - 0x46 -- Background 0x66
      11'h331: dout  = 8'b11101010; //  817 : 234 - 0xea
      11'h332: dout  = 8'b01110000; //  818 : 112 - 0x70
      11'h333: dout  = 8'b00111010; //  819 :  58 - 0x3a
      11'h334: dout  = 8'b01101100; //  820 : 108 - 0x6c
      11'h335: dout  = 8'b10111000; //  821 : 184 - 0xb8
      11'h336: dout  = 8'b00011100; //  822 :  28 - 0x1c
      11'h337: dout  = 8'b10101110; //  823 : 174 - 0xae
      11'h338: dout  = 8'b00000000; //  824 :   0 - 0x0 -- Background 0x67
      11'h339: dout  = 8'b01111111; //  825 : 127 - 0x7f
      11'h33A: dout  = 8'b01111111; //  826 : 127 - 0x7f
      11'h33B: dout  = 8'b00110011; //  827 :  51 - 0x33
      11'h33C: dout  = 8'b00000000; //  828 :   0 - 0x0
      11'h33D: dout  = 8'b00000000; //  829 :   0 - 0x0
      11'h33E: dout  = 8'b00000000; //  830 :   0 - 0x0
      11'h33F: dout  = 8'b00000000; //  831 :   0 - 0x0
      11'h340: dout  = 8'b00000000; //  832 :   0 - 0x0 -- Background 0x68
      11'h341: dout  = 8'b11111111; //  833 : 255 - 0xff
      11'h342: dout  = 8'b11111111; //  834 : 255 - 0xff
      11'h343: dout  = 8'b11111111; //  835 : 255 - 0xff
      11'h344: dout  = 8'b11001100; //  836 : 204 - 0xcc
      11'h345: dout  = 8'b00000000; //  837 :   0 - 0x0
      11'h346: dout  = 8'b00000000; //  838 :   0 - 0x0
      11'h347: dout  = 8'b00000000; //  839 :   0 - 0x0
      11'h348: dout  = 8'b00000000; //  840 :   0 - 0x0 -- Background 0x69
      11'h349: dout  = 8'b11111110; //  841 : 254 - 0xfe
      11'h34A: dout  = 8'b11111110; //  842 : 254 - 0xfe
      11'h34B: dout  = 8'b11110000; //  843 : 240 - 0xf0
      11'h34C: dout  = 8'b11000000; //  844 : 192 - 0xc0
      11'h34D: dout  = 8'b00000000; //  845 :   0 - 0x0
      11'h34E: dout  = 8'b00000000; //  846 :   0 - 0x0
      11'h34F: dout  = 8'b00000000; //  847 :   0 - 0x0
      11'h350: dout  = 8'b00000000; //  848 :   0 - 0x0 -- Background 0x6a
      11'h351: dout  = 8'b00000000; //  849 :   0 - 0x0
      11'h352: dout  = 8'b00000000; //  850 :   0 - 0x0
      11'h353: dout  = 8'b00000000; //  851 :   0 - 0x0
      11'h354: dout  = 8'b00000000; //  852 :   0 - 0x0
      11'h355: dout  = 8'b00000000; //  853 :   0 - 0x0
      11'h356: dout  = 8'b00000000; //  854 :   0 - 0x0
      11'h357: dout  = 8'b00000000; //  855 :   0 - 0x0
      11'h358: dout  = 8'b00111101; //  856 :  61 - 0x3d -- Background 0x6b
      11'h359: dout  = 8'b01111111; //  857 : 127 - 0x7f
      11'h35A: dout  = 8'b01111111; //  858 : 127 - 0x7f
      11'h35B: dout  = 8'b01111111; //  859 : 127 - 0x7f
      11'h35C: dout  = 8'b00111111; //  860 :  63 - 0x3f
      11'h35D: dout  = 8'b00001111; //  861 :  15 - 0xf
      11'h35E: dout  = 8'b00000000; //  862 :   0 - 0x0
      11'h35F: dout  = 8'b00000000; //  863 :   0 - 0x0
      11'h360: dout  = 8'b11111111; //  864 : 255 - 0xff -- Background 0x6c
      11'h361: dout  = 8'b11111111; //  865 : 255 - 0xff
      11'h362: dout  = 8'b11111111; //  866 : 255 - 0xff
      11'h363: dout  = 8'b11111111; //  867 : 255 - 0xff
      11'h364: dout  = 8'b11111111; //  868 : 255 - 0xff
      11'h365: dout  = 8'b11111111; //  869 : 255 - 0xff
      11'h366: dout  = 8'b11111110; //  870 : 254 - 0xfe
      11'h367: dout  = 8'b00000000; //  871 :   0 - 0x0
      11'h368: dout  = 8'b00000000; //  872 :   0 - 0x0 -- Background 0x6d
      11'h369: dout  = 8'b00000000; //  873 :   0 - 0x0
      11'h36A: dout  = 8'b00000000; //  874 :   0 - 0x0
      11'h36B: dout  = 8'b00000000; //  875 :   0 - 0x0
      11'h36C: dout  = 8'b00000000; //  876 :   0 - 0x0
      11'h36D: dout  = 8'b00000000; //  877 :   0 - 0x0
      11'h36E: dout  = 8'b00000000; //  878 :   0 - 0x0
      11'h36F: dout  = 8'b00000000; //  879 :   0 - 0x0
      11'h370: dout  = 8'b00000000; //  880 :   0 - 0x0 -- Background 0x6e
      11'h371: dout  = 8'b00000000; //  881 :   0 - 0x0
      11'h372: dout  = 8'b00000000; //  882 :   0 - 0x0
      11'h373: dout  = 8'b00000000; //  883 :   0 - 0x0
      11'h374: dout  = 8'b00000000; //  884 :   0 - 0x0
      11'h375: dout  = 8'b00000000; //  885 :   0 - 0x0
      11'h376: dout  = 8'b00000000; //  886 :   0 - 0x0
      11'h377: dout  = 8'b00000000; //  887 :   0 - 0x0
      11'h378: dout  = 8'b10111000; //  888 : 184 - 0xb8 -- Background 0x6f
      11'h379: dout  = 8'b11111100; //  889 : 252 - 0xfc
      11'h37A: dout  = 8'b11111110; //  890 : 254 - 0xfe
      11'h37B: dout  = 8'b11111110; //  891 : 254 - 0xfe
      11'h37C: dout  = 8'b11111100; //  892 : 252 - 0xfc
      11'h37D: dout  = 8'b11110000; //  893 : 240 - 0xf0
      11'h37E: dout  = 8'b00000000; //  894 :   0 - 0x0
      11'h37F: dout  = 8'b00000000; //  895 :   0 - 0x0
      11'h380: dout  = 8'b00000000; //  896 :   0 - 0x0 -- Background 0x70
      11'h381: dout  = 8'b00111111; //  897 :  63 - 0x3f
      11'h382: dout  = 8'b01111111; //  898 : 127 - 0x7f
      11'h383: dout  = 8'b01111111; //  899 : 127 - 0x7f
      11'h384: dout  = 8'b00011100; //  900 :  28 - 0x1c
      11'h385: dout  = 8'b00000000; //  901 :   0 - 0x0
      11'h386: dout  = 8'b00000000; //  902 :   0 - 0x0
      11'h387: dout  = 8'b00000000; //  903 :   0 - 0x0
      11'h388: dout  = 8'b00000000; //  904 :   0 - 0x0 -- Background 0x71
      11'h389: dout  = 8'b11111111; //  905 : 255 - 0xff
      11'h38A: dout  = 8'b11111111; //  906 : 255 - 0xff
      11'h38B: dout  = 8'b11111111; //  907 : 255 - 0xff
      11'h38C: dout  = 8'b11111111; //  908 : 255 - 0xff
      11'h38D: dout  = 8'b00111100; //  909 :  60 - 0x3c
      11'h38E: dout  = 8'b00000000; //  910 :   0 - 0x0
      11'h38F: dout  = 8'b00000000; //  911 :   0 - 0x0
      11'h390: dout  = 8'b00000000; //  912 :   0 - 0x0 -- Background 0x72
      11'h391: dout  = 8'b11111100; //  913 : 252 - 0xfc
      11'h392: dout  = 8'b11111110; //  914 : 254 - 0xfe
      11'h393: dout  = 8'b11111110; //  915 : 254 - 0xfe
      11'h394: dout  = 8'b00111000; //  916 :  56 - 0x38
      11'h395: dout  = 8'b00000000; //  917 :   0 - 0x0
      11'h396: dout  = 8'b00000000; //  918 :   0 - 0x0
      11'h397: dout  = 8'b00000000; //  919 :   0 - 0x0
      11'h398: dout  = 8'b11111111; //  920 : 255 - 0xff -- Background 0x73
      11'h399: dout  = 8'b11111111; //  921 : 255 - 0xff
      11'h39A: dout  = 8'b11111101; //  922 : 253 - 0xfd
      11'h39B: dout  = 8'b11111111; //  923 : 255 - 0xff
      11'h39C: dout  = 8'b10111111; //  924 : 191 - 0xbf
      11'h39D: dout  = 8'b11111111; //  925 : 255 - 0xff
      11'h39E: dout  = 8'b11111111; //  926 : 255 - 0xff
      11'h39F: dout  = 8'b11110111; //  927 : 247 - 0xf7
      11'h3A0: dout  = 8'b01000110; //  928 :  70 - 0x46 -- Background 0x74
      11'h3A1: dout  = 8'b01101011; //  929 : 107 - 0x6b
      11'h3A2: dout  = 8'b01110001; //  930 : 113 - 0x71
      11'h3A3: dout  = 8'b00111010; //  931 :  58 - 0x3a
      11'h3A4: dout  = 8'b01101101; //  932 : 109 - 0x6d
      11'h3A5: dout  = 8'b00111000; //  933 :  56 - 0x38
      11'h3A6: dout  = 8'b00011101; //  934 :  29 - 0x1d
      11'h3A7: dout  = 8'b00000000; //  935 :   0 - 0x0
      11'h3A8: dout  = 8'b01000110; //  936 :  70 - 0x46 -- Background 0x75
      11'h3A9: dout  = 8'b11101011; //  937 : 235 - 0xeb
      11'h3AA: dout  = 8'b01110001; //  938 : 113 - 0x71
      11'h3AB: dout  = 8'b00111010; //  939 :  58 - 0x3a
      11'h3AC: dout  = 8'b01101101; //  940 : 109 - 0x6d
      11'h3AD: dout  = 8'b10111000; //  941 : 184 - 0xb8
      11'h3AE: dout  = 8'b00011101; //  942 :  29 - 0x1d
      11'h3AF: dout  = 8'b00000000; //  943 :   0 - 0x0
      11'h3B0: dout  = 8'b01000110; //  944 :  70 - 0x46 -- Background 0x76
      11'h3B1: dout  = 8'b11101010; //  945 : 234 - 0xea
      11'h3B2: dout  = 8'b01110000; //  946 : 112 - 0x70
      11'h3B3: dout  = 8'b00111010; //  947 :  58 - 0x3a
      11'h3B4: dout  = 8'b01101100; //  948 : 108 - 0x6c
      11'h3B5: dout  = 8'b10111000; //  949 : 184 - 0xb8
      11'h3B6: dout  = 8'b00011100; //  950 :  28 - 0x1c
      11'h3B7: dout  = 8'b00000000; //  951 :   0 - 0x0
      11'h3B8: dout  = 8'b10000001; //  952 : 129 - 0x81 -- Background 0x77
      11'h3B9: dout  = 8'b11111111; //  953 : 255 - 0xff
      11'h3BA: dout  = 8'b11111101; //  954 : 253 - 0xfd
      11'h3BB: dout  = 8'b11111111; //  955 : 255 - 0xff
      11'h3BC: dout  = 8'b10111111; //  956 : 191 - 0xbf
      11'h3BD: dout  = 8'b11111111; //  957 : 255 - 0xff
      11'h3BE: dout  = 8'b11111111; //  958 : 255 - 0xff
      11'h3BF: dout  = 8'b11110111; //  959 : 247 - 0xf7
      11'h3C0: dout  = 8'b00000000; //  960 :   0 - 0x0 -- Background 0x78
      11'h3C1: dout  = 8'b00000000; //  961 :   0 - 0x0
      11'h3C2: dout  = 8'b00000000; //  962 :   0 - 0x0
      11'h3C3: dout  = 8'b00000000; //  963 :   0 - 0x0
      11'h3C4: dout  = 8'b00000000; //  964 :   0 - 0x0
      11'h3C5: dout  = 8'b00000000; //  965 :   0 - 0x0
      11'h3C6: dout  = 8'b00000000; //  966 :   0 - 0x0
      11'h3C7: dout  = 8'b00000000; //  967 :   0 - 0x0
      11'h3C8: dout  = 8'b00000000; //  968 :   0 - 0x0 -- Background 0x79
      11'h3C9: dout  = 8'b00000000; //  969 :   0 - 0x0
      11'h3CA: dout  = 8'b00000000; //  970 :   0 - 0x0
      11'h3CB: dout  = 8'b00000000; //  971 :   0 - 0x0
      11'h3CC: dout  = 8'b00000000; //  972 :   0 - 0x0
      11'h3CD: dout  = 8'b00000000; //  973 :   0 - 0x0
      11'h3CE: dout  = 8'b00000000; //  974 :   0 - 0x0
      11'h3CF: dout  = 8'b00000000; //  975 :   0 - 0x0
      11'h3D0: dout  = 8'b00000000; //  976 :   0 - 0x0 -- Background 0x7a
      11'h3D1: dout  = 8'b00000000; //  977 :   0 - 0x0
      11'h3D2: dout  = 8'b00000000; //  978 :   0 - 0x0
      11'h3D3: dout  = 8'b00000000; //  979 :   0 - 0x0
      11'h3D4: dout  = 8'b00000000; //  980 :   0 - 0x0
      11'h3D5: dout  = 8'b00000000; //  981 :   0 - 0x0
      11'h3D6: dout  = 8'b00000000; //  982 :   0 - 0x0
      11'h3D7: dout  = 8'b00000000; //  983 :   0 - 0x0
      11'h3D8: dout  = 8'b00000000; //  984 :   0 - 0x0 -- Background 0x7b
      11'h3D9: dout  = 8'b00000000; //  985 :   0 - 0x0
      11'h3DA: dout  = 8'b00000000; //  986 :   0 - 0x0
      11'h3DB: dout  = 8'b00000000; //  987 :   0 - 0x0
      11'h3DC: dout  = 8'b00000000; //  988 :   0 - 0x0
      11'h3DD: dout  = 8'b00000000; //  989 :   0 - 0x0
      11'h3DE: dout  = 8'b00000000; //  990 :   0 - 0x0
      11'h3DF: dout  = 8'b00000000; //  991 :   0 - 0x0
      11'h3E0: dout  = 8'b00000000; //  992 :   0 - 0x0 -- Background 0x7c
      11'h3E1: dout  = 8'b00100010; //  993 :  34 - 0x22
      11'h3E2: dout  = 8'b01110111; //  994 : 119 - 0x77
      11'h3E3: dout  = 8'b11111111; //  995 : 255 - 0xff
      11'h3E4: dout  = 8'b11111011; //  996 : 251 - 0xfb
      11'h3E5: dout  = 8'b11110101; //  997 : 245 - 0xf5
      11'h3E6: dout  = 8'b11101111; //  998 : 239 - 0xef
      11'h3E7: dout  = 8'b11111111; //  999 : 255 - 0xff
      11'h3E8: dout  = 8'b00000000; // 1000 :   0 - 0x0 -- Background 0x7d
      11'h3E9: dout  = 8'b01110011; // 1001 : 115 - 0x73
      11'h3EA: dout  = 8'b11111111; // 1002 : 255 - 0xff
      11'h3EB: dout  = 8'b11111111; // 1003 : 255 - 0xff
      11'h3EC: dout  = 8'b11111011; // 1004 : 251 - 0xfb
      11'h3ED: dout  = 8'b11111101; // 1005 : 253 - 0xfd
      11'h3EE: dout  = 8'b11101111; // 1006 : 239 - 0xef
      11'h3EF: dout  = 8'b11111111; // 1007 : 255 - 0xff
      11'h3F0: dout  = 8'b11011111; // 1008 : 223 - 0xdf -- Background 0x7e
      11'h3F1: dout  = 8'b10101111; // 1009 : 175 - 0xaf
      11'h3F2: dout  = 8'b01111111; // 1010 : 127 - 0x7f
      11'h3F3: dout  = 8'b11111111; // 1011 : 255 - 0xff
      11'h3F4: dout  = 8'b11111011; // 1012 : 251 - 0xfb
      11'h3F5: dout  = 8'b11110101; // 1013 : 245 - 0xf5
      11'h3F6: dout  = 8'b11101111; // 1014 : 239 - 0xef
      11'h3F7: dout  = 8'b11111111; // 1015 : 255 - 0xff
      11'h3F8: dout  = 8'b00000000; // 1016 :   0 - 0x0 -- Background 0x7f
      11'h3F9: dout  = 8'b10101111; // 1017 : 175 - 0xaf
      11'h3FA: dout  = 8'b01111111; // 1018 : 127 - 0x7f
      11'h3FB: dout  = 8'b11111111; // 1019 : 255 - 0xff
      11'h3FC: dout  = 8'b11111011; // 1020 : 251 - 0xfb
      11'h3FD: dout  = 8'b11110101; // 1021 : 245 - 0xf5
      11'h3FE: dout  = 8'b11101111; // 1022 : 239 - 0xef
      11'h3FF: dout  = 8'b11111111; // 1023 : 255 - 0xff
      11'h400: dout  = 8'b00000000; // 1024 :   0 - 0x0 -- Background 0x80
      11'h401: dout  = 8'b01111111; // 1025 : 127 - 0x7f
      11'h402: dout  = 8'b00110000; // 1026 :  48 - 0x30
      11'h403: dout  = 8'b00110000; // 1027 :  48 - 0x30
      11'h404: dout  = 8'b00110000; // 1028 :  48 - 0x30
      11'h405: dout  = 8'b01111111; // 1029 : 127 - 0x7f
      11'h406: dout  = 8'b00110000; // 1030 :  48 - 0x30
      11'h407: dout  = 8'b00110000; // 1031 :  48 - 0x30
      11'h408: dout  = 8'b00000000; // 1032 :   0 - 0x0 -- Background 0x81
      11'h409: dout  = 8'b01111111; // 1033 : 127 - 0x7f
      11'h40A: dout  = 8'b00000000; // 1034 :   0 - 0x0
      11'h40B: dout  = 8'b01111111; // 1035 : 127 - 0x7f
      11'h40C: dout  = 8'b01111111; // 1036 : 127 - 0x7f
      11'h40D: dout  = 8'b00100000; // 1037 :  32 - 0x20
      11'h40E: dout  = 8'b01000000; // 1038 :  64 - 0x40
      11'h40F: dout  = 8'b00000000; // 1039 :   0 - 0x0
      11'h410: dout  = 8'b00000000; // 1040 :   0 - 0x0 -- Background 0x82
      11'h411: dout  = 8'b11111110; // 1041 : 254 - 0xfe
      11'h412: dout  = 8'b00001100; // 1042 :  12 - 0xc
      11'h413: dout  = 8'b00001100; // 1043 :  12 - 0xc
      11'h414: dout  = 8'b00001100; // 1044 :  12 - 0xc
      11'h415: dout  = 8'b11111110; // 1045 : 254 - 0xfe
      11'h416: dout  = 8'b00001100; // 1046 :  12 - 0xc
      11'h417: dout  = 8'b00001100; // 1047 :  12 - 0xc
      11'h418: dout  = 8'b00000000; // 1048 :   0 - 0x0 -- Background 0x83
      11'h419: dout  = 8'b11111111; // 1049 : 255 - 0xff
      11'h41A: dout  = 8'b00000000; // 1050 :   0 - 0x0
      11'h41B: dout  = 8'b11111111; // 1051 : 255 - 0xff
      11'h41C: dout  = 8'b11111111; // 1052 : 255 - 0xff
      11'h41D: dout  = 8'b00000000; // 1053 :   0 - 0x0
      11'h41E: dout  = 8'b00000000; // 1054 :   0 - 0x0
      11'h41F: dout  = 8'b00000000; // 1055 :   0 - 0x0
      11'h420: dout  = 8'b00000000; // 1056 :   0 - 0x0 -- Background 0x84
      11'h421: dout  = 8'b11111111; // 1057 : 255 - 0xff
      11'h422: dout  = 8'b11111111; // 1058 : 255 - 0xff
      11'h423: dout  = 8'b11111111; // 1059 : 255 - 0xff
      11'h424: dout  = 8'b11111111; // 1060 : 255 - 0xff
      11'h425: dout  = 8'b11101111; // 1061 : 239 - 0xef
      11'h426: dout  = 8'b10111011; // 1062 : 187 - 0xbb
      11'h427: dout  = 8'b00000000; // 1063 :   0 - 0x0
      11'h428: dout  = 8'b00000000; // 1064 :   0 - 0x0 -- Background 0x85
      11'h429: dout  = 8'b11111110; // 1065 : 254 - 0xfe
      11'h42A: dout  = 8'b00000000; // 1066 :   0 - 0x0
      11'h42B: dout  = 8'b11111110; // 1067 : 254 - 0xfe
      11'h42C: dout  = 8'b11111110; // 1068 : 254 - 0xfe
      11'h42D: dout  = 8'b00001100; // 1069 :  12 - 0xc
      11'h42E: dout  = 8'b00000010; // 1070 :   2 - 0x2
      11'h42F: dout  = 8'b00000000; // 1071 :   0 - 0x0
      11'h430: dout  = 8'b00000000; // 1072 :   0 - 0x0 -- Background 0x86
      11'h431: dout  = 8'b00000000; // 1073 :   0 - 0x0
      11'h432: dout  = 8'b00000000; // 1074 :   0 - 0x0
      11'h433: dout  = 8'b00000000; // 1075 :   0 - 0x0
      11'h434: dout  = 8'b00000000; // 1076 :   0 - 0x0
      11'h435: dout  = 8'b00000000; // 1077 :   0 - 0x0
      11'h436: dout  = 8'b00000000; // 1078 :   0 - 0x0
      11'h437: dout  = 8'b00000000; // 1079 :   0 - 0x0
      11'h438: dout  = 8'b00000000; // 1080 :   0 - 0x0 -- Background 0x87
      11'h439: dout  = 8'b00000000; // 1081 :   0 - 0x0
      11'h43A: dout  = 8'b00000000; // 1082 :   0 - 0x0
      11'h43B: dout  = 8'b00000000; // 1083 :   0 - 0x0
      11'h43C: dout  = 8'b00000000; // 1084 :   0 - 0x0
      11'h43D: dout  = 8'b00000000; // 1085 :   0 - 0x0
      11'h43E: dout  = 8'b00000000; // 1086 :   0 - 0x0
      11'h43F: dout  = 8'b00000000; // 1087 :   0 - 0x0
      11'h440: dout  = 8'b00000000; // 1088 :   0 - 0x0 -- Background 0x88
      11'h441: dout  = 8'b00000111; // 1089 :   7 - 0x7
      11'h442: dout  = 8'b00011111; // 1090 :  31 - 0x1f
      11'h443: dout  = 8'b00111100; // 1091 :  60 - 0x3c
      11'h444: dout  = 8'b00110001; // 1092 :  49 - 0x31
      11'h445: dout  = 8'b01110100; // 1093 : 116 - 0x74
      11'h446: dout  = 8'b01100101; // 1094 : 101 - 0x65
      11'h447: dout  = 8'b01101010; // 1095 : 106 - 0x6a
      11'h448: dout  = 8'b01100100; // 1096 : 100 - 0x64 -- Background 0x89
      11'h449: dout  = 8'b01101101; // 1097 : 109 - 0x6d
      11'h44A: dout  = 8'b01110010; // 1098 : 114 - 0x72
      11'h44B: dout  = 8'b00110000; // 1099 :  48 - 0x30
      11'h44C: dout  = 8'b00111100; // 1100 :  60 - 0x3c
      11'h44D: dout  = 8'b00011111; // 1101 :  31 - 0x1f
      11'h44E: dout  = 8'b00000111; // 1102 :   7 - 0x7
      11'h44F: dout  = 8'b00000000; // 1103 :   0 - 0x0
      11'h450: dout  = 8'b00000000; // 1104 :   0 - 0x0 -- Background 0x8a
      11'h451: dout  = 8'b11100000; // 1105 : 224 - 0xe0
      11'h452: dout  = 8'b11111000; // 1106 : 248 - 0xf8
      11'h453: dout  = 8'b00111100; // 1107 :  60 - 0x3c
      11'h454: dout  = 8'b01001100; // 1108 :  76 - 0x4c
      11'h455: dout  = 8'b01101110; // 1109 : 110 - 0x6e
      11'h456: dout  = 8'b00100110; // 1110 :  38 - 0x26
      11'h457: dout  = 8'b01000110; // 1111 :  70 - 0x46
      11'h458: dout  = 8'b10010110; // 1112 : 150 - 0x96 -- Background 0x8b
      11'h459: dout  = 8'b01100110; // 1113 : 102 - 0x66
      11'h45A: dout  = 8'b10101110; // 1114 : 174 - 0xae
      11'h45B: dout  = 8'b01001100; // 1115 :  76 - 0x4c
      11'h45C: dout  = 8'b00111100; // 1116 :  60 - 0x3c
      11'h45D: dout  = 8'b11111000; // 1117 : 248 - 0xf8
      11'h45E: dout  = 8'b11100000; // 1118 : 224 - 0xe0
      11'h45F: dout  = 8'b00000000; // 1119 :   0 - 0x0
      11'h460: dout  = 8'b00000000; // 1120 :   0 - 0x0 -- Background 0x8c
      11'h461: dout  = 8'b00000111; // 1121 :   7 - 0x7
      11'h462: dout  = 8'b00011111; // 1122 :  31 - 0x1f
      11'h463: dout  = 8'b00111111; // 1123 :  63 - 0x3f
      11'h464: dout  = 8'b00111111; // 1124 :  63 - 0x3f
      11'h465: dout  = 8'b01111111; // 1125 : 127 - 0x7f
      11'h466: dout  = 8'b01111111; // 1126 : 127 - 0x7f
      11'h467: dout  = 8'b01111111; // 1127 : 127 - 0x7f
      11'h468: dout  = 8'b01111111; // 1128 : 127 - 0x7f -- Background 0x8d
      11'h469: dout  = 8'b01111111; // 1129 : 127 - 0x7f
      11'h46A: dout  = 8'b01111111; // 1130 : 127 - 0x7f
      11'h46B: dout  = 8'b00111111; // 1131 :  63 - 0x3f
      11'h46C: dout  = 8'b00111111; // 1132 :  63 - 0x3f
      11'h46D: dout  = 8'b00011111; // 1133 :  31 - 0x1f
      11'h46E: dout  = 8'b00000111; // 1134 :   7 - 0x7
      11'h46F: dout  = 8'b00000000; // 1135 :   0 - 0x0
      11'h470: dout  = 8'b00000000; // 1136 :   0 - 0x0 -- Background 0x8e
      11'h471: dout  = 8'b11100000; // 1137 : 224 - 0xe0
      11'h472: dout  = 8'b11111000; // 1138 : 248 - 0xf8
      11'h473: dout  = 8'b11111100; // 1139 : 252 - 0xfc
      11'h474: dout  = 8'b11111100; // 1140 : 252 - 0xfc
      11'h475: dout  = 8'b11111110; // 1141 : 254 - 0xfe
      11'h476: dout  = 8'b11111110; // 1142 : 254 - 0xfe
      11'h477: dout  = 8'b11111110; // 1143 : 254 - 0xfe
      11'h478: dout  = 8'b11111110; // 1144 : 254 - 0xfe -- Background 0x8f
      11'h479: dout  = 8'b11111110; // 1145 : 254 - 0xfe
      11'h47A: dout  = 8'b11111110; // 1146 : 254 - 0xfe
      11'h47B: dout  = 8'b11111100; // 1147 : 252 - 0xfc
      11'h47C: dout  = 8'b11111100; // 1148 : 252 - 0xfc
      11'h47D: dout  = 8'b11111000; // 1149 : 248 - 0xf8
      11'h47E: dout  = 8'b11100000; // 1150 : 224 - 0xe0
      11'h47F: dout  = 8'b00000000; // 1151 :   0 - 0x0
      11'h480: dout  = 8'b00000000; // 1152 :   0 - 0x0 -- Background 0x90
      11'h481: dout  = 8'b00000000; // 1153 :   0 - 0x0
      11'h482: dout  = 8'b00000000; // 1154 :   0 - 0x0
      11'h483: dout  = 8'b00000000; // 1155 :   0 - 0x0
      11'h484: dout  = 8'b00010000; // 1156 :  16 - 0x10
      11'h485: dout  = 8'b00011100; // 1157 :  28 - 0x1c
      11'h486: dout  = 8'b00001110; // 1158 :  14 - 0xe
      11'h487: dout  = 8'b00000111; // 1159 :   7 - 0x7
      11'h488: dout  = 8'b00000011; // 1160 :   3 - 0x3 -- Background 0x91
      11'h489: dout  = 8'b00000001; // 1161 :   1 - 0x1
      11'h48A: dout  = 8'b00110000; // 1162 :  48 - 0x30
      11'h48B: dout  = 8'b00001111; // 1163 :  15 - 0xf
      11'h48C: dout  = 8'b00000011; // 1164 :   3 - 0x3
      11'h48D: dout  = 8'b00000000; // 1165 :   0 - 0x0
      11'h48E: dout  = 8'b01111111; // 1166 : 127 - 0x7f
      11'h48F: dout  = 8'b00000000; // 1167 :   0 - 0x0
      11'h490: dout  = 8'b00000000; // 1168 :   0 - 0x0 -- Background 0x92
      11'h491: dout  = 8'b01000010; // 1169 :  66 - 0x42
      11'h492: dout  = 8'b01000010; // 1170 :  66 - 0x42
      11'h493: dout  = 8'b01100110; // 1171 : 102 - 0x66
      11'h494: dout  = 8'b01100110; // 1172 : 102 - 0x66
      11'h495: dout  = 8'b01100110; // 1173 : 102 - 0x66
      11'h496: dout  = 8'b11111110; // 1174 : 254 - 0xfe
      11'h497: dout  = 8'b11111111; // 1175 : 255 - 0xff
      11'h498: dout  = 8'b01111110; // 1176 : 126 - 0x7e -- Background 0x93
      11'h499: dout  = 8'b01111110; // 1177 : 126 - 0x7e
      11'h49A: dout  = 8'b01111110; // 1178 : 126 - 0x7e
      11'h49B: dout  = 8'b01111110; // 1179 : 126 - 0x7e
      11'h49C: dout  = 8'b01111110; // 1180 : 126 - 0x7e
      11'h49D: dout  = 8'b01111110; // 1181 : 126 - 0x7e
      11'h49E: dout  = 8'b01111110; // 1182 : 126 - 0x7e
      11'h49F: dout  = 8'b01111110; // 1183 : 126 - 0x7e
      11'h4A0: dout  = 8'b00000000; // 1184 :   0 - 0x0 -- Background 0x94
      11'h4A1: dout  = 8'b00000000; // 1185 :   0 - 0x0
      11'h4A2: dout  = 8'b00000000; // 1186 :   0 - 0x0
      11'h4A3: dout  = 8'b00000000; // 1187 :   0 - 0x0
      11'h4A4: dout  = 8'b00001000; // 1188 :   8 - 0x8
      11'h4A5: dout  = 8'b00111000; // 1189 :  56 - 0x38
      11'h4A6: dout  = 8'b01110000; // 1190 : 112 - 0x70
      11'h4A7: dout  = 8'b11100000; // 1191 : 224 - 0xe0
      11'h4A8: dout  = 8'b11000000; // 1192 : 192 - 0xc0 -- Background 0x95
      11'h4A9: dout  = 8'b10000000; // 1193 : 128 - 0x80
      11'h4AA: dout  = 8'b00001100; // 1194 :  12 - 0xc
      11'h4AB: dout  = 8'b11110000; // 1195 : 240 - 0xf0
      11'h4AC: dout  = 8'b11000000; // 1196 : 192 - 0xc0
      11'h4AD: dout  = 8'b00000000; // 1197 :   0 - 0x0
      11'h4AE: dout  = 8'b11111110; // 1198 : 254 - 0xfe
      11'h4AF: dout  = 8'b00000000; // 1199 :   0 - 0x0
      11'h4B0: dout  = 8'b00000000; // 1200 :   0 - 0x0 -- Background 0x96
      11'h4B1: dout  = 8'b00111111; // 1201 :  63 - 0x3f
      11'h4B2: dout  = 8'b01111111; // 1202 : 127 - 0x7f
      11'h4B3: dout  = 8'b01111111; // 1203 : 127 - 0x7f
      11'h4B4: dout  = 8'b01111111; // 1204 : 127 - 0x7f
      11'h4B5: dout  = 8'b01111111; // 1205 : 127 - 0x7f
      11'h4B6: dout  = 8'b01111111; // 1206 : 127 - 0x7f
      11'h4B7: dout  = 8'b01111111; // 1207 : 127 - 0x7f
      11'h4B8: dout  = 8'b01111111; // 1208 : 127 - 0x7f -- Background 0x97
      11'h4B9: dout  = 8'b01111111; // 1209 : 127 - 0x7f
      11'h4BA: dout  = 8'b00111111; // 1210 :  63 - 0x3f
      11'h4BB: dout  = 8'b01111111; // 1211 : 127 - 0x7f
      11'h4BC: dout  = 8'b01111111; // 1212 : 127 - 0x7f
      11'h4BD: dout  = 8'b01111111; // 1213 : 127 - 0x7f
      11'h4BE: dout  = 8'b01111111; // 1214 : 127 - 0x7f
      11'h4BF: dout  = 8'b01111111; // 1215 : 127 - 0x7f
      11'h4C0: dout  = 8'b00000000; // 1216 :   0 - 0x0 -- Background 0x98
      11'h4C1: dout  = 8'b11011111; // 1217 : 223 - 0xdf
      11'h4C2: dout  = 8'b11111111; // 1218 : 255 - 0xff
      11'h4C3: dout  = 8'b11111111; // 1219 : 255 - 0xff
      11'h4C4: dout  = 8'b11111111; // 1220 : 255 - 0xff
      11'h4C5: dout  = 8'b11111111; // 1221 : 255 - 0xff
      11'h4C6: dout  = 8'b11111111; // 1222 : 255 - 0xff
      11'h4C7: dout  = 8'b11111111; // 1223 : 255 - 0xff
      11'h4C8: dout  = 8'b11111111; // 1224 : 255 - 0xff -- Background 0x99
      11'h4C9: dout  = 8'b11111111; // 1225 : 255 - 0xff
      11'h4CA: dout  = 8'b10111111; // 1226 : 191 - 0xbf
      11'h4CB: dout  = 8'b11111111; // 1227 : 255 - 0xff
      11'h4CC: dout  = 8'b11111111; // 1228 : 255 - 0xff
      11'h4CD: dout  = 8'b11111111; // 1229 : 255 - 0xff
      11'h4CE: dout  = 8'b11111111; // 1230 : 255 - 0xff
      11'h4CF: dout  = 8'b11111111; // 1231 : 255 - 0xff
      11'h4D0: dout  = 8'b00000000; // 1232 :   0 - 0x0 -- Background 0x9a
      11'h4D1: dout  = 8'b10111100; // 1233 : 188 - 0xbc
      11'h4D2: dout  = 8'b11111110; // 1234 : 254 - 0xfe
      11'h4D3: dout  = 8'b11111110; // 1235 : 254 - 0xfe
      11'h4D4: dout  = 8'b11111110; // 1236 : 254 - 0xfe
      11'h4D5: dout  = 8'b11111110; // 1237 : 254 - 0xfe
      11'h4D6: dout  = 8'b11111110; // 1238 : 254 - 0xfe
      11'h4D7: dout  = 8'b11111110; // 1239 : 254 - 0xfe
      11'h4D8: dout  = 8'b11111110; // 1240 : 254 - 0xfe -- Background 0x9b
      11'h4D9: dout  = 8'b11111110; // 1241 : 254 - 0xfe
      11'h4DA: dout  = 8'b10111110; // 1242 : 190 - 0xbe
      11'h4DB: dout  = 8'b11111110; // 1243 : 254 - 0xfe
      11'h4DC: dout  = 8'b11111110; // 1244 : 254 - 0xfe
      11'h4DD: dout  = 8'b11111110; // 1245 : 254 - 0xfe
      11'h4DE: dout  = 8'b11111110; // 1246 : 254 - 0xfe
      11'h4DF: dout  = 8'b11111110; // 1247 : 254 - 0xfe
      11'h4E0: dout  = 8'b00000000; // 1248 :   0 - 0x0 -- Background 0x9c
      11'h4E1: dout  = 8'b00111111; // 1249 :  63 - 0x3f
      11'h4E2: dout  = 8'b01011111; // 1250 :  95 - 0x5f
      11'h4E3: dout  = 8'b01101111; // 1251 : 111 - 0x6f
      11'h4E4: dout  = 8'b01110111; // 1252 : 119 - 0x77
      11'h4E5: dout  = 8'b01111011; // 1253 : 123 - 0x7b
      11'h4E6: dout  = 8'b00010101; // 1254 :  21 - 0x15
      11'h4E7: dout  = 8'b00000000; // 1255 :   0 - 0x0
      11'h4E8: dout  = 8'b00000000; // 1256 :   0 - 0x0 -- Background 0x9d
      11'h4E9: dout  = 8'b10111110; // 1257 : 190 - 0xbe
      11'h4EA: dout  = 8'b11011110; // 1258 : 222 - 0xde
      11'h4EB: dout  = 8'b11101110; // 1259 : 238 - 0xee
      11'h4EC: dout  = 8'b11110110; // 1260 : 246 - 0xf6
      11'h4ED: dout  = 8'b11111010; // 1261 : 250 - 0xfa
      11'h4EE: dout  = 8'b01010100; // 1262 :  84 - 0x54
      11'h4EF: dout  = 8'b00000000; // 1263 :   0 - 0x0
      11'h4F0: dout  = 8'b00000000; // 1264 :   0 - 0x0 -- Background 0x9e
      11'h4F1: dout  = 8'b10111111; // 1265 : 191 - 0xbf
      11'h4F2: dout  = 8'b11011111; // 1266 : 223 - 0xdf
      11'h4F3: dout  = 8'b11101111; // 1267 : 239 - 0xef
      11'h4F4: dout  = 8'b11110111; // 1268 : 247 - 0xf7
      11'h4F5: dout  = 8'b11111011; // 1269 : 251 - 0xfb
      11'h4F6: dout  = 8'b01010101; // 1270 :  85 - 0x55
      11'h4F7: dout  = 8'b00000000; // 1271 :   0 - 0x0
      11'h4F8: dout  = 8'b00000000; // 1272 :   0 - 0x0 -- Background 0x9f
      11'h4F9: dout  = 8'b00000000; // 1273 :   0 - 0x0
      11'h4FA: dout  = 8'b00000000; // 1274 :   0 - 0x0
      11'h4FB: dout  = 8'b00000000; // 1275 :   0 - 0x0
      11'h4FC: dout  = 8'b00000000; // 1276 :   0 - 0x0
      11'h4FD: dout  = 8'b00000000; // 1277 :   0 - 0x0
      11'h4FE: dout  = 8'b00000000; // 1278 :   0 - 0x0
      11'h4FF: dout  = 8'b00000000; // 1279 :   0 - 0x0
      11'h500: dout  = 8'b00000000; // 1280 :   0 - 0x0 -- Background 0xa0
      11'h501: dout  = 8'b01111111; // 1281 : 127 - 0x7f
      11'h502: dout  = 8'b00000000; // 1282 :   0 - 0x0
      11'h503: dout  = 8'b00000001; // 1283 :   1 - 0x1
      11'h504: dout  = 8'b00000001; // 1284 :   1 - 0x1
      11'h505: dout  = 8'b00000001; // 1285 :   1 - 0x1
      11'h506: dout  = 8'b00000001; // 1286 :   1 - 0x1
      11'h507: dout  = 8'b00000001; // 1287 :   1 - 0x1
      11'h508: dout  = 8'b00000001; // 1288 :   1 - 0x1 -- Background 0xa1
      11'h509: dout  = 8'b00000001; // 1289 :   1 - 0x1
      11'h50A: dout  = 8'b00000001; // 1290 :   1 - 0x1
      11'h50B: dout  = 8'b00000001; // 1291 :   1 - 0x1
      11'h50C: dout  = 8'b00000001; // 1292 :   1 - 0x1
      11'h50D: dout  = 8'b00000001; // 1293 :   1 - 0x1
      11'h50E: dout  = 8'b00000001; // 1294 :   1 - 0x1
      11'h50F: dout  = 8'b00000001; // 1295 :   1 - 0x1
      11'h510: dout  = 8'b00000000; // 1296 :   0 - 0x0 -- Background 0xa2
      11'h511: dout  = 8'b11111110; // 1297 : 254 - 0xfe
      11'h512: dout  = 8'b00000000; // 1298 :   0 - 0x0
      11'h513: dout  = 8'b10000000; // 1299 : 128 - 0x80
      11'h514: dout  = 8'b10000000; // 1300 : 128 - 0x80
      11'h515: dout  = 8'b10000000; // 1301 : 128 - 0x80
      11'h516: dout  = 8'b10000000; // 1302 : 128 - 0x80
      11'h517: dout  = 8'b10000000; // 1303 : 128 - 0x80
      11'h518: dout  = 8'b10000000; // 1304 : 128 - 0x80 -- Background 0xa3
      11'h519: dout  = 8'b10000000; // 1305 : 128 - 0x80
      11'h51A: dout  = 8'b10000000; // 1306 : 128 - 0x80
      11'h51B: dout  = 8'b10000000; // 1307 : 128 - 0x80
      11'h51C: dout  = 8'b10000000; // 1308 : 128 - 0x80
      11'h51D: dout  = 8'b10000000; // 1309 : 128 - 0x80
      11'h51E: dout  = 8'b10000000; // 1310 : 128 - 0x80
      11'h51F: dout  = 8'b10000000; // 1311 : 128 - 0x80
      11'h520: dout  = 8'b00000000; // 1312 :   0 - 0x0 -- Background 0xa4
      11'h521: dout  = 8'b00110000; // 1313 :  48 - 0x30
      11'h522: dout  = 8'b00111000; // 1314 :  56 - 0x38
      11'h523: dout  = 8'b01111000; // 1315 : 120 - 0x78
      11'h524: dout  = 8'b01111100; // 1316 : 124 - 0x7c
      11'h525: dout  = 8'b01111101; // 1317 : 125 - 0x7d
      11'h526: dout  = 8'b00011101; // 1318 :  29 - 0x1d
      11'h527: dout  = 8'b00001101; // 1319 :  13 - 0xd
      11'h528: dout  = 8'b00001101; // 1320 :  13 - 0xd -- Background 0xa5
      11'h529: dout  = 8'b00011101; // 1321 :  29 - 0x1d
      11'h52A: dout  = 8'b00111101; // 1322 :  61 - 0x3d
      11'h52B: dout  = 8'b00111111; // 1323 :  63 - 0x3f
      11'h52C: dout  = 8'b00111111; // 1324 :  63 - 0x3f
      11'h52D: dout  = 8'b00011111; // 1325 :  31 - 0x1f
      11'h52E: dout  = 8'b00000001; // 1326 :   1 - 0x1
      11'h52F: dout  = 8'b00000000; // 1327 :   0 - 0x0
      11'h530: dout  = 8'b00000000; // 1328 :   0 - 0x0 -- Background 0xa6
      11'h531: dout  = 8'b00000000; // 1329 :   0 - 0x0
      11'h532: dout  = 8'b11100000; // 1330 : 224 - 0xe0
      11'h533: dout  = 8'b11111000; // 1331 : 248 - 0xf8
      11'h534: dout  = 8'b11111000; // 1332 : 248 - 0xf8
      11'h535: dout  = 8'b11110000; // 1333 : 240 - 0xf0
      11'h536: dout  = 8'b11000000; // 1334 : 192 - 0xc0
      11'h537: dout  = 8'b11000000; // 1335 : 192 - 0xc0
      11'h538: dout  = 8'b11000000; // 1336 : 192 - 0xc0 -- Background 0xa7
      11'h539: dout  = 8'b11110000; // 1337 : 240 - 0xf0
      11'h53A: dout  = 8'b11110000; // 1338 : 240 - 0xf0
      11'h53B: dout  = 8'b11000000; // 1339 : 192 - 0xc0
      11'h53C: dout  = 8'b11000000; // 1340 : 192 - 0xc0
      11'h53D: dout  = 8'b11000000; // 1341 : 192 - 0xc0
      11'h53E: dout  = 8'b11000000; // 1342 : 192 - 0xc0
      11'h53F: dout  = 8'b00000000; // 1343 :   0 - 0x0
      11'h540: dout  = 8'b00000000; // 1344 :   0 - 0x0 -- Background 0xa8
      11'h541: dout  = 8'b01100000; // 1345 :  96 - 0x60
      11'h542: dout  = 8'b01100000; // 1346 :  96 - 0x60
      11'h543: dout  = 8'b01100000; // 1347 :  96 - 0x60
      11'h544: dout  = 8'b01100000; // 1348 :  96 - 0x60
      11'h545: dout  = 8'b01100000; // 1349 :  96 - 0x60
      11'h546: dout  = 8'b01100000; // 1350 :  96 - 0x60
      11'h547: dout  = 8'b01100000; // 1351 :  96 - 0x60
      11'h548: dout  = 8'b01100000; // 1352 :  96 - 0x60 -- Background 0xa9
      11'h549: dout  = 8'b01100000; // 1353 :  96 - 0x60
      11'h54A: dout  = 8'b01100000; // 1354 :  96 - 0x60
      11'h54B: dout  = 8'b01100000; // 1355 :  96 - 0x60
      11'h54C: dout  = 8'b01100000; // 1356 :  96 - 0x60
      11'h54D: dout  = 8'b01100000; // 1357 :  96 - 0x60
      11'h54E: dout  = 8'b01100000; // 1358 :  96 - 0x60
      11'h54F: dout  = 8'b00000000; // 1359 :   0 - 0x0
      11'h550: dout  = 8'b00000000; // 1360 :   0 - 0x0 -- Background 0xaa
      11'h551: dout  = 8'b00000000; // 1361 :   0 - 0x0
      11'h552: dout  = 8'b00000000; // 1362 :   0 - 0x0
      11'h553: dout  = 8'b00000000; // 1363 :   0 - 0x0
      11'h554: dout  = 8'b00000000; // 1364 :   0 - 0x0
      11'h555: dout  = 8'b00000000; // 1365 :   0 - 0x0
      11'h556: dout  = 8'b00000000; // 1366 :   0 - 0x0
      11'h557: dout  = 8'b00000000; // 1367 :   0 - 0x0
      11'h558: dout  = 8'b00000000; // 1368 :   0 - 0x0 -- Background 0xab
      11'h559: dout  = 8'b00000000; // 1369 :   0 - 0x0
      11'h55A: dout  = 8'b00000000; // 1370 :   0 - 0x0
      11'h55B: dout  = 8'b00000000; // 1371 :   0 - 0x0
      11'h55C: dout  = 8'b00000000; // 1372 :   0 - 0x0
      11'h55D: dout  = 8'b00000000; // 1373 :   0 - 0x0
      11'h55E: dout  = 8'b00000000; // 1374 :   0 - 0x0
      11'h55F: dout  = 8'b00000000; // 1375 :   0 - 0x0
      11'h560: dout  = 8'b00000000; // 1376 :   0 - 0x0 -- Background 0xac
      11'h561: dout  = 8'b00000110; // 1377 :   6 - 0x6
      11'h562: dout  = 8'b00000110; // 1378 :   6 - 0x6
      11'h563: dout  = 8'b00000110; // 1379 :   6 - 0x6
      11'h564: dout  = 8'b00000110; // 1380 :   6 - 0x6
      11'h565: dout  = 8'b00000110; // 1381 :   6 - 0x6
      11'h566: dout  = 8'b00000110; // 1382 :   6 - 0x6
      11'h567: dout  = 8'b00000110; // 1383 :   6 - 0x6
      11'h568: dout  = 8'b00000110; // 1384 :   6 - 0x6 -- Background 0xad
      11'h569: dout  = 8'b00000110; // 1385 :   6 - 0x6
      11'h56A: dout  = 8'b00000110; // 1386 :   6 - 0x6
      11'h56B: dout  = 8'b00000110; // 1387 :   6 - 0x6
      11'h56C: dout  = 8'b00000110; // 1388 :   6 - 0x6
      11'h56D: dout  = 8'b00000110; // 1389 :   6 - 0x6
      11'h56E: dout  = 8'b00000110; // 1390 :   6 - 0x6
      11'h56F: dout  = 8'b00000000; // 1391 :   0 - 0x0
      11'h570: dout  = 8'b00000000; // 1392 :   0 - 0x0 -- Background 0xae
      11'h571: dout  = 8'b00000001; // 1393 :   1 - 0x1
      11'h572: dout  = 8'b00000011; // 1394 :   3 - 0x3
      11'h573: dout  = 8'b00000010; // 1395 :   2 - 0x2
      11'h574: dout  = 8'b00000010; // 1396 :   2 - 0x2
      11'h575: dout  = 8'b00000000; // 1397 :   0 - 0x0
      11'h576: dout  = 8'b00000011; // 1398 :   3 - 0x3
      11'h577: dout  = 8'b00000010; // 1399 :   2 - 0x2
      11'h578: dout  = 8'b00000001; // 1400 :   1 - 0x1 -- Background 0xaf
      11'h579: dout  = 8'b00000011; // 1401 :   3 - 0x3
      11'h57A: dout  = 8'b00000101; // 1402 :   5 - 0x5
      11'h57B: dout  = 8'b00000100; // 1403 :   4 - 0x4
      11'h57C: dout  = 8'b00000101; // 1404 :   5 - 0x5
      11'h57D: dout  = 8'b00001101; // 1405 :  13 - 0xd
      11'h57E: dout  = 8'b00001100; // 1406 :  12 - 0xc
      11'h57F: dout  = 8'b00000001; // 1407 :   1 - 0x1
      11'h580: dout  = 8'b00000000; // 1408 :   0 - 0x0 -- Background 0xb0
      11'h581: dout  = 8'b00000000; // 1409 :   0 - 0x0
      11'h582: dout  = 8'b01000000; // 1410 :  64 - 0x40
      11'h583: dout  = 8'b11110000; // 1411 : 240 - 0xf0
      11'h584: dout  = 8'b11101000; // 1412 : 232 - 0xe8
      11'h585: dout  = 8'b10010000; // 1413 : 144 - 0x90
      11'h586: dout  = 8'b01010000; // 1414 :  80 - 0x50
      11'h587: dout  = 8'b11010000; // 1415 : 208 - 0xd0
      11'h588: dout  = 8'b11111000; // 1416 : 248 - 0xf8 -- Background 0xb1
      11'h589: dout  = 8'b11000000; // 1417 : 192 - 0xc0
      11'h58A: dout  = 8'b11100000; // 1418 : 224 - 0xe0
      11'h58B: dout  = 8'b01000000; // 1419 :  64 - 0x40
      11'h58C: dout  = 8'b10000000; // 1420 : 128 - 0x80
      11'h58D: dout  = 8'b11000000; // 1421 : 192 - 0xc0
      11'h58E: dout  = 8'b11100000; // 1422 : 224 - 0xe0
      11'h58F: dout  = 8'b01110000; // 1423 : 112 - 0x70
      11'h590: dout  = 8'b00000001; // 1424 :   1 - 0x1 -- Background 0xb2
      11'h591: dout  = 8'b00001101; // 1425 :  13 - 0xd
      11'h592: dout  = 8'b00001101; // 1426 :  13 - 0xd
      11'h593: dout  = 8'b00000011; // 1427 :   3 - 0x3
      11'h594: dout  = 8'b00000011; // 1428 :   3 - 0x3
      11'h595: dout  = 8'b00000111; // 1429 :   7 - 0x7
      11'h596: dout  = 8'b00000111; // 1430 :   7 - 0x7
      11'h597: dout  = 8'b00000000; // 1431 :   0 - 0x0
      11'h598: dout  = 8'b00111111; // 1432 :  63 - 0x3f -- Background 0xb3
      11'h599: dout  = 8'b00111111; // 1433 :  63 - 0x3f
      11'h59A: dout  = 8'b00111111; // 1434 :  63 - 0x3f
      11'h59B: dout  = 8'b00111111; // 1435 :  63 - 0x3f
      11'h59C: dout  = 8'b00111111; // 1436 :  63 - 0x3f
      11'h59D: dout  = 8'b00111111; // 1437 :  63 - 0x3f
      11'h59E: dout  = 8'b00110101; // 1438 :  53 - 0x35
      11'h59F: dout  = 8'b00000000; // 1439 :   0 - 0x0
      11'h5A0: dout  = 8'b10110000; // 1440 : 176 - 0xb0 -- Background 0xb4
      11'h5A1: dout  = 8'b11000000; // 1441 : 192 - 0xc0
      11'h5A2: dout  = 8'b11100000; // 1442 : 224 - 0xe0
      11'h5A3: dout  = 8'b11100000; // 1443 : 224 - 0xe0
      11'h5A4: dout  = 8'b11110000; // 1444 : 240 - 0xf0
      11'h5A5: dout  = 8'b11110000; // 1445 : 240 - 0xf0
      11'h5A6: dout  = 8'b11110000; // 1446 : 240 - 0xf0
      11'h5A7: dout  = 8'b00000000; // 1447 :   0 - 0x0
      11'h5A8: dout  = 8'b11111100; // 1448 : 252 - 0xfc -- Background 0xb5
      11'h5A9: dout  = 8'b11111000; // 1449 : 248 - 0xf8
      11'h5AA: dout  = 8'b11111100; // 1450 : 252 - 0xfc
      11'h5AB: dout  = 8'b11111000; // 1451 : 248 - 0xf8
      11'h5AC: dout  = 8'b11111100; // 1452 : 252 - 0xfc
      11'h5AD: dout  = 8'b11111000; // 1453 : 248 - 0xf8
      11'h5AE: dout  = 8'b01010100; // 1454 :  84 - 0x54
      11'h5AF: dout  = 8'b00000000; // 1455 :   0 - 0x0
      11'h5B0: dout  = 8'b00000000; // 1456 :   0 - 0x0 -- Background 0xb6
      11'h5B1: dout  = 8'b01111111; // 1457 : 127 - 0x7f
      11'h5B2: dout  = 8'b01111111; // 1458 : 127 - 0x7f
      11'h5B3: dout  = 8'b01111111; // 1459 : 127 - 0x7f
      11'h5B4: dout  = 8'b01111111; // 1460 : 127 - 0x7f
      11'h5B5: dout  = 8'b01111111; // 1461 : 127 - 0x7f
      11'h5B6: dout  = 8'b01101010; // 1462 : 106 - 0x6a
      11'h5B7: dout  = 8'b00000000; // 1463 :   0 - 0x0
      11'h5B8: dout  = 8'b00000000; // 1464 :   0 - 0x0 -- Background 0xb7
      11'h5B9: dout  = 8'b01111011; // 1465 : 123 - 0x7b
      11'h5BA: dout  = 8'b01110011; // 1466 : 115 - 0x73
      11'h5BB: dout  = 8'b01111011; // 1467 : 123 - 0x7b
      11'h5BC: dout  = 8'b01110011; // 1468 : 115 - 0x73
      11'h5BD: dout  = 8'b01111011; // 1469 : 123 - 0x7b
      11'h5BE: dout  = 8'b01010011; // 1470 :  83 - 0x53
      11'h5BF: dout  = 8'b00000000; // 1471 :   0 - 0x0
      11'h5C0: dout  = 8'b00000000; // 1472 :   0 - 0x0 -- Background 0xb8
      11'h5C1: dout  = 8'b11011110; // 1473 : 222 - 0xde
      11'h5C2: dout  = 8'b10011110; // 1474 : 158 - 0x9e
      11'h5C3: dout  = 8'b11011100; // 1475 : 220 - 0xdc
      11'h5C4: dout  = 8'b10011110; // 1476 : 158 - 0x9e
      11'h5C5: dout  = 8'b11011100; // 1477 : 220 - 0xdc
      11'h5C6: dout  = 8'b10011010; // 1478 : 154 - 0x9a
      11'h5C7: dout  = 8'b00000000; // 1479 :   0 - 0x0
      11'h5C8: dout  = 8'b00000000; // 1480 :   0 - 0x0 -- Background 0xb9
      11'h5C9: dout  = 8'b11111110; // 1481 : 254 - 0xfe
      11'h5CA: dout  = 8'b11111100; // 1482 : 252 - 0xfc
      11'h5CB: dout  = 8'b11111110; // 1483 : 254 - 0xfe
      11'h5CC: dout  = 8'b11111100; // 1484 : 252 - 0xfc
      11'h5CD: dout  = 8'b11111110; // 1485 : 254 - 0xfe
      11'h5CE: dout  = 8'b01010100; // 1486 :  84 - 0x54
      11'h5CF: dout  = 8'b00000000; // 1487 :   0 - 0x0
      11'h5D0: dout  = 8'b00000000; // 1488 :   0 - 0x0 -- Background 0xba
      11'h5D1: dout  = 8'b01111111; // 1489 : 127 - 0x7f
      11'h5D2: dout  = 8'b01111111; // 1490 : 127 - 0x7f
      11'h5D3: dout  = 8'b00000000; // 1491 :   0 - 0x0
      11'h5D4: dout  = 8'b01111111; // 1492 : 127 - 0x7f
      11'h5D5: dout  = 8'b01111111; // 1493 : 127 - 0x7f
      11'h5D6: dout  = 8'b01101010; // 1494 : 106 - 0x6a
      11'h5D7: dout  = 8'b00000000; // 1495 :   0 - 0x0
      11'h5D8: dout  = 8'b00000000; // 1496 :   0 - 0x0 -- Background 0xbb
      11'h5D9: dout  = 8'b00000000; // 1497 :   0 - 0x0
      11'h5DA: dout  = 8'b00000000; // 1498 :   0 - 0x0
      11'h5DB: dout  = 8'b00000000; // 1499 :   0 - 0x0
      11'h5DC: dout  = 8'b00000000; // 1500 :   0 - 0x0
      11'h5DD: dout  = 8'b00000000; // 1501 :   0 - 0x0
      11'h5DE: dout  = 8'b00000000; // 1502 :   0 - 0x0
      11'h5DF: dout  = 8'b00000000; // 1503 :   0 - 0x0
      11'h5E0: dout  = 8'b00000000; // 1504 :   0 - 0x0 -- Background 0xbc
      11'h5E1: dout  = 8'b11111110; // 1505 : 254 - 0xfe
      11'h5E2: dout  = 8'b11111110; // 1506 : 254 - 0xfe
      11'h5E3: dout  = 8'b00000000; // 1507 :   0 - 0x0
      11'h5E4: dout  = 8'b10011110; // 1508 : 158 - 0x9e
      11'h5E5: dout  = 8'b11011100; // 1509 : 220 - 0xdc
      11'h5E6: dout  = 8'b10011010; // 1510 : 154 - 0x9a
      11'h5E7: dout  = 8'b00000000; // 1511 :   0 - 0x0
      11'h5E8: dout  = 8'b00000000; // 1512 :   0 - 0x0 -- Background 0xbd
      11'h5E9: dout  = 8'b00000000; // 1513 :   0 - 0x0
      11'h5EA: dout  = 8'b00000000; // 1514 :   0 - 0x0
      11'h5EB: dout  = 8'b00000000; // 1515 :   0 - 0x0
      11'h5EC: dout  = 8'b00000000; // 1516 :   0 - 0x0
      11'h5ED: dout  = 8'b00000000; // 1517 :   0 - 0x0
      11'h5EE: dout  = 8'b00000000; // 1518 :   0 - 0x0
      11'h5EF: dout  = 8'b00000000; // 1519 :   0 - 0x0
      11'h5F0: dout  = 8'b00000000; // 1520 :   0 - 0x0 -- Background 0xbe
      11'h5F1: dout  = 8'b00000000; // 1521 :   0 - 0x0
      11'h5F2: dout  = 8'b00000000; // 1522 :   0 - 0x0
      11'h5F3: dout  = 8'b00000000; // 1523 :   0 - 0x0
      11'h5F4: dout  = 8'b00000000; // 1524 :   0 - 0x0
      11'h5F5: dout  = 8'b00000000; // 1525 :   0 - 0x0
      11'h5F6: dout  = 8'b00000000; // 1526 :   0 - 0x0
      11'h5F7: dout  = 8'b00000000; // 1527 :   0 - 0x0
      11'h5F8: dout  = 8'b00000000; // 1528 :   0 - 0x0 -- Background 0xbf
      11'h5F9: dout  = 8'b00000000; // 1529 :   0 - 0x0
      11'h5FA: dout  = 8'b00000000; // 1530 :   0 - 0x0
      11'h5FB: dout  = 8'b00000000; // 1531 :   0 - 0x0
      11'h5FC: dout  = 8'b00000000; // 1532 :   0 - 0x0
      11'h5FD: dout  = 8'b00000000; // 1533 :   0 - 0x0
      11'h5FE: dout  = 8'b00000000; // 1534 :   0 - 0x0
      11'h5FF: dout  = 8'b00000000; // 1535 :   0 - 0x0
      11'h600: dout  = 8'b00000000; // 1536 :   0 - 0x0 -- Background 0xc0
      11'h601: dout  = 8'b00000000; // 1537 :   0 - 0x0
      11'h602: dout  = 8'b00000000; // 1538 :   0 - 0x0
      11'h603: dout  = 8'b00000000; // 1539 :   0 - 0x0
      11'h604: dout  = 8'b00000000; // 1540 :   0 - 0x0
      11'h605: dout  = 8'b00000000; // 1541 :   0 - 0x0
      11'h606: dout  = 8'b00000000; // 1542 :   0 - 0x0
      11'h607: dout  = 8'b00000000; // 1543 :   0 - 0x0
      11'h608: dout  = 8'b00000000; // 1544 :   0 - 0x0 -- Background 0xc1
      11'h609: dout  = 8'b00000000; // 1545 :   0 - 0x0
      11'h60A: dout  = 8'b00000000; // 1546 :   0 - 0x0
      11'h60B: dout  = 8'b00000000; // 1547 :   0 - 0x0
      11'h60C: dout  = 8'b00000000; // 1548 :   0 - 0x0
      11'h60D: dout  = 8'b00000000; // 1549 :   0 - 0x0
      11'h60E: dout  = 8'b00000000; // 1550 :   0 - 0x0
      11'h60F: dout  = 8'b00000000; // 1551 :   0 - 0x0
      11'h610: dout  = 8'b00000000; // 1552 :   0 - 0x0 -- Background 0xc2
      11'h611: dout  = 8'b00000000; // 1553 :   0 - 0x0
      11'h612: dout  = 8'b00000000; // 1554 :   0 - 0x0
      11'h613: dout  = 8'b00000000; // 1555 :   0 - 0x0
      11'h614: dout  = 8'b00000000; // 1556 :   0 - 0x0
      11'h615: dout  = 8'b00000000; // 1557 :   0 - 0x0
      11'h616: dout  = 8'b00000000; // 1558 :   0 - 0x0
      11'h617: dout  = 8'b00000000; // 1559 :   0 - 0x0
      11'h618: dout  = 8'b00000000; // 1560 :   0 - 0x0 -- Background 0xc3
      11'h619: dout  = 8'b00000000; // 1561 :   0 - 0x0
      11'h61A: dout  = 8'b00000000; // 1562 :   0 - 0x0
      11'h61B: dout  = 8'b00000000; // 1563 :   0 - 0x0
      11'h61C: dout  = 8'b00000000; // 1564 :   0 - 0x0
      11'h61D: dout  = 8'b00000000; // 1565 :   0 - 0x0
      11'h61E: dout  = 8'b00000000; // 1566 :   0 - 0x0
      11'h61F: dout  = 8'b00000000; // 1567 :   0 - 0x0
      11'h620: dout  = 8'b00000000; // 1568 :   0 - 0x0 -- Background 0xc4
      11'h621: dout  = 8'b00000000; // 1569 :   0 - 0x0
      11'h622: dout  = 8'b00000000; // 1570 :   0 - 0x0
      11'h623: dout  = 8'b00000000; // 1571 :   0 - 0x0
      11'h624: dout  = 8'b00000000; // 1572 :   0 - 0x0
      11'h625: dout  = 8'b00000000; // 1573 :   0 - 0x0
      11'h626: dout  = 8'b00000000; // 1574 :   0 - 0x0
      11'h627: dout  = 8'b00000000; // 1575 :   0 - 0x0
      11'h628: dout  = 8'b00000000; // 1576 :   0 - 0x0 -- Background 0xc5
      11'h629: dout  = 8'b00000000; // 1577 :   0 - 0x0
      11'h62A: dout  = 8'b00000000; // 1578 :   0 - 0x0
      11'h62B: dout  = 8'b00000001; // 1579 :   1 - 0x1
      11'h62C: dout  = 8'b00000111; // 1580 :   7 - 0x7
      11'h62D: dout  = 8'b00001111; // 1581 :  15 - 0xf
      11'h62E: dout  = 8'b00001111; // 1582 :  15 - 0xf
      11'h62F: dout  = 8'b00011111; // 1583 :  31 - 0x1f
      11'h630: dout  = 8'b00000000; // 1584 :   0 - 0x0 -- Background 0xc6
      11'h631: dout  = 8'b00011111; // 1585 :  31 - 0x1f
      11'h632: dout  = 8'b01111111; // 1586 : 127 - 0x7f
      11'h633: dout  = 8'b11111111; // 1587 : 255 - 0xff
      11'h634: dout  = 8'b11111111; // 1588 : 255 - 0xff
      11'h635: dout  = 8'b11111111; // 1589 : 255 - 0xff
      11'h636: dout  = 8'b11111111; // 1590 : 255 - 0xff
      11'h637: dout  = 8'b11111111; // 1591 : 255 - 0xff
      11'h638: dout  = 8'b00011111; // 1592 :  31 - 0x1f -- Background 0xc7
      11'h639: dout  = 8'b00111111; // 1593 :  63 - 0x3f
      11'h63A: dout  = 8'b00111111; // 1594 :  63 - 0x3f
      11'h63B: dout  = 8'b01111111; // 1595 : 127 - 0x7f
      11'h63C: dout  = 8'b01111111; // 1596 : 127 - 0x7f
      11'h63D: dout  = 8'b01111111; // 1597 : 127 - 0x7f
      11'h63E: dout  = 8'b01111111; // 1598 : 127 - 0x7f
      11'h63F: dout  = 8'b01111111; // 1599 : 127 - 0x7f
      11'h640: dout  = 8'b00000000; // 1600 :   0 - 0x0 -- Background 0xc8
      11'h641: dout  = 8'b11111111; // 1601 : 255 - 0xff
      11'h642: dout  = 8'b11111111; // 1602 : 255 - 0xff
      11'h643: dout  = 8'b11111111; // 1603 : 255 - 0xff
      11'h644: dout  = 8'b11111111; // 1604 : 255 - 0xff
      11'h645: dout  = 8'b11111111; // 1605 : 255 - 0xff
      11'h646: dout  = 8'b11111111; // 1606 : 255 - 0xff
      11'h647: dout  = 8'b11111111; // 1607 : 255 - 0xff
      11'h648: dout  = 8'b11101000; // 1608 : 232 - 0xe8 -- Background 0xc9
      11'h649: dout  = 8'b11010100; // 1609 : 212 - 0xd4
      11'h64A: dout  = 8'b11101000; // 1610 : 232 - 0xe8
      11'h64B: dout  = 8'b11010100; // 1611 : 212 - 0xd4
      11'h64C: dout  = 8'b11101010; // 1612 : 234 - 0xea
      11'h64D: dout  = 8'b11010100; // 1613 : 212 - 0xd4
      11'h64E: dout  = 8'b11101010; // 1614 : 234 - 0xea
      11'h64F: dout  = 8'b11010100; // 1615 : 212 - 0xd4
      11'h650: dout  = 8'b00000000; // 1616 :   0 - 0x0 -- Background 0xca
      11'h651: dout  = 8'b00000000; // 1617 :   0 - 0x0
      11'h652: dout  = 8'b00000000; // 1618 :   0 - 0x0
      11'h653: dout  = 8'b00000000; // 1619 :   0 - 0x0
      11'h654: dout  = 8'b00000000; // 1620 :   0 - 0x0
      11'h655: dout  = 8'b00000000; // 1621 :   0 - 0x0
      11'h656: dout  = 8'b00000000; // 1622 :   0 - 0x0
      11'h657: dout  = 8'b00000000; // 1623 :   0 - 0x0
      11'h658: dout  = 8'b00000000; // 1624 :   0 - 0x0 -- Background 0xcb
      11'h659: dout  = 8'b00000000; // 1625 :   0 - 0x0
      11'h65A: dout  = 8'b00000000; // 1626 :   0 - 0x0
      11'h65B: dout  = 8'b00000000; // 1627 :   0 - 0x0
      11'h65C: dout  = 8'b00000000; // 1628 :   0 - 0x0
      11'h65D: dout  = 8'b00000000; // 1629 :   0 - 0x0
      11'h65E: dout  = 8'b00000000; // 1630 :   0 - 0x0
      11'h65F: dout  = 8'b00000000; // 1631 :   0 - 0x0
      11'h660: dout  = 8'b00000000; // 1632 :   0 - 0x0 -- Background 0xcc
      11'h661: dout  = 8'b00000000; // 1633 :   0 - 0x0
      11'h662: dout  = 8'b00000000; // 1634 :   0 - 0x0
      11'h663: dout  = 8'b00000000; // 1635 :   0 - 0x0
      11'h664: dout  = 8'b00000101; // 1636 :   5 - 0x5
      11'h665: dout  = 8'b00000010; // 1637 :   2 - 0x2
      11'h666: dout  = 8'b00000001; // 1638 :   1 - 0x1
      11'h667: dout  = 8'b00000000; // 1639 :   0 - 0x0
      11'h668: dout  = 8'b00000000; // 1640 :   0 - 0x0 -- Background 0xcd
      11'h669: dout  = 8'b00000000; // 1641 :   0 - 0x0
      11'h66A: dout  = 8'b00000000; // 1642 :   0 - 0x0
      11'h66B: dout  = 8'b10000000; // 1643 : 128 - 0x80
      11'h66C: dout  = 8'b01010000; // 1644 :  80 - 0x50
      11'h66D: dout  = 8'b10100000; // 1645 : 160 - 0xa0
      11'h66E: dout  = 8'b01000000; // 1646 :  64 - 0x40
      11'h66F: dout  = 8'b10000000; // 1647 : 128 - 0x80
      11'h670: dout  = 8'b00000000; // 1648 :   0 - 0x0 -- Background 0xce
      11'h671: dout  = 8'b00000000; // 1649 :   0 - 0x0
      11'h672: dout  = 8'b00000000; // 1650 :   0 - 0x0
      11'h673: dout  = 8'b00000000; // 1651 :   0 - 0x0
      11'h674: dout  = 8'b00110000; // 1652 :  48 - 0x30
      11'h675: dout  = 8'b01111111; // 1653 : 127 - 0x7f
      11'h676: dout  = 8'b00110000; // 1654 :  48 - 0x30
      11'h677: dout  = 8'b00110000; // 1655 :  48 - 0x30
      11'h678: dout  = 8'b00000000; // 1656 :   0 - 0x0 -- Background 0xcf
      11'h679: dout  = 8'b00000000; // 1657 :   0 - 0x0
      11'h67A: dout  = 8'b00000000; // 1658 :   0 - 0x0
      11'h67B: dout  = 8'b00000000; // 1659 :   0 - 0x0
      11'h67C: dout  = 8'b00001100; // 1660 :  12 - 0xc
      11'h67D: dout  = 8'b11111110; // 1661 : 254 - 0xfe
      11'h67E: dout  = 8'b00001100; // 1662 :  12 - 0xc
      11'h67F: dout  = 8'b00001100; // 1663 :  12 - 0xc
      11'h680: dout  = 8'b00000000; // 1664 :   0 - 0x0 -- Background 0xd0
      11'h681: dout  = 8'b00000000; // 1665 :   0 - 0x0
      11'h682: dout  = 8'b00000000; // 1666 :   0 - 0x0
      11'h683: dout  = 8'b00000000; // 1667 :   0 - 0x0
      11'h684: dout  = 8'b00000000; // 1668 :   0 - 0x0
      11'h685: dout  = 8'b00000000; // 1669 :   0 - 0x0
      11'h686: dout  = 8'b00000000; // 1670 :   0 - 0x0
      11'h687: dout  = 8'b00000000; // 1671 :   0 - 0x0
      11'h688: dout  = 8'b00000000; // 1672 :   0 - 0x0 -- Background 0xd1
      11'h689: dout  = 8'b00000000; // 1673 :   0 - 0x0
      11'h68A: dout  = 8'b00000000; // 1674 :   0 - 0x0
      11'h68B: dout  = 8'b00000000; // 1675 :   0 - 0x0
      11'h68C: dout  = 8'b00000000; // 1676 :   0 - 0x0
      11'h68D: dout  = 8'b00000000; // 1677 :   0 - 0x0
      11'h68E: dout  = 8'b00000000; // 1678 :   0 - 0x0
      11'h68F: dout  = 8'b00000000; // 1679 :   0 - 0x0
      11'h690: dout  = 8'b00000111; // 1680 :   7 - 0x7 -- Background 0xd2
      11'h691: dout  = 8'b00000111; // 1681 :   7 - 0x7
      11'h692: dout  = 8'b00000111; // 1682 :   7 - 0x7
      11'h693: dout  = 8'b00000111; // 1683 :   7 - 0x7
      11'h694: dout  = 8'b00000111; // 1684 :   7 - 0x7
      11'h695: dout  = 8'b00000111; // 1685 :   7 - 0x7
      11'h696: dout  = 8'b00000111; // 1686 :   7 - 0x7
      11'h697: dout  = 8'b00000111; // 1687 :   7 - 0x7
      11'h698: dout  = 8'b11100000; // 1688 : 224 - 0xe0 -- Background 0xd3
      11'h699: dout  = 8'b11100000; // 1689 : 224 - 0xe0
      11'h69A: dout  = 8'b11000000; // 1690 : 192 - 0xc0
      11'h69B: dout  = 8'b11100000; // 1691 : 224 - 0xe0
      11'h69C: dout  = 8'b10100000; // 1692 : 160 - 0xa0
      11'h69D: dout  = 8'b11100000; // 1693 : 224 - 0xe0
      11'h69E: dout  = 8'b11000000; // 1694 : 192 - 0xc0
      11'h69F: dout  = 8'b11100000; // 1695 : 224 - 0xe0
      11'h6A0: dout  = 8'b00000000; // 1696 :   0 - 0x0 -- Background 0xd4
      11'h6A1: dout  = 8'b00000000; // 1697 :   0 - 0x0
      11'h6A2: dout  = 8'b00000000; // 1698 :   0 - 0x0
      11'h6A3: dout  = 8'b00000000; // 1699 :   0 - 0x0
      11'h6A4: dout  = 8'b00000000; // 1700 :   0 - 0x0
      11'h6A5: dout  = 8'b00000000; // 1701 :   0 - 0x0
      11'h6A6: dout  = 8'b00000000; // 1702 :   0 - 0x0
      11'h6A7: dout  = 8'b00000000; // 1703 :   0 - 0x0
      11'h6A8: dout  = 8'b00000000; // 1704 :   0 - 0x0 -- Background 0xd5
      11'h6A9: dout  = 8'b11111000; // 1705 : 248 - 0xf8
      11'h6AA: dout  = 8'b11111110; // 1706 : 254 - 0xfe
      11'h6AB: dout  = 8'b11111111; // 1707 : 255 - 0xff
      11'h6AC: dout  = 8'b11111111; // 1708 : 255 - 0xff
      11'h6AD: dout  = 8'b11111111; // 1709 : 255 - 0xff
      11'h6AE: dout  = 8'b11111111; // 1710 : 255 - 0xff
      11'h6AF: dout  = 8'b11111111; // 1711 : 255 - 0xff
      11'h6B0: dout  = 8'b00000000; // 1712 :   0 - 0x0 -- Background 0xd6
      11'h6B1: dout  = 8'b00000000; // 1713 :   0 - 0x0
      11'h6B2: dout  = 8'b00000000; // 1714 :   0 - 0x0
      11'h6B3: dout  = 8'b10000000; // 1715 : 128 - 0x80
      11'h6B4: dout  = 8'b10100000; // 1716 : 160 - 0xa0
      11'h6B5: dout  = 8'b01010000; // 1717 :  80 - 0x50
      11'h6B6: dout  = 8'b10100000; // 1718 : 160 - 0xa0
      11'h6B7: dout  = 8'b11010000; // 1719 : 208 - 0xd0
      11'h6B8: dout  = 8'b01111111; // 1720 : 127 - 0x7f -- Background 0xd7
      11'h6B9: dout  = 8'b01111111; // 1721 : 127 - 0x7f
      11'h6BA: dout  = 8'b01111111; // 1722 : 127 - 0x7f
      11'h6BB: dout  = 8'b00111111; // 1723 :  63 - 0x3f
      11'h6BC: dout  = 8'b00111111; // 1724 :  63 - 0x3f
      11'h6BD: dout  = 8'b00001111; // 1725 :  15 - 0xf
      11'h6BE: dout  = 8'b00000111; // 1726 :   7 - 0x7
      11'h6BF: dout  = 8'b00000000; // 1727 :   0 - 0x0
      11'h6C0: dout  = 8'b11111111; // 1728 : 255 - 0xff -- Background 0xd8
      11'h6C1: dout  = 8'b11111111; // 1729 : 255 - 0xff
      11'h6C2: dout  = 8'b11111111; // 1730 : 255 - 0xff
      11'h6C3: dout  = 8'b11111111; // 1731 : 255 - 0xff
      11'h6C4: dout  = 8'b11111111; // 1732 : 255 - 0xff
      11'h6C5: dout  = 8'b11111111; // 1733 : 255 - 0xff
      11'h6C6: dout  = 8'b11111111; // 1734 : 255 - 0xff
      11'h6C7: dout  = 8'b00000000; // 1735 :   0 - 0x0
      11'h6C8: dout  = 8'b11101010; // 1736 : 234 - 0xea -- Background 0xd9
      11'h6C9: dout  = 8'b11010100; // 1737 : 212 - 0xd4
      11'h6CA: dout  = 8'b11101010; // 1738 : 234 - 0xea
      11'h6CB: dout  = 8'b11010100; // 1739 : 212 - 0xd4
      11'h6CC: dout  = 8'b10101000; // 1740 : 168 - 0xa8
      11'h6CD: dout  = 8'b01010000; // 1741 :  80 - 0x50
      11'h6CE: dout  = 8'b10100000; // 1742 : 160 - 0xa0
      11'h6CF: dout  = 8'b00000000; // 1743 :   0 - 0x0
      11'h6D0: dout  = 8'b00000000; // 1744 :   0 - 0x0 -- Background 0xda
      11'h6D1: dout  = 8'b00000000; // 1745 :   0 - 0x0
      11'h6D2: dout  = 8'b00001100; // 1746 :  12 - 0xc
      11'h6D3: dout  = 8'b00000000; // 1747 :   0 - 0x0
      11'h6D4: dout  = 8'b00000000; // 1748 :   0 - 0x0
      11'h6D5: dout  = 8'b00000000; // 1749 :   0 - 0x0
      11'h6D6: dout  = 8'b00000000; // 1750 :   0 - 0x0
      11'h6D7: dout  = 8'b00000000; // 1751 :   0 - 0x0
      11'h6D8: dout  = 8'b00000000; // 1752 :   0 - 0x0 -- Background 0xdb
      11'h6D9: dout  = 8'b10000000; // 1753 : 128 - 0x80
      11'h6DA: dout  = 8'b10000000; // 1754 : 128 - 0x80
      11'h6DB: dout  = 8'b10000000; // 1755 : 128 - 0x80
      11'h6DC: dout  = 8'b10011000; // 1756 : 152 - 0x98
      11'h6DD: dout  = 8'b10000000; // 1757 : 128 - 0x80
      11'h6DE: dout  = 8'b10000000; // 1758 : 128 - 0x80
      11'h6DF: dout  = 8'b10000000; // 1759 : 128 - 0x80
      11'h6E0: dout  = 8'b00000000; // 1760 :   0 - 0x0 -- Background 0xdc
      11'h6E1: dout  = 8'b00000000; // 1761 :   0 - 0x0
      11'h6E2: dout  = 8'b00000000; // 1762 :   0 - 0x0
      11'h6E3: dout  = 8'b00000000; // 1763 :   0 - 0x0
      11'h6E4: dout  = 8'b00000010; // 1764 :   2 - 0x2
      11'h6E5: dout  = 8'b00000011; // 1765 :   3 - 0x3
      11'h6E6: dout  = 8'b00000011; // 1766 :   3 - 0x3
      11'h6E7: dout  = 8'b00000001; // 1767 :   1 - 0x1
      11'h6E8: dout  = 8'b00000000; // 1768 :   0 - 0x0 -- Background 0xdd
      11'h6E9: dout  = 8'b00000000; // 1769 :   0 - 0x0
      11'h6EA: dout  = 8'b00000000; // 1770 :   0 - 0x0
      11'h6EB: dout  = 8'b00000000; // 1771 :   0 - 0x0
      11'h6EC: dout  = 8'b10100000; // 1772 : 160 - 0xa0
      11'h6ED: dout  = 8'b11100000; // 1773 : 224 - 0xe0
      11'h6EE: dout  = 8'b11100000; // 1774 : 224 - 0xe0
      11'h6EF: dout  = 8'b11000000; // 1775 : 192 - 0xc0
      11'h6F0: dout  = 8'b00110000; // 1776 :  48 - 0x30 -- Background 0xde
      11'h6F1: dout  = 8'b01111111; // 1777 : 127 - 0x7f
      11'h6F2: dout  = 8'b00110000; // 1778 :  48 - 0x30
      11'h6F3: dout  = 8'b00110000; // 1779 :  48 - 0x30
      11'h6F4: dout  = 8'b00110000; // 1780 :  48 - 0x30
      11'h6F5: dout  = 8'b00110000; // 1781 :  48 - 0x30
      11'h6F6: dout  = 8'b00110000; // 1782 :  48 - 0x30
      11'h6F7: dout  = 8'b00110000; // 1783 :  48 - 0x30
      11'h6F8: dout  = 8'b00001100; // 1784 :  12 - 0xc -- Background 0xdf
      11'h6F9: dout  = 8'b11111110; // 1785 : 254 - 0xfe
      11'h6FA: dout  = 8'b00001100; // 1786 :  12 - 0xc
      11'h6FB: dout  = 8'b00001100; // 1787 :  12 - 0xc
      11'h6FC: dout  = 8'b00001100; // 1788 :  12 - 0xc
      11'h6FD: dout  = 8'b00001100; // 1789 :  12 - 0xc
      11'h6FE: dout  = 8'b00001100; // 1790 :  12 - 0xc
      11'h6FF: dout  = 8'b00001100; // 1791 :  12 - 0xc
      11'h700: dout  = 8'b00000000; // 1792 :   0 - 0x0 -- Background 0xe0
      11'h701: dout  = 8'b00000000; // 1793 :   0 - 0x0
      11'h702: dout  = 8'b00000000; // 1794 :   0 - 0x0
      11'h703: dout  = 8'b00000000; // 1795 :   0 - 0x0
      11'h704: dout  = 8'b00000000; // 1796 :   0 - 0x0
      11'h705: dout  = 8'b00000000; // 1797 :   0 - 0x0
      11'h706: dout  = 8'b00000000; // 1798 :   0 - 0x0
      11'h707: dout  = 8'b00000000; // 1799 :   0 - 0x0
      11'h708: dout  = 8'b00000000; // 1800 :   0 - 0x0 -- Background 0xe1
      11'h709: dout  = 8'b00000000; // 1801 :   0 - 0x0
      11'h70A: dout  = 8'b00000000; // 1802 :   0 - 0x0
      11'h70B: dout  = 8'b00000000; // 1803 :   0 - 0x0
      11'h70C: dout  = 8'b00000000; // 1804 :   0 - 0x0
      11'h70D: dout  = 8'b00000000; // 1805 :   0 - 0x0
      11'h70E: dout  = 8'b00000000; // 1806 :   0 - 0x0
      11'h70F: dout  = 8'b00000000; // 1807 :   0 - 0x0
      11'h710: dout  = 8'b00000000; // 1808 :   0 - 0x0 -- Background 0xe2
      11'h711: dout  = 8'b00000000; // 1809 :   0 - 0x0
      11'h712: dout  = 8'b00000000; // 1810 :   0 - 0x0
      11'h713: dout  = 8'b00000000; // 1811 :   0 - 0x0
      11'h714: dout  = 8'b00000000; // 1812 :   0 - 0x0
      11'h715: dout  = 8'b00000000; // 1813 :   0 - 0x0
      11'h716: dout  = 8'b00000000; // 1814 :   0 - 0x0
      11'h717: dout  = 8'b00000000; // 1815 :   0 - 0x0
      11'h718: dout  = 8'b00000000; // 1816 :   0 - 0x0 -- Background 0xe3
      11'h719: dout  = 8'b00000000; // 1817 :   0 - 0x0
      11'h71A: dout  = 8'b00000000; // 1818 :   0 - 0x0
      11'h71B: dout  = 8'b00000000; // 1819 :   0 - 0x0
      11'h71C: dout  = 8'b00000000; // 1820 :   0 - 0x0
      11'h71D: dout  = 8'b00000000; // 1821 :   0 - 0x0
      11'h71E: dout  = 8'b00000000; // 1822 :   0 - 0x0
      11'h71F: dout  = 8'b00000000; // 1823 :   0 - 0x0
      11'h720: dout  = 8'b00000000; // 1824 :   0 - 0x0 -- Background 0xe4
      11'h721: dout  = 8'b00000000; // 1825 :   0 - 0x0
      11'h722: dout  = 8'b00000000; // 1826 :   0 - 0x0
      11'h723: dout  = 8'b00000000; // 1827 :   0 - 0x0
      11'h724: dout  = 8'b00000000; // 1828 :   0 - 0x0
      11'h725: dout  = 8'b00000000; // 1829 :   0 - 0x0
      11'h726: dout  = 8'b00000000; // 1830 :   0 - 0x0
      11'h727: dout  = 8'b00000000; // 1831 :   0 - 0x0
      11'h728: dout  = 8'b00000000; // 1832 :   0 - 0x0 -- Background 0xe5
      11'h729: dout  = 8'b00000000; // 1833 :   0 - 0x0
      11'h72A: dout  = 8'b00000000; // 1834 :   0 - 0x0
      11'h72B: dout  = 8'b00000000; // 1835 :   0 - 0x0
      11'h72C: dout  = 8'b00000000; // 1836 :   0 - 0x0
      11'h72D: dout  = 8'b00000000; // 1837 :   0 - 0x0
      11'h72E: dout  = 8'b00000000; // 1838 :   0 - 0x0
      11'h72F: dout  = 8'b00000000; // 1839 :   0 - 0x0
      11'h730: dout  = 8'b00000000; // 1840 :   0 - 0x0 -- Background 0xe6
      11'h731: dout  = 8'b00000000; // 1841 :   0 - 0x0
      11'h732: dout  = 8'b00000000; // 1842 :   0 - 0x0
      11'h733: dout  = 8'b00000000; // 1843 :   0 - 0x0
      11'h734: dout  = 8'b00000000; // 1844 :   0 - 0x0
      11'h735: dout  = 8'b00000000; // 1845 :   0 - 0x0
      11'h736: dout  = 8'b00000000; // 1846 :   0 - 0x0
      11'h737: dout  = 8'b00000000; // 1847 :   0 - 0x0
      11'h738: dout  = 8'b00000000; // 1848 :   0 - 0x0 -- Background 0xe7
      11'h739: dout  = 8'b00000000; // 1849 :   0 - 0x0
      11'h73A: dout  = 8'b00000000; // 1850 :   0 - 0x0
      11'h73B: dout  = 8'b00000000; // 1851 :   0 - 0x0
      11'h73C: dout  = 8'b00000000; // 1852 :   0 - 0x0
      11'h73D: dout  = 8'b00000000; // 1853 :   0 - 0x0
      11'h73E: dout  = 8'b00000000; // 1854 :   0 - 0x0
      11'h73F: dout  = 8'b00000000; // 1855 :   0 - 0x0
      11'h740: dout  = 8'b00000000; // 1856 :   0 - 0x0 -- Background 0xe8
      11'h741: dout  = 8'b00000000; // 1857 :   0 - 0x0
      11'h742: dout  = 8'b00000000; // 1858 :   0 - 0x0
      11'h743: dout  = 8'b00000000; // 1859 :   0 - 0x0
      11'h744: dout  = 8'b00000000; // 1860 :   0 - 0x0
      11'h745: dout  = 8'b00000000; // 1861 :   0 - 0x0
      11'h746: dout  = 8'b00000000; // 1862 :   0 - 0x0
      11'h747: dout  = 8'b00000000; // 1863 :   0 - 0x0
      11'h748: dout  = 8'b00000000; // 1864 :   0 - 0x0 -- Background 0xe9
      11'h749: dout  = 8'b00000000; // 1865 :   0 - 0x0
      11'h74A: dout  = 8'b00000000; // 1866 :   0 - 0x0
      11'h74B: dout  = 8'b00000000; // 1867 :   0 - 0x0
      11'h74C: dout  = 8'b00000000; // 1868 :   0 - 0x0
      11'h74D: dout  = 8'b00000000; // 1869 :   0 - 0x0
      11'h74E: dout  = 8'b00000000; // 1870 :   0 - 0x0
      11'h74F: dout  = 8'b00000000; // 1871 :   0 - 0x0
      11'h750: dout  = 8'b00000000; // 1872 :   0 - 0x0 -- Background 0xea
      11'h751: dout  = 8'b00000000; // 1873 :   0 - 0x0
      11'h752: dout  = 8'b00000000; // 1874 :   0 - 0x0
      11'h753: dout  = 8'b00000000; // 1875 :   0 - 0x0
      11'h754: dout  = 8'b00000000; // 1876 :   0 - 0x0
      11'h755: dout  = 8'b00000000; // 1877 :   0 - 0x0
      11'h756: dout  = 8'b00000000; // 1878 :   0 - 0x0
      11'h757: dout  = 8'b00000000; // 1879 :   0 - 0x0
      11'h758: dout  = 8'b00000000; // 1880 :   0 - 0x0 -- Background 0xeb
      11'h759: dout  = 8'b00000000; // 1881 :   0 - 0x0
      11'h75A: dout  = 8'b00000000; // 1882 :   0 - 0x0
      11'h75B: dout  = 8'b00000000; // 1883 :   0 - 0x0
      11'h75C: dout  = 8'b00000000; // 1884 :   0 - 0x0
      11'h75D: dout  = 8'b00000000; // 1885 :   0 - 0x0
      11'h75E: dout  = 8'b00000000; // 1886 :   0 - 0x0
      11'h75F: dout  = 8'b00000000; // 1887 :   0 - 0x0
      11'h760: dout  = 8'b00000000; // 1888 :   0 - 0x0 -- Background 0xec
      11'h761: dout  = 8'b00000000; // 1889 :   0 - 0x0
      11'h762: dout  = 8'b00000000; // 1890 :   0 - 0x0
      11'h763: dout  = 8'b00000000; // 1891 :   0 - 0x0
      11'h764: dout  = 8'b00000000; // 1892 :   0 - 0x0
      11'h765: dout  = 8'b00000000; // 1893 :   0 - 0x0
      11'h766: dout  = 8'b00000000; // 1894 :   0 - 0x0
      11'h767: dout  = 8'b00000000; // 1895 :   0 - 0x0
      11'h768: dout  = 8'b00000000; // 1896 :   0 - 0x0 -- Background 0xed
      11'h769: dout  = 8'b00000000; // 1897 :   0 - 0x0
      11'h76A: dout  = 8'b00000000; // 1898 :   0 - 0x0
      11'h76B: dout  = 8'b00000000; // 1899 :   0 - 0x0
      11'h76C: dout  = 8'b00000000; // 1900 :   0 - 0x0
      11'h76D: dout  = 8'b00000000; // 1901 :   0 - 0x0
      11'h76E: dout  = 8'b00000000; // 1902 :   0 - 0x0
      11'h76F: dout  = 8'b00000000; // 1903 :   0 - 0x0
      11'h770: dout  = 8'b00000000; // 1904 :   0 - 0x0 -- Background 0xee
      11'h771: dout  = 8'b00000000; // 1905 :   0 - 0x0
      11'h772: dout  = 8'b00000000; // 1906 :   0 - 0x0
      11'h773: dout  = 8'b00000000; // 1907 :   0 - 0x0
      11'h774: dout  = 8'b00000000; // 1908 :   0 - 0x0
      11'h775: dout  = 8'b00000000; // 1909 :   0 - 0x0
      11'h776: dout  = 8'b00000000; // 1910 :   0 - 0x0
      11'h777: dout  = 8'b00000000; // 1911 :   0 - 0x0
      11'h778: dout  = 8'b00000000; // 1912 :   0 - 0x0 -- Background 0xef
      11'h779: dout  = 8'b00000000; // 1913 :   0 - 0x0
      11'h77A: dout  = 8'b00000000; // 1914 :   0 - 0x0
      11'h77B: dout  = 8'b00000000; // 1915 :   0 - 0x0
      11'h77C: dout  = 8'b00000000; // 1916 :   0 - 0x0
      11'h77D: dout  = 8'b00000000; // 1917 :   0 - 0x0
      11'h77E: dout  = 8'b00000000; // 1918 :   0 - 0x0
      11'h77F: dout  = 8'b00000000; // 1919 :   0 - 0x0
      11'h780: dout  = 8'b00000000; // 1920 :   0 - 0x0 -- Background 0xf0
      11'h781: dout  = 8'b00000000; // 1921 :   0 - 0x0
      11'h782: dout  = 8'b00000000; // 1922 :   0 - 0x0
      11'h783: dout  = 8'b00000000; // 1923 :   0 - 0x0
      11'h784: dout  = 8'b00000000; // 1924 :   0 - 0x0
      11'h785: dout  = 8'b00000000; // 1925 :   0 - 0x0
      11'h786: dout  = 8'b00000000; // 1926 :   0 - 0x0
      11'h787: dout  = 8'b00000000; // 1927 :   0 - 0x0
      11'h788: dout  = 8'b00000000; // 1928 :   0 - 0x0 -- Background 0xf1
      11'h789: dout  = 8'b00000000; // 1929 :   0 - 0x0
      11'h78A: dout  = 8'b00000000; // 1930 :   0 - 0x0
      11'h78B: dout  = 8'b00000000; // 1931 :   0 - 0x0
      11'h78C: dout  = 8'b00000000; // 1932 :   0 - 0x0
      11'h78D: dout  = 8'b00000000; // 1933 :   0 - 0x0
      11'h78E: dout  = 8'b00000000; // 1934 :   0 - 0x0
      11'h78F: dout  = 8'b00000000; // 1935 :   0 - 0x0
      11'h790: dout  = 8'b00000000; // 1936 :   0 - 0x0 -- Background 0xf2
      11'h791: dout  = 8'b00000000; // 1937 :   0 - 0x0
      11'h792: dout  = 8'b00000000; // 1938 :   0 - 0x0
      11'h793: dout  = 8'b00000000; // 1939 :   0 - 0x0
      11'h794: dout  = 8'b00000000; // 1940 :   0 - 0x0
      11'h795: dout  = 8'b00000000; // 1941 :   0 - 0x0
      11'h796: dout  = 8'b00000000; // 1942 :   0 - 0x0
      11'h797: dout  = 8'b00000000; // 1943 :   0 - 0x0
      11'h798: dout  = 8'b00000000; // 1944 :   0 - 0x0 -- Background 0xf3
      11'h799: dout  = 8'b00000000; // 1945 :   0 - 0x0
      11'h79A: dout  = 8'b00000000; // 1946 :   0 - 0x0
      11'h79B: dout  = 8'b00000000; // 1947 :   0 - 0x0
      11'h79C: dout  = 8'b00000000; // 1948 :   0 - 0x0
      11'h79D: dout  = 8'b00000000; // 1949 :   0 - 0x0
      11'h79E: dout  = 8'b00000000; // 1950 :   0 - 0x0
      11'h79F: dout  = 8'b00000000; // 1951 :   0 - 0x0
      11'h7A0: dout  = 8'b00000000; // 1952 :   0 - 0x0 -- Background 0xf4
      11'h7A1: dout  = 8'b00000000; // 1953 :   0 - 0x0
      11'h7A2: dout  = 8'b00000000; // 1954 :   0 - 0x0
      11'h7A3: dout  = 8'b00000000; // 1955 :   0 - 0x0
      11'h7A4: dout  = 8'b00000000; // 1956 :   0 - 0x0
      11'h7A5: dout  = 8'b00000000; // 1957 :   0 - 0x0
      11'h7A6: dout  = 8'b00000000; // 1958 :   0 - 0x0
      11'h7A7: dout  = 8'b00000000; // 1959 :   0 - 0x0
      11'h7A8: dout  = 8'b00000000; // 1960 :   0 - 0x0 -- Background 0xf5
      11'h7A9: dout  = 8'b00000000; // 1961 :   0 - 0x0
      11'h7AA: dout  = 8'b00000000; // 1962 :   0 - 0x0
      11'h7AB: dout  = 8'b00000000; // 1963 :   0 - 0x0
      11'h7AC: dout  = 8'b00000000; // 1964 :   0 - 0x0
      11'h7AD: dout  = 8'b00000000; // 1965 :   0 - 0x0
      11'h7AE: dout  = 8'b00000000; // 1966 :   0 - 0x0
      11'h7AF: dout  = 8'b00000000; // 1967 :   0 - 0x0
      11'h7B0: dout  = 8'b00000000; // 1968 :   0 - 0x0 -- Background 0xf6
      11'h7B1: dout  = 8'b00000000; // 1969 :   0 - 0x0
      11'h7B2: dout  = 8'b00000000; // 1970 :   0 - 0x0
      11'h7B3: dout  = 8'b00000000; // 1971 :   0 - 0x0
      11'h7B4: dout  = 8'b00000000; // 1972 :   0 - 0x0
      11'h7B5: dout  = 8'b00000000; // 1973 :   0 - 0x0
      11'h7B6: dout  = 8'b00000000; // 1974 :   0 - 0x0
      11'h7B7: dout  = 8'b00000000; // 1975 :   0 - 0x0
      11'h7B8: dout  = 8'b00000000; // 1976 :   0 - 0x0 -- Background 0xf7
      11'h7B9: dout  = 8'b00000000; // 1977 :   0 - 0x0
      11'h7BA: dout  = 8'b00000000; // 1978 :   0 - 0x0
      11'h7BB: dout  = 8'b00000000; // 1979 :   0 - 0x0
      11'h7BC: dout  = 8'b00000000; // 1980 :   0 - 0x0
      11'h7BD: dout  = 8'b00000000; // 1981 :   0 - 0x0
      11'h7BE: dout  = 8'b00000000; // 1982 :   0 - 0x0
      11'h7BF: dout  = 8'b00000000; // 1983 :   0 - 0x0
      11'h7C0: dout  = 8'b00000000; // 1984 :   0 - 0x0 -- Background 0xf8
      11'h7C1: dout  = 8'b00000000; // 1985 :   0 - 0x0
      11'h7C2: dout  = 8'b00000000; // 1986 :   0 - 0x0
      11'h7C3: dout  = 8'b00000000; // 1987 :   0 - 0x0
      11'h7C4: dout  = 8'b00000000; // 1988 :   0 - 0x0
      11'h7C5: dout  = 8'b00000000; // 1989 :   0 - 0x0
      11'h7C6: dout  = 8'b00000000; // 1990 :   0 - 0x0
      11'h7C7: dout  = 8'b00000000; // 1991 :   0 - 0x0
      11'h7C8: dout  = 8'b00000000; // 1992 :   0 - 0x0 -- Background 0xf9
      11'h7C9: dout  = 8'b00000000; // 1993 :   0 - 0x0
      11'h7CA: dout  = 8'b00000000; // 1994 :   0 - 0x0
      11'h7CB: dout  = 8'b00000000; // 1995 :   0 - 0x0
      11'h7CC: dout  = 8'b00000000; // 1996 :   0 - 0x0
      11'h7CD: dout  = 8'b00000000; // 1997 :   0 - 0x0
      11'h7CE: dout  = 8'b00000000; // 1998 :   0 - 0x0
      11'h7CF: dout  = 8'b00000000; // 1999 :   0 - 0x0
      11'h7D0: dout  = 8'b00000000; // 2000 :   0 - 0x0 -- Background 0xfa
      11'h7D1: dout  = 8'b00000000; // 2001 :   0 - 0x0
      11'h7D2: dout  = 8'b00000000; // 2002 :   0 - 0x0
      11'h7D3: dout  = 8'b00000000; // 2003 :   0 - 0x0
      11'h7D4: dout  = 8'b00000000; // 2004 :   0 - 0x0
      11'h7D5: dout  = 8'b00000000; // 2005 :   0 - 0x0
      11'h7D6: dout  = 8'b00000000; // 2006 :   0 - 0x0
      11'h7D7: dout  = 8'b00000000; // 2007 :   0 - 0x0
      11'h7D8: dout  = 8'b00000000; // 2008 :   0 - 0x0 -- Background 0xfb
      11'h7D9: dout  = 8'b00000000; // 2009 :   0 - 0x0
      11'h7DA: dout  = 8'b00000000; // 2010 :   0 - 0x0
      11'h7DB: dout  = 8'b00000000; // 2011 :   0 - 0x0
      11'h7DC: dout  = 8'b00000000; // 2012 :   0 - 0x0
      11'h7DD: dout  = 8'b00000000; // 2013 :   0 - 0x0
      11'h7DE: dout  = 8'b00000000; // 2014 :   0 - 0x0
      11'h7DF: dout  = 8'b00000000; // 2015 :   0 - 0x0
      11'h7E0: dout  = 8'b00000000; // 2016 :   0 - 0x0 -- Background 0xfc
      11'h7E1: dout  = 8'b00000000; // 2017 :   0 - 0x0
      11'h7E2: dout  = 8'b00000000; // 2018 :   0 - 0x0
      11'h7E3: dout  = 8'b00000000; // 2019 :   0 - 0x0
      11'h7E4: dout  = 8'b00000000; // 2020 :   0 - 0x0
      11'h7E5: dout  = 8'b00000000; // 2021 :   0 - 0x0
      11'h7E6: dout  = 8'b00000000; // 2022 :   0 - 0x0
      11'h7E7: dout  = 8'b00000000; // 2023 :   0 - 0x0
      11'h7E8: dout  = 8'b00000000; // 2024 :   0 - 0x0 -- Background 0xfd
      11'h7E9: dout  = 8'b00000000; // 2025 :   0 - 0x0
      11'h7EA: dout  = 8'b00000000; // 2026 :   0 - 0x0
      11'h7EB: dout  = 8'b00000000; // 2027 :   0 - 0x0
      11'h7EC: dout  = 8'b00000000; // 2028 :   0 - 0x0
      11'h7ED: dout  = 8'b00000000; // 2029 :   0 - 0x0
      11'h7EE: dout  = 8'b00000000; // 2030 :   0 - 0x0
      11'h7EF: dout  = 8'b00000000; // 2031 :   0 - 0x0
      11'h7F0: dout  = 8'b00000000; // 2032 :   0 - 0x0 -- Background 0xfe
      11'h7F1: dout  = 8'b00000000; // 2033 :   0 - 0x0
      11'h7F2: dout  = 8'b00000000; // 2034 :   0 - 0x0
      11'h7F3: dout  = 8'b00000000; // 2035 :   0 - 0x0
      11'h7F4: dout  = 8'b00000000; // 2036 :   0 - 0x0
      11'h7F5: dout  = 8'b00000000; // 2037 :   0 - 0x0
      11'h7F6: dout  = 8'b00000000; // 2038 :   0 - 0x0
      11'h7F7: dout  = 8'b00000000; // 2039 :   0 - 0x0
      11'h7F8: dout  = 8'b00000000; // 2040 :   0 - 0x0 -- Background 0xff
      11'h7F9: dout  = 8'b00000000; // 2041 :   0 - 0x0
      11'h7FA: dout  = 8'b00000000; // 2042 :   0 - 0x0
      11'h7FB: dout  = 8'b00000000; // 2043 :   0 - 0x0
      11'h7FC: dout  = 8'b00000000; // 2044 :   0 - 0x0
      11'h7FD: dout  = 8'b00000000; // 2045 :   0 - 0x0
      11'h7FE: dout  = 8'b00000000; // 2046 :   0 - 0x0
      11'h7FF: dout  = 8'b00000000; // 2047 :   0 - 0x0
    endcase
  end

endmodule
