//- Autcmatically generated verilog ROM from a NES memory file----
//-   NAME TABLE
// https://wiki.nesdev.com/w/index.php/PPU_nametables


//-  Original memory dump file name: nova_ntable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_NTABLE_NOVA_00
  (
     //input     clk,   // clock
     input      [11-1:0] addr,  //2048 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
     //----- Name Table 0---------
      11'h0: dout  = 8'b00110000; //    0 :  48 - 0x30 -- line 0x0
      11'h1: dout  = 8'b00111111; //    1 :  63 - 0x3f
      11'h2: dout  = 8'b00110000; //    2 :  48 - 0x30
      11'h3: dout  = 8'b00111111; //    3 :  63 - 0x3f
      11'h4: dout  = 8'b00110000; //    4 :  48 - 0x30
      11'h5: dout  = 8'b00111111; //    5 :  63 - 0x3f
      11'h6: dout  = 8'b00110000; //    6 :  48 - 0x30
      11'h7: dout  = 8'b00111111; //    7 :  63 - 0x3f
      11'h8: dout  = 8'b00110000; //    8 :  48 - 0x30
      11'h9: dout  = 8'b00111111; //    9 :  63 - 0x3f
      11'hA: dout  = 8'b00110000; //   10 :  48 - 0x30
      11'hB: dout  = 8'b00111111; //   11 :  63 - 0x3f
      11'hC: dout  = 8'b00110000; //   12 :  48 - 0x30
      11'hD: dout  = 8'b00111111; //   13 :  63 - 0x3f
      11'hE: dout  = 8'b00110000; //   14 :  48 - 0x30
      11'hF: dout  = 8'b00111111; //   15 :  63 - 0x3f
      11'h10: dout  = 8'b00110000; //   16 :  48 - 0x30
      11'h11: dout  = 8'b00111111; //   17 :  63 - 0x3f
      11'h12: dout  = 8'b00110000; //   18 :  48 - 0x30
      11'h13: dout  = 8'b00111111; //   19 :  63 - 0x3f
      11'h14: dout  = 8'b01110000; //   20 : 112 - 0x70
      11'h15: dout  = 8'b01110001; //   21 : 113 - 0x71
      11'h16: dout  = 8'b01110001; //   22 : 113 - 0x71
      11'h17: dout  = 8'b01110001; //   23 : 113 - 0x71
      11'h18: dout  = 8'b01110001; //   24 : 113 - 0x71
      11'h19: dout  = 8'b01110001; //   25 : 113 - 0x71
      11'h1A: dout  = 8'b01110001; //   26 : 113 - 0x71
      11'h1B: dout  = 8'b01110001; //   27 : 113 - 0x71
      11'h1C: dout  = 8'b01110001; //   28 : 113 - 0x71
      11'h1D: dout  = 8'b01110001; //   29 : 113 - 0x71
      11'h1E: dout  = 8'b01110001; //   30 : 113 - 0x71
      11'h1F: dout  = 8'b01110001; //   31 : 113 - 0x71
      11'h20: dout  = 8'b00111111; //   32 :  63 - 0x3f -- line 0x1
      11'h21: dout  = 8'b00110000; //   33 :  48 - 0x30
      11'h22: dout  = 8'b00111111; //   34 :  63 - 0x3f
      11'h23: dout  = 8'b00110000; //   35 :  48 - 0x30
      11'h24: dout  = 8'b00111111; //   36 :  63 - 0x3f
      11'h25: dout  = 8'b00110000; //   37 :  48 - 0x30
      11'h26: dout  = 8'b00111111; //   38 :  63 - 0x3f
      11'h27: dout  = 8'b00110000; //   39 :  48 - 0x30
      11'h28: dout  = 8'b00111111; //   40 :  63 - 0x3f
      11'h29: dout  = 8'b00110000; //   41 :  48 - 0x30
      11'h2A: dout  = 8'b00111111; //   42 :  63 - 0x3f
      11'h2B: dout  = 8'b00110000; //   43 :  48 - 0x30
      11'h2C: dout  = 8'b00111111; //   44 :  63 - 0x3f
      11'h2D: dout  = 8'b00110000; //   45 :  48 - 0x30
      11'h2E: dout  = 8'b00111111; //   46 :  63 - 0x3f
      11'h2F: dout  = 8'b00110000; //   47 :  48 - 0x30
      11'h30: dout  = 8'b00111111; //   48 :  63 - 0x3f
      11'h31: dout  = 8'b00110000; //   49 :  48 - 0x30
      11'h32: dout  = 8'b00111111; //   50 :  63 - 0x3f
      11'h33: dout  = 8'b00110000; //   51 :  48 - 0x30
      11'h34: dout  = 8'b01100000; //   52 :  96 - 0x60
      11'h35: dout  = 8'b01110111; //   53 : 119 - 0x77
      11'h36: dout  = 8'b01110111; //   54 : 119 - 0x77
      11'h37: dout  = 8'b01110111; //   55 : 119 - 0x77
      11'h38: dout  = 8'b01110111; //   56 : 119 - 0x77
      11'h39: dout  = 8'b01110111; //   57 : 119 - 0x77
      11'h3A: dout  = 8'b01110111; //   58 : 119 - 0x77
      11'h3B: dout  = 8'b01110111; //   59 : 119 - 0x77
      11'h3C: dout  = 8'b01110111; //   60 : 119 - 0x77
      11'h3D: dout  = 8'b01110111; //   61 : 119 - 0x77
      11'h3E: dout  = 8'b01110111; //   62 : 119 - 0x77
      11'h3F: dout  = 8'b01110111; //   63 : 119 - 0x77
      11'h40: dout  = 8'b00110000; //   64 :  48 - 0x30 -- line 0x2
      11'h41: dout  = 8'b00111111; //   65 :  63 - 0x3f
      11'h42: dout  = 8'b00110000; //   66 :  48 - 0x30
      11'h43: dout  = 8'b00111111; //   67 :  63 - 0x3f
      11'h44: dout  = 8'b00110000; //   68 :  48 - 0x30
      11'h45: dout  = 8'b00111111; //   69 :  63 - 0x3f
      11'h46: dout  = 8'b00110000; //   70 :  48 - 0x30
      11'h47: dout  = 8'b00111111; //   71 :  63 - 0x3f
      11'h48: dout  = 8'b00110000; //   72 :  48 - 0x30
      11'h49: dout  = 8'b00111111; //   73 :  63 - 0x3f
      11'h4A: dout  = 8'b00110000; //   74 :  48 - 0x30
      11'h4B: dout  = 8'b00111111; //   75 :  63 - 0x3f
      11'h4C: dout  = 8'b00110000; //   76 :  48 - 0x30
      11'h4D: dout  = 8'b00111111; //   77 :  63 - 0x3f
      11'h4E: dout  = 8'b00110000; //   78 :  48 - 0x30
      11'h4F: dout  = 8'b00111111; //   79 :  63 - 0x3f
      11'h50: dout  = 8'b00110000; //   80 :  48 - 0x30
      11'h51: dout  = 8'b00111111; //   81 :  63 - 0x3f
      11'h52: dout  = 8'b00110000; //   82 :  48 - 0x30
      11'h53: dout  = 8'b00111111; //   83 :  63 - 0x3f
      11'h54: dout  = 8'b00111001; //   84 :  57 - 0x39
      11'h55: dout  = 8'b00111001; //   85 :  57 - 0x39
      11'h56: dout  = 8'b00111001; //   86 :  57 - 0x39
      11'h57: dout  = 8'b00111001; //   87 :  57 - 0x39
      11'h58: dout  = 8'b00111001; //   88 :  57 - 0x39
      11'h59: dout  = 8'b00111001; //   89 :  57 - 0x39
      11'h5A: dout  = 8'b00111001; //   90 :  57 - 0x39
      11'h5B: dout  = 8'b00111001; //   91 :  57 - 0x39
      11'h5C: dout  = 8'b00111001; //   92 :  57 - 0x39
      11'h5D: dout  = 8'b00111001; //   93 :  57 - 0x39
      11'h5E: dout  = 8'b00111001; //   94 :  57 - 0x39
      11'h5F: dout  = 8'b00111001; //   95 :  57 - 0x39
      11'h60: dout  = 8'b00111111; //   96 :  63 - 0x3f -- line 0x3
      11'h61: dout  = 8'b00110000; //   97 :  48 - 0x30
      11'h62: dout  = 8'b00111111; //   98 :  63 - 0x3f
      11'h63: dout  = 8'b00110000; //   99 :  48 - 0x30
      11'h64: dout  = 8'b00111111; //  100 :  63 - 0x3f
      11'h65: dout  = 8'b00110000; //  101 :  48 - 0x30
      11'h66: dout  = 8'b00111111; //  102 :  63 - 0x3f
      11'h67: dout  = 8'b00110000; //  103 :  48 - 0x30
      11'h68: dout  = 8'b00111111; //  104 :  63 - 0x3f
      11'h69: dout  = 8'b00110000; //  105 :  48 - 0x30
      11'h6A: dout  = 8'b00111111; //  106 :  63 - 0x3f
      11'h6B: dout  = 8'b00110000; //  107 :  48 - 0x30
      11'h6C: dout  = 8'b00111111; //  108 :  63 - 0x3f
      11'h6D: dout  = 8'b00110000; //  109 :  48 - 0x30
      11'h6E: dout  = 8'b00111111; //  110 :  63 - 0x3f
      11'h6F: dout  = 8'b00110000; //  111 :  48 - 0x30
      11'h70: dout  = 8'b00111111; //  112 :  63 - 0x3f
      11'h71: dout  = 8'b00110000; //  113 :  48 - 0x30
      11'h72: dout  = 8'b00111111; //  114 :  63 - 0x3f
      11'h73: dout  = 8'b00110000; //  115 :  48 - 0x30
      11'h74: dout  = 8'b00111111; //  116 :  63 - 0x3f
      11'h75: dout  = 8'b00111111; //  117 :  63 - 0x3f
      11'h76: dout  = 8'b00111111; //  118 :  63 - 0x3f
      11'h77: dout  = 8'b00111111; //  119 :  63 - 0x3f
      11'h78: dout  = 8'b00111111; //  120 :  63 - 0x3f
      11'h79: dout  = 8'b00111111; //  121 :  63 - 0x3f
      11'h7A: dout  = 8'b00111111; //  122 :  63 - 0x3f
      11'h7B: dout  = 8'b00111111; //  123 :  63 - 0x3f
      11'h7C: dout  = 8'b00111111; //  124 :  63 - 0x3f
      11'h7D: dout  = 8'b00111111; //  125 :  63 - 0x3f
      11'h7E: dout  = 8'b00111111; //  126 :  63 - 0x3f
      11'h7F: dout  = 8'b00111111; //  127 :  63 - 0x3f
      11'h80: dout  = 8'b00111111; //  128 :  63 - 0x3f -- line 0x4
      11'h81: dout  = 8'b00111111; //  129 :  63 - 0x3f
      11'h82: dout  = 8'b00111111; //  130 :  63 - 0x3f
      11'h83: dout  = 8'b00111111; //  131 :  63 - 0x3f
      11'h84: dout  = 8'b00111111; //  132 :  63 - 0x3f
      11'h85: dout  = 8'b00111111; //  133 :  63 - 0x3f
      11'h86: dout  = 8'b00111111; //  134 :  63 - 0x3f
      11'h87: dout  = 8'b00111111; //  135 :  63 - 0x3f
      11'h88: dout  = 8'b00111111; //  136 :  63 - 0x3f
      11'h89: dout  = 8'b00111111; //  137 :  63 - 0x3f
      11'h8A: dout  = 8'b00111111; //  138 :  63 - 0x3f
      11'h8B: dout  = 8'b00111111; //  139 :  63 - 0x3f
      11'h8C: dout  = 8'b00111111; //  140 :  63 - 0x3f
      11'h8D: dout  = 8'b00111111; //  141 :  63 - 0x3f
      11'h8E: dout  = 8'b00111111; //  142 :  63 - 0x3f
      11'h8F: dout  = 8'b00111111; //  143 :  63 - 0x3f
      11'h90: dout  = 8'b00111111; //  144 :  63 - 0x3f
      11'h91: dout  = 8'b00111111; //  145 :  63 - 0x3f
      11'h92: dout  = 8'b00111111; //  146 :  63 - 0x3f
      11'h93: dout  = 8'b00111111; //  147 :  63 - 0x3f
      11'h94: dout  = 8'b00111111; //  148 :  63 - 0x3f
      11'h95: dout  = 8'b00111111; //  149 :  63 - 0x3f
      11'h96: dout  = 8'b00111111; //  150 :  63 - 0x3f
      11'h97: dout  = 8'b00111111; //  151 :  63 - 0x3f
      11'h98: dout  = 8'b00111111; //  152 :  63 - 0x3f
      11'h99: dout  = 8'b00111111; //  153 :  63 - 0x3f
      11'h9A: dout  = 8'b00000100; //  154 :   4 - 0x4
      11'h9B: dout  = 8'b00000110; //  155 :   6 - 0x6
      11'h9C: dout  = 8'b00111111; //  156 :  63 - 0x3f
      11'h9D: dout  = 8'b00111111; //  157 :  63 - 0x3f
      11'h9E: dout  = 8'b00010100; //  158 :  20 - 0x14
      11'h9F: dout  = 8'b00010110; //  159 :  22 - 0x16
      11'hA0: dout  = 8'b00111111; //  160 :  63 - 0x3f -- line 0x5
      11'hA1: dout  = 8'b00111111; //  161 :  63 - 0x3f
      11'hA2: dout  = 8'b00111111; //  162 :  63 - 0x3f
      11'hA3: dout  = 8'b00111111; //  163 :  63 - 0x3f
      11'hA4: dout  = 8'b00111111; //  164 :  63 - 0x3f
      11'hA5: dout  = 8'b00111111; //  165 :  63 - 0x3f
      11'hA6: dout  = 8'b00111111; //  166 :  63 - 0x3f
      11'hA7: dout  = 8'b00111111; //  167 :  63 - 0x3f
      11'hA8: dout  = 8'b00111111; //  168 :  63 - 0x3f
      11'hA9: dout  = 8'b00111111; //  169 :  63 - 0x3f
      11'hAA: dout  = 8'b00111111; //  170 :  63 - 0x3f
      11'hAB: dout  = 8'b00111111; //  171 :  63 - 0x3f
      11'hAC: dout  = 8'b00111111; //  172 :  63 - 0x3f
      11'hAD: dout  = 8'b00111111; //  173 :  63 - 0x3f
      11'hAE: dout  = 8'b00111111; //  174 :  63 - 0x3f
      11'hAF: dout  = 8'b00111111; //  175 :  63 - 0x3f
      11'hB0: dout  = 8'b00111111; //  176 :  63 - 0x3f
      11'hB1: dout  = 8'b00111111; //  177 :  63 - 0x3f
      11'hB2: dout  = 8'b00111111; //  178 :  63 - 0x3f
      11'hB3: dout  = 8'b00111111; //  179 :  63 - 0x3f
      11'hB4: dout  = 8'b00111111; //  180 :  63 - 0x3f
      11'hB5: dout  = 8'b00111111; //  181 :  63 - 0x3f
      11'hB6: dout  = 8'b00111111; //  182 :  63 - 0x3f
      11'hB7: dout  = 8'b00111111; //  183 :  63 - 0x3f
      11'hB8: dout  = 8'b00111111; //  184 :  63 - 0x3f
      11'hB9: dout  = 8'b00111111; //  185 :  63 - 0x3f
      11'hBA: dout  = 8'b00000101; //  186 :   5 - 0x5
      11'hBB: dout  = 8'b00000111; //  187 :   7 - 0x7
      11'hBC: dout  = 8'b00111111; //  188 :  63 - 0x3f
      11'hBD: dout  = 8'b00111111; //  189 :  63 - 0x3f
      11'hBE: dout  = 8'b00010101; //  190 :  21 - 0x15
      11'hBF: dout  = 8'b00010111; //  191 :  23 - 0x17
      11'hC0: dout  = 8'b00111111; //  192 :  63 - 0x3f -- line 0x6
      11'hC1: dout  = 8'b00111111; //  193 :  63 - 0x3f
      11'hC2: dout  = 8'b00111111; //  194 :  63 - 0x3f
      11'hC3: dout  = 8'b00111111; //  195 :  63 - 0x3f
      11'hC4: dout  = 8'b00111111; //  196 :  63 - 0x3f
      11'hC5: dout  = 8'b00111111; //  197 :  63 - 0x3f
      11'hC6: dout  = 8'b00111111; //  198 :  63 - 0x3f
      11'hC7: dout  = 8'b00111111; //  199 :  63 - 0x3f
      11'hC8: dout  = 8'b00111111; //  200 :  63 - 0x3f
      11'hC9: dout  = 8'b00111111; //  201 :  63 - 0x3f
      11'hCA: dout  = 8'b00111111; //  202 :  63 - 0x3f
      11'hCB: dout  = 8'b00111111; //  203 :  63 - 0x3f
      11'hCC: dout  = 8'b00111111; //  204 :  63 - 0x3f
      11'hCD: dout  = 8'b00111111; //  205 :  63 - 0x3f
      11'hCE: dout  = 8'b00111111; //  206 :  63 - 0x3f
      11'hCF: dout  = 8'b00111111; //  207 :  63 - 0x3f
      11'hD0: dout  = 8'b00111111; //  208 :  63 - 0x3f
      11'hD1: dout  = 8'b00111111; //  209 :  63 - 0x3f
      11'hD2: dout  = 8'b00111111; //  210 :  63 - 0x3f
      11'hD3: dout  = 8'b00111111; //  211 :  63 - 0x3f
      11'hD4: dout  = 8'b00111111; //  212 :  63 - 0x3f
      11'hD5: dout  = 8'b00111111; //  213 :  63 - 0x3f
      11'hD6: dout  = 8'b00111111; //  214 :  63 - 0x3f
      11'hD7: dout  = 8'b00111111; //  215 :  63 - 0x3f
      11'hD8: dout  = 8'b00111111; //  216 :  63 - 0x3f
      11'hD9: dout  = 8'b00111111; //  217 :  63 - 0x3f
      11'hDA: dout  = 8'b00111111; //  218 :  63 - 0x3f
      11'hDB: dout  = 8'b00111111; //  219 :  63 - 0x3f
      11'hDC: dout  = 8'b00111111; //  220 :  63 - 0x3f
      11'hDD: dout  = 8'b00111111; //  221 :  63 - 0x3f
      11'hDE: dout  = 8'b00111111; //  222 :  63 - 0x3f
      11'hDF: dout  = 8'b00111111; //  223 :  63 - 0x3f
      11'hE0: dout  = 8'b00111111; //  224 :  63 - 0x3f -- line 0x7
      11'hE1: dout  = 8'b00111111; //  225 :  63 - 0x3f
      11'hE2: dout  = 8'b00111111; //  226 :  63 - 0x3f
      11'hE3: dout  = 8'b00111111; //  227 :  63 - 0x3f
      11'hE4: dout  = 8'b00111111; //  228 :  63 - 0x3f
      11'hE5: dout  = 8'b00111111; //  229 :  63 - 0x3f
      11'hE6: dout  = 8'b00111111; //  230 :  63 - 0x3f
      11'hE7: dout  = 8'b00111111; //  231 :  63 - 0x3f
      11'hE8: dout  = 8'b00111111; //  232 :  63 - 0x3f
      11'hE9: dout  = 8'b00111111; //  233 :  63 - 0x3f
      11'hEA: dout  = 8'b00111111; //  234 :  63 - 0x3f
      11'hEB: dout  = 8'b00111111; //  235 :  63 - 0x3f
      11'hEC: dout  = 8'b00111111; //  236 :  63 - 0x3f
      11'hED: dout  = 8'b00111111; //  237 :  63 - 0x3f
      11'hEE: dout  = 8'b00111111; //  238 :  63 - 0x3f
      11'hEF: dout  = 8'b00111111; //  239 :  63 - 0x3f
      11'hF0: dout  = 8'b00111111; //  240 :  63 - 0x3f
      11'hF1: dout  = 8'b00111111; //  241 :  63 - 0x3f
      11'hF2: dout  = 8'b00111111; //  242 :  63 - 0x3f
      11'hF3: dout  = 8'b00111111; //  243 :  63 - 0x3f
      11'hF4: dout  = 8'b00111111; //  244 :  63 - 0x3f
      11'hF5: dout  = 8'b00111111; //  245 :  63 - 0x3f
      11'hF6: dout  = 8'b00111111; //  246 :  63 - 0x3f
      11'hF7: dout  = 8'b00111111; //  247 :  63 - 0x3f
      11'hF8: dout  = 8'b00111111; //  248 :  63 - 0x3f
      11'hF9: dout  = 8'b00111111; //  249 :  63 - 0x3f
      11'hFA: dout  = 8'b00111111; //  250 :  63 - 0x3f
      11'hFB: dout  = 8'b00111111; //  251 :  63 - 0x3f
      11'hFC: dout  = 8'b00111111; //  252 :  63 - 0x3f
      11'hFD: dout  = 8'b00111111; //  253 :  63 - 0x3f
      11'hFE: dout  = 8'b00111111; //  254 :  63 - 0x3f
      11'hFF: dout  = 8'b00111111; //  255 :  63 - 0x3f
      11'h100: dout  = 8'b00111111; //  256 :  63 - 0x3f -- line 0x8
      11'h101: dout  = 8'b00111111; //  257 :  63 - 0x3f
      11'h102: dout  = 8'b00111111; //  258 :  63 - 0x3f
      11'h103: dout  = 8'b00111111; //  259 :  63 - 0x3f
      11'h104: dout  = 8'b00111111; //  260 :  63 - 0x3f
      11'h105: dout  = 8'b00111111; //  261 :  63 - 0x3f
      11'h106: dout  = 8'b00111111; //  262 :  63 - 0x3f
      11'h107: dout  = 8'b00111111; //  263 :  63 - 0x3f
      11'h108: dout  = 8'b00111111; //  264 :  63 - 0x3f
      11'h109: dout  = 8'b00111111; //  265 :  63 - 0x3f
      11'h10A: dout  = 8'b00111111; //  266 :  63 - 0x3f
      11'h10B: dout  = 8'b00111111; //  267 :  63 - 0x3f
      11'h10C: dout  = 8'b00111111; //  268 :  63 - 0x3f
      11'h10D: dout  = 8'b00111111; //  269 :  63 - 0x3f
      11'h10E: dout  = 8'b00111111; //  270 :  63 - 0x3f
      11'h10F: dout  = 8'b00111111; //  271 :  63 - 0x3f
      11'h110: dout  = 8'b00111111; //  272 :  63 - 0x3f
      11'h111: dout  = 8'b00111111; //  273 :  63 - 0x3f
      11'h112: dout  = 8'b00111111; //  274 :  63 - 0x3f
      11'h113: dout  = 8'b00111111; //  275 :  63 - 0x3f
      11'h114: dout  = 8'b00001100; //  276 :  12 - 0xc
      11'h115: dout  = 8'b00001110; //  277 :  14 - 0xe
      11'h116: dout  = 8'b00111111; //  278 :  63 - 0x3f
      11'h117: dout  = 8'b00111111; //  279 :  63 - 0x3f
      11'h118: dout  = 8'b00111111; //  280 :  63 - 0x3f
      11'h119: dout  = 8'b00111111; //  281 :  63 - 0x3f
      11'h11A: dout  = 8'b00111111; //  282 :  63 - 0x3f
      11'h11B: dout  = 8'b00111111; //  283 :  63 - 0x3f
      11'h11C: dout  = 8'b00111111; //  284 :  63 - 0x3f
      11'h11D: dout  = 8'b00111111; //  285 :  63 - 0x3f
      11'h11E: dout  = 8'b00111111; //  286 :  63 - 0x3f
      11'h11F: dout  = 8'b00111111; //  287 :  63 - 0x3f
      11'h120: dout  = 8'b00111111; //  288 :  63 - 0x3f -- line 0x9
      11'h121: dout  = 8'b00111111; //  289 :  63 - 0x3f
      11'h122: dout  = 8'b00111111; //  290 :  63 - 0x3f
      11'h123: dout  = 8'b00111111; //  291 :  63 - 0x3f
      11'h124: dout  = 8'b00111111; //  292 :  63 - 0x3f
      11'h125: dout  = 8'b00111111; //  293 :  63 - 0x3f
      11'h126: dout  = 8'b00111111; //  294 :  63 - 0x3f
      11'h127: dout  = 8'b00111111; //  295 :  63 - 0x3f
      11'h128: dout  = 8'b00111111; //  296 :  63 - 0x3f
      11'h129: dout  = 8'b00111111; //  297 :  63 - 0x3f
      11'h12A: dout  = 8'b00111111; //  298 :  63 - 0x3f
      11'h12B: dout  = 8'b00111111; //  299 :  63 - 0x3f
      11'h12C: dout  = 8'b00111111; //  300 :  63 - 0x3f
      11'h12D: dout  = 8'b00111111; //  301 :  63 - 0x3f
      11'h12E: dout  = 8'b00111111; //  302 :  63 - 0x3f
      11'h12F: dout  = 8'b00111111; //  303 :  63 - 0x3f
      11'h130: dout  = 8'b00111111; //  304 :  63 - 0x3f
      11'h131: dout  = 8'b00111111; //  305 :  63 - 0x3f
      11'h132: dout  = 8'b00111111; //  306 :  63 - 0x3f
      11'h133: dout  = 8'b00111111; //  307 :  63 - 0x3f
      11'h134: dout  = 8'b00001101; //  308 :  13 - 0xd
      11'h135: dout  = 8'b00001111; //  309 :  15 - 0xf
      11'h136: dout  = 8'b00111111; //  310 :  63 - 0x3f
      11'h137: dout  = 8'b00111111; //  311 :  63 - 0x3f
      11'h138: dout  = 8'b00111111; //  312 :  63 - 0x3f
      11'h139: dout  = 8'b00111111; //  313 :  63 - 0x3f
      11'h13A: dout  = 8'b00111111; //  314 :  63 - 0x3f
      11'h13B: dout  = 8'b00111111; //  315 :  63 - 0x3f
      11'h13C: dout  = 8'b00111111; //  316 :  63 - 0x3f
      11'h13D: dout  = 8'b00111111; //  317 :  63 - 0x3f
      11'h13E: dout  = 8'b00111111; //  318 :  63 - 0x3f
      11'h13F: dout  = 8'b00111111; //  319 :  63 - 0x3f
      11'h140: dout  = 8'b00111111; //  320 :  63 - 0x3f -- line 0xa
      11'h141: dout  = 8'b00111111; //  321 :  63 - 0x3f
      11'h142: dout  = 8'b00111111; //  322 :  63 - 0x3f
      11'h143: dout  = 8'b00111111; //  323 :  63 - 0x3f
      11'h144: dout  = 8'b00111111; //  324 :  63 - 0x3f
      11'h145: dout  = 8'b00111111; //  325 :  63 - 0x3f
      11'h146: dout  = 8'b00111111; //  326 :  63 - 0x3f
      11'h147: dout  = 8'b00111111; //  327 :  63 - 0x3f
      11'h148: dout  = 8'b00111111; //  328 :  63 - 0x3f
      11'h149: dout  = 8'b00111111; //  329 :  63 - 0x3f
      11'h14A: dout  = 8'b00111111; //  330 :  63 - 0x3f
      11'h14B: dout  = 8'b00111111; //  331 :  63 - 0x3f
      11'h14C: dout  = 8'b00111111; //  332 :  63 - 0x3f
      11'h14D: dout  = 8'b00111111; //  333 :  63 - 0x3f
      11'h14E: dout  = 8'b00111111; //  334 :  63 - 0x3f
      11'h14F: dout  = 8'b00111111; //  335 :  63 - 0x3f
      11'h150: dout  = 8'b00111111; //  336 :  63 - 0x3f
      11'h151: dout  = 8'b00111111; //  337 :  63 - 0x3f
      11'h152: dout  = 8'b00111111; //  338 :  63 - 0x3f
      11'h153: dout  = 8'b00111111; //  339 :  63 - 0x3f
      11'h154: dout  = 8'b01010111; //  340 :  87 - 0x57
      11'h155: dout  = 8'b01011000; //  341 :  88 - 0x58
      11'h156: dout  = 8'b01011000; //  342 :  88 - 0x58
      11'h157: dout  = 8'b01011000; //  343 :  88 - 0x58
      11'h158: dout  = 8'b01011000; //  344 :  88 - 0x58
      11'h159: dout  = 8'b01011000; //  345 :  88 - 0x58
      11'h15A: dout  = 8'b01011000; //  346 :  88 - 0x58
      11'h15B: dout  = 8'b01011000; //  347 :  88 - 0x58
      11'h15C: dout  = 8'b01011000; //  348 :  88 - 0x58
      11'h15D: dout  = 8'b01011000; //  349 :  88 - 0x58
      11'h15E: dout  = 8'b01011000; //  350 :  88 - 0x58
      11'h15F: dout  = 8'b01011000; //  351 :  88 - 0x58
      11'h160: dout  = 8'b00111111; //  352 :  63 - 0x3f -- line 0xb
      11'h161: dout  = 8'b00111111; //  353 :  63 - 0x3f
      11'h162: dout  = 8'b00111111; //  354 :  63 - 0x3f
      11'h163: dout  = 8'b00111111; //  355 :  63 - 0x3f
      11'h164: dout  = 8'b00111111; //  356 :  63 - 0x3f
      11'h165: dout  = 8'b00111111; //  357 :  63 - 0x3f
      11'h166: dout  = 8'b00111111; //  358 :  63 - 0x3f
      11'h167: dout  = 8'b00111111; //  359 :  63 - 0x3f
      11'h168: dout  = 8'b00111111; //  360 :  63 - 0x3f
      11'h169: dout  = 8'b00111111; //  361 :  63 - 0x3f
      11'h16A: dout  = 8'b00111111; //  362 :  63 - 0x3f
      11'h16B: dout  = 8'b00111111; //  363 :  63 - 0x3f
      11'h16C: dout  = 8'b00111111; //  364 :  63 - 0x3f
      11'h16D: dout  = 8'b00111111; //  365 :  63 - 0x3f
      11'h16E: dout  = 8'b00111111; //  366 :  63 - 0x3f
      11'h16F: dout  = 8'b00111111; //  367 :  63 - 0x3f
      11'h170: dout  = 8'b00111111; //  368 :  63 - 0x3f
      11'h171: dout  = 8'b00111111; //  369 :  63 - 0x3f
      11'h172: dout  = 8'b00111111; //  370 :  63 - 0x3f
      11'h173: dout  = 8'b00111111; //  371 :  63 - 0x3f
      11'h174: dout  = 8'b00111111; //  372 :  63 - 0x3f
      11'h175: dout  = 8'b00111111; //  373 :  63 - 0x3f
      11'h176: dout  = 8'b00111111; //  374 :  63 - 0x3f
      11'h177: dout  = 8'b00111111; //  375 :  63 - 0x3f
      11'h178: dout  = 8'b00111111; //  376 :  63 - 0x3f
      11'h179: dout  = 8'b00111111; //  377 :  63 - 0x3f
      11'h17A: dout  = 8'b00111111; //  378 :  63 - 0x3f
      11'h17B: dout  = 8'b00111111; //  379 :  63 - 0x3f
      11'h17C: dout  = 8'b00111111; //  380 :  63 - 0x3f
      11'h17D: dout  = 8'b00111111; //  381 :  63 - 0x3f
      11'h17E: dout  = 8'b00111111; //  382 :  63 - 0x3f
      11'h17F: dout  = 8'b00111111; //  383 :  63 - 0x3f
      11'h180: dout  = 8'b00111111; //  384 :  63 - 0x3f -- line 0xc
      11'h181: dout  = 8'b00111111; //  385 :  63 - 0x3f
      11'h182: dout  = 8'b00111111; //  386 :  63 - 0x3f
      11'h183: dout  = 8'b00111111; //  387 :  63 - 0x3f
      11'h184: dout  = 8'b00111111; //  388 :  63 - 0x3f
      11'h185: dout  = 8'b00111111; //  389 :  63 - 0x3f
      11'h186: dout  = 8'b00111111; //  390 :  63 - 0x3f
      11'h187: dout  = 8'b00111111; //  391 :  63 - 0x3f
      11'h188: dout  = 8'b00111111; //  392 :  63 - 0x3f
      11'h189: dout  = 8'b00111111; //  393 :  63 - 0x3f
      11'h18A: dout  = 8'b00111111; //  394 :  63 - 0x3f
      11'h18B: dout  = 8'b00111111; //  395 :  63 - 0x3f
      11'h18C: dout  = 8'b00111111; //  396 :  63 - 0x3f
      11'h18D: dout  = 8'b00111111; //  397 :  63 - 0x3f
      11'h18E: dout  = 8'b00111111; //  398 :  63 - 0x3f
      11'h18F: dout  = 8'b00111111; //  399 :  63 - 0x3f
      11'h190: dout  = 8'b00111111; //  400 :  63 - 0x3f
      11'h191: dout  = 8'b00111111; //  401 :  63 - 0x3f
      11'h192: dout  = 8'b00111111; //  402 :  63 - 0x3f
      11'h193: dout  = 8'b00111111; //  403 :  63 - 0x3f
      11'h194: dout  = 8'b00111111; //  404 :  63 - 0x3f
      11'h195: dout  = 8'b00111111; //  405 :  63 - 0x3f
      11'h196: dout  = 8'b00111111; //  406 :  63 - 0x3f
      11'h197: dout  = 8'b00111111; //  407 :  63 - 0x3f
      11'h198: dout  = 8'b00111111; //  408 :  63 - 0x3f
      11'h199: dout  = 8'b00111111; //  409 :  63 - 0x3f
      11'h19A: dout  = 8'b00111111; //  410 :  63 - 0x3f
      11'h19B: dout  = 8'b00111111; //  411 :  63 - 0x3f
      11'h19C: dout  = 8'b00111111; //  412 :  63 - 0x3f
      11'h19D: dout  = 8'b00111111; //  413 :  63 - 0x3f
      11'h19E: dout  = 8'b00111111; //  414 :  63 - 0x3f
      11'h19F: dout  = 8'b00111111; //  415 :  63 - 0x3f
      11'h1A0: dout  = 8'b00111111; //  416 :  63 - 0x3f -- line 0xd
      11'h1A1: dout  = 8'b00111111; //  417 :  63 - 0x3f
      11'h1A2: dout  = 8'b00111111; //  418 :  63 - 0x3f
      11'h1A3: dout  = 8'b00111111; //  419 :  63 - 0x3f
      11'h1A4: dout  = 8'b00111111; //  420 :  63 - 0x3f
      11'h1A5: dout  = 8'b00111111; //  421 :  63 - 0x3f
      11'h1A6: dout  = 8'b00111111; //  422 :  63 - 0x3f
      11'h1A7: dout  = 8'b00111111; //  423 :  63 - 0x3f
      11'h1A8: dout  = 8'b00111111; //  424 :  63 - 0x3f
      11'h1A9: dout  = 8'b00111111; //  425 :  63 - 0x3f
      11'h1AA: dout  = 8'b00111111; //  426 :  63 - 0x3f
      11'h1AB: dout  = 8'b00111111; //  427 :  63 - 0x3f
      11'h1AC: dout  = 8'b00111111; //  428 :  63 - 0x3f
      11'h1AD: dout  = 8'b00111111; //  429 :  63 - 0x3f
      11'h1AE: dout  = 8'b00111111; //  430 :  63 - 0x3f
      11'h1AF: dout  = 8'b00111111; //  431 :  63 - 0x3f
      11'h1B0: dout  = 8'b00111111; //  432 :  63 - 0x3f
      11'h1B1: dout  = 8'b00111111; //  433 :  63 - 0x3f
      11'h1B2: dout  = 8'b00111111; //  434 :  63 - 0x3f
      11'h1B3: dout  = 8'b00111111; //  435 :  63 - 0x3f
      11'h1B4: dout  = 8'b00111111; //  436 :  63 - 0x3f
      11'h1B5: dout  = 8'b00111111; //  437 :  63 - 0x3f
      11'h1B6: dout  = 8'b00111111; //  438 :  63 - 0x3f
      11'h1B7: dout  = 8'b00111111; //  439 :  63 - 0x3f
      11'h1B8: dout  = 8'b00111111; //  440 :  63 - 0x3f
      11'h1B9: dout  = 8'b00111111; //  441 :  63 - 0x3f
      11'h1BA: dout  = 8'b00111111; //  442 :  63 - 0x3f
      11'h1BB: dout  = 8'b00111111; //  443 :  63 - 0x3f
      11'h1BC: dout  = 8'b00111111; //  444 :  63 - 0x3f
      11'h1BD: dout  = 8'b00111111; //  445 :  63 - 0x3f
      11'h1BE: dout  = 8'b00111111; //  446 :  63 - 0x3f
      11'h1BF: dout  = 8'b00111111; //  447 :  63 - 0x3f
      11'h1C0: dout  = 8'b00111111; //  448 :  63 - 0x3f -- line 0xe
      11'h1C1: dout  = 8'b00111111; //  449 :  63 - 0x3f
      11'h1C2: dout  = 8'b00111111; //  450 :  63 - 0x3f
      11'h1C3: dout  = 8'b00111111; //  451 :  63 - 0x3f
      11'h1C4: dout  = 8'b00111111; //  452 :  63 - 0x3f
      11'h1C5: dout  = 8'b00111111; //  453 :  63 - 0x3f
      11'h1C6: dout  = 8'b00111111; //  454 :  63 - 0x3f
      11'h1C7: dout  = 8'b00111111; //  455 :  63 - 0x3f
      11'h1C8: dout  = 8'b00111111; //  456 :  63 - 0x3f
      11'h1C9: dout  = 8'b00111111; //  457 :  63 - 0x3f
      11'h1CA: dout  = 8'b00111111; //  458 :  63 - 0x3f
      11'h1CB: dout  = 8'b00111111; //  459 :  63 - 0x3f
      11'h1CC: dout  = 8'b00111111; //  460 :  63 - 0x3f
      11'h1CD: dout  = 8'b00111111; //  461 :  63 - 0x3f
      11'h1CE: dout  = 8'b00111111; //  462 :  63 - 0x3f
      11'h1CF: dout  = 8'b00111111; //  463 :  63 - 0x3f
      11'h1D0: dout  = 8'b00111111; //  464 :  63 - 0x3f
      11'h1D1: dout  = 8'b00111111; //  465 :  63 - 0x3f
      11'h1D2: dout  = 8'b00111111; //  466 :  63 - 0x3f
      11'h1D3: dout  = 8'b00111111; //  467 :  63 - 0x3f
      11'h1D4: dout  = 8'b00111111; //  468 :  63 - 0x3f
      11'h1D5: dout  = 8'b00111111; //  469 :  63 - 0x3f
      11'h1D6: dout  = 8'b00111111; //  470 :  63 - 0x3f
      11'h1D7: dout  = 8'b00111111; //  471 :  63 - 0x3f
      11'h1D8: dout  = 8'b00111111; //  472 :  63 - 0x3f
      11'h1D9: dout  = 8'b00111111; //  473 :  63 - 0x3f
      11'h1DA: dout  = 8'b00111111; //  474 :  63 - 0x3f
      11'h1DB: dout  = 8'b00111111; //  475 :  63 - 0x3f
      11'h1DC: dout  = 8'b00111111; //  476 :  63 - 0x3f
      11'h1DD: dout  = 8'b00111111; //  477 :  63 - 0x3f
      11'h1DE: dout  = 8'b00111111; //  478 :  63 - 0x3f
      11'h1DF: dout  = 8'b00111111; //  479 :  63 - 0x3f
      11'h1E0: dout  = 8'b00111111; //  480 :  63 - 0x3f -- line 0xf
      11'h1E1: dout  = 8'b00111111; //  481 :  63 - 0x3f
      11'h1E2: dout  = 8'b00111111; //  482 :  63 - 0x3f
      11'h1E3: dout  = 8'b00111111; //  483 :  63 - 0x3f
      11'h1E4: dout  = 8'b00111111; //  484 :  63 - 0x3f
      11'h1E5: dout  = 8'b00111111; //  485 :  63 - 0x3f
      11'h1E6: dout  = 8'b00111111; //  486 :  63 - 0x3f
      11'h1E7: dout  = 8'b00111111; //  487 :  63 - 0x3f
      11'h1E8: dout  = 8'b00111111; //  488 :  63 - 0x3f
      11'h1E9: dout  = 8'b00111111; //  489 :  63 - 0x3f
      11'h1EA: dout  = 8'b00111111; //  490 :  63 - 0x3f
      11'h1EB: dout  = 8'b00111111; //  491 :  63 - 0x3f
      11'h1EC: dout  = 8'b00111111; //  492 :  63 - 0x3f
      11'h1ED: dout  = 8'b00111111; //  493 :  63 - 0x3f
      11'h1EE: dout  = 8'b00111111; //  494 :  63 - 0x3f
      11'h1EF: dout  = 8'b00111111; //  495 :  63 - 0x3f
      11'h1F0: dout  = 8'b00111111; //  496 :  63 - 0x3f
      11'h1F1: dout  = 8'b00111111; //  497 :  63 - 0x3f
      11'h1F2: dout  = 8'b00111111; //  498 :  63 - 0x3f
      11'h1F3: dout  = 8'b00111111; //  499 :  63 - 0x3f
      11'h1F4: dout  = 8'b00111111; //  500 :  63 - 0x3f
      11'h1F5: dout  = 8'b00111111; //  501 :  63 - 0x3f
      11'h1F6: dout  = 8'b00111111; //  502 :  63 - 0x3f
      11'h1F7: dout  = 8'b00111111; //  503 :  63 - 0x3f
      11'h1F8: dout  = 8'b00111111; //  504 :  63 - 0x3f
      11'h1F9: dout  = 8'b00111111; //  505 :  63 - 0x3f
      11'h1FA: dout  = 8'b00111111; //  506 :  63 - 0x3f
      11'h1FB: dout  = 8'b00111111; //  507 :  63 - 0x3f
      11'h1FC: dout  = 8'b00111111; //  508 :  63 - 0x3f
      11'h1FD: dout  = 8'b00111111; //  509 :  63 - 0x3f
      11'h1FE: dout  = 8'b00111111; //  510 :  63 - 0x3f
      11'h1FF: dout  = 8'b00111111; //  511 :  63 - 0x3f
      11'h200: dout  = 8'b00111111; //  512 :  63 - 0x3f -- line 0x10
      11'h201: dout  = 8'b00111111; //  513 :  63 - 0x3f
      11'h202: dout  = 8'b00111111; //  514 :  63 - 0x3f
      11'h203: dout  = 8'b00111111; //  515 :  63 - 0x3f
      11'h204: dout  = 8'b00111111; //  516 :  63 - 0x3f
      11'h205: dout  = 8'b00111111; //  517 :  63 - 0x3f
      11'h206: dout  = 8'b00111111; //  518 :  63 - 0x3f
      11'h207: dout  = 8'b00111111; //  519 :  63 - 0x3f
      11'h208: dout  = 8'b00111111; //  520 :  63 - 0x3f
      11'h209: dout  = 8'b00111111; //  521 :  63 - 0x3f
      11'h20A: dout  = 8'b00111111; //  522 :  63 - 0x3f
      11'h20B: dout  = 8'b00111111; //  523 :  63 - 0x3f
      11'h20C: dout  = 8'b00111111; //  524 :  63 - 0x3f
      11'h20D: dout  = 8'b00111111; //  525 :  63 - 0x3f
      11'h20E: dout  = 8'b00111111; //  526 :  63 - 0x3f
      11'h20F: dout  = 8'b00111111; //  527 :  63 - 0x3f
      11'h210: dout  = 8'b00111111; //  528 :  63 - 0x3f
      11'h211: dout  = 8'b00111111; //  529 :  63 - 0x3f
      11'h212: dout  = 8'b00111111; //  530 :  63 - 0x3f
      11'h213: dout  = 8'b00111111; //  531 :  63 - 0x3f
      11'h214: dout  = 8'b00111111; //  532 :  63 - 0x3f
      11'h215: dout  = 8'b00111111; //  533 :  63 - 0x3f
      11'h216: dout  = 8'b00111111; //  534 :  63 - 0x3f
      11'h217: dout  = 8'b00111111; //  535 :  63 - 0x3f
      11'h218: dout  = 8'b00111111; //  536 :  63 - 0x3f
      11'h219: dout  = 8'b00111111; //  537 :  63 - 0x3f
      11'h21A: dout  = 8'b00111111; //  538 :  63 - 0x3f
      11'h21B: dout  = 8'b00111111; //  539 :  63 - 0x3f
      11'h21C: dout  = 8'b00111111; //  540 :  63 - 0x3f
      11'h21D: dout  = 8'b00111111; //  541 :  63 - 0x3f
      11'h21E: dout  = 8'b00111111; //  542 :  63 - 0x3f
      11'h21F: dout  = 8'b00111111; //  543 :  63 - 0x3f
      11'h220: dout  = 8'b00111111; //  544 :  63 - 0x3f -- line 0x11
      11'h221: dout  = 8'b00111111; //  545 :  63 - 0x3f
      11'h222: dout  = 8'b00111111; //  546 :  63 - 0x3f
      11'h223: dout  = 8'b00111111; //  547 :  63 - 0x3f
      11'h224: dout  = 8'b00111111; //  548 :  63 - 0x3f
      11'h225: dout  = 8'b00111111; //  549 :  63 - 0x3f
      11'h226: dout  = 8'b00111111; //  550 :  63 - 0x3f
      11'h227: dout  = 8'b00111111; //  551 :  63 - 0x3f
      11'h228: dout  = 8'b00111111; //  552 :  63 - 0x3f
      11'h229: dout  = 8'b00111111; //  553 :  63 - 0x3f
      11'h22A: dout  = 8'b00111111; //  554 :  63 - 0x3f
      11'h22B: dout  = 8'b00111111; //  555 :  63 - 0x3f
      11'h22C: dout  = 8'b00111111; //  556 :  63 - 0x3f
      11'h22D: dout  = 8'b00111111; //  557 :  63 - 0x3f
      11'h22E: dout  = 8'b00111111; //  558 :  63 - 0x3f
      11'h22F: dout  = 8'b00111111; //  559 :  63 - 0x3f
      11'h230: dout  = 8'b00111111; //  560 :  63 - 0x3f
      11'h231: dout  = 8'b00111111; //  561 :  63 - 0x3f
      11'h232: dout  = 8'b00111111; //  562 :  63 - 0x3f
      11'h233: dout  = 8'b00111111; //  563 :  63 - 0x3f
      11'h234: dout  = 8'b00111111; //  564 :  63 - 0x3f
      11'h235: dout  = 8'b00111111; //  565 :  63 - 0x3f
      11'h236: dout  = 8'b00111111; //  566 :  63 - 0x3f
      11'h237: dout  = 8'b00111111; //  567 :  63 - 0x3f
      11'h238: dout  = 8'b00111111; //  568 :  63 - 0x3f
      11'h239: dout  = 8'b00111111; //  569 :  63 - 0x3f
      11'h23A: dout  = 8'b00111111; //  570 :  63 - 0x3f
      11'h23B: dout  = 8'b00111111; //  571 :  63 - 0x3f
      11'h23C: dout  = 8'b00111111; //  572 :  63 - 0x3f
      11'h23D: dout  = 8'b00111111; //  573 :  63 - 0x3f
      11'h23E: dout  = 8'b00111111; //  574 :  63 - 0x3f
      11'h23F: dout  = 8'b00111111; //  575 :  63 - 0x3f
      11'h240: dout  = 8'b00111111; //  576 :  63 - 0x3f -- line 0x12
      11'h241: dout  = 8'b00111111; //  577 :  63 - 0x3f
      11'h242: dout  = 8'b00111111; //  578 :  63 - 0x3f
      11'h243: dout  = 8'b00111111; //  579 :  63 - 0x3f
      11'h244: dout  = 8'b00111111; //  580 :  63 - 0x3f
      11'h245: dout  = 8'b00111111; //  581 :  63 - 0x3f
      11'h246: dout  = 8'b00111111; //  582 :  63 - 0x3f
      11'h247: dout  = 8'b00111111; //  583 :  63 - 0x3f
      11'h248: dout  = 8'b00111111; //  584 :  63 - 0x3f
      11'h249: dout  = 8'b00111111; //  585 :  63 - 0x3f
      11'h24A: dout  = 8'b00111111; //  586 :  63 - 0x3f
      11'h24B: dout  = 8'b00111111; //  587 :  63 - 0x3f
      11'h24C: dout  = 8'b00111111; //  588 :  63 - 0x3f
      11'h24D: dout  = 8'b00111111; //  589 :  63 - 0x3f
      11'h24E: dout  = 8'b00111111; //  590 :  63 - 0x3f
      11'h24F: dout  = 8'b00111111; //  591 :  63 - 0x3f
      11'h250: dout  = 8'b00000000; //  592 :   0 - 0x0
      11'h251: dout  = 8'b00000010; //  593 :   2 - 0x2
      11'h252: dout  = 8'b00000000; //  594 :   0 - 0x0
      11'h253: dout  = 8'b00000010; //  595 :   2 - 0x2
      11'h254: dout  = 8'b00000000; //  596 :   0 - 0x0
      11'h255: dout  = 8'b00000010; //  597 :   2 - 0x2
      11'h256: dout  = 8'b00000100; //  598 :   4 - 0x4
      11'h257: dout  = 8'b00000110; //  599 :   6 - 0x6
      11'h258: dout  = 8'b00000000; //  600 :   0 - 0x0
      11'h259: dout  = 8'b00000010; //  601 :   2 - 0x2
      11'h25A: dout  = 8'b00000000; //  602 :   0 - 0x0
      11'h25B: dout  = 8'b00000010; //  603 :   2 - 0x2
      11'h25C: dout  = 8'b00000100; //  604 :   4 - 0x4
      11'h25D: dout  = 8'b00000110; //  605 :   6 - 0x6
      11'h25E: dout  = 8'b00000000; //  606 :   0 - 0x0
      11'h25F: dout  = 8'b00000010; //  607 :   2 - 0x2
      11'h260: dout  = 8'b00111111; //  608 :  63 - 0x3f -- line 0x13
      11'h261: dout  = 8'b00111111; //  609 :  63 - 0x3f
      11'h262: dout  = 8'b00111111; //  610 :  63 - 0x3f
      11'h263: dout  = 8'b00111111; //  611 :  63 - 0x3f
      11'h264: dout  = 8'b00111111; //  612 :  63 - 0x3f
      11'h265: dout  = 8'b00111111; //  613 :  63 - 0x3f
      11'h266: dout  = 8'b00111111; //  614 :  63 - 0x3f
      11'h267: dout  = 8'b00111111; //  615 :  63 - 0x3f
      11'h268: dout  = 8'b00111111; //  616 :  63 - 0x3f
      11'h269: dout  = 8'b00111111; //  617 :  63 - 0x3f
      11'h26A: dout  = 8'b00111111; //  618 :  63 - 0x3f
      11'h26B: dout  = 8'b00111111; //  619 :  63 - 0x3f
      11'h26C: dout  = 8'b00111111; //  620 :  63 - 0x3f
      11'h26D: dout  = 8'b00111111; //  621 :  63 - 0x3f
      11'h26E: dout  = 8'b00111111; //  622 :  63 - 0x3f
      11'h26F: dout  = 8'b00111111; //  623 :  63 - 0x3f
      11'h270: dout  = 8'b00000001; //  624 :   1 - 0x1
      11'h271: dout  = 8'b00000011; //  625 :   3 - 0x3
      11'h272: dout  = 8'b00000001; //  626 :   1 - 0x1
      11'h273: dout  = 8'b00000011; //  627 :   3 - 0x3
      11'h274: dout  = 8'b00000001; //  628 :   1 - 0x1
      11'h275: dout  = 8'b00000011; //  629 :   3 - 0x3
      11'h276: dout  = 8'b00000101; //  630 :   5 - 0x5
      11'h277: dout  = 8'b00000111; //  631 :   7 - 0x7
      11'h278: dout  = 8'b00000001; //  632 :   1 - 0x1
      11'h279: dout  = 8'b00000011; //  633 :   3 - 0x3
      11'h27A: dout  = 8'b00000001; //  634 :   1 - 0x1
      11'h27B: dout  = 8'b00000011; //  635 :   3 - 0x3
      11'h27C: dout  = 8'b00000101; //  636 :   5 - 0x5
      11'h27D: dout  = 8'b00000111; //  637 :   7 - 0x7
      11'h27E: dout  = 8'b00000001; //  638 :   1 - 0x1
      11'h27F: dout  = 8'b00000011; //  639 :   3 - 0x3
      11'h280: dout  = 8'b00111111; //  640 :  63 - 0x3f -- line 0x14
      11'h281: dout  = 8'b00111111; //  641 :  63 - 0x3f
      11'h282: dout  = 8'b00111111; //  642 :  63 - 0x3f
      11'h283: dout  = 8'b00111111; //  643 :  63 - 0x3f
      11'h284: dout  = 8'b00111111; //  644 :  63 - 0x3f
      11'h285: dout  = 8'b00111111; //  645 :  63 - 0x3f
      11'h286: dout  = 8'b00111111; //  646 :  63 - 0x3f
      11'h287: dout  = 8'b00111111; //  647 :  63 - 0x3f
      11'h288: dout  = 8'b00111111; //  648 :  63 - 0x3f
      11'h289: dout  = 8'b00111111; //  649 :  63 - 0x3f
      11'h28A: dout  = 8'b00111111; //  650 :  63 - 0x3f
      11'h28B: dout  = 8'b00111111; //  651 :  63 - 0x3f
      11'h28C: dout  = 8'b00111111; //  652 :  63 - 0x3f
      11'h28D: dout  = 8'b00111111; //  653 :  63 - 0x3f
      11'h28E: dout  = 8'b00111111; //  654 :  63 - 0x3f
      11'h28F: dout  = 8'b00111111; //  655 :  63 - 0x3f
      11'h290: dout  = 8'b00111111; //  656 :  63 - 0x3f
      11'h291: dout  = 8'b00111111; //  657 :  63 - 0x3f
      11'h292: dout  = 8'b00111111; //  658 :  63 - 0x3f
      11'h293: dout  = 8'b00111111; //  659 :  63 - 0x3f
      11'h294: dout  = 8'b00111111; //  660 :  63 - 0x3f
      11'h295: dout  = 8'b00111111; //  661 :  63 - 0x3f
      11'h296: dout  = 8'b00111111; //  662 :  63 - 0x3f
      11'h297: dout  = 8'b00111111; //  663 :  63 - 0x3f
      11'h298: dout  = 8'b00111111; //  664 :  63 - 0x3f
      11'h299: dout  = 8'b00111111; //  665 :  63 - 0x3f
      11'h29A: dout  = 8'b00111111; //  666 :  63 - 0x3f
      11'h29B: dout  = 8'b00111111; //  667 :  63 - 0x3f
      11'h29C: dout  = 8'b00111111; //  668 :  63 - 0x3f
      11'h29D: dout  = 8'b00111111; //  669 :  63 - 0x3f
      11'h29E: dout  = 8'b00111111; //  670 :  63 - 0x3f
      11'h29F: dout  = 8'b00111111; //  671 :  63 - 0x3f
      11'h2A0: dout  = 8'b00111111; //  672 :  63 - 0x3f -- line 0x15
      11'h2A1: dout  = 8'b00111111; //  673 :  63 - 0x3f
      11'h2A2: dout  = 8'b00111111; //  674 :  63 - 0x3f
      11'h2A3: dout  = 8'b00111111; //  675 :  63 - 0x3f
      11'h2A4: dout  = 8'b00111111; //  676 :  63 - 0x3f
      11'h2A5: dout  = 8'b00111111; //  677 :  63 - 0x3f
      11'h2A6: dout  = 8'b00111111; //  678 :  63 - 0x3f
      11'h2A7: dout  = 8'b00111111; //  679 :  63 - 0x3f
      11'h2A8: dout  = 8'b00111111; //  680 :  63 - 0x3f
      11'h2A9: dout  = 8'b00111111; //  681 :  63 - 0x3f
      11'h2AA: dout  = 8'b00111111; //  682 :  63 - 0x3f
      11'h2AB: dout  = 8'b00111111; //  683 :  63 - 0x3f
      11'h2AC: dout  = 8'b00111111; //  684 :  63 - 0x3f
      11'h2AD: dout  = 8'b00111111; //  685 :  63 - 0x3f
      11'h2AE: dout  = 8'b00111111; //  686 :  63 - 0x3f
      11'h2AF: dout  = 8'b00111111; //  687 :  63 - 0x3f
      11'h2B0: dout  = 8'b00111111; //  688 :  63 - 0x3f
      11'h2B1: dout  = 8'b00111111; //  689 :  63 - 0x3f
      11'h2B2: dout  = 8'b00111111; //  690 :  63 - 0x3f
      11'h2B3: dout  = 8'b00111111; //  691 :  63 - 0x3f
      11'h2B4: dout  = 8'b00111111; //  692 :  63 - 0x3f
      11'h2B5: dout  = 8'b00111111; //  693 :  63 - 0x3f
      11'h2B6: dout  = 8'b00111111; //  694 :  63 - 0x3f
      11'h2B7: dout  = 8'b00111111; //  695 :  63 - 0x3f
      11'h2B8: dout  = 8'b00111111; //  696 :  63 - 0x3f
      11'h2B9: dout  = 8'b00111111; //  697 :  63 - 0x3f
      11'h2BA: dout  = 8'b00111111; //  698 :  63 - 0x3f
      11'h2BB: dout  = 8'b00111111; //  699 :  63 - 0x3f
      11'h2BC: dout  = 8'b00111111; //  700 :  63 - 0x3f
      11'h2BD: dout  = 8'b00111111; //  701 :  63 - 0x3f
      11'h2BE: dout  = 8'b00111111; //  702 :  63 - 0x3f
      11'h2BF: dout  = 8'b00111111; //  703 :  63 - 0x3f
      11'h2C0: dout  = 8'b00111111; //  704 :  63 - 0x3f -- line 0x16
      11'h2C1: dout  = 8'b00111111; //  705 :  63 - 0x3f
      11'h2C2: dout  = 8'b00111111; //  706 :  63 - 0x3f
      11'h2C3: dout  = 8'b00111111; //  707 :  63 - 0x3f
      11'h2C4: dout  = 8'b00111111; //  708 :  63 - 0x3f
      11'h2C5: dout  = 8'b00111111; //  709 :  63 - 0x3f
      11'h2C6: dout  = 8'b00111111; //  710 :  63 - 0x3f
      11'h2C7: dout  = 8'b00111111; //  711 :  63 - 0x3f
      11'h2C8: dout  = 8'b00111111; //  712 :  63 - 0x3f
      11'h2C9: dout  = 8'b00111111; //  713 :  63 - 0x3f
      11'h2CA: dout  = 8'b00111111; //  714 :  63 - 0x3f
      11'h2CB: dout  = 8'b00111111; //  715 :  63 - 0x3f
      11'h2CC: dout  = 8'b00111111; //  716 :  63 - 0x3f
      11'h2CD: dout  = 8'b00111111; //  717 :  63 - 0x3f
      11'h2CE: dout  = 8'b00111111; //  718 :  63 - 0x3f
      11'h2CF: dout  = 8'b00111111; //  719 :  63 - 0x3f
      11'h2D0: dout  = 8'b00111111; //  720 :  63 - 0x3f
      11'h2D1: dout  = 8'b00111111; //  721 :  63 - 0x3f
      11'h2D2: dout  = 8'b00111111; //  722 :  63 - 0x3f
      11'h2D3: dout  = 8'b00111111; //  723 :  63 - 0x3f
      11'h2D4: dout  = 8'b00111111; //  724 :  63 - 0x3f
      11'h2D5: dout  = 8'b00111111; //  725 :  63 - 0x3f
      11'h2D6: dout  = 8'b00111111; //  726 :  63 - 0x3f
      11'h2D7: dout  = 8'b00111111; //  727 :  63 - 0x3f
      11'h2D8: dout  = 8'b00111111; //  728 :  63 - 0x3f
      11'h2D9: dout  = 8'b00111111; //  729 :  63 - 0x3f
      11'h2DA: dout  = 8'b00111111; //  730 :  63 - 0x3f
      11'h2DB: dout  = 8'b00111111; //  731 :  63 - 0x3f
      11'h2DC: dout  = 8'b00111111; //  732 :  63 - 0x3f
      11'h2DD: dout  = 8'b00111111; //  733 :  63 - 0x3f
      11'h2DE: dout  = 8'b00111111; //  734 :  63 - 0x3f
      11'h2DF: dout  = 8'b00111111; //  735 :  63 - 0x3f
      11'h2E0: dout  = 8'b00111111; //  736 :  63 - 0x3f -- line 0x17
      11'h2E1: dout  = 8'b00111111; //  737 :  63 - 0x3f
      11'h2E2: dout  = 8'b00111111; //  738 :  63 - 0x3f
      11'h2E3: dout  = 8'b00111111; //  739 :  63 - 0x3f
      11'h2E4: dout  = 8'b00111111; //  740 :  63 - 0x3f
      11'h2E5: dout  = 8'b00111111; //  741 :  63 - 0x3f
      11'h2E6: dout  = 8'b00111111; //  742 :  63 - 0x3f
      11'h2E7: dout  = 8'b00111111; //  743 :  63 - 0x3f
      11'h2E8: dout  = 8'b00111111; //  744 :  63 - 0x3f
      11'h2E9: dout  = 8'b00111111; //  745 :  63 - 0x3f
      11'h2EA: dout  = 8'b00111111; //  746 :  63 - 0x3f
      11'h2EB: dout  = 8'b00111111; //  747 :  63 - 0x3f
      11'h2EC: dout  = 8'b00111111; //  748 :  63 - 0x3f
      11'h2ED: dout  = 8'b00111111; //  749 :  63 - 0x3f
      11'h2EE: dout  = 8'b00111111; //  750 :  63 - 0x3f
      11'h2EF: dout  = 8'b00111111; //  751 :  63 - 0x3f
      11'h2F0: dout  = 8'b11000101; //  752 : 197 - 0xc5
      11'h2F1: dout  = 8'b11010110; //  753 : 214 - 0xd6
      11'h2F2: dout  = 8'b11000101; //  754 : 197 - 0xc5
      11'h2F3: dout  = 8'b11010110; //  755 : 214 - 0xd6
      11'h2F4: dout  = 8'b11000101; //  756 : 197 - 0xc5
      11'h2F5: dout  = 8'b11010110; //  757 : 214 - 0xd6
      11'h2F6: dout  = 8'b11000101; //  758 : 197 - 0xc5
      11'h2F7: dout  = 8'b11010110; //  759 : 214 - 0xd6
      11'h2F8: dout  = 8'b11000101; //  760 : 197 - 0xc5
      11'h2F9: dout  = 8'b11010110; //  761 : 214 - 0xd6
      11'h2FA: dout  = 8'b11000101; //  762 : 197 - 0xc5
      11'h2FB: dout  = 8'b11010110; //  763 : 214 - 0xd6
      11'h2FC: dout  = 8'b11000101; //  764 : 197 - 0xc5
      11'h2FD: dout  = 8'b11010110; //  765 : 214 - 0xd6
      11'h2FE: dout  = 8'b11000101; //  766 : 197 - 0xc5
      11'h2FF: dout  = 8'b11010110; //  767 : 214 - 0xd6
      11'h300: dout  = 8'b00111111; //  768 :  63 - 0x3f -- line 0x18
      11'h301: dout  = 8'b00111111; //  769 :  63 - 0x3f
      11'h302: dout  = 8'b00111111; //  770 :  63 - 0x3f
      11'h303: dout  = 8'b00111111; //  771 :  63 - 0x3f
      11'h304: dout  = 8'b00011100; //  772 :  28 - 0x1c
      11'h305: dout  = 8'b00011110; //  773 :  30 - 0x1e
      11'h306: dout  = 8'b00111111; //  774 :  63 - 0x3f
      11'h307: dout  = 8'b00111111; //  775 :  63 - 0x3f
      11'h308: dout  = 8'b00111111; //  776 :  63 - 0x3f
      11'h309: dout  = 8'b00111111; //  777 :  63 - 0x3f
      11'h30A: dout  = 8'b00111111; //  778 :  63 - 0x3f
      11'h30B: dout  = 8'b00111111; //  779 :  63 - 0x3f
      11'h30C: dout  = 8'b00111111; //  780 :  63 - 0x3f
      11'h30D: dout  = 8'b00111111; //  781 :  63 - 0x3f
      11'h30E: dout  = 8'b00111111; //  782 :  63 - 0x3f
      11'h30F: dout  = 8'b00111111; //  783 :  63 - 0x3f
      11'h310: dout  = 8'b11000111; //  784 : 199 - 0xc7
      11'h311: dout  = 8'b11001001; //  785 : 201 - 0xc9
      11'h312: dout  = 8'b11000111; //  786 : 199 - 0xc7
      11'h313: dout  = 8'b11001001; //  787 : 201 - 0xc9
      11'h314: dout  = 8'b11000111; //  788 : 199 - 0xc7
      11'h315: dout  = 8'b11001001; //  789 : 201 - 0xc9
      11'h316: dout  = 8'b11000111; //  790 : 199 - 0xc7
      11'h317: dout  = 8'b11001001; //  791 : 201 - 0xc9
      11'h318: dout  = 8'b11000111; //  792 : 199 - 0xc7
      11'h319: dout  = 8'b11001001; //  793 : 201 - 0xc9
      11'h31A: dout  = 8'b11000111; //  794 : 199 - 0xc7
      11'h31B: dout  = 8'b11001001; //  795 : 201 - 0xc9
      11'h31C: dout  = 8'b11000111; //  796 : 199 - 0xc7
      11'h31D: dout  = 8'b11001001; //  797 : 201 - 0xc9
      11'h31E: dout  = 8'b11000111; //  798 : 199 - 0xc7
      11'h31F: dout  = 8'b11001001; //  799 : 201 - 0xc9
      11'h320: dout  = 8'b00111111; //  800 :  63 - 0x3f -- line 0x19
      11'h321: dout  = 8'b00111111; //  801 :  63 - 0x3f
      11'h322: dout  = 8'b00111111; //  802 :  63 - 0x3f
      11'h323: dout  = 8'b00111111; //  803 :  63 - 0x3f
      11'h324: dout  = 8'b00011101; //  804 :  29 - 0x1d
      11'h325: dout  = 8'b00011111; //  805 :  31 - 0x1f
      11'h326: dout  = 8'b00111111; //  806 :  63 - 0x3f
      11'h327: dout  = 8'b00111111; //  807 :  63 - 0x3f
      11'h328: dout  = 8'b00111111; //  808 :  63 - 0x3f
      11'h329: dout  = 8'b00111111; //  809 :  63 - 0x3f
      11'h32A: dout  = 8'b00111111; //  810 :  63 - 0x3f
      11'h32B: dout  = 8'b00111111; //  811 :  63 - 0x3f
      11'h32C: dout  = 8'b00111111; //  812 :  63 - 0x3f
      11'h32D: dout  = 8'b00111111; //  813 :  63 - 0x3f
      11'h32E: dout  = 8'b00111111; //  814 :  63 - 0x3f
      11'h32F: dout  = 8'b00111111; //  815 :  63 - 0x3f
      11'h330: dout  = 8'b11010111; //  816 : 215 - 0xd7
      11'h331: dout  = 8'b11011001; //  817 : 217 - 0xd9
      11'h332: dout  = 8'b11010111; //  818 : 215 - 0xd7
      11'h333: dout  = 8'b11011001; //  819 : 217 - 0xd9
      11'h334: dout  = 8'b11010111; //  820 : 215 - 0xd7
      11'h335: dout  = 8'b11011001; //  821 : 217 - 0xd9
      11'h336: dout  = 8'b11010111; //  822 : 215 - 0xd7
      11'h337: dout  = 8'b11011001; //  823 : 217 - 0xd9
      11'h338: dout  = 8'b11010111; //  824 : 215 - 0xd7
      11'h339: dout  = 8'b11011001; //  825 : 217 - 0xd9
      11'h33A: dout  = 8'b11010111; //  826 : 215 - 0xd7
      11'h33B: dout  = 8'b11011001; //  827 : 217 - 0xd9
      11'h33C: dout  = 8'b11010111; //  828 : 215 - 0xd7
      11'h33D: dout  = 8'b11011001; //  829 : 217 - 0xd9
      11'h33E: dout  = 8'b11010111; //  830 : 215 - 0xd7
      11'h33F: dout  = 8'b11011001; //  831 : 217 - 0xd9
      11'h340: dout  = 8'b01110000; //  832 : 112 - 0x70 -- line 0x1a
      11'h341: dout  = 8'b01110001; //  833 : 113 - 0x71
      11'h342: dout  = 8'b01110001; //  834 : 113 - 0x71
      11'h343: dout  = 8'b01110001; //  835 : 113 - 0x71
      11'h344: dout  = 8'b01110001; //  836 : 113 - 0x71
      11'h345: dout  = 8'b01110001; //  837 : 113 - 0x71
      11'h346: dout  = 8'b01110001; //  838 : 113 - 0x71
      11'h347: dout  = 8'b01110001; //  839 : 113 - 0x71
      11'h348: dout  = 8'b01110001; //  840 : 113 - 0x71
      11'h349: dout  = 8'b01110001; //  841 : 113 - 0x71
      11'h34A: dout  = 8'b01110001; //  842 : 113 - 0x71
      11'h34B: dout  = 8'b01110001; //  843 : 113 - 0x71
      11'h34C: dout  = 8'b01110001; //  844 : 113 - 0x71
      11'h34D: dout  = 8'b01110001; //  845 : 113 - 0x71
      11'h34E: dout  = 8'b01110001; //  846 : 113 - 0x71
      11'h34F: dout  = 8'b01110001; //  847 : 113 - 0x71
      11'h350: dout  = 8'b01110001; //  848 : 113 - 0x71
      11'h351: dout  = 8'b01110001; //  849 : 113 - 0x71
      11'h352: dout  = 8'b01110001; //  850 : 113 - 0x71
      11'h353: dout  = 8'b01110001; //  851 : 113 - 0x71
      11'h354: dout  = 8'b01110001; //  852 : 113 - 0x71
      11'h355: dout  = 8'b01110001; //  853 : 113 - 0x71
      11'h356: dout  = 8'b01110001; //  854 : 113 - 0x71
      11'h357: dout  = 8'b01110001; //  855 : 113 - 0x71
      11'h358: dout  = 8'b01110001; //  856 : 113 - 0x71
      11'h359: dout  = 8'b01110001; //  857 : 113 - 0x71
      11'h35A: dout  = 8'b01110001; //  858 : 113 - 0x71
      11'h35B: dout  = 8'b01110001; //  859 : 113 - 0x71
      11'h35C: dout  = 8'b01110001; //  860 : 113 - 0x71
      11'h35D: dout  = 8'b01110001; //  861 : 113 - 0x71
      11'h35E: dout  = 8'b01110001; //  862 : 113 - 0x71
      11'h35F: dout  = 8'b01110001; //  863 : 113 - 0x71
      11'h360: dout  = 8'b01100000; //  864 :  96 - 0x60 -- line 0x1b
      11'h361: dout  = 8'b01110111; //  865 : 119 - 0x77
      11'h362: dout  = 8'b01110111; //  866 : 119 - 0x77
      11'h363: dout  = 8'b01110111; //  867 : 119 - 0x77
      11'h364: dout  = 8'b01110111; //  868 : 119 - 0x77
      11'h365: dout  = 8'b01110111; //  869 : 119 - 0x77
      11'h366: dout  = 8'b01110111; //  870 : 119 - 0x77
      11'h367: dout  = 8'b01110111; //  871 : 119 - 0x77
      11'h368: dout  = 8'b01110111; //  872 : 119 - 0x77
      11'h369: dout  = 8'b01110111; //  873 : 119 - 0x77
      11'h36A: dout  = 8'b01110111; //  874 : 119 - 0x77
      11'h36B: dout  = 8'b01110111; //  875 : 119 - 0x77
      11'h36C: dout  = 8'b01110111; //  876 : 119 - 0x77
      11'h36D: dout  = 8'b01110111; //  877 : 119 - 0x77
      11'h36E: dout  = 8'b01110111; //  878 : 119 - 0x77
      11'h36F: dout  = 8'b01110111; //  879 : 119 - 0x77
      11'h370: dout  = 8'b01110111; //  880 : 119 - 0x77
      11'h371: dout  = 8'b01110111; //  881 : 119 - 0x77
      11'h372: dout  = 8'b01110111; //  882 : 119 - 0x77
      11'h373: dout  = 8'b01110111; //  883 : 119 - 0x77
      11'h374: dout  = 8'b01110111; //  884 : 119 - 0x77
      11'h375: dout  = 8'b01110111; //  885 : 119 - 0x77
      11'h376: dout  = 8'b01110111; //  886 : 119 - 0x77
      11'h377: dout  = 8'b01110111; //  887 : 119 - 0x77
      11'h378: dout  = 8'b01110111; //  888 : 119 - 0x77
      11'h379: dout  = 8'b01110111; //  889 : 119 - 0x77
      11'h37A: dout  = 8'b01110111; //  890 : 119 - 0x77
      11'h37B: dout  = 8'b01110111; //  891 : 119 - 0x77
      11'h37C: dout  = 8'b01110111; //  892 : 119 - 0x77
      11'h37D: dout  = 8'b01110111; //  893 : 119 - 0x77
      11'h37E: dout  = 8'b01110111; //  894 : 119 - 0x77
      11'h37F: dout  = 8'b01110111; //  895 : 119 - 0x77
      11'h380: dout  = 8'b01100000; //  896 :  96 - 0x60 -- line 0x1c
      11'h381: dout  = 8'b01110011; //  897 : 115 - 0x73
      11'h382: dout  = 8'b01110011; //  898 : 115 - 0x73
      11'h383: dout  = 8'b01110011; //  899 : 115 - 0x73
      11'h384: dout  = 8'b01110011; //  900 : 115 - 0x73
      11'h385: dout  = 8'b01110011; //  901 : 115 - 0x73
      11'h386: dout  = 8'b01110011; //  902 : 115 - 0x73
      11'h387: dout  = 8'b01110011; //  903 : 115 - 0x73
      11'h388: dout  = 8'b01110011; //  904 : 115 - 0x73
      11'h389: dout  = 8'b01110011; //  905 : 115 - 0x73
      11'h38A: dout  = 8'b01110011; //  906 : 115 - 0x73
      11'h38B: dout  = 8'b01110011; //  907 : 115 - 0x73
      11'h38C: dout  = 8'b01110011; //  908 : 115 - 0x73
      11'h38D: dout  = 8'b01110011; //  909 : 115 - 0x73
      11'h38E: dout  = 8'b01110011; //  910 : 115 - 0x73
      11'h38F: dout  = 8'b01110011; //  911 : 115 - 0x73
      11'h390: dout  = 8'b01110011; //  912 : 115 - 0x73
      11'h391: dout  = 8'b01110011; //  913 : 115 - 0x73
      11'h392: dout  = 8'b01110011; //  914 : 115 - 0x73
      11'h393: dout  = 8'b01110011; //  915 : 115 - 0x73
      11'h394: dout  = 8'b01110011; //  916 : 115 - 0x73
      11'h395: dout  = 8'b01110011; //  917 : 115 - 0x73
      11'h396: dout  = 8'b01110011; //  918 : 115 - 0x73
      11'h397: dout  = 8'b01110011; //  919 : 115 - 0x73
      11'h398: dout  = 8'b01110011; //  920 : 115 - 0x73
      11'h399: dout  = 8'b01110011; //  921 : 115 - 0x73
      11'h39A: dout  = 8'b01110011; //  922 : 115 - 0x73
      11'h39B: dout  = 8'b01110011; //  923 : 115 - 0x73
      11'h39C: dout  = 8'b01110011; //  924 : 115 - 0x73
      11'h39D: dout  = 8'b01110011; //  925 : 115 - 0x73
      11'h39E: dout  = 8'b01110011; //  926 : 115 - 0x73
      11'h39F: dout  = 8'b01110011; //  927 : 115 - 0x73
      11'h3A0: dout  = 8'b01100000; //  928 :  96 - 0x60 -- line 0x1d
      11'h3A1: dout  = 8'b01110011; //  929 : 115 - 0x73
      11'h3A2: dout  = 8'b01110011; //  930 : 115 - 0x73
      11'h3A3: dout  = 8'b01110011; //  931 : 115 - 0x73
      11'h3A4: dout  = 8'b01110011; //  932 : 115 - 0x73
      11'h3A5: dout  = 8'b01110011; //  933 : 115 - 0x73
      11'h3A6: dout  = 8'b01110011; //  934 : 115 - 0x73
      11'h3A7: dout  = 8'b01110011; //  935 : 115 - 0x73
      11'h3A8: dout  = 8'b01110011; //  936 : 115 - 0x73
      11'h3A9: dout  = 8'b01110011; //  937 : 115 - 0x73
      11'h3AA: dout  = 8'b01110011; //  938 : 115 - 0x73
      11'h3AB: dout  = 8'b01110011; //  939 : 115 - 0x73
      11'h3AC: dout  = 8'b01110011; //  940 : 115 - 0x73
      11'h3AD: dout  = 8'b01110011; //  941 : 115 - 0x73
      11'h3AE: dout  = 8'b01110011; //  942 : 115 - 0x73
      11'h3AF: dout  = 8'b01110011; //  943 : 115 - 0x73
      11'h3B0: dout  = 8'b01110011; //  944 : 115 - 0x73
      11'h3B1: dout  = 8'b01110011; //  945 : 115 - 0x73
      11'h3B2: dout  = 8'b01110011; //  946 : 115 - 0x73
      11'h3B3: dout  = 8'b01110011; //  947 : 115 - 0x73
      11'h3B4: dout  = 8'b01110011; //  948 : 115 - 0x73
      11'h3B5: dout  = 8'b01110011; //  949 : 115 - 0x73
      11'h3B6: dout  = 8'b01110011; //  950 : 115 - 0x73
      11'h3B7: dout  = 8'b01110011; //  951 : 115 - 0x73
      11'h3B8: dout  = 8'b01110011; //  952 : 115 - 0x73
      11'h3B9: dout  = 8'b01110011; //  953 : 115 - 0x73
      11'h3BA: dout  = 8'b01110011; //  954 : 115 - 0x73
      11'h3BB: dout  = 8'b01110011; //  955 : 115 - 0x73
      11'h3BC: dout  = 8'b01110011; //  956 : 115 - 0x73
      11'h3BD: dout  = 8'b01110011; //  957 : 115 - 0x73
      11'h3BE: dout  = 8'b01110011; //  958 : 115 - 0x73
      11'h3BF: dout  = 8'b01110011; //  959 : 115 - 0x73
        //-- Attribute Table 0----
      11'h3C0: dout  = 8'b00000000; //  960 :   0 - 0x0
      11'h3C1: dout  = 8'b00000000; //  961 :   0 - 0x0
      11'h3C2: dout  = 8'b00000000; //  962 :   0 - 0x0
      11'h3C3: dout  = 8'b00000000; //  963 :   0 - 0x0
      11'h3C4: dout  = 8'b00000000; //  964 :   0 - 0x0
      11'h3C5: dout  = 8'b00000000; //  965 :   0 - 0x0
      11'h3C6: dout  = 8'b00000000; //  966 :   0 - 0x0
      11'h3C7: dout  = 8'b00000000; //  967 :   0 - 0x0
      11'h3C8: dout  = 8'b00000000; //  968 :   0 - 0x0
      11'h3C9: dout  = 8'b00000000; //  969 :   0 - 0x0
      11'h3CA: dout  = 8'b00000000; //  970 :   0 - 0x0
      11'h3CB: dout  = 8'b00000000; //  971 :   0 - 0x0
      11'h3CC: dout  = 8'b00000000; //  972 :   0 - 0x0
      11'h3CD: dout  = 8'b00000000; //  973 :   0 - 0x0
      11'h3CE: dout  = 8'b00001000; //  974 :   8 - 0x8
      11'h3CF: dout  = 8'b00001000; //  975 :   8 - 0x8
      11'h3D0: dout  = 8'b00000000; //  976 :   0 - 0x0
      11'h3D1: dout  = 8'b00000000; //  977 :   0 - 0x0
      11'h3D2: dout  = 8'b00000000; //  978 :   0 - 0x0
      11'h3D3: dout  = 8'b00000000; //  979 :   0 - 0x0
      11'h3D4: dout  = 8'b00000000; //  980 :   0 - 0x0
      11'h3D5: dout  = 8'b01010001; //  981 :  81 - 0x51
      11'h3D6: dout  = 8'b01010000; //  982 :  80 - 0x50
      11'h3D7: dout  = 8'b01010000; //  983 :  80 - 0x50
      11'h3D8: dout  = 8'b00000000; //  984 :   0 - 0x0
      11'h3D9: dout  = 8'b00000000; //  985 :   0 - 0x0
      11'h3DA: dout  = 8'b00000000; //  986 :   0 - 0x0
      11'h3DB: dout  = 8'b00000000; //  987 :   0 - 0x0
      11'h3DC: dout  = 8'b00000000; //  988 :   0 - 0x0
      11'h3DD: dout  = 8'b00000000; //  989 :   0 - 0x0
      11'h3DE: dout  = 8'b00000000; //  990 :   0 - 0x0
      11'h3DF: dout  = 8'b00000000; //  991 :   0 - 0x0
      11'h3E0: dout  = 8'b00000000; //  992 :   0 - 0x0
      11'h3E1: dout  = 8'b00000000; //  993 :   0 - 0x0
      11'h3E2: dout  = 8'b00000000; //  994 :   0 - 0x0
      11'h3E3: dout  = 8'b00000000; //  995 :   0 - 0x0
      11'h3E4: dout  = 8'b10100000; //  996 : 160 - 0xa0
      11'h3E5: dout  = 8'b10100000; //  997 : 160 - 0xa0
      11'h3E6: dout  = 8'b10100000; //  998 : 160 - 0xa0
      11'h3E7: dout  = 8'b10100000; //  999 : 160 - 0xa0
      11'h3E8: dout  = 8'b00000000; // 1000 :   0 - 0x0
      11'h3E9: dout  = 8'b00000000; // 1001 :   0 - 0x0
      11'h3EA: dout  = 8'b00000000; // 1002 :   0 - 0x0
      11'h3EB: dout  = 8'b00000000; // 1003 :   0 - 0x0
      11'h3EC: dout  = 8'b00000000; // 1004 :   0 - 0x0
      11'h3ED: dout  = 8'b00000000; // 1005 :   0 - 0x0
      11'h3EE: dout  = 8'b00000000; // 1006 :   0 - 0x0
      11'h3EF: dout  = 8'b00000000; // 1007 :   0 - 0x0
      11'h3F0: dout  = 8'b00000000; // 1008 :   0 - 0x0
      11'h3F1: dout  = 8'b00000010; // 1009 :   2 - 0x2
      11'h3F2: dout  = 8'b00000000; // 1010 :   0 - 0x0
      11'h3F3: dout  = 8'b00000000; // 1011 :   0 - 0x0
      11'h3F4: dout  = 8'b00000000; // 1012 :   0 - 0x0
      11'h3F5: dout  = 8'b00000000; // 1013 :   0 - 0x0
      11'h3F6: dout  = 8'b00000000; // 1014 :   0 - 0x0
      11'h3F7: dout  = 8'b00000000; // 1015 :   0 - 0x0
      11'h3F8: dout  = 8'b00000000; // 1016 :   0 - 0x0
      11'h3F9: dout  = 8'b00000000; // 1017 :   0 - 0x0
      11'h3FA: dout  = 8'b00000000; // 1018 :   0 - 0x0
      11'h3FB: dout  = 8'b00000000; // 1019 :   0 - 0x0
      11'h3FC: dout  = 8'b00000000; // 1020 :   0 - 0x0
      11'h3FD: dout  = 8'b00000000; // 1021 :   0 - 0x0
      11'h3FE: dout  = 8'b00000000; // 1022 :   0 - 0x0
      11'h3FF: dout  = 8'b00000000; // 1023 :   0 - 0x0
     //----- Name Table 1---------
      11'h400: dout  = 8'b01110001; // 1024 : 113 - 0x71 -- line 0x0
      11'h401: dout  = 8'b01110001; // 1025 : 113 - 0x71
      11'h402: dout  = 8'b01110001; // 1026 : 113 - 0x71
      11'h403: dout  = 8'b01110001; // 1027 : 113 - 0x71
      11'h404: dout  = 8'b01110001; // 1028 : 113 - 0x71
      11'h405: dout  = 8'b01110001; // 1029 : 113 - 0x71
      11'h406: dout  = 8'b01110001; // 1030 : 113 - 0x71
      11'h407: dout  = 8'b01110001; // 1031 : 113 - 0x71
      11'h408: dout  = 8'b01110001; // 1032 : 113 - 0x71
      11'h409: dout  = 8'b01110010; // 1033 : 114 - 0x72
      11'h40A: dout  = 8'b00010000; // 1034 :  16 - 0x10
      11'h40B: dout  = 8'b00010001; // 1035 :  17 - 0x11
      11'h40C: dout  = 8'b00001100; // 1036 :  12 - 0xc
      11'h40D: dout  = 8'b00001110; // 1037 :  14 - 0xe
      11'h40E: dout  = 8'b00110000; // 1038 :  48 - 0x30
      11'h40F: dout  = 8'b00111111; // 1039 :  63 - 0x3f
      11'h410: dout  = 8'b00110000; // 1040 :  48 - 0x30
      11'h411: dout  = 8'b00111111; // 1041 :  63 - 0x3f
      11'h412: dout  = 8'b00110000; // 1042 :  48 - 0x30
      11'h413: dout  = 8'b00111111; // 1043 :  63 - 0x3f
      11'h414: dout  = 8'b00110000; // 1044 :  48 - 0x30
      11'h415: dout  = 8'b00111111; // 1045 :  63 - 0x3f
      11'h416: dout  = 8'b00110000; // 1046 :  48 - 0x30
      11'h417: dout  = 8'b00111111; // 1047 :  63 - 0x3f
      11'h418: dout  = 8'b00110000; // 1048 :  48 - 0x30
      11'h419: dout  = 8'b00111111; // 1049 :  63 - 0x3f
      11'h41A: dout  = 8'b00110000; // 1050 :  48 - 0x30
      11'h41B: dout  = 8'b00111111; // 1051 :  63 - 0x3f
      11'h41C: dout  = 8'b00110000; // 1052 :  48 - 0x30
      11'h41D: dout  = 8'b00111111; // 1053 :  63 - 0x3f
      11'h41E: dout  = 8'b00110000; // 1054 :  48 - 0x30
      11'h41F: dout  = 8'b00111111; // 1055 :  63 - 0x3f
      11'h420: dout  = 8'b01110111; // 1056 : 119 - 0x77 -- line 0x1
      11'h421: dout  = 8'b01110111; // 1057 : 119 - 0x77
      11'h422: dout  = 8'b01110111; // 1058 : 119 - 0x77
      11'h423: dout  = 8'b01110111; // 1059 : 119 - 0x77
      11'h424: dout  = 8'b01110111; // 1060 : 119 - 0x77
      11'h425: dout  = 8'b01110111; // 1061 : 119 - 0x77
      11'h426: dout  = 8'b01110111; // 1062 : 119 - 0x77
      11'h427: dout  = 8'b01110111; // 1063 : 119 - 0x77
      11'h428: dout  = 8'b01110111; // 1064 : 119 - 0x77
      11'h429: dout  = 8'b01100001; // 1065 :  97 - 0x61
      11'h42A: dout  = 8'b00010000; // 1066 :  16 - 0x10
      11'h42B: dout  = 8'b00010001; // 1067 :  17 - 0x11
      11'h42C: dout  = 8'b00001101; // 1068 :  13 - 0xd
      11'h42D: dout  = 8'b00001111; // 1069 :  15 - 0xf
      11'h42E: dout  = 8'b00111111; // 1070 :  63 - 0x3f
      11'h42F: dout  = 8'b00110000; // 1071 :  48 - 0x30
      11'h430: dout  = 8'b00111111; // 1072 :  63 - 0x3f
      11'h431: dout  = 8'b00110000; // 1073 :  48 - 0x30
      11'h432: dout  = 8'b00111111; // 1074 :  63 - 0x3f
      11'h433: dout  = 8'b00110000; // 1075 :  48 - 0x30
      11'h434: dout  = 8'b00111111; // 1076 :  63 - 0x3f
      11'h435: dout  = 8'b00110000; // 1077 :  48 - 0x30
      11'h436: dout  = 8'b00111111; // 1078 :  63 - 0x3f
      11'h437: dout  = 8'b00110000; // 1079 :  48 - 0x30
      11'h438: dout  = 8'b00111111; // 1080 :  63 - 0x3f
      11'h439: dout  = 8'b00110000; // 1081 :  48 - 0x30
      11'h43A: dout  = 8'b00111111; // 1082 :  63 - 0x3f
      11'h43B: dout  = 8'b00110000; // 1083 :  48 - 0x30
      11'h43C: dout  = 8'b00111111; // 1084 :  63 - 0x3f
      11'h43D: dout  = 8'b00110000; // 1085 :  48 - 0x30
      11'h43E: dout  = 8'b00111111; // 1086 :  63 - 0x3f
      11'h43F: dout  = 8'b00110000; // 1087 :  48 - 0x30
      11'h440: dout  = 8'b00111001; // 1088 :  57 - 0x39 -- line 0x2
      11'h441: dout  = 8'b00111001; // 1089 :  57 - 0x39
      11'h442: dout  = 8'b00111001; // 1090 :  57 - 0x39
      11'h443: dout  = 8'b00111001; // 1091 :  57 - 0x39
      11'h444: dout  = 8'b00111001; // 1092 :  57 - 0x39
      11'h445: dout  = 8'b00111001; // 1093 :  57 - 0x39
      11'h446: dout  = 8'b00111001; // 1094 :  57 - 0x39
      11'h447: dout  = 8'b00111001; // 1095 :  57 - 0x39
      11'h448: dout  = 8'b00111001; // 1096 :  57 - 0x39
      11'h449: dout  = 8'b00111001; // 1097 :  57 - 0x39
      11'h44A: dout  = 8'b00010000; // 1098 :  16 - 0x10
      11'h44B: dout  = 8'b00010001; // 1099 :  17 - 0x11
      11'h44C: dout  = 8'b00001100; // 1100 :  12 - 0xc
      11'h44D: dout  = 8'b00001110; // 1101 :  14 - 0xe
      11'h44E: dout  = 8'b00110000; // 1102 :  48 - 0x30
      11'h44F: dout  = 8'b00111111; // 1103 :  63 - 0x3f
      11'h450: dout  = 8'b00110000; // 1104 :  48 - 0x30
      11'h451: dout  = 8'b00111111; // 1105 :  63 - 0x3f
      11'h452: dout  = 8'b00110000; // 1106 :  48 - 0x30
      11'h453: dout  = 8'b00111111; // 1107 :  63 - 0x3f
      11'h454: dout  = 8'b00110000; // 1108 :  48 - 0x30
      11'h455: dout  = 8'b00111111; // 1109 :  63 - 0x3f
      11'h456: dout  = 8'b00110000; // 1110 :  48 - 0x30
      11'h457: dout  = 8'b00111111; // 1111 :  63 - 0x3f
      11'h458: dout  = 8'b00110000; // 1112 :  48 - 0x30
      11'h459: dout  = 8'b00111111; // 1113 :  63 - 0x3f
      11'h45A: dout  = 8'b00110000; // 1114 :  48 - 0x30
      11'h45B: dout  = 8'b00111111; // 1115 :  63 - 0x3f
      11'h45C: dout  = 8'b00110000; // 1116 :  48 - 0x30
      11'h45D: dout  = 8'b00111111; // 1117 :  63 - 0x3f
      11'h45E: dout  = 8'b00110000; // 1118 :  48 - 0x30
      11'h45F: dout  = 8'b00111111; // 1119 :  63 - 0x3f
      11'h460: dout  = 8'b00111111; // 1120 :  63 - 0x3f -- line 0x3
      11'h461: dout  = 8'b00111111; // 1121 :  63 - 0x3f
      11'h462: dout  = 8'b00111111; // 1122 :  63 - 0x3f
      11'h463: dout  = 8'b00111111; // 1123 :  63 - 0x3f
      11'h464: dout  = 8'b00111111; // 1124 :  63 - 0x3f
      11'h465: dout  = 8'b00111111; // 1125 :  63 - 0x3f
      11'h466: dout  = 8'b00111111; // 1126 :  63 - 0x3f
      11'h467: dout  = 8'b00111111; // 1127 :  63 - 0x3f
      11'h468: dout  = 8'b00111111; // 1128 :  63 - 0x3f
      11'h469: dout  = 8'b00111111; // 1129 :  63 - 0x3f
      11'h46A: dout  = 8'b00010000; // 1130 :  16 - 0x10
      11'h46B: dout  = 8'b00010001; // 1131 :  17 - 0x11
      11'h46C: dout  = 8'b00001101; // 1132 :  13 - 0xd
      11'h46D: dout  = 8'b00001111; // 1133 :  15 - 0xf
      11'h46E: dout  = 8'b00111111; // 1134 :  63 - 0x3f
      11'h46F: dout  = 8'b00110000; // 1135 :  48 - 0x30
      11'h470: dout  = 8'b00111111; // 1136 :  63 - 0x3f
      11'h471: dout  = 8'b00110000; // 1137 :  48 - 0x30
      11'h472: dout  = 8'b00111111; // 1138 :  63 - 0x3f
      11'h473: dout  = 8'b00110000; // 1139 :  48 - 0x30
      11'h474: dout  = 8'b00111111; // 1140 :  63 - 0x3f
      11'h475: dout  = 8'b00110000; // 1141 :  48 - 0x30
      11'h476: dout  = 8'b00111111; // 1142 :  63 - 0x3f
      11'h477: dout  = 8'b00110000; // 1143 :  48 - 0x30
      11'h478: dout  = 8'b00111111; // 1144 :  63 - 0x3f
      11'h479: dout  = 8'b00110000; // 1145 :  48 - 0x30
      11'h47A: dout  = 8'b00111111; // 1146 :  63 - 0x3f
      11'h47B: dout  = 8'b00110000; // 1147 :  48 - 0x30
      11'h47C: dout  = 8'b00111111; // 1148 :  63 - 0x3f
      11'h47D: dout  = 8'b00110000; // 1149 :  48 - 0x30
      11'h47E: dout  = 8'b00111111; // 1150 :  63 - 0x3f
      11'h47F: dout  = 8'b00110000; // 1151 :  48 - 0x30
      11'h480: dout  = 8'b00010100; // 1152 :  20 - 0x14 -- line 0x4
      11'h481: dout  = 8'b00010110; // 1153 :  22 - 0x16
      11'h482: dout  = 8'b00010100; // 1154 :  20 - 0x14
      11'h483: dout  = 8'b00010110; // 1155 :  22 - 0x16
      11'h484: dout  = 8'b00010100; // 1156 :  20 - 0x14
      11'h485: dout  = 8'b00010110; // 1157 :  22 - 0x16
      11'h486: dout  = 8'b00111111; // 1158 :  63 - 0x3f
      11'h487: dout  = 8'b00111111; // 1159 :  63 - 0x3f
      11'h488: dout  = 8'b00111111; // 1160 :  63 - 0x3f
      11'h489: dout  = 8'b00111111; // 1161 :  63 - 0x3f
      11'h48A: dout  = 8'b00010000; // 1162 :  16 - 0x10
      11'h48B: dout  = 8'b00010001; // 1163 :  17 - 0x11
      11'h48C: dout  = 8'b00001100; // 1164 :  12 - 0xc
      11'h48D: dout  = 8'b00001110; // 1165 :  14 - 0xe
      11'h48E: dout  = 8'b00111111; // 1166 :  63 - 0x3f
      11'h48F: dout  = 8'b00111111; // 1167 :  63 - 0x3f
      11'h490: dout  = 8'b00111111; // 1168 :  63 - 0x3f
      11'h491: dout  = 8'b00111111; // 1169 :  63 - 0x3f
      11'h492: dout  = 8'b00111111; // 1170 :  63 - 0x3f
      11'h493: dout  = 8'b00111111; // 1171 :  63 - 0x3f
      11'h494: dout  = 8'b00111111; // 1172 :  63 - 0x3f
      11'h495: dout  = 8'b00111111; // 1173 :  63 - 0x3f
      11'h496: dout  = 8'b00111111; // 1174 :  63 - 0x3f
      11'h497: dout  = 8'b00111111; // 1175 :  63 - 0x3f
      11'h498: dout  = 8'b00111111; // 1176 :  63 - 0x3f
      11'h499: dout  = 8'b00111111; // 1177 :  63 - 0x3f
      11'h49A: dout  = 8'b00111111; // 1178 :  63 - 0x3f
      11'h49B: dout  = 8'b00111111; // 1179 :  63 - 0x3f
      11'h49C: dout  = 8'b00111111; // 1180 :  63 - 0x3f
      11'h49D: dout  = 8'b00111111; // 1181 :  63 - 0x3f
      11'h49E: dout  = 8'b00111111; // 1182 :  63 - 0x3f
      11'h49F: dout  = 8'b00111111; // 1183 :  63 - 0x3f
      11'h4A0: dout  = 8'b00010101; // 1184 :  21 - 0x15 -- line 0x5
      11'h4A1: dout  = 8'b00010111; // 1185 :  23 - 0x17
      11'h4A2: dout  = 8'b00010101; // 1186 :  21 - 0x15
      11'h4A3: dout  = 8'b00010111; // 1187 :  23 - 0x17
      11'h4A4: dout  = 8'b00010101; // 1188 :  21 - 0x15
      11'h4A5: dout  = 8'b00010111; // 1189 :  23 - 0x17
      11'h4A6: dout  = 8'b00111111; // 1190 :  63 - 0x3f
      11'h4A7: dout  = 8'b00111111; // 1191 :  63 - 0x3f
      11'h4A8: dout  = 8'b00111111; // 1192 :  63 - 0x3f
      11'h4A9: dout  = 8'b00111111; // 1193 :  63 - 0x3f
      11'h4AA: dout  = 8'b00010000; // 1194 :  16 - 0x10
      11'h4AB: dout  = 8'b00010001; // 1195 :  17 - 0x11
      11'h4AC: dout  = 8'b00001101; // 1196 :  13 - 0xd
      11'h4AD: dout  = 8'b00001111; // 1197 :  15 - 0xf
      11'h4AE: dout  = 8'b00111111; // 1198 :  63 - 0x3f
      11'h4AF: dout  = 8'b00111111; // 1199 :  63 - 0x3f
      11'h4B0: dout  = 8'b00111111; // 1200 :  63 - 0x3f
      11'h4B1: dout  = 8'b00111111; // 1201 :  63 - 0x3f
      11'h4B2: dout  = 8'b00111111; // 1202 :  63 - 0x3f
      11'h4B3: dout  = 8'b00111111; // 1203 :  63 - 0x3f
      11'h4B4: dout  = 8'b00111111; // 1204 :  63 - 0x3f
      11'h4B5: dout  = 8'b00111111; // 1205 :  63 - 0x3f
      11'h4B6: dout  = 8'b00111111; // 1206 :  63 - 0x3f
      11'h4B7: dout  = 8'b00111111; // 1207 :  63 - 0x3f
      11'h4B8: dout  = 8'b00111111; // 1208 :  63 - 0x3f
      11'h4B9: dout  = 8'b00111111; // 1209 :  63 - 0x3f
      11'h4BA: dout  = 8'b00111111; // 1210 :  63 - 0x3f
      11'h4BB: dout  = 8'b00111111; // 1211 :  63 - 0x3f
      11'h4BC: dout  = 8'b00111111; // 1212 :  63 - 0x3f
      11'h4BD: dout  = 8'b00111111; // 1213 :  63 - 0x3f
      11'h4BE: dout  = 8'b00111111; // 1214 :  63 - 0x3f
      11'h4BF: dout  = 8'b00111111; // 1215 :  63 - 0x3f
      11'h4C0: dout  = 8'b00111111; // 1216 :  63 - 0x3f -- line 0x6
      11'h4C1: dout  = 8'b00111111; // 1217 :  63 - 0x3f
      11'h4C2: dout  = 8'b00111111; // 1218 :  63 - 0x3f
      11'h4C3: dout  = 8'b00111111; // 1219 :  63 - 0x3f
      11'h4C4: dout  = 8'b00111111; // 1220 :  63 - 0x3f
      11'h4C5: dout  = 8'b00111111; // 1221 :  63 - 0x3f
      11'h4C6: dout  = 8'b00111111; // 1222 :  63 - 0x3f
      11'h4C7: dout  = 8'b00111111; // 1223 :  63 - 0x3f
      11'h4C8: dout  = 8'b00111111; // 1224 :  63 - 0x3f
      11'h4C9: dout  = 8'b00111111; // 1225 :  63 - 0x3f
      11'h4CA: dout  = 8'b00010000; // 1226 :  16 - 0x10
      11'h4CB: dout  = 8'b00010001; // 1227 :  17 - 0x11
      11'h4CC: dout  = 8'b00001100; // 1228 :  12 - 0xc
      11'h4CD: dout  = 8'b00001110; // 1229 :  14 - 0xe
      11'h4CE: dout  = 8'b00111111; // 1230 :  63 - 0x3f
      11'h4CF: dout  = 8'b00111111; // 1231 :  63 - 0x3f
      11'h4D0: dout  = 8'b00111111; // 1232 :  63 - 0x3f
      11'h4D1: dout  = 8'b00111111; // 1233 :  63 - 0x3f
      11'h4D2: dout  = 8'b00111111; // 1234 :  63 - 0x3f
      11'h4D3: dout  = 8'b00111111; // 1235 :  63 - 0x3f
      11'h4D4: dout  = 8'b00111111; // 1236 :  63 - 0x3f
      11'h4D5: dout  = 8'b00111111; // 1237 :  63 - 0x3f
      11'h4D6: dout  = 8'b00111111; // 1238 :  63 - 0x3f
      11'h4D7: dout  = 8'b00111111; // 1239 :  63 - 0x3f
      11'h4D8: dout  = 8'b00111111; // 1240 :  63 - 0x3f
      11'h4D9: dout  = 8'b00111111; // 1241 :  63 - 0x3f
      11'h4DA: dout  = 8'b00111111; // 1242 :  63 - 0x3f
      11'h4DB: dout  = 8'b00111111; // 1243 :  63 - 0x3f
      11'h4DC: dout  = 8'b00111111; // 1244 :  63 - 0x3f
      11'h4DD: dout  = 8'b00111111; // 1245 :  63 - 0x3f
      11'h4DE: dout  = 8'b00111111; // 1246 :  63 - 0x3f
      11'h4DF: dout  = 8'b00111111; // 1247 :  63 - 0x3f
      11'h4E0: dout  = 8'b00111111; // 1248 :  63 - 0x3f -- line 0x7
      11'h4E1: dout  = 8'b00111111; // 1249 :  63 - 0x3f
      11'h4E2: dout  = 8'b00111111; // 1250 :  63 - 0x3f
      11'h4E3: dout  = 8'b00111111; // 1251 :  63 - 0x3f
      11'h4E4: dout  = 8'b00111111; // 1252 :  63 - 0x3f
      11'h4E5: dout  = 8'b00111111; // 1253 :  63 - 0x3f
      11'h4E6: dout  = 8'b00111111; // 1254 :  63 - 0x3f
      11'h4E7: dout  = 8'b00111111; // 1255 :  63 - 0x3f
      11'h4E8: dout  = 8'b00111111; // 1256 :  63 - 0x3f
      11'h4E9: dout  = 8'b00111111; // 1257 :  63 - 0x3f
      11'h4EA: dout  = 8'b00010000; // 1258 :  16 - 0x10
      11'h4EB: dout  = 8'b00010001; // 1259 :  17 - 0x11
      11'h4EC: dout  = 8'b00001101; // 1260 :  13 - 0xd
      11'h4ED: dout  = 8'b00001111; // 1261 :  15 - 0xf
      11'h4EE: dout  = 8'b00111111; // 1262 :  63 - 0x3f
      11'h4EF: dout  = 8'b00111111; // 1263 :  63 - 0x3f
      11'h4F0: dout  = 8'b00111111; // 1264 :  63 - 0x3f
      11'h4F1: dout  = 8'b00111111; // 1265 :  63 - 0x3f
      11'h4F2: dout  = 8'b00111111; // 1266 :  63 - 0x3f
      11'h4F3: dout  = 8'b00111111; // 1267 :  63 - 0x3f
      11'h4F4: dout  = 8'b00111111; // 1268 :  63 - 0x3f
      11'h4F5: dout  = 8'b00111111; // 1269 :  63 - 0x3f
      11'h4F6: dout  = 8'b00111111; // 1270 :  63 - 0x3f
      11'h4F7: dout  = 8'b00111111; // 1271 :  63 - 0x3f
      11'h4F8: dout  = 8'b00111111; // 1272 :  63 - 0x3f
      11'h4F9: dout  = 8'b00111111; // 1273 :  63 - 0x3f
      11'h4FA: dout  = 8'b00111111; // 1274 :  63 - 0x3f
      11'h4FB: dout  = 8'b00111111; // 1275 :  63 - 0x3f
      11'h4FC: dout  = 8'b00111111; // 1276 :  63 - 0x3f
      11'h4FD: dout  = 8'b00111111; // 1277 :  63 - 0x3f
      11'h4FE: dout  = 8'b00111111; // 1278 :  63 - 0x3f
      11'h4FF: dout  = 8'b00111111; // 1279 :  63 - 0x3f
      11'h500: dout  = 8'b00111111; // 1280 :  63 - 0x3f -- line 0x8
      11'h501: dout  = 8'b00111111; // 1281 :  63 - 0x3f
      11'h502: dout  = 8'b00001100; // 1282 :  12 - 0xc
      11'h503: dout  = 8'b00001110; // 1283 :  14 - 0xe
      11'h504: dout  = 8'b00001100; // 1284 :  12 - 0xc
      11'h505: dout  = 8'b00001110; // 1285 :  14 - 0xe
      11'h506: dout  = 8'b00001100; // 1286 :  12 - 0xc
      11'h507: dout  = 8'b00001110; // 1287 :  14 - 0xe
      11'h508: dout  = 8'b00001100; // 1288 :  12 - 0xc
      11'h509: dout  = 8'b00001110; // 1289 :  14 - 0xe
      11'h50A: dout  = 8'b00001100; // 1290 :  12 - 0xc
      11'h50B: dout  = 8'b00001110; // 1291 :  14 - 0xe
      11'h50C: dout  = 8'b00001100; // 1292 :  12 - 0xc
      11'h50D: dout  = 8'b00001110; // 1293 :  14 - 0xe
      11'h50E: dout  = 8'b00111111; // 1294 :  63 - 0x3f
      11'h50F: dout  = 8'b00111111; // 1295 :  63 - 0x3f
      11'h510: dout  = 8'b00111111; // 1296 :  63 - 0x3f
      11'h511: dout  = 8'b00111111; // 1297 :  63 - 0x3f
      11'h512: dout  = 8'b00111111; // 1298 :  63 - 0x3f
      11'h513: dout  = 8'b00111111; // 1299 :  63 - 0x3f
      11'h514: dout  = 8'b00111111; // 1300 :  63 - 0x3f
      11'h515: dout  = 8'b00111111; // 1301 :  63 - 0x3f
      11'h516: dout  = 8'b00111111; // 1302 :  63 - 0x3f
      11'h517: dout  = 8'b00111111; // 1303 :  63 - 0x3f
      11'h518: dout  = 8'b00111111; // 1304 :  63 - 0x3f
      11'h519: dout  = 8'b00111111; // 1305 :  63 - 0x3f
      11'h51A: dout  = 8'b00111111; // 1306 :  63 - 0x3f
      11'h51B: dout  = 8'b00111111; // 1307 :  63 - 0x3f
      11'h51C: dout  = 8'b00111111; // 1308 :  63 - 0x3f
      11'h51D: dout  = 8'b00111111; // 1309 :  63 - 0x3f
      11'h51E: dout  = 8'b00111111; // 1310 :  63 - 0x3f
      11'h51F: dout  = 8'b00111111; // 1311 :  63 - 0x3f
      11'h520: dout  = 8'b00111111; // 1312 :  63 - 0x3f -- line 0x9
      11'h521: dout  = 8'b00111111; // 1313 :  63 - 0x3f
      11'h522: dout  = 8'b00001101; // 1314 :  13 - 0xd
      11'h523: dout  = 8'b00001111; // 1315 :  15 - 0xf
      11'h524: dout  = 8'b00001101; // 1316 :  13 - 0xd
      11'h525: dout  = 8'b00001111; // 1317 :  15 - 0xf
      11'h526: dout  = 8'b00001101; // 1318 :  13 - 0xd
      11'h527: dout  = 8'b00001111; // 1319 :  15 - 0xf
      11'h528: dout  = 8'b00001101; // 1320 :  13 - 0xd
      11'h529: dout  = 8'b00001111; // 1321 :  15 - 0xf
      11'h52A: dout  = 8'b00001101; // 1322 :  13 - 0xd
      11'h52B: dout  = 8'b00001111; // 1323 :  15 - 0xf
      11'h52C: dout  = 8'b00001101; // 1324 :  13 - 0xd
      11'h52D: dout  = 8'b00001111; // 1325 :  15 - 0xf
      11'h52E: dout  = 8'b00111111; // 1326 :  63 - 0x3f
      11'h52F: dout  = 8'b00111111; // 1327 :  63 - 0x3f
      11'h530: dout  = 8'b00111111; // 1328 :  63 - 0x3f
      11'h531: dout  = 8'b00111111; // 1329 :  63 - 0x3f
      11'h532: dout  = 8'b00111111; // 1330 :  63 - 0x3f
      11'h533: dout  = 8'b00111111; // 1331 :  63 - 0x3f
      11'h534: dout  = 8'b00111111; // 1332 :  63 - 0x3f
      11'h535: dout  = 8'b00111111; // 1333 :  63 - 0x3f
      11'h536: dout  = 8'b00111111; // 1334 :  63 - 0x3f
      11'h537: dout  = 8'b00111111; // 1335 :  63 - 0x3f
      11'h538: dout  = 8'b00111111; // 1336 :  63 - 0x3f
      11'h539: dout  = 8'b00111111; // 1337 :  63 - 0x3f
      11'h53A: dout  = 8'b00111111; // 1338 :  63 - 0x3f
      11'h53B: dout  = 8'b00111111; // 1339 :  63 - 0x3f
      11'h53C: dout  = 8'b00111111; // 1340 :  63 - 0x3f
      11'h53D: dout  = 8'b00111111; // 1341 :  63 - 0x3f
      11'h53E: dout  = 8'b00111111; // 1342 :  63 - 0x3f
      11'h53F: dout  = 8'b00111111; // 1343 :  63 - 0x3f
      11'h540: dout  = 8'b01011000; // 1344 :  88 - 0x58 -- line 0xa
      11'h541: dout  = 8'b01011000; // 1345 :  88 - 0x58
      11'h542: dout  = 8'b01011000; // 1346 :  88 - 0x58
      11'h543: dout  = 8'b01011001; // 1347 :  89 - 0x59
      11'h544: dout  = 8'b00111111; // 1348 :  63 - 0x3f
      11'h545: dout  = 8'b00111111; // 1349 :  63 - 0x3f
      11'h546: dout  = 8'b00111111; // 1350 :  63 - 0x3f
      11'h547: dout  = 8'b00111111; // 1351 :  63 - 0x3f
      11'h548: dout  = 8'b00111111; // 1352 :  63 - 0x3f
      11'h549: dout  = 8'b00111111; // 1353 :  63 - 0x3f
      11'h54A: dout  = 8'b00111111; // 1354 :  63 - 0x3f
      11'h54B: dout  = 8'b00111111; // 1355 :  63 - 0x3f
      11'h54C: dout  = 8'b00111111; // 1356 :  63 - 0x3f
      11'h54D: dout  = 8'b00111111; // 1357 :  63 - 0x3f
      11'h54E: dout  = 8'b00111111; // 1358 :  63 - 0x3f
      11'h54F: dout  = 8'b00111111; // 1359 :  63 - 0x3f
      11'h550: dout  = 8'b00111111; // 1360 :  63 - 0x3f
      11'h551: dout  = 8'b00111111; // 1361 :  63 - 0x3f
      11'h552: dout  = 8'b00111111; // 1362 :  63 - 0x3f
      11'h553: dout  = 8'b00111111; // 1363 :  63 - 0x3f
      11'h554: dout  = 8'b00111111; // 1364 :  63 - 0x3f
      11'h555: dout  = 8'b00111111; // 1365 :  63 - 0x3f
      11'h556: dout  = 8'b00111111; // 1366 :  63 - 0x3f
      11'h557: dout  = 8'b00111111; // 1367 :  63 - 0x3f
      11'h558: dout  = 8'b00111111; // 1368 :  63 - 0x3f
      11'h559: dout  = 8'b00111111; // 1369 :  63 - 0x3f
      11'h55A: dout  = 8'b00010100; // 1370 :  20 - 0x14
      11'h55B: dout  = 8'b00010110; // 1371 :  22 - 0x16
      11'h55C: dout  = 8'b00010100; // 1372 :  20 - 0x14
      11'h55D: dout  = 8'b00010110; // 1373 :  22 - 0x16
      11'h55E: dout  = 8'b00010100; // 1374 :  20 - 0x14
      11'h55F: dout  = 8'b00010110; // 1375 :  22 - 0x16
      11'h560: dout  = 8'b00111111; // 1376 :  63 - 0x3f -- line 0xb
      11'h561: dout  = 8'b00111111; // 1377 :  63 - 0x3f
      11'h562: dout  = 8'b00111111; // 1378 :  63 - 0x3f
      11'h563: dout  = 8'b00111111; // 1379 :  63 - 0x3f
      11'h564: dout  = 8'b00111111; // 1380 :  63 - 0x3f
      11'h565: dout  = 8'b00111111; // 1381 :  63 - 0x3f
      11'h566: dout  = 8'b00111111; // 1382 :  63 - 0x3f
      11'h567: dout  = 8'b00111111; // 1383 :  63 - 0x3f
      11'h568: dout  = 8'b00111111; // 1384 :  63 - 0x3f
      11'h569: dout  = 8'b00111111; // 1385 :  63 - 0x3f
      11'h56A: dout  = 8'b00111111; // 1386 :  63 - 0x3f
      11'h56B: dout  = 8'b00111111; // 1387 :  63 - 0x3f
      11'h56C: dout  = 8'b00111111; // 1388 :  63 - 0x3f
      11'h56D: dout  = 8'b00111111; // 1389 :  63 - 0x3f
      11'h56E: dout  = 8'b00111111; // 1390 :  63 - 0x3f
      11'h56F: dout  = 8'b00111111; // 1391 :  63 - 0x3f
      11'h570: dout  = 8'b00111111; // 1392 :  63 - 0x3f
      11'h571: dout  = 8'b00111111; // 1393 :  63 - 0x3f
      11'h572: dout  = 8'b00111111; // 1394 :  63 - 0x3f
      11'h573: dout  = 8'b00111111; // 1395 :  63 - 0x3f
      11'h574: dout  = 8'b00111111; // 1396 :  63 - 0x3f
      11'h575: dout  = 8'b00111111; // 1397 :  63 - 0x3f
      11'h576: dout  = 8'b00111111; // 1398 :  63 - 0x3f
      11'h577: dout  = 8'b00111111; // 1399 :  63 - 0x3f
      11'h578: dout  = 8'b00111111; // 1400 :  63 - 0x3f
      11'h579: dout  = 8'b00111111; // 1401 :  63 - 0x3f
      11'h57A: dout  = 8'b00010101; // 1402 :  21 - 0x15
      11'h57B: dout  = 8'b00010111; // 1403 :  23 - 0x17
      11'h57C: dout  = 8'b00010101; // 1404 :  21 - 0x15
      11'h57D: dout  = 8'b00010111; // 1405 :  23 - 0x17
      11'h57E: dout  = 8'b00010101; // 1406 :  21 - 0x15
      11'h57F: dout  = 8'b00010111; // 1407 :  23 - 0x17
      11'h580: dout  = 8'b00111111; // 1408 :  63 - 0x3f -- line 0xc
      11'h581: dout  = 8'b00111111; // 1409 :  63 - 0x3f
      11'h582: dout  = 8'b00111111; // 1410 :  63 - 0x3f
      11'h583: dout  = 8'b00111111; // 1411 :  63 - 0x3f
      11'h584: dout  = 8'b00111111; // 1412 :  63 - 0x3f
      11'h585: dout  = 8'b00111111; // 1413 :  63 - 0x3f
      11'h586: dout  = 8'b00111111; // 1414 :  63 - 0x3f
      11'h587: dout  = 8'b00111111; // 1415 :  63 - 0x3f
      11'h588: dout  = 8'b00111111; // 1416 :  63 - 0x3f
      11'h589: dout  = 8'b00111111; // 1417 :  63 - 0x3f
      11'h58A: dout  = 8'b00111111; // 1418 :  63 - 0x3f
      11'h58B: dout  = 8'b00111111; // 1419 :  63 - 0x3f
      11'h58C: dout  = 8'b00111111; // 1420 :  63 - 0x3f
      11'h58D: dout  = 8'b00111111; // 1421 :  63 - 0x3f
      11'h58E: dout  = 8'b00111111; // 1422 :  63 - 0x3f
      11'h58F: dout  = 8'b00111111; // 1423 :  63 - 0x3f
      11'h590: dout  = 8'b00111111; // 1424 :  63 - 0x3f
      11'h591: dout  = 8'b00111111; // 1425 :  63 - 0x3f
      11'h592: dout  = 8'b00111111; // 1426 :  63 - 0x3f
      11'h593: dout  = 8'b00111111; // 1427 :  63 - 0x3f
      11'h594: dout  = 8'b00111111; // 1428 :  63 - 0x3f
      11'h595: dout  = 8'b00111111; // 1429 :  63 - 0x3f
      11'h596: dout  = 8'b00111111; // 1430 :  63 - 0x3f
      11'h597: dout  = 8'b00111111; // 1431 :  63 - 0x3f
      11'h598: dout  = 8'b00111111; // 1432 :  63 - 0x3f
      11'h599: dout  = 8'b00111111; // 1433 :  63 - 0x3f
      11'h59A: dout  = 8'b00111111; // 1434 :  63 - 0x3f
      11'h59B: dout  = 8'b00111111; // 1435 :  63 - 0x3f
      11'h59C: dout  = 8'b00111111; // 1436 :  63 - 0x3f
      11'h59D: dout  = 8'b00111111; // 1437 :  63 - 0x3f
      11'h59E: dout  = 8'b00111111; // 1438 :  63 - 0x3f
      11'h59F: dout  = 8'b00111111; // 1439 :  63 - 0x3f
      11'h5A0: dout  = 8'b00111111; // 1440 :  63 - 0x3f -- line 0xd
      11'h5A1: dout  = 8'b00111111; // 1441 :  63 - 0x3f
      11'h5A2: dout  = 8'b00111111; // 1442 :  63 - 0x3f
      11'h5A3: dout  = 8'b00111111; // 1443 :  63 - 0x3f
      11'h5A4: dout  = 8'b00111111; // 1444 :  63 - 0x3f
      11'h5A5: dout  = 8'b00111111; // 1445 :  63 - 0x3f
      11'h5A6: dout  = 8'b00111111; // 1446 :  63 - 0x3f
      11'h5A7: dout  = 8'b00111111; // 1447 :  63 - 0x3f
      11'h5A8: dout  = 8'b00111111; // 1448 :  63 - 0x3f
      11'h5A9: dout  = 8'b00111111; // 1449 :  63 - 0x3f
      11'h5AA: dout  = 8'b00111111; // 1450 :  63 - 0x3f
      11'h5AB: dout  = 8'b00111111; // 1451 :  63 - 0x3f
      11'h5AC: dout  = 8'b00111111; // 1452 :  63 - 0x3f
      11'h5AD: dout  = 8'b00111111; // 1453 :  63 - 0x3f
      11'h5AE: dout  = 8'b00111111; // 1454 :  63 - 0x3f
      11'h5AF: dout  = 8'b00111111; // 1455 :  63 - 0x3f
      11'h5B0: dout  = 8'b00111111; // 1456 :  63 - 0x3f
      11'h5B1: dout  = 8'b00111111; // 1457 :  63 - 0x3f
      11'h5B2: dout  = 8'b00111111; // 1458 :  63 - 0x3f
      11'h5B3: dout  = 8'b00111111; // 1459 :  63 - 0x3f
      11'h5B4: dout  = 8'b00111111; // 1460 :  63 - 0x3f
      11'h5B5: dout  = 8'b00111111; // 1461 :  63 - 0x3f
      11'h5B6: dout  = 8'b00111111; // 1462 :  63 - 0x3f
      11'h5B7: dout  = 8'b00111111; // 1463 :  63 - 0x3f
      11'h5B8: dout  = 8'b00111111; // 1464 :  63 - 0x3f
      11'h5B9: dout  = 8'b00111111; // 1465 :  63 - 0x3f
      11'h5BA: dout  = 8'b00111111; // 1466 :  63 - 0x3f
      11'h5BB: dout  = 8'b00111111; // 1467 :  63 - 0x3f
      11'h5BC: dout  = 8'b00111111; // 1468 :  63 - 0x3f
      11'h5BD: dout  = 8'b00111111; // 1469 :  63 - 0x3f
      11'h5BE: dout  = 8'b00111111; // 1470 :  63 - 0x3f
      11'h5BF: dout  = 8'b00111111; // 1471 :  63 - 0x3f
      11'h5C0: dout  = 8'b00111111; // 1472 :  63 - 0x3f -- line 0xe
      11'h5C1: dout  = 8'b00111111; // 1473 :  63 - 0x3f
      11'h5C2: dout  = 8'b00111111; // 1474 :  63 - 0x3f
      11'h5C3: dout  = 8'b00111111; // 1475 :  63 - 0x3f
      11'h5C4: dout  = 8'b00111111; // 1476 :  63 - 0x3f
      11'h5C5: dout  = 8'b00111111; // 1477 :  63 - 0x3f
      11'h5C6: dout  = 8'b00111111; // 1478 :  63 - 0x3f
      11'h5C7: dout  = 8'b00111111; // 1479 :  63 - 0x3f
      11'h5C8: dout  = 8'b00111111; // 1480 :  63 - 0x3f
      11'h5C9: dout  = 8'b00111111; // 1481 :  63 - 0x3f
      11'h5CA: dout  = 8'b00111111; // 1482 :  63 - 0x3f
      11'h5CB: dout  = 8'b00111111; // 1483 :  63 - 0x3f
      11'h5CC: dout  = 8'b00111111; // 1484 :  63 - 0x3f
      11'h5CD: dout  = 8'b00111111; // 1485 :  63 - 0x3f
      11'h5CE: dout  = 8'b00111111; // 1486 :  63 - 0x3f
      11'h5CF: dout  = 8'b00111111; // 1487 :  63 - 0x3f
      11'h5D0: dout  = 8'b00111111; // 1488 :  63 - 0x3f
      11'h5D1: dout  = 8'b00111111; // 1489 :  63 - 0x3f
      11'h5D2: dout  = 8'b00111111; // 1490 :  63 - 0x3f
      11'h5D3: dout  = 8'b00111111; // 1491 :  63 - 0x3f
      11'h5D4: dout  = 8'b00111111; // 1492 :  63 - 0x3f
      11'h5D5: dout  = 8'b00111111; // 1493 :  63 - 0x3f
      11'h5D6: dout  = 8'b00111111; // 1494 :  63 - 0x3f
      11'h5D7: dout  = 8'b00111111; // 1495 :  63 - 0x3f
      11'h5D8: dout  = 8'b01010111; // 1496 :  87 - 0x57
      11'h5D9: dout  = 8'b01011000; // 1497 :  88 - 0x58
      11'h5DA: dout  = 8'b01011000; // 1498 :  88 - 0x58
      11'h5DB: dout  = 8'b01011000; // 1499 :  88 - 0x58
      11'h5DC: dout  = 8'b01011000; // 1500 :  88 - 0x58
      11'h5DD: dout  = 8'b01011000; // 1501 :  88 - 0x58
      11'h5DE: dout  = 8'b01011000; // 1502 :  88 - 0x58
      11'h5DF: dout  = 8'b01011000; // 1503 :  88 - 0x58
      11'h5E0: dout  = 8'b00111111; // 1504 :  63 - 0x3f -- line 0xf
      11'h5E1: dout  = 8'b00111111; // 1505 :  63 - 0x3f
      11'h5E2: dout  = 8'b00111111; // 1506 :  63 - 0x3f
      11'h5E3: dout  = 8'b00111111; // 1507 :  63 - 0x3f
      11'h5E4: dout  = 8'b00111111; // 1508 :  63 - 0x3f
      11'h5E5: dout  = 8'b00111111; // 1509 :  63 - 0x3f
      11'h5E6: dout  = 8'b00111111; // 1510 :  63 - 0x3f
      11'h5E7: dout  = 8'b00111111; // 1511 :  63 - 0x3f
      11'h5E8: dout  = 8'b00111111; // 1512 :  63 - 0x3f
      11'h5E9: dout  = 8'b00111111; // 1513 :  63 - 0x3f
      11'h5EA: dout  = 8'b00111111; // 1514 :  63 - 0x3f
      11'h5EB: dout  = 8'b00111111; // 1515 :  63 - 0x3f
      11'h5EC: dout  = 8'b00111111; // 1516 :  63 - 0x3f
      11'h5ED: dout  = 8'b00111111; // 1517 :  63 - 0x3f
      11'h5EE: dout  = 8'b00111111; // 1518 :  63 - 0x3f
      11'h5EF: dout  = 8'b00111111; // 1519 :  63 - 0x3f
      11'h5F0: dout  = 8'b00111111; // 1520 :  63 - 0x3f
      11'h5F1: dout  = 8'b00111111; // 1521 :  63 - 0x3f
      11'h5F2: dout  = 8'b00111111; // 1522 :  63 - 0x3f
      11'h5F3: dout  = 8'b00111111; // 1523 :  63 - 0x3f
      11'h5F4: dout  = 8'b00111111; // 1524 :  63 - 0x3f
      11'h5F5: dout  = 8'b00111111; // 1525 :  63 - 0x3f
      11'h5F6: dout  = 8'b00111111; // 1526 :  63 - 0x3f
      11'h5F7: dout  = 8'b00111111; // 1527 :  63 - 0x3f
      11'h5F8: dout  = 8'b00111111; // 1528 :  63 - 0x3f
      11'h5F9: dout  = 8'b00111111; // 1529 :  63 - 0x3f
      11'h5FA: dout  = 8'b00111111; // 1530 :  63 - 0x3f
      11'h5FB: dout  = 8'b00111111; // 1531 :  63 - 0x3f
      11'h5FC: dout  = 8'b00111111; // 1532 :  63 - 0x3f
      11'h5FD: dout  = 8'b00111111; // 1533 :  63 - 0x3f
      11'h5FE: dout  = 8'b00111111; // 1534 :  63 - 0x3f
      11'h5FF: dout  = 8'b00111111; // 1535 :  63 - 0x3f
      11'h600: dout  = 8'b00111111; // 1536 :  63 - 0x3f -- line 0x10
      11'h601: dout  = 8'b00111111; // 1537 :  63 - 0x3f
      11'h602: dout  = 8'b00111111; // 1538 :  63 - 0x3f
      11'h603: dout  = 8'b00111111; // 1539 :  63 - 0x3f
      11'h604: dout  = 8'b00111111; // 1540 :  63 - 0x3f
      11'h605: dout  = 8'b00111111; // 1541 :  63 - 0x3f
      11'h606: dout  = 8'b00111111; // 1542 :  63 - 0x3f
      11'h607: dout  = 8'b00111111; // 1543 :  63 - 0x3f
      11'h608: dout  = 8'b00111111; // 1544 :  63 - 0x3f
      11'h609: dout  = 8'b00111111; // 1545 :  63 - 0x3f
      11'h60A: dout  = 8'b00111111; // 1546 :  63 - 0x3f
      11'h60B: dout  = 8'b00111111; // 1547 :  63 - 0x3f
      11'h60C: dout  = 8'b00111111; // 1548 :  63 - 0x3f
      11'h60D: dout  = 8'b00111111; // 1549 :  63 - 0x3f
      11'h60E: dout  = 8'b00111111; // 1550 :  63 - 0x3f
      11'h60F: dout  = 8'b00111111; // 1551 :  63 - 0x3f
      11'h610: dout  = 8'b00111111; // 1552 :  63 - 0x3f
      11'h611: dout  = 8'b00111111; // 1553 :  63 - 0x3f
      11'h612: dout  = 8'b00111111; // 1554 :  63 - 0x3f
      11'h613: dout  = 8'b00111111; // 1555 :  63 - 0x3f
      11'h614: dout  = 8'b00111111; // 1556 :  63 - 0x3f
      11'h615: dout  = 8'b00111111; // 1557 :  63 - 0x3f
      11'h616: dout  = 8'b00111111; // 1558 :  63 - 0x3f
      11'h617: dout  = 8'b00111111; // 1559 :  63 - 0x3f
      11'h618: dout  = 8'b00111111; // 1560 :  63 - 0x3f
      11'h619: dout  = 8'b00111111; // 1561 :  63 - 0x3f
      11'h61A: dout  = 8'b00111111; // 1562 :  63 - 0x3f
      11'h61B: dout  = 8'b00111111; // 1563 :  63 - 0x3f
      11'h61C: dout  = 8'b00111111; // 1564 :  63 - 0x3f
      11'h61D: dout  = 8'b00111111; // 1565 :  63 - 0x3f
      11'h61E: dout  = 8'b00111111; // 1566 :  63 - 0x3f
      11'h61F: dout  = 8'b00111111; // 1567 :  63 - 0x3f
      11'h620: dout  = 8'b00111111; // 1568 :  63 - 0x3f -- line 0x11
      11'h621: dout  = 8'b00111111; // 1569 :  63 - 0x3f
      11'h622: dout  = 8'b00111111; // 1570 :  63 - 0x3f
      11'h623: dout  = 8'b00111111; // 1571 :  63 - 0x3f
      11'h624: dout  = 8'b00111111; // 1572 :  63 - 0x3f
      11'h625: dout  = 8'b00111111; // 1573 :  63 - 0x3f
      11'h626: dout  = 8'b00111111; // 1574 :  63 - 0x3f
      11'h627: dout  = 8'b00111111; // 1575 :  63 - 0x3f
      11'h628: dout  = 8'b00111111; // 1576 :  63 - 0x3f
      11'h629: dout  = 8'b00111111; // 1577 :  63 - 0x3f
      11'h62A: dout  = 8'b00111111; // 1578 :  63 - 0x3f
      11'h62B: dout  = 8'b00111111; // 1579 :  63 - 0x3f
      11'h62C: dout  = 8'b00111111; // 1580 :  63 - 0x3f
      11'h62D: dout  = 8'b00111111; // 1581 :  63 - 0x3f
      11'h62E: dout  = 8'b00111111; // 1582 :  63 - 0x3f
      11'h62F: dout  = 8'b00111111; // 1583 :  63 - 0x3f
      11'h630: dout  = 8'b00111111; // 1584 :  63 - 0x3f
      11'h631: dout  = 8'b00111111; // 1585 :  63 - 0x3f
      11'h632: dout  = 8'b00111111; // 1586 :  63 - 0x3f
      11'h633: dout  = 8'b00111111; // 1587 :  63 - 0x3f
      11'h634: dout  = 8'b00111111; // 1588 :  63 - 0x3f
      11'h635: dout  = 8'b00111111; // 1589 :  63 - 0x3f
      11'h636: dout  = 8'b00111111; // 1590 :  63 - 0x3f
      11'h637: dout  = 8'b00111111; // 1591 :  63 - 0x3f
      11'h638: dout  = 8'b00111111; // 1592 :  63 - 0x3f
      11'h639: dout  = 8'b00111111; // 1593 :  63 - 0x3f
      11'h63A: dout  = 8'b00111111; // 1594 :  63 - 0x3f
      11'h63B: dout  = 8'b00111111; // 1595 :  63 - 0x3f
      11'h63C: dout  = 8'b00111111; // 1596 :  63 - 0x3f
      11'h63D: dout  = 8'b00111111; // 1597 :  63 - 0x3f
      11'h63E: dout  = 8'b00111111; // 1598 :  63 - 0x3f
      11'h63F: dout  = 8'b00111111; // 1599 :  63 - 0x3f
      11'h640: dout  = 8'b00111111; // 1600 :  63 - 0x3f -- line 0x12
      11'h641: dout  = 8'b00111111; // 1601 :  63 - 0x3f
      11'h642: dout  = 8'b00111111; // 1602 :  63 - 0x3f
      11'h643: dout  = 8'b00111111; // 1603 :  63 - 0x3f
      11'h644: dout  = 8'b00111111; // 1604 :  63 - 0x3f
      11'h645: dout  = 8'b00111111; // 1605 :  63 - 0x3f
      11'h646: dout  = 8'b00111111; // 1606 :  63 - 0x3f
      11'h647: dout  = 8'b00111111; // 1607 :  63 - 0x3f
      11'h648: dout  = 8'b00111111; // 1608 :  63 - 0x3f
      11'h649: dout  = 8'b00111111; // 1609 :  63 - 0x3f
      11'h64A: dout  = 8'b00111111; // 1610 :  63 - 0x3f
      11'h64B: dout  = 8'b00111111; // 1611 :  63 - 0x3f
      11'h64C: dout  = 8'b11011100; // 1612 : 220 - 0xdc
      11'h64D: dout  = 8'b11011101; // 1613 : 221 - 0xdd
      11'h64E: dout  = 8'b11001100; // 1614 : 204 - 0xcc
      11'h64F: dout  = 8'b11001101; // 1615 : 205 - 0xcd
      11'h650: dout  = 8'b00111111; // 1616 :  63 - 0x3f
      11'h651: dout  = 8'b00111111; // 1617 :  63 - 0x3f
      11'h652: dout  = 8'b00111111; // 1618 :  63 - 0x3f
      11'h653: dout  = 8'b00111111; // 1619 :  63 - 0x3f
      11'h654: dout  = 8'b00111111; // 1620 :  63 - 0x3f
      11'h655: dout  = 8'b00111111; // 1621 :  63 - 0x3f
      11'h656: dout  = 8'b00111111; // 1622 :  63 - 0x3f
      11'h657: dout  = 8'b00111111; // 1623 :  63 - 0x3f
      11'h658: dout  = 8'b00111111; // 1624 :  63 - 0x3f
      11'h659: dout  = 8'b00111111; // 1625 :  63 - 0x3f
      11'h65A: dout  = 8'b00111111; // 1626 :  63 - 0x3f
      11'h65B: dout  = 8'b00111111; // 1627 :  63 - 0x3f
      11'h65C: dout  = 8'b00111111; // 1628 :  63 - 0x3f
      11'h65D: dout  = 8'b00111111; // 1629 :  63 - 0x3f
      11'h65E: dout  = 8'b00111111; // 1630 :  63 - 0x3f
      11'h65F: dout  = 8'b00111111; // 1631 :  63 - 0x3f
      11'h660: dout  = 8'b00111111; // 1632 :  63 - 0x3f -- line 0x13
      11'h661: dout  = 8'b00111111; // 1633 :  63 - 0x3f
      11'h662: dout  = 8'b00111111; // 1634 :  63 - 0x3f
      11'h663: dout  = 8'b00111111; // 1635 :  63 - 0x3f
      11'h664: dout  = 8'b00111111; // 1636 :  63 - 0x3f
      11'h665: dout  = 8'b00111111; // 1637 :  63 - 0x3f
      11'h666: dout  = 8'b00111111; // 1638 :  63 - 0x3f
      11'h667: dout  = 8'b00111111; // 1639 :  63 - 0x3f
      11'h668: dout  = 8'b00111111; // 1640 :  63 - 0x3f
      11'h669: dout  = 8'b00111111; // 1641 :  63 - 0x3f
      11'h66A: dout  = 8'b00111111; // 1642 :  63 - 0x3f
      11'h66B: dout  = 8'b00111111; // 1643 :  63 - 0x3f
      11'h66C: dout  = 8'b11011010; // 1644 : 218 - 0xda
      11'h66D: dout  = 8'b11011011; // 1645 : 219 - 0xdb
      11'h66E: dout  = 8'b11011010; // 1646 : 218 - 0xda
      11'h66F: dout  = 8'b11011011; // 1647 : 219 - 0xdb
      11'h670: dout  = 8'b00111111; // 1648 :  63 - 0x3f
      11'h671: dout  = 8'b00111111; // 1649 :  63 - 0x3f
      11'h672: dout  = 8'b00011000; // 1650 :  24 - 0x18
      11'h673: dout  = 8'b00011001; // 1651 :  25 - 0x19
      11'h674: dout  = 8'b00111111; // 1652 :  63 - 0x3f
      11'h675: dout  = 8'b00111111; // 1653 :  63 - 0x3f
      11'h676: dout  = 8'b00111111; // 1654 :  63 - 0x3f
      11'h677: dout  = 8'b00111111; // 1655 :  63 - 0x3f
      11'h678: dout  = 8'b00111111; // 1656 :  63 - 0x3f
      11'h679: dout  = 8'b00111111; // 1657 :  63 - 0x3f
      11'h67A: dout  = 8'b00111111; // 1658 :  63 - 0x3f
      11'h67B: dout  = 8'b00111111; // 1659 :  63 - 0x3f
      11'h67C: dout  = 8'b00111111; // 1660 :  63 - 0x3f
      11'h67D: dout  = 8'b00111111; // 1661 :  63 - 0x3f
      11'h67E: dout  = 8'b00111111; // 1662 :  63 - 0x3f
      11'h67F: dout  = 8'b00111111; // 1663 :  63 - 0x3f
      11'h680: dout  = 8'b00111111; // 1664 :  63 - 0x3f -- line 0x14
      11'h681: dout  = 8'b00111111; // 1665 :  63 - 0x3f
      11'h682: dout  = 8'b00111111; // 1666 :  63 - 0x3f
      11'h683: dout  = 8'b00111111; // 1667 :  63 - 0x3f
      11'h684: dout  = 8'b00111111; // 1668 :  63 - 0x3f
      11'h685: dout  = 8'b00111111; // 1669 :  63 - 0x3f
      11'h686: dout  = 8'b00111111; // 1670 :  63 - 0x3f
      11'h687: dout  = 8'b00111111; // 1671 :  63 - 0x3f
      11'h688: dout  = 8'b00111111; // 1672 :  63 - 0x3f
      11'h689: dout  = 8'b00111111; // 1673 :  63 - 0x3f
      11'h68A: dout  = 8'b01110000; // 1674 : 112 - 0x70
      11'h68B: dout  = 8'b01110001; // 1675 : 113 - 0x71
      11'h68C: dout  = 8'b01110001; // 1676 : 113 - 0x71
      11'h68D: dout  = 8'b01110001; // 1677 : 113 - 0x71
      11'h68E: dout  = 8'b01110001; // 1678 : 113 - 0x71
      11'h68F: dout  = 8'b01110001; // 1679 : 113 - 0x71
      11'h690: dout  = 8'b01110001; // 1680 : 113 - 0x71
      11'h691: dout  = 8'b01110001; // 1681 : 113 - 0x71
      11'h692: dout  = 8'b01110001; // 1682 : 113 - 0x71
      11'h693: dout  = 8'b01110001; // 1683 : 113 - 0x71
      11'h694: dout  = 8'b01110001; // 1684 : 113 - 0x71
      11'h695: dout  = 8'b01110010; // 1685 : 114 - 0x72
      11'h696: dout  = 8'b00111111; // 1686 :  63 - 0x3f
      11'h697: dout  = 8'b00111111; // 1687 :  63 - 0x3f
      11'h698: dout  = 8'b00111111; // 1688 :  63 - 0x3f
      11'h699: dout  = 8'b00111111; // 1689 :  63 - 0x3f
      11'h69A: dout  = 8'b00111111; // 1690 :  63 - 0x3f
      11'h69B: dout  = 8'b00111111; // 1691 :  63 - 0x3f
      11'h69C: dout  = 8'b00111111; // 1692 :  63 - 0x3f
      11'h69D: dout  = 8'b00111111; // 1693 :  63 - 0x3f
      11'h69E: dout  = 8'b00111111; // 1694 :  63 - 0x3f
      11'h69F: dout  = 8'b00111111; // 1695 :  63 - 0x3f
      11'h6A0: dout  = 8'b00111111; // 1696 :  63 - 0x3f -- line 0x15
      11'h6A1: dout  = 8'b00111111; // 1697 :  63 - 0x3f
      11'h6A2: dout  = 8'b00111111; // 1698 :  63 - 0x3f
      11'h6A3: dout  = 8'b00111111; // 1699 :  63 - 0x3f
      11'h6A4: dout  = 8'b00111111; // 1700 :  63 - 0x3f
      11'h6A5: dout  = 8'b00111111; // 1701 :  63 - 0x3f
      11'h6A6: dout  = 8'b00111111; // 1702 :  63 - 0x3f
      11'h6A7: dout  = 8'b00111111; // 1703 :  63 - 0x3f
      11'h6A8: dout  = 8'b00111111; // 1704 :  63 - 0x3f
      11'h6A9: dout  = 8'b00111111; // 1705 :  63 - 0x3f
      11'h6AA: dout  = 8'b01100000; // 1706 :  96 - 0x60
      11'h6AB: dout  = 8'b01110111; // 1707 : 119 - 0x77
      11'h6AC: dout  = 8'b01110111; // 1708 : 119 - 0x77
      11'h6AD: dout  = 8'b01110111; // 1709 : 119 - 0x77
      11'h6AE: dout  = 8'b01110111; // 1710 : 119 - 0x77
      11'h6AF: dout  = 8'b01110111; // 1711 : 119 - 0x77
      11'h6B0: dout  = 8'b01110111; // 1712 : 119 - 0x77
      11'h6B1: dout  = 8'b01110111; // 1713 : 119 - 0x77
      11'h6B2: dout  = 8'b01110111; // 1714 : 119 - 0x77
      11'h6B3: dout  = 8'b01110111; // 1715 : 119 - 0x77
      11'h6B4: dout  = 8'b01110111; // 1716 : 119 - 0x77
      11'h6B5: dout  = 8'b01100001; // 1717 :  97 - 0x61
      11'h6B6: dout  = 8'b00111111; // 1718 :  63 - 0x3f
      11'h6B7: dout  = 8'b00111111; // 1719 :  63 - 0x3f
      11'h6B8: dout  = 8'b00111111; // 1720 :  63 - 0x3f
      11'h6B9: dout  = 8'b00111111; // 1721 :  63 - 0x3f
      11'h6BA: dout  = 8'b00111111; // 1722 :  63 - 0x3f
      11'h6BB: dout  = 8'b00111111; // 1723 :  63 - 0x3f
      11'h6BC: dout  = 8'b00111111; // 1724 :  63 - 0x3f
      11'h6BD: dout  = 8'b00111111; // 1725 :  63 - 0x3f
      11'h6BE: dout  = 8'b00111111; // 1726 :  63 - 0x3f
      11'h6BF: dout  = 8'b00111111; // 1727 :  63 - 0x3f
      11'h6C0: dout  = 8'b00111111; // 1728 :  63 - 0x3f -- line 0x16
      11'h6C1: dout  = 8'b00111111; // 1729 :  63 - 0x3f
      11'h6C2: dout  = 8'b00111111; // 1730 :  63 - 0x3f
      11'h6C3: dout  = 8'b00111111; // 1731 :  63 - 0x3f
      11'h6C4: dout  = 8'b00111111; // 1732 :  63 - 0x3f
      11'h6C5: dout  = 8'b00111111; // 1733 :  63 - 0x3f
      11'h6C6: dout  = 8'b00111111; // 1734 :  63 - 0x3f
      11'h6C7: dout  = 8'b00111111; // 1735 :  63 - 0x3f
      11'h6C8: dout  = 8'b00111111; // 1736 :  63 - 0x3f
      11'h6C9: dout  = 8'b00111111; // 1737 :  63 - 0x3f
      11'h6CA: dout  = 8'b01100000; // 1738 :  96 - 0x60
      11'h6CB: dout  = 8'b01110011; // 1739 : 115 - 0x73
      11'h6CC: dout  = 8'b01110011; // 1740 : 115 - 0x73
      11'h6CD: dout  = 8'b01110011; // 1741 : 115 - 0x73
      11'h6CE: dout  = 8'b01110011; // 1742 : 115 - 0x73
      11'h6CF: dout  = 8'b01110011; // 1743 : 115 - 0x73
      11'h6D0: dout  = 8'b01110011; // 1744 : 115 - 0x73
      11'h6D1: dout  = 8'b01110011; // 1745 : 115 - 0x73
      11'h6D2: dout  = 8'b01110011; // 1746 : 115 - 0x73
      11'h6D3: dout  = 8'b01110011; // 1747 : 115 - 0x73
      11'h6D4: dout  = 8'b01110011; // 1748 : 115 - 0x73
      11'h6D5: dout  = 8'b01100001; // 1749 :  97 - 0x61
      11'h6D6: dout  = 8'b00111111; // 1750 :  63 - 0x3f
      11'h6D7: dout  = 8'b00111111; // 1751 :  63 - 0x3f
      11'h6D8: dout  = 8'b00111111; // 1752 :  63 - 0x3f
      11'h6D9: dout  = 8'b00111111; // 1753 :  63 - 0x3f
      11'h6DA: dout  = 8'b00111111; // 1754 :  63 - 0x3f
      11'h6DB: dout  = 8'b00111111; // 1755 :  63 - 0x3f
      11'h6DC: dout  = 8'b00111111; // 1756 :  63 - 0x3f
      11'h6DD: dout  = 8'b00111111; // 1757 :  63 - 0x3f
      11'h6DE: dout  = 8'b00111111; // 1758 :  63 - 0x3f
      11'h6DF: dout  = 8'b00111111; // 1759 :  63 - 0x3f
      11'h6E0: dout  = 8'b11000101; // 1760 : 197 - 0xc5 -- line 0x17
      11'h6E1: dout  = 8'b11010110; // 1761 : 214 - 0xd6
      11'h6E2: dout  = 8'b00111111; // 1762 :  63 - 0x3f
      11'h6E3: dout  = 8'b00111111; // 1763 :  63 - 0x3f
      11'h6E4: dout  = 8'b00111111; // 1764 :  63 - 0x3f
      11'h6E5: dout  = 8'b00111111; // 1765 :  63 - 0x3f
      11'h6E6: dout  = 8'b00111111; // 1766 :  63 - 0x3f
      11'h6E7: dout  = 8'b00111111; // 1767 :  63 - 0x3f
      11'h6E8: dout  = 8'b00111111; // 1768 :  63 - 0x3f
      11'h6E9: dout  = 8'b00111111; // 1769 :  63 - 0x3f
      11'h6EA: dout  = 8'b01100000; // 1770 :  96 - 0x60
      11'h6EB: dout  = 8'b01110011; // 1771 : 115 - 0x73
      11'h6EC: dout  = 8'b01110011; // 1772 : 115 - 0x73
      11'h6ED: dout  = 8'b01110011; // 1773 : 115 - 0x73
      11'h6EE: dout  = 8'b01110011; // 1774 : 115 - 0x73
      11'h6EF: dout  = 8'b01110011; // 1775 : 115 - 0x73
      11'h6F0: dout  = 8'b01110011; // 1776 : 115 - 0x73
      11'h6F1: dout  = 8'b01110011; // 1777 : 115 - 0x73
      11'h6F2: dout  = 8'b01110011; // 1778 : 115 - 0x73
      11'h6F3: dout  = 8'b01110011; // 1779 : 115 - 0x73
      11'h6F4: dout  = 8'b01110011; // 1780 : 115 - 0x73
      11'h6F5: dout  = 8'b01100001; // 1781 :  97 - 0x61
      11'h6F6: dout  = 8'b00111111; // 1782 :  63 - 0x3f
      11'h6F7: dout  = 8'b00111111; // 1783 :  63 - 0x3f
      11'h6F8: dout  = 8'b00111111; // 1784 :  63 - 0x3f
      11'h6F9: dout  = 8'b00111111; // 1785 :  63 - 0x3f
      11'h6FA: dout  = 8'b00111111; // 1786 :  63 - 0x3f
      11'h6FB: dout  = 8'b00111111; // 1787 :  63 - 0x3f
      11'h6FC: dout  = 8'b00111111; // 1788 :  63 - 0x3f
      11'h6FD: dout  = 8'b00111111; // 1789 :  63 - 0x3f
      11'h6FE: dout  = 8'b00111111; // 1790 :  63 - 0x3f
      11'h6FF: dout  = 8'b00111111; // 1791 :  63 - 0x3f
      11'h700: dout  = 8'b11000111; // 1792 : 199 - 0xc7 -- line 0x18
      11'h701: dout  = 8'b11001001; // 1793 : 201 - 0xc9
      11'h702: dout  = 8'b00111111; // 1794 :  63 - 0x3f
      11'h703: dout  = 8'b00111111; // 1795 :  63 - 0x3f
      11'h704: dout  = 8'b00111111; // 1796 :  63 - 0x3f
      11'h705: dout  = 8'b00111111; // 1797 :  63 - 0x3f
      11'h706: dout  = 8'b00111111; // 1798 :  63 - 0x3f
      11'h707: dout  = 8'b00111111; // 1799 :  63 - 0x3f
      11'h708: dout  = 8'b00111111; // 1800 :  63 - 0x3f
      11'h709: dout  = 8'b00111111; // 1801 :  63 - 0x3f
      11'h70A: dout  = 8'b01100000; // 1802 :  96 - 0x60
      11'h70B: dout  = 8'b01110011; // 1803 : 115 - 0x73
      11'h70C: dout  = 8'b01110011; // 1804 : 115 - 0x73
      11'h70D: dout  = 8'b01110011; // 1805 : 115 - 0x73
      11'h70E: dout  = 8'b01110011; // 1806 : 115 - 0x73
      11'h70F: dout  = 8'b01110011; // 1807 : 115 - 0x73
      11'h710: dout  = 8'b01110011; // 1808 : 115 - 0x73
      11'h711: dout  = 8'b01110011; // 1809 : 115 - 0x73
      11'h712: dout  = 8'b01110011; // 1810 : 115 - 0x73
      11'h713: dout  = 8'b01110011; // 1811 : 115 - 0x73
      11'h714: dout  = 8'b01110011; // 1812 : 115 - 0x73
      11'h715: dout  = 8'b01100001; // 1813 :  97 - 0x61
      11'h716: dout  = 8'b00111111; // 1814 :  63 - 0x3f
      11'h717: dout  = 8'b00111111; // 1815 :  63 - 0x3f
      11'h718: dout  = 8'b00111111; // 1816 :  63 - 0x3f
      11'h719: dout  = 8'b00111111; // 1817 :  63 - 0x3f
      11'h71A: dout  = 8'b00111111; // 1818 :  63 - 0x3f
      11'h71B: dout  = 8'b00111111; // 1819 :  63 - 0x3f
      11'h71C: dout  = 8'b00111111; // 1820 :  63 - 0x3f
      11'h71D: dout  = 8'b00111111; // 1821 :  63 - 0x3f
      11'h71E: dout  = 8'b00111111; // 1822 :  63 - 0x3f
      11'h71F: dout  = 8'b00111111; // 1823 :  63 - 0x3f
      11'h720: dout  = 8'b11010111; // 1824 : 215 - 0xd7 -- line 0x19
      11'h721: dout  = 8'b11011001; // 1825 : 217 - 0xd9
      11'h722: dout  = 8'b00111111; // 1826 :  63 - 0x3f
      11'h723: dout  = 8'b00111111; // 1827 :  63 - 0x3f
      11'h724: dout  = 8'b00111111; // 1828 :  63 - 0x3f
      11'h725: dout  = 8'b00111111; // 1829 :  63 - 0x3f
      11'h726: dout  = 8'b00111111; // 1830 :  63 - 0x3f
      11'h727: dout  = 8'b00111111; // 1831 :  63 - 0x3f
      11'h728: dout  = 8'b00011000; // 1832 :  24 - 0x18
      11'h729: dout  = 8'b00011001; // 1833 :  25 - 0x19
      11'h72A: dout  = 8'b01100000; // 1834 :  96 - 0x60
      11'h72B: dout  = 8'b01110011; // 1835 : 115 - 0x73
      11'h72C: dout  = 8'b01110011; // 1836 : 115 - 0x73
      11'h72D: dout  = 8'b01110011; // 1837 : 115 - 0x73
      11'h72E: dout  = 8'b01110011; // 1838 : 115 - 0x73
      11'h72F: dout  = 8'b01110011; // 1839 : 115 - 0x73
      11'h730: dout  = 8'b01110011; // 1840 : 115 - 0x73
      11'h731: dout  = 8'b01110011; // 1841 : 115 - 0x73
      11'h732: dout  = 8'b01110011; // 1842 : 115 - 0x73
      11'h733: dout  = 8'b01110011; // 1843 : 115 - 0x73
      11'h734: dout  = 8'b01110011; // 1844 : 115 - 0x73
      11'h735: dout  = 8'b01100001; // 1845 :  97 - 0x61
      11'h736: dout  = 8'b00111111; // 1846 :  63 - 0x3f
      11'h737: dout  = 8'b00111111; // 1847 :  63 - 0x3f
      11'h738: dout  = 8'b00111111; // 1848 :  63 - 0x3f
      11'h739: dout  = 8'b00111111; // 1849 :  63 - 0x3f
      11'h73A: dout  = 8'b00111111; // 1850 :  63 - 0x3f
      11'h73B: dout  = 8'b00111111; // 1851 :  63 - 0x3f
      11'h73C: dout  = 8'b00111111; // 1852 :  63 - 0x3f
      11'h73D: dout  = 8'b00111111; // 1853 :  63 - 0x3f
      11'h73E: dout  = 8'b00111111; // 1854 :  63 - 0x3f
      11'h73F: dout  = 8'b00111111; // 1855 :  63 - 0x3f
      11'h740: dout  = 8'b01110001; // 1856 : 113 - 0x71 -- line 0x1a
      11'h741: dout  = 8'b01110001; // 1857 : 113 - 0x71
      11'h742: dout  = 8'b01110001; // 1858 : 113 - 0x71
      11'h743: dout  = 8'b01110001; // 1859 : 113 - 0x71
      11'h744: dout  = 8'b01110001; // 1860 : 113 - 0x71
      11'h745: dout  = 8'b01110001; // 1861 : 113 - 0x71
      11'h746: dout  = 8'b01110001; // 1862 : 113 - 0x71
      11'h747: dout  = 8'b01110001; // 1863 : 113 - 0x71
      11'h748: dout  = 8'b01110001; // 1864 : 113 - 0x71
      11'h749: dout  = 8'b01110001; // 1865 : 113 - 0x71
      11'h74A: dout  = 8'b01100000; // 1866 :  96 - 0x60
      11'h74B: dout  = 8'b01110011; // 1867 : 115 - 0x73
      11'h74C: dout  = 8'b01110011; // 1868 : 115 - 0x73
      11'h74D: dout  = 8'b01110011; // 1869 : 115 - 0x73
      11'h74E: dout  = 8'b01110011; // 1870 : 115 - 0x73
      11'h74F: dout  = 8'b01110011; // 1871 : 115 - 0x73
      11'h750: dout  = 8'b01110011; // 1872 : 115 - 0x73
      11'h751: dout  = 8'b01110011; // 1873 : 115 - 0x73
      11'h752: dout  = 8'b01110011; // 1874 : 115 - 0x73
      11'h753: dout  = 8'b01110011; // 1875 : 115 - 0x73
      11'h754: dout  = 8'b01110011; // 1876 : 115 - 0x73
      11'h755: dout  = 8'b01100001; // 1877 :  97 - 0x61
      11'h756: dout  = 8'b00111111; // 1878 :  63 - 0x3f
      11'h757: dout  = 8'b00111111; // 1879 :  63 - 0x3f
      11'h758: dout  = 8'b00111111; // 1880 :  63 - 0x3f
      11'h759: dout  = 8'b00111111; // 1881 :  63 - 0x3f
      11'h75A: dout  = 8'b00111111; // 1882 :  63 - 0x3f
      11'h75B: dout  = 8'b00111111; // 1883 :  63 - 0x3f
      11'h75C: dout  = 8'b00111111; // 1884 :  63 - 0x3f
      11'h75D: dout  = 8'b00111111; // 1885 :  63 - 0x3f
      11'h75E: dout  = 8'b00111111; // 1886 :  63 - 0x3f
      11'h75F: dout  = 8'b00111111; // 1887 :  63 - 0x3f
      11'h760: dout  = 8'b01110111; // 1888 : 119 - 0x77 -- line 0x1b
      11'h761: dout  = 8'b01110111; // 1889 : 119 - 0x77
      11'h762: dout  = 8'b01110111; // 1890 : 119 - 0x77
      11'h763: dout  = 8'b01110111; // 1891 : 119 - 0x77
      11'h764: dout  = 8'b01110111; // 1892 : 119 - 0x77
      11'h765: dout  = 8'b01110111; // 1893 : 119 - 0x77
      11'h766: dout  = 8'b01110111; // 1894 : 119 - 0x77
      11'h767: dout  = 8'b01110111; // 1895 : 119 - 0x77
      11'h768: dout  = 8'b01110111; // 1896 : 119 - 0x77
      11'h769: dout  = 8'b01110111; // 1897 : 119 - 0x77
      11'h76A: dout  = 8'b01110011; // 1898 : 115 - 0x73
      11'h76B: dout  = 8'b01110011; // 1899 : 115 - 0x73
      11'h76C: dout  = 8'b01110011; // 1900 : 115 - 0x73
      11'h76D: dout  = 8'b01110011; // 1901 : 115 - 0x73
      11'h76E: dout  = 8'b01110011; // 1902 : 115 - 0x73
      11'h76F: dout  = 8'b01110011; // 1903 : 115 - 0x73
      11'h770: dout  = 8'b01110011; // 1904 : 115 - 0x73
      11'h771: dout  = 8'b01110011; // 1905 : 115 - 0x73
      11'h772: dout  = 8'b01110011; // 1906 : 115 - 0x73
      11'h773: dout  = 8'b01110011; // 1907 : 115 - 0x73
      11'h774: dout  = 8'b01110011; // 1908 : 115 - 0x73
      11'h775: dout  = 8'b01100001; // 1909 :  97 - 0x61
      11'h776: dout  = 8'b00111111; // 1910 :  63 - 0x3f
      11'h777: dout  = 8'b00111111; // 1911 :  63 - 0x3f
      11'h778: dout  = 8'b00111111; // 1912 :  63 - 0x3f
      11'h779: dout  = 8'b00111111; // 1913 :  63 - 0x3f
      11'h77A: dout  = 8'b00111111; // 1914 :  63 - 0x3f
      11'h77B: dout  = 8'b00111111; // 1915 :  63 - 0x3f
      11'h77C: dout  = 8'b00111111; // 1916 :  63 - 0x3f
      11'h77D: dout  = 8'b00111111; // 1917 :  63 - 0x3f
      11'h77E: dout  = 8'b00111111; // 1918 :  63 - 0x3f
      11'h77F: dout  = 8'b00111111; // 1919 :  63 - 0x3f
      11'h780: dout  = 8'b01110011; // 1920 : 115 - 0x73 -- line 0x1c
      11'h781: dout  = 8'b01110011; // 1921 : 115 - 0x73
      11'h782: dout  = 8'b01110011; // 1922 : 115 - 0x73
      11'h783: dout  = 8'b01110011; // 1923 : 115 - 0x73
      11'h784: dout  = 8'b01110011; // 1924 : 115 - 0x73
      11'h785: dout  = 8'b01110011; // 1925 : 115 - 0x73
      11'h786: dout  = 8'b01110011; // 1926 : 115 - 0x73
      11'h787: dout  = 8'b01110011; // 1927 : 115 - 0x73
      11'h788: dout  = 8'b01110011; // 1928 : 115 - 0x73
      11'h789: dout  = 8'b01110011; // 1929 : 115 - 0x73
      11'h78A: dout  = 8'b01110011; // 1930 : 115 - 0x73
      11'h78B: dout  = 8'b01110011; // 1931 : 115 - 0x73
      11'h78C: dout  = 8'b01110011; // 1932 : 115 - 0x73
      11'h78D: dout  = 8'b01110011; // 1933 : 115 - 0x73
      11'h78E: dout  = 8'b01110011; // 1934 : 115 - 0x73
      11'h78F: dout  = 8'b01110011; // 1935 : 115 - 0x73
      11'h790: dout  = 8'b01110011; // 1936 : 115 - 0x73
      11'h791: dout  = 8'b01110011; // 1937 : 115 - 0x73
      11'h792: dout  = 8'b01110011; // 1938 : 115 - 0x73
      11'h793: dout  = 8'b01110011; // 1939 : 115 - 0x73
      11'h794: dout  = 8'b01110011; // 1940 : 115 - 0x73
      11'h795: dout  = 8'b01100001; // 1941 :  97 - 0x61
      11'h796: dout  = 8'b00111111; // 1942 :  63 - 0x3f
      11'h797: dout  = 8'b00111111; // 1943 :  63 - 0x3f
      11'h798: dout  = 8'b00111111; // 1944 :  63 - 0x3f
      11'h799: dout  = 8'b00111111; // 1945 :  63 - 0x3f
      11'h79A: dout  = 8'b00111111; // 1946 :  63 - 0x3f
      11'h79B: dout  = 8'b00111111; // 1947 :  63 - 0x3f
      11'h79C: dout  = 8'b00111111; // 1948 :  63 - 0x3f
      11'h79D: dout  = 8'b00111111; // 1949 :  63 - 0x3f
      11'h79E: dout  = 8'b00111111; // 1950 :  63 - 0x3f
      11'h79F: dout  = 8'b00111111; // 1951 :  63 - 0x3f
      11'h7A0: dout  = 8'b01110011; // 1952 : 115 - 0x73 -- line 0x1d
      11'h7A1: dout  = 8'b01110011; // 1953 : 115 - 0x73
      11'h7A2: dout  = 8'b01110011; // 1954 : 115 - 0x73
      11'h7A3: dout  = 8'b01110011; // 1955 : 115 - 0x73
      11'h7A4: dout  = 8'b01110011; // 1956 : 115 - 0x73
      11'h7A5: dout  = 8'b01110011; // 1957 : 115 - 0x73
      11'h7A6: dout  = 8'b01110011; // 1958 : 115 - 0x73
      11'h7A7: dout  = 8'b01110011; // 1959 : 115 - 0x73
      11'h7A8: dout  = 8'b01110011; // 1960 : 115 - 0x73
      11'h7A9: dout  = 8'b01110011; // 1961 : 115 - 0x73
      11'h7AA: dout  = 8'b01110011; // 1962 : 115 - 0x73
      11'h7AB: dout  = 8'b01110011; // 1963 : 115 - 0x73
      11'h7AC: dout  = 8'b01110011; // 1964 : 115 - 0x73
      11'h7AD: dout  = 8'b01110011; // 1965 : 115 - 0x73
      11'h7AE: dout  = 8'b01110011; // 1966 : 115 - 0x73
      11'h7AF: dout  = 8'b01110011; // 1967 : 115 - 0x73
      11'h7B0: dout  = 8'b01110011; // 1968 : 115 - 0x73
      11'h7B1: dout  = 8'b01110011; // 1969 : 115 - 0x73
      11'h7B2: dout  = 8'b01110011; // 1970 : 115 - 0x73
      11'h7B3: dout  = 8'b01110011; // 1971 : 115 - 0x73
      11'h7B4: dout  = 8'b01110011; // 1972 : 115 - 0x73
      11'h7B5: dout  = 8'b01100001; // 1973 :  97 - 0x61
      11'h7B6: dout  = 8'b00111111; // 1974 :  63 - 0x3f
      11'h7B7: dout  = 8'b00111111; // 1975 :  63 - 0x3f
      11'h7B8: dout  = 8'b00111111; // 1976 :  63 - 0x3f
      11'h7B9: dout  = 8'b00111111; // 1977 :  63 - 0x3f
      11'h7BA: dout  = 8'b00111111; // 1978 :  63 - 0x3f
      11'h7BB: dout  = 8'b00111111; // 1979 :  63 - 0x3f
      11'h7BC: dout  = 8'b00111111; // 1980 :  63 - 0x3f
      11'h7BD: dout  = 8'b00111111; // 1981 :  63 - 0x3f
      11'h7BE: dout  = 8'b00111111; // 1982 :  63 - 0x3f
      11'h7BF: dout  = 8'b00111111; // 1983 :  63 - 0x3f
        //-- Attribute Table 1----
      11'h7C0: dout  = 8'b00000000; // 1984 :   0 - 0x0
      11'h7C1: dout  = 8'b00000000; // 1985 :   0 - 0x0
      11'h7C2: dout  = 8'b10001000; // 1986 : 136 - 0x88
      11'h7C3: dout  = 8'b00010001; // 1987 :  17 - 0x11
      11'h7C4: dout  = 8'b00000000; // 1988 :   0 - 0x0
      11'h7C5: dout  = 8'b00000000; // 1989 :   0 - 0x0
      11'h7C6: dout  = 8'b00000000; // 1990 :   0 - 0x0
      11'h7C7: dout  = 8'b00000000; // 1991 :   0 - 0x0
      11'h7C8: dout  = 8'b00001010; // 1992 :  10 - 0xa
      11'h7C9: dout  = 8'b00000010; // 1993 :   2 - 0x2
      11'h7CA: dout  = 8'b10001000; // 1994 : 136 - 0x88
      11'h7CB: dout  = 8'b00010001; // 1995 :  17 - 0x11
      11'h7CC: dout  = 8'b00000000; // 1996 :   0 - 0x0
      11'h7CD: dout  = 8'b00000000; // 1997 :   0 - 0x0
      11'h7CE: dout  = 8'b00000000; // 1998 :   0 - 0x0
      11'h7CF: dout  = 8'b00000000; // 1999 :   0 - 0x0
      11'h7D0: dout  = 8'b01010100; // 2000 :  84 - 0x54
      11'h7D1: dout  = 8'b00000101; // 2001 :   5 - 0x5
      11'h7D2: dout  = 8'b00000101; // 2002 :   5 - 0x5
      11'h7D3: dout  = 8'b00000001; // 2003 :   1 - 0x1
      11'h7D4: dout  = 8'b00000000; // 2004 :   0 - 0x0
      11'h7D5: dout  = 8'b00000000; // 2005 :   0 - 0x0
      11'h7D6: dout  = 8'b10000000; // 2006 : 128 - 0x80
      11'h7D7: dout  = 8'b10100000; // 2007 : 160 - 0xa0
      11'h7D8: dout  = 8'b00000000; // 2008 :   0 - 0x0
      11'h7D9: dout  = 8'b00000000; // 2009 :   0 - 0x0
      11'h7DA: dout  = 8'b00000000; // 2010 :   0 - 0x0
      11'h7DB: dout  = 8'b00000000; // 2011 :   0 - 0x0
      11'h7DC: dout  = 8'b00000000; // 2012 :   0 - 0x0
      11'h7DD: dout  = 8'b00000000; // 2013 :   0 - 0x0
      11'h7DE: dout  = 8'b01010000; // 2014 :  80 - 0x50
      11'h7DF: dout  = 8'b01010000; // 2015 :  80 - 0x50
      11'h7E0: dout  = 8'b00000000; // 2016 :   0 - 0x0
      11'h7E1: dout  = 8'b00000000; // 2017 :   0 - 0x0
      11'h7E2: dout  = 8'b00000000; // 2018 :   0 - 0x0
      11'h7E3: dout  = 8'b00000000; // 2019 :   0 - 0x0
      11'h7E4: dout  = 8'b10000000; // 2020 : 128 - 0x80
      11'h7E5: dout  = 8'b00000000; // 2021 :   0 - 0x0
      11'h7E6: dout  = 8'b00000000; // 2022 :   0 - 0x0
      11'h7E7: dout  = 8'b00000000; // 2023 :   0 - 0x0
      11'h7E8: dout  = 8'b00000000; // 2024 :   0 - 0x0
      11'h7E9: dout  = 8'b00000000; // 2025 :   0 - 0x0
      11'h7EA: dout  = 8'b00000000; // 2026 :   0 - 0x0
      11'h7EB: dout  = 8'b00000000; // 2027 :   0 - 0x0
      11'h7EC: dout  = 8'b00000000; // 2028 :   0 - 0x0
      11'h7ED: dout  = 8'b00000000; // 2029 :   0 - 0x0
      11'h7EE: dout  = 8'b00000000; // 2030 :   0 - 0x0
      11'h7EF: dout  = 8'b00000000; // 2031 :   0 - 0x0
      11'h7F0: dout  = 8'b00000000; // 2032 :   0 - 0x0
      11'h7F1: dout  = 8'b00000000; // 2033 :   0 - 0x0
      11'h7F2: dout  = 8'b00000010; // 2034 :   2 - 0x2
      11'h7F3: dout  = 8'b00000000; // 2035 :   0 - 0x0
      11'h7F4: dout  = 8'b00000000; // 2036 :   0 - 0x0
      11'h7F5: dout  = 8'b00000000; // 2037 :   0 - 0x0
      11'h7F6: dout  = 8'b00000000; // 2038 :   0 - 0x0
      11'h7F7: dout  = 8'b00000000; // 2039 :   0 - 0x0
      11'h7F8: dout  = 8'b00000000; // 2040 :   0 - 0x0
      11'h7F9: dout  = 8'b00000000; // 2041 :   0 - 0x0
      11'h7FA: dout  = 8'b00000000; // 2042 :   0 - 0x0
      11'h7FB: dout  = 8'b00000000; // 2043 :   0 - 0x0
      11'h7FC: dout  = 8'b00000000; // 2044 :   0 - 0x0
      11'h7FD: dout  = 8'b00000000; // 2045 :   0 - 0x0
      11'h7FE: dout  = 8'b00000000; // 2046 :   0 - 0x0
      11'h7FF: dout  = 8'b00000000; // 2047 :   0 - 0x0
    endcase
  end

endmodule
