------- ROM creada automaticamente por ppm2rom -----------
------- Felipe Machado -----------------------------------
------- Departamento de Tecnologia Electronica -----------
------- Universidad Rey Juan Carlos ----------------------
------- http://gtebim.es ---------------------------------
----------------------------------------------------------
--------Datos de la imagen -------------------------------
--- Fichero original    : mario32x32.ppm 
--- Filas    : 32 
--- Columnas : 32 
----------------------------------------------------------
--------Codificacion de la memoria------------------------
--- Palabras de 9 bits
--- De cada palabra hay 3 bits para cada color : "RRRGGGBBB" 512 colores



------ Puertos -------------------------------------------
-- Entradas ----------------------------------------------
--    clk  :  senal de reloj
--    addr :  direccion de la memoria
-- Salidas  ----------------------------------------------
--    dout :  dato de 9 bits de la direccion addr (un ciclo despues)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;
entity ROM_RGB_9b_mario32x32 is
  port (
    clk  : in  std_logic;   -- reloj
    addr : in  std_logic_vector(10-1 downto 0);
    dout : out std_logic_vector(9-1 downto 0) 
  );
end ROM_RGB_9b_mario32x32;


architecture BEHAVIORAL of ROM_RGB_9b_mario32x32 is
  signal addr_int  : natural range 0 to 2**10-1;
  type memostruct is array (natural range<>) of std_logic_vector(9-1 downto 0);
  constant filaimg : memostruct := (
     --"RRRGGGBBB"
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111110110",
       "111100100",
       "111010010",
       "111100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111101101",
       "111001001",
       "111000000",
       "111000000",
       "111000000",
       "111100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "110010010",
       "111000000",
       "111000000",
       "111000001",
       "111001001",
       "111000000",
       "111000000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "110011100",
       "110000000",
       "111001001",
       "111000001",
       "111000001",
       "111001001",
       "111001001",
       "111000000",
       "111100100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111110110",
       "101000000",
       "111001001",
       "111000001",
       "111000001",
       "111000001",
       "111000001",
       "111001001",
       "111000000",
       "110001001",
       "111100101",
       "111011011",
       "111001010",
       "100000000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "101000000",
       "110000000",
       "111000001",
       "111000001",
       "111000001",
       "111000001",
       "111001001",
       "111001001",
       "111000001",
       "111000000",
       "111000000",
       "110000000",
       "010000000",
       "100001001",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111101101",
       "101000000",
       "110001001",
       "111000001",
       "111000001",
       "111000001",
       "111000001",
       "111000001",
       "111000000",
       "111000000",
       "010000000",
       "011001001",
       "010000000",
       "100001001",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "101001001",
       "101000000",
       "110001001",
       "111000001",
       "111001001",
       "111001001",
       "111000001",
       "110000000",
       "110001001",
       "110011010",
       "110101100",
       "110101100",
       "101011011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "101000000",
       "101000001",
       "110000001",
       "110000000",
       "110000000",
       "110000001",
       "101000000",
       "110100011",
       "111111110",
       "111111101",
       "111111111",
       "011100101",
       "111111111",
       "111111111",
       "111110110",
       "111111110",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111110110",
       "100000000",
       "101000000",
       "101001001",
       "100000000",
       "100000000",
       "101011011",
       "011000000",
       "010000000",
       "101001000",
       "110101100",
       "111111110",
       "111111111",
       "010011101",
       "111111110",
       "111101100",
       "111101100",
       "111111110",
       "111111110",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "101000000",
       "101000000",
       "101001001",
       "100000000",
       "100000000",
       "111111110",
       "111111110",
       "111110101",
       "010000000",
       "001000000",
       "011000000",
       "111111110",
       "111111101",
       "001001001",
       "101100011",
       "111100011",
       "111101100",
       "111110101",
       "111110100",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "101000000",
       "101000000",
       "101001001",
       "100000000",
       "101010001",
       "111111111",
       "111110100",
       "111100011",
       "110101100",
       "010000000",
       "110101100",
       "111111111",
       "111111110",
       "001000000",
       "000000000",
       "000000000",
       "101011010",
       "111100011",
       "111101101",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111110110",
       "101000000",
       "101000000",
       "100000000",
       "010000000",
       "111111110",
       "111111111",
       "111111101",
       "111111110",
       "111110101",
       "111111101",
       "111110101",
       "111111101",
       "111111101",
       "100010010",
       "000000000",
       "000000000",
       "110110110",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111110110",
       "101001001",
       "010000000",
       "010000000",
       "100001001",
       "111111101",
       "111111110",
       "111101100",
       "111100011",
       "111101100",
       "111101100",
       "111101100",
       "111101100",
       "111110100",
       "111101100",
       "101101101",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "101101101",
       "011001001",
       "001000000",
       "001000000",
       "001000000",
       "100001000",
       "111011010",
       "111100010",
       "111100011",
       "110100011",
       "111100100",
       "111100011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "110000001",
       "110000000",
       "100001000",
       "100001001",
       "010001010",
       "100010001",
       "111010000",
       "111011001",
       "111110101",
       "111111111",
       "111111111",
       "110111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "101110110",
       "110110111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111110110",
       "111000000",
       "111001001",
       "111000001",
       "101000001",
       "000010110",
       "000010111",
       "100000001",
       "011000001",
       "111000000",
       "111101101",
       "101110111",
       "111111111",
       "110111111",
       "101110110",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100101101",
       "100101110",
       "101110111",
       "110111111",
       "111111111",
       "111111111",
       "111111111",
       "110111111",
       "110000000",
       "111001001",
       "111001001",
       "111001000",
       "111000000",
       "000010111",
       "011110111",
       "010100111",
       "010001101",
       "111110011",
       "101110111",
       "111111111",
       "101101110",
       "100101110",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100101101",
       "011100101",
       "100101110",
       "100101110",
       "110111111",
       "100101110",
       "111111111",
       "101100100",
       "101000000",
       "100001001",
       "101000000",
       "111000000",
       "111000000",
       "001001101",
       "111111010",
       "111111000",
       "000100111",
       "010011100",
       "011100100",
       "110111111",
       "111111111",
       "011101101",
       "100101110",
       "110111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100101110",
       "011100101",
       "100101101",
       "101110110",
       "100101101",
       "111111111",
       "100011100",
       "010000000",
       "101000000",
       "111000000",
       "110001010",
       "010010110",
       "000011111",
       "000010101",
       "110101000",
       "001011111",
       "000001110",
       "011011011",
       "010100101",
       "100101110",
       "100100100",
       "011011011",
       "101110111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100101110",
       "011100101",
       "101110111",
       "111111111",
       "111111111",
       "000000101",
       "000010101",
       "000010110",
       "000011111",
       "000011111",
       "000011111",
       "000010111",
       "000001111",
       "000001111",
       "001011110",
       "111111111",
       "111111111",
       "101101100",
       "111011000",
       "111011000",
       "101011010",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "110110110",
       "111111110",
       "111111111",
       "000000101",
       "000010101",
       "000010101",
       "000010110",
       "000010110",
       "000010110",
       "000010110",
       "000011111",
       "000011111",
       "000010111",
       "101110111",
       "101110111",
       "101010000",
       "110011001",
       "101011001",
       "010000000",
       "111111110",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001000000",
       "000000000",
       "000000100",
       "000010110",
       "000001100",
       "000010101",
       "000010110",
       "000010101",
       "000010110",
       "000011111",
       "000011111",
       "000011111",
       "000011111",
       "000010111",
       "000000101",
       "101010000",
       "101011001",
       "011001000",
       "100010000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "110101101",
       "001000000",
       "011010001",
       "000001100",
       "000010110",
       "000010101",
       "000001100",
       "000010101",
       "000010110",
       "000010110",
       "000010110",
       "000010110",
       "000011110",
       "000011110",
       "000011111",
       "000010111",
       "101010000",
       "100010001",
       "001000000",
       "111110101",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011010010",
       "010000000",
       "001010100",
       "000000011",
       "000010101",
       "000010110",
       "000010101",
       "000010101",
       "000010101",
       "000010101",
       "000010101",
       "000010110",
       "000010110",
       "000010110",
       "000010110",
       "000010111",
       "100010000",
       "010001000",
       "010001000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "011010001",
       "011000000",
       "000010101",
       "000001100",
       "000001011",
       "000001100",
       "000010101",
       "000010101",
       "000010101",
       "000001101",
       "000001100",
       "000001101",
       "000010101",
       "000010101",
       "000010110",
       "000010110",
       "100010000",
       "001000000",
       "110110101",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "001000000",
       "100001000",
       "000001101",
       "000010101",
       "000010101",
       "000001100",
       "000001011",
       "000001011",
       "000000011",
       "010011101",
       "010011110",
       "000000101",
       "000000100",
       "000001100",
       "000010110",
       "001010100",
       "011001000",
       "010000000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "101100011",
       "001000000",
       "100010000",
       "001001011",
       "000010110",
       "000001100",
       "000000100",
       "000000100",
       "000000100",
       "011100101",
       "111111111",
       "111111111",
       "111111111",
       "101110111",
       "001010101",
       "000000101",
       "011001001",
       "001000000",
       "110101101",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "010001000",
       "010000000",
       "100010000",
       "011001000",
       "000000101",
       "010011110",
       "100100110",
       "101110111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100100101",
       "001000000",
       "001000000",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "000000000",
       "011001000",
       "100010001",
       "011000000",
       "110110110",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "100011010",
       "011000000",
       "100001000",
       "101100011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "101100011",
       "101100011",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111",
       "111111111"
        );

begin

  addr_int <= TO_INTEGER(unsigned(addr));

  P_ROM: process (clk)
  begin
    if clk'event and clk='1' then
      dout <= filaimg(addr_int);
    end if;
  end process;

end BEHAVIORAL;

