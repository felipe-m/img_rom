--- Autcmatically generated VHDL ROM from a NES memory file----
---   ATTRIBUTE TABLE SEPARATED FROM NAME TABLE
-- https://wiki.nesdev.com/w/index.php/PPU_attribute_tables


---  Original memory dump file name: pacman_ntable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_ATABLE_PACMAN_00 is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(7-1 downto 0);  --128 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_ATABLE_PACMAN_00;

architecture BEHAVIORAL of ROM_ATABLE_PACMAN_00 is
  signal addr_int  : natural range 0 to 2**7-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
    "01010101", --    0 -  0x0  :   85 - 0x55
    "01010101", --    1 -  0x1  :   85 - 0x55
    "01010101", --    2 -  0x2  :   85 - 0x55
    "01010101", --    3 -  0x3  :   85 - 0x55
    "01010101", --    4 -  0x4  :   85 - 0x55
    "00010001", --    5 -  0x5  :   17 - 0x11
    "00000000", --    6 -  0x6  :    0 - 0x0
    "00000000", --    7 -  0x7  :    0 - 0x0
    "01010101", --    8 -  0x8  :   85 - 0x55
    "01010101", --    9 -  0x9  :   85 - 0x55
    "01010101", --   10 -  0xa  :   85 - 0x55
    "01010101", --   11 -  0xb  :   85 - 0x55
    "01010101", --   12 -  0xc  :   85 - 0x55
    "00010001", --   13 -  0xd  :   17 - 0x11
    "00000000", --   14 -  0xe  :    0 - 0x0
    "00000000", --   15 -  0xf  :    0 - 0x0
    "01010101", --   16 - 0x10  :   85 - 0x55
    "01010101", --   17 - 0x11  :   85 - 0x55
    "01010101", --   18 - 0x12  :   85 - 0x55
    "01010101", --   19 - 0x13  :   85 - 0x55
    "01010101", --   20 - 0x14  :   85 - 0x55
    "00010001", --   21 - 0x15  :   17 - 0x11
    "00000000", --   22 - 0x16  :    0 - 0x0
    "00000000", --   23 - 0x17  :    0 - 0x0
    "01010101", --   24 - 0x18  :   85 - 0x55
    "01010101", --   25 - 0x19  :   85 - 0x55
    "01010101", --   26 - 0x1a  :   85 - 0x55
    "01010101", --   27 - 0x1b  :   85 - 0x55
    "01010101", --   28 - 0x1c  :   85 - 0x55
    "01010001", --   29 - 0x1d  :   81 - 0x51
    "01010000", --   30 - 0x1e  :   80 - 0x50
    "01010000", --   31 - 0x1f  :   80 - 0x50
    "01010101", --   32 - 0x20  :   85 - 0x55
    "01010101", --   33 - 0x21  :   85 - 0x55
    "01010101", --   34 - 0x22  :   85 - 0x55
    "01010101", --   35 - 0x23  :   85 - 0x55
    "01010101", --   36 - 0x24  :   85 - 0x55
    "10010101", --   37 - 0x25  :  149 - 0x95
    "00000101", --   38 - 0x26  :    5 - 0x5
    "00000101", --   39 - 0x27  :    5 - 0x5
    "01010101", --   40 - 0x28  :   85 - 0x55
    "01010101", --   41 - 0x29  :   85 - 0x55
    "01010101", --   42 - 0x2a  :   85 - 0x55
    "01010101", --   43 - 0x2b  :   85 - 0x55
    "01010101", --   44 - 0x2c  :   85 - 0x55
    "00010001", --   45 - 0x2d  :   17 - 0x11
    "00000000", --   46 - 0x2e  :    0 - 0x0
    "00000000", --   47 - 0x2f  :    0 - 0x0
    "01010101", --   48 - 0x30  :   85 - 0x55
    "01010101", --   49 - 0x31  :   85 - 0x55
    "01010101", --   50 - 0x32  :   85 - 0x55
    "01010101", --   51 - 0x33  :   85 - 0x55
    "01010101", --   52 - 0x34  :   85 - 0x55
    "01010101", --   53 - 0x35  :   85 - 0x55
    "01010101", --   54 - 0x36  :   85 - 0x55
    "01010101", --   55 - 0x37  :   85 - 0x55
    "01010101", --   56 - 0x38  :   85 - 0x55
    "01010101", --   57 - 0x39  :   85 - 0x55
    "01010101", --   58 - 0x3a  :   85 - 0x55
    "01010101", --   59 - 0x3b  :   85 - 0x55
    "01010101", --   60 - 0x3c  :   85 - 0x55
    "01010101", --   61 - 0x3d  :   85 - 0x55
    "01010101", --   62 - 0x3e  :   85 - 0x55
    "01010101", --   63 - 0x3f  :   85 - 0x55
    "01010101", --   64 - 0x40  :   85 - 0x55
    "01010101", --   65 - 0x41  :   85 - 0x55
    "01010101", --   66 - 0x42  :   85 - 0x55
    "01010101", --   67 - 0x43  :   85 - 0x55
    "01010101", --   68 - 0x44  :   85 - 0x55
    "00010001", --   69 - 0x45  :   17 - 0x11
    "00000000", --   70 - 0x46  :    0 - 0x0
    "00000000", --   71 - 0x47  :    0 - 0x0
    "01010101", --   72 - 0x48  :   85 - 0x55
    "01010101", --   73 - 0x49  :   85 - 0x55
    "01010101", --   74 - 0x4a  :   85 - 0x55
    "01010101", --   75 - 0x4b  :   85 - 0x55
    "01010101", --   76 - 0x4c  :   85 - 0x55
    "00010001", --   77 - 0x4d  :   17 - 0x11
    "00000000", --   78 - 0x4e  :    0 - 0x0
    "00000000", --   79 - 0x4f  :    0 - 0x0
    "01010101", --   80 - 0x50  :   85 - 0x55
    "01010101", --   81 - 0x51  :   85 - 0x55
    "01010101", --   82 - 0x52  :   85 - 0x55
    "01010101", --   83 - 0x53  :   85 - 0x55
    "01010101", --   84 - 0x54  :   85 - 0x55
    "00010001", --   85 - 0x55  :   17 - 0x11
    "00000000", --   86 - 0x56  :    0 - 0x0
    "00000000", --   87 - 0x57  :    0 - 0x0
    "01010101", --   88 - 0x58  :   85 - 0x55
    "01010101", --   89 - 0x59  :   85 - 0x55
    "01010101", --   90 - 0x5a  :   85 - 0x55
    "01010101", --   91 - 0x5b  :   85 - 0x55
    "01010101", --   92 - 0x5c  :   85 - 0x55
    "01010001", --   93 - 0x5d  :   81 - 0x51
    "01010000", --   94 - 0x5e  :   80 - 0x50
    "01010000", --   95 - 0x5f  :   80 - 0x50
    "01010101", --   96 - 0x60  :   85 - 0x55
    "01010101", --   97 - 0x61  :   85 - 0x55
    "01010101", --   98 - 0x62  :   85 - 0x55
    "01010101", --   99 - 0x63  :   85 - 0x55
    "01010101", --  100 - 0x64  :   85 - 0x55
    "00010001", --  101 - 0x65  :   17 - 0x11
    "00000101", --  102 - 0x66  :    5 - 0x5
    "00000101", --  103 - 0x67  :    5 - 0x5
    "01010101", --  104 - 0x68  :   85 - 0x55
    "01010101", --  105 - 0x69  :   85 - 0x55
    "01010101", --  106 - 0x6a  :   85 - 0x55
    "01010101", --  107 - 0x6b  :   85 - 0x55
    "01010101", --  108 - 0x6c  :   85 - 0x55
    "00010001", --  109 - 0x6d  :   17 - 0x11
    "00000000", --  110 - 0x6e  :    0 - 0x0
    "00000000", --  111 - 0x6f  :    0 - 0x0
    "01010101", --  112 - 0x70  :   85 - 0x55
    "01010101", --  113 - 0x71  :   85 - 0x55
    "01010101", --  114 - 0x72  :   85 - 0x55
    "01010101", --  115 - 0x73  :   85 - 0x55
    "01010101", --  116 - 0x74  :   85 - 0x55
    "01010101", --  117 - 0x75  :   85 - 0x55
    "01010101", --  118 - 0x76  :   85 - 0x55
    "01010101", --  119 - 0x77  :   85 - 0x55
    "01010101", --  120 - 0x78  :   85 - 0x55
    "01010101", --  121 - 0x79  :   85 - 0x55
    "01010101", --  122 - 0x7a  :   85 - 0x55
    "01010101", --  123 - 0x7b  :   85 - 0x55
    "01010101", --  124 - 0x7c  :   85 - 0x55
    "01010101", --  125 - 0x7d  :   85 - 0x55
    "01010101", --  126 - 0x7e  :   85 - 0x55
    "01010101"  --  127 - 0x7f  :   85 - 0x55
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
