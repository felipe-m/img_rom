//- Autcmatically generated verilog ROM from a NES memory file----
//-   PATTERN TABLE WITH ONLY ONE COLOR PLANE
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


//-  Original memory dump file name: nova_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_PTABLE_NOVA_color1
  (
     //input     clk,   // clock
     input      [12-1:0] addr,  //4096 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                              //  address:   value 
                              //    dec  : dec - hex
          // Sprite pattern Table
      12'h0: dout  = 8'b00000000; //    0 :   0 - 0x0 -- Sprite 0x0
      12'h1: dout  = 8'b00000000; //    1 :   0 - 0x0
      12'h2: dout  = 8'b00000011; //    2 :   3 - 0x3
      12'h3: dout  = 8'b00000001; //    3 :   1 - 0x1
      12'h4: dout  = 8'b00000001; //    4 :   1 - 0x1
      12'h5: dout  = 8'b00000000; //    5 :   0 - 0x0
      12'h6: dout  = 8'b00000011; //    6 :   3 - 0x3
      12'h7: dout  = 8'b00000001; //    7 :   1 - 0x1
      12'h8: dout  = 8'b00000000; //    8 :   0 - 0x0 -- Sprite 0x1
      12'h9: dout  = 8'b00000000; //    9 :   0 - 0x0
      12'hA: dout  = 8'b00111000; //   10 :  56 - 0x38
      12'hB: dout  = 8'b10110100; //   11 : 180 - 0xb4
      12'hC: dout  = 8'b10101000; //   12 : 168 - 0xa8
      12'hD: dout  = 8'b11010100; //   13 : 212 - 0xd4
      12'hE: dout  = 8'b01110100; //   14 : 116 - 0x74
      12'hF: dout  = 8'b01111110; //   15 : 126 - 0x7e
      12'h10: dout  = 8'b00111000; //   16 :  56 - 0x38 -- Sprite 0x2
      12'h11: dout  = 8'b01111000; //   17 : 120 - 0x78
      12'h12: dout  = 8'b01111100; //   18 : 124 - 0x7c
      12'h13: dout  = 8'b01111110; //   19 : 126 - 0x7e
      12'h14: dout  = 8'b01111110; //   20 : 126 - 0x7e
      12'h15: dout  = 8'b01111110; //   21 : 126 - 0x7e
      12'h16: dout  = 8'b00111110; //   22 :  62 - 0x3e
      12'h17: dout  = 8'b00011110; //   23 :  30 - 0x1e
      12'h18: dout  = 8'b11110110; //   24 : 246 - 0xf6 -- Sprite 0x3
      12'h19: dout  = 8'b11110000; //   25 : 240 - 0xf0
      12'h1A: dout  = 8'b00111000; //   26 :  56 - 0x38
      12'h1B: dout  = 8'b11010000; //   27 : 208 - 0xd0
      12'h1C: dout  = 8'b11100000; //   28 : 224 - 0xe0
      12'h1D: dout  = 8'b01110000; //   29 : 112 - 0x70
      12'h1E: dout  = 8'b10111000; //   30 : 184 - 0xb8
      12'h1F: dout  = 8'b01000000; //   31 :  64 - 0x40
      12'h20: dout  = 8'b00011100; //   32 :  28 - 0x1c -- Sprite 0x4
      12'h21: dout  = 8'b00011100; //   33 :  28 - 0x1c
      12'h22: dout  = 8'b00011110; //   34 :  30 - 0x1e
      12'h23: dout  = 8'b00011111; //   35 :  31 - 0x1f
      12'h24: dout  = 8'b00001100; //   36 :  12 - 0xc
      12'h25: dout  = 8'b00000000; //   37 :   0 - 0x0
      12'h26: dout  = 8'b00000000; //   38 :   0 - 0x0
      12'h27: dout  = 8'b00000000; //   39 :   0 - 0x0
      12'h28: dout  = 8'b10101000; //   40 : 168 - 0xa8 -- Sprite 0x5
      12'h29: dout  = 8'b01010000; //   41 :  80 - 0x50
      12'h2A: dout  = 8'b10101000; //   42 : 168 - 0xa8
      12'h2B: dout  = 8'b00000000; //   43 :   0 - 0x0
      12'h2C: dout  = 8'b01100000; //   44 :  96 - 0x60
      12'h2D: dout  = 8'b01100000; //   45 :  96 - 0x60
      12'h2E: dout  = 8'b01110000; //   46 : 112 - 0x70
      12'h2F: dout  = 8'b00000000; //   47 :   0 - 0x0
      12'h30: dout  = 8'b00011100; //   48 :  28 - 0x1c -- Sprite 0x6
      12'h31: dout  = 8'b00011100; //   49 :  28 - 0x1c
      12'h32: dout  = 8'b00011110; //   50 :  30 - 0x1e
      12'h33: dout  = 8'b00011111; //   51 :  31 - 0x1f
      12'h34: dout  = 8'b00001100; //   52 :  12 - 0xc
      12'h35: dout  = 8'b00000000; //   53 :   0 - 0x0
      12'h36: dout  = 8'b00000001; //   54 :   1 - 0x1
      12'h37: dout  = 8'b00000000; //   55 :   0 - 0x0
      12'h38: dout  = 8'b10101000; //   56 : 168 - 0xa8 -- Sprite 0x7
      12'h39: dout  = 8'b01010000; //   57 :  80 - 0x50
      12'h3A: dout  = 8'b10101000; //   58 : 168 - 0xa8
      12'h3B: dout  = 8'b00000000; //   59 :   0 - 0x0
      12'h3C: dout  = 8'b01011000; //   60 :  88 - 0x58
      12'h3D: dout  = 8'b11011000; //   61 : 216 - 0xd8
      12'h3E: dout  = 8'b10001100; //   62 : 140 - 0x8c
      12'h3F: dout  = 8'b00000000; //   63 :   0 - 0x0
      12'h40: dout  = 8'b00011100; //   64 :  28 - 0x1c -- Sprite 0x8
      12'h41: dout  = 8'b00011100; //   65 :  28 - 0x1c
      12'h42: dout  = 8'b00011110; //   66 :  30 - 0x1e
      12'h43: dout  = 8'b00011111; //   67 :  31 - 0x1f
      12'h44: dout  = 8'b00001100; //   68 :  12 - 0xc
      12'h45: dout  = 8'b00000000; //   69 :   0 - 0x0
      12'h46: dout  = 8'b00000000; //   70 :   0 - 0x0
      12'h47: dout  = 8'b00000000; //   71 :   0 - 0x0
      12'h48: dout  = 8'b10101000; //   72 : 168 - 0xa8 -- Sprite 0x9
      12'h49: dout  = 8'b01010100; //   73 :  84 - 0x54
      12'h4A: dout  = 8'b10101000; //   74 : 168 - 0xa8
      12'h4B: dout  = 8'b00000000; //   75 :   0 - 0x0
      12'h4C: dout  = 8'b01101110; //   76 : 110 - 0x6e
      12'h4D: dout  = 8'b11000000; //   77 : 192 - 0xc0
      12'h4E: dout  = 8'b10000000; //   78 : 128 - 0x80
      12'h4F: dout  = 8'b00000000; //   79 :   0 - 0x0
      12'h50: dout  = 8'b00011100; //   80 :  28 - 0x1c -- Sprite 0xa
      12'h51: dout  = 8'b00011100; //   81 :  28 - 0x1c
      12'h52: dout  = 8'b00011110; //   82 :  30 - 0x1e
      12'h53: dout  = 8'b00011111; //   83 :  31 - 0x1f
      12'h54: dout  = 8'b00001100; //   84 :  12 - 0xc
      12'h55: dout  = 8'b00000001; //   85 :   1 - 0x1
      12'h56: dout  = 8'b00000000; //   86 :   0 - 0x0
      12'h57: dout  = 8'b00000000; //   87 :   0 - 0x0
      12'h58: dout  = 8'b10101000; //   88 : 168 - 0xa8 -- Sprite 0xb
      12'h59: dout  = 8'b01010100; //   89 :  84 - 0x54
      12'h5A: dout  = 8'b10101000; //   90 : 168 - 0xa8
      12'h5B: dout  = 8'b00000000; //   91 :   0 - 0x0
      12'h5C: dout  = 8'b11011000; //   92 : 216 - 0xd8
      12'h5D: dout  = 8'b11011100; //   93 : 220 - 0xdc
      12'h5E: dout  = 8'b00001100; //   94 :  12 - 0xc
      12'h5F: dout  = 8'b00000000; //   95 :   0 - 0x0
      12'h60: dout  = 8'b11110110; //   96 : 246 - 0xf6 -- Sprite 0xc
      12'h61: dout  = 8'b11110000; //   97 : 240 - 0xf0
      12'h62: dout  = 8'b00000000; //   98 :   0 - 0x0
      12'h63: dout  = 8'b11111100; //   99 : 252 - 0xfc
      12'h64: dout  = 8'b11111000; //  100 : 248 - 0xf8
      12'h65: dout  = 8'b00000000; //  101 :   0 - 0x0
      12'h66: dout  = 8'b10101000; //  102 : 168 - 0xa8
      12'h67: dout  = 8'b01010100; //  103 :  84 - 0x54
      12'h68: dout  = 8'b00111000; //  104 :  56 - 0x38 -- Sprite 0xd
      12'h69: dout  = 8'b01111000; //  105 : 120 - 0x78
      12'h6A: dout  = 8'b01111100; //  106 : 124 - 0x7c
      12'h6B: dout  = 8'b01111101; //  107 : 125 - 0x7d
      12'h6C: dout  = 8'b01111101; //  108 : 125 - 0x7d
      12'h6D: dout  = 8'b01111011; //  109 : 123 - 0x7b
      12'h6E: dout  = 8'b00111011; //  110 :  59 - 0x3b
      12'h6F: dout  = 8'b00011011; //  111 :  27 - 0x1b
      12'h70: dout  = 8'b11110110; //  112 : 246 - 0xf6 -- Sprite 0xe
      12'h71: dout  = 8'b11110000; //  113 : 240 - 0xf0
      12'h72: dout  = 8'b01111000; //  114 : 120 - 0x78
      12'h73: dout  = 8'b01110000; //  115 : 112 - 0x70
      12'h74: dout  = 8'b10100000; //  116 : 160 - 0xa0
      12'h75: dout  = 8'b10010000; //  117 : 144 - 0x90
      12'h76: dout  = 8'b00101000; //  118 :  40 - 0x28
      12'h77: dout  = 8'b01010100; //  119 :  84 - 0x54
      12'h78: dout  = 8'b00000000; //  120 :   0 - 0x0 -- Sprite 0xf
      12'h79: dout  = 8'b00000000; //  121 :   0 - 0x0
      12'h7A: dout  = 8'b00000011; //  122 :   3 - 0x3
      12'h7B: dout  = 8'b00000001; //  123 :   1 - 0x1
      12'h7C: dout  = 8'b00000001; //  124 :   1 - 0x1
      12'h7D: dout  = 8'b00000000; //  125 :   0 - 0x0
      12'h7E: dout  = 8'b00000011; //  126 :   3 - 0x3
      12'h7F: dout  = 8'b00000001; //  127 :   1 - 0x1
      12'h80: dout  = 8'b00000000; //  128 :   0 - 0x0 -- Sprite 0x10
      12'h81: dout  = 8'b00000011; //  129 :   3 - 0x3
      12'h82: dout  = 8'b00001111; //  130 :  15 - 0xf
      12'h83: dout  = 8'b00001111; //  131 :  15 - 0xf
      12'h84: dout  = 8'b00001111; //  132 :  15 - 0xf
      12'h85: dout  = 8'b00011111; //  133 :  31 - 0x1f
      12'h86: dout  = 8'b00011111; //  134 :  31 - 0x1f
      12'h87: dout  = 8'b00011110; //  135 :  30 - 0x1e
      12'h88: dout  = 8'b00110110; //  136 :  54 - 0x36 -- Sprite 0x11
      12'h89: dout  = 8'b10110000; //  137 : 176 - 0xb0
      12'h8A: dout  = 8'b10111000; //  138 : 184 - 0xb8
      12'h8B: dout  = 8'b10010000; //  139 : 144 - 0x90
      12'h8C: dout  = 8'b10100000; //  140 : 160 - 0xa0
      12'h8D: dout  = 8'b01110000; //  141 : 112 - 0x70
      12'h8E: dout  = 8'b00111000; //  142 :  56 - 0x38
      12'h8F: dout  = 8'b01000000; //  143 :  64 - 0x40
      12'h90: dout  = 8'b00011100; //  144 :  28 - 0x1c -- Sprite 0x12
      12'h91: dout  = 8'b00011100; //  145 :  28 - 0x1c
      12'h92: dout  = 8'b00011110; //  146 :  30 - 0x1e
      12'h93: dout  = 8'b00011111; //  147 :  31 - 0x1f
      12'h94: dout  = 8'b00001100; //  148 :  12 - 0xc
      12'h95: dout  = 8'b00000000; //  149 :   0 - 0x0
      12'h96: dout  = 8'b00000000; //  150 :   0 - 0x0
      12'h97: dout  = 8'b00000000; //  151 :   0 - 0x0
      12'h98: dout  = 8'b00000000; //  152 :   0 - 0x0 -- Sprite 0x13
      12'h99: dout  = 8'b00000000; //  153 :   0 - 0x0
      12'h9A: dout  = 8'b00000000; //  154 :   0 - 0x0
      12'h9B: dout  = 8'b00000011; //  155 :   3 - 0x3
      12'h9C: dout  = 8'b00000111; //  156 :   7 - 0x7
      12'h9D: dout  = 8'b00001111; //  157 :  15 - 0xf
      12'h9E: dout  = 8'b00001111; //  158 :  15 - 0xf
      12'h9F: dout  = 8'b00011111; //  159 :  31 - 0x1f
      12'hA0: dout  = 8'b11110110; //  160 : 246 - 0xf6 -- Sprite 0x14
      12'hA1: dout  = 8'b00000000; //  161 :   0 - 0x0
      12'hA2: dout  = 8'b11111000; //  162 : 248 - 0xf8
      12'hA3: dout  = 8'b11111110; //  163 : 254 - 0xfe
      12'hA4: dout  = 8'b11111110; //  164 : 254 - 0xfe
      12'hA5: dout  = 8'b11111110; //  165 : 254 - 0xfe
      12'hA6: dout  = 8'b11111000; //  166 : 248 - 0xf8
      12'hA7: dout  = 8'b00000000; //  167 :   0 - 0x0
      12'hA8: dout  = 8'b00000011; //  168 :   3 - 0x3 -- Sprite 0x15
      12'hA9: dout  = 8'b00000011; //  169 :   3 - 0x3
      12'hAA: dout  = 8'b00000000; //  170 :   0 - 0x0
      12'hAB: dout  = 8'b00000011; //  171 :   3 - 0x3
      12'hAC: dout  = 8'b00000011; //  172 :   3 - 0x3
      12'hAD: dout  = 8'b00000000; //  173 :   0 - 0x0
      12'hAE: dout  = 8'b00001111; //  174 :  15 - 0xf
      12'hAF: dout  = 8'b00111111; //  175 :  63 - 0x3f
      12'hB0: dout  = 8'b11011000; //  176 : 216 - 0xd8 -- Sprite 0x16
      12'hB1: dout  = 8'b11000000; //  177 : 192 - 0xc0
      12'hB2: dout  = 8'b11100000; //  178 : 224 - 0xe0
      12'hB3: dout  = 8'b01000000; //  179 :  64 - 0x40
      12'hB4: dout  = 8'b10000000; //  180 : 128 - 0x80
      12'hB5: dout  = 8'b00000000; //  181 :   0 - 0x0
      12'hB6: dout  = 8'b11100000; //  182 : 224 - 0xe0
      12'hB7: dout  = 8'b11111100; //  183 : 252 - 0xfc
      12'hB8: dout  = 8'b01111111; //  184 : 127 - 0x7f -- Sprite 0x17
      12'hB9: dout  = 8'b01111111; //  185 : 127 - 0x7f
      12'hBA: dout  = 8'b01111111; //  186 : 127 - 0x7f
      12'hBB: dout  = 8'b01111100; //  187 : 124 - 0x7c
      12'hBC: dout  = 8'b00110000; //  188 :  48 - 0x30
      12'hBD: dout  = 8'b00000001; //  189 :   1 - 0x1
      12'hBE: dout  = 8'b00000001; //  190 :   1 - 0x1
      12'hBF: dout  = 8'b00000000; //  191 :   0 - 0x0
      12'hC0: dout  = 8'b11111100; //  192 : 252 - 0xfc -- Sprite 0x18
      12'hC1: dout  = 8'b11111110; //  193 : 254 - 0xfe
      12'hC2: dout  = 8'b11111100; //  194 : 252 - 0xfc
      12'hC3: dout  = 8'b00000000; //  195 :   0 - 0x0
      12'hC4: dout  = 8'b00000000; //  196 :   0 - 0x0
      12'hC5: dout  = 8'b10000000; //  197 : 128 - 0x80
      12'hC6: dout  = 8'b11000000; //  198 : 192 - 0xc0
      12'hC7: dout  = 8'b00000000; //  199 :   0 - 0x0
      12'hC8: dout  = 8'b00000111; //  200 :   7 - 0x7 -- Sprite 0x19
      12'hC9: dout  = 8'b00000111; //  201 :   7 - 0x7
      12'hCA: dout  = 8'b00000001; //  202 :   1 - 0x1
      12'hCB: dout  = 8'b00000110; //  203 :   6 - 0x6
      12'hCC: dout  = 8'b00000111; //  204 :   7 - 0x7
      12'hCD: dout  = 8'b00000110; //  205 :   6 - 0x6
      12'hCE: dout  = 8'b00000000; //  206 :   0 - 0x0
      12'hCF: dout  = 8'b00001111; //  207 :  15 - 0xf
      12'hD0: dout  = 8'b10110000; //  208 : 176 - 0xb0 -- Sprite 0x1a
      12'hD1: dout  = 8'b10000000; //  209 : 128 - 0x80
      12'hD2: dout  = 8'b11000000; //  210 : 192 - 0xc0
      12'hD3: dout  = 8'b10000000; //  211 : 128 - 0x80
      12'hD4: dout  = 8'b00000000; //  212 :   0 - 0x0
      12'hD5: dout  = 8'b00000000; //  213 :   0 - 0x0
      12'hD6: dout  = 8'b00000000; //  214 :   0 - 0x0
      12'hD7: dout  = 8'b11100000; //  215 : 224 - 0xe0
      12'hD8: dout  = 8'b00111111; //  216 :  63 - 0x3f -- Sprite 0x1b
      12'hD9: dout  = 8'b00111111; //  217 :  63 - 0x3f
      12'hDA: dout  = 8'b01111111; //  218 : 127 - 0x7f
      12'hDB: dout  = 8'b01111111; //  219 : 127 - 0x7f
      12'hDC: dout  = 8'b00111111; //  220 :  63 - 0x3f
      12'hDD: dout  = 8'b00000000; //  221 :   0 - 0x0
      12'hDE: dout  = 8'b00000011; //  222 :   3 - 0x3
      12'hDF: dout  = 8'b00000000; //  223 :   0 - 0x0
      12'hE0: dout  = 8'b11111111; //  224 : 255 - 0xff -- Sprite 0x1c
      12'hE1: dout  = 8'b11111111; //  225 : 255 - 0xff
      12'hE2: dout  = 8'b11111111; //  226 : 255 - 0xff
      12'hE3: dout  = 8'b11111111; //  227 : 255 - 0xff
      12'hE4: dout  = 8'b11111111; //  228 : 255 - 0xff
      12'hE5: dout  = 8'b00000000; //  229 :   0 - 0x0
      12'hE6: dout  = 8'b10000000; //  230 : 128 - 0x80
      12'hE7: dout  = 8'b00000000; //  231 :   0 - 0x0
      12'hE8: dout  = 8'b00000000; //  232 :   0 - 0x0 -- Sprite 0x1d
      12'hE9: dout  = 8'b11000000; //  233 : 192 - 0xc0
      12'hEA: dout  = 8'b11000000; //  234 : 192 - 0xc0
      12'hEB: dout  = 8'b11000000; //  235 : 192 - 0xc0
      12'hEC: dout  = 8'b10000000; //  236 : 128 - 0x80
      12'hED: dout  = 8'b00000000; //  237 :   0 - 0x0
      12'hEE: dout  = 8'b00000000; //  238 :   0 - 0x0
      12'hEF: dout  = 8'b00000000; //  239 :   0 - 0x0
      12'hF0: dout  = 8'b11100000; //  240 : 224 - 0xe0 -- Sprite 0x1e
      12'hF1: dout  = 8'b10011100; //  241 : 156 - 0x9c
      12'hF2: dout  = 8'b00111000; //  242 :  56 - 0x38
      12'hF3: dout  = 8'b11100000; //  243 : 224 - 0xe0
      12'hF4: dout  = 8'b11001000; //  244 : 200 - 0xc8
      12'hF5: dout  = 8'b00010100; //  245 :  20 - 0x14
      12'hF6: dout  = 8'b10101000; //  246 : 168 - 0xa8
      12'hF7: dout  = 8'b01010100; //  247 :  84 - 0x54
      12'hF8: dout  = 8'b00000000; //  248 :   0 - 0x0 -- Sprite 0x1f
      12'hF9: dout  = 8'b00000000; //  249 :   0 - 0x0
      12'hFA: dout  = 8'b00111000; //  250 :  56 - 0x38
      12'hFB: dout  = 8'b10110100; //  251 : 180 - 0xb4
      12'hFC: dout  = 8'b10101000; //  252 : 168 - 0xa8
      12'hFD: dout  = 8'b11010100; //  253 : 212 - 0xd4
      12'hFE: dout  = 8'b01110100; //  254 : 116 - 0x74
      12'hFF: dout  = 8'b00011110; //  255 :  30 - 0x1e
      12'h100: dout  = 8'b00000000; //  256 :   0 - 0x0 -- Sprite 0x20
      12'h101: dout  = 8'b00000000; //  257 :   0 - 0x0
      12'h102: dout  = 8'b00001100; //  258 :  12 - 0xc
      12'h103: dout  = 8'b00000111; //  259 :   7 - 0x7
      12'h104: dout  = 8'b00001111; //  260 :  15 - 0xf
      12'h105: dout  = 8'b00000111; //  261 :   7 - 0x7
      12'h106: dout  = 8'b00001111; //  262 :  15 - 0xf
      12'h107: dout  = 8'b00001111; //  263 :  15 - 0xf
      12'h108: dout  = 8'b00000000; //  264 :   0 - 0x0 -- Sprite 0x21
      12'h109: dout  = 8'b00000000; //  265 :   0 - 0x0
      12'h10A: dout  = 8'b00110000; //  266 :  48 - 0x30
      12'h10B: dout  = 8'b11100000; //  267 : 224 - 0xe0
      12'h10C: dout  = 8'b11110000; //  268 : 240 - 0xf0
      12'h10D: dout  = 8'b11100000; //  269 : 224 - 0xe0
      12'h10E: dout  = 8'b11110000; //  270 : 240 - 0xf0
      12'h10F: dout  = 8'b11110000; //  271 : 240 - 0xf0
      12'h110: dout  = 8'b00000111; //  272 :   7 - 0x7 -- Sprite 0x22
      12'h111: dout  = 8'b00000011; //  273 :   3 - 0x3
      12'h112: dout  = 8'b00011000; //  274 :  24 - 0x18
      12'h113: dout  = 8'b00010101; //  275 :  21 - 0x15
      12'h114: dout  = 8'b00000010; //  276 :   2 - 0x2
      12'h115: dout  = 8'b00000101; //  277 :   5 - 0x5
      12'h116: dout  = 8'b00000010; //  278 :   2 - 0x2
      12'h117: dout  = 8'b00000100; //  279 :   4 - 0x4
      12'h118: dout  = 8'b11100000; //  280 : 224 - 0xe0 -- Sprite 0x23
      12'h119: dout  = 8'b11000000; //  281 : 192 - 0xc0
      12'h11A: dout  = 8'b00111100; //  282 :  60 - 0x3c
      12'h11B: dout  = 8'b01111100; //  283 : 124 - 0x7c
      12'h11C: dout  = 8'b01111100; //  284 : 124 - 0x7c
      12'h11D: dout  = 8'b01111100; //  285 : 124 - 0x7c
      12'h11E: dout  = 8'b11101100; //  286 : 236 - 0xec
      12'h11F: dout  = 8'b11100000; //  287 : 224 - 0xe0
      12'h120: dout  = 8'b00000010; //  288 :   2 - 0x2 -- Sprite 0x24
      12'h121: dout  = 8'b00000101; //  289 :   5 - 0x5
      12'h122: dout  = 8'b00001011; //  290 :  11 - 0xb
      12'h123: dout  = 8'b00001011; //  291 :  11 - 0xb
      12'h124: dout  = 8'b00001101; //  292 :  13 - 0xd
      12'h125: dout  = 8'b00011000; //  293 :  24 - 0x18
      12'h126: dout  = 8'b00111000; //  294 :  56 - 0x38
      12'h127: dout  = 8'b00000000; //  295 :   0 - 0x0
      12'h128: dout  = 8'b11100000; //  296 : 224 - 0xe0 -- Sprite 0x25
      12'h129: dout  = 8'b11100000; //  297 : 224 - 0xe0
      12'h12A: dout  = 8'b11100000; //  298 : 224 - 0xe0
      12'h12B: dout  = 8'b11010000; //  299 : 208 - 0xd0
      12'h12C: dout  = 8'b10111000; //  300 : 184 - 0xb8
      12'h12D: dout  = 8'b00111000; //  301 :  56 - 0x38
      12'h12E: dout  = 8'b00000000; //  302 :   0 - 0x0
      12'h12F: dout  = 8'b00000000; //  303 :   0 - 0x0
      12'h130: dout  = 8'b00000000; //  304 :   0 - 0x0 -- Sprite 0x26
      12'h131: dout  = 8'b00000000; //  305 :   0 - 0x0
      12'h132: dout  = 8'b00000000; //  306 :   0 - 0x0
      12'h133: dout  = 8'b00000000; //  307 :   0 - 0x0
      12'h134: dout  = 8'b00000000; //  308 :   0 - 0x0
      12'h135: dout  = 8'b00000000; //  309 :   0 - 0x0
      12'h136: dout  = 8'b00000000; //  310 :   0 - 0x0
      12'h137: dout  = 8'b00000000; //  311 :   0 - 0x0
      12'h138: dout  = 8'b00000000; //  312 :   0 - 0x0 -- Sprite 0x27
      12'h139: dout  = 8'b00000000; //  313 :   0 - 0x0
      12'h13A: dout  = 8'b00000000; //  314 :   0 - 0x0
      12'h13B: dout  = 8'b00000000; //  315 :   0 - 0x0
      12'h13C: dout  = 8'b00000000; //  316 :   0 - 0x0
      12'h13D: dout  = 8'b00000000; //  317 :   0 - 0x0
      12'h13E: dout  = 8'b00000000; //  318 :   0 - 0x0
      12'h13F: dout  = 8'b00000000; //  319 :   0 - 0x0
      12'h140: dout  = 8'b00000000; //  320 :   0 - 0x0 -- Sprite 0x28
      12'h141: dout  = 8'b00000000; //  321 :   0 - 0x0
      12'h142: dout  = 8'b00000000; //  322 :   0 - 0x0
      12'h143: dout  = 8'b00000000; //  323 :   0 - 0x0
      12'h144: dout  = 8'b00000000; //  324 :   0 - 0x0
      12'h145: dout  = 8'b00000000; //  325 :   0 - 0x0
      12'h146: dout  = 8'b00000000; //  326 :   0 - 0x0
      12'h147: dout  = 8'b00000000; //  327 :   0 - 0x0
      12'h148: dout  = 8'b00011111; //  328 :  31 - 0x1f -- Sprite 0x29
      12'h149: dout  = 8'b00011111; //  329 :  31 - 0x1f
      12'h14A: dout  = 8'b00011111; //  330 :  31 - 0x1f
      12'h14B: dout  = 8'b00011111; //  331 :  31 - 0x1f
      12'h14C: dout  = 8'b00001100; //  332 :  12 - 0xc
      12'h14D: dout  = 8'b00000000; //  333 :   0 - 0x0
      12'h14E: dout  = 8'b00000001; //  334 :   1 - 0x1
      12'h14F: dout  = 8'b00000000; //  335 :   0 - 0x0
      12'h150: dout  = 8'b00011111; //  336 :  31 - 0x1f -- Sprite 0x2a
      12'h151: dout  = 8'b00011111; //  337 :  31 - 0x1f
      12'h152: dout  = 8'b00011111; //  338 :  31 - 0x1f
      12'h153: dout  = 8'b00011111; //  339 :  31 - 0x1f
      12'h154: dout  = 8'b00001100; //  340 :  12 - 0xc
      12'h155: dout  = 8'b00000000; //  341 :   0 - 0x0
      12'h156: dout  = 8'b00000000; //  342 :   0 - 0x0
      12'h157: dout  = 8'b00000000; //  343 :   0 - 0x0
      12'h158: dout  = 8'b00000000; //  344 :   0 - 0x0 -- Sprite 0x2b
      12'h159: dout  = 8'b00000000; //  345 :   0 - 0x0
      12'h15A: dout  = 8'b00000000; //  346 :   0 - 0x0
      12'h15B: dout  = 8'b00000000; //  347 :   0 - 0x0
      12'h15C: dout  = 8'b00000000; //  348 :   0 - 0x0
      12'h15D: dout  = 8'b00000000; //  349 :   0 - 0x0
      12'h15E: dout  = 8'b00000000; //  350 :   0 - 0x0
      12'h15F: dout  = 8'b00000000; //  351 :   0 - 0x0
      12'h160: dout  = 8'b00000000; //  352 :   0 - 0x0 -- Sprite 0x2c
      12'h161: dout  = 8'b00000000; //  353 :   0 - 0x0
      12'h162: dout  = 8'b00000000; //  354 :   0 - 0x0
      12'h163: dout  = 8'b00000000; //  355 :   0 - 0x0
      12'h164: dout  = 8'b00000000; //  356 :   0 - 0x0
      12'h165: dout  = 8'b00000000; //  357 :   0 - 0x0
      12'h166: dout  = 8'b00000000; //  358 :   0 - 0x0
      12'h167: dout  = 8'b00000000; //  359 :   0 - 0x0
      12'h168: dout  = 8'b00000000; //  360 :   0 - 0x0 -- Sprite 0x2d
      12'h169: dout  = 8'b01111110; //  361 : 126 - 0x7e
      12'h16A: dout  = 8'b01000010; //  362 :  66 - 0x42
      12'h16B: dout  = 8'b01000010; //  363 :  66 - 0x42
      12'h16C: dout  = 8'b01000010; //  364 :  66 - 0x42
      12'h16D: dout  = 8'b01000010; //  365 :  66 - 0x42
      12'h16E: dout  = 8'b01111110; //  366 : 126 - 0x7e
      12'h16F: dout  = 8'b00000000; //  367 :   0 - 0x0
      12'h170: dout  = 8'b00000000; //  368 :   0 - 0x0 -- Sprite 0x2e
      12'h171: dout  = 8'b00000000; //  369 :   0 - 0x0
      12'h172: dout  = 8'b00000000; //  370 :   0 - 0x0
      12'h173: dout  = 8'b00000000; //  371 :   0 - 0x0
      12'h174: dout  = 8'b00000000; //  372 :   0 - 0x0
      12'h175: dout  = 8'b00000000; //  373 :   0 - 0x0
      12'h176: dout  = 8'b00000000; //  374 :   0 - 0x0
      12'h177: dout  = 8'b00000000; //  375 :   0 - 0x0
      12'h178: dout  = 8'b01100110; //  376 : 102 - 0x66 -- Sprite 0x2f
      12'h179: dout  = 8'b01100000; //  377 :  96 - 0x60
      12'h17A: dout  = 8'b01101000; //  378 : 104 - 0x68
      12'h17B: dout  = 8'b11100000; //  379 : 224 - 0xe0
      12'h17C: dout  = 8'b11000000; //  380 : 192 - 0xc0
      12'h17D: dout  = 8'b00010000; //  381 :  16 - 0x10
      12'h17E: dout  = 8'b00101000; //  382 :  40 - 0x28
      12'h17F: dout  = 8'b01010000; //  383 :  80 - 0x50
      12'h180: dout  = 8'b11110110; //  384 : 246 - 0xf6 -- Sprite 0x30
      12'h181: dout  = 8'b11110000; //  385 : 240 - 0xf0
      12'h182: dout  = 8'b00111000; //  386 :  56 - 0x38
      12'h183: dout  = 8'b11010000; //  387 : 208 - 0xd0
      12'h184: dout  = 8'b11000000; //  388 : 192 - 0xc0
      12'h185: dout  = 8'b11111000; //  389 : 248 - 0xf8
      12'h186: dout  = 8'b01111000; //  390 : 120 - 0x78
      12'h187: dout  = 8'b00000000; //  391 :   0 - 0x0
      12'h188: dout  = 8'b11110110; //  392 : 246 - 0xf6 -- Sprite 0x31
      12'h189: dout  = 8'b11110000; //  393 : 240 - 0xf0
      12'h18A: dout  = 8'b00111000; //  394 :  56 - 0x38
      12'h18B: dout  = 8'b11010000; //  395 : 208 - 0xd0
      12'h18C: dout  = 8'b11000000; //  396 : 192 - 0xc0
      12'h18D: dout  = 8'b11100000; //  397 : 224 - 0xe0
      12'h18E: dout  = 8'b01111000; //  398 : 120 - 0x78
      12'h18F: dout  = 8'b00111000; //  399 :  56 - 0x38
      12'h190: dout  = 8'b11110110; //  400 : 246 - 0xf6 -- Sprite 0x32
      12'h191: dout  = 8'b11110000; //  401 : 240 - 0xf0
      12'h192: dout  = 8'b00111000; //  402 :  56 - 0x38
      12'h193: dout  = 8'b11000000; //  403 : 192 - 0xc0
      12'h194: dout  = 8'b11011000; //  404 : 216 - 0xd8
      12'h195: dout  = 8'b11111000; //  405 : 248 - 0xf8
      12'h196: dout  = 8'b01100000; //  406 :  96 - 0x60
      12'h197: dout  = 8'b00010000; //  407 :  16 - 0x10
      12'h198: dout  = 8'b00011100; //  408 :  28 - 0x1c -- Sprite 0x33
      12'h199: dout  = 8'b00011100; //  409 :  28 - 0x1c
      12'h19A: dout  = 8'b00011110; //  410 :  30 - 0x1e
      12'h19B: dout  = 8'b00011111; //  411 :  31 - 0x1f
      12'h19C: dout  = 8'b00001100; //  412 :  12 - 0xc
      12'h19D: dout  = 8'b00000000; //  413 :   0 - 0x0
      12'h19E: dout  = 8'b00000000; //  414 :   0 - 0x0
      12'h19F: dout  = 8'b00000000; //  415 :   0 - 0x0
      12'h1A0: dout  = 8'b10000000; //  416 : 128 - 0x80 -- Sprite 0x34
      12'h1A1: dout  = 8'b01010000; //  417 :  80 - 0x50
      12'h1A2: dout  = 8'b10101000; //  418 : 168 - 0xa8
      12'h1A3: dout  = 8'b00000000; //  419 :   0 - 0x0
      12'h1A4: dout  = 8'b01011000; //  420 :  88 - 0x58
      12'h1A5: dout  = 8'b11011000; //  421 : 216 - 0xd8
      12'h1A6: dout  = 8'b11101100; //  422 : 236 - 0xec
      12'h1A7: dout  = 8'b00000000; //  423 :   0 - 0x0
      12'h1A8: dout  = 8'b00011100; //  424 :  28 - 0x1c -- Sprite 0x35
      12'h1A9: dout  = 8'b00011100; //  425 :  28 - 0x1c
      12'h1AA: dout  = 8'b00011110; //  426 :  30 - 0x1e
      12'h1AB: dout  = 8'b00011111; //  427 :  31 - 0x1f
      12'h1AC: dout  = 8'b00001100; //  428 :  12 - 0xc
      12'h1AD: dout  = 8'b00000001; //  429 :   1 - 0x1
      12'h1AE: dout  = 8'b00000001; //  430 :   1 - 0x1
      12'h1AF: dout  = 8'b00000000; //  431 :   0 - 0x0
      12'h1B0: dout  = 8'b10101000; //  432 : 168 - 0xa8 -- Sprite 0x36
      12'h1B1: dout  = 8'b01010000; //  433 :  80 - 0x50
      12'h1B2: dout  = 8'b10101000; //  434 : 168 - 0xa8
      12'h1B3: dout  = 8'b00000000; //  435 :   0 - 0x0
      12'h1B4: dout  = 8'b01011000; //  436 :  88 - 0x58
      12'h1B5: dout  = 8'b11001110; //  437 : 206 - 0xce
      12'h1B6: dout  = 8'b10000110; //  438 : 134 - 0x86
      12'h1B7: dout  = 8'b00000000; //  439 :   0 - 0x0
      12'h1B8: dout  = 8'b10101000; //  440 : 168 - 0xa8 -- Sprite 0x37
      12'h1B9: dout  = 8'b01010000; //  441 :  80 - 0x50
      12'h1BA: dout  = 8'b10101000; //  442 : 168 - 0xa8
      12'h1BB: dout  = 8'b00000000; //  443 :   0 - 0x0
      12'h1BC: dout  = 8'b01011000; //  444 :  88 - 0x58
      12'h1BD: dout  = 8'b11011000; //  445 : 216 - 0xd8
      12'h1BE: dout  = 8'b11101100; //  446 : 236 - 0xec
      12'h1BF: dout  = 8'b00000000; //  447 :   0 - 0x0
      12'h1C0: dout  = 8'b00000000; //  448 :   0 - 0x0 -- Sprite 0x38
      12'h1C1: dout  = 8'b00000000; //  449 :   0 - 0x0
      12'h1C2: dout  = 8'b00000000; //  450 :   0 - 0x0
      12'h1C3: dout  = 8'b00000000; //  451 :   0 - 0x0
      12'h1C4: dout  = 8'b00000000; //  452 :   0 - 0x0
      12'h1C5: dout  = 8'b00000000; //  453 :   0 - 0x0
      12'h1C6: dout  = 8'b00000000; //  454 :   0 - 0x0
      12'h1C7: dout  = 8'b00000000; //  455 :   0 - 0x0
      12'h1C8: dout  = 8'b00000000; //  456 :   0 - 0x0 -- Sprite 0x39
      12'h1C9: dout  = 8'b00000000; //  457 :   0 - 0x0
      12'h1CA: dout  = 8'b00000000; //  458 :   0 - 0x0
      12'h1CB: dout  = 8'b00000000; //  459 :   0 - 0x0
      12'h1CC: dout  = 8'b00000000; //  460 :   0 - 0x0
      12'h1CD: dout  = 8'b00000000; //  461 :   0 - 0x0
      12'h1CE: dout  = 8'b00000000; //  462 :   0 - 0x0
      12'h1CF: dout  = 8'b00000000; //  463 :   0 - 0x0
      12'h1D0: dout  = 8'b00000000; //  464 :   0 - 0x0 -- Sprite 0x3a
      12'h1D1: dout  = 8'b00000000; //  465 :   0 - 0x0
      12'h1D2: dout  = 8'b00000000; //  466 :   0 - 0x0
      12'h1D3: dout  = 8'b00000000; //  467 :   0 - 0x0
      12'h1D4: dout  = 8'b00000000; //  468 :   0 - 0x0
      12'h1D5: dout  = 8'b00000000; //  469 :   0 - 0x0
      12'h1D6: dout  = 8'b00000000; //  470 :   0 - 0x0
      12'h1D7: dout  = 8'b00000000; //  471 :   0 - 0x0
      12'h1D8: dout  = 8'b00000000; //  472 :   0 - 0x0 -- Sprite 0x3b
      12'h1D9: dout  = 8'b00000000; //  473 :   0 - 0x0
      12'h1DA: dout  = 8'b00000000; //  474 :   0 - 0x0
      12'h1DB: dout  = 8'b00000000; //  475 :   0 - 0x0
      12'h1DC: dout  = 8'b00000000; //  476 :   0 - 0x0
      12'h1DD: dout  = 8'b00000000; //  477 :   0 - 0x0
      12'h1DE: dout  = 8'b00000000; //  478 :   0 - 0x0
      12'h1DF: dout  = 8'b00000000; //  479 :   0 - 0x0
      12'h1E0: dout  = 8'b00000000; //  480 :   0 - 0x0 -- Sprite 0x3c
      12'h1E1: dout  = 8'b00000000; //  481 :   0 - 0x0
      12'h1E2: dout  = 8'b00000000; //  482 :   0 - 0x0
      12'h1E3: dout  = 8'b00000000; //  483 :   0 - 0x0
      12'h1E4: dout  = 8'b00000000; //  484 :   0 - 0x0
      12'h1E5: dout  = 8'b00000000; //  485 :   0 - 0x0
      12'h1E6: dout  = 8'b00000000; //  486 :   0 - 0x0
      12'h1E7: dout  = 8'b00000000; //  487 :   0 - 0x0
      12'h1E8: dout  = 8'b00000000; //  488 :   0 - 0x0 -- Sprite 0x3d
      12'h1E9: dout  = 8'b00000000; //  489 :   0 - 0x0
      12'h1EA: dout  = 8'b00000000; //  490 :   0 - 0x0
      12'h1EB: dout  = 8'b00000000; //  491 :   0 - 0x0
      12'h1EC: dout  = 8'b00000000; //  492 :   0 - 0x0
      12'h1ED: dout  = 8'b00000000; //  493 :   0 - 0x0
      12'h1EE: dout  = 8'b00000000; //  494 :   0 - 0x0
      12'h1EF: dout  = 8'b00000000; //  495 :   0 - 0x0
      12'h1F0: dout  = 8'b00000000; //  496 :   0 - 0x0 -- Sprite 0x3e
      12'h1F1: dout  = 8'b00000000; //  497 :   0 - 0x0
      12'h1F2: dout  = 8'b00000000; //  498 :   0 - 0x0
      12'h1F3: dout  = 8'b00000000; //  499 :   0 - 0x0
      12'h1F4: dout  = 8'b00000000; //  500 :   0 - 0x0
      12'h1F5: dout  = 8'b00000000; //  501 :   0 - 0x0
      12'h1F6: dout  = 8'b00000000; //  502 :   0 - 0x0
      12'h1F7: dout  = 8'b00000000; //  503 :   0 - 0x0
      12'h1F8: dout  = 8'b00000000; //  504 :   0 - 0x0 -- Sprite 0x3f
      12'h1F9: dout  = 8'b00000000; //  505 :   0 - 0x0
      12'h1FA: dout  = 8'b00000000; //  506 :   0 - 0x0
      12'h1FB: dout  = 8'b00000000; //  507 :   0 - 0x0
      12'h1FC: dout  = 8'b00000000; //  508 :   0 - 0x0
      12'h1FD: dout  = 8'b00000000; //  509 :   0 - 0x0
      12'h1FE: dout  = 8'b00000000; //  510 :   0 - 0x0
      12'h1FF: dout  = 8'b00000000; //  511 :   0 - 0x0
      12'h200: dout  = 8'b00111100; //  512 :  60 - 0x3c -- Sprite 0x40
      12'h201: dout  = 8'b01111100; //  513 : 124 - 0x7c
      12'h202: dout  = 8'b11100110; //  514 : 230 - 0xe6
      12'h203: dout  = 8'b11101110; //  515 : 238 - 0xee
      12'h204: dout  = 8'b11110110; //  516 : 246 - 0xf6
      12'h205: dout  = 8'b11100110; //  517 : 230 - 0xe6
      12'h206: dout  = 8'b00111100; //  518 :  60 - 0x3c
      12'h207: dout  = 8'b00000000; //  519 :   0 - 0x0
      12'h208: dout  = 8'b00111000; //  520 :  56 - 0x38 -- Sprite 0x41
      12'h209: dout  = 8'b01111000; //  521 : 120 - 0x78
      12'h20A: dout  = 8'b00111000; //  522 :  56 - 0x38
      12'h20B: dout  = 8'b00111000; //  523 :  56 - 0x38
      12'h20C: dout  = 8'b00111000; //  524 :  56 - 0x38
      12'h20D: dout  = 8'b00111000; //  525 :  56 - 0x38
      12'h20E: dout  = 8'b00111000; //  526 :  56 - 0x38
      12'h20F: dout  = 8'b00000000; //  527 :   0 - 0x0
      12'h210: dout  = 8'b01111100; //  528 : 124 - 0x7c -- Sprite 0x42
      12'h211: dout  = 8'b11111110; //  529 : 254 - 0xfe
      12'h212: dout  = 8'b11100110; //  530 : 230 - 0xe6
      12'h213: dout  = 8'b00011110; //  531 :  30 - 0x1e
      12'h214: dout  = 8'b01111100; //  532 : 124 - 0x7c
      12'h215: dout  = 8'b11100000; //  533 : 224 - 0xe0
      12'h216: dout  = 8'b11111110; //  534 : 254 - 0xfe
      12'h217: dout  = 8'b00000000; //  535 :   0 - 0x0
      12'h218: dout  = 8'b01111100; //  536 : 124 - 0x7c -- Sprite 0x43
      12'h219: dout  = 8'b11111100; //  537 : 252 - 0xfc
      12'h21A: dout  = 8'b11100110; //  538 : 230 - 0xe6
      12'h21B: dout  = 8'b00011100; //  539 :  28 - 0x1c
      12'h21C: dout  = 8'b01100110; //  540 : 102 - 0x66
      12'h21D: dout  = 8'b11101110; //  541 : 238 - 0xee
      12'h21E: dout  = 8'b11111100; //  542 : 252 - 0xfc
      12'h21F: dout  = 8'b00000000; //  543 :   0 - 0x0
      12'h220: dout  = 8'b00001100; //  544 :  12 - 0xc -- Sprite 0x44
      12'h221: dout  = 8'b00011100; //  545 :  28 - 0x1c
      12'h222: dout  = 8'b00111100; //  546 :  60 - 0x3c
      12'h223: dout  = 8'b01111100; //  547 : 124 - 0x7c
      12'h224: dout  = 8'b11101100; //  548 : 236 - 0xec
      12'h225: dout  = 8'b11111110; //  549 : 254 - 0xfe
      12'h226: dout  = 8'b00001100; //  550 :  12 - 0xc
      12'h227: dout  = 8'b00000000; //  551 :   0 - 0x0
      12'h228: dout  = 8'b11111110; //  552 : 254 - 0xfe -- Sprite 0x45
      12'h229: dout  = 8'b11111110; //  553 : 254 - 0xfe
      12'h22A: dout  = 8'b11100000; //  554 : 224 - 0xe0
      12'h22B: dout  = 8'b11111110; //  555 : 254 - 0xfe
      12'h22C: dout  = 8'b00000110; //  556 :   6 - 0x6
      12'h22D: dout  = 8'b11101110; //  557 : 238 - 0xee
      12'h22E: dout  = 8'b11111100; //  558 : 252 - 0xfc
      12'h22F: dout  = 8'b00000000; //  559 :   0 - 0x0
      12'h230: dout  = 8'b00111100; //  560 :  60 - 0x3c -- Sprite 0x46
      12'h231: dout  = 8'b01111100; //  561 : 124 - 0x7c
      12'h232: dout  = 8'b11100000; //  562 : 224 - 0xe0
      12'h233: dout  = 8'b11111110; //  563 : 254 - 0xfe
      12'h234: dout  = 8'b11100110; //  564 : 230 - 0xe6
      12'h235: dout  = 8'b11101110; //  565 : 238 - 0xee
      12'h236: dout  = 8'b00111100; //  566 :  60 - 0x3c
      12'h237: dout  = 8'b00000000; //  567 :   0 - 0x0
      12'h238: dout  = 8'b11111110; //  568 : 254 - 0xfe -- Sprite 0x47
      12'h239: dout  = 8'b11111100; //  569 : 252 - 0xfc
      12'h23A: dout  = 8'b00001100; //  570 :  12 - 0xc
      12'h23B: dout  = 8'b00111000; //  571 :  56 - 0x38
      12'h23C: dout  = 8'b00111000; //  572 :  56 - 0x38
      12'h23D: dout  = 8'b01110000; //  573 : 112 - 0x70
      12'h23E: dout  = 8'b01110000; //  574 : 112 - 0x70
      12'h23F: dout  = 8'b00000000; //  575 :   0 - 0x0
      12'h240: dout  = 8'b00111110; //  576 :  62 - 0x3e -- Sprite 0x48
      12'h241: dout  = 8'b01111100; //  577 : 124 - 0x7c
      12'h242: dout  = 8'b11100110; //  578 : 230 - 0xe6
      12'h243: dout  = 8'b10111100; //  579 : 188 - 0xbc
      12'h244: dout  = 8'b11100110; //  580 : 230 - 0xe6
      12'h245: dout  = 8'b11101110; //  581 : 238 - 0xee
      12'h246: dout  = 8'b00111100; //  582 :  60 - 0x3c
      12'h247: dout  = 8'b00000000; //  583 :   0 - 0x0
      12'h248: dout  = 8'b00111100; //  584 :  60 - 0x3c -- Sprite 0x49
      12'h249: dout  = 8'b01111100; //  585 : 124 - 0x7c
      12'h24A: dout  = 8'b11100110; //  586 : 230 - 0xe6
      12'h24B: dout  = 8'b11101110; //  587 : 238 - 0xee
      12'h24C: dout  = 8'b11111110; //  588 : 254 - 0xfe
      12'h24D: dout  = 8'b10000110; //  589 : 134 - 0x86
      12'h24E: dout  = 8'b01111100; //  590 : 124 - 0x7c
      12'h24F: dout  = 8'b01000000; //  591 :  64 - 0x40
      12'h250: dout  = 8'b11101110; //  592 : 238 - 0xee -- Sprite 0x4a
      12'h251: dout  = 8'b11101110; //  593 : 238 - 0xee
      12'h252: dout  = 8'b11101110; //  594 : 238 - 0xee
      12'h253: dout  = 8'b11101110; //  595 : 238 - 0xee
      12'h254: dout  = 8'b11101110; //  596 : 238 - 0xee
      12'h255: dout  = 8'b11101110; //  597 : 238 - 0xee
      12'h256: dout  = 8'b11101110; //  598 : 238 - 0xee
      12'h257: dout  = 8'b10001000; //  599 : 136 - 0x88
      12'h258: dout  = 8'b11100000; //  600 : 224 - 0xe0 -- Sprite 0x4b
      12'h259: dout  = 8'b11100000; //  601 : 224 - 0xe0
      12'h25A: dout  = 8'b11100000; //  602 : 224 - 0xe0
      12'h25B: dout  = 8'b11100000; //  603 : 224 - 0xe0
      12'h25C: dout  = 8'b11100000; //  604 : 224 - 0xe0
      12'h25D: dout  = 8'b11100000; //  605 : 224 - 0xe0
      12'h25E: dout  = 8'b11100000; //  606 : 224 - 0xe0
      12'h25F: dout  = 8'b10000000; //  607 : 128 - 0x80
      12'h260: dout  = 8'b00000000; //  608 :   0 - 0x0 -- Sprite 0x4c
      12'h261: dout  = 8'b01111111; //  609 : 127 - 0x7f
      12'h262: dout  = 8'b01111111; //  610 : 127 - 0x7f
      12'h263: dout  = 8'b01111111; //  611 : 127 - 0x7f
      12'h264: dout  = 8'b01111111; //  612 : 127 - 0x7f
      12'h265: dout  = 8'b01111111; //  613 : 127 - 0x7f
      12'h266: dout  = 8'b01111111; //  614 : 127 - 0x7f
      12'h267: dout  = 8'b01111111; //  615 : 127 - 0x7f
      12'h268: dout  = 8'b01111111; //  616 : 127 - 0x7f -- Sprite 0x4d
      12'h269: dout  = 8'b01111111; //  617 : 127 - 0x7f
      12'h26A: dout  = 8'b01111111; //  618 : 127 - 0x7f
      12'h26B: dout  = 8'b01111111; //  619 : 127 - 0x7f
      12'h26C: dout  = 8'b01111111; //  620 : 127 - 0x7f
      12'h26D: dout  = 8'b01111111; //  621 : 127 - 0x7f
      12'h26E: dout  = 8'b01111111; //  622 : 127 - 0x7f
      12'h26F: dout  = 8'b00000000; //  623 :   0 - 0x0
      12'h270: dout  = 8'b00000000; //  624 :   0 - 0x0 -- Sprite 0x4e
      12'h271: dout  = 8'b11111110; //  625 : 254 - 0xfe
      12'h272: dout  = 8'b11111110; //  626 : 254 - 0xfe
      12'h273: dout  = 8'b11111110; //  627 : 254 - 0xfe
      12'h274: dout  = 8'b11111110; //  628 : 254 - 0xfe
      12'h275: dout  = 8'b11111110; //  629 : 254 - 0xfe
      12'h276: dout  = 8'b11111110; //  630 : 254 - 0xfe
      12'h277: dout  = 8'b11111110; //  631 : 254 - 0xfe
      12'h278: dout  = 8'b11111110; //  632 : 254 - 0xfe -- Sprite 0x4f
      12'h279: dout  = 8'b11111110; //  633 : 254 - 0xfe
      12'h27A: dout  = 8'b11111110; //  634 : 254 - 0xfe
      12'h27B: dout  = 8'b11111110; //  635 : 254 - 0xfe
      12'h27C: dout  = 8'b11111110; //  636 : 254 - 0xfe
      12'h27D: dout  = 8'b11111110; //  637 : 254 - 0xfe
      12'h27E: dout  = 8'b11111110; //  638 : 254 - 0xfe
      12'h27F: dout  = 8'b00000000; //  639 :   0 - 0x0
      12'h280: dout  = 8'b00000000; //  640 :   0 - 0x0 -- Sprite 0x50
      12'h281: dout  = 8'b00000000; //  641 :   0 - 0x0
      12'h282: dout  = 8'b00000000; //  642 :   0 - 0x0
      12'h283: dout  = 8'b00000000; //  643 :   0 - 0x0
      12'h284: dout  = 8'b00000000; //  644 :   0 - 0x0
      12'h285: dout  = 8'b00000000; //  645 :   0 - 0x0
      12'h286: dout  = 8'b00000000; //  646 :   0 - 0x0
      12'h287: dout  = 8'b00000000; //  647 :   0 - 0x0
      12'h288: dout  = 8'b00000000; //  648 :   0 - 0x0 -- Sprite 0x51
      12'h289: dout  = 8'b00010000; //  649 :  16 - 0x10
      12'h28A: dout  = 8'b00010000; //  650 :  16 - 0x10
      12'h28B: dout  = 8'b01111100; //  651 : 124 - 0x7c
      12'h28C: dout  = 8'b00111000; //  652 :  56 - 0x38
      12'h28D: dout  = 8'b00111000; //  653 :  56 - 0x38
      12'h28E: dout  = 8'b01101100; //  654 : 108 - 0x6c
      12'h28F: dout  = 8'b00000000; //  655 :   0 - 0x0
      12'h290: dout  = 8'b00000000; //  656 :   0 - 0x0 -- Sprite 0x52
      12'h291: dout  = 8'b00010000; //  657 :  16 - 0x10
      12'h292: dout  = 8'b00010000; //  658 :  16 - 0x10
      12'h293: dout  = 8'b01111100; //  659 : 124 - 0x7c
      12'h294: dout  = 8'b00111000; //  660 :  56 - 0x38
      12'h295: dout  = 8'b00111000; //  661 :  56 - 0x38
      12'h296: dout  = 8'b01101100; //  662 : 108 - 0x6c
      12'h297: dout  = 8'b00000000; //  663 :   0 - 0x0
      12'h298: dout  = 8'b00000000; //  664 :   0 - 0x0 -- Sprite 0x53
      12'h299: dout  = 8'b00000000; //  665 :   0 - 0x0
      12'h29A: dout  = 8'b00000000; //  666 :   0 - 0x0
      12'h29B: dout  = 8'b00000000; //  667 :   0 - 0x0
      12'h29C: dout  = 8'b00000000; //  668 :   0 - 0x0
      12'h29D: dout  = 8'b00000000; //  669 :   0 - 0x0
      12'h29E: dout  = 8'b00000000; //  670 :   0 - 0x0
      12'h29F: dout  = 8'b00000000; //  671 :   0 - 0x0
      12'h2A0: dout  = 8'b11111111; //  672 : 255 - 0xff -- Sprite 0x54
      12'h2A1: dout  = 8'b11111111; //  673 : 255 - 0xff
      12'h2A2: dout  = 8'b11111111; //  674 : 255 - 0xff
      12'h2A3: dout  = 8'b11111111; //  675 : 255 - 0xff
      12'h2A4: dout  = 8'b11111111; //  676 : 255 - 0xff
      12'h2A5: dout  = 8'b11111111; //  677 : 255 - 0xff
      12'h2A6: dout  = 8'b11111111; //  678 : 255 - 0xff
      12'h2A7: dout  = 8'b11111111; //  679 : 255 - 0xff
      12'h2A8: dout  = 8'b11111111; //  680 : 255 - 0xff -- Sprite 0x55
      12'h2A9: dout  = 8'b11111111; //  681 : 255 - 0xff
      12'h2AA: dout  = 8'b11111111; //  682 : 255 - 0xff
      12'h2AB: dout  = 8'b11111111; //  683 : 255 - 0xff
      12'h2AC: dout  = 8'b11111111; //  684 : 255 - 0xff
      12'h2AD: dout  = 8'b11111111; //  685 : 255 - 0xff
      12'h2AE: dout  = 8'b11111111; //  686 : 255 - 0xff
      12'h2AF: dout  = 8'b11111111; //  687 : 255 - 0xff
      12'h2B0: dout  = 8'b00000010; //  688 :   2 - 0x2 -- Sprite 0x56
      12'h2B1: dout  = 8'b00000101; //  689 :   5 - 0x5
      12'h2B2: dout  = 8'b10101010; //  690 : 170 - 0xaa
      12'h2B3: dout  = 8'b01010001; //  691 :  81 - 0x51
      12'h2B4: dout  = 8'b10101010; //  692 : 170 - 0xaa
      12'h2B5: dout  = 8'b01010001; //  693 :  81 - 0x51
      12'h2B6: dout  = 8'b10100010; //  694 : 162 - 0xa2
      12'h2B7: dout  = 8'b00000100; //  695 :   4 - 0x4
      12'h2B8: dout  = 8'b00001000; //  696 :   8 - 0x8 -- Sprite 0x57
      12'h2B9: dout  = 8'b01010101; //  697 :  85 - 0x55
      12'h2BA: dout  = 8'b00101010; //  698 :  42 - 0x2a
      12'h2BB: dout  = 8'b01010101; //  699 :  85 - 0x55
      12'h2BC: dout  = 8'b00101010; //  700 :  42 - 0x2a
      12'h2BD: dout  = 8'b01000101; //  701 :  69 - 0x45
      12'h2BE: dout  = 8'b00001010; //  702 :  10 - 0xa
      12'h2BF: dout  = 8'b00010000; //  703 :  16 - 0x10
      12'h2C0: dout  = 8'b00000000; //  704 :   0 - 0x0 -- Sprite 0x58
      12'h2C1: dout  = 8'b00111111; //  705 :  63 - 0x3f
      12'h2C2: dout  = 8'b01011111; //  706 :  95 - 0x5f
      12'h2C3: dout  = 8'b01101111; //  707 : 111 - 0x6f
      12'h2C4: dout  = 8'b01110000; //  708 : 112 - 0x70
      12'h2C5: dout  = 8'b01110111; //  709 : 119 - 0x77
      12'h2C6: dout  = 8'b01110111; //  710 : 119 - 0x77
      12'h2C7: dout  = 8'b01110111; //  711 : 119 - 0x77
      12'h2C8: dout  = 8'b01110111; //  712 : 119 - 0x77 -- Sprite 0x59
      12'h2C9: dout  = 8'b01110111; //  713 : 119 - 0x77
      12'h2CA: dout  = 8'b01110111; //  714 : 119 - 0x77
      12'h2CB: dout  = 8'b01110000; //  715 : 112 - 0x70
      12'h2CC: dout  = 8'b01101111; //  716 : 111 - 0x6f
      12'h2CD: dout  = 8'b01011111; //  717 :  95 - 0x5f
      12'h2CE: dout  = 8'b00010101; //  718 :  21 - 0x15
      12'h2CF: dout  = 8'b00000000; //  719 :   0 - 0x0
      12'h2D0: dout  = 8'b00000000; //  720 :   0 - 0x0 -- Sprite 0x5a
      12'h2D1: dout  = 8'b11111100; //  721 : 252 - 0xfc
      12'h2D2: dout  = 8'b11111000; //  722 : 248 - 0xf8
      12'h2D3: dout  = 8'b11110110; //  723 : 246 - 0xf6
      12'h2D4: dout  = 8'b00001100; //  724 :  12 - 0xc
      12'h2D5: dout  = 8'b11101110; //  725 : 238 - 0xee
      12'h2D6: dout  = 8'b11101100; //  726 : 236 - 0xec
      12'h2D7: dout  = 8'b11101110; //  727 : 238 - 0xee
      12'h2D8: dout  = 8'b11101100; //  728 : 236 - 0xec -- Sprite 0x5b
      12'h2D9: dout  = 8'b11101110; //  729 : 238 - 0xee
      12'h2DA: dout  = 8'b11101100; //  730 : 236 - 0xec
      12'h2DB: dout  = 8'b00001110; //  731 :  14 - 0xe
      12'h2DC: dout  = 8'b11110100; //  732 : 244 - 0xf4
      12'h2DD: dout  = 8'b11111010; //  733 : 250 - 0xfa
      12'h2DE: dout  = 8'b01010100; //  734 :  84 - 0x54
      12'h2DF: dout  = 8'b00000000; //  735 :   0 - 0x0
      12'h2E0: dout  = 8'b00000000; //  736 :   0 - 0x0 -- Sprite 0x5c
      12'h2E1: dout  = 8'b00011100; //  737 :  28 - 0x1c
      12'h2E2: dout  = 8'b00111110; //  738 :  62 - 0x3e
      12'h2E3: dout  = 8'b00111110; //  739 :  62 - 0x3e
      12'h2E4: dout  = 8'b00111110; //  740 :  62 - 0x3e
      12'h2E5: dout  = 8'b00011100; //  741 :  28 - 0x1c
      12'h2E6: dout  = 8'b00011100; //  742 :  28 - 0x1c
      12'h2E7: dout  = 8'b00000000; //  743 :   0 - 0x0
      12'h2E8: dout  = 8'b00000000; //  744 :   0 - 0x0 -- Sprite 0x5d
      12'h2E9: dout  = 8'b00000000; //  745 :   0 - 0x0
      12'h2EA: dout  = 8'b00000000; //  746 :   0 - 0x0
      12'h2EB: dout  = 8'b00000000; //  747 :   0 - 0x0
      12'h2EC: dout  = 8'b00000000; //  748 :   0 - 0x0
      12'h2ED: dout  = 8'b00000000; //  749 :   0 - 0x0
      12'h2EE: dout  = 8'b00000000; //  750 :   0 - 0x0
      12'h2EF: dout  = 8'b00000000; //  751 :   0 - 0x0
      12'h2F0: dout  = 8'b00000000; //  752 :   0 - 0x0 -- Sprite 0x5e
      12'h2F1: dout  = 8'b00010100; //  753 :  20 - 0x14
      12'h2F2: dout  = 8'b00110110; //  754 :  54 - 0x36
      12'h2F3: dout  = 8'b00111110; //  755 :  62 - 0x3e
      12'h2F4: dout  = 8'b00111110; //  756 :  62 - 0x3e
      12'h2F5: dout  = 8'b00011100; //  757 :  28 - 0x1c
      12'h2F6: dout  = 8'b00001000; //  758 :   8 - 0x8
      12'h2F7: dout  = 8'b00000000; //  759 :   0 - 0x0
      12'h2F8: dout  = 8'b00000000; //  760 :   0 - 0x0 -- Sprite 0x5f
      12'h2F9: dout  = 8'b00010100; //  761 :  20 - 0x14
      12'h2FA: dout  = 8'b00011100; //  762 :  28 - 0x1c
      12'h2FB: dout  = 8'b00011100; //  763 :  28 - 0x1c
      12'h2FC: dout  = 8'b00011100; //  764 :  28 - 0x1c
      12'h2FD: dout  = 8'b00011100; //  765 :  28 - 0x1c
      12'h2FE: dout  = 8'b00011100; //  766 :  28 - 0x1c
      12'h2FF: dout  = 8'b00000000; //  767 :   0 - 0x0
      12'h300: dout  = 8'b00000000; //  768 :   0 - 0x0 -- Sprite 0x60
      12'h301: dout  = 8'b01111111; //  769 : 127 - 0x7f
      12'h302: dout  = 8'b01111111; //  770 : 127 - 0x7f
      12'h303: dout  = 8'b01111111; //  771 : 127 - 0x7f
      12'h304: dout  = 8'b01111111; //  772 : 127 - 0x7f
      12'h305: dout  = 8'b01111111; //  773 : 127 - 0x7f
      12'h306: dout  = 8'b00101010; //  774 :  42 - 0x2a
      12'h307: dout  = 8'b00000000; //  775 :   0 - 0x0
      12'h308: dout  = 8'b00000000; //  776 :   0 - 0x0 -- Sprite 0x61
      12'h309: dout  = 8'b11111111; //  777 : 255 - 0xff
      12'h30A: dout  = 8'b11111111; //  778 : 255 - 0xff
      12'h30B: dout  = 8'b11111111; //  779 : 255 - 0xff
      12'h30C: dout  = 8'b11111111; //  780 : 255 - 0xff
      12'h30D: dout  = 8'b11111111; //  781 : 255 - 0xff
      12'h30E: dout  = 8'b10101010; //  782 : 170 - 0xaa
      12'h30F: dout  = 8'b00000000; //  783 :   0 - 0x0
      12'h310: dout  = 8'b00000000; //  784 :   0 - 0x0 -- Sprite 0x62
      12'h311: dout  = 8'b11111110; //  785 : 254 - 0xfe
      12'h312: dout  = 8'b11111110; //  786 : 254 - 0xfe
      12'h313: dout  = 8'b11111110; //  787 : 254 - 0xfe
      12'h314: dout  = 8'b11111110; //  788 : 254 - 0xfe
      12'h315: dout  = 8'b11111110; //  789 : 254 - 0xfe
      12'h316: dout  = 8'b10101010; //  790 : 170 - 0xaa
      12'h317: dout  = 8'b00000000; //  791 :   0 - 0x0
      12'h318: dout  = 8'b00000000; //  792 :   0 - 0x0 -- Sprite 0x63
      12'h319: dout  = 8'b00000000; //  793 :   0 - 0x0
      12'h31A: dout  = 8'b00000000; //  794 :   0 - 0x0
      12'h31B: dout  = 8'b00000000; //  795 :   0 - 0x0
      12'h31C: dout  = 8'b00000000; //  796 :   0 - 0x0
      12'h31D: dout  = 8'b00000000; //  797 :   0 - 0x0
      12'h31E: dout  = 8'b00000000; //  798 :   0 - 0x0
      12'h31F: dout  = 8'b00000000; //  799 :   0 - 0x0
      12'h320: dout  = 8'b00000000; //  800 :   0 - 0x0 -- Sprite 0x64
      12'h321: dout  = 8'b00000000; //  801 :   0 - 0x0
      12'h322: dout  = 8'b00000001; //  802 :   1 - 0x1
      12'h323: dout  = 8'b00000001; //  803 :   1 - 0x1
      12'h324: dout  = 8'b00000011; //  804 :   3 - 0x3
      12'h325: dout  = 8'b00000011; //  805 :   3 - 0x3
      12'h326: dout  = 8'b00000111; //  806 :   7 - 0x7
      12'h327: dout  = 8'b00000111; //  807 :   7 - 0x7
      12'h328: dout  = 8'b00001111; //  808 :  15 - 0xf -- Sprite 0x65
      12'h329: dout  = 8'b00001111; //  809 :  15 - 0xf
      12'h32A: dout  = 8'b00011111; //  810 :  31 - 0x1f
      12'h32B: dout  = 8'b00011111; //  811 :  31 - 0x1f
      12'h32C: dout  = 8'b00111111; //  812 :  63 - 0x3f
      12'h32D: dout  = 8'b00111111; //  813 :  63 - 0x3f
      12'h32E: dout  = 8'b01010101; //  814 :  85 - 0x55
      12'h32F: dout  = 8'b00000000; //  815 :   0 - 0x0
      12'h330: dout  = 8'b00000000; //  816 :   0 - 0x0 -- Sprite 0x66
      12'h331: dout  = 8'b00000000; //  817 :   0 - 0x0
      12'h332: dout  = 8'b00000000; //  818 :   0 - 0x0
      12'h333: dout  = 8'b10000000; //  819 : 128 - 0x80
      12'h334: dout  = 8'b01000000; //  820 :  64 - 0x40
      12'h335: dout  = 8'b10000000; //  821 : 128 - 0x80
      12'h336: dout  = 8'b11000000; //  822 : 192 - 0xc0
      12'h337: dout  = 8'b11100000; //  823 : 224 - 0xe0
      12'h338: dout  = 8'b11010000; //  824 : 208 - 0xd0 -- Sprite 0x67
      12'h339: dout  = 8'b11100000; //  825 : 224 - 0xe0
      12'h33A: dout  = 8'b11110000; //  826 : 240 - 0xf0
      12'h33B: dout  = 8'b11101000; //  827 : 232 - 0xe8
      12'h33C: dout  = 8'b11110100; //  828 : 244 - 0xf4
      12'h33D: dout  = 8'b11111000; //  829 : 248 - 0xf8
      12'h33E: dout  = 8'b01010100; //  830 :  84 - 0x54
      12'h33F: dout  = 8'b00000000; //  831 :   0 - 0x0
      12'h340: dout  = 8'b00000000; //  832 :   0 - 0x0 -- Sprite 0x68
      12'h341: dout  = 8'b00000000; //  833 :   0 - 0x0
      12'h342: dout  = 8'b00000000; //  834 :   0 - 0x0
      12'h343: dout  = 8'b00000000; //  835 :   0 - 0x0
      12'h344: dout  = 8'b00000000; //  836 :   0 - 0x0
      12'h345: dout  = 8'b00000000; //  837 :   0 - 0x0
      12'h346: dout  = 8'b00000000; //  838 :   0 - 0x0
      12'h347: dout  = 8'b00000000; //  839 :   0 - 0x0
      12'h348: dout  = 8'b00000000; //  840 :   0 - 0x0 -- Sprite 0x69
      12'h349: dout  = 8'b00000000; //  841 :   0 - 0x0
      12'h34A: dout  = 8'b00000000; //  842 :   0 - 0x0
      12'h34B: dout  = 8'b00000000; //  843 :   0 - 0x0
      12'h34C: dout  = 8'b00000000; //  844 :   0 - 0x0
      12'h34D: dout  = 8'b00000000; //  845 :   0 - 0x0
      12'h34E: dout  = 8'b00000000; //  846 :   0 - 0x0
      12'h34F: dout  = 8'b00000000; //  847 :   0 - 0x0
      12'h350: dout  = 8'b00000000; //  848 :   0 - 0x0 -- Sprite 0x6a
      12'h351: dout  = 8'b00000000; //  849 :   0 - 0x0
      12'h352: dout  = 8'b00000000; //  850 :   0 - 0x0
      12'h353: dout  = 8'b00000000; //  851 :   0 - 0x0
      12'h354: dout  = 8'b00000000; //  852 :   0 - 0x0
      12'h355: dout  = 8'b00000000; //  853 :   0 - 0x0
      12'h356: dout  = 8'b00000000; //  854 :   0 - 0x0
      12'h357: dout  = 8'b00000000; //  855 :   0 - 0x0
      12'h358: dout  = 8'b00000000; //  856 :   0 - 0x0 -- Sprite 0x6b
      12'h359: dout  = 8'b00000000; //  857 :   0 - 0x0
      12'h35A: dout  = 8'b00000000; //  858 :   0 - 0x0
      12'h35B: dout  = 8'b00000000; //  859 :   0 - 0x0
      12'h35C: dout  = 8'b00000000; //  860 :   0 - 0x0
      12'h35D: dout  = 8'b00000000; //  861 :   0 - 0x0
      12'h35E: dout  = 8'b00000000; //  862 :   0 - 0x0
      12'h35F: dout  = 8'b00000000; //  863 :   0 - 0x0
      12'h360: dout  = 8'b00000000; //  864 :   0 - 0x0 -- Sprite 0x6c
      12'h361: dout  = 8'b00000000; //  865 :   0 - 0x0
      12'h362: dout  = 8'b00000000; //  866 :   0 - 0x0
      12'h363: dout  = 8'b00000000; //  867 :   0 - 0x0
      12'h364: dout  = 8'b00000000; //  868 :   0 - 0x0
      12'h365: dout  = 8'b00000000; //  869 :   0 - 0x0
      12'h366: dout  = 8'b00000000; //  870 :   0 - 0x0
      12'h367: dout  = 8'b00000000; //  871 :   0 - 0x0
      12'h368: dout  = 8'b00000000; //  872 :   0 - 0x0 -- Sprite 0x6d
      12'h369: dout  = 8'b00000000; //  873 :   0 - 0x0
      12'h36A: dout  = 8'b00000000; //  874 :   0 - 0x0
      12'h36B: dout  = 8'b00000000; //  875 :   0 - 0x0
      12'h36C: dout  = 8'b00000000; //  876 :   0 - 0x0
      12'h36D: dout  = 8'b00000000; //  877 :   0 - 0x0
      12'h36E: dout  = 8'b00000000; //  878 :   0 - 0x0
      12'h36F: dout  = 8'b00000000; //  879 :   0 - 0x0
      12'h370: dout  = 8'b00000000; //  880 :   0 - 0x0 -- Sprite 0x6e
      12'h371: dout  = 8'b00000000; //  881 :   0 - 0x0
      12'h372: dout  = 8'b00000000; //  882 :   0 - 0x0
      12'h373: dout  = 8'b00000000; //  883 :   0 - 0x0
      12'h374: dout  = 8'b00000000; //  884 :   0 - 0x0
      12'h375: dout  = 8'b00000000; //  885 :   0 - 0x0
      12'h376: dout  = 8'b00000000; //  886 :   0 - 0x0
      12'h377: dout  = 8'b00000000; //  887 :   0 - 0x0
      12'h378: dout  = 8'b00000000; //  888 :   0 - 0x0 -- Sprite 0x6f
      12'h379: dout  = 8'b00000000; //  889 :   0 - 0x0
      12'h37A: dout  = 8'b00000000; //  890 :   0 - 0x0
      12'h37B: dout  = 8'b00000000; //  891 :   0 - 0x0
      12'h37C: dout  = 8'b00000000; //  892 :   0 - 0x0
      12'h37D: dout  = 8'b00000000; //  893 :   0 - 0x0
      12'h37E: dout  = 8'b00000000; //  894 :   0 - 0x0
      12'h37F: dout  = 8'b00000000; //  895 :   0 - 0x0
      12'h380: dout  = 8'b00000000; //  896 :   0 - 0x0 -- Sprite 0x70
      12'h381: dout  = 8'b00000000; //  897 :   0 - 0x0
      12'h382: dout  = 8'b00000000; //  898 :   0 - 0x0
      12'h383: dout  = 8'b00000000; //  899 :   0 - 0x0
      12'h384: dout  = 8'b00000000; //  900 :   0 - 0x0
      12'h385: dout  = 8'b00000000; //  901 :   0 - 0x0
      12'h386: dout  = 8'b00000000; //  902 :   0 - 0x0
      12'h387: dout  = 8'b00000000; //  903 :   0 - 0x0
      12'h388: dout  = 8'b00000000; //  904 :   0 - 0x0 -- Sprite 0x71
      12'h389: dout  = 8'b00000000; //  905 :   0 - 0x0
      12'h38A: dout  = 8'b00000000; //  906 :   0 - 0x0
      12'h38B: dout  = 8'b00000000; //  907 :   0 - 0x0
      12'h38C: dout  = 8'b00000000; //  908 :   0 - 0x0
      12'h38D: dout  = 8'b00000000; //  909 :   0 - 0x0
      12'h38E: dout  = 8'b00000000; //  910 :   0 - 0x0
      12'h38F: dout  = 8'b00000000; //  911 :   0 - 0x0
      12'h390: dout  = 8'b00000000; //  912 :   0 - 0x0 -- Sprite 0x72
      12'h391: dout  = 8'b00000000; //  913 :   0 - 0x0
      12'h392: dout  = 8'b00000000; //  914 :   0 - 0x0
      12'h393: dout  = 8'b00000000; //  915 :   0 - 0x0
      12'h394: dout  = 8'b00000000; //  916 :   0 - 0x0
      12'h395: dout  = 8'b00000000; //  917 :   0 - 0x0
      12'h396: dout  = 8'b00000000; //  918 :   0 - 0x0
      12'h397: dout  = 8'b00000000; //  919 :   0 - 0x0
      12'h398: dout  = 8'b00000000; //  920 :   0 - 0x0 -- Sprite 0x73
      12'h399: dout  = 8'b00000000; //  921 :   0 - 0x0
      12'h39A: dout  = 8'b00000000; //  922 :   0 - 0x0
      12'h39B: dout  = 8'b00000000; //  923 :   0 - 0x0
      12'h39C: dout  = 8'b00000000; //  924 :   0 - 0x0
      12'h39D: dout  = 8'b00000000; //  925 :   0 - 0x0
      12'h39E: dout  = 8'b00000000; //  926 :   0 - 0x0
      12'h39F: dout  = 8'b00000000; //  927 :   0 - 0x0
      12'h3A0: dout  = 8'b00000000; //  928 :   0 - 0x0 -- Sprite 0x74
      12'h3A1: dout  = 8'b00000000; //  929 :   0 - 0x0
      12'h3A2: dout  = 8'b00000000; //  930 :   0 - 0x0
      12'h3A3: dout  = 8'b00000000; //  931 :   0 - 0x0
      12'h3A4: dout  = 8'b00000000; //  932 :   0 - 0x0
      12'h3A5: dout  = 8'b00000000; //  933 :   0 - 0x0
      12'h3A6: dout  = 8'b00000000; //  934 :   0 - 0x0
      12'h3A7: dout  = 8'b00000000; //  935 :   0 - 0x0
      12'h3A8: dout  = 8'b00000000; //  936 :   0 - 0x0 -- Sprite 0x75
      12'h3A9: dout  = 8'b00000000; //  937 :   0 - 0x0
      12'h3AA: dout  = 8'b00000000; //  938 :   0 - 0x0
      12'h3AB: dout  = 8'b00000000; //  939 :   0 - 0x0
      12'h3AC: dout  = 8'b00000000; //  940 :   0 - 0x0
      12'h3AD: dout  = 8'b00000000; //  941 :   0 - 0x0
      12'h3AE: dout  = 8'b00000000; //  942 :   0 - 0x0
      12'h3AF: dout  = 8'b00000000; //  943 :   0 - 0x0
      12'h3B0: dout  = 8'b00000000; //  944 :   0 - 0x0 -- Sprite 0x76
      12'h3B1: dout  = 8'b00000000; //  945 :   0 - 0x0
      12'h3B2: dout  = 8'b00000000; //  946 :   0 - 0x0
      12'h3B3: dout  = 8'b00000000; //  947 :   0 - 0x0
      12'h3B4: dout  = 8'b00000000; //  948 :   0 - 0x0
      12'h3B5: dout  = 8'b00000000; //  949 :   0 - 0x0
      12'h3B6: dout  = 8'b00000000; //  950 :   0 - 0x0
      12'h3B7: dout  = 8'b00000000; //  951 :   0 - 0x0
      12'h3B8: dout  = 8'b00000000; //  952 :   0 - 0x0 -- Sprite 0x77
      12'h3B9: dout  = 8'b00000000; //  953 :   0 - 0x0
      12'h3BA: dout  = 8'b00000000; //  954 :   0 - 0x0
      12'h3BB: dout  = 8'b00000000; //  955 :   0 - 0x0
      12'h3BC: dout  = 8'b00000000; //  956 :   0 - 0x0
      12'h3BD: dout  = 8'b00000000; //  957 :   0 - 0x0
      12'h3BE: dout  = 8'b00000000; //  958 :   0 - 0x0
      12'h3BF: dout  = 8'b00000000; //  959 :   0 - 0x0
      12'h3C0: dout  = 8'b00000000; //  960 :   0 - 0x0 -- Sprite 0x78
      12'h3C1: dout  = 8'b00000000; //  961 :   0 - 0x0
      12'h3C2: dout  = 8'b00000000; //  962 :   0 - 0x0
      12'h3C3: dout  = 8'b00000000; //  963 :   0 - 0x0
      12'h3C4: dout  = 8'b00000000; //  964 :   0 - 0x0
      12'h3C5: dout  = 8'b00000000; //  965 :   0 - 0x0
      12'h3C6: dout  = 8'b00000000; //  966 :   0 - 0x0
      12'h3C7: dout  = 8'b00000000; //  967 :   0 - 0x0
      12'h3C8: dout  = 8'b00000000; //  968 :   0 - 0x0 -- Sprite 0x79
      12'h3C9: dout  = 8'b00000000; //  969 :   0 - 0x0
      12'h3CA: dout  = 8'b00000000; //  970 :   0 - 0x0
      12'h3CB: dout  = 8'b00000000; //  971 :   0 - 0x0
      12'h3CC: dout  = 8'b00000000; //  972 :   0 - 0x0
      12'h3CD: dout  = 8'b00000000; //  973 :   0 - 0x0
      12'h3CE: dout  = 8'b00000000; //  974 :   0 - 0x0
      12'h3CF: dout  = 8'b00000000; //  975 :   0 - 0x0
      12'h3D0: dout  = 8'b00000000; //  976 :   0 - 0x0 -- Sprite 0x7a
      12'h3D1: dout  = 8'b00000000; //  977 :   0 - 0x0
      12'h3D2: dout  = 8'b00000000; //  978 :   0 - 0x0
      12'h3D3: dout  = 8'b00000000; //  979 :   0 - 0x0
      12'h3D4: dout  = 8'b00000000; //  980 :   0 - 0x0
      12'h3D5: dout  = 8'b00000000; //  981 :   0 - 0x0
      12'h3D6: dout  = 8'b00000000; //  982 :   0 - 0x0
      12'h3D7: dout  = 8'b00000000; //  983 :   0 - 0x0
      12'h3D8: dout  = 8'b00000000; //  984 :   0 - 0x0 -- Sprite 0x7b
      12'h3D9: dout  = 8'b00000000; //  985 :   0 - 0x0
      12'h3DA: dout  = 8'b00000000; //  986 :   0 - 0x0
      12'h3DB: dout  = 8'b00000000; //  987 :   0 - 0x0
      12'h3DC: dout  = 8'b00000000; //  988 :   0 - 0x0
      12'h3DD: dout  = 8'b00000000; //  989 :   0 - 0x0
      12'h3DE: dout  = 8'b00000000; //  990 :   0 - 0x0
      12'h3DF: dout  = 8'b00000000; //  991 :   0 - 0x0
      12'h3E0: dout  = 8'b00000000; //  992 :   0 - 0x0 -- Sprite 0x7c
      12'h3E1: dout  = 8'b00000000; //  993 :   0 - 0x0
      12'h3E2: dout  = 8'b00000000; //  994 :   0 - 0x0
      12'h3E3: dout  = 8'b00000000; //  995 :   0 - 0x0
      12'h3E4: dout  = 8'b00000000; //  996 :   0 - 0x0
      12'h3E5: dout  = 8'b00000000; //  997 :   0 - 0x0
      12'h3E6: dout  = 8'b00000000; //  998 :   0 - 0x0
      12'h3E7: dout  = 8'b00000000; //  999 :   0 - 0x0
      12'h3E8: dout  = 8'b00000000; // 1000 :   0 - 0x0 -- Sprite 0x7d
      12'h3E9: dout  = 8'b00000000; // 1001 :   0 - 0x0
      12'h3EA: dout  = 8'b00000000; // 1002 :   0 - 0x0
      12'h3EB: dout  = 8'b00000000; // 1003 :   0 - 0x0
      12'h3EC: dout  = 8'b00000000; // 1004 :   0 - 0x0
      12'h3ED: dout  = 8'b00000000; // 1005 :   0 - 0x0
      12'h3EE: dout  = 8'b00000000; // 1006 :   0 - 0x0
      12'h3EF: dout  = 8'b00000000; // 1007 :   0 - 0x0
      12'h3F0: dout  = 8'b00000000; // 1008 :   0 - 0x0 -- Sprite 0x7e
      12'h3F1: dout  = 8'b00000000; // 1009 :   0 - 0x0
      12'h3F2: dout  = 8'b00000000; // 1010 :   0 - 0x0
      12'h3F3: dout  = 8'b00000000; // 1011 :   0 - 0x0
      12'h3F4: dout  = 8'b00000000; // 1012 :   0 - 0x0
      12'h3F5: dout  = 8'b00000000; // 1013 :   0 - 0x0
      12'h3F6: dout  = 8'b00000000; // 1014 :   0 - 0x0
      12'h3F7: dout  = 8'b00000000; // 1015 :   0 - 0x0
      12'h3F8: dout  = 8'b00000000; // 1016 :   0 - 0x0 -- Sprite 0x7f
      12'h3F9: dout  = 8'b00000000; // 1017 :   0 - 0x0
      12'h3FA: dout  = 8'b00000000; // 1018 :   0 - 0x0
      12'h3FB: dout  = 8'b00000000; // 1019 :   0 - 0x0
      12'h3FC: dout  = 8'b00000000; // 1020 :   0 - 0x0
      12'h3FD: dout  = 8'b00000000; // 1021 :   0 - 0x0
      12'h3FE: dout  = 8'b00000000; // 1022 :   0 - 0x0
      12'h3FF: dout  = 8'b00000000; // 1023 :   0 - 0x0
      12'h400: dout  = 8'b00000000; // 1024 :   0 - 0x0 -- Sprite 0x80
      12'h401: dout  = 8'b00000011; // 1025 :   3 - 0x3
      12'h402: dout  = 8'b00001111; // 1026 :  15 - 0xf
      12'h403: dout  = 8'b00011111; // 1027 :  31 - 0x1f
      12'h404: dout  = 8'b00011111; // 1028 :  31 - 0x1f
      12'h405: dout  = 8'b00111111; // 1029 :  63 - 0x3f
      12'h406: dout  = 8'b00111111; // 1030 :  63 - 0x3f
      12'h407: dout  = 8'b00000000; // 1031 :   0 - 0x0
      12'h408: dout  = 8'b00000000; // 1032 :   0 - 0x0 -- Sprite 0x81
      12'h409: dout  = 8'b00000000; // 1033 :   0 - 0x0
      12'h40A: dout  = 8'b00000000; // 1034 :   0 - 0x0
      12'h40B: dout  = 8'b00000000; // 1035 :   0 - 0x0
      12'h40C: dout  = 8'b00000000; // 1036 :   0 - 0x0
      12'h40D: dout  = 8'b00000000; // 1037 :   0 - 0x0
      12'h40E: dout  = 8'b00000000; // 1038 :   0 - 0x0
      12'h40F: dout  = 8'b00000000; // 1039 :   0 - 0x0
      12'h410: dout  = 8'b00000000; // 1040 :   0 - 0x0 -- Sprite 0x82
      12'h411: dout  = 8'b11000000; // 1041 : 192 - 0xc0
      12'h412: dout  = 8'b11110000; // 1042 : 240 - 0xf0
      12'h413: dout  = 8'b11110000; // 1043 : 240 - 0xf0
      12'h414: dout  = 8'b11101100; // 1044 : 236 - 0xec
      12'h415: dout  = 8'b11100000; // 1045 : 224 - 0xe0
      12'h416: dout  = 8'b11111100; // 1046 : 252 - 0xfc
      12'h417: dout  = 8'b00000000; // 1047 :   0 - 0x0
      12'h418: dout  = 8'b00000000; // 1048 :   0 - 0x0 -- Sprite 0x83
      12'h419: dout  = 8'b00000000; // 1049 :   0 - 0x0
      12'h41A: dout  = 8'b00000000; // 1050 :   0 - 0x0
      12'h41B: dout  = 8'b00000000; // 1051 :   0 - 0x0
      12'h41C: dout  = 8'b00000000; // 1052 :   0 - 0x0
      12'h41D: dout  = 8'b00000000; // 1053 :   0 - 0x0
      12'h41E: dout  = 8'b11100000; // 1054 : 224 - 0xe0
      12'h41F: dout  = 8'b00000000; // 1055 :   0 - 0x0
      12'h420: dout  = 8'b00000000; // 1056 :   0 - 0x0 -- Sprite 0x84
      12'h421: dout  = 8'b00000011; // 1057 :   3 - 0x3
      12'h422: dout  = 8'b00001111; // 1058 :  15 - 0xf
      12'h423: dout  = 8'b00011111; // 1059 :  31 - 0x1f
      12'h424: dout  = 8'b00011111; // 1060 :  31 - 0x1f
      12'h425: dout  = 8'b00111111; // 1061 :  63 - 0x3f
      12'h426: dout  = 8'b00111111; // 1062 :  63 - 0x3f
      12'h427: dout  = 8'b00000000; // 1063 :   0 - 0x0
      12'h428: dout  = 8'b00000000; // 1064 :   0 - 0x0 -- Sprite 0x85
      12'h429: dout  = 8'b00000000; // 1065 :   0 - 0x0
      12'h42A: dout  = 8'b00000000; // 1066 :   0 - 0x0
      12'h42B: dout  = 8'b00000000; // 1067 :   0 - 0x0
      12'h42C: dout  = 8'b00000000; // 1068 :   0 - 0x0
      12'h42D: dout  = 8'b00001000; // 1069 :   8 - 0x8
      12'h42E: dout  = 8'b00001110; // 1070 :  14 - 0xe
      12'h42F: dout  = 8'b00000000; // 1071 :   0 - 0x0
      12'h430: dout  = 8'b00000000; // 1072 :   0 - 0x0 -- Sprite 0x86
      12'h431: dout  = 8'b11000000; // 1073 : 192 - 0xc0
      12'h432: dout  = 8'b11110000; // 1074 : 240 - 0xf0
      12'h433: dout  = 8'b11110000; // 1075 : 240 - 0xf0
      12'h434: dout  = 8'b11101100; // 1076 : 236 - 0xec
      12'h435: dout  = 8'b11100000; // 1077 : 224 - 0xe0
      12'h436: dout  = 8'b11111100; // 1078 : 252 - 0xfc
      12'h437: dout  = 8'b00000000; // 1079 :   0 - 0x0
      12'h438: dout  = 8'b00000000; // 1080 :   0 - 0x0 -- Sprite 0x87
      12'h439: dout  = 8'b00000000; // 1081 :   0 - 0x0
      12'h43A: dout  = 8'b00000000; // 1082 :   0 - 0x0
      12'h43B: dout  = 8'b00000000; // 1083 :   0 - 0x0
      12'h43C: dout  = 8'b00000000; // 1084 :   0 - 0x0
      12'h43D: dout  = 8'b00000110; // 1085 :   6 - 0x6
      12'h43E: dout  = 8'b00001100; // 1086 :  12 - 0xc
      12'h43F: dout  = 8'b00000000; // 1087 :   0 - 0x0
      12'h440: dout  = 8'b00000000; // 1088 :   0 - 0x0 -- Sprite 0x88
      12'h441: dout  = 8'b00000011; // 1089 :   3 - 0x3
      12'h442: dout  = 8'b00000011; // 1090 :   3 - 0x3
      12'h443: dout  = 8'b00000100; // 1091 :   4 - 0x4
      12'h444: dout  = 8'b00001111; // 1092 :  15 - 0xf
      12'h445: dout  = 8'b00011111; // 1093 :  31 - 0x1f
      12'h446: dout  = 8'b01101111; // 1094 : 111 - 0x6f
      12'h447: dout  = 8'b01101111; // 1095 : 111 - 0x6f
      12'h448: dout  = 8'b01101111; // 1096 : 111 - 0x6f -- Sprite 0x89
      12'h449: dout  = 8'b01101111; // 1097 : 111 - 0x6f
      12'h44A: dout  = 8'b00011111; // 1098 :  31 - 0x1f
      12'h44B: dout  = 8'b00001111; // 1099 :  15 - 0xf
      12'h44C: dout  = 8'b00000100; // 1100 :   4 - 0x4
      12'h44D: dout  = 8'b00000011; // 1101 :   3 - 0x3
      12'h44E: dout  = 8'b00000011; // 1102 :   3 - 0x3
      12'h44F: dout  = 8'b00000000; // 1103 :   0 - 0x0
      12'h450: dout  = 8'b00000000; // 1104 :   0 - 0x0 -- Sprite 0x8a
      12'h451: dout  = 8'b00000000; // 1105 :   0 - 0x0
      12'h452: dout  = 8'b00011000; // 1106 :  24 - 0x18
      12'h453: dout  = 8'b00110111; // 1107 :  55 - 0x37
      12'h454: dout  = 8'b00101111; // 1108 :  47 - 0x2f
      12'h455: dout  = 8'b00011111; // 1109 :  31 - 0x1f
      12'h456: dout  = 8'b00011111; // 1110 :  31 - 0x1f
      12'h457: dout  = 8'b00011111; // 1111 :  31 - 0x1f
      12'h458: dout  = 8'b00011111; // 1112 :  31 - 0x1f -- Sprite 0x8b
      12'h459: dout  = 8'b00011111; // 1113 :  31 - 0x1f
      12'h45A: dout  = 8'b00011111; // 1114 :  31 - 0x1f
      12'h45B: dout  = 8'b00101111; // 1115 :  47 - 0x2f
      12'h45C: dout  = 8'b00110111; // 1116 :  55 - 0x37
      12'h45D: dout  = 8'b00011000; // 1117 :  24 - 0x18
      12'h45E: dout  = 8'b00000000; // 1118 :   0 - 0x0
      12'h45F: dout  = 8'b00000000; // 1119 :   0 - 0x0
      12'h460: dout  = 8'b00000000; // 1120 :   0 - 0x0 -- Sprite 0x8c
      12'h461: dout  = 8'b00000011; // 1121 :   3 - 0x3
      12'h462: dout  = 8'b00000001; // 1122 :   1 - 0x1
      12'h463: dout  = 8'b00011001; // 1123 :  25 - 0x19
      12'h464: dout  = 8'b00111001; // 1124 :  57 - 0x39
      12'h465: dout  = 8'b00011011; // 1125 :  27 - 0x1b
      12'h466: dout  = 8'b00001111; // 1126 :  15 - 0xf
      12'h467: dout  = 8'b00001111; // 1127 :  15 - 0xf
      12'h468: dout  = 8'b01111111; // 1128 : 127 - 0x7f -- Sprite 0x8d
      12'h469: dout  = 8'b01111111; // 1129 : 127 - 0x7f
      12'h46A: dout  = 8'b00111111; // 1130 :  63 - 0x3f
      12'h46B: dout  = 8'b00010111; // 1131 :  23 - 0x17
      12'h46C: dout  = 8'b00000110; // 1132 :   6 - 0x6
      12'h46D: dout  = 8'b00000100; // 1133 :   4 - 0x4
      12'h46E: dout  = 8'b00000111; // 1134 :   7 - 0x7
      12'h46F: dout  = 8'b00000000; // 1135 :   0 - 0x0
      12'h470: dout  = 8'b00000000; // 1136 :   0 - 0x0 -- Sprite 0x8e
      12'h471: dout  = 8'b11000000; // 1137 : 192 - 0xc0
      12'h472: dout  = 8'b11110000; // 1138 : 240 - 0xf0
      12'h473: dout  = 8'b10111000; // 1139 : 184 - 0xb8
      12'h474: dout  = 8'b10011100; // 1140 : 156 - 0x9c
      12'h475: dout  = 8'b11111100; // 1141 : 252 - 0xfc
      12'h476: dout  = 8'b11111110; // 1142 : 254 - 0xfe
      12'h477: dout  = 8'b11000000; // 1143 : 192 - 0xc0
      12'h478: dout  = 8'b11111110; // 1144 : 254 - 0xfe -- Sprite 0x8f
      12'h479: dout  = 8'b11111110; // 1145 : 254 - 0xfe
      12'h47A: dout  = 8'b11111000; // 1146 : 248 - 0xf8
      12'h47B: dout  = 8'b11110000; // 1147 : 240 - 0xf0
      12'h47C: dout  = 8'b11000000; // 1148 : 192 - 0xc0
      12'h47D: dout  = 8'b00000000; // 1149 :   0 - 0x0
      12'h47E: dout  = 8'b00000000; // 1150 :   0 - 0x0
      12'h47F: dout  = 8'b10000000; // 1151 : 128 - 0x80
      12'h480: dout  = 8'b00000000; // 1152 :   0 - 0x0 -- Sprite 0x90
      12'h481: dout  = 8'b00000001; // 1153 :   1 - 0x1
      12'h482: dout  = 8'b00001001; // 1154 :   9 - 0x9
      12'h483: dout  = 8'b00011001; // 1155 :  25 - 0x19
      12'h484: dout  = 8'b00011100; // 1156 :  28 - 0x1c
      12'h485: dout  = 8'b00001101; // 1157 :  13 - 0xd
      12'h486: dout  = 8'b00001111; // 1158 :  15 - 0xf
      12'h487: dout  = 8'b00101111; // 1159 :  47 - 0x2f
      12'h488: dout  = 8'b01111111; // 1160 : 127 - 0x7f -- Sprite 0x91
      12'h489: dout  = 8'b01111111; // 1161 : 127 - 0x7f
      12'h48A: dout  = 8'b00111111; // 1162 :  63 - 0x3f
      12'h48B: dout  = 8'b00011011; // 1163 :  27 - 0x1b
      12'h48C: dout  = 8'b00000011; // 1164 :   3 - 0x3
      12'h48D: dout  = 8'b00000011; // 1165 :   3 - 0x3
      12'h48E: dout  = 8'b00000001; // 1166 :   1 - 0x1
      12'h48F: dout  = 8'b00000000; // 1167 :   0 - 0x0
      12'h490: dout  = 8'b00000000; // 1168 :   0 - 0x0 -- Sprite 0x92
      12'h491: dout  = 8'b11000000; // 1169 : 192 - 0xc0
      12'h492: dout  = 8'b11110000; // 1170 : 240 - 0xf0
      12'h493: dout  = 8'b11011000; // 1171 : 216 - 0xd8
      12'h494: dout  = 8'b11001100; // 1172 : 204 - 0xcc
      12'h495: dout  = 8'b11111100; // 1173 : 252 - 0xfc
      12'h496: dout  = 8'b11111110; // 1174 : 254 - 0xfe
      12'h497: dout  = 8'b11100000; // 1175 : 224 - 0xe0
      12'h498: dout  = 8'b11111110; // 1176 : 254 - 0xfe -- Sprite 0x93
      12'h499: dout  = 8'b11111110; // 1177 : 254 - 0xfe
      12'h49A: dout  = 8'b11111000; // 1178 : 248 - 0xf8
      12'h49B: dout  = 8'b01110000; // 1179 : 112 - 0x70
      12'h49C: dout  = 8'b01000000; // 1180 :  64 - 0x40
      12'h49D: dout  = 8'b00000000; // 1181 :   0 - 0x0
      12'h49E: dout  = 8'b11000000; // 1182 : 192 - 0xc0
      12'h49F: dout  = 8'b00100000; // 1183 :  32 - 0x20
      12'h4A0: dout  = 8'b00000000; // 1184 :   0 - 0x0 -- Sprite 0x94
      12'h4A1: dout  = 8'b00000000; // 1185 :   0 - 0x0
      12'h4A2: dout  = 8'b00001100; // 1186 :  12 - 0xc
      12'h4A3: dout  = 8'b00001110; // 1187 :  14 - 0xe
      12'h4A4: dout  = 8'b00000110; // 1188 :   6 - 0x6
      12'h4A5: dout  = 8'b00100110; // 1189 :  38 - 0x26
      12'h4A6: dout  = 8'b00110111; // 1190 :  55 - 0x37
      12'h4A7: dout  = 8'b00110011; // 1191 :  51 - 0x33
      12'h4A8: dout  = 8'b01111111; // 1192 : 127 - 0x7f -- Sprite 0x95
      12'h4A9: dout  = 8'b01111111; // 1193 : 127 - 0x7f
      12'h4AA: dout  = 8'b00111111; // 1194 :  63 - 0x3f
      12'h4AB: dout  = 8'b00011111; // 1195 :  31 - 0x1f
      12'h4AC: dout  = 8'b00001110; // 1196 :  14 - 0xe
      12'h4AD: dout  = 8'b00000000; // 1197 :   0 - 0x0
      12'h4AE: dout  = 8'b00000000; // 1198 :   0 - 0x0
      12'h4AF: dout  = 8'b00000000; // 1199 :   0 - 0x0
      12'h4B0: dout  = 8'b00000000; // 1200 :   0 - 0x0 -- Sprite 0x96
      12'h4B1: dout  = 8'b11000000; // 1201 : 192 - 0xc0
      12'h4B2: dout  = 8'b11110000; // 1202 : 240 - 0xf0
      12'h4B3: dout  = 8'b01101000; // 1203 : 104 - 0x68
      12'h4B4: dout  = 8'b01100100; // 1204 : 100 - 0x64
      12'h4B5: dout  = 8'b11111100; // 1205 : 252 - 0xfc
      12'h4B6: dout  = 8'b11111110; // 1206 : 254 - 0xfe
      12'h4B7: dout  = 8'b11110000; // 1207 : 240 - 0xf0
      12'h4B8: dout  = 8'b11111111; // 1208 : 255 - 0xff -- Sprite 0x97
      12'h4B9: dout  = 8'b11111110; // 1209 : 254 - 0xfe
      12'h4BA: dout  = 8'b11111100; // 1210 : 252 - 0xfc
      12'h4BB: dout  = 8'b10110000; // 1211 : 176 - 0xb0
      12'h4BC: dout  = 8'b11000000; // 1212 : 192 - 0xc0
      12'h4BD: dout  = 8'b11000000; // 1213 : 192 - 0xc0
      12'h4BE: dout  = 8'b01110000; // 1214 : 112 - 0x70
      12'h4BF: dout  = 8'b00001000; // 1215 :   8 - 0x8
      12'h4C0: dout  = 8'b00000000; // 1216 :   0 - 0x0 -- Sprite 0x98
      12'h4C1: dout  = 8'b00000001; // 1217 :   1 - 0x1
      12'h4C2: dout  = 8'b00000000; // 1218 :   0 - 0x0
      12'h4C3: dout  = 8'b00000000; // 1219 :   0 - 0x0
      12'h4C4: dout  = 8'b00000000; // 1220 :   0 - 0x0
      12'h4C5: dout  = 8'b00000000; // 1221 :   0 - 0x0
      12'h4C6: dout  = 8'b00000001; // 1222 :   1 - 0x1
      12'h4C7: dout  = 8'b00000011; // 1223 :   3 - 0x3
      12'h4C8: dout  = 8'b00000111; // 1224 :   7 - 0x7 -- Sprite 0x99
      12'h4C9: dout  = 8'b00010111; // 1225 :  23 - 0x17
      12'h4CA: dout  = 8'b00101111; // 1226 :  47 - 0x2f
      12'h4CB: dout  = 8'b00011110; // 1227 :  30 - 0x1e
      12'h4CC: dout  = 8'b00010001; // 1228 :  17 - 0x11
      12'h4CD: dout  = 8'b00000000; // 1229 :   0 - 0x0
      12'h4CE: dout  = 8'b00000001; // 1230 :   1 - 0x1
      12'h4CF: dout  = 8'b00000000; // 1231 :   0 - 0x0
      12'h4D0: dout  = 8'b00000000; // 1232 :   0 - 0x0 -- Sprite 0x9a
      12'h4D1: dout  = 8'b00010000; // 1233 :  16 - 0x10
      12'h4D2: dout  = 8'b01111000; // 1234 : 120 - 0x78
      12'h4D3: dout  = 8'b01110100; // 1235 : 116 - 0x74
      12'h4D4: dout  = 8'b11111110; // 1236 : 254 - 0xfe
      12'h4D5: dout  = 8'b11111000; // 1237 : 248 - 0xf8
      12'h4D6: dout  = 8'b11111100; // 1238 : 252 - 0xfc
      12'h4D7: dout  = 8'b11111000; // 1239 : 248 - 0xf8
      12'h4D8: dout  = 8'b11111000; // 1240 : 248 - 0xf8 -- Sprite 0x9b
      12'h4D9: dout  = 8'b11010000; // 1241 : 208 - 0xd0
      12'h4DA: dout  = 8'b00110000; // 1242 :  48 - 0x30
      12'h4DB: dout  = 8'b01100000; // 1243 :  96 - 0x60
      12'h4DC: dout  = 8'b10000000; // 1244 : 128 - 0x80
      12'h4DD: dout  = 8'b00000000; // 1245 :   0 - 0x0
      12'h4DE: dout  = 8'b00000000; // 1246 :   0 - 0x0
      12'h4DF: dout  = 8'b00000000; // 1247 :   0 - 0x0
      12'h4E0: dout  = 8'b00000000; // 1248 :   0 - 0x0 -- Sprite 0x9c
      12'h4E1: dout  = 8'b00000001; // 1249 :   1 - 0x1
      12'h4E2: dout  = 8'b00000000; // 1250 :   0 - 0x0
      12'h4E3: dout  = 8'b00000000; // 1251 :   0 - 0x0
      12'h4E4: dout  = 8'b00000000; // 1252 :   0 - 0x0
      12'h4E5: dout  = 8'b00000000; // 1253 :   0 - 0x0
      12'h4E6: dout  = 8'b00000001; // 1254 :   1 - 0x1
      12'h4E7: dout  = 8'b00000011; // 1255 :   3 - 0x3
      12'h4E8: dout  = 8'b00000111; // 1256 :   7 - 0x7 -- Sprite 0x9d
      12'h4E9: dout  = 8'b00010111; // 1257 :  23 - 0x17
      12'h4EA: dout  = 8'b00101111; // 1258 :  47 - 0x2f
      12'h4EB: dout  = 8'b00011110; // 1259 :  30 - 0x1e
      12'h4EC: dout  = 8'b00010000; // 1260 :  16 - 0x10
      12'h4ED: dout  = 8'b00000100; // 1261 :   4 - 0x4
      12'h4EE: dout  = 8'b00000000; // 1262 :   0 - 0x0
      12'h4EF: dout  = 8'b00000000; // 1263 :   0 - 0x0
      12'h4F0: dout  = 8'b00000000; // 1264 :   0 - 0x0 -- Sprite 0x9e
      12'h4F1: dout  = 8'b00010000; // 1265 :  16 - 0x10
      12'h4F2: dout  = 8'b01111000; // 1266 : 120 - 0x78
      12'h4F3: dout  = 8'b01110100; // 1267 : 116 - 0x74
      12'h4F4: dout  = 8'b11111110; // 1268 : 254 - 0xfe
      12'h4F5: dout  = 8'b11111000; // 1269 : 248 - 0xf8
      12'h4F6: dout  = 8'b11111100; // 1270 : 252 - 0xfc
      12'h4F7: dout  = 8'b11111000; // 1271 : 248 - 0xf8
      12'h4F8: dout  = 8'b11111000; // 1272 : 248 - 0xf8 -- Sprite 0x9f
      12'h4F9: dout  = 8'b11010000; // 1273 : 208 - 0xd0
      12'h4FA: dout  = 8'b00110000; // 1274 :  48 - 0x30
      12'h4FB: dout  = 8'b11000000; // 1275 : 192 - 0xc0
      12'h4FC: dout  = 8'b00000000; // 1276 :   0 - 0x0
      12'h4FD: dout  = 8'b00000000; // 1277 :   0 - 0x0
      12'h4FE: dout  = 8'b00000000; // 1278 :   0 - 0x0
      12'h4FF: dout  = 8'b00000000; // 1279 :   0 - 0x0
      12'h500: dout  = 8'b00000000; // 1280 :   0 - 0x0 -- Sprite 0xa0
      12'h501: dout  = 8'b00000011; // 1281 :   3 - 0x3
      12'h502: dout  = 8'b00001111; // 1282 :  15 - 0xf
      12'h503: dout  = 8'b00011111; // 1283 :  31 - 0x1f
      12'h504: dout  = 8'b00111111; // 1284 :  63 - 0x3f
      12'h505: dout  = 8'b00111111; // 1285 :  63 - 0x3f
      12'h506: dout  = 8'b01111111; // 1286 : 127 - 0x7f
      12'h507: dout  = 8'b01111111; // 1287 : 127 - 0x7f
      12'h508: dout  = 8'b01111111; // 1288 : 127 - 0x7f -- Sprite 0xa1
      12'h509: dout  = 8'b01111111; // 1289 : 127 - 0x7f
      12'h50A: dout  = 8'b00111111; // 1290 :  63 - 0x3f
      12'h50B: dout  = 8'b00111111; // 1291 :  63 - 0x3f
      12'h50C: dout  = 8'b00011111; // 1292 :  31 - 0x1f
      12'h50D: dout  = 8'b00000101; // 1293 :   5 - 0x5
      12'h50E: dout  = 8'b00000010; // 1294 :   2 - 0x2
      12'h50F: dout  = 8'b00000000; // 1295 :   0 - 0x0
      12'h510: dout  = 8'b00000000; // 1296 :   0 - 0x0 -- Sprite 0xa2
      12'h511: dout  = 8'b11000000; // 1297 : 192 - 0xc0
      12'h512: dout  = 8'b11110000; // 1298 : 240 - 0xf0
      12'h513: dout  = 8'b11111000; // 1299 : 248 - 0xf8
      12'h514: dout  = 8'b11111000; // 1300 : 248 - 0xf8
      12'h515: dout  = 8'b11111100; // 1301 : 252 - 0xfc
      12'h516: dout  = 8'b11111010; // 1302 : 250 - 0xfa
      12'h517: dout  = 8'b11111100; // 1303 : 252 - 0xfc
      12'h518: dout  = 8'b11111010; // 1304 : 250 - 0xfa -- Sprite 0xa3
      12'h519: dout  = 8'b11110100; // 1305 : 244 - 0xf4
      12'h51A: dout  = 8'b11101000; // 1306 : 232 - 0xe8
      12'h51B: dout  = 8'b11010100; // 1307 : 212 - 0xd4
      12'h51C: dout  = 8'b10101000; // 1308 : 168 - 0xa8
      12'h51D: dout  = 8'b01010000; // 1309 :  80 - 0x50
      12'h51E: dout  = 8'b10000000; // 1310 : 128 - 0x80
      12'h51F: dout  = 8'b00000000; // 1311 :   0 - 0x0
      12'h520: dout  = 8'b00000000; // 1312 :   0 - 0x0 -- Sprite 0xa4
      12'h521: dout  = 8'b00000000; // 1313 :   0 - 0x0
      12'h522: dout  = 8'b00000000; // 1314 :   0 - 0x0
      12'h523: dout  = 8'b00001110; // 1315 :  14 - 0xe
      12'h524: dout  = 8'b00000000; // 1316 :   0 - 0x0
      12'h525: dout  = 8'b00001010; // 1317 :  10 - 0xa
      12'h526: dout  = 8'b01001010; // 1318 :  74 - 0x4a
      12'h527: dout  = 8'b01100000; // 1319 :  96 - 0x60
      12'h528: dout  = 8'b01111111; // 1320 : 127 - 0x7f -- Sprite 0xa5
      12'h529: dout  = 8'b01111000; // 1321 : 120 - 0x78
      12'h52A: dout  = 8'b00110111; // 1322 :  55 - 0x37
      12'h52B: dout  = 8'b00111011; // 1323 :  59 - 0x3b
      12'h52C: dout  = 8'b00111100; // 1324 :  60 - 0x3c
      12'h52D: dout  = 8'b00011111; // 1325 :  31 - 0x1f
      12'h52E: dout  = 8'b00000111; // 1326 :   7 - 0x7
      12'h52F: dout  = 8'b00000000; // 1327 :   0 - 0x0
      12'h530: dout  = 8'b00000000; // 1328 :   0 - 0x0 -- Sprite 0xa6
      12'h531: dout  = 8'b00000000; // 1329 :   0 - 0x0
      12'h532: dout  = 8'b00000000; // 1330 :   0 - 0x0
      12'h533: dout  = 8'b01110000; // 1331 : 112 - 0x70
      12'h534: dout  = 8'b00000000; // 1332 :   0 - 0x0
      12'h535: dout  = 8'b01010000; // 1333 :  80 - 0x50
      12'h536: dout  = 8'b01010010; // 1334 :  82 - 0x52
      12'h537: dout  = 8'b00000110; // 1335 :   6 - 0x6
      12'h538: dout  = 8'b11111100; // 1336 : 252 - 0xfc -- Sprite 0xa7
      12'h539: dout  = 8'b00011010; // 1337 :  26 - 0x1a
      12'h53A: dout  = 8'b11101100; // 1338 : 236 - 0xec
      12'h53B: dout  = 8'b11011000; // 1339 : 216 - 0xd8
      12'h53C: dout  = 8'b00110100; // 1340 :  52 - 0x34
      12'h53D: dout  = 8'b11101000; // 1341 : 232 - 0xe8
      12'h53E: dout  = 8'b11000000; // 1342 : 192 - 0xc0
      12'h53F: dout  = 8'b00000000; // 1343 :   0 - 0x0
      12'h540: dout  = 8'b00000000; // 1344 :   0 - 0x0 -- Sprite 0xa8
      12'h541: dout  = 8'b00000000; // 1345 :   0 - 0x0
      12'h542: dout  = 8'b00000000; // 1346 :   0 - 0x0
      12'h543: dout  = 8'b00001110; // 1347 :  14 - 0xe
      12'h544: dout  = 8'b00000000; // 1348 :   0 - 0x0
      12'h545: dout  = 8'b00001110; // 1349 :  14 - 0xe
      12'h546: dout  = 8'b01001010; // 1350 :  74 - 0x4a
      12'h547: dout  = 8'b01100000; // 1351 :  96 - 0x60
      12'h548: dout  = 8'b01111111; // 1352 : 127 - 0x7f -- Sprite 0xa9
      12'h549: dout  = 8'b01111100; // 1353 : 124 - 0x7c
      12'h54A: dout  = 8'b01111011; // 1354 : 123 - 0x7b
      12'h54B: dout  = 8'b01110111; // 1355 : 119 - 0x77
      12'h54C: dout  = 8'b01111000; // 1356 : 120 - 0x78
      12'h54D: dout  = 8'b01111111; // 1357 : 127 - 0x7f
      12'h54E: dout  = 8'b01111111; // 1358 : 127 - 0x7f
      12'h54F: dout  = 8'b00000000; // 1359 :   0 - 0x0
      12'h550: dout  = 8'b00000000; // 1360 :   0 - 0x0 -- Sprite 0xaa
      12'h551: dout  = 8'b00000000; // 1361 :   0 - 0x0
      12'h552: dout  = 8'b00000000; // 1362 :   0 - 0x0
      12'h553: dout  = 8'b01110000; // 1363 : 112 - 0x70
      12'h554: dout  = 8'b00000000; // 1364 :   0 - 0x0
      12'h555: dout  = 8'b01110000; // 1365 : 112 - 0x70
      12'h556: dout  = 8'b01010010; // 1366 :  82 - 0x52
      12'h557: dout  = 8'b00000110; // 1367 :   6 - 0x6
      12'h558: dout  = 8'b11111100; // 1368 : 252 - 0xfc -- Sprite 0xab
      12'h559: dout  = 8'b00111010; // 1369 :  58 - 0x3a
      12'h55A: dout  = 8'b11011100; // 1370 : 220 - 0xdc
      12'h55B: dout  = 8'b11101010; // 1371 : 234 - 0xea
      12'h55C: dout  = 8'b00011100; // 1372 :  28 - 0x1c
      12'h55D: dout  = 8'b11111010; // 1373 : 250 - 0xfa
      12'h55E: dout  = 8'b11110100; // 1374 : 244 - 0xf4
      12'h55F: dout  = 8'b00000000; // 1375 :   0 - 0x0
      12'h560: dout  = 8'b00000000; // 1376 :   0 - 0x0 -- Sprite 0xac
      12'h561: dout  = 8'b00000011; // 1377 :   3 - 0x3
      12'h562: dout  = 8'b00001111; // 1378 :  15 - 0xf
      12'h563: dout  = 8'b00001111; // 1379 :  15 - 0xf
      12'h564: dout  = 8'b00011111; // 1380 :  31 - 0x1f
      12'h565: dout  = 8'b01011111; // 1381 :  95 - 0x5f
      12'h566: dout  = 8'b01010000; // 1382 :  80 - 0x50
      12'h567: dout  = 8'b00010000; // 1383 :  16 - 0x10
      12'h568: dout  = 8'b00000000; // 1384 :   0 - 0x0 -- Sprite 0xad
      12'h569: dout  = 8'b11111010; // 1385 : 250 - 0xfa
      12'h56A: dout  = 8'b11111010; // 1386 : 250 - 0xfa
      12'h56B: dout  = 8'b11111010; // 1387 : 250 - 0xfa
      12'h56C: dout  = 8'b10111010; // 1388 : 186 - 0xba
      12'h56D: dout  = 8'b10011010; // 1389 : 154 - 0x9a
      12'h56E: dout  = 8'b00001010; // 1390 :  10 - 0xa
      12'h56F: dout  = 8'b00000010; // 1391 :   2 - 0x2
      12'h570: dout  = 8'b00000000; // 1392 :   0 - 0x0 -- Sprite 0xae
      12'h571: dout  = 8'b00000011; // 1393 :   3 - 0x3
      12'h572: dout  = 8'b00001111; // 1394 :  15 - 0xf
      12'h573: dout  = 8'b00001111; // 1395 :  15 - 0xf
      12'h574: dout  = 8'b00011111; // 1396 :  31 - 0x1f
      12'h575: dout  = 8'b01011111; // 1397 :  95 - 0x5f
      12'h576: dout  = 8'b01010000; // 1398 :  80 - 0x50
      12'h577: dout  = 8'b00010111; // 1399 :  23 - 0x17
      12'h578: dout  = 8'b00000000; // 1400 :   0 - 0x0 -- Sprite 0xaf
      12'h579: dout  = 8'b11111010; // 1401 : 250 - 0xfa
      12'h57A: dout  = 8'b11111010; // 1402 : 250 - 0xfa
      12'h57B: dout  = 8'b11111010; // 1403 : 250 - 0xfa
      12'h57C: dout  = 8'b00111010; // 1404 :  58 - 0x3a
      12'h57D: dout  = 8'b01011010; // 1405 :  90 - 0x5a
      12'h57E: dout  = 8'b01101010; // 1406 : 106 - 0x6a
      12'h57F: dout  = 8'b11110010; // 1407 : 242 - 0xf2
      12'h580: dout  = 8'b00000000; // 1408 :   0 - 0x0 -- Sprite 0xb0
      12'h581: dout  = 8'b00000000; // 1409 :   0 - 0x0
      12'h582: dout  = 8'b00000011; // 1410 :   3 - 0x3
      12'h583: dout  = 8'b00001111; // 1411 :  15 - 0xf
      12'h584: dout  = 8'b00111011; // 1412 :  59 - 0x3b
      12'h585: dout  = 8'b00111111; // 1413 :  63 - 0x3f
      12'h586: dout  = 8'b01101111; // 1414 : 111 - 0x6f
      12'h587: dout  = 8'b01111101; // 1415 : 125 - 0x7d
      12'h588: dout  = 8'b00001111; // 1416 :  15 - 0xf -- Sprite 0xb1
      12'h589: dout  = 8'b01110000; // 1417 : 112 - 0x70
      12'h58A: dout  = 8'b01111111; // 1418 : 127 - 0x7f
      12'h58B: dout  = 8'b00001111; // 1419 :  15 - 0xf
      12'h58C: dout  = 8'b01110000; // 1420 : 112 - 0x70
      12'h58D: dout  = 8'b01111111; // 1421 : 127 - 0x7f
      12'h58E: dout  = 8'b00001111; // 1422 :  15 - 0xf
      12'h58F: dout  = 8'b00000000; // 1423 :   0 - 0x0
      12'h590: dout  = 8'b00000000; // 1424 :   0 - 0x0 -- Sprite 0xb2
      12'h591: dout  = 8'b00000000; // 1425 :   0 - 0x0
      12'h592: dout  = 8'b11000000; // 1426 : 192 - 0xc0
      12'h593: dout  = 8'b11110000; // 1427 : 240 - 0xf0
      12'h594: dout  = 8'b10111100; // 1428 : 188 - 0xbc
      12'h595: dout  = 8'b11110100; // 1429 : 244 - 0xf4
      12'h596: dout  = 8'b11111110; // 1430 : 254 - 0xfe
      12'h597: dout  = 8'b11011110; // 1431 : 222 - 0xde
      12'h598: dout  = 8'b11110000; // 1432 : 240 - 0xf0 -- Sprite 0xb3
      12'h599: dout  = 8'b00001110; // 1433 :  14 - 0xe
      12'h59A: dout  = 8'b11111110; // 1434 : 254 - 0xfe
      12'h59B: dout  = 8'b11110000; // 1435 : 240 - 0xf0
      12'h59C: dout  = 8'b00001110; // 1436 :  14 - 0xe
      12'h59D: dout  = 8'b11111110; // 1437 : 254 - 0xfe
      12'h59E: dout  = 8'b11110000; // 1438 : 240 - 0xf0
      12'h59F: dout  = 8'b00000000; // 1439 :   0 - 0x0
      12'h5A0: dout  = 8'b00000000; // 1440 :   0 - 0x0 -- Sprite 0xb4
      12'h5A1: dout  = 8'b00000000; // 1441 :   0 - 0x0
      12'h5A2: dout  = 8'b00000011; // 1442 :   3 - 0x3
      12'h5A3: dout  = 8'b00001111; // 1443 :  15 - 0xf
      12'h5A4: dout  = 8'b00111011; // 1444 :  59 - 0x3b
      12'h5A5: dout  = 8'b00111111; // 1445 :  63 - 0x3f
      12'h5A6: dout  = 8'b01101111; // 1446 : 111 - 0x6f
      12'h5A7: dout  = 8'b01111101; // 1447 : 125 - 0x7d
      12'h5A8: dout  = 8'b00001111; // 1448 :  15 - 0xf -- Sprite 0xb5
      12'h5A9: dout  = 8'b01110000; // 1449 : 112 - 0x70
      12'h5AA: dout  = 8'b01111111; // 1450 : 127 - 0x7f
      12'h5AB: dout  = 8'b00001111; // 1451 :  15 - 0xf
      12'h5AC: dout  = 8'b01110000; // 1452 : 112 - 0x70
      12'h5AD: dout  = 8'b01111111; // 1453 : 127 - 0x7f
      12'h5AE: dout  = 8'b00001111; // 1454 :  15 - 0xf
      12'h5AF: dout  = 8'b00000000; // 1455 :   0 - 0x0
      12'h5B0: dout  = 8'b00000000; // 1456 :   0 - 0x0 -- Sprite 0xb6
      12'h5B1: dout  = 8'b00000000; // 1457 :   0 - 0x0
      12'h5B2: dout  = 8'b11000000; // 1458 : 192 - 0xc0
      12'h5B3: dout  = 8'b11110000; // 1459 : 240 - 0xf0
      12'h5B4: dout  = 8'b10111100; // 1460 : 188 - 0xbc
      12'h5B5: dout  = 8'b11110100; // 1461 : 244 - 0xf4
      12'h5B6: dout  = 8'b11111110; // 1462 : 254 - 0xfe
      12'h5B7: dout  = 8'b11011110; // 1463 : 222 - 0xde
      12'h5B8: dout  = 8'b11110000; // 1464 : 240 - 0xf0 -- Sprite 0xb7
      12'h5B9: dout  = 8'b00001110; // 1465 :  14 - 0xe
      12'h5BA: dout  = 8'b11111110; // 1466 : 254 - 0xfe
      12'h5BB: dout  = 8'b11110000; // 1467 : 240 - 0xf0
      12'h5BC: dout  = 8'b00001110; // 1468 :  14 - 0xe
      12'h5BD: dout  = 8'b11111110; // 1469 : 254 - 0xfe
      12'h5BE: dout  = 8'b11110000; // 1470 : 240 - 0xf0
      12'h5BF: dout  = 8'b00000000; // 1471 :   0 - 0x0
      12'h5C0: dout  = 8'b00000000; // 1472 :   0 - 0x0 -- Sprite 0xb8
      12'h5C1: dout  = 8'b00000000; // 1473 :   0 - 0x0
      12'h5C2: dout  = 8'b00000011; // 1474 :   3 - 0x3
      12'h5C3: dout  = 8'b00001111; // 1475 :  15 - 0xf
      12'h5C4: dout  = 8'b00111011; // 1476 :  59 - 0x3b
      12'h5C5: dout  = 8'b00111111; // 1477 :  63 - 0x3f
      12'h5C6: dout  = 8'b01101111; // 1478 : 111 - 0x6f
      12'h5C7: dout  = 8'b01111101; // 1479 : 125 - 0x7d
      12'h5C8: dout  = 8'b00001111; // 1480 :  15 - 0xf -- Sprite 0xb9
      12'h5C9: dout  = 8'b00100000; // 1481 :  32 - 0x20
      12'h5CA: dout  = 8'b01010101; // 1482 :  85 - 0x55
      12'h5CB: dout  = 8'b00001010; // 1483 :  10 - 0xa
      12'h5CC: dout  = 8'b01110000; // 1484 : 112 - 0x70
      12'h5CD: dout  = 8'b01111111; // 1485 : 127 - 0x7f
      12'h5CE: dout  = 8'b00001111; // 1486 :  15 - 0xf
      12'h5CF: dout  = 8'b00000000; // 1487 :   0 - 0x0
      12'h5D0: dout  = 8'b00000000; // 1488 :   0 - 0x0 -- Sprite 0xba
      12'h5D1: dout  = 8'b00000000; // 1489 :   0 - 0x0
      12'h5D2: dout  = 8'b11000000; // 1490 : 192 - 0xc0
      12'h5D3: dout  = 8'b11110000; // 1491 : 240 - 0xf0
      12'h5D4: dout  = 8'b10111100; // 1492 : 188 - 0xbc
      12'h5D5: dout  = 8'b11110100; // 1493 : 244 - 0xf4
      12'h5D6: dout  = 8'b11111110; // 1494 : 254 - 0xfe
      12'h5D7: dout  = 8'b11011110; // 1495 : 222 - 0xde
      12'h5D8: dout  = 8'b11110000; // 1496 : 240 - 0xf0 -- Sprite 0xbb
      12'h5D9: dout  = 8'b00001010; // 1497 :  10 - 0xa
      12'h5DA: dout  = 8'b01010100; // 1498 :  84 - 0x54
      12'h5DB: dout  = 8'b10100000; // 1499 : 160 - 0xa0
      12'h5DC: dout  = 8'b00001110; // 1500 :  14 - 0xe
      12'h5DD: dout  = 8'b11111110; // 1501 : 254 - 0xfe
      12'h5DE: dout  = 8'b11110000; // 1502 : 240 - 0xf0
      12'h5DF: dout  = 8'b00000000; // 1503 :   0 - 0x0
      12'h5E0: dout  = 8'b00000000; // 1504 :   0 - 0x0 -- Sprite 0xbc
      12'h5E1: dout  = 8'b01110011; // 1505 : 115 - 0x73
      12'h5E2: dout  = 8'b01111011; // 1506 : 123 - 0x7b
      12'h5E3: dout  = 8'b01111111; // 1507 : 127 - 0x7f
      12'h5E4: dout  = 8'b00111111; // 1508 :  63 - 0x3f
      12'h5E5: dout  = 8'b00011100; // 1509 :  28 - 0x1c
      12'h5E6: dout  = 8'b01111011; // 1510 : 123 - 0x7b
      12'h5E7: dout  = 8'b01111011; // 1511 : 123 - 0x7b
      12'h5E8: dout  = 8'b01111011; // 1512 : 123 - 0x7b -- Sprite 0xbd
      12'h5E9: dout  = 8'b01111011; // 1513 : 123 - 0x7b
      12'h5EA: dout  = 8'b00011100; // 1514 :  28 - 0x1c
      12'h5EB: dout  = 8'b00111111; // 1515 :  63 - 0x3f
      12'h5EC: dout  = 8'b01111111; // 1516 : 127 - 0x7f
      12'h5ED: dout  = 8'b01111011; // 1517 : 123 - 0x7b
      12'h5EE: dout  = 8'b01110011; // 1518 : 115 - 0x73
      12'h5EF: dout  = 8'b00000000; // 1519 :   0 - 0x0
      12'h5F0: dout  = 8'b00000000; // 1520 :   0 - 0x0 -- Sprite 0xbe
      12'h5F1: dout  = 8'b11001110; // 1521 : 206 - 0xce
      12'h5F2: dout  = 8'b11011110; // 1522 : 222 - 0xde
      12'h5F3: dout  = 8'b11111110; // 1523 : 254 - 0xfe
      12'h5F4: dout  = 8'b11111100; // 1524 : 252 - 0xfc
      12'h5F5: dout  = 8'b00111000; // 1525 :  56 - 0x38
      12'h5F6: dout  = 8'b11011110; // 1526 : 222 - 0xde
      12'h5F7: dout  = 8'b11011110; // 1527 : 222 - 0xde
      12'h5F8: dout  = 8'b11011110; // 1528 : 222 - 0xde -- Sprite 0xbf
      12'h5F9: dout  = 8'b11011110; // 1529 : 222 - 0xde
      12'h5FA: dout  = 8'b00111000; // 1530 :  56 - 0x38
      12'h5FB: dout  = 8'b11111100; // 1531 : 252 - 0xfc
      12'h5FC: dout  = 8'b11111110; // 1532 : 254 - 0xfe
      12'h5FD: dout  = 8'b11011110; // 1533 : 222 - 0xde
      12'h5FE: dout  = 8'b11001110; // 1534 : 206 - 0xce
      12'h5FF: dout  = 8'b00000000; // 1535 :   0 - 0x0
      12'h600: dout  = 8'b00000000; // 1536 :   0 - 0x0 -- Sprite 0xc0
      12'h601: dout  = 8'b00000000; // 1537 :   0 - 0x0
      12'h602: dout  = 8'b01000000; // 1538 :  64 - 0x40
      12'h603: dout  = 8'b01100000; // 1539 :  96 - 0x60
      12'h604: dout  = 8'b01100001; // 1540 :  97 - 0x61
      12'h605: dout  = 8'b00000010; // 1541 :   2 - 0x2
      12'h606: dout  = 8'b00000010; // 1542 :   2 - 0x2
      12'h607: dout  = 8'b00000111; // 1543 :   7 - 0x7
      12'h608: dout  = 8'b00000111; // 1544 :   7 - 0x7 -- Sprite 0xc1
      12'h609: dout  = 8'b00000100; // 1545 :   4 - 0x4
      12'h60A: dout  = 8'b00000111; // 1546 :   7 - 0x7
      12'h60B: dout  = 8'b00000001; // 1547 :   1 - 0x1
      12'h60C: dout  = 8'b00000000; // 1548 :   0 - 0x0
      12'h60D: dout  = 8'b00010000; // 1549 :  16 - 0x10
      12'h60E: dout  = 8'b00101000; // 1550 :  40 - 0x28
      12'h60F: dout  = 8'b00000000; // 1551 :   0 - 0x0
      12'h610: dout  = 8'b00000000; // 1552 :   0 - 0x0 -- Sprite 0xc2
      12'h611: dout  = 8'b00000000; // 1553 :   0 - 0x0
      12'h612: dout  = 8'b00000010; // 1554 :   2 - 0x2
      12'h613: dout  = 8'b00000110; // 1555 :   6 - 0x6
      12'h614: dout  = 8'b11100110; // 1556 : 230 - 0xe6
      12'h615: dout  = 8'b10100000; // 1557 : 160 - 0xa0
      12'h616: dout  = 8'b10100000; // 1558 : 160 - 0xa0
      12'h617: dout  = 8'b11110000; // 1559 : 240 - 0xf0
      12'h618: dout  = 8'b11110000; // 1560 : 240 - 0xf0 -- Sprite 0xc3
      12'h619: dout  = 8'b00110000; // 1561 :  48 - 0x30
      12'h61A: dout  = 8'b11000000; // 1562 : 192 - 0xc0
      12'h61B: dout  = 8'b10000000; // 1563 : 128 - 0x80
      12'h61C: dout  = 8'b00000000; // 1564 :   0 - 0x0
      12'h61D: dout  = 8'b00001000; // 1565 :   8 - 0x8
      12'h61E: dout  = 8'b00010100; // 1566 :  20 - 0x14
      12'h61F: dout  = 8'b00000000; // 1567 :   0 - 0x0
      12'h620: dout  = 8'b00000000; // 1568 :   0 - 0x0 -- Sprite 0xc4
      12'h621: dout  = 8'b00000101; // 1569 :   5 - 0x5
      12'h622: dout  = 8'b00000111; // 1570 :   7 - 0x7
      12'h623: dout  = 8'b00000000; // 1571 :   0 - 0x0
      12'h624: dout  = 8'b00000000; // 1572 :   0 - 0x0
      12'h625: dout  = 8'b00000000; // 1573 :   0 - 0x0
      12'h626: dout  = 8'b00000000; // 1574 :   0 - 0x0
      12'h627: dout  = 8'b00000001; // 1575 :   1 - 0x1
      12'h628: dout  = 8'b00000010; // 1576 :   2 - 0x2 -- Sprite 0xc5
      12'h629: dout  = 8'b00000111; // 1577 :   7 - 0x7
      12'h62A: dout  = 8'b00100111; // 1578 :  39 - 0x27
      12'h62B: dout  = 8'b01010011; // 1579 :  83 - 0x53
      12'h62C: dout  = 8'b00000000; // 1580 :   0 - 0x0
      12'h62D: dout  = 8'b00000010; // 1581 :   2 - 0x2
      12'h62E: dout  = 8'b00000101; // 1582 :   5 - 0x5
      12'h62F: dout  = 8'b00000000; // 1583 :   0 - 0x0
      12'h630: dout  = 8'b00000000; // 1584 :   0 - 0x0 -- Sprite 0xc6
      12'h631: dout  = 8'b00000000; // 1585 :   0 - 0x0
      12'h632: dout  = 8'b00000000; // 1586 :   0 - 0x0
      12'h633: dout  = 8'b00000000; // 1587 :   0 - 0x0
      12'h634: dout  = 8'b00000000; // 1588 :   0 - 0x0
      12'h635: dout  = 8'b01100000; // 1589 :  96 - 0x60
      12'h636: dout  = 8'b11011000; // 1590 : 216 - 0xd8
      12'h637: dout  = 8'b10110000; // 1591 : 176 - 0xb0
      12'h638: dout  = 8'b11101000; // 1592 : 232 - 0xe8 -- Sprite 0xc7
      12'h639: dout  = 8'b01111000; // 1593 : 120 - 0x78
      12'h63A: dout  = 8'b10110110; // 1594 : 182 - 0xb6
      12'h63B: dout  = 8'b11100100; // 1595 : 228 - 0xe4
      12'h63C: dout  = 8'b00000110; // 1596 :   6 - 0x6
      12'h63D: dout  = 8'b00000000; // 1597 :   0 - 0x0
      12'h63E: dout  = 8'b00000000; // 1598 :   0 - 0x0
      12'h63F: dout  = 8'b00000000; // 1599 :   0 - 0x0
      12'h640: dout  = 8'b00000000; // 1600 :   0 - 0x0 -- Sprite 0xc8
      12'h641: dout  = 8'b00000000; // 1601 :   0 - 0x0
      12'h642: dout  = 8'b01000000; // 1602 :  64 - 0x40
      12'h643: dout  = 8'b00100000; // 1603 :  32 - 0x20
      12'h644: dout  = 8'b01000000; // 1604 :  64 - 0x40
      12'h645: dout  = 8'b00000111; // 1605 :   7 - 0x7
      12'h646: dout  = 8'b00000101; // 1606 :   5 - 0x5
      12'h647: dout  = 8'b00001101; // 1607 :  13 - 0xd
      12'h648: dout  = 8'b00001101; // 1608 :  13 - 0xd -- Sprite 0xc9
      12'h649: dout  = 8'b00000101; // 1609 :   5 - 0x5
      12'h64A: dout  = 8'b00000011; // 1610 :   3 - 0x3
      12'h64B: dout  = 8'b01000011; // 1611 :  67 - 0x43
      12'h64C: dout  = 8'b00100000; // 1612 :  32 - 0x20
      12'h64D: dout  = 8'b01000000; // 1613 :  64 - 0x40
      12'h64E: dout  = 8'b00000000; // 1614 :   0 - 0x0
      12'h64F: dout  = 8'b00000000; // 1615 :   0 - 0x0
      12'h650: dout  = 8'b00000000; // 1616 :   0 - 0x0 -- Sprite 0xca
      12'h651: dout  = 8'b00011100; // 1617 :  28 - 0x1c
      12'h652: dout  = 8'b00011000; // 1618 :  24 - 0x18
      12'h653: dout  = 8'b00000000; // 1619 :   0 - 0x0
      12'h654: dout  = 8'b00000000; // 1620 :   0 - 0x0
      12'h655: dout  = 8'b10000000; // 1621 : 128 - 0x80
      12'h656: dout  = 8'b11100000; // 1622 : 224 - 0xe0
      12'h657: dout  = 8'b10010000; // 1623 : 144 - 0x90
      12'h658: dout  = 8'b11110000; // 1624 : 240 - 0xf0 -- Sprite 0xcb
      12'h659: dout  = 8'b10010000; // 1625 : 144 - 0x90
      12'h65A: dout  = 8'b11110000; // 1626 : 240 - 0xf0
      12'h65B: dout  = 8'b10000000; // 1627 : 128 - 0x80
      12'h65C: dout  = 8'b00000000; // 1628 :   0 - 0x0
      12'h65D: dout  = 8'b00011000; // 1629 :  24 - 0x18
      12'h65E: dout  = 8'b00011100; // 1630 :  28 - 0x1c
      12'h65F: dout  = 8'b00000000; // 1631 :   0 - 0x0
      12'h660: dout  = 8'b00000000; // 1632 :   0 - 0x0 -- Sprite 0xcc
      12'h661: dout  = 8'b00001000; // 1633 :   8 - 0x8
      12'h662: dout  = 8'b00000100; // 1634 :   4 - 0x4
      12'h663: dout  = 8'b00001000; // 1635 :   8 - 0x8
      12'h664: dout  = 8'b00000000; // 1636 :   0 - 0x0
      12'h665: dout  = 8'b01000110; // 1637 :  70 - 0x46
      12'h666: dout  = 8'b00101111; // 1638 :  47 - 0x2f
      12'h667: dout  = 8'b01001110; // 1639 :  78 - 0x4e
      12'h668: dout  = 8'b00001101; // 1640 :  13 - 0xd -- Sprite 0xcd
      12'h669: dout  = 8'b00001011; // 1641 :  11 - 0xb
      12'h66A: dout  = 8'b00001111; // 1642 :  15 - 0xf
      12'h66B: dout  = 8'b00000110; // 1643 :   6 - 0x6
      12'h66C: dout  = 8'b00000011; // 1644 :   3 - 0x3
      12'h66D: dout  = 8'b00011100; // 1645 :  28 - 0x1c
      12'h66E: dout  = 8'b00010100; // 1646 :  20 - 0x14
      12'h66F: dout  = 8'b00000000; // 1647 :   0 - 0x0
      12'h670: dout  = 8'b00000000; // 1648 :   0 - 0x0 -- Sprite 0xce
      12'h671: dout  = 8'b00000000; // 1649 :   0 - 0x0
      12'h672: dout  = 8'b00000000; // 1650 :   0 - 0x0
      12'h673: dout  = 8'b00000000; // 1651 :   0 - 0x0
      12'h674: dout  = 8'b00000000; // 1652 :   0 - 0x0
      12'h675: dout  = 8'b00000110; // 1653 :   6 - 0x6
      12'h676: dout  = 8'b00000100; // 1654 :   4 - 0x4
      12'h677: dout  = 8'b10000110; // 1655 : 134 - 0x86
      12'h678: dout  = 8'b11000000; // 1656 : 192 - 0xc0 -- Sprite 0xcf
      12'h679: dout  = 8'b01100000; // 1657 :  96 - 0x60
      12'h67A: dout  = 8'b10100000; // 1658 : 160 - 0xa0
      12'h67B: dout  = 8'b11000000; // 1659 : 192 - 0xc0
      12'h67C: dout  = 8'b01000000; // 1660 :  64 - 0x40
      12'h67D: dout  = 8'b00000000; // 1661 :   0 - 0x0
      12'h67E: dout  = 8'b00000000; // 1662 :   0 - 0x0
      12'h67F: dout  = 8'b00000000; // 1663 :   0 - 0x0
      12'h680: dout  = 8'b00000000; // 1664 :   0 - 0x0 -- Sprite 0xd0
      12'h681: dout  = 8'b00000000; // 1665 :   0 - 0x0
      12'h682: dout  = 8'b00000000; // 1666 :   0 - 0x0
      12'h683: dout  = 8'b00000000; // 1667 :   0 - 0x0
      12'h684: dout  = 8'b00000100; // 1668 :   4 - 0x4
      12'h685: dout  = 8'b00001110; // 1669 :  14 - 0xe
      12'h686: dout  = 8'b00111111; // 1670 :  63 - 0x3f
      12'h687: dout  = 8'b00111001; // 1671 :  57 - 0x39
      12'h688: dout  = 8'b01110000; // 1672 : 112 - 0x70 -- Sprite 0xd1
      12'h689: dout  = 8'b01111000; // 1673 : 120 - 0x78
      12'h68A: dout  = 8'b00111111; // 1674 :  63 - 0x3f
      12'h68B: dout  = 8'b00111111; // 1675 :  63 - 0x3f
      12'h68C: dout  = 8'b00000011; // 1676 :   3 - 0x3
      12'h68D: dout  = 8'b00001100; // 1677 :  12 - 0xc
      12'h68E: dout  = 8'b00001110; // 1678 :  14 - 0xe
      12'h68F: dout  = 8'b00000000; // 1679 :   0 - 0x0
      12'h690: dout  = 8'b00000000; // 1680 :   0 - 0x0 -- Sprite 0xd2
      12'h691: dout  = 8'b00000000; // 1681 :   0 - 0x0
      12'h692: dout  = 8'b00000000; // 1682 :   0 - 0x0
      12'h693: dout  = 8'b00001000; // 1683 :   8 - 0x8
      12'h694: dout  = 8'b11011000; // 1684 : 216 - 0xd8
      12'h695: dout  = 8'b11111100; // 1685 : 252 - 0xfc
      12'h696: dout  = 8'b11111100; // 1686 : 252 - 0xfc
      12'h697: dout  = 8'b10011100; // 1687 : 156 - 0x9c
      12'h698: dout  = 8'b00001100; // 1688 :  12 - 0xc -- Sprite 0xd3
      12'h699: dout  = 8'b10011100; // 1689 : 156 - 0x9c
      12'h69A: dout  = 8'b11111000; // 1690 : 248 - 0xf8
      12'h69B: dout  = 8'b01111000; // 1691 : 120 - 0x78
      12'h69C: dout  = 8'b10001000; // 1692 : 136 - 0x88
      12'h69D: dout  = 8'b00110000; // 1693 :  48 - 0x30
      12'h69E: dout  = 8'b00111000; // 1694 :  56 - 0x38
      12'h69F: dout  = 8'b00000000; // 1695 :   0 - 0x0
      12'h6A0: dout  = 8'b00000000; // 1696 :   0 - 0x0 -- Sprite 0xd4
      12'h6A1: dout  = 8'b00000000; // 1697 :   0 - 0x0
      12'h6A2: dout  = 8'b00000000; // 1698 :   0 - 0x0
      12'h6A3: dout  = 8'b00000000; // 1699 :   0 - 0x0
      12'h6A4: dout  = 8'b00000001; // 1700 :   1 - 0x1
      12'h6A5: dout  = 8'b00001011; // 1701 :  11 - 0xb
      12'h6A6: dout  = 8'b00011111; // 1702 :  31 - 0x1f
      12'h6A7: dout  = 8'b00111001; // 1703 :  57 - 0x39
      12'h6A8: dout  = 8'b01110000; // 1704 : 112 - 0x70 -- Sprite 0xd5
      12'h6A9: dout  = 8'b01111000; // 1705 : 120 - 0x78
      12'h6AA: dout  = 8'b00111111; // 1706 :  63 - 0x3f
      12'h6AB: dout  = 8'b00111111; // 1707 :  63 - 0x3f
      12'h6AC: dout  = 8'b00000011; // 1708 :   3 - 0x3
      12'h6AD: dout  = 8'b00111000; // 1709 :  56 - 0x38
      12'h6AE: dout  = 8'b00011100; // 1710 :  28 - 0x1c
      12'h6AF: dout  = 8'b00000000; // 1711 :   0 - 0x0
      12'h6B0: dout  = 8'b00000000; // 1712 :   0 - 0x0 -- Sprite 0xd6
      12'h6B1: dout  = 8'b00000000; // 1713 :   0 - 0x0
      12'h6B2: dout  = 8'b00000000; // 1714 :   0 - 0x0
      12'h6B3: dout  = 8'b11000000; // 1715 : 192 - 0xc0
      12'h6B4: dout  = 8'b11001000; // 1716 : 200 - 0xc8
      12'h6B5: dout  = 8'b11111000; // 1717 : 248 - 0xf8
      12'h6B6: dout  = 8'b11111100; // 1718 : 252 - 0xfc
      12'h6B7: dout  = 8'b10011100; // 1719 : 156 - 0x9c
      12'h6B8: dout  = 8'b00001100; // 1720 :  12 - 0xc -- Sprite 0xd7
      12'h6B9: dout  = 8'b10011100; // 1721 : 156 - 0x9c
      12'h6BA: dout  = 8'b11111000; // 1722 : 248 - 0xf8
      12'h6BB: dout  = 8'b01111000; // 1723 : 120 - 0x78
      12'h6BC: dout  = 8'b11100010; // 1724 : 226 - 0xe2
      12'h6BD: dout  = 8'b00011110; // 1725 :  30 - 0x1e
      12'h6BE: dout  = 8'b00001100; // 1726 :  12 - 0xc
      12'h6BF: dout  = 8'b00000000; // 1727 :   0 - 0x0
      12'h6C0: dout  = 8'b00000000; // 1728 :   0 - 0x0 -- Sprite 0xd8
      12'h6C1: dout  = 8'b00110000; // 1729 :  48 - 0x30
      12'h6C2: dout  = 8'b00111100; // 1730 :  60 - 0x3c
      12'h6C3: dout  = 8'b01111100; // 1731 : 124 - 0x7c
      12'h6C4: dout  = 8'b01111100; // 1732 : 124 - 0x7c
      12'h6C5: dout  = 8'b00111110; // 1733 :  62 - 0x3e
      12'h6C6: dout  = 8'b00011100; // 1734 :  28 - 0x1c
      12'h6C7: dout  = 8'b00000000; // 1735 :   0 - 0x0
      12'h6C8: dout  = 8'b00000000; // 1736 :   0 - 0x0 -- Sprite 0xd9
      12'h6C9: dout  = 8'b00001110; // 1737 :  14 - 0xe
      12'h6CA: dout  = 8'b00111110; // 1738 :  62 - 0x3e
      12'h6CB: dout  = 8'b01111110; // 1739 : 126 - 0x7e
      12'h6CC: dout  = 8'b01111110; // 1740 : 126 - 0x7e
      12'h6CD: dout  = 8'b00111100; // 1741 :  60 - 0x3c
      12'h6CE: dout  = 8'b00001100; // 1742 :  12 - 0xc
      12'h6CF: dout  = 8'b00000000; // 1743 :   0 - 0x0
      12'h6D0: dout  = 8'b00000000; // 1744 :   0 - 0x0 -- Sprite 0xda
      12'h6D1: dout  = 8'b00100000; // 1745 :  32 - 0x20
      12'h6D2: dout  = 8'b01111110; // 1746 : 126 - 0x7e
      12'h6D3: dout  = 8'b01111110; // 1747 : 126 - 0x7e
      12'h6D4: dout  = 8'b01111110; // 1748 : 126 - 0x7e
      12'h6D5: dout  = 8'b00111100; // 1749 :  60 - 0x3c
      12'h6D6: dout  = 8'b00111000; // 1750 :  56 - 0x38
      12'h6D7: dout  = 8'b00000000; // 1751 :   0 - 0x0
      12'h6D8: dout  = 8'b00000000; // 1752 :   0 - 0x0 -- Sprite 0xdb
      12'h6D9: dout  = 8'b00011100; // 1753 :  28 - 0x1c
      12'h6DA: dout  = 8'b00111110; // 1754 :  62 - 0x3e
      12'h6DB: dout  = 8'b01111110; // 1755 : 126 - 0x7e
      12'h6DC: dout  = 8'b01111110; // 1756 : 126 - 0x7e
      12'h6DD: dout  = 8'b00111100; // 1757 :  60 - 0x3c
      12'h6DE: dout  = 8'b00010000; // 1758 :  16 - 0x10
      12'h6DF: dout  = 8'b00000000; // 1759 :   0 - 0x0
      12'h6E0: dout  = 8'b00000000; // 1760 :   0 - 0x0 -- Sprite 0xdc
      12'h6E1: dout  = 8'b00000000; // 1761 :   0 - 0x0
      12'h6E2: dout  = 8'b00000000; // 1762 :   0 - 0x0
      12'h6E3: dout  = 8'b00000001; // 1763 :   1 - 0x1
      12'h6E4: dout  = 8'b00000011; // 1764 :   3 - 0x3
      12'h6E5: dout  = 8'b00000001; // 1765 :   1 - 0x1
      12'h6E6: dout  = 8'b00000001; // 1766 :   1 - 0x1
      12'h6E7: dout  = 8'b00001111; // 1767 :  15 - 0xf
      12'h6E8: dout  = 8'b00000111; // 1768 :   7 - 0x7 -- Sprite 0xdd
      12'h6E9: dout  = 8'b00000111; // 1769 :   7 - 0x7
      12'h6EA: dout  = 8'b00000111; // 1770 :   7 - 0x7
      12'h6EB: dout  = 8'b00011111; // 1771 :  31 - 0x1f
      12'h6EC: dout  = 8'b00001111; // 1772 :  15 - 0xf
      12'h6ED: dout  = 8'b00000111; // 1773 :   7 - 0x7
      12'h6EE: dout  = 8'b00000011; // 1774 :   3 - 0x3
      12'h6EF: dout  = 8'b00000000; // 1775 :   0 - 0x0
      12'h6F0: dout  = 8'b00000000; // 1776 :   0 - 0x0 -- Sprite 0xde
      12'h6F1: dout  = 8'b00000000; // 1777 :   0 - 0x0
      12'h6F2: dout  = 8'b00000000; // 1778 :   0 - 0x0
      12'h6F3: dout  = 8'b00000000; // 1779 :   0 - 0x0
      12'h6F4: dout  = 8'b10000000; // 1780 : 128 - 0x80
      12'h6F5: dout  = 8'b10000000; // 1781 : 128 - 0x80
      12'h6F6: dout  = 8'b10010000; // 1782 : 144 - 0x90
      12'h6F7: dout  = 8'b11110000; // 1783 : 240 - 0xf0
      12'h6F8: dout  = 8'b11100000; // 1784 : 224 - 0xe0 -- Sprite 0xdf
      12'h6F9: dout  = 8'b11100000; // 1785 : 224 - 0xe0
      12'h6FA: dout  = 8'b11110000; // 1786 : 240 - 0xf0
      12'h6FB: dout  = 8'b11110000; // 1787 : 240 - 0xf0
      12'h6FC: dout  = 8'b11100000; // 1788 : 224 - 0xe0
      12'h6FD: dout  = 8'b11000000; // 1789 : 192 - 0xc0
      12'h6FE: dout  = 8'b11000000; // 1790 : 192 - 0xc0
      12'h6FF: dout  = 8'b00000000; // 1791 :   0 - 0x0
      12'h700: dout  = 8'b00001111; // 1792 :  15 - 0xf -- Sprite 0xe0
      12'h701: dout  = 8'b00011111; // 1793 :  31 - 0x1f
      12'h702: dout  = 8'b00011111; // 1794 :  31 - 0x1f
      12'h703: dout  = 8'b00111111; // 1795 :  63 - 0x3f
      12'h704: dout  = 8'b01111111; // 1796 : 127 - 0x7f
      12'h705: dout  = 8'b11111111; // 1797 : 255 - 0xff
      12'h706: dout  = 8'b11111111; // 1798 : 255 - 0xff
      12'h707: dout  = 8'b11111111; // 1799 : 255 - 0xff
      12'h708: dout  = 8'b11111111; // 1800 : 255 - 0xff -- Sprite 0xe1
      12'h709: dout  = 8'b11111111; // 1801 : 255 - 0xff
      12'h70A: dout  = 8'b01111111; // 1802 : 127 - 0x7f
      12'h70B: dout  = 8'b00111111; // 1803 :  63 - 0x3f
      12'h70C: dout  = 8'b00111111; // 1804 :  63 - 0x3f
      12'h70D: dout  = 8'b00011111; // 1805 :  31 - 0x1f
      12'h70E: dout  = 8'b00001111; // 1806 :  15 - 0xf
      12'h70F: dout  = 8'b00000111; // 1807 :   7 - 0x7
      12'h710: dout  = 8'b11111110; // 1808 : 254 - 0xfe -- Sprite 0xe2
      12'h711: dout  = 8'b11111111; // 1809 : 255 - 0xff
      12'h712: dout  = 8'b11111111; // 1810 : 255 - 0xff
      12'h713: dout  = 8'b00001111; // 1811 :  15 - 0xf
      12'h714: dout  = 8'b10111111; // 1812 : 191 - 0xbf
      12'h715: dout  = 8'b10100011; // 1813 : 163 - 0xa3
      12'h716: dout  = 8'b11110111; // 1814 : 247 - 0xf7
      12'h717: dout  = 8'b11110111; // 1815 : 247 - 0xf7
      12'h718: dout  = 8'b11111111; // 1816 : 255 - 0xff -- Sprite 0xe3
      12'h719: dout  = 8'b11111111; // 1817 : 255 - 0xff
      12'h71A: dout  = 8'b00111111; // 1818 :  63 - 0x3f
      12'h71B: dout  = 8'b00011111; // 1819 :  31 - 0x1f
      12'h71C: dout  = 8'b11111110; // 1820 : 254 - 0xfe
      12'h71D: dout  = 8'b11111100; // 1821 : 252 - 0xfc
      12'h71E: dout  = 8'b11111000; // 1822 : 248 - 0xf8
      12'h71F: dout  = 8'b11110000; // 1823 : 240 - 0xf0
      12'h720: dout  = 8'b00001111; // 1824 :  15 - 0xf -- Sprite 0xe4
      12'h721: dout  = 8'b00011111; // 1825 :  31 - 0x1f
      12'h722: dout  = 8'b00011111; // 1826 :  31 - 0x1f
      12'h723: dout  = 8'b00111111; // 1827 :  63 - 0x3f
      12'h724: dout  = 8'b01111111; // 1828 : 127 - 0x7f
      12'h725: dout  = 8'b11111111; // 1829 : 255 - 0xff
      12'h726: dout  = 8'b11111111; // 1830 : 255 - 0xff
      12'h727: dout  = 8'b11111111; // 1831 : 255 - 0xff
      12'h728: dout  = 8'b11111111; // 1832 : 255 - 0xff -- Sprite 0xe5
      12'h729: dout  = 8'b11111111; // 1833 : 255 - 0xff
      12'h72A: dout  = 8'b01111110; // 1834 : 126 - 0x7e
      12'h72B: dout  = 8'b00111111; // 1835 :  63 - 0x3f
      12'h72C: dout  = 8'b00111111; // 1836 :  63 - 0x3f
      12'h72D: dout  = 8'b00011111; // 1837 :  31 - 0x1f
      12'h72E: dout  = 8'b00001111; // 1838 :  15 - 0xf
      12'h72F: dout  = 8'b00000111; // 1839 :   7 - 0x7
      12'h730: dout  = 8'b11111110; // 1840 : 254 - 0xfe -- Sprite 0xe6
      12'h731: dout  = 8'b11111111; // 1841 : 255 - 0xff
      12'h732: dout  = 8'b11111111; // 1842 : 255 - 0xff
      12'h733: dout  = 8'b11100011; // 1843 : 227 - 0xe3
      12'h734: dout  = 8'b00010111; // 1844 :  23 - 0x17
      12'h735: dout  = 8'b10110111; // 1845 : 183 - 0xb7
      12'h736: dout  = 8'b10111111; // 1846 : 191 - 0xbf
      12'h737: dout  = 8'b11111111; // 1847 : 255 - 0xff
      12'h738: dout  = 8'b11111111; // 1848 : 255 - 0xff -- Sprite 0xe7
      12'h739: dout  = 8'b11111111; // 1849 : 255 - 0xff
      12'h73A: dout  = 8'b00111111; // 1850 :  63 - 0x3f
      12'h73B: dout  = 8'b00001111; // 1851 :  15 - 0xf
      12'h73C: dout  = 8'b00001110; // 1852 :  14 - 0xe
      12'h73D: dout  = 8'b11111100; // 1853 : 252 - 0xfc
      12'h73E: dout  = 8'b11111000; // 1854 : 248 - 0xf8
      12'h73F: dout  = 8'b11110000; // 1855 : 240 - 0xf0
      12'h740: dout  = 8'b00000000; // 1856 :   0 - 0x0 -- Sprite 0xe8
      12'h741: dout  = 8'b00000101; // 1857 :   5 - 0x5
      12'h742: dout  = 8'b00000111; // 1858 :   7 - 0x7
      12'h743: dout  = 8'b00000011; // 1859 :   3 - 0x3
      12'h744: dout  = 8'b00000000; // 1860 :   0 - 0x0
      12'h745: dout  = 8'b00000000; // 1861 :   0 - 0x0
      12'h746: dout  = 8'b00000000; // 1862 :   0 - 0x0
      12'h747: dout  = 8'b00000000; // 1863 :   0 - 0x0
      12'h748: dout  = 8'b00000000; // 1864 :   0 - 0x0 -- Sprite 0xe9
      12'h749: dout  = 8'b00000000; // 1865 :   0 - 0x0
      12'h74A: dout  = 8'b00000000; // 1866 :   0 - 0x0
      12'h74B: dout  = 8'b00000000; // 1867 :   0 - 0x0
      12'h74C: dout  = 8'b00000000; // 1868 :   0 - 0x0
      12'h74D: dout  = 8'b00000000; // 1869 :   0 - 0x0
      12'h74E: dout  = 8'b00000000; // 1870 :   0 - 0x0
      12'h74F: dout  = 8'b00000000; // 1871 :   0 - 0x0
      12'h750: dout  = 8'b00000011; // 1872 :   3 - 0x3 -- Sprite 0xea
      12'h751: dout  = 8'b10011110; // 1873 : 158 - 0x9e
      12'h752: dout  = 8'b00001110; // 1874 :  14 - 0xe
      12'h753: dout  = 8'b00000000; // 1875 :   0 - 0x0
      12'h754: dout  = 8'b00000000; // 1876 :   0 - 0x0
      12'h755: dout  = 8'b00000000; // 1877 :   0 - 0x0
      12'h756: dout  = 8'b00000000; // 1878 :   0 - 0x0
      12'h757: dout  = 8'b00000000; // 1879 :   0 - 0x0
      12'h758: dout  = 8'b00000000; // 1880 :   0 - 0x0 -- Sprite 0xeb
      12'h759: dout  = 8'b00000000; // 1881 :   0 - 0x0
      12'h75A: dout  = 8'b00000000; // 1882 :   0 - 0x0
      12'h75B: dout  = 8'b00000000; // 1883 :   0 - 0x0
      12'h75C: dout  = 8'b00000000; // 1884 :   0 - 0x0
      12'h75D: dout  = 8'b00000000; // 1885 :   0 - 0x0
      12'h75E: dout  = 8'b00000000; // 1886 :   0 - 0x0
      12'h75F: dout  = 8'b00000000; // 1887 :   0 - 0x0
      12'h760: dout  = 8'b00000000; // 1888 :   0 - 0x0 -- Sprite 0xec
      12'h761: dout  = 8'b00000000; // 1889 :   0 - 0x0
      12'h762: dout  = 8'b00000000; // 1890 :   0 - 0x0
      12'h763: dout  = 8'b00000000; // 1891 :   0 - 0x0
      12'h764: dout  = 8'b00000100; // 1892 :   4 - 0x4
      12'h765: dout  = 8'b00001110; // 1893 :  14 - 0xe
      12'h766: dout  = 8'b00001111; // 1894 :  15 - 0xf
      12'h767: dout  = 8'b00001011; // 1895 :  11 - 0xb
      12'h768: dout  = 8'b00001111; // 1896 :  15 - 0xf -- Sprite 0xed
      12'h769: dout  = 8'b00001100; // 1897 :  12 - 0xc
      12'h76A: dout  = 8'b00001111; // 1898 :  15 - 0xf
      12'h76B: dout  = 8'b00001111; // 1899 :  15 - 0xf
      12'h76C: dout  = 8'b00000000; // 1900 :   0 - 0x0
      12'h76D: dout  = 8'b01111111; // 1901 : 127 - 0x7f
      12'h76E: dout  = 8'b11010101; // 1902 : 213 - 0xd5
      12'h76F: dout  = 8'b01111111; // 1903 : 127 - 0x7f
      12'h770: dout  = 8'b00000000; // 1904 :   0 - 0x0 -- Sprite 0xee
      12'h771: dout  = 8'b00000000; // 1905 :   0 - 0x0
      12'h772: dout  = 8'b00000000; // 1906 :   0 - 0x0
      12'h773: dout  = 8'b00000000; // 1907 :   0 - 0x0
      12'h774: dout  = 8'b00100000; // 1908 :  32 - 0x20
      12'h775: dout  = 8'b01110000; // 1909 : 112 - 0x70
      12'h776: dout  = 8'b11110000; // 1910 : 240 - 0xf0
      12'h777: dout  = 8'b11100000; // 1911 : 224 - 0xe0
      12'h778: dout  = 8'b11110000; // 1912 : 240 - 0xf0 -- Sprite 0xef
      12'h779: dout  = 8'b00110000; // 1913 :  48 - 0x30
      12'h77A: dout  = 8'b11110000; // 1914 : 240 - 0xf0
      12'h77B: dout  = 8'b11110000; // 1915 : 240 - 0xf0
      12'h77C: dout  = 8'b00000000; // 1916 :   0 - 0x0
      12'h77D: dout  = 8'b11111110; // 1917 : 254 - 0xfe
      12'h77E: dout  = 8'b01010101; // 1918 :  85 - 0x55
      12'h77F: dout  = 8'b11111110; // 1919 : 254 - 0xfe
      12'h780: dout  = 8'b00000000; // 1920 :   0 - 0x0 -- Sprite 0xf0
      12'h781: dout  = 8'b00000000; // 1921 :   0 - 0x0
      12'h782: dout  = 8'b00000000; // 1922 :   0 - 0x0
      12'h783: dout  = 8'b00000000; // 1923 :   0 - 0x0
      12'h784: dout  = 8'b00000100; // 1924 :   4 - 0x4
      12'h785: dout  = 8'b00001110; // 1925 :  14 - 0xe
      12'h786: dout  = 8'b00001111; // 1926 :  15 - 0xf
      12'h787: dout  = 8'b00001011; // 1927 :  11 - 0xb
      12'h788: dout  = 8'b00001111; // 1928 :  15 - 0xf -- Sprite 0xf1
      12'h789: dout  = 8'b00001100; // 1929 :  12 - 0xc
      12'h78A: dout  = 8'b00001111; // 1930 :  15 - 0xf
      12'h78B: dout  = 8'b00001111; // 1931 :  15 - 0xf
      12'h78C: dout  = 8'b00000000; // 1932 :   0 - 0x0
      12'h78D: dout  = 8'b01111111; // 1933 : 127 - 0x7f
      12'h78E: dout  = 8'b10101010; // 1934 : 170 - 0xaa
      12'h78F: dout  = 8'b01111111; // 1935 : 127 - 0x7f
      12'h790: dout  = 8'b00000000; // 1936 :   0 - 0x0 -- Sprite 0xf2
      12'h791: dout  = 8'b00000000; // 1937 :   0 - 0x0
      12'h792: dout  = 8'b00000000; // 1938 :   0 - 0x0
      12'h793: dout  = 8'b00000000; // 1939 :   0 - 0x0
      12'h794: dout  = 8'b00100000; // 1940 :  32 - 0x20
      12'h795: dout  = 8'b01110000; // 1941 : 112 - 0x70
      12'h796: dout  = 8'b11110000; // 1942 : 240 - 0xf0
      12'h797: dout  = 8'b11100000; // 1943 : 224 - 0xe0
      12'h798: dout  = 8'b11110000; // 1944 : 240 - 0xf0 -- Sprite 0xf3
      12'h799: dout  = 8'b00110000; // 1945 :  48 - 0x30
      12'h79A: dout  = 8'b11110000; // 1946 : 240 - 0xf0
      12'h79B: dout  = 8'b11110000; // 1947 : 240 - 0xf0
      12'h79C: dout  = 8'b00000000; // 1948 :   0 - 0x0
      12'h79D: dout  = 8'b11111110; // 1949 : 254 - 0xfe
      12'h79E: dout  = 8'b10101011; // 1950 : 171 - 0xab
      12'h79F: dout  = 8'b11111110; // 1951 : 254 - 0xfe
      12'h7A0: dout  = 8'b00000000; // 1952 :   0 - 0x0 -- Sprite 0xf4
      12'h7A1: dout  = 8'b00010101; // 1953 :  21 - 0x15
      12'h7A2: dout  = 8'b00001010; // 1954 :  10 - 0xa
      12'h7A3: dout  = 8'b00000101; // 1955 :   5 - 0x5
      12'h7A4: dout  = 8'b00000010; // 1956 :   2 - 0x2
      12'h7A5: dout  = 8'b00000101; // 1957 :   5 - 0x5
      12'h7A6: dout  = 8'b00000111; // 1958 :   7 - 0x7
      12'h7A7: dout  = 8'b00000111; // 1959 :   7 - 0x7
      12'h7A8: dout  = 8'b00111100; // 1960 :  60 - 0x3c -- Sprite 0xf5
      12'h7A9: dout  = 8'b01111011; // 1961 : 123 - 0x7b
      12'h7AA: dout  = 8'b01111011; // 1962 : 123 - 0x7b
      12'h7AB: dout  = 8'b01111111; // 1963 : 127 - 0x7f
      12'h7AC: dout  = 8'b01111110; // 1964 : 126 - 0x7e
      12'h7AD: dout  = 8'b01111111; // 1965 : 127 - 0x7f
      12'h7AE: dout  = 8'b00111110; // 1966 :  62 - 0x3e
      12'h7AF: dout  = 8'b00000000; // 1967 :   0 - 0x0
      12'h7B0: dout  = 8'b00000000; // 1968 :   0 - 0x0 -- Sprite 0xf6
      12'h7B1: dout  = 8'b01010000; // 1969 :  80 - 0x50
      12'h7B2: dout  = 8'b10100000; // 1970 : 160 - 0xa0
      12'h7B3: dout  = 8'b01000000; // 1971 :  64 - 0x40
      12'h7B4: dout  = 8'b10100000; // 1972 : 160 - 0xa0
      12'h7B5: dout  = 8'b01000000; // 1973 :  64 - 0x40
      12'h7B6: dout  = 8'b11100000; // 1974 : 224 - 0xe0
      12'h7B7: dout  = 8'b11100000; // 1975 : 224 - 0xe0
      12'h7B8: dout  = 8'b01111000; // 1976 : 120 - 0x78 -- Sprite 0xf7
      12'h7B9: dout  = 8'b10111100; // 1977 : 188 - 0xbc
      12'h7BA: dout  = 8'b10111000; // 1978 : 184 - 0xb8
      12'h7BB: dout  = 8'b10111110; // 1979 : 190 - 0xbe
      12'h7BC: dout  = 8'b01111100; // 1980 : 124 - 0x7c
      12'h7BD: dout  = 8'b11111110; // 1981 : 254 - 0xfe
      12'h7BE: dout  = 8'b01111000; // 1982 : 120 - 0x78
      12'h7BF: dout  = 8'b00000000; // 1983 :   0 - 0x0
      12'h7C0: dout  = 8'b00000011; // 1984 :   3 - 0x3 -- Sprite 0xf8
      12'h7C1: dout  = 8'b00000011; // 1985 :   3 - 0x3
      12'h7C2: dout  = 8'b00000000; // 1986 :   0 - 0x0
      12'h7C3: dout  = 8'b00000011; // 1987 :   3 - 0x3
      12'h7C4: dout  = 8'b00000111; // 1988 :   7 - 0x7
      12'h7C5: dout  = 8'b00000110; // 1989 :   6 - 0x6
      12'h7C6: dout  = 8'b00000111; // 1990 :   7 - 0x7
      12'h7C7: dout  = 8'b00000000; // 1991 :   0 - 0x0
      12'h7C8: dout  = 8'b00000000; // 1992 :   0 - 0x0 -- Sprite 0xf9
      12'h7C9: dout  = 8'b00011111; // 1993 :  31 - 0x1f
      12'h7CA: dout  = 8'b00011111; // 1994 :  31 - 0x1f
      12'h7CB: dout  = 8'b00001111; // 1995 :  15 - 0xf
      12'h7CC: dout  = 8'b00000011; // 1996 :   3 - 0x3
      12'h7CD: dout  = 8'b00000000; // 1997 :   0 - 0x0
      12'h7CE: dout  = 8'b00000000; // 1998 :   0 - 0x0
      12'h7CF: dout  = 8'b00000000; // 1999 :   0 - 0x0
      12'h7D0: dout  = 8'b11100000; // 2000 : 224 - 0xe0 -- Sprite 0xfa
      12'h7D1: dout  = 8'b11100000; // 2001 : 224 - 0xe0
      12'h7D2: dout  = 8'b00000000; // 2002 :   0 - 0x0
      12'h7D3: dout  = 8'b00110000; // 2003 :  48 - 0x30
      12'h7D4: dout  = 8'b01110000; // 2004 : 112 - 0x70
      12'h7D5: dout  = 8'b01100000; // 2005 :  96 - 0x60
      12'h7D6: dout  = 8'b01110000; // 2006 : 112 - 0x70
      12'h7D7: dout  = 8'b00000000; // 2007 :   0 - 0x0
      12'h7D8: dout  = 8'b00000000; // 2008 :   0 - 0x0 -- Sprite 0xfb
      12'h7D9: dout  = 8'b11111000; // 2009 : 248 - 0xf8
      12'h7DA: dout  = 8'b11111000; // 2010 : 248 - 0xf8
      12'h7DB: dout  = 8'b11110000; // 2011 : 240 - 0xf0
      12'h7DC: dout  = 8'b11000000; // 2012 : 192 - 0xc0
      12'h7DD: dout  = 8'b00000000; // 2013 :   0 - 0x0
      12'h7DE: dout  = 8'b00000000; // 2014 :   0 - 0x0
      12'h7DF: dout  = 8'b00000000; // 2015 :   0 - 0x0
      12'h7E0: dout  = 8'b00111000; // 2016 :  56 - 0x38 -- Sprite 0xfc
      12'h7E1: dout  = 8'b00111000; // 2017 :  56 - 0x38
      12'h7E2: dout  = 8'b00000000; // 2018 :   0 - 0x0
      12'h7E3: dout  = 8'b01111100; // 2019 : 124 - 0x7c
      12'h7E4: dout  = 8'b00000000; // 2020 :   0 - 0x0
      12'h7E5: dout  = 8'b00111000; // 2021 :  56 - 0x38
      12'h7E6: dout  = 8'b00111000; // 2022 :  56 - 0x38
      12'h7E7: dout  = 8'b01111100; // 2023 : 124 - 0x7c
      12'h7E8: dout  = 8'b01111100; // 2024 : 124 - 0x7c -- Sprite 0xfd
      12'h7E9: dout  = 8'b01111100; // 2025 : 124 - 0x7c
      12'h7EA: dout  = 8'b01111100; // 2026 : 124 - 0x7c
      12'h7EB: dout  = 8'b00111000; // 2027 :  56 - 0x38
      12'h7EC: dout  = 8'b00000000; // 2028 :   0 - 0x0
      12'h7ED: dout  = 8'b01111100; // 2029 : 124 - 0x7c
      12'h7EE: dout  = 8'b01111100; // 2030 : 124 - 0x7c
      12'h7EF: dout  = 8'b00000000; // 2031 :   0 - 0x0
      12'h7F0: dout  = 8'b00000000; // 2032 :   0 - 0x0 -- Sprite 0xfe
      12'h7F1: dout  = 8'b00000000; // 2033 :   0 - 0x0
      12'h7F2: dout  = 8'b00010001; // 2034 :  17 - 0x11
      12'h7F3: dout  = 8'b11010111; // 2035 : 215 - 0xd7
      12'h7F4: dout  = 8'b11010111; // 2036 : 215 - 0xd7
      12'h7F5: dout  = 8'b11010111; // 2037 : 215 - 0xd7
      12'h7F6: dout  = 8'b00010001; // 2038 :  17 - 0x11
      12'h7F7: dout  = 8'b00000000; // 2039 :   0 - 0x0
      12'h7F8: dout  = 8'b00000000; // 2040 :   0 - 0x0 -- Sprite 0xff
      12'h7F9: dout  = 8'b00000000; // 2041 :   0 - 0x0
      12'h7FA: dout  = 8'b11100110; // 2042 : 230 - 0xe6
      12'h7FB: dout  = 8'b11110110; // 2043 : 246 - 0xf6
      12'h7FC: dout  = 8'b11110110; // 2044 : 246 - 0xf6
      12'h7FD: dout  = 8'b11110110; // 2045 : 246 - 0xf6
      12'h7FE: dout  = 8'b11100110; // 2046 : 230 - 0xe6
      12'h7FF: dout  = 8'b00000000; // 2047 :   0 - 0x0
          // Background pattern Table
      12'h800: dout  = 8'b00000000; // 2048 :   0 - 0x0 -- Background 0x0
      12'h801: dout  = 8'b01111111; // 2049 : 127 - 0x7f
      12'h802: dout  = 8'b01111111; // 2050 : 127 - 0x7f
      12'h803: dout  = 8'b01111111; // 2051 : 127 - 0x7f
      12'h804: dout  = 8'b01111111; // 2052 : 127 - 0x7f
      12'h805: dout  = 8'b01111111; // 2053 : 127 - 0x7f
      12'h806: dout  = 8'b01101010; // 2054 : 106 - 0x6a
      12'h807: dout  = 8'b00000000; // 2055 :   0 - 0x0
      12'h808: dout  = 8'b00000000; // 2056 :   0 - 0x0 -- Background 0x1
      12'h809: dout  = 8'b01111011; // 2057 : 123 - 0x7b
      12'h80A: dout  = 8'b01110011; // 2058 : 115 - 0x73
      12'h80B: dout  = 8'b01111011; // 2059 : 123 - 0x7b
      12'h80C: dout  = 8'b01110011; // 2060 : 115 - 0x73
      12'h80D: dout  = 8'b01111011; // 2061 : 123 - 0x7b
      12'h80E: dout  = 8'b01010011; // 2062 :  83 - 0x53
      12'h80F: dout  = 8'b00000000; // 2063 :   0 - 0x0
      12'h810: dout  = 8'b00000000; // 2064 :   0 - 0x0 -- Background 0x2
      12'h811: dout  = 8'b11011110; // 2065 : 222 - 0xde
      12'h812: dout  = 8'b10011110; // 2066 : 158 - 0x9e
      12'h813: dout  = 8'b11011100; // 2067 : 220 - 0xdc
      12'h814: dout  = 8'b10011110; // 2068 : 158 - 0x9e
      12'h815: dout  = 8'b11011100; // 2069 : 220 - 0xdc
      12'h816: dout  = 8'b10011010; // 2070 : 154 - 0x9a
      12'h817: dout  = 8'b00000000; // 2071 :   0 - 0x0
      12'h818: dout  = 8'b00000000; // 2072 :   0 - 0x0 -- Background 0x3
      12'h819: dout  = 8'b11111110; // 2073 : 254 - 0xfe
      12'h81A: dout  = 8'b11111100; // 2074 : 252 - 0xfc
      12'h81B: dout  = 8'b11111110; // 2075 : 254 - 0xfe
      12'h81C: dout  = 8'b11111100; // 2076 : 252 - 0xfc
      12'h81D: dout  = 8'b11111110; // 2077 : 254 - 0xfe
      12'h81E: dout  = 8'b01010100; // 2078 :  84 - 0x54
      12'h81F: dout  = 8'b00000000; // 2079 :   0 - 0x0
      12'h820: dout  = 8'b00000000; // 2080 :   0 - 0x0 -- Background 0x4
      12'h821: dout  = 8'b01111111; // 2081 : 127 - 0x7f
      12'h822: dout  = 8'b01011111; // 2082 :  95 - 0x5f
      12'h823: dout  = 8'b01111001; // 2083 : 121 - 0x79
      12'h824: dout  = 8'b01111001; // 2084 : 121 - 0x79
      12'h825: dout  = 8'b01001001; // 2085 :  73 - 0x49
      12'h826: dout  = 8'b01001111; // 2086 :  79 - 0x4f
      12'h827: dout  = 8'b01001110; // 2087 :  78 - 0x4e
      12'h828: dout  = 8'b01111000; // 2088 : 120 - 0x78 -- Background 0x5
      12'h829: dout  = 8'b01110000; // 2089 : 112 - 0x70
      12'h82A: dout  = 8'b01100000; // 2090 :  96 - 0x60
      12'h82B: dout  = 8'b01100000; // 2091 :  96 - 0x60
      12'h82C: dout  = 8'b01110001; // 2092 : 113 - 0x71
      12'h82D: dout  = 8'b01011111; // 2093 :  95 - 0x5f
      12'h82E: dout  = 8'b01111111; // 2094 : 127 - 0x7f
      12'h82F: dout  = 8'b00000000; // 2095 :   0 - 0x0
      12'h830: dout  = 8'b00000000; // 2096 :   0 - 0x0 -- Background 0x6
      12'h831: dout  = 8'b11111110; // 2097 : 254 - 0xfe
      12'h832: dout  = 8'b11111010; // 2098 : 250 - 0xfa
      12'h833: dout  = 8'b10011110; // 2099 : 158 - 0x9e
      12'h834: dout  = 8'b10011110; // 2100 : 158 - 0x9e
      12'h835: dout  = 8'b10010010; // 2101 : 146 - 0x92
      12'h836: dout  = 8'b11110010; // 2102 : 242 - 0xf2
      12'h837: dout  = 8'b01110010; // 2103 : 114 - 0x72
      12'h838: dout  = 8'b00011110; // 2104 :  30 - 0x1e -- Background 0x7
      12'h839: dout  = 8'b00001110; // 2105 :  14 - 0xe
      12'h83A: dout  = 8'b00000110; // 2106 :   6 - 0x6
      12'h83B: dout  = 8'b00000110; // 2107 :   6 - 0x6
      12'h83C: dout  = 8'b10001110; // 2108 : 142 - 0x8e
      12'h83D: dout  = 8'b11111010; // 2109 : 250 - 0xfa
      12'h83E: dout  = 8'b11111110; // 2110 : 254 - 0xfe
      12'h83F: dout  = 8'b00000000; // 2111 :   0 - 0x0
      12'h840: dout  = 8'b00000000; // 2112 :   0 - 0x0 -- Background 0x8
      12'h841: dout  = 8'b01111111; // 2113 : 127 - 0x7f
      12'h842: dout  = 8'b01011111; // 2114 :  95 - 0x5f
      12'h843: dout  = 8'b01111111; // 2115 : 127 - 0x7f
      12'h844: dout  = 8'b01111111; // 2116 : 127 - 0x7f
      12'h845: dout  = 8'b01111111; // 2117 : 127 - 0x7f
      12'h846: dout  = 8'b01111111; // 2118 : 127 - 0x7f
      12'h847: dout  = 8'b01111111; // 2119 : 127 - 0x7f
      12'h848: dout  = 8'b01111111; // 2120 : 127 - 0x7f -- Background 0x9
      12'h849: dout  = 8'b01111111; // 2121 : 127 - 0x7f
      12'h84A: dout  = 8'b01111111; // 2122 : 127 - 0x7f
      12'h84B: dout  = 8'b01111111; // 2123 : 127 - 0x7f
      12'h84C: dout  = 8'b01111111; // 2124 : 127 - 0x7f
      12'h84D: dout  = 8'b01011111; // 2125 :  95 - 0x5f
      12'h84E: dout  = 8'b01111111; // 2126 : 127 - 0x7f
      12'h84F: dout  = 8'b00000000; // 2127 :   0 - 0x0
      12'h850: dout  = 8'b00000000; // 2128 :   0 - 0x0 -- Background 0xa
      12'h851: dout  = 8'b11111110; // 2129 : 254 - 0xfe
      12'h852: dout  = 8'b11111010; // 2130 : 250 - 0xfa
      12'h853: dout  = 8'b11111110; // 2131 : 254 - 0xfe
      12'h854: dout  = 8'b11111110; // 2132 : 254 - 0xfe
      12'h855: dout  = 8'b11111110; // 2133 : 254 - 0xfe
      12'h856: dout  = 8'b11111110; // 2134 : 254 - 0xfe
      12'h857: dout  = 8'b11111110; // 2135 : 254 - 0xfe
      12'h858: dout  = 8'b11111110; // 2136 : 254 - 0xfe -- Background 0xb
      12'h859: dout  = 8'b11111110; // 2137 : 254 - 0xfe
      12'h85A: dout  = 8'b11111110; // 2138 : 254 - 0xfe
      12'h85B: dout  = 8'b11111110; // 2139 : 254 - 0xfe
      12'h85C: dout  = 8'b11111110; // 2140 : 254 - 0xfe
      12'h85D: dout  = 8'b11111010; // 2141 : 250 - 0xfa
      12'h85E: dout  = 8'b11111110; // 2142 : 254 - 0xfe
      12'h85F: dout  = 8'b00000000; // 2143 :   0 - 0x0
      12'h860: dout  = 8'b00000000; // 2144 :   0 - 0x0 -- Background 0xc
      12'h861: dout  = 8'b00111111; // 2145 :  63 - 0x3f
      12'h862: dout  = 8'b01011111; // 2146 :  95 - 0x5f
      12'h863: dout  = 8'b01101111; // 2147 : 111 - 0x6f
      12'h864: dout  = 8'b01110000; // 2148 : 112 - 0x70
      12'h865: dout  = 8'b01110111; // 2149 : 119 - 0x77
      12'h866: dout  = 8'b01110111; // 2150 : 119 - 0x77
      12'h867: dout  = 8'b01110111; // 2151 : 119 - 0x77
      12'h868: dout  = 8'b01110111; // 2152 : 119 - 0x77 -- Background 0xd
      12'h869: dout  = 8'b01110111; // 2153 : 119 - 0x77
      12'h86A: dout  = 8'b01110111; // 2154 : 119 - 0x77
      12'h86B: dout  = 8'b01110000; // 2155 : 112 - 0x70
      12'h86C: dout  = 8'b01101111; // 2156 : 111 - 0x6f
      12'h86D: dout  = 8'b01011111; // 2157 :  95 - 0x5f
      12'h86E: dout  = 8'b00010101; // 2158 :  21 - 0x15
      12'h86F: dout  = 8'b00000000; // 2159 :   0 - 0x0
      12'h870: dout  = 8'b00000000; // 2160 :   0 - 0x0 -- Background 0xe
      12'h871: dout  = 8'b11111100; // 2161 : 252 - 0xfc
      12'h872: dout  = 8'b11111000; // 2162 : 248 - 0xf8
      12'h873: dout  = 8'b11110110; // 2163 : 246 - 0xf6
      12'h874: dout  = 8'b00001100; // 2164 :  12 - 0xc
      12'h875: dout  = 8'b11101110; // 2165 : 238 - 0xee
      12'h876: dout  = 8'b11101100; // 2166 : 236 - 0xec
      12'h877: dout  = 8'b11101110; // 2167 : 238 - 0xee
      12'h878: dout  = 8'b11101100; // 2168 : 236 - 0xec -- Background 0xf
      12'h879: dout  = 8'b11101110; // 2169 : 238 - 0xee
      12'h87A: dout  = 8'b11101100; // 2170 : 236 - 0xec
      12'h87B: dout  = 8'b00001110; // 2171 :  14 - 0xe
      12'h87C: dout  = 8'b11110100; // 2172 : 244 - 0xf4
      12'h87D: dout  = 8'b11111010; // 2173 : 250 - 0xfa
      12'h87E: dout  = 8'b01010100; // 2174 :  84 - 0x54
      12'h87F: dout  = 8'b00000000; // 2175 :   0 - 0x0
      12'h880: dout  = 8'b01100000; // 2176 :  96 - 0x60 -- Background 0x10
      12'h881: dout  = 8'b01100000; // 2177 :  96 - 0x60
      12'h882: dout  = 8'b01100000; // 2178 :  96 - 0x60
      12'h883: dout  = 8'b01101111; // 2179 : 111 - 0x6f
      12'h884: dout  = 8'b01101010; // 2180 : 106 - 0x6a
      12'h885: dout  = 8'b01100000; // 2181 :  96 - 0x60
      12'h886: dout  = 8'b01100000; // 2182 :  96 - 0x60
      12'h887: dout  = 8'b01100000; // 2183 :  96 - 0x60
      12'h888: dout  = 8'b00000110; // 2184 :   6 - 0x6 -- Background 0x11
      12'h889: dout  = 8'b00000100; // 2185 :   4 - 0x4
      12'h88A: dout  = 8'b00000110; // 2186 :   6 - 0x6
      12'h88B: dout  = 8'b11110100; // 2187 : 244 - 0xf4
      12'h88C: dout  = 8'b10100110; // 2188 : 166 - 0xa6
      12'h88D: dout  = 8'b00000100; // 2189 :   4 - 0x4
      12'h88E: dout  = 8'b00000110; // 2190 :   6 - 0x6
      12'h88F: dout  = 8'b00000100; // 2191 :   4 - 0x4
      12'h890: dout  = 8'b00000000; // 2192 :   0 - 0x0 -- Background 0x12
      12'h891: dout  = 8'b00001000; // 2193 :   8 - 0x8
      12'h892: dout  = 8'b00001000; // 2194 :   8 - 0x8
      12'h893: dout  = 8'b00011100; // 2195 :  28 - 0x1c
      12'h894: dout  = 8'b00011100; // 2196 :  28 - 0x1c
      12'h895: dout  = 8'b00111100; // 2197 :  60 - 0x3c
      12'h896: dout  = 8'b00111100; // 2198 :  60 - 0x3c
      12'h897: dout  = 8'b00111100; // 2199 :  60 - 0x3c
      12'h898: dout  = 8'b00111100; // 2200 :  60 - 0x3c -- Background 0x13
      12'h899: dout  = 8'b01111110; // 2201 : 126 - 0x7e
      12'h89A: dout  = 8'b01111110; // 2202 : 126 - 0x7e
      12'h89B: dout  = 8'b01111110; // 2203 : 126 - 0x7e
      12'h89C: dout  = 8'b01111110; // 2204 : 126 - 0x7e
      12'h89D: dout  = 8'b01111110; // 2205 : 126 - 0x7e
      12'h89E: dout  = 8'b01111110; // 2206 : 126 - 0x7e
      12'h89F: dout  = 8'b00000000; // 2207 :   0 - 0x0
      12'h8A0: dout  = 8'b00000000; // 2208 :   0 - 0x0 -- Background 0x14
      12'h8A1: dout  = 8'b00000000; // 2209 :   0 - 0x0
      12'h8A2: dout  = 8'b00000101; // 2210 :   5 - 0x5
      12'h8A3: dout  = 8'b00000011; // 2211 :   3 - 0x3
      12'h8A4: dout  = 8'b00000000; // 2212 :   0 - 0x0
      12'h8A5: dout  = 8'b00000000; // 2213 :   0 - 0x0
      12'h8A6: dout  = 8'b00000010; // 2214 :   2 - 0x2
      12'h8A7: dout  = 8'b00001111; // 2215 :  15 - 0xf
      12'h8A8: dout  = 8'b00011100; // 2216 :  28 - 0x1c -- Background 0x15
      12'h8A9: dout  = 8'b00111010; // 2217 :  58 - 0x3a
      12'h8AA: dout  = 8'b00111100; // 2218 :  60 - 0x3c
      12'h8AB: dout  = 8'b00111111; // 2219 :  63 - 0x3f
      12'h8AC: dout  = 8'b00111000; // 2220 :  56 - 0x38
      12'h8AD: dout  = 8'b00011110; // 2221 :  30 - 0x1e
      12'h8AE: dout  = 8'b00001111; // 2222 :  15 - 0xf
      12'h8AF: dout  = 8'b00000000; // 2223 :   0 - 0x0
      12'h8B0: dout  = 8'b00000000; // 2224 :   0 - 0x0 -- Background 0x16
      12'h8B1: dout  = 8'b00000000; // 2225 :   0 - 0x0
      12'h8B2: dout  = 8'b01000000; // 2226 :  64 - 0x40
      12'h8B3: dout  = 8'b11000000; // 2227 : 192 - 0xc0
      12'h8B4: dout  = 8'b00000000; // 2228 :   0 - 0x0
      12'h8B5: dout  = 8'b10000000; // 2229 : 128 - 0x80
      12'h8B6: dout  = 8'b11000000; // 2230 : 192 - 0xc0
      12'h8B7: dout  = 8'b01110000; // 2231 : 112 - 0x70
      12'h8B8: dout  = 8'b00011000; // 2232 :  24 - 0x18 -- Background 0x17
      12'h8B9: dout  = 8'b11111100; // 2233 : 252 - 0xfc
      12'h8BA: dout  = 8'b00111100; // 2234 :  60 - 0x3c
      12'h8BB: dout  = 8'b01011100; // 2235 :  92 - 0x5c
      12'h8BC: dout  = 8'b00111100; // 2236 :  60 - 0x3c
      12'h8BD: dout  = 8'b11111000; // 2237 : 248 - 0xf8
      12'h8BE: dout  = 8'b11110000; // 2238 : 240 - 0xf0
      12'h8BF: dout  = 8'b00000000; // 2239 :   0 - 0x0
      12'h8C0: dout  = 8'b00000000; // 2240 :   0 - 0x0 -- Background 0x18
      12'h8C1: dout  = 8'b00111111; // 2241 :  63 - 0x3f
      12'h8C2: dout  = 8'b00111111; // 2242 :  63 - 0x3f
      12'h8C3: dout  = 8'b01111111; // 2243 : 127 - 0x7f
      12'h8C4: dout  = 8'b01111111; // 2244 : 127 - 0x7f
      12'h8C5: dout  = 8'b00000000; // 2245 :   0 - 0x0
      12'h8C6: dout  = 8'b00000000; // 2246 :   0 - 0x0
      12'h8C7: dout  = 8'b00000000; // 2247 :   0 - 0x0
      12'h8C8: dout  = 8'b00000000; // 2248 :   0 - 0x0 -- Background 0x19
      12'h8C9: dout  = 8'b11111100; // 2249 : 252 - 0xfc
      12'h8CA: dout  = 8'b11111100; // 2250 : 252 - 0xfc
      12'h8CB: dout  = 8'b11111110; // 2251 : 254 - 0xfe
      12'h8CC: dout  = 8'b11111110; // 2252 : 254 - 0xfe
      12'h8CD: dout  = 8'b00000000; // 2253 :   0 - 0x0
      12'h8CE: dout  = 8'b00000000; // 2254 :   0 - 0x0
      12'h8CF: dout  = 8'b00000000; // 2255 :   0 - 0x0
      12'h8D0: dout  = 8'b00000000; // 2256 :   0 - 0x0 -- Background 0x1a
      12'h8D1: dout  = 8'b00000000; // 2257 :   0 - 0x0
      12'h8D2: dout  = 8'b00000000; // 2258 :   0 - 0x0
      12'h8D3: dout  = 8'b00111111; // 2259 :  63 - 0x3f
      12'h8D4: dout  = 8'b00111111; // 2260 :  63 - 0x3f
      12'h8D5: dout  = 8'b01111111; // 2261 : 127 - 0x7f
      12'h8D6: dout  = 8'b01111111; // 2262 : 127 - 0x7f
      12'h8D7: dout  = 8'b00000000; // 2263 :   0 - 0x0
      12'h8D8: dout  = 8'b00000000; // 2264 :   0 - 0x0 -- Background 0x1b
      12'h8D9: dout  = 8'b00000000; // 2265 :   0 - 0x0
      12'h8DA: dout  = 8'b00000000; // 2266 :   0 - 0x0
      12'h8DB: dout  = 8'b11111100; // 2267 : 252 - 0xfc
      12'h8DC: dout  = 8'b11111100; // 2268 : 252 - 0xfc
      12'h8DD: dout  = 8'b11111110; // 2269 : 254 - 0xfe
      12'h8DE: dout  = 8'b11111110; // 2270 : 254 - 0xfe
      12'h8DF: dout  = 8'b00000000; // 2271 :   0 - 0x0
      12'h8E0: dout  = 8'b00000000; // 2272 :   0 - 0x0 -- Background 0x1c
      12'h8E1: dout  = 8'b01111111; // 2273 : 127 - 0x7f
      12'h8E2: dout  = 8'b01111111; // 2274 : 127 - 0x7f
      12'h8E3: dout  = 8'b01111111; // 2275 : 127 - 0x7f
      12'h8E4: dout  = 8'b01100100; // 2276 : 100 - 0x64
      12'h8E5: dout  = 8'b01011011; // 2277 :  91 - 0x5b
      12'h8E6: dout  = 8'b01011001; // 2278 :  89 - 0x59
      12'h8E7: dout  = 8'b01111111; // 2279 : 127 - 0x7f
      12'h8E8: dout  = 8'b01111111; // 2280 : 127 - 0x7f -- Background 0x1d
      12'h8E9: dout  = 8'b00000000; // 2281 :   0 - 0x0
      12'h8EA: dout  = 8'b00000001; // 2282 :   1 - 0x1
      12'h8EB: dout  = 8'b00000001; // 2283 :   1 - 0x1
      12'h8EC: dout  = 8'b00000001; // 2284 :   1 - 0x1
      12'h8ED: dout  = 8'b00000001; // 2285 :   1 - 0x1
      12'h8EE: dout  = 8'b00000001; // 2286 :   1 - 0x1
      12'h8EF: dout  = 8'b00000000; // 2287 :   0 - 0x0
      12'h8F0: dout  = 8'b00000000; // 2288 :   0 - 0x0 -- Background 0x1e
      12'h8F1: dout  = 8'b11111110; // 2289 : 254 - 0xfe
      12'h8F2: dout  = 8'b11111110; // 2290 : 254 - 0xfe
      12'h8F3: dout  = 8'b11111110; // 2291 : 254 - 0xfe
      12'h8F4: dout  = 8'b10111110; // 2292 : 190 - 0xbe
      12'h8F5: dout  = 8'b00001010; // 2293 :  10 - 0xa
      12'h8F6: dout  = 8'b11100010; // 2294 : 226 - 0xe2
      12'h8F7: dout  = 8'b11111110; // 2295 : 254 - 0xfe
      12'h8F8: dout  = 8'b11111110; // 2296 : 254 - 0xfe -- Background 0x1f
      12'h8F9: dout  = 8'b00000000; // 2297 :   0 - 0x0
      12'h8FA: dout  = 8'b10000000; // 2298 : 128 - 0x80
      12'h8FB: dout  = 8'b10000000; // 2299 : 128 - 0x80
      12'h8FC: dout  = 8'b10000000; // 2300 : 128 - 0x80
      12'h8FD: dout  = 8'b10000000; // 2301 : 128 - 0x80
      12'h8FE: dout  = 8'b10000000; // 2302 : 128 - 0x80
      12'h8FF: dout  = 8'b00000000; // 2303 :   0 - 0x0
      12'h900: dout  = 8'b00000000; // 2304 :   0 - 0x0 -- Background 0x20
      12'h901: dout  = 8'b00000000; // 2305 :   0 - 0x0
      12'h902: dout  = 8'b00000000; // 2306 :   0 - 0x0
      12'h903: dout  = 8'b00000000; // 2307 :   0 - 0x0
      12'h904: dout  = 8'b00000000; // 2308 :   0 - 0x0
      12'h905: dout  = 8'b00000000; // 2309 :   0 - 0x0
      12'h906: dout  = 8'b00000000; // 2310 :   0 - 0x0
      12'h907: dout  = 8'b00000000; // 2311 :   0 - 0x0
      12'h908: dout  = 8'b00000000; // 2312 :   0 - 0x0 -- Background 0x21
      12'h909: dout  = 8'b00000000; // 2313 :   0 - 0x0
      12'h90A: dout  = 8'b00000000; // 2314 :   0 - 0x0
      12'h90B: dout  = 8'b00000000; // 2315 :   0 - 0x0
      12'h90C: dout  = 8'b00000000; // 2316 :   0 - 0x0
      12'h90D: dout  = 8'b00000000; // 2317 :   0 - 0x0
      12'h90E: dout  = 8'b00000000; // 2318 :   0 - 0x0
      12'h90F: dout  = 8'b00000000; // 2319 :   0 - 0x0
      12'h910: dout  = 8'b00000000; // 2320 :   0 - 0x0 -- Background 0x22
      12'h911: dout  = 8'b00000000; // 2321 :   0 - 0x0
      12'h912: dout  = 8'b00011000; // 2322 :  24 - 0x18
      12'h913: dout  = 8'b00010000; // 2323 :  16 - 0x10
      12'h914: dout  = 8'b00011010; // 2324 :  26 - 0x1a
      12'h915: dout  = 8'b00010001; // 2325 :  17 - 0x11
      12'h916: dout  = 8'b00011010; // 2326 :  26 - 0x1a
      12'h917: dout  = 8'b00000000; // 2327 :   0 - 0x0
      12'h918: dout  = 8'b00000000; // 2328 :   0 - 0x0 -- Background 0x23
      12'h919: dout  = 8'b00000000; // 2329 :   0 - 0x0
      12'h91A: dout  = 8'b00000000; // 2330 :   0 - 0x0
      12'h91B: dout  = 8'b00101000; // 2331 :  40 - 0x28
      12'h91C: dout  = 8'b10001100; // 2332 : 140 - 0x8c
      12'h91D: dout  = 8'b00101000; // 2333 :  40 - 0x28
      12'h91E: dout  = 8'b10101100; // 2334 : 172 - 0xac
      12'h91F: dout  = 8'b00000000; // 2335 :   0 - 0x0
      12'h920: dout  = 8'b00000000; // 2336 :   0 - 0x0 -- Background 0x24
      12'h921: dout  = 8'b00000000; // 2337 :   0 - 0x0
      12'h922: dout  = 8'b00000000; // 2338 :   0 - 0x0
      12'h923: dout  = 8'b00000000; // 2339 :   0 - 0x0
      12'h924: dout  = 8'b00000000; // 2340 :   0 - 0x0
      12'h925: dout  = 8'b00000000; // 2341 :   0 - 0x0
      12'h926: dout  = 8'b00000000; // 2342 :   0 - 0x0
      12'h927: dout  = 8'b00000000; // 2343 :   0 - 0x0
      12'h928: dout  = 8'b00011100; // 2344 :  28 - 0x1c -- Background 0x25
      12'h929: dout  = 8'b00111001; // 2345 :  57 - 0x39
      12'h92A: dout  = 8'b00111111; // 2346 :  63 - 0x3f
      12'h92B: dout  = 8'b00111110; // 2347 :  62 - 0x3e
      12'h92C: dout  = 8'b00111111; // 2348 :  63 - 0x3f
      12'h92D: dout  = 8'b00011110; // 2349 :  30 - 0x1e
      12'h92E: dout  = 8'b00001111; // 2350 :  15 - 0xf
      12'h92F: dout  = 8'b00000000; // 2351 :   0 - 0x0
      12'h930: dout  = 8'b00000000; // 2352 :   0 - 0x0 -- Background 0x26
      12'h931: dout  = 8'b00000000; // 2353 :   0 - 0x0
      12'h932: dout  = 8'b01000000; // 2354 :  64 - 0x40
      12'h933: dout  = 8'b11000000; // 2355 : 192 - 0xc0
      12'h934: dout  = 8'b00000000; // 2356 :   0 - 0x0
      12'h935: dout  = 8'b10000000; // 2357 : 128 - 0x80
      12'h936: dout  = 8'b11000000; // 2358 : 192 - 0xc0
      12'h937: dout  = 8'b11110000; // 2359 : 240 - 0xf0
      12'h938: dout  = 8'b00111000; // 2360 :  56 - 0x38 -- Background 0x27
      12'h939: dout  = 8'b10011100; // 2361 : 156 - 0x9c
      12'h93A: dout  = 8'b10011100; // 2362 : 156 - 0x9c
      12'h93B: dout  = 8'b00111100; // 2363 :  60 - 0x3c
      12'h93C: dout  = 8'b11111100; // 2364 : 252 - 0xfc
      12'h93D: dout  = 8'b01111000; // 2365 : 120 - 0x78
      12'h93E: dout  = 8'b11110000; // 2366 : 240 - 0xf0
      12'h93F: dout  = 8'b00000000; // 2367 :   0 - 0x0
      12'h940: dout  = 8'b00000000; // 2368 :   0 - 0x0 -- Background 0x28
      12'h941: dout  = 8'b00111110; // 2369 :  62 - 0x3e
      12'h942: dout  = 8'b01011101; // 2370 :  93 - 0x5d
      12'h943: dout  = 8'b01101011; // 2371 : 107 - 0x6b
      12'h944: dout  = 8'b01110101; // 2372 : 117 - 0x75
      12'h945: dout  = 8'b01110001; // 2373 : 113 - 0x71
      12'h946: dout  = 8'b01110101; // 2374 : 117 - 0x75
      12'h947: dout  = 8'b01110100; // 2375 : 116 - 0x74
      12'h948: dout  = 8'b01110000; // 2376 : 112 - 0x70 -- Background 0x29
      12'h949: dout  = 8'b01110111; // 2377 : 119 - 0x77
      12'h94A: dout  = 8'b01110111; // 2378 : 119 - 0x77
      12'h94B: dout  = 8'b01110000; // 2379 : 112 - 0x70
      12'h94C: dout  = 8'b01101111; // 2380 : 111 - 0x6f
      12'h94D: dout  = 8'b01011111; // 2381 :  95 - 0x5f
      12'h94E: dout  = 8'b00010101; // 2382 :  21 - 0x15
      12'h94F: dout  = 8'b00000000; // 2383 :   0 - 0x0
      12'h950: dout  = 8'b00000000; // 2384 :   0 - 0x0 -- Background 0x2a
      12'h951: dout  = 8'b01111100; // 2385 : 124 - 0x7c
      12'h952: dout  = 8'b10111000; // 2386 : 184 - 0xb8
      12'h953: dout  = 8'b11010110; // 2387 : 214 - 0xd6
      12'h954: dout  = 8'b10101100; // 2388 : 172 - 0xac
      12'h955: dout  = 8'b10001110; // 2389 : 142 - 0x8e
      12'h956: dout  = 8'b10101100; // 2390 : 172 - 0xac
      12'h957: dout  = 8'b00101110; // 2391 :  46 - 0x2e
      12'h958: dout  = 8'b00001100; // 2392 :  12 - 0xc -- Background 0x2b
      12'h959: dout  = 8'b11101110; // 2393 : 238 - 0xee
      12'h95A: dout  = 8'b11101100; // 2394 : 236 - 0xec
      12'h95B: dout  = 8'b00001110; // 2395 :  14 - 0xe
      12'h95C: dout  = 8'b11110100; // 2396 : 244 - 0xf4
      12'h95D: dout  = 8'b11111010; // 2397 : 250 - 0xfa
      12'h95E: dout  = 8'b01010100; // 2398 :  84 - 0x54
      12'h95F: dout  = 8'b00000000; // 2399 :   0 - 0x0
      12'h960: dout  = 8'b00000000; // 2400 :   0 - 0x0 -- Background 0x2c
      12'h961: dout  = 8'b00000000; // 2401 :   0 - 0x0
      12'h962: dout  = 8'b00000000; // 2402 :   0 - 0x0
      12'h963: dout  = 8'b00000000; // 2403 :   0 - 0x0
      12'h964: dout  = 8'b00000000; // 2404 :   0 - 0x0
      12'h965: dout  = 8'b00000000; // 2405 :   0 - 0x0
      12'h966: dout  = 8'b00000000; // 2406 :   0 - 0x0
      12'h967: dout  = 8'b00000000; // 2407 :   0 - 0x0
      12'h968: dout  = 8'b00011110; // 2408 :  30 - 0x1e -- Background 0x2d
      12'h969: dout  = 8'b00111110; // 2409 :  62 - 0x3e
      12'h96A: dout  = 8'b00111110; // 2410 :  62 - 0x3e
      12'h96B: dout  = 8'b00111110; // 2411 :  62 - 0x3e
      12'h96C: dout  = 8'b00111111; // 2412 :  63 - 0x3f
      12'h96D: dout  = 8'b00011110; // 2413 :  30 - 0x1e
      12'h96E: dout  = 8'b00001111; // 2414 :  15 - 0xf
      12'h96F: dout  = 8'b00000000; // 2415 :   0 - 0x0
      12'h970: dout  = 8'b00000000; // 2416 :   0 - 0x0 -- Background 0x2e
      12'h971: dout  = 8'b00000000; // 2417 :   0 - 0x0
      12'h972: dout  = 8'b00000000; // 2418 :   0 - 0x0
      12'h973: dout  = 8'b00000000; // 2419 :   0 - 0x0
      12'h974: dout  = 8'b00000000; // 2420 :   0 - 0x0
      12'h975: dout  = 8'b00000000; // 2421 :   0 - 0x0
      12'h976: dout  = 8'b00000000; // 2422 :   0 - 0x0
      12'h977: dout  = 8'b00000000; // 2423 :   0 - 0x0
      12'h978: dout  = 8'b01111000; // 2424 : 120 - 0x78 -- Background 0x2f
      12'h979: dout  = 8'b01111100; // 2425 : 124 - 0x7c
      12'h97A: dout  = 8'b01111100; // 2426 : 124 - 0x7c
      12'h97B: dout  = 8'b01111100; // 2427 : 124 - 0x7c
      12'h97C: dout  = 8'b11111100; // 2428 : 252 - 0xfc
      12'h97D: dout  = 8'b01111000; // 2429 : 120 - 0x78
      12'h97E: dout  = 8'b11110000; // 2430 : 240 - 0xf0
      12'h97F: dout  = 8'b00000000; // 2431 :   0 - 0x0
      12'h980: dout  = 8'b00000000; // 2432 :   0 - 0x0 -- Background 0x30
      12'h981: dout  = 8'b00011000; // 2433 :  24 - 0x18
      12'h982: dout  = 8'b00111100; // 2434 :  60 - 0x3c
      12'h983: dout  = 8'b01011010; // 2435 :  90 - 0x5a
      12'h984: dout  = 8'b00011000; // 2436 :  24 - 0x18
      12'h985: dout  = 8'b00011000; // 2437 :  24 - 0x18
      12'h986: dout  = 8'b00011000; // 2438 :  24 - 0x18
      12'h987: dout  = 8'b00000000; // 2439 :   0 - 0x0
      12'h988: dout  = 8'b00000000; // 2440 :   0 - 0x0 -- Background 0x31
      12'h989: dout  = 8'b00011000; // 2441 :  24 - 0x18
      12'h98A: dout  = 8'b00011000; // 2442 :  24 - 0x18
      12'h98B: dout  = 8'b00011000; // 2443 :  24 - 0x18
      12'h98C: dout  = 8'b01011010; // 2444 :  90 - 0x5a
      12'h98D: dout  = 8'b00111100; // 2445 :  60 - 0x3c
      12'h98E: dout  = 8'b00011000; // 2446 :  24 - 0x18
      12'h98F: dout  = 8'b00000000; // 2447 :   0 - 0x0
      12'h990: dout  = 8'b00000001; // 2448 :   1 - 0x1 -- Background 0x32
      12'h991: dout  = 8'b00000001; // 2449 :   1 - 0x1
      12'h992: dout  = 8'b00000000; // 2450 :   0 - 0x0
      12'h993: dout  = 8'b00000001; // 2451 :   1 - 0x1
      12'h994: dout  = 8'b00000001; // 2452 :   1 - 0x1
      12'h995: dout  = 8'b00000001; // 2453 :   1 - 0x1
      12'h996: dout  = 8'b00000000; // 2454 :   0 - 0x0
      12'h997: dout  = 8'b00000001; // 2455 :   1 - 0x1
      12'h998: dout  = 8'b10000000; // 2456 : 128 - 0x80 -- Background 0x33
      12'h999: dout  = 8'b00000000; // 2457 :   0 - 0x0
      12'h99A: dout  = 8'b10000000; // 2458 : 128 - 0x80
      12'h99B: dout  = 8'b10000000; // 2459 : 128 - 0x80
      12'h99C: dout  = 8'b10000000; // 2460 : 128 - 0x80
      12'h99D: dout  = 8'b00000000; // 2461 :   0 - 0x0
      12'h99E: dout  = 8'b10000000; // 2462 : 128 - 0x80
      12'h99F: dout  = 8'b10000000; // 2463 : 128 - 0x80
      12'h9A0: dout  = 8'b00000000; // 2464 :   0 - 0x0 -- Background 0x34
      12'h9A1: dout  = 8'b00000000; // 2465 :   0 - 0x0
      12'h9A2: dout  = 8'b00011000; // 2466 :  24 - 0x18
      12'h9A3: dout  = 8'b00111100; // 2467 :  60 - 0x3c
      12'h9A4: dout  = 8'b00111110; // 2468 :  62 - 0x3e
      12'h9A5: dout  = 8'b01111111; // 2469 : 127 - 0x7f
      12'h9A6: dout  = 8'b01111111; // 2470 : 127 - 0x7f
      12'h9A7: dout  = 8'b01111111; // 2471 : 127 - 0x7f
      12'h9A8: dout  = 8'b00111111; // 2472 :  63 - 0x3f -- Background 0x35
      12'h9A9: dout  = 8'b00111111; // 2473 :  63 - 0x3f
      12'h9AA: dout  = 8'b00011111; // 2474 :  31 - 0x1f
      12'h9AB: dout  = 8'b00001111; // 2475 :  15 - 0xf
      12'h9AC: dout  = 8'b00000111; // 2476 :   7 - 0x7
      12'h9AD: dout  = 8'b00000011; // 2477 :   3 - 0x3
      12'h9AE: dout  = 8'b00000001; // 2478 :   1 - 0x1
      12'h9AF: dout  = 8'b00000000; // 2479 :   0 - 0x0
      12'h9B0: dout  = 8'b00000000; // 2480 :   0 - 0x0 -- Background 0x36
      12'h9B1: dout  = 8'b00000000; // 2481 :   0 - 0x0
      12'h9B2: dout  = 8'b00011000; // 2482 :  24 - 0x18
      12'h9B3: dout  = 8'b00111100; // 2483 :  60 - 0x3c
      12'h9B4: dout  = 8'b01111100; // 2484 : 124 - 0x7c
      12'h9B5: dout  = 8'b11111110; // 2485 : 254 - 0xfe
      12'h9B6: dout  = 8'b11111110; // 2486 : 254 - 0xfe
      12'h9B7: dout  = 8'b11111110; // 2487 : 254 - 0xfe
      12'h9B8: dout  = 8'b11111100; // 2488 : 252 - 0xfc -- Background 0x37
      12'h9B9: dout  = 8'b11111100; // 2489 : 252 - 0xfc
      12'h9BA: dout  = 8'b11111000; // 2490 : 248 - 0xf8
      12'h9BB: dout  = 8'b11110000; // 2491 : 240 - 0xf0
      12'h9BC: dout  = 8'b11100000; // 2492 : 224 - 0xe0
      12'h9BD: dout  = 8'b11000000; // 2493 : 192 - 0xc0
      12'h9BE: dout  = 8'b10000000; // 2494 : 128 - 0x80
      12'h9BF: dout  = 8'b00000000; // 2495 :   0 - 0x0
      12'h9C0: dout  = 8'b00000000; // 2496 :   0 - 0x0 -- Background 0x38
      12'h9C1: dout  = 8'b00000000; // 2497 :   0 - 0x0
      12'h9C2: dout  = 8'b00000110; // 2498 :   6 - 0x6
      12'h9C3: dout  = 8'b00000111; // 2499 :   7 - 0x7
      12'h9C4: dout  = 8'b00000111; // 2500 :   7 - 0x7
      12'h9C5: dout  = 8'b00000011; // 2501 :   3 - 0x3
      12'h9C6: dout  = 8'b00000001; // 2502 :   1 - 0x1
      12'h9C7: dout  = 8'b00000000; // 2503 :   0 - 0x0
      12'h9C8: dout  = 8'b00000000; // 2504 :   0 - 0x0 -- Background 0x39
      12'h9C9: dout  = 8'b00000000; // 2505 :   0 - 0x0
      12'h9CA: dout  = 8'b00000000; // 2506 :   0 - 0x0
      12'h9CB: dout  = 8'b00000000; // 2507 :   0 - 0x0
      12'h9CC: dout  = 8'b00000000; // 2508 :   0 - 0x0
      12'h9CD: dout  = 8'b00000000; // 2509 :   0 - 0x0
      12'h9CE: dout  = 8'b00000000; // 2510 :   0 - 0x0
      12'h9CF: dout  = 8'b00000000; // 2511 :   0 - 0x0
      12'h9D0: dout  = 8'b00000000; // 2512 :   0 - 0x0 -- Background 0x3a
      12'h9D1: dout  = 8'b00000000; // 2513 :   0 - 0x0
      12'h9D2: dout  = 8'b01100000; // 2514 :  96 - 0x60
      12'h9D3: dout  = 8'b11100000; // 2515 : 224 - 0xe0
      12'h9D4: dout  = 8'b11100000; // 2516 : 224 - 0xe0
      12'h9D5: dout  = 8'b11000000; // 2517 : 192 - 0xc0
      12'h9D6: dout  = 8'b10000000; // 2518 : 128 - 0x80
      12'h9D7: dout  = 8'b00000000; // 2519 :   0 - 0x0
      12'h9D8: dout  = 8'b00000000; // 2520 :   0 - 0x0 -- Background 0x3b
      12'h9D9: dout  = 8'b00101010; // 2521 :  42 - 0x2a
      12'h9DA: dout  = 8'b01000000; // 2522 :  64 - 0x40
      12'h9DB: dout  = 8'b00000010; // 2523 :   2 - 0x2
      12'h9DC: dout  = 8'b01000000; // 2524 :  64 - 0x40
      12'h9DD: dout  = 8'b00000010; // 2525 :   2 - 0x2
      12'h9DE: dout  = 8'b01010100; // 2526 :  84 - 0x54
      12'h9DF: dout  = 8'b00000000; // 2527 :   0 - 0x0
      12'h9E0: dout  = 8'b00000000; // 2528 :   0 - 0x0 -- Background 0x3c
      12'h9E1: dout  = 8'b00000000; // 2529 :   0 - 0x0
      12'h9E2: dout  = 8'b00000000; // 2530 :   0 - 0x0
      12'h9E3: dout  = 8'b00000000; // 2531 :   0 - 0x0
      12'h9E4: dout  = 8'b00000000; // 2532 :   0 - 0x0
      12'h9E5: dout  = 8'b00000000; // 2533 :   0 - 0x0
      12'h9E6: dout  = 8'b00000000; // 2534 :   0 - 0x0
      12'h9E7: dout  = 8'b00000000; // 2535 :   0 - 0x0
      12'h9E8: dout  = 8'b11111111; // 2536 : 255 - 0xff -- Background 0x3d
      12'h9E9: dout  = 8'b11111111; // 2537 : 255 - 0xff
      12'h9EA: dout  = 8'b11111111; // 2538 : 255 - 0xff
      12'h9EB: dout  = 8'b11111111; // 2539 : 255 - 0xff
      12'h9EC: dout  = 8'b11111111; // 2540 : 255 - 0xff
      12'h9ED: dout  = 8'b11111111; // 2541 : 255 - 0xff
      12'h9EE: dout  = 8'b11111111; // 2542 : 255 - 0xff
      12'h9EF: dout  = 8'b11111111; // 2543 : 255 - 0xff
      12'h9F0: dout  = 8'b11111111; // 2544 : 255 - 0xff -- Background 0x3e
      12'h9F1: dout  = 8'b11111111; // 2545 : 255 - 0xff
      12'h9F2: dout  = 8'b11111111; // 2546 : 255 - 0xff
      12'h9F3: dout  = 8'b11111111; // 2547 : 255 - 0xff
      12'h9F4: dout  = 8'b11111111; // 2548 : 255 - 0xff
      12'h9F5: dout  = 8'b11111111; // 2549 : 255 - 0xff
      12'h9F6: dout  = 8'b11111111; // 2550 : 255 - 0xff
      12'h9F7: dout  = 8'b11111111; // 2551 : 255 - 0xff
      12'h9F8: dout  = 8'b00000000; // 2552 :   0 - 0x0 -- Background 0x3f
      12'h9F9: dout  = 8'b00000000; // 2553 :   0 - 0x0
      12'h9FA: dout  = 8'b00000000; // 2554 :   0 - 0x0
      12'h9FB: dout  = 8'b00000000; // 2555 :   0 - 0x0
      12'h9FC: dout  = 8'b00000000; // 2556 :   0 - 0x0
      12'h9FD: dout  = 8'b00000000; // 2557 :   0 - 0x0
      12'h9FE: dout  = 8'b00000000; // 2558 :   0 - 0x0
      12'h9FF: dout  = 8'b00000000; // 2559 :   0 - 0x0
      12'hA00: dout  = 8'b00000000; // 2560 :   0 - 0x0 -- Background 0x40
      12'hA01: dout  = 8'b00000000; // 2561 :   0 - 0x0
      12'hA02: dout  = 8'b00000000; // 2562 :   0 - 0x0
      12'hA03: dout  = 8'b00000000; // 2563 :   0 - 0x0
      12'hA04: dout  = 8'b00000000; // 2564 :   0 - 0x0
      12'hA05: dout  = 8'b00000000; // 2565 :   0 - 0x0
      12'hA06: dout  = 8'b00000000; // 2566 :   0 - 0x0
      12'hA07: dout  = 8'b00000000; // 2567 :   0 - 0x0
      12'hA08: dout  = 8'b00000000; // 2568 :   0 - 0x0 -- Background 0x41
      12'hA09: dout  = 8'b00000000; // 2569 :   0 - 0x0
      12'hA0A: dout  = 8'b00000000; // 2570 :   0 - 0x0
      12'hA0B: dout  = 8'b00000000; // 2571 :   0 - 0x0
      12'hA0C: dout  = 8'b00000000; // 2572 :   0 - 0x0
      12'hA0D: dout  = 8'b00000000; // 2573 :   0 - 0x0
      12'hA0E: dout  = 8'b00000000; // 2574 :   0 - 0x0
      12'hA0F: dout  = 8'b00000000; // 2575 :   0 - 0x0
      12'hA10: dout  = 8'b00000000; // 2576 :   0 - 0x0 -- Background 0x42
      12'hA11: dout  = 8'b00000000; // 2577 :   0 - 0x0
      12'hA12: dout  = 8'b00000000; // 2578 :   0 - 0x0
      12'hA13: dout  = 8'b00000000; // 2579 :   0 - 0x0
      12'hA14: dout  = 8'b00000000; // 2580 :   0 - 0x0
      12'hA15: dout  = 8'b00000000; // 2581 :   0 - 0x0
      12'hA16: dout  = 8'b00000000; // 2582 :   0 - 0x0
      12'hA17: dout  = 8'b00000000; // 2583 :   0 - 0x0
      12'hA18: dout  = 8'b00000000; // 2584 :   0 - 0x0 -- Background 0x43
      12'hA19: dout  = 8'b00000000; // 2585 :   0 - 0x0
      12'hA1A: dout  = 8'b00000000; // 2586 :   0 - 0x0
      12'hA1B: dout  = 8'b00000000; // 2587 :   0 - 0x0
      12'hA1C: dout  = 8'b00000000; // 2588 :   0 - 0x0
      12'hA1D: dout  = 8'b00000000; // 2589 :   0 - 0x0
      12'hA1E: dout  = 8'b00000000; // 2590 :   0 - 0x0
      12'hA1F: dout  = 8'b00000000; // 2591 :   0 - 0x0
      12'hA20: dout  = 8'b00000000; // 2592 :   0 - 0x0 -- Background 0x44
      12'hA21: dout  = 8'b00000000; // 2593 :   0 - 0x0
      12'hA22: dout  = 8'b00000000; // 2594 :   0 - 0x0
      12'hA23: dout  = 8'b00000000; // 2595 :   0 - 0x0
      12'hA24: dout  = 8'b00000000; // 2596 :   0 - 0x0
      12'hA25: dout  = 8'b00000000; // 2597 :   0 - 0x0
      12'hA26: dout  = 8'b00000000; // 2598 :   0 - 0x0
      12'hA27: dout  = 8'b00000000; // 2599 :   0 - 0x0
      12'hA28: dout  = 8'b00000000; // 2600 :   0 - 0x0 -- Background 0x45
      12'hA29: dout  = 8'b00000000; // 2601 :   0 - 0x0
      12'hA2A: dout  = 8'b00000000; // 2602 :   0 - 0x0
      12'hA2B: dout  = 8'b00000000; // 2603 :   0 - 0x0
      12'hA2C: dout  = 8'b00000000; // 2604 :   0 - 0x0
      12'hA2D: dout  = 8'b00000000; // 2605 :   0 - 0x0
      12'hA2E: dout  = 8'b00000000; // 2606 :   0 - 0x0
      12'hA2F: dout  = 8'b00000000; // 2607 :   0 - 0x0
      12'hA30: dout  = 8'b00000000; // 2608 :   0 - 0x0 -- Background 0x46
      12'hA31: dout  = 8'b00000000; // 2609 :   0 - 0x0
      12'hA32: dout  = 8'b00000000; // 2610 :   0 - 0x0
      12'hA33: dout  = 8'b00000000; // 2611 :   0 - 0x0
      12'hA34: dout  = 8'b00000000; // 2612 :   0 - 0x0
      12'hA35: dout  = 8'b00000000; // 2613 :   0 - 0x0
      12'hA36: dout  = 8'b00000000; // 2614 :   0 - 0x0
      12'hA37: dout  = 8'b00000000; // 2615 :   0 - 0x0
      12'hA38: dout  = 8'b00000000; // 2616 :   0 - 0x0 -- Background 0x47
      12'hA39: dout  = 8'b00000000; // 2617 :   0 - 0x0
      12'hA3A: dout  = 8'b00000000; // 2618 :   0 - 0x0
      12'hA3B: dout  = 8'b00000000; // 2619 :   0 - 0x0
      12'hA3C: dout  = 8'b00000000; // 2620 :   0 - 0x0
      12'hA3D: dout  = 8'b00000000; // 2621 :   0 - 0x0
      12'hA3E: dout  = 8'b00000000; // 2622 :   0 - 0x0
      12'hA3F: dout  = 8'b00000000; // 2623 :   0 - 0x0
      12'hA40: dout  = 8'b00000000; // 2624 :   0 - 0x0 -- Background 0x48
      12'hA41: dout  = 8'b00000000; // 2625 :   0 - 0x0
      12'hA42: dout  = 8'b00000000; // 2626 :   0 - 0x0
      12'hA43: dout  = 8'b00000000; // 2627 :   0 - 0x0
      12'hA44: dout  = 8'b00000000; // 2628 :   0 - 0x0
      12'hA45: dout  = 8'b00000000; // 2629 :   0 - 0x0
      12'hA46: dout  = 8'b00000000; // 2630 :   0 - 0x0
      12'hA47: dout  = 8'b00000000; // 2631 :   0 - 0x0
      12'hA48: dout  = 8'b00000000; // 2632 :   0 - 0x0 -- Background 0x49
      12'hA49: dout  = 8'b00000000; // 2633 :   0 - 0x0
      12'hA4A: dout  = 8'b00000000; // 2634 :   0 - 0x0
      12'hA4B: dout  = 8'b00000000; // 2635 :   0 - 0x0
      12'hA4C: dout  = 8'b00000000; // 2636 :   0 - 0x0
      12'hA4D: dout  = 8'b00000000; // 2637 :   0 - 0x0
      12'hA4E: dout  = 8'b00000000; // 2638 :   0 - 0x0
      12'hA4F: dout  = 8'b00000000; // 2639 :   0 - 0x0
      12'hA50: dout  = 8'b00000000; // 2640 :   0 - 0x0 -- Background 0x4a
      12'hA51: dout  = 8'b00000000; // 2641 :   0 - 0x0
      12'hA52: dout  = 8'b00000000; // 2642 :   0 - 0x0
      12'hA53: dout  = 8'b00000000; // 2643 :   0 - 0x0
      12'hA54: dout  = 8'b00000000; // 2644 :   0 - 0x0
      12'hA55: dout  = 8'b00000000; // 2645 :   0 - 0x0
      12'hA56: dout  = 8'b00000000; // 2646 :   0 - 0x0
      12'hA57: dout  = 8'b00000000; // 2647 :   0 - 0x0
      12'hA58: dout  = 8'b00000000; // 2648 :   0 - 0x0 -- Background 0x4b
      12'hA59: dout  = 8'b00000000; // 2649 :   0 - 0x0
      12'hA5A: dout  = 8'b00000000; // 2650 :   0 - 0x0
      12'hA5B: dout  = 8'b00000000; // 2651 :   0 - 0x0
      12'hA5C: dout  = 8'b00000000; // 2652 :   0 - 0x0
      12'hA5D: dout  = 8'b00000000; // 2653 :   0 - 0x0
      12'hA5E: dout  = 8'b00000000; // 2654 :   0 - 0x0
      12'hA5F: dout  = 8'b00000000; // 2655 :   0 - 0x0
      12'hA60: dout  = 8'b00000000; // 2656 :   0 - 0x0 -- Background 0x4c
      12'hA61: dout  = 8'b00000000; // 2657 :   0 - 0x0
      12'hA62: dout  = 8'b00000000; // 2658 :   0 - 0x0
      12'hA63: dout  = 8'b00000000; // 2659 :   0 - 0x0
      12'hA64: dout  = 8'b00000000; // 2660 :   0 - 0x0
      12'hA65: dout  = 8'b00000000; // 2661 :   0 - 0x0
      12'hA66: dout  = 8'b00000000; // 2662 :   0 - 0x0
      12'hA67: dout  = 8'b00000000; // 2663 :   0 - 0x0
      12'hA68: dout  = 8'b00000000; // 2664 :   0 - 0x0 -- Background 0x4d
      12'hA69: dout  = 8'b00000000; // 2665 :   0 - 0x0
      12'hA6A: dout  = 8'b00000000; // 2666 :   0 - 0x0
      12'hA6B: dout  = 8'b00000000; // 2667 :   0 - 0x0
      12'hA6C: dout  = 8'b00000000; // 2668 :   0 - 0x0
      12'hA6D: dout  = 8'b00000000; // 2669 :   0 - 0x0
      12'hA6E: dout  = 8'b00000000; // 2670 :   0 - 0x0
      12'hA6F: dout  = 8'b00000000; // 2671 :   0 - 0x0
      12'hA70: dout  = 8'b00000000; // 2672 :   0 - 0x0 -- Background 0x4e
      12'hA71: dout  = 8'b00000000; // 2673 :   0 - 0x0
      12'hA72: dout  = 8'b00000000; // 2674 :   0 - 0x0
      12'hA73: dout  = 8'b00000000; // 2675 :   0 - 0x0
      12'hA74: dout  = 8'b00000000; // 2676 :   0 - 0x0
      12'hA75: dout  = 8'b00000000; // 2677 :   0 - 0x0
      12'hA76: dout  = 8'b00000000; // 2678 :   0 - 0x0
      12'hA77: dout  = 8'b00000000; // 2679 :   0 - 0x0
      12'hA78: dout  = 8'b00000000; // 2680 :   0 - 0x0 -- Background 0x4f
      12'hA79: dout  = 8'b00000000; // 2681 :   0 - 0x0
      12'hA7A: dout  = 8'b00000000; // 2682 :   0 - 0x0
      12'hA7B: dout  = 8'b00000000; // 2683 :   0 - 0x0
      12'hA7C: dout  = 8'b00000000; // 2684 :   0 - 0x0
      12'hA7D: dout  = 8'b00000000; // 2685 :   0 - 0x0
      12'hA7E: dout  = 8'b00000000; // 2686 :   0 - 0x0
      12'hA7F: dout  = 8'b00000000; // 2687 :   0 - 0x0
      12'hA80: dout  = 8'b00000000; // 2688 :   0 - 0x0 -- Background 0x50
      12'hA81: dout  = 8'b00111111; // 2689 :  63 - 0x3f
      12'hA82: dout  = 8'b01111111; // 2690 : 127 - 0x7f
      12'hA83: dout  = 8'b01111111; // 2691 : 127 - 0x7f
      12'hA84: dout  = 8'b01111111; // 2692 : 127 - 0x7f
      12'hA85: dout  = 8'b00111100; // 2693 :  60 - 0x3c
      12'hA86: dout  = 8'b00000000; // 2694 :   0 - 0x0
      12'hA87: dout  = 8'b01000000; // 2695 :  64 - 0x40
      12'hA88: dout  = 8'b00000000; // 2696 :   0 - 0x0 -- Background 0x51
      12'hA89: dout  = 8'b11111100; // 2697 : 252 - 0xfc
      12'hA8A: dout  = 8'b11111110; // 2698 : 254 - 0xfe
      12'hA8B: dout  = 8'b11111110; // 2699 : 254 - 0xfe
      12'hA8C: dout  = 8'b11111110; // 2700 : 254 - 0xfe
      12'hA8D: dout  = 8'b00111100; // 2701 :  60 - 0x3c
      12'hA8E: dout  = 8'b00000000; // 2702 :   0 - 0x0
      12'hA8F: dout  = 8'b00000010; // 2703 :   2 - 0x2
      12'hA90: dout  = 8'b00000000; // 2704 :   0 - 0x0 -- Background 0x52
      12'hA91: dout  = 8'b00000000; // 2705 :   0 - 0x0
      12'hA92: dout  = 8'b00000011; // 2706 :   3 - 0x3
      12'hA93: dout  = 8'b00000111; // 2707 :   7 - 0x7
      12'hA94: dout  = 8'b00001111; // 2708 :  15 - 0xf
      12'hA95: dout  = 8'b00011111; // 2709 :  31 - 0x1f
      12'hA96: dout  = 8'b00111111; // 2710 :  63 - 0x3f
      12'hA97: dout  = 8'b00110000; // 2711 :  48 - 0x30
      12'hA98: dout  = 8'b00000000; // 2712 :   0 - 0x0 -- Background 0x53
      12'hA99: dout  = 8'b00000000; // 2713 :   0 - 0x0
      12'hA9A: dout  = 8'b10100000; // 2714 : 160 - 0xa0
      12'hA9B: dout  = 8'b10110000; // 2715 : 176 - 0xb0
      12'hA9C: dout  = 8'b10110000; // 2716 : 176 - 0xb0
      12'hA9D: dout  = 8'b10111000; // 2717 : 184 - 0xb8
      12'hA9E: dout  = 8'b01111100; // 2718 : 124 - 0x7c
      12'hA9F: dout  = 8'b01111100; // 2719 : 124 - 0x7c
      12'hAA0: dout  = 8'b00000000; // 2720 :   0 - 0x0 -- Background 0x54
      12'hAA1: dout  = 8'b00100001; // 2721 :  33 - 0x21
      12'hAA2: dout  = 8'b01110001; // 2722 : 113 - 0x71
      12'hAA3: dout  = 8'b00111010; // 2723 :  58 - 0x3a
      12'hAA4: dout  = 8'b01101101; // 2724 : 109 - 0x6d
      12'hAA5: dout  = 8'b00111000; // 2725 :  56 - 0x38
      12'hAA6: dout  = 8'b00011101; // 2726 :  29 - 0x1d
      12'hAA7: dout  = 8'b00101111; // 2727 :  47 - 0x2f
      12'hAA8: dout  = 8'b00000000; // 2728 :   0 - 0x0 -- Background 0x55
      12'hAA9: dout  = 8'b00100001; // 2729 :  33 - 0x21
      12'hAAA: dout  = 8'b01110001; // 2730 : 113 - 0x71
      12'hAAB: dout  = 8'b00111010; // 2731 :  58 - 0x3a
      12'hAAC: dout  = 8'b01101101; // 2732 : 109 - 0x6d
      12'hAAD: dout  = 8'b10111000; // 2733 : 184 - 0xb8
      12'hAAE: dout  = 8'b00011101; // 2734 :  29 - 0x1d
      12'hAAF: dout  = 8'b10101111; // 2735 : 175 - 0xaf
      12'hAB0: dout  = 8'b00000000; // 2736 :   0 - 0x0 -- Background 0x56
      12'hAB1: dout  = 8'b00100000; // 2737 :  32 - 0x20
      12'hAB2: dout  = 8'b01110000; // 2738 : 112 - 0x70
      12'hAB3: dout  = 8'b00111010; // 2739 :  58 - 0x3a
      12'hAB4: dout  = 8'b01101100; // 2740 : 108 - 0x6c
      12'hAB5: dout  = 8'b10111000; // 2741 : 184 - 0xb8
      12'hAB6: dout  = 8'b00011100; // 2742 :  28 - 0x1c
      12'hAB7: dout  = 8'b10101110; // 2743 : 174 - 0xae
      12'hAB8: dout  = 8'b00000000; // 2744 :   0 - 0x0 -- Background 0x57
      12'hAB9: dout  = 8'b01111111; // 2745 : 127 - 0x7f
      12'hABA: dout  = 8'b01001100; // 2746 :  76 - 0x4c
      12'hABB: dout  = 8'b00110011; // 2747 :  51 - 0x33
      12'hABC: dout  = 8'b00000000; // 2748 :   0 - 0x0
      12'hABD: dout  = 8'b00000000; // 2749 :   0 - 0x0
      12'hABE: dout  = 8'b00000000; // 2750 :   0 - 0x0
      12'hABF: dout  = 8'b00000000; // 2751 :   0 - 0x0
      12'hAC0: dout  = 8'b00000000; // 2752 :   0 - 0x0 -- Background 0x58
      12'hAC1: dout  = 8'b11111111; // 2753 : 255 - 0xff
      12'hAC2: dout  = 8'b11001100; // 2754 : 204 - 0xcc
      12'hAC3: dout  = 8'b00110011; // 2755 :  51 - 0x33
      12'hAC4: dout  = 8'b11001100; // 2756 : 204 - 0xcc
      12'hAC5: dout  = 8'b00000000; // 2757 :   0 - 0x0
      12'hAC6: dout  = 8'b00000000; // 2758 :   0 - 0x0
      12'hAC7: dout  = 8'b00000000; // 2759 :   0 - 0x0
      12'hAC8: dout  = 8'b00000000; // 2760 :   0 - 0x0 -- Background 0x59
      12'hAC9: dout  = 8'b11111110; // 2761 : 254 - 0xfe
      12'hACA: dout  = 8'b11001100; // 2762 : 204 - 0xcc
      12'hACB: dout  = 8'b00110000; // 2763 :  48 - 0x30
      12'hACC: dout  = 8'b11000000; // 2764 : 192 - 0xc0
      12'hACD: dout  = 8'b00000000; // 2765 :   0 - 0x0
      12'hACE: dout  = 8'b00000000; // 2766 :   0 - 0x0
      12'hACF: dout  = 8'b00000000; // 2767 :   0 - 0x0
      12'hAD0: dout  = 8'b00000000; // 2768 :   0 - 0x0 -- Background 0x5a
      12'hAD1: dout  = 8'b00000000; // 2769 :   0 - 0x0
      12'hAD2: dout  = 8'b00000000; // 2770 :   0 - 0x0
      12'hAD3: dout  = 8'b00000000; // 2771 :   0 - 0x0
      12'hAD4: dout  = 8'b00000000; // 2772 :   0 - 0x0
      12'hAD5: dout  = 8'b00000000; // 2773 :   0 - 0x0
      12'hAD6: dout  = 8'b00000000; // 2774 :   0 - 0x0
      12'hAD7: dout  = 8'b00000000; // 2775 :   0 - 0x0
      12'hAD8: dout  = 8'b00000000; // 2776 :   0 - 0x0 -- Background 0x5b
      12'hAD9: dout  = 8'b00000000; // 2777 :   0 - 0x0
      12'hADA: dout  = 8'b00000000; // 2778 :   0 - 0x0
      12'hADB: dout  = 8'b00000000; // 2779 :   0 - 0x0
      12'hADC: dout  = 8'b00000001; // 2780 :   1 - 0x1
      12'hADD: dout  = 8'b00000001; // 2781 :   1 - 0x1
      12'hADE: dout  = 8'b00000011; // 2782 :   3 - 0x3
      12'hADF: dout  = 8'b00000011; // 2783 :   3 - 0x3
      12'hAE0: dout  = 8'b00000000; // 2784 :   0 - 0x0 -- Background 0x5c
      12'hAE1: dout  = 8'b00000000; // 2785 :   0 - 0x0
      12'hAE2: dout  = 8'b00000001; // 2786 :   1 - 0x1
      12'hAE3: dout  = 8'b01111110; // 2787 : 126 - 0x7e
      12'hAE4: dout  = 8'b11111111; // 2788 : 255 - 0xff
      12'hAE5: dout  = 8'b11111111; // 2789 : 255 - 0xff
      12'hAE6: dout  = 8'b11111111; // 2790 : 255 - 0xff
      12'hAE7: dout  = 8'b11111111; // 2791 : 255 - 0xff
      12'hAE8: dout  = 8'b00000000; // 2792 :   0 - 0x0 -- Background 0x5d
      12'hAE9: dout  = 8'b11111111; // 2793 : 255 - 0xff
      12'hAEA: dout  = 8'b11111111; // 2794 : 255 - 0xff
      12'hAEB: dout  = 8'b11111111; // 2795 : 255 - 0xff
      12'hAEC: dout  = 8'b01111111; // 2796 : 127 - 0x7f
      12'hAED: dout  = 8'b11111111; // 2797 : 255 - 0xff
      12'hAEE: dout  = 8'b11111111; // 2798 : 255 - 0xff
      12'hAEF: dout  = 8'b11111111; // 2799 : 255 - 0xff
      12'hAF0: dout  = 8'b00000000; // 2800 :   0 - 0x0 -- Background 0x5e
      12'hAF1: dout  = 8'b00000000; // 2801 :   0 - 0x0
      12'hAF2: dout  = 8'b10000000; // 2802 : 128 - 0x80
      12'hAF3: dout  = 8'b01111110; // 2803 : 126 - 0x7e
      12'hAF4: dout  = 8'b10111111; // 2804 : 191 - 0xbf
      12'hAF5: dout  = 8'b11111111; // 2805 : 255 - 0xff
      12'hAF6: dout  = 8'b11111111; // 2806 : 255 - 0xff
      12'hAF7: dout  = 8'b11111111; // 2807 : 255 - 0xff
      12'hAF8: dout  = 8'b00000000; // 2808 :   0 - 0x0 -- Background 0x5f
      12'hAF9: dout  = 8'b00000000; // 2809 :   0 - 0x0
      12'hAFA: dout  = 8'b00000000; // 2810 :   0 - 0x0
      12'hAFB: dout  = 8'b00000000; // 2811 :   0 - 0x0
      12'hAFC: dout  = 8'b10000000; // 2812 : 128 - 0x80
      12'hAFD: dout  = 8'b10000000; // 2813 : 128 - 0x80
      12'hAFE: dout  = 8'b11000000; // 2814 : 192 - 0xc0
      12'hAFF: dout  = 8'b11000000; // 2815 : 192 - 0xc0
      12'hB00: dout  = 8'b01111111; // 2816 : 127 - 0x7f -- Background 0x60
      12'hB01: dout  = 8'b01111111; // 2817 : 127 - 0x7f
      12'hB02: dout  = 8'b01111101; // 2818 : 125 - 0x7d
      12'hB03: dout  = 8'b01111111; // 2819 : 127 - 0x7f
      12'hB04: dout  = 8'b00111111; // 2820 :  63 - 0x3f
      12'hB05: dout  = 8'b01111111; // 2821 : 127 - 0x7f
      12'hB06: dout  = 8'b01111111; // 2822 : 127 - 0x7f
      12'hB07: dout  = 8'b01110111; // 2823 : 119 - 0x77
      12'hB08: dout  = 8'b11111110; // 2824 : 254 - 0xfe -- Background 0x61
      12'hB09: dout  = 8'b11111110; // 2825 : 254 - 0xfe
      12'hB0A: dout  = 8'b11111100; // 2826 : 252 - 0xfc
      12'hB0B: dout  = 8'b11111110; // 2827 : 254 - 0xfe
      12'hB0C: dout  = 8'b10111110; // 2828 : 190 - 0xbe
      12'hB0D: dout  = 8'b11111110; // 2829 : 254 - 0xfe
      12'hB0E: dout  = 8'b11111110; // 2830 : 254 - 0xfe
      12'hB0F: dout  = 8'b11110110; // 2831 : 246 - 0xf6
      12'hB10: dout  = 8'b00000111; // 2832 :   7 - 0x7 -- Background 0x62
      12'hB11: dout  = 8'b00011111; // 2833 :  31 - 0x1f
      12'hB12: dout  = 8'b00111111; // 2834 :  63 - 0x3f
      12'hB13: dout  = 8'b00111111; // 2835 :  63 - 0x3f
      12'hB14: dout  = 8'b00111111; // 2836 :  63 - 0x3f
      12'hB15: dout  = 8'b00011111; // 2837 :  31 - 0x1f
      12'hB16: dout  = 8'b00001111; // 2838 :  15 - 0xf
      12'hB17: dout  = 8'b00000000; // 2839 :   0 - 0x0
      12'hB18: dout  = 8'b01111110; // 2840 : 126 - 0x7e -- Background 0x63
      12'hB19: dout  = 8'b01111100; // 2841 : 124 - 0x7c
      12'hB1A: dout  = 8'b00111110; // 2842 :  62 - 0x3e
      12'hB1B: dout  = 8'b10111100; // 2843 : 188 - 0xbc
      12'hB1C: dout  = 8'b10111110; // 2844 : 190 - 0xbe
      12'hB1D: dout  = 8'b10011100; // 2845 : 156 - 0x9c
      12'hB1E: dout  = 8'b11011000; // 2846 : 216 - 0xd8
      12'hB1F: dout  = 8'b00000000; // 2847 :   0 - 0x0
      12'hB20: dout  = 8'b01000110; // 2848 :  70 - 0x46 -- Background 0x64
      12'hB21: dout  = 8'b01101011; // 2849 : 107 - 0x6b
      12'hB22: dout  = 8'b01110001; // 2850 : 113 - 0x71
      12'hB23: dout  = 8'b00111010; // 2851 :  58 - 0x3a
      12'hB24: dout  = 8'b01101101; // 2852 : 109 - 0x6d
      12'hB25: dout  = 8'b00111000; // 2853 :  56 - 0x38
      12'hB26: dout  = 8'b00011101; // 2854 :  29 - 0x1d
      12'hB27: dout  = 8'b00101111; // 2855 :  47 - 0x2f
      12'hB28: dout  = 8'b01000110; // 2856 :  70 - 0x46 -- Background 0x65
      12'hB29: dout  = 8'b11101011; // 2857 : 235 - 0xeb
      12'hB2A: dout  = 8'b01110001; // 2858 : 113 - 0x71
      12'hB2B: dout  = 8'b00111010; // 2859 :  58 - 0x3a
      12'hB2C: dout  = 8'b01101101; // 2860 : 109 - 0x6d
      12'hB2D: dout  = 8'b10111000; // 2861 : 184 - 0xb8
      12'hB2E: dout  = 8'b00011101; // 2862 :  29 - 0x1d
      12'hB2F: dout  = 8'b10101111; // 2863 : 175 - 0xaf
      12'hB30: dout  = 8'b01000110; // 2864 :  70 - 0x46 -- Background 0x66
      12'hB31: dout  = 8'b11101010; // 2865 : 234 - 0xea
      12'hB32: dout  = 8'b01110000; // 2866 : 112 - 0x70
      12'hB33: dout  = 8'b00111010; // 2867 :  58 - 0x3a
      12'hB34: dout  = 8'b01101100; // 2868 : 108 - 0x6c
      12'hB35: dout  = 8'b10111000; // 2869 : 184 - 0xb8
      12'hB36: dout  = 8'b00011100; // 2870 :  28 - 0x1c
      12'hB37: dout  = 8'b10101110; // 2871 : 174 - 0xae
      12'hB38: dout  = 8'b00000000; // 2872 :   0 - 0x0 -- Background 0x67
      12'hB39: dout  = 8'b01111111; // 2873 : 127 - 0x7f
      12'hB3A: dout  = 8'b01111111; // 2874 : 127 - 0x7f
      12'hB3B: dout  = 8'b00110011; // 2875 :  51 - 0x33
      12'hB3C: dout  = 8'b00000000; // 2876 :   0 - 0x0
      12'hB3D: dout  = 8'b00000000; // 2877 :   0 - 0x0
      12'hB3E: dout  = 8'b00000000; // 2878 :   0 - 0x0
      12'hB3F: dout  = 8'b00000000; // 2879 :   0 - 0x0
      12'hB40: dout  = 8'b00000000; // 2880 :   0 - 0x0 -- Background 0x68
      12'hB41: dout  = 8'b11111111; // 2881 : 255 - 0xff
      12'hB42: dout  = 8'b11111111; // 2882 : 255 - 0xff
      12'hB43: dout  = 8'b11111111; // 2883 : 255 - 0xff
      12'hB44: dout  = 8'b11001100; // 2884 : 204 - 0xcc
      12'hB45: dout  = 8'b00000000; // 2885 :   0 - 0x0
      12'hB46: dout  = 8'b00000000; // 2886 :   0 - 0x0
      12'hB47: dout  = 8'b00000000; // 2887 :   0 - 0x0
      12'hB48: dout  = 8'b00000000; // 2888 :   0 - 0x0 -- Background 0x69
      12'hB49: dout  = 8'b11111110; // 2889 : 254 - 0xfe
      12'hB4A: dout  = 8'b11111110; // 2890 : 254 - 0xfe
      12'hB4B: dout  = 8'b11110000; // 2891 : 240 - 0xf0
      12'hB4C: dout  = 8'b11000000; // 2892 : 192 - 0xc0
      12'hB4D: dout  = 8'b00000000; // 2893 :   0 - 0x0
      12'hB4E: dout  = 8'b00000000; // 2894 :   0 - 0x0
      12'hB4F: dout  = 8'b00000000; // 2895 :   0 - 0x0
      12'hB50: dout  = 8'b00000000; // 2896 :   0 - 0x0 -- Background 0x6a
      12'hB51: dout  = 8'b00000000; // 2897 :   0 - 0x0
      12'hB52: dout  = 8'b00000000; // 2898 :   0 - 0x0
      12'hB53: dout  = 8'b00000000; // 2899 :   0 - 0x0
      12'hB54: dout  = 8'b00000000; // 2900 :   0 - 0x0
      12'hB55: dout  = 8'b00000000; // 2901 :   0 - 0x0
      12'hB56: dout  = 8'b00000000; // 2902 :   0 - 0x0
      12'hB57: dout  = 8'b00000000; // 2903 :   0 - 0x0
      12'hB58: dout  = 8'b00111101; // 2904 :  61 - 0x3d -- Background 0x6b
      12'hB59: dout  = 8'b01111111; // 2905 : 127 - 0x7f
      12'hB5A: dout  = 8'b01111111; // 2906 : 127 - 0x7f
      12'hB5B: dout  = 8'b01111111; // 2907 : 127 - 0x7f
      12'hB5C: dout  = 8'b00111111; // 2908 :  63 - 0x3f
      12'hB5D: dout  = 8'b00001111; // 2909 :  15 - 0xf
      12'hB5E: dout  = 8'b00000000; // 2910 :   0 - 0x0
      12'hB5F: dout  = 8'b00000000; // 2911 :   0 - 0x0
      12'hB60: dout  = 8'b11111111; // 2912 : 255 - 0xff -- Background 0x6c
      12'hB61: dout  = 8'b11111111; // 2913 : 255 - 0xff
      12'hB62: dout  = 8'b11111111; // 2914 : 255 - 0xff
      12'hB63: dout  = 8'b11111111; // 2915 : 255 - 0xff
      12'hB64: dout  = 8'b11111111; // 2916 : 255 - 0xff
      12'hB65: dout  = 8'b11111111; // 2917 : 255 - 0xff
      12'hB66: dout  = 8'b11111110; // 2918 : 254 - 0xfe
      12'hB67: dout  = 8'b00000000; // 2919 :   0 - 0x0
      12'hB68: dout  = 8'b00000000; // 2920 :   0 - 0x0 -- Background 0x6d
      12'hB69: dout  = 8'b00000000; // 2921 :   0 - 0x0
      12'hB6A: dout  = 8'b00000000; // 2922 :   0 - 0x0
      12'hB6B: dout  = 8'b00000000; // 2923 :   0 - 0x0
      12'hB6C: dout  = 8'b00000000; // 2924 :   0 - 0x0
      12'hB6D: dout  = 8'b00000000; // 2925 :   0 - 0x0
      12'hB6E: dout  = 8'b00000000; // 2926 :   0 - 0x0
      12'hB6F: dout  = 8'b00000000; // 2927 :   0 - 0x0
      12'hB70: dout  = 8'b00000000; // 2928 :   0 - 0x0 -- Background 0x6e
      12'hB71: dout  = 8'b00000000; // 2929 :   0 - 0x0
      12'hB72: dout  = 8'b00000000; // 2930 :   0 - 0x0
      12'hB73: dout  = 8'b00000000; // 2931 :   0 - 0x0
      12'hB74: dout  = 8'b00000000; // 2932 :   0 - 0x0
      12'hB75: dout  = 8'b00000000; // 2933 :   0 - 0x0
      12'hB76: dout  = 8'b00000000; // 2934 :   0 - 0x0
      12'hB77: dout  = 8'b00000000; // 2935 :   0 - 0x0
      12'hB78: dout  = 8'b10111000; // 2936 : 184 - 0xb8 -- Background 0x6f
      12'hB79: dout  = 8'b11111100; // 2937 : 252 - 0xfc
      12'hB7A: dout  = 8'b11111110; // 2938 : 254 - 0xfe
      12'hB7B: dout  = 8'b11111110; // 2939 : 254 - 0xfe
      12'hB7C: dout  = 8'b11111100; // 2940 : 252 - 0xfc
      12'hB7D: dout  = 8'b11110000; // 2941 : 240 - 0xf0
      12'hB7E: dout  = 8'b00000000; // 2942 :   0 - 0x0
      12'hB7F: dout  = 8'b00000000; // 2943 :   0 - 0x0
      12'hB80: dout  = 8'b00000000; // 2944 :   0 - 0x0 -- Background 0x70
      12'hB81: dout  = 8'b00111111; // 2945 :  63 - 0x3f
      12'hB82: dout  = 8'b01111111; // 2946 : 127 - 0x7f
      12'hB83: dout  = 8'b01111111; // 2947 : 127 - 0x7f
      12'hB84: dout  = 8'b00011100; // 2948 :  28 - 0x1c
      12'hB85: dout  = 8'b00000000; // 2949 :   0 - 0x0
      12'hB86: dout  = 8'b00000000; // 2950 :   0 - 0x0
      12'hB87: dout  = 8'b00000000; // 2951 :   0 - 0x0
      12'hB88: dout  = 8'b00000000; // 2952 :   0 - 0x0 -- Background 0x71
      12'hB89: dout  = 8'b11111111; // 2953 : 255 - 0xff
      12'hB8A: dout  = 8'b11111111; // 2954 : 255 - 0xff
      12'hB8B: dout  = 8'b11111111; // 2955 : 255 - 0xff
      12'hB8C: dout  = 8'b11111111; // 2956 : 255 - 0xff
      12'hB8D: dout  = 8'b00111100; // 2957 :  60 - 0x3c
      12'hB8E: dout  = 8'b00000000; // 2958 :   0 - 0x0
      12'hB8F: dout  = 8'b00000000; // 2959 :   0 - 0x0
      12'hB90: dout  = 8'b00000000; // 2960 :   0 - 0x0 -- Background 0x72
      12'hB91: dout  = 8'b11111100; // 2961 : 252 - 0xfc
      12'hB92: dout  = 8'b11111110; // 2962 : 254 - 0xfe
      12'hB93: dout  = 8'b11111110; // 2963 : 254 - 0xfe
      12'hB94: dout  = 8'b00111000; // 2964 :  56 - 0x38
      12'hB95: dout  = 8'b00000000; // 2965 :   0 - 0x0
      12'hB96: dout  = 8'b00000000; // 2966 :   0 - 0x0
      12'hB97: dout  = 8'b00000000; // 2967 :   0 - 0x0
      12'hB98: dout  = 8'b11111111; // 2968 : 255 - 0xff -- Background 0x73
      12'hB99: dout  = 8'b11111111; // 2969 : 255 - 0xff
      12'hB9A: dout  = 8'b11111101; // 2970 : 253 - 0xfd
      12'hB9B: dout  = 8'b11111111; // 2971 : 255 - 0xff
      12'hB9C: dout  = 8'b10111111; // 2972 : 191 - 0xbf
      12'hB9D: dout  = 8'b11111111; // 2973 : 255 - 0xff
      12'hB9E: dout  = 8'b11111111; // 2974 : 255 - 0xff
      12'hB9F: dout  = 8'b11110111; // 2975 : 247 - 0xf7
      12'hBA0: dout  = 8'b01000110; // 2976 :  70 - 0x46 -- Background 0x74
      12'hBA1: dout  = 8'b01101011; // 2977 : 107 - 0x6b
      12'hBA2: dout  = 8'b01110001; // 2978 : 113 - 0x71
      12'hBA3: dout  = 8'b00111010; // 2979 :  58 - 0x3a
      12'hBA4: dout  = 8'b01101101; // 2980 : 109 - 0x6d
      12'hBA5: dout  = 8'b00111000; // 2981 :  56 - 0x38
      12'hBA6: dout  = 8'b00011101; // 2982 :  29 - 0x1d
      12'hBA7: dout  = 8'b00000000; // 2983 :   0 - 0x0
      12'hBA8: dout  = 8'b01000110; // 2984 :  70 - 0x46 -- Background 0x75
      12'hBA9: dout  = 8'b11101011; // 2985 : 235 - 0xeb
      12'hBAA: dout  = 8'b01110001; // 2986 : 113 - 0x71
      12'hBAB: dout  = 8'b00111010; // 2987 :  58 - 0x3a
      12'hBAC: dout  = 8'b01101101; // 2988 : 109 - 0x6d
      12'hBAD: dout  = 8'b10111000; // 2989 : 184 - 0xb8
      12'hBAE: dout  = 8'b00011101; // 2990 :  29 - 0x1d
      12'hBAF: dout  = 8'b00000000; // 2991 :   0 - 0x0
      12'hBB0: dout  = 8'b01000110; // 2992 :  70 - 0x46 -- Background 0x76
      12'hBB1: dout  = 8'b11101010; // 2993 : 234 - 0xea
      12'hBB2: dout  = 8'b01110000; // 2994 : 112 - 0x70
      12'hBB3: dout  = 8'b00111010; // 2995 :  58 - 0x3a
      12'hBB4: dout  = 8'b01101100; // 2996 : 108 - 0x6c
      12'hBB5: dout  = 8'b10111000; // 2997 : 184 - 0xb8
      12'hBB6: dout  = 8'b00011100; // 2998 :  28 - 0x1c
      12'hBB7: dout  = 8'b00000000; // 2999 :   0 - 0x0
      12'hBB8: dout  = 8'b10000001; // 3000 : 129 - 0x81 -- Background 0x77
      12'hBB9: dout  = 8'b11111111; // 3001 : 255 - 0xff
      12'hBBA: dout  = 8'b11111101; // 3002 : 253 - 0xfd
      12'hBBB: dout  = 8'b11111111; // 3003 : 255 - 0xff
      12'hBBC: dout  = 8'b10111111; // 3004 : 191 - 0xbf
      12'hBBD: dout  = 8'b11111111; // 3005 : 255 - 0xff
      12'hBBE: dout  = 8'b11111111; // 3006 : 255 - 0xff
      12'hBBF: dout  = 8'b11110111; // 3007 : 247 - 0xf7
      12'hBC0: dout  = 8'b00000000; // 3008 :   0 - 0x0 -- Background 0x78
      12'hBC1: dout  = 8'b00000000; // 3009 :   0 - 0x0
      12'hBC2: dout  = 8'b00000000; // 3010 :   0 - 0x0
      12'hBC3: dout  = 8'b00000000; // 3011 :   0 - 0x0
      12'hBC4: dout  = 8'b00000000; // 3012 :   0 - 0x0
      12'hBC5: dout  = 8'b00000000; // 3013 :   0 - 0x0
      12'hBC6: dout  = 8'b00000000; // 3014 :   0 - 0x0
      12'hBC7: dout  = 8'b00000000; // 3015 :   0 - 0x0
      12'hBC8: dout  = 8'b00000000; // 3016 :   0 - 0x0 -- Background 0x79
      12'hBC9: dout  = 8'b00000000; // 3017 :   0 - 0x0
      12'hBCA: dout  = 8'b00000000; // 3018 :   0 - 0x0
      12'hBCB: dout  = 8'b00000000; // 3019 :   0 - 0x0
      12'hBCC: dout  = 8'b00000000; // 3020 :   0 - 0x0
      12'hBCD: dout  = 8'b00000000; // 3021 :   0 - 0x0
      12'hBCE: dout  = 8'b00000000; // 3022 :   0 - 0x0
      12'hBCF: dout  = 8'b00000000; // 3023 :   0 - 0x0
      12'hBD0: dout  = 8'b00000000; // 3024 :   0 - 0x0 -- Background 0x7a
      12'hBD1: dout  = 8'b00000000; // 3025 :   0 - 0x0
      12'hBD2: dout  = 8'b00000000; // 3026 :   0 - 0x0
      12'hBD3: dout  = 8'b00000000; // 3027 :   0 - 0x0
      12'hBD4: dout  = 8'b00000000; // 3028 :   0 - 0x0
      12'hBD5: dout  = 8'b00000000; // 3029 :   0 - 0x0
      12'hBD6: dout  = 8'b00000000; // 3030 :   0 - 0x0
      12'hBD7: dout  = 8'b00000000; // 3031 :   0 - 0x0
      12'hBD8: dout  = 8'b00000000; // 3032 :   0 - 0x0 -- Background 0x7b
      12'hBD9: dout  = 8'b00000000; // 3033 :   0 - 0x0
      12'hBDA: dout  = 8'b00000000; // 3034 :   0 - 0x0
      12'hBDB: dout  = 8'b00000000; // 3035 :   0 - 0x0
      12'hBDC: dout  = 8'b00000000; // 3036 :   0 - 0x0
      12'hBDD: dout  = 8'b00000000; // 3037 :   0 - 0x0
      12'hBDE: dout  = 8'b00000000; // 3038 :   0 - 0x0
      12'hBDF: dout  = 8'b00000000; // 3039 :   0 - 0x0
      12'hBE0: dout  = 8'b00000000; // 3040 :   0 - 0x0 -- Background 0x7c
      12'hBE1: dout  = 8'b00100010; // 3041 :  34 - 0x22
      12'hBE2: dout  = 8'b01110111; // 3042 : 119 - 0x77
      12'hBE3: dout  = 8'b11111111; // 3043 : 255 - 0xff
      12'hBE4: dout  = 8'b11111011; // 3044 : 251 - 0xfb
      12'hBE5: dout  = 8'b11110101; // 3045 : 245 - 0xf5
      12'hBE6: dout  = 8'b11101111; // 3046 : 239 - 0xef
      12'hBE7: dout  = 8'b11111111; // 3047 : 255 - 0xff
      12'hBE8: dout  = 8'b00000000; // 3048 :   0 - 0x0 -- Background 0x7d
      12'hBE9: dout  = 8'b01110011; // 3049 : 115 - 0x73
      12'hBEA: dout  = 8'b11111111; // 3050 : 255 - 0xff
      12'hBEB: dout  = 8'b11111111; // 3051 : 255 - 0xff
      12'hBEC: dout  = 8'b11111011; // 3052 : 251 - 0xfb
      12'hBED: dout  = 8'b11111101; // 3053 : 253 - 0xfd
      12'hBEE: dout  = 8'b11101111; // 3054 : 239 - 0xef
      12'hBEF: dout  = 8'b11111111; // 3055 : 255 - 0xff
      12'hBF0: dout  = 8'b11011111; // 3056 : 223 - 0xdf -- Background 0x7e
      12'hBF1: dout  = 8'b10101111; // 3057 : 175 - 0xaf
      12'hBF2: dout  = 8'b01111111; // 3058 : 127 - 0x7f
      12'hBF3: dout  = 8'b11111111; // 3059 : 255 - 0xff
      12'hBF4: dout  = 8'b11111011; // 3060 : 251 - 0xfb
      12'hBF5: dout  = 8'b11110101; // 3061 : 245 - 0xf5
      12'hBF6: dout  = 8'b11101111; // 3062 : 239 - 0xef
      12'hBF7: dout  = 8'b11111111; // 3063 : 255 - 0xff
      12'hBF8: dout  = 8'b00000000; // 3064 :   0 - 0x0 -- Background 0x7f
      12'hBF9: dout  = 8'b10101111; // 3065 : 175 - 0xaf
      12'hBFA: dout  = 8'b01111111; // 3066 : 127 - 0x7f
      12'hBFB: dout  = 8'b11111111; // 3067 : 255 - 0xff
      12'hBFC: dout  = 8'b11111011; // 3068 : 251 - 0xfb
      12'hBFD: dout  = 8'b11110101; // 3069 : 245 - 0xf5
      12'hBFE: dout  = 8'b11101111; // 3070 : 239 - 0xef
      12'hBFF: dout  = 8'b11111111; // 3071 : 255 - 0xff
      12'hC00: dout  = 8'b00000000; // 3072 :   0 - 0x0 -- Background 0x80
      12'hC01: dout  = 8'b01111111; // 3073 : 127 - 0x7f
      12'hC02: dout  = 8'b00110000; // 3074 :  48 - 0x30
      12'hC03: dout  = 8'b00110000; // 3075 :  48 - 0x30
      12'hC04: dout  = 8'b00110000; // 3076 :  48 - 0x30
      12'hC05: dout  = 8'b01111111; // 3077 : 127 - 0x7f
      12'hC06: dout  = 8'b00110000; // 3078 :  48 - 0x30
      12'hC07: dout  = 8'b00110000; // 3079 :  48 - 0x30
      12'hC08: dout  = 8'b00000000; // 3080 :   0 - 0x0 -- Background 0x81
      12'hC09: dout  = 8'b01111111; // 3081 : 127 - 0x7f
      12'hC0A: dout  = 8'b00000000; // 3082 :   0 - 0x0
      12'hC0B: dout  = 8'b01111111; // 3083 : 127 - 0x7f
      12'hC0C: dout  = 8'b01111111; // 3084 : 127 - 0x7f
      12'hC0D: dout  = 8'b00100000; // 3085 :  32 - 0x20
      12'hC0E: dout  = 8'b01000000; // 3086 :  64 - 0x40
      12'hC0F: dout  = 8'b00000000; // 3087 :   0 - 0x0
      12'hC10: dout  = 8'b00000000; // 3088 :   0 - 0x0 -- Background 0x82
      12'hC11: dout  = 8'b11111110; // 3089 : 254 - 0xfe
      12'hC12: dout  = 8'b00001100; // 3090 :  12 - 0xc
      12'hC13: dout  = 8'b00001100; // 3091 :  12 - 0xc
      12'hC14: dout  = 8'b00001100; // 3092 :  12 - 0xc
      12'hC15: dout  = 8'b11111110; // 3093 : 254 - 0xfe
      12'hC16: dout  = 8'b00001100; // 3094 :  12 - 0xc
      12'hC17: dout  = 8'b00001100; // 3095 :  12 - 0xc
      12'hC18: dout  = 8'b00000000; // 3096 :   0 - 0x0 -- Background 0x83
      12'hC19: dout  = 8'b11111111; // 3097 : 255 - 0xff
      12'hC1A: dout  = 8'b00000000; // 3098 :   0 - 0x0
      12'hC1B: dout  = 8'b11111111; // 3099 : 255 - 0xff
      12'hC1C: dout  = 8'b11111111; // 3100 : 255 - 0xff
      12'hC1D: dout  = 8'b00000000; // 3101 :   0 - 0x0
      12'hC1E: dout  = 8'b00000000; // 3102 :   0 - 0x0
      12'hC1F: dout  = 8'b00000000; // 3103 :   0 - 0x0
      12'hC20: dout  = 8'b00000000; // 3104 :   0 - 0x0 -- Background 0x84
      12'hC21: dout  = 8'b11111111; // 3105 : 255 - 0xff
      12'hC22: dout  = 8'b11111111; // 3106 : 255 - 0xff
      12'hC23: dout  = 8'b11111111; // 3107 : 255 - 0xff
      12'hC24: dout  = 8'b11111111; // 3108 : 255 - 0xff
      12'hC25: dout  = 8'b11101111; // 3109 : 239 - 0xef
      12'hC26: dout  = 8'b10111011; // 3110 : 187 - 0xbb
      12'hC27: dout  = 8'b00000000; // 3111 :   0 - 0x0
      12'hC28: dout  = 8'b00000000; // 3112 :   0 - 0x0 -- Background 0x85
      12'hC29: dout  = 8'b11111110; // 3113 : 254 - 0xfe
      12'hC2A: dout  = 8'b00000000; // 3114 :   0 - 0x0
      12'hC2B: dout  = 8'b11111110; // 3115 : 254 - 0xfe
      12'hC2C: dout  = 8'b11111110; // 3116 : 254 - 0xfe
      12'hC2D: dout  = 8'b00001100; // 3117 :  12 - 0xc
      12'hC2E: dout  = 8'b00000010; // 3118 :   2 - 0x2
      12'hC2F: dout  = 8'b00000000; // 3119 :   0 - 0x0
      12'hC30: dout  = 8'b00000000; // 3120 :   0 - 0x0 -- Background 0x86
      12'hC31: dout  = 8'b00000000; // 3121 :   0 - 0x0
      12'hC32: dout  = 8'b00000000; // 3122 :   0 - 0x0
      12'hC33: dout  = 8'b00000000; // 3123 :   0 - 0x0
      12'hC34: dout  = 8'b00000000; // 3124 :   0 - 0x0
      12'hC35: dout  = 8'b00000000; // 3125 :   0 - 0x0
      12'hC36: dout  = 8'b00000000; // 3126 :   0 - 0x0
      12'hC37: dout  = 8'b00000000; // 3127 :   0 - 0x0
      12'hC38: dout  = 8'b00000000; // 3128 :   0 - 0x0 -- Background 0x87
      12'hC39: dout  = 8'b00000000; // 3129 :   0 - 0x0
      12'hC3A: dout  = 8'b00000000; // 3130 :   0 - 0x0
      12'hC3B: dout  = 8'b00000000; // 3131 :   0 - 0x0
      12'hC3C: dout  = 8'b00000000; // 3132 :   0 - 0x0
      12'hC3D: dout  = 8'b00000000; // 3133 :   0 - 0x0
      12'hC3E: dout  = 8'b00000000; // 3134 :   0 - 0x0
      12'hC3F: dout  = 8'b00000000; // 3135 :   0 - 0x0
      12'hC40: dout  = 8'b00000000; // 3136 :   0 - 0x0 -- Background 0x88
      12'hC41: dout  = 8'b00000111; // 3137 :   7 - 0x7
      12'hC42: dout  = 8'b00011111; // 3138 :  31 - 0x1f
      12'hC43: dout  = 8'b00111100; // 3139 :  60 - 0x3c
      12'hC44: dout  = 8'b00110001; // 3140 :  49 - 0x31
      12'hC45: dout  = 8'b01110100; // 3141 : 116 - 0x74
      12'hC46: dout  = 8'b01100101; // 3142 : 101 - 0x65
      12'hC47: dout  = 8'b01101010; // 3143 : 106 - 0x6a
      12'hC48: dout  = 8'b01100100; // 3144 : 100 - 0x64 -- Background 0x89
      12'hC49: dout  = 8'b01101101; // 3145 : 109 - 0x6d
      12'hC4A: dout  = 8'b01110010; // 3146 : 114 - 0x72
      12'hC4B: dout  = 8'b00110000; // 3147 :  48 - 0x30
      12'hC4C: dout  = 8'b00111100; // 3148 :  60 - 0x3c
      12'hC4D: dout  = 8'b00011111; // 3149 :  31 - 0x1f
      12'hC4E: dout  = 8'b00000111; // 3150 :   7 - 0x7
      12'hC4F: dout  = 8'b00000000; // 3151 :   0 - 0x0
      12'hC50: dout  = 8'b00000000; // 3152 :   0 - 0x0 -- Background 0x8a
      12'hC51: dout  = 8'b11100000; // 3153 : 224 - 0xe0
      12'hC52: dout  = 8'b11111000; // 3154 : 248 - 0xf8
      12'hC53: dout  = 8'b00111100; // 3155 :  60 - 0x3c
      12'hC54: dout  = 8'b01001100; // 3156 :  76 - 0x4c
      12'hC55: dout  = 8'b01101110; // 3157 : 110 - 0x6e
      12'hC56: dout  = 8'b00100110; // 3158 :  38 - 0x26
      12'hC57: dout  = 8'b01000110; // 3159 :  70 - 0x46
      12'hC58: dout  = 8'b10010110; // 3160 : 150 - 0x96 -- Background 0x8b
      12'hC59: dout  = 8'b01100110; // 3161 : 102 - 0x66
      12'hC5A: dout  = 8'b10101110; // 3162 : 174 - 0xae
      12'hC5B: dout  = 8'b01001100; // 3163 :  76 - 0x4c
      12'hC5C: dout  = 8'b00111100; // 3164 :  60 - 0x3c
      12'hC5D: dout  = 8'b11111000; // 3165 : 248 - 0xf8
      12'hC5E: dout  = 8'b11100000; // 3166 : 224 - 0xe0
      12'hC5F: dout  = 8'b00000000; // 3167 :   0 - 0x0
      12'hC60: dout  = 8'b00000000; // 3168 :   0 - 0x0 -- Background 0x8c
      12'hC61: dout  = 8'b00000111; // 3169 :   7 - 0x7
      12'hC62: dout  = 8'b00011111; // 3170 :  31 - 0x1f
      12'hC63: dout  = 8'b00111111; // 3171 :  63 - 0x3f
      12'hC64: dout  = 8'b00111111; // 3172 :  63 - 0x3f
      12'hC65: dout  = 8'b01111111; // 3173 : 127 - 0x7f
      12'hC66: dout  = 8'b01111111; // 3174 : 127 - 0x7f
      12'hC67: dout  = 8'b01111111; // 3175 : 127 - 0x7f
      12'hC68: dout  = 8'b01111111; // 3176 : 127 - 0x7f -- Background 0x8d
      12'hC69: dout  = 8'b01111111; // 3177 : 127 - 0x7f
      12'hC6A: dout  = 8'b01111111; // 3178 : 127 - 0x7f
      12'hC6B: dout  = 8'b00111111; // 3179 :  63 - 0x3f
      12'hC6C: dout  = 8'b00111111; // 3180 :  63 - 0x3f
      12'hC6D: dout  = 8'b00011111; // 3181 :  31 - 0x1f
      12'hC6E: dout  = 8'b00000111; // 3182 :   7 - 0x7
      12'hC6F: dout  = 8'b00000000; // 3183 :   0 - 0x0
      12'hC70: dout  = 8'b00000000; // 3184 :   0 - 0x0 -- Background 0x8e
      12'hC71: dout  = 8'b11100000; // 3185 : 224 - 0xe0
      12'hC72: dout  = 8'b11111000; // 3186 : 248 - 0xf8
      12'hC73: dout  = 8'b11111100; // 3187 : 252 - 0xfc
      12'hC74: dout  = 8'b11111100; // 3188 : 252 - 0xfc
      12'hC75: dout  = 8'b11111110; // 3189 : 254 - 0xfe
      12'hC76: dout  = 8'b11111110; // 3190 : 254 - 0xfe
      12'hC77: dout  = 8'b11111110; // 3191 : 254 - 0xfe
      12'hC78: dout  = 8'b11111110; // 3192 : 254 - 0xfe -- Background 0x8f
      12'hC79: dout  = 8'b11111110; // 3193 : 254 - 0xfe
      12'hC7A: dout  = 8'b11111110; // 3194 : 254 - 0xfe
      12'hC7B: dout  = 8'b11111100; // 3195 : 252 - 0xfc
      12'hC7C: dout  = 8'b11111100; // 3196 : 252 - 0xfc
      12'hC7D: dout  = 8'b11111000; // 3197 : 248 - 0xf8
      12'hC7E: dout  = 8'b11100000; // 3198 : 224 - 0xe0
      12'hC7F: dout  = 8'b00000000; // 3199 :   0 - 0x0
      12'hC80: dout  = 8'b00000000; // 3200 :   0 - 0x0 -- Background 0x90
      12'hC81: dout  = 8'b00000000; // 3201 :   0 - 0x0
      12'hC82: dout  = 8'b00000000; // 3202 :   0 - 0x0
      12'hC83: dout  = 8'b00000000; // 3203 :   0 - 0x0
      12'hC84: dout  = 8'b00010000; // 3204 :  16 - 0x10
      12'hC85: dout  = 8'b00011100; // 3205 :  28 - 0x1c
      12'hC86: dout  = 8'b00001110; // 3206 :  14 - 0xe
      12'hC87: dout  = 8'b00000111; // 3207 :   7 - 0x7
      12'hC88: dout  = 8'b00000011; // 3208 :   3 - 0x3 -- Background 0x91
      12'hC89: dout  = 8'b00000001; // 3209 :   1 - 0x1
      12'hC8A: dout  = 8'b00110000; // 3210 :  48 - 0x30
      12'hC8B: dout  = 8'b00001111; // 3211 :  15 - 0xf
      12'hC8C: dout  = 8'b00000011; // 3212 :   3 - 0x3
      12'hC8D: dout  = 8'b00000000; // 3213 :   0 - 0x0
      12'hC8E: dout  = 8'b01111111; // 3214 : 127 - 0x7f
      12'hC8F: dout  = 8'b00000000; // 3215 :   0 - 0x0
      12'hC90: dout  = 8'b00000000; // 3216 :   0 - 0x0 -- Background 0x92
      12'hC91: dout  = 8'b01000010; // 3217 :  66 - 0x42
      12'hC92: dout  = 8'b01000010; // 3218 :  66 - 0x42
      12'hC93: dout  = 8'b01100110; // 3219 : 102 - 0x66
      12'hC94: dout  = 8'b01100110; // 3220 : 102 - 0x66
      12'hC95: dout  = 8'b01100110; // 3221 : 102 - 0x66
      12'hC96: dout  = 8'b11111110; // 3222 : 254 - 0xfe
      12'hC97: dout  = 8'b11111111; // 3223 : 255 - 0xff
      12'hC98: dout  = 8'b01111110; // 3224 : 126 - 0x7e -- Background 0x93
      12'hC99: dout  = 8'b01111110; // 3225 : 126 - 0x7e
      12'hC9A: dout  = 8'b01111110; // 3226 : 126 - 0x7e
      12'hC9B: dout  = 8'b01111110; // 3227 : 126 - 0x7e
      12'hC9C: dout  = 8'b01111110; // 3228 : 126 - 0x7e
      12'hC9D: dout  = 8'b01111110; // 3229 : 126 - 0x7e
      12'hC9E: dout  = 8'b01111110; // 3230 : 126 - 0x7e
      12'hC9F: dout  = 8'b01111110; // 3231 : 126 - 0x7e
      12'hCA0: dout  = 8'b00000000; // 3232 :   0 - 0x0 -- Background 0x94
      12'hCA1: dout  = 8'b00000000; // 3233 :   0 - 0x0
      12'hCA2: dout  = 8'b00000000; // 3234 :   0 - 0x0
      12'hCA3: dout  = 8'b00000000; // 3235 :   0 - 0x0
      12'hCA4: dout  = 8'b00001000; // 3236 :   8 - 0x8
      12'hCA5: dout  = 8'b00111000; // 3237 :  56 - 0x38
      12'hCA6: dout  = 8'b01110000; // 3238 : 112 - 0x70
      12'hCA7: dout  = 8'b11100000; // 3239 : 224 - 0xe0
      12'hCA8: dout  = 8'b11000000; // 3240 : 192 - 0xc0 -- Background 0x95
      12'hCA9: dout  = 8'b10000000; // 3241 : 128 - 0x80
      12'hCAA: dout  = 8'b00001100; // 3242 :  12 - 0xc
      12'hCAB: dout  = 8'b11110000; // 3243 : 240 - 0xf0
      12'hCAC: dout  = 8'b11000000; // 3244 : 192 - 0xc0
      12'hCAD: dout  = 8'b00000000; // 3245 :   0 - 0x0
      12'hCAE: dout  = 8'b11111110; // 3246 : 254 - 0xfe
      12'hCAF: dout  = 8'b00000000; // 3247 :   0 - 0x0
      12'hCB0: dout  = 8'b00000000; // 3248 :   0 - 0x0 -- Background 0x96
      12'hCB1: dout  = 8'b00111111; // 3249 :  63 - 0x3f
      12'hCB2: dout  = 8'b01111111; // 3250 : 127 - 0x7f
      12'hCB3: dout  = 8'b01111111; // 3251 : 127 - 0x7f
      12'hCB4: dout  = 8'b01111111; // 3252 : 127 - 0x7f
      12'hCB5: dout  = 8'b01111111; // 3253 : 127 - 0x7f
      12'hCB6: dout  = 8'b01111111; // 3254 : 127 - 0x7f
      12'hCB7: dout  = 8'b01111111; // 3255 : 127 - 0x7f
      12'hCB8: dout  = 8'b01111111; // 3256 : 127 - 0x7f -- Background 0x97
      12'hCB9: dout  = 8'b01111111; // 3257 : 127 - 0x7f
      12'hCBA: dout  = 8'b00111111; // 3258 :  63 - 0x3f
      12'hCBB: dout  = 8'b01111111; // 3259 : 127 - 0x7f
      12'hCBC: dout  = 8'b01111111; // 3260 : 127 - 0x7f
      12'hCBD: dout  = 8'b01111111; // 3261 : 127 - 0x7f
      12'hCBE: dout  = 8'b01111111; // 3262 : 127 - 0x7f
      12'hCBF: dout  = 8'b01111111; // 3263 : 127 - 0x7f
      12'hCC0: dout  = 8'b00000000; // 3264 :   0 - 0x0 -- Background 0x98
      12'hCC1: dout  = 8'b11011111; // 3265 : 223 - 0xdf
      12'hCC2: dout  = 8'b11111111; // 3266 : 255 - 0xff
      12'hCC3: dout  = 8'b11111111; // 3267 : 255 - 0xff
      12'hCC4: dout  = 8'b11111111; // 3268 : 255 - 0xff
      12'hCC5: dout  = 8'b11111111; // 3269 : 255 - 0xff
      12'hCC6: dout  = 8'b11111111; // 3270 : 255 - 0xff
      12'hCC7: dout  = 8'b11111111; // 3271 : 255 - 0xff
      12'hCC8: dout  = 8'b11111111; // 3272 : 255 - 0xff -- Background 0x99
      12'hCC9: dout  = 8'b11111111; // 3273 : 255 - 0xff
      12'hCCA: dout  = 8'b10111111; // 3274 : 191 - 0xbf
      12'hCCB: dout  = 8'b11111111; // 3275 : 255 - 0xff
      12'hCCC: dout  = 8'b11111111; // 3276 : 255 - 0xff
      12'hCCD: dout  = 8'b11111111; // 3277 : 255 - 0xff
      12'hCCE: dout  = 8'b11111111; // 3278 : 255 - 0xff
      12'hCCF: dout  = 8'b11111111; // 3279 : 255 - 0xff
      12'hCD0: dout  = 8'b00000000; // 3280 :   0 - 0x0 -- Background 0x9a
      12'hCD1: dout  = 8'b10111100; // 3281 : 188 - 0xbc
      12'hCD2: dout  = 8'b11111110; // 3282 : 254 - 0xfe
      12'hCD3: dout  = 8'b11111110; // 3283 : 254 - 0xfe
      12'hCD4: dout  = 8'b11111110; // 3284 : 254 - 0xfe
      12'hCD5: dout  = 8'b11111110; // 3285 : 254 - 0xfe
      12'hCD6: dout  = 8'b11111110; // 3286 : 254 - 0xfe
      12'hCD7: dout  = 8'b11111110; // 3287 : 254 - 0xfe
      12'hCD8: dout  = 8'b11111110; // 3288 : 254 - 0xfe -- Background 0x9b
      12'hCD9: dout  = 8'b11111110; // 3289 : 254 - 0xfe
      12'hCDA: dout  = 8'b10111110; // 3290 : 190 - 0xbe
      12'hCDB: dout  = 8'b11111110; // 3291 : 254 - 0xfe
      12'hCDC: dout  = 8'b11111110; // 3292 : 254 - 0xfe
      12'hCDD: dout  = 8'b11111110; // 3293 : 254 - 0xfe
      12'hCDE: dout  = 8'b11111110; // 3294 : 254 - 0xfe
      12'hCDF: dout  = 8'b11111110; // 3295 : 254 - 0xfe
      12'hCE0: dout  = 8'b00000000; // 3296 :   0 - 0x0 -- Background 0x9c
      12'hCE1: dout  = 8'b00111111; // 3297 :  63 - 0x3f
      12'hCE2: dout  = 8'b01011111; // 3298 :  95 - 0x5f
      12'hCE3: dout  = 8'b01101111; // 3299 : 111 - 0x6f
      12'hCE4: dout  = 8'b01110111; // 3300 : 119 - 0x77
      12'hCE5: dout  = 8'b01111011; // 3301 : 123 - 0x7b
      12'hCE6: dout  = 8'b00010101; // 3302 :  21 - 0x15
      12'hCE7: dout  = 8'b00000000; // 3303 :   0 - 0x0
      12'hCE8: dout  = 8'b00000000; // 3304 :   0 - 0x0 -- Background 0x9d
      12'hCE9: dout  = 8'b10111110; // 3305 : 190 - 0xbe
      12'hCEA: dout  = 8'b11011110; // 3306 : 222 - 0xde
      12'hCEB: dout  = 8'b11101110; // 3307 : 238 - 0xee
      12'hCEC: dout  = 8'b11110110; // 3308 : 246 - 0xf6
      12'hCED: dout  = 8'b11111010; // 3309 : 250 - 0xfa
      12'hCEE: dout  = 8'b01010100; // 3310 :  84 - 0x54
      12'hCEF: dout  = 8'b00000000; // 3311 :   0 - 0x0
      12'hCF0: dout  = 8'b00000000; // 3312 :   0 - 0x0 -- Background 0x9e
      12'hCF1: dout  = 8'b10111111; // 3313 : 191 - 0xbf
      12'hCF2: dout  = 8'b11011111; // 3314 : 223 - 0xdf
      12'hCF3: dout  = 8'b11101111; // 3315 : 239 - 0xef
      12'hCF4: dout  = 8'b11110111; // 3316 : 247 - 0xf7
      12'hCF5: dout  = 8'b11111011; // 3317 : 251 - 0xfb
      12'hCF6: dout  = 8'b01010101; // 3318 :  85 - 0x55
      12'hCF7: dout  = 8'b00000000; // 3319 :   0 - 0x0
      12'hCF8: dout  = 8'b00000000; // 3320 :   0 - 0x0 -- Background 0x9f
      12'hCF9: dout  = 8'b00000000; // 3321 :   0 - 0x0
      12'hCFA: dout  = 8'b00000000; // 3322 :   0 - 0x0
      12'hCFB: dout  = 8'b00000000; // 3323 :   0 - 0x0
      12'hCFC: dout  = 8'b00000000; // 3324 :   0 - 0x0
      12'hCFD: dout  = 8'b00000000; // 3325 :   0 - 0x0
      12'hCFE: dout  = 8'b00000000; // 3326 :   0 - 0x0
      12'hCFF: dout  = 8'b00000000; // 3327 :   0 - 0x0
      12'hD00: dout  = 8'b00000000; // 3328 :   0 - 0x0 -- Background 0xa0
      12'hD01: dout  = 8'b01111111; // 3329 : 127 - 0x7f
      12'hD02: dout  = 8'b00000000; // 3330 :   0 - 0x0
      12'hD03: dout  = 8'b00000001; // 3331 :   1 - 0x1
      12'hD04: dout  = 8'b00000001; // 3332 :   1 - 0x1
      12'hD05: dout  = 8'b00000001; // 3333 :   1 - 0x1
      12'hD06: dout  = 8'b00000001; // 3334 :   1 - 0x1
      12'hD07: dout  = 8'b00000001; // 3335 :   1 - 0x1
      12'hD08: dout  = 8'b00000001; // 3336 :   1 - 0x1 -- Background 0xa1
      12'hD09: dout  = 8'b00000001; // 3337 :   1 - 0x1
      12'hD0A: dout  = 8'b00000001; // 3338 :   1 - 0x1
      12'hD0B: dout  = 8'b00000001; // 3339 :   1 - 0x1
      12'hD0C: dout  = 8'b00000001; // 3340 :   1 - 0x1
      12'hD0D: dout  = 8'b00000001; // 3341 :   1 - 0x1
      12'hD0E: dout  = 8'b00000001; // 3342 :   1 - 0x1
      12'hD0F: dout  = 8'b00000001; // 3343 :   1 - 0x1
      12'hD10: dout  = 8'b00000000; // 3344 :   0 - 0x0 -- Background 0xa2
      12'hD11: dout  = 8'b11111110; // 3345 : 254 - 0xfe
      12'hD12: dout  = 8'b00000000; // 3346 :   0 - 0x0
      12'hD13: dout  = 8'b10000000; // 3347 : 128 - 0x80
      12'hD14: dout  = 8'b10000000; // 3348 : 128 - 0x80
      12'hD15: dout  = 8'b10000000; // 3349 : 128 - 0x80
      12'hD16: dout  = 8'b10000000; // 3350 : 128 - 0x80
      12'hD17: dout  = 8'b10000000; // 3351 : 128 - 0x80
      12'hD18: dout  = 8'b10000000; // 3352 : 128 - 0x80 -- Background 0xa3
      12'hD19: dout  = 8'b10000000; // 3353 : 128 - 0x80
      12'hD1A: dout  = 8'b10000000; // 3354 : 128 - 0x80
      12'hD1B: dout  = 8'b10000000; // 3355 : 128 - 0x80
      12'hD1C: dout  = 8'b10000000; // 3356 : 128 - 0x80
      12'hD1D: dout  = 8'b10000000; // 3357 : 128 - 0x80
      12'hD1E: dout  = 8'b10000000; // 3358 : 128 - 0x80
      12'hD1F: dout  = 8'b10000000; // 3359 : 128 - 0x80
      12'hD20: dout  = 8'b00000000; // 3360 :   0 - 0x0 -- Background 0xa4
      12'hD21: dout  = 8'b00110000; // 3361 :  48 - 0x30
      12'hD22: dout  = 8'b00111000; // 3362 :  56 - 0x38
      12'hD23: dout  = 8'b01111000; // 3363 : 120 - 0x78
      12'hD24: dout  = 8'b01111100; // 3364 : 124 - 0x7c
      12'hD25: dout  = 8'b01111101; // 3365 : 125 - 0x7d
      12'hD26: dout  = 8'b00011101; // 3366 :  29 - 0x1d
      12'hD27: dout  = 8'b00001101; // 3367 :  13 - 0xd
      12'hD28: dout  = 8'b00001101; // 3368 :  13 - 0xd -- Background 0xa5
      12'hD29: dout  = 8'b00011101; // 3369 :  29 - 0x1d
      12'hD2A: dout  = 8'b00111101; // 3370 :  61 - 0x3d
      12'hD2B: dout  = 8'b00111111; // 3371 :  63 - 0x3f
      12'hD2C: dout  = 8'b00111111; // 3372 :  63 - 0x3f
      12'hD2D: dout  = 8'b00011111; // 3373 :  31 - 0x1f
      12'hD2E: dout  = 8'b00000001; // 3374 :   1 - 0x1
      12'hD2F: dout  = 8'b00000000; // 3375 :   0 - 0x0
      12'hD30: dout  = 8'b00000000; // 3376 :   0 - 0x0 -- Background 0xa6
      12'hD31: dout  = 8'b00000000; // 3377 :   0 - 0x0
      12'hD32: dout  = 8'b11100000; // 3378 : 224 - 0xe0
      12'hD33: dout  = 8'b11111000; // 3379 : 248 - 0xf8
      12'hD34: dout  = 8'b11111000; // 3380 : 248 - 0xf8
      12'hD35: dout  = 8'b11110000; // 3381 : 240 - 0xf0
      12'hD36: dout  = 8'b11000000; // 3382 : 192 - 0xc0
      12'hD37: dout  = 8'b11000000; // 3383 : 192 - 0xc0
      12'hD38: dout  = 8'b11000000; // 3384 : 192 - 0xc0 -- Background 0xa7
      12'hD39: dout  = 8'b11110000; // 3385 : 240 - 0xf0
      12'hD3A: dout  = 8'b11110000; // 3386 : 240 - 0xf0
      12'hD3B: dout  = 8'b11000000; // 3387 : 192 - 0xc0
      12'hD3C: dout  = 8'b11000000; // 3388 : 192 - 0xc0
      12'hD3D: dout  = 8'b11000000; // 3389 : 192 - 0xc0
      12'hD3E: dout  = 8'b11000000; // 3390 : 192 - 0xc0
      12'hD3F: dout  = 8'b00000000; // 3391 :   0 - 0x0
      12'hD40: dout  = 8'b00000000; // 3392 :   0 - 0x0 -- Background 0xa8
      12'hD41: dout  = 8'b01100000; // 3393 :  96 - 0x60
      12'hD42: dout  = 8'b01100000; // 3394 :  96 - 0x60
      12'hD43: dout  = 8'b01100000; // 3395 :  96 - 0x60
      12'hD44: dout  = 8'b01100000; // 3396 :  96 - 0x60
      12'hD45: dout  = 8'b01100000; // 3397 :  96 - 0x60
      12'hD46: dout  = 8'b01100000; // 3398 :  96 - 0x60
      12'hD47: dout  = 8'b01100000; // 3399 :  96 - 0x60
      12'hD48: dout  = 8'b01100000; // 3400 :  96 - 0x60 -- Background 0xa9
      12'hD49: dout  = 8'b01100000; // 3401 :  96 - 0x60
      12'hD4A: dout  = 8'b01100000; // 3402 :  96 - 0x60
      12'hD4B: dout  = 8'b01100000; // 3403 :  96 - 0x60
      12'hD4C: dout  = 8'b01100000; // 3404 :  96 - 0x60
      12'hD4D: dout  = 8'b01100000; // 3405 :  96 - 0x60
      12'hD4E: dout  = 8'b01100000; // 3406 :  96 - 0x60
      12'hD4F: dout  = 8'b00000000; // 3407 :   0 - 0x0
      12'hD50: dout  = 8'b00000000; // 3408 :   0 - 0x0 -- Background 0xaa
      12'hD51: dout  = 8'b00000000; // 3409 :   0 - 0x0
      12'hD52: dout  = 8'b00000000; // 3410 :   0 - 0x0
      12'hD53: dout  = 8'b00000000; // 3411 :   0 - 0x0
      12'hD54: dout  = 8'b00000000; // 3412 :   0 - 0x0
      12'hD55: dout  = 8'b00000000; // 3413 :   0 - 0x0
      12'hD56: dout  = 8'b00000000; // 3414 :   0 - 0x0
      12'hD57: dout  = 8'b00000000; // 3415 :   0 - 0x0
      12'hD58: dout  = 8'b00000000; // 3416 :   0 - 0x0 -- Background 0xab
      12'hD59: dout  = 8'b00000000; // 3417 :   0 - 0x0
      12'hD5A: dout  = 8'b00000000; // 3418 :   0 - 0x0
      12'hD5B: dout  = 8'b00000000; // 3419 :   0 - 0x0
      12'hD5C: dout  = 8'b00000000; // 3420 :   0 - 0x0
      12'hD5D: dout  = 8'b00000000; // 3421 :   0 - 0x0
      12'hD5E: dout  = 8'b00000000; // 3422 :   0 - 0x0
      12'hD5F: dout  = 8'b00000000; // 3423 :   0 - 0x0
      12'hD60: dout  = 8'b00000000; // 3424 :   0 - 0x0 -- Background 0xac
      12'hD61: dout  = 8'b00000110; // 3425 :   6 - 0x6
      12'hD62: dout  = 8'b00000110; // 3426 :   6 - 0x6
      12'hD63: dout  = 8'b00000110; // 3427 :   6 - 0x6
      12'hD64: dout  = 8'b00000110; // 3428 :   6 - 0x6
      12'hD65: dout  = 8'b00000110; // 3429 :   6 - 0x6
      12'hD66: dout  = 8'b00000110; // 3430 :   6 - 0x6
      12'hD67: dout  = 8'b00000110; // 3431 :   6 - 0x6
      12'hD68: dout  = 8'b00000110; // 3432 :   6 - 0x6 -- Background 0xad
      12'hD69: dout  = 8'b00000110; // 3433 :   6 - 0x6
      12'hD6A: dout  = 8'b00000110; // 3434 :   6 - 0x6
      12'hD6B: dout  = 8'b00000110; // 3435 :   6 - 0x6
      12'hD6C: dout  = 8'b00000110; // 3436 :   6 - 0x6
      12'hD6D: dout  = 8'b00000110; // 3437 :   6 - 0x6
      12'hD6E: dout  = 8'b00000110; // 3438 :   6 - 0x6
      12'hD6F: dout  = 8'b00000000; // 3439 :   0 - 0x0
      12'hD70: dout  = 8'b00000000; // 3440 :   0 - 0x0 -- Background 0xae
      12'hD71: dout  = 8'b00000001; // 3441 :   1 - 0x1
      12'hD72: dout  = 8'b00000011; // 3442 :   3 - 0x3
      12'hD73: dout  = 8'b00000010; // 3443 :   2 - 0x2
      12'hD74: dout  = 8'b00000010; // 3444 :   2 - 0x2
      12'hD75: dout  = 8'b00000000; // 3445 :   0 - 0x0
      12'hD76: dout  = 8'b00000011; // 3446 :   3 - 0x3
      12'hD77: dout  = 8'b00000010; // 3447 :   2 - 0x2
      12'hD78: dout  = 8'b00000001; // 3448 :   1 - 0x1 -- Background 0xaf
      12'hD79: dout  = 8'b00000011; // 3449 :   3 - 0x3
      12'hD7A: dout  = 8'b00000101; // 3450 :   5 - 0x5
      12'hD7B: dout  = 8'b00000100; // 3451 :   4 - 0x4
      12'hD7C: dout  = 8'b00000101; // 3452 :   5 - 0x5
      12'hD7D: dout  = 8'b00001101; // 3453 :  13 - 0xd
      12'hD7E: dout  = 8'b00001100; // 3454 :  12 - 0xc
      12'hD7F: dout  = 8'b00000001; // 3455 :   1 - 0x1
      12'hD80: dout  = 8'b00000000; // 3456 :   0 - 0x0 -- Background 0xb0
      12'hD81: dout  = 8'b00000000; // 3457 :   0 - 0x0
      12'hD82: dout  = 8'b01000000; // 3458 :  64 - 0x40
      12'hD83: dout  = 8'b11110000; // 3459 : 240 - 0xf0
      12'hD84: dout  = 8'b11101000; // 3460 : 232 - 0xe8
      12'hD85: dout  = 8'b10010000; // 3461 : 144 - 0x90
      12'hD86: dout  = 8'b01010000; // 3462 :  80 - 0x50
      12'hD87: dout  = 8'b11010000; // 3463 : 208 - 0xd0
      12'hD88: dout  = 8'b11111000; // 3464 : 248 - 0xf8 -- Background 0xb1
      12'hD89: dout  = 8'b11000000; // 3465 : 192 - 0xc0
      12'hD8A: dout  = 8'b11100000; // 3466 : 224 - 0xe0
      12'hD8B: dout  = 8'b01000000; // 3467 :  64 - 0x40
      12'hD8C: dout  = 8'b10000000; // 3468 : 128 - 0x80
      12'hD8D: dout  = 8'b11000000; // 3469 : 192 - 0xc0
      12'hD8E: dout  = 8'b11100000; // 3470 : 224 - 0xe0
      12'hD8F: dout  = 8'b01110000; // 3471 : 112 - 0x70
      12'hD90: dout  = 8'b00000001; // 3472 :   1 - 0x1 -- Background 0xb2
      12'hD91: dout  = 8'b00001101; // 3473 :  13 - 0xd
      12'hD92: dout  = 8'b00001101; // 3474 :  13 - 0xd
      12'hD93: dout  = 8'b00000011; // 3475 :   3 - 0x3
      12'hD94: dout  = 8'b00000011; // 3476 :   3 - 0x3
      12'hD95: dout  = 8'b00000111; // 3477 :   7 - 0x7
      12'hD96: dout  = 8'b00000111; // 3478 :   7 - 0x7
      12'hD97: dout  = 8'b00000000; // 3479 :   0 - 0x0
      12'hD98: dout  = 8'b00111111; // 3480 :  63 - 0x3f -- Background 0xb3
      12'hD99: dout  = 8'b00111111; // 3481 :  63 - 0x3f
      12'hD9A: dout  = 8'b00111111; // 3482 :  63 - 0x3f
      12'hD9B: dout  = 8'b00111111; // 3483 :  63 - 0x3f
      12'hD9C: dout  = 8'b00111111; // 3484 :  63 - 0x3f
      12'hD9D: dout  = 8'b00111111; // 3485 :  63 - 0x3f
      12'hD9E: dout  = 8'b00110101; // 3486 :  53 - 0x35
      12'hD9F: dout  = 8'b00000000; // 3487 :   0 - 0x0
      12'hDA0: dout  = 8'b10110000; // 3488 : 176 - 0xb0 -- Background 0xb4
      12'hDA1: dout  = 8'b11000000; // 3489 : 192 - 0xc0
      12'hDA2: dout  = 8'b11100000; // 3490 : 224 - 0xe0
      12'hDA3: dout  = 8'b11100000; // 3491 : 224 - 0xe0
      12'hDA4: dout  = 8'b11110000; // 3492 : 240 - 0xf0
      12'hDA5: dout  = 8'b11110000; // 3493 : 240 - 0xf0
      12'hDA6: dout  = 8'b11110000; // 3494 : 240 - 0xf0
      12'hDA7: dout  = 8'b00000000; // 3495 :   0 - 0x0
      12'hDA8: dout  = 8'b11111100; // 3496 : 252 - 0xfc -- Background 0xb5
      12'hDA9: dout  = 8'b11111000; // 3497 : 248 - 0xf8
      12'hDAA: dout  = 8'b11111100; // 3498 : 252 - 0xfc
      12'hDAB: dout  = 8'b11111000; // 3499 : 248 - 0xf8
      12'hDAC: dout  = 8'b11111100; // 3500 : 252 - 0xfc
      12'hDAD: dout  = 8'b11111000; // 3501 : 248 - 0xf8
      12'hDAE: dout  = 8'b01010100; // 3502 :  84 - 0x54
      12'hDAF: dout  = 8'b00000000; // 3503 :   0 - 0x0
      12'hDB0: dout  = 8'b00000000; // 3504 :   0 - 0x0 -- Background 0xb6
      12'hDB1: dout  = 8'b01111111; // 3505 : 127 - 0x7f
      12'hDB2: dout  = 8'b01111111; // 3506 : 127 - 0x7f
      12'hDB3: dout  = 8'b01111111; // 3507 : 127 - 0x7f
      12'hDB4: dout  = 8'b01111111; // 3508 : 127 - 0x7f
      12'hDB5: dout  = 8'b01111111; // 3509 : 127 - 0x7f
      12'hDB6: dout  = 8'b01101010; // 3510 : 106 - 0x6a
      12'hDB7: dout  = 8'b00000000; // 3511 :   0 - 0x0
      12'hDB8: dout  = 8'b00000000; // 3512 :   0 - 0x0 -- Background 0xb7
      12'hDB9: dout  = 8'b01111011; // 3513 : 123 - 0x7b
      12'hDBA: dout  = 8'b01110011; // 3514 : 115 - 0x73
      12'hDBB: dout  = 8'b01111011; // 3515 : 123 - 0x7b
      12'hDBC: dout  = 8'b01110011; // 3516 : 115 - 0x73
      12'hDBD: dout  = 8'b01111011; // 3517 : 123 - 0x7b
      12'hDBE: dout  = 8'b01010011; // 3518 :  83 - 0x53
      12'hDBF: dout  = 8'b00000000; // 3519 :   0 - 0x0
      12'hDC0: dout  = 8'b00000000; // 3520 :   0 - 0x0 -- Background 0xb8
      12'hDC1: dout  = 8'b11011110; // 3521 : 222 - 0xde
      12'hDC2: dout  = 8'b10011110; // 3522 : 158 - 0x9e
      12'hDC3: dout  = 8'b11011100; // 3523 : 220 - 0xdc
      12'hDC4: dout  = 8'b10011110; // 3524 : 158 - 0x9e
      12'hDC5: dout  = 8'b11011100; // 3525 : 220 - 0xdc
      12'hDC6: dout  = 8'b10011010; // 3526 : 154 - 0x9a
      12'hDC7: dout  = 8'b00000000; // 3527 :   0 - 0x0
      12'hDC8: dout  = 8'b00000000; // 3528 :   0 - 0x0 -- Background 0xb9
      12'hDC9: dout  = 8'b11111110; // 3529 : 254 - 0xfe
      12'hDCA: dout  = 8'b11111100; // 3530 : 252 - 0xfc
      12'hDCB: dout  = 8'b11111110; // 3531 : 254 - 0xfe
      12'hDCC: dout  = 8'b11111100; // 3532 : 252 - 0xfc
      12'hDCD: dout  = 8'b11111110; // 3533 : 254 - 0xfe
      12'hDCE: dout  = 8'b01010100; // 3534 :  84 - 0x54
      12'hDCF: dout  = 8'b00000000; // 3535 :   0 - 0x0
      12'hDD0: dout  = 8'b00000000; // 3536 :   0 - 0x0 -- Background 0xba
      12'hDD1: dout  = 8'b01111111; // 3537 : 127 - 0x7f
      12'hDD2: dout  = 8'b01111111; // 3538 : 127 - 0x7f
      12'hDD3: dout  = 8'b00000000; // 3539 :   0 - 0x0
      12'hDD4: dout  = 8'b01111111; // 3540 : 127 - 0x7f
      12'hDD5: dout  = 8'b01111111; // 3541 : 127 - 0x7f
      12'hDD6: dout  = 8'b01101010; // 3542 : 106 - 0x6a
      12'hDD7: dout  = 8'b00000000; // 3543 :   0 - 0x0
      12'hDD8: dout  = 8'b00000000; // 3544 :   0 - 0x0 -- Background 0xbb
      12'hDD9: dout  = 8'b00000000; // 3545 :   0 - 0x0
      12'hDDA: dout  = 8'b00000000; // 3546 :   0 - 0x0
      12'hDDB: dout  = 8'b00000000; // 3547 :   0 - 0x0
      12'hDDC: dout  = 8'b00000000; // 3548 :   0 - 0x0
      12'hDDD: dout  = 8'b00000000; // 3549 :   0 - 0x0
      12'hDDE: dout  = 8'b00000000; // 3550 :   0 - 0x0
      12'hDDF: dout  = 8'b00000000; // 3551 :   0 - 0x0
      12'hDE0: dout  = 8'b00000000; // 3552 :   0 - 0x0 -- Background 0xbc
      12'hDE1: dout  = 8'b11111110; // 3553 : 254 - 0xfe
      12'hDE2: dout  = 8'b11111110; // 3554 : 254 - 0xfe
      12'hDE3: dout  = 8'b00000000; // 3555 :   0 - 0x0
      12'hDE4: dout  = 8'b10011110; // 3556 : 158 - 0x9e
      12'hDE5: dout  = 8'b11011100; // 3557 : 220 - 0xdc
      12'hDE6: dout  = 8'b10011010; // 3558 : 154 - 0x9a
      12'hDE7: dout  = 8'b00000000; // 3559 :   0 - 0x0
      12'hDE8: dout  = 8'b00000000; // 3560 :   0 - 0x0 -- Background 0xbd
      12'hDE9: dout  = 8'b00000000; // 3561 :   0 - 0x0
      12'hDEA: dout  = 8'b00000000; // 3562 :   0 - 0x0
      12'hDEB: dout  = 8'b00000000; // 3563 :   0 - 0x0
      12'hDEC: dout  = 8'b00000000; // 3564 :   0 - 0x0
      12'hDED: dout  = 8'b00000000; // 3565 :   0 - 0x0
      12'hDEE: dout  = 8'b00000000; // 3566 :   0 - 0x0
      12'hDEF: dout  = 8'b00000000; // 3567 :   0 - 0x0
      12'hDF0: dout  = 8'b00000000; // 3568 :   0 - 0x0 -- Background 0xbe
      12'hDF1: dout  = 8'b00000000; // 3569 :   0 - 0x0
      12'hDF2: dout  = 8'b00000000; // 3570 :   0 - 0x0
      12'hDF3: dout  = 8'b00000000; // 3571 :   0 - 0x0
      12'hDF4: dout  = 8'b00000000; // 3572 :   0 - 0x0
      12'hDF5: dout  = 8'b00000000; // 3573 :   0 - 0x0
      12'hDF6: dout  = 8'b00000000; // 3574 :   0 - 0x0
      12'hDF7: dout  = 8'b00000000; // 3575 :   0 - 0x0
      12'hDF8: dout  = 8'b00000000; // 3576 :   0 - 0x0 -- Background 0xbf
      12'hDF9: dout  = 8'b00000000; // 3577 :   0 - 0x0
      12'hDFA: dout  = 8'b00000000; // 3578 :   0 - 0x0
      12'hDFB: dout  = 8'b00000000; // 3579 :   0 - 0x0
      12'hDFC: dout  = 8'b00000000; // 3580 :   0 - 0x0
      12'hDFD: dout  = 8'b00000000; // 3581 :   0 - 0x0
      12'hDFE: dout  = 8'b00000000; // 3582 :   0 - 0x0
      12'hDFF: dout  = 8'b00000000; // 3583 :   0 - 0x0
      12'hE00: dout  = 8'b00000000; // 3584 :   0 - 0x0 -- Background 0xc0
      12'hE01: dout  = 8'b00000000; // 3585 :   0 - 0x0
      12'hE02: dout  = 8'b00000000; // 3586 :   0 - 0x0
      12'hE03: dout  = 8'b00000000; // 3587 :   0 - 0x0
      12'hE04: dout  = 8'b00000000; // 3588 :   0 - 0x0
      12'hE05: dout  = 8'b00000000; // 3589 :   0 - 0x0
      12'hE06: dout  = 8'b00000000; // 3590 :   0 - 0x0
      12'hE07: dout  = 8'b00000000; // 3591 :   0 - 0x0
      12'hE08: dout  = 8'b00000000; // 3592 :   0 - 0x0 -- Background 0xc1
      12'hE09: dout  = 8'b00000000; // 3593 :   0 - 0x0
      12'hE0A: dout  = 8'b00000000; // 3594 :   0 - 0x0
      12'hE0B: dout  = 8'b00000000; // 3595 :   0 - 0x0
      12'hE0C: dout  = 8'b00000000; // 3596 :   0 - 0x0
      12'hE0D: dout  = 8'b00000000; // 3597 :   0 - 0x0
      12'hE0E: dout  = 8'b00000000; // 3598 :   0 - 0x0
      12'hE0F: dout  = 8'b00000000; // 3599 :   0 - 0x0
      12'hE10: dout  = 8'b00000000; // 3600 :   0 - 0x0 -- Background 0xc2
      12'hE11: dout  = 8'b00000000; // 3601 :   0 - 0x0
      12'hE12: dout  = 8'b00000000; // 3602 :   0 - 0x0
      12'hE13: dout  = 8'b00000000; // 3603 :   0 - 0x0
      12'hE14: dout  = 8'b00000000; // 3604 :   0 - 0x0
      12'hE15: dout  = 8'b00000000; // 3605 :   0 - 0x0
      12'hE16: dout  = 8'b00000000; // 3606 :   0 - 0x0
      12'hE17: dout  = 8'b00000000; // 3607 :   0 - 0x0
      12'hE18: dout  = 8'b00000000; // 3608 :   0 - 0x0 -- Background 0xc3
      12'hE19: dout  = 8'b00000000; // 3609 :   0 - 0x0
      12'hE1A: dout  = 8'b00000000; // 3610 :   0 - 0x0
      12'hE1B: dout  = 8'b00000000; // 3611 :   0 - 0x0
      12'hE1C: dout  = 8'b00000000; // 3612 :   0 - 0x0
      12'hE1D: dout  = 8'b00000000; // 3613 :   0 - 0x0
      12'hE1E: dout  = 8'b00000000; // 3614 :   0 - 0x0
      12'hE1F: dout  = 8'b00000000; // 3615 :   0 - 0x0
      12'hE20: dout  = 8'b00000000; // 3616 :   0 - 0x0 -- Background 0xc4
      12'hE21: dout  = 8'b00000000; // 3617 :   0 - 0x0
      12'hE22: dout  = 8'b00000000; // 3618 :   0 - 0x0
      12'hE23: dout  = 8'b00000000; // 3619 :   0 - 0x0
      12'hE24: dout  = 8'b00000000; // 3620 :   0 - 0x0
      12'hE25: dout  = 8'b00000000; // 3621 :   0 - 0x0
      12'hE26: dout  = 8'b00000000; // 3622 :   0 - 0x0
      12'hE27: dout  = 8'b00000000; // 3623 :   0 - 0x0
      12'hE28: dout  = 8'b00000000; // 3624 :   0 - 0x0 -- Background 0xc5
      12'hE29: dout  = 8'b00000000; // 3625 :   0 - 0x0
      12'hE2A: dout  = 8'b00000000; // 3626 :   0 - 0x0
      12'hE2B: dout  = 8'b00000001; // 3627 :   1 - 0x1
      12'hE2C: dout  = 8'b00000111; // 3628 :   7 - 0x7
      12'hE2D: dout  = 8'b00001111; // 3629 :  15 - 0xf
      12'hE2E: dout  = 8'b00001111; // 3630 :  15 - 0xf
      12'hE2F: dout  = 8'b00011111; // 3631 :  31 - 0x1f
      12'hE30: dout  = 8'b00000000; // 3632 :   0 - 0x0 -- Background 0xc6
      12'hE31: dout  = 8'b00011111; // 3633 :  31 - 0x1f
      12'hE32: dout  = 8'b01111111; // 3634 : 127 - 0x7f
      12'hE33: dout  = 8'b11111111; // 3635 : 255 - 0xff
      12'hE34: dout  = 8'b11111111; // 3636 : 255 - 0xff
      12'hE35: dout  = 8'b11111111; // 3637 : 255 - 0xff
      12'hE36: dout  = 8'b11111111; // 3638 : 255 - 0xff
      12'hE37: dout  = 8'b11111111; // 3639 : 255 - 0xff
      12'hE38: dout  = 8'b00011111; // 3640 :  31 - 0x1f -- Background 0xc7
      12'hE39: dout  = 8'b00111111; // 3641 :  63 - 0x3f
      12'hE3A: dout  = 8'b00111111; // 3642 :  63 - 0x3f
      12'hE3B: dout  = 8'b01111111; // 3643 : 127 - 0x7f
      12'hE3C: dout  = 8'b01111111; // 3644 : 127 - 0x7f
      12'hE3D: dout  = 8'b01111111; // 3645 : 127 - 0x7f
      12'hE3E: dout  = 8'b01111111; // 3646 : 127 - 0x7f
      12'hE3F: dout  = 8'b01111111; // 3647 : 127 - 0x7f
      12'hE40: dout  = 8'b00000000; // 3648 :   0 - 0x0 -- Background 0xc8
      12'hE41: dout  = 8'b11111111; // 3649 : 255 - 0xff
      12'hE42: dout  = 8'b11111111; // 3650 : 255 - 0xff
      12'hE43: dout  = 8'b11111111; // 3651 : 255 - 0xff
      12'hE44: dout  = 8'b11111111; // 3652 : 255 - 0xff
      12'hE45: dout  = 8'b11111111; // 3653 : 255 - 0xff
      12'hE46: dout  = 8'b11111111; // 3654 : 255 - 0xff
      12'hE47: dout  = 8'b11111111; // 3655 : 255 - 0xff
      12'hE48: dout  = 8'b11101000; // 3656 : 232 - 0xe8 -- Background 0xc9
      12'hE49: dout  = 8'b11010100; // 3657 : 212 - 0xd4
      12'hE4A: dout  = 8'b11101000; // 3658 : 232 - 0xe8
      12'hE4B: dout  = 8'b11010100; // 3659 : 212 - 0xd4
      12'hE4C: dout  = 8'b11101010; // 3660 : 234 - 0xea
      12'hE4D: dout  = 8'b11010100; // 3661 : 212 - 0xd4
      12'hE4E: dout  = 8'b11101010; // 3662 : 234 - 0xea
      12'hE4F: dout  = 8'b11010100; // 3663 : 212 - 0xd4
      12'hE50: dout  = 8'b00000000; // 3664 :   0 - 0x0 -- Background 0xca
      12'hE51: dout  = 8'b00000000; // 3665 :   0 - 0x0
      12'hE52: dout  = 8'b00000000; // 3666 :   0 - 0x0
      12'hE53: dout  = 8'b00000000; // 3667 :   0 - 0x0
      12'hE54: dout  = 8'b00000000; // 3668 :   0 - 0x0
      12'hE55: dout  = 8'b00000000; // 3669 :   0 - 0x0
      12'hE56: dout  = 8'b00000000; // 3670 :   0 - 0x0
      12'hE57: dout  = 8'b00000000; // 3671 :   0 - 0x0
      12'hE58: dout  = 8'b00000000; // 3672 :   0 - 0x0 -- Background 0xcb
      12'hE59: dout  = 8'b00000000; // 3673 :   0 - 0x0
      12'hE5A: dout  = 8'b00000000; // 3674 :   0 - 0x0
      12'hE5B: dout  = 8'b00000000; // 3675 :   0 - 0x0
      12'hE5C: dout  = 8'b00000000; // 3676 :   0 - 0x0
      12'hE5D: dout  = 8'b00000000; // 3677 :   0 - 0x0
      12'hE5E: dout  = 8'b00000000; // 3678 :   0 - 0x0
      12'hE5F: dout  = 8'b00000000; // 3679 :   0 - 0x0
      12'hE60: dout  = 8'b00000000; // 3680 :   0 - 0x0 -- Background 0xcc
      12'hE61: dout  = 8'b00000000; // 3681 :   0 - 0x0
      12'hE62: dout  = 8'b00000000; // 3682 :   0 - 0x0
      12'hE63: dout  = 8'b00000000; // 3683 :   0 - 0x0
      12'hE64: dout  = 8'b00000101; // 3684 :   5 - 0x5
      12'hE65: dout  = 8'b00000010; // 3685 :   2 - 0x2
      12'hE66: dout  = 8'b00000001; // 3686 :   1 - 0x1
      12'hE67: dout  = 8'b00000000; // 3687 :   0 - 0x0
      12'hE68: dout  = 8'b00000000; // 3688 :   0 - 0x0 -- Background 0xcd
      12'hE69: dout  = 8'b00000000; // 3689 :   0 - 0x0
      12'hE6A: dout  = 8'b00000000; // 3690 :   0 - 0x0
      12'hE6B: dout  = 8'b10000000; // 3691 : 128 - 0x80
      12'hE6C: dout  = 8'b01010000; // 3692 :  80 - 0x50
      12'hE6D: dout  = 8'b10100000; // 3693 : 160 - 0xa0
      12'hE6E: dout  = 8'b01000000; // 3694 :  64 - 0x40
      12'hE6F: dout  = 8'b10000000; // 3695 : 128 - 0x80
      12'hE70: dout  = 8'b00000000; // 3696 :   0 - 0x0 -- Background 0xce
      12'hE71: dout  = 8'b00000000; // 3697 :   0 - 0x0
      12'hE72: dout  = 8'b00000000; // 3698 :   0 - 0x0
      12'hE73: dout  = 8'b00000000; // 3699 :   0 - 0x0
      12'hE74: dout  = 8'b00110000; // 3700 :  48 - 0x30
      12'hE75: dout  = 8'b01111111; // 3701 : 127 - 0x7f
      12'hE76: dout  = 8'b00110000; // 3702 :  48 - 0x30
      12'hE77: dout  = 8'b00110000; // 3703 :  48 - 0x30
      12'hE78: dout  = 8'b00000000; // 3704 :   0 - 0x0 -- Background 0xcf
      12'hE79: dout  = 8'b00000000; // 3705 :   0 - 0x0
      12'hE7A: dout  = 8'b00000000; // 3706 :   0 - 0x0
      12'hE7B: dout  = 8'b00000000; // 3707 :   0 - 0x0
      12'hE7C: dout  = 8'b00001100; // 3708 :  12 - 0xc
      12'hE7D: dout  = 8'b11111110; // 3709 : 254 - 0xfe
      12'hE7E: dout  = 8'b00001100; // 3710 :  12 - 0xc
      12'hE7F: dout  = 8'b00001100; // 3711 :  12 - 0xc
      12'hE80: dout  = 8'b00000000; // 3712 :   0 - 0x0 -- Background 0xd0
      12'hE81: dout  = 8'b00000000; // 3713 :   0 - 0x0
      12'hE82: dout  = 8'b00000000; // 3714 :   0 - 0x0
      12'hE83: dout  = 8'b00000000; // 3715 :   0 - 0x0
      12'hE84: dout  = 8'b00000000; // 3716 :   0 - 0x0
      12'hE85: dout  = 8'b00000000; // 3717 :   0 - 0x0
      12'hE86: dout  = 8'b00000000; // 3718 :   0 - 0x0
      12'hE87: dout  = 8'b00000000; // 3719 :   0 - 0x0
      12'hE88: dout  = 8'b00000000; // 3720 :   0 - 0x0 -- Background 0xd1
      12'hE89: dout  = 8'b00000000; // 3721 :   0 - 0x0
      12'hE8A: dout  = 8'b00000000; // 3722 :   0 - 0x0
      12'hE8B: dout  = 8'b00000000; // 3723 :   0 - 0x0
      12'hE8C: dout  = 8'b00000000; // 3724 :   0 - 0x0
      12'hE8D: dout  = 8'b00000000; // 3725 :   0 - 0x0
      12'hE8E: dout  = 8'b00000000; // 3726 :   0 - 0x0
      12'hE8F: dout  = 8'b00000000; // 3727 :   0 - 0x0
      12'hE90: dout  = 8'b00000111; // 3728 :   7 - 0x7 -- Background 0xd2
      12'hE91: dout  = 8'b00000111; // 3729 :   7 - 0x7
      12'hE92: dout  = 8'b00000111; // 3730 :   7 - 0x7
      12'hE93: dout  = 8'b00000111; // 3731 :   7 - 0x7
      12'hE94: dout  = 8'b00000111; // 3732 :   7 - 0x7
      12'hE95: dout  = 8'b00000111; // 3733 :   7 - 0x7
      12'hE96: dout  = 8'b00000111; // 3734 :   7 - 0x7
      12'hE97: dout  = 8'b00000111; // 3735 :   7 - 0x7
      12'hE98: dout  = 8'b11100000; // 3736 : 224 - 0xe0 -- Background 0xd3
      12'hE99: dout  = 8'b11100000; // 3737 : 224 - 0xe0
      12'hE9A: dout  = 8'b11000000; // 3738 : 192 - 0xc0
      12'hE9B: dout  = 8'b11100000; // 3739 : 224 - 0xe0
      12'hE9C: dout  = 8'b10100000; // 3740 : 160 - 0xa0
      12'hE9D: dout  = 8'b11100000; // 3741 : 224 - 0xe0
      12'hE9E: dout  = 8'b11000000; // 3742 : 192 - 0xc0
      12'hE9F: dout  = 8'b11100000; // 3743 : 224 - 0xe0
      12'hEA0: dout  = 8'b00000000; // 3744 :   0 - 0x0 -- Background 0xd4
      12'hEA1: dout  = 8'b00000000; // 3745 :   0 - 0x0
      12'hEA2: dout  = 8'b00000000; // 3746 :   0 - 0x0
      12'hEA3: dout  = 8'b00000000; // 3747 :   0 - 0x0
      12'hEA4: dout  = 8'b00000000; // 3748 :   0 - 0x0
      12'hEA5: dout  = 8'b00000000; // 3749 :   0 - 0x0
      12'hEA6: dout  = 8'b00000000; // 3750 :   0 - 0x0
      12'hEA7: dout  = 8'b00000000; // 3751 :   0 - 0x0
      12'hEA8: dout  = 8'b00000000; // 3752 :   0 - 0x0 -- Background 0xd5
      12'hEA9: dout  = 8'b11111000; // 3753 : 248 - 0xf8
      12'hEAA: dout  = 8'b11111110; // 3754 : 254 - 0xfe
      12'hEAB: dout  = 8'b11111111; // 3755 : 255 - 0xff
      12'hEAC: dout  = 8'b11111111; // 3756 : 255 - 0xff
      12'hEAD: dout  = 8'b11111111; // 3757 : 255 - 0xff
      12'hEAE: dout  = 8'b11111111; // 3758 : 255 - 0xff
      12'hEAF: dout  = 8'b11111111; // 3759 : 255 - 0xff
      12'hEB0: dout  = 8'b00000000; // 3760 :   0 - 0x0 -- Background 0xd6
      12'hEB1: dout  = 8'b00000000; // 3761 :   0 - 0x0
      12'hEB2: dout  = 8'b00000000; // 3762 :   0 - 0x0
      12'hEB3: dout  = 8'b10000000; // 3763 : 128 - 0x80
      12'hEB4: dout  = 8'b10100000; // 3764 : 160 - 0xa0
      12'hEB5: dout  = 8'b01010000; // 3765 :  80 - 0x50
      12'hEB6: dout  = 8'b10100000; // 3766 : 160 - 0xa0
      12'hEB7: dout  = 8'b11010000; // 3767 : 208 - 0xd0
      12'hEB8: dout  = 8'b01111111; // 3768 : 127 - 0x7f -- Background 0xd7
      12'hEB9: dout  = 8'b01111111; // 3769 : 127 - 0x7f
      12'hEBA: dout  = 8'b01111111; // 3770 : 127 - 0x7f
      12'hEBB: dout  = 8'b00111111; // 3771 :  63 - 0x3f
      12'hEBC: dout  = 8'b00111111; // 3772 :  63 - 0x3f
      12'hEBD: dout  = 8'b00001111; // 3773 :  15 - 0xf
      12'hEBE: dout  = 8'b00000111; // 3774 :   7 - 0x7
      12'hEBF: dout  = 8'b00000000; // 3775 :   0 - 0x0
      12'hEC0: dout  = 8'b11111111; // 3776 : 255 - 0xff -- Background 0xd8
      12'hEC1: dout  = 8'b11111111; // 3777 : 255 - 0xff
      12'hEC2: dout  = 8'b11111111; // 3778 : 255 - 0xff
      12'hEC3: dout  = 8'b11111111; // 3779 : 255 - 0xff
      12'hEC4: dout  = 8'b11111111; // 3780 : 255 - 0xff
      12'hEC5: dout  = 8'b11111111; // 3781 : 255 - 0xff
      12'hEC6: dout  = 8'b11111111; // 3782 : 255 - 0xff
      12'hEC7: dout  = 8'b00000000; // 3783 :   0 - 0x0
      12'hEC8: dout  = 8'b11101010; // 3784 : 234 - 0xea -- Background 0xd9
      12'hEC9: dout  = 8'b11010100; // 3785 : 212 - 0xd4
      12'hECA: dout  = 8'b11101010; // 3786 : 234 - 0xea
      12'hECB: dout  = 8'b11010100; // 3787 : 212 - 0xd4
      12'hECC: dout  = 8'b10101000; // 3788 : 168 - 0xa8
      12'hECD: dout  = 8'b01010000; // 3789 :  80 - 0x50
      12'hECE: dout  = 8'b10100000; // 3790 : 160 - 0xa0
      12'hECF: dout  = 8'b00000000; // 3791 :   0 - 0x0
      12'hED0: dout  = 8'b00000000; // 3792 :   0 - 0x0 -- Background 0xda
      12'hED1: dout  = 8'b00000000; // 3793 :   0 - 0x0
      12'hED2: dout  = 8'b00001100; // 3794 :  12 - 0xc
      12'hED3: dout  = 8'b00000000; // 3795 :   0 - 0x0
      12'hED4: dout  = 8'b00000000; // 3796 :   0 - 0x0
      12'hED5: dout  = 8'b00000000; // 3797 :   0 - 0x0
      12'hED6: dout  = 8'b00000000; // 3798 :   0 - 0x0
      12'hED7: dout  = 8'b00000000; // 3799 :   0 - 0x0
      12'hED8: dout  = 8'b00000000; // 3800 :   0 - 0x0 -- Background 0xdb
      12'hED9: dout  = 8'b10000000; // 3801 : 128 - 0x80
      12'hEDA: dout  = 8'b10000000; // 3802 : 128 - 0x80
      12'hEDB: dout  = 8'b10000000; // 3803 : 128 - 0x80
      12'hEDC: dout  = 8'b10011000; // 3804 : 152 - 0x98
      12'hEDD: dout  = 8'b10000000; // 3805 : 128 - 0x80
      12'hEDE: dout  = 8'b10000000; // 3806 : 128 - 0x80
      12'hEDF: dout  = 8'b10000000; // 3807 : 128 - 0x80
      12'hEE0: dout  = 8'b00000000; // 3808 :   0 - 0x0 -- Background 0xdc
      12'hEE1: dout  = 8'b00000000; // 3809 :   0 - 0x0
      12'hEE2: dout  = 8'b00000000; // 3810 :   0 - 0x0
      12'hEE3: dout  = 8'b00000000; // 3811 :   0 - 0x0
      12'hEE4: dout  = 8'b00000010; // 3812 :   2 - 0x2
      12'hEE5: dout  = 8'b00000011; // 3813 :   3 - 0x3
      12'hEE6: dout  = 8'b00000011; // 3814 :   3 - 0x3
      12'hEE7: dout  = 8'b00000001; // 3815 :   1 - 0x1
      12'hEE8: dout  = 8'b00000000; // 3816 :   0 - 0x0 -- Background 0xdd
      12'hEE9: dout  = 8'b00000000; // 3817 :   0 - 0x0
      12'hEEA: dout  = 8'b00000000; // 3818 :   0 - 0x0
      12'hEEB: dout  = 8'b00000000; // 3819 :   0 - 0x0
      12'hEEC: dout  = 8'b10100000; // 3820 : 160 - 0xa0
      12'hEED: dout  = 8'b11100000; // 3821 : 224 - 0xe0
      12'hEEE: dout  = 8'b11100000; // 3822 : 224 - 0xe0
      12'hEEF: dout  = 8'b11000000; // 3823 : 192 - 0xc0
      12'hEF0: dout  = 8'b00110000; // 3824 :  48 - 0x30 -- Background 0xde
      12'hEF1: dout  = 8'b01111111; // 3825 : 127 - 0x7f
      12'hEF2: dout  = 8'b00110000; // 3826 :  48 - 0x30
      12'hEF3: dout  = 8'b00110000; // 3827 :  48 - 0x30
      12'hEF4: dout  = 8'b00110000; // 3828 :  48 - 0x30
      12'hEF5: dout  = 8'b00110000; // 3829 :  48 - 0x30
      12'hEF6: dout  = 8'b00110000; // 3830 :  48 - 0x30
      12'hEF7: dout  = 8'b00110000; // 3831 :  48 - 0x30
      12'hEF8: dout  = 8'b00001100; // 3832 :  12 - 0xc -- Background 0xdf
      12'hEF9: dout  = 8'b11111110; // 3833 : 254 - 0xfe
      12'hEFA: dout  = 8'b00001100; // 3834 :  12 - 0xc
      12'hEFB: dout  = 8'b00001100; // 3835 :  12 - 0xc
      12'hEFC: dout  = 8'b00001100; // 3836 :  12 - 0xc
      12'hEFD: dout  = 8'b00001100; // 3837 :  12 - 0xc
      12'hEFE: dout  = 8'b00001100; // 3838 :  12 - 0xc
      12'hEFF: dout  = 8'b00001100; // 3839 :  12 - 0xc
      12'hF00: dout  = 8'b00000000; // 3840 :   0 - 0x0 -- Background 0xe0
      12'hF01: dout  = 8'b00000000; // 3841 :   0 - 0x0
      12'hF02: dout  = 8'b00000000; // 3842 :   0 - 0x0
      12'hF03: dout  = 8'b00000000; // 3843 :   0 - 0x0
      12'hF04: dout  = 8'b00000000; // 3844 :   0 - 0x0
      12'hF05: dout  = 8'b00000000; // 3845 :   0 - 0x0
      12'hF06: dout  = 8'b00000000; // 3846 :   0 - 0x0
      12'hF07: dout  = 8'b00000000; // 3847 :   0 - 0x0
      12'hF08: dout  = 8'b00000000; // 3848 :   0 - 0x0 -- Background 0xe1
      12'hF09: dout  = 8'b00000000; // 3849 :   0 - 0x0
      12'hF0A: dout  = 8'b00000000; // 3850 :   0 - 0x0
      12'hF0B: dout  = 8'b00000000; // 3851 :   0 - 0x0
      12'hF0C: dout  = 8'b00000000; // 3852 :   0 - 0x0
      12'hF0D: dout  = 8'b00000000; // 3853 :   0 - 0x0
      12'hF0E: dout  = 8'b00000000; // 3854 :   0 - 0x0
      12'hF0F: dout  = 8'b00000000; // 3855 :   0 - 0x0
      12'hF10: dout  = 8'b00000000; // 3856 :   0 - 0x0 -- Background 0xe2
      12'hF11: dout  = 8'b00000000; // 3857 :   0 - 0x0
      12'hF12: dout  = 8'b00000000; // 3858 :   0 - 0x0
      12'hF13: dout  = 8'b00000000; // 3859 :   0 - 0x0
      12'hF14: dout  = 8'b00000000; // 3860 :   0 - 0x0
      12'hF15: dout  = 8'b00000000; // 3861 :   0 - 0x0
      12'hF16: dout  = 8'b00000000; // 3862 :   0 - 0x0
      12'hF17: dout  = 8'b00000000; // 3863 :   0 - 0x0
      12'hF18: dout  = 8'b00000000; // 3864 :   0 - 0x0 -- Background 0xe3
      12'hF19: dout  = 8'b00000000; // 3865 :   0 - 0x0
      12'hF1A: dout  = 8'b00000000; // 3866 :   0 - 0x0
      12'hF1B: dout  = 8'b00000000; // 3867 :   0 - 0x0
      12'hF1C: dout  = 8'b00000000; // 3868 :   0 - 0x0
      12'hF1D: dout  = 8'b00000000; // 3869 :   0 - 0x0
      12'hF1E: dout  = 8'b00000000; // 3870 :   0 - 0x0
      12'hF1F: dout  = 8'b00000000; // 3871 :   0 - 0x0
      12'hF20: dout  = 8'b00000000; // 3872 :   0 - 0x0 -- Background 0xe4
      12'hF21: dout  = 8'b00000000; // 3873 :   0 - 0x0
      12'hF22: dout  = 8'b00000000; // 3874 :   0 - 0x0
      12'hF23: dout  = 8'b00000000; // 3875 :   0 - 0x0
      12'hF24: dout  = 8'b00000000; // 3876 :   0 - 0x0
      12'hF25: dout  = 8'b00000000; // 3877 :   0 - 0x0
      12'hF26: dout  = 8'b00000000; // 3878 :   0 - 0x0
      12'hF27: dout  = 8'b00000000; // 3879 :   0 - 0x0
      12'hF28: dout  = 8'b00000000; // 3880 :   0 - 0x0 -- Background 0xe5
      12'hF29: dout  = 8'b00000000; // 3881 :   0 - 0x0
      12'hF2A: dout  = 8'b00000000; // 3882 :   0 - 0x0
      12'hF2B: dout  = 8'b00000000; // 3883 :   0 - 0x0
      12'hF2C: dout  = 8'b00000000; // 3884 :   0 - 0x0
      12'hF2D: dout  = 8'b00000000; // 3885 :   0 - 0x0
      12'hF2E: dout  = 8'b00000000; // 3886 :   0 - 0x0
      12'hF2F: dout  = 8'b00000000; // 3887 :   0 - 0x0
      12'hF30: dout  = 8'b00000000; // 3888 :   0 - 0x0 -- Background 0xe6
      12'hF31: dout  = 8'b00000000; // 3889 :   0 - 0x0
      12'hF32: dout  = 8'b00000000; // 3890 :   0 - 0x0
      12'hF33: dout  = 8'b00000000; // 3891 :   0 - 0x0
      12'hF34: dout  = 8'b00000000; // 3892 :   0 - 0x0
      12'hF35: dout  = 8'b00000000; // 3893 :   0 - 0x0
      12'hF36: dout  = 8'b00000000; // 3894 :   0 - 0x0
      12'hF37: dout  = 8'b00000000; // 3895 :   0 - 0x0
      12'hF38: dout  = 8'b00000000; // 3896 :   0 - 0x0 -- Background 0xe7
      12'hF39: dout  = 8'b00000000; // 3897 :   0 - 0x0
      12'hF3A: dout  = 8'b00000000; // 3898 :   0 - 0x0
      12'hF3B: dout  = 8'b00000000; // 3899 :   0 - 0x0
      12'hF3C: dout  = 8'b00000000; // 3900 :   0 - 0x0
      12'hF3D: dout  = 8'b00000000; // 3901 :   0 - 0x0
      12'hF3E: dout  = 8'b00000000; // 3902 :   0 - 0x0
      12'hF3F: dout  = 8'b00000000; // 3903 :   0 - 0x0
      12'hF40: dout  = 8'b00000000; // 3904 :   0 - 0x0 -- Background 0xe8
      12'hF41: dout  = 8'b00000000; // 3905 :   0 - 0x0
      12'hF42: dout  = 8'b00000000; // 3906 :   0 - 0x0
      12'hF43: dout  = 8'b00000000; // 3907 :   0 - 0x0
      12'hF44: dout  = 8'b00000000; // 3908 :   0 - 0x0
      12'hF45: dout  = 8'b00000000; // 3909 :   0 - 0x0
      12'hF46: dout  = 8'b00000000; // 3910 :   0 - 0x0
      12'hF47: dout  = 8'b00000000; // 3911 :   0 - 0x0
      12'hF48: dout  = 8'b00000000; // 3912 :   0 - 0x0 -- Background 0xe9
      12'hF49: dout  = 8'b00000000; // 3913 :   0 - 0x0
      12'hF4A: dout  = 8'b00000000; // 3914 :   0 - 0x0
      12'hF4B: dout  = 8'b00000000; // 3915 :   0 - 0x0
      12'hF4C: dout  = 8'b00000000; // 3916 :   0 - 0x0
      12'hF4D: dout  = 8'b00000000; // 3917 :   0 - 0x0
      12'hF4E: dout  = 8'b00000000; // 3918 :   0 - 0x0
      12'hF4F: dout  = 8'b00000000; // 3919 :   0 - 0x0
      12'hF50: dout  = 8'b00000000; // 3920 :   0 - 0x0 -- Background 0xea
      12'hF51: dout  = 8'b00000000; // 3921 :   0 - 0x0
      12'hF52: dout  = 8'b00000000; // 3922 :   0 - 0x0
      12'hF53: dout  = 8'b00000000; // 3923 :   0 - 0x0
      12'hF54: dout  = 8'b00000000; // 3924 :   0 - 0x0
      12'hF55: dout  = 8'b00000000; // 3925 :   0 - 0x0
      12'hF56: dout  = 8'b00000000; // 3926 :   0 - 0x0
      12'hF57: dout  = 8'b00000000; // 3927 :   0 - 0x0
      12'hF58: dout  = 8'b00000000; // 3928 :   0 - 0x0 -- Background 0xeb
      12'hF59: dout  = 8'b00000000; // 3929 :   0 - 0x0
      12'hF5A: dout  = 8'b00000000; // 3930 :   0 - 0x0
      12'hF5B: dout  = 8'b00000000; // 3931 :   0 - 0x0
      12'hF5C: dout  = 8'b00000000; // 3932 :   0 - 0x0
      12'hF5D: dout  = 8'b00000000; // 3933 :   0 - 0x0
      12'hF5E: dout  = 8'b00000000; // 3934 :   0 - 0x0
      12'hF5F: dout  = 8'b00000000; // 3935 :   0 - 0x0
      12'hF60: dout  = 8'b00000000; // 3936 :   0 - 0x0 -- Background 0xec
      12'hF61: dout  = 8'b00000000; // 3937 :   0 - 0x0
      12'hF62: dout  = 8'b00000000; // 3938 :   0 - 0x0
      12'hF63: dout  = 8'b00000000; // 3939 :   0 - 0x0
      12'hF64: dout  = 8'b00000000; // 3940 :   0 - 0x0
      12'hF65: dout  = 8'b00000000; // 3941 :   0 - 0x0
      12'hF66: dout  = 8'b00000000; // 3942 :   0 - 0x0
      12'hF67: dout  = 8'b00000000; // 3943 :   0 - 0x0
      12'hF68: dout  = 8'b00000000; // 3944 :   0 - 0x0 -- Background 0xed
      12'hF69: dout  = 8'b00000000; // 3945 :   0 - 0x0
      12'hF6A: dout  = 8'b00000000; // 3946 :   0 - 0x0
      12'hF6B: dout  = 8'b00000000; // 3947 :   0 - 0x0
      12'hF6C: dout  = 8'b00000000; // 3948 :   0 - 0x0
      12'hF6D: dout  = 8'b00000000; // 3949 :   0 - 0x0
      12'hF6E: dout  = 8'b00000000; // 3950 :   0 - 0x0
      12'hF6F: dout  = 8'b00000000; // 3951 :   0 - 0x0
      12'hF70: dout  = 8'b00000000; // 3952 :   0 - 0x0 -- Background 0xee
      12'hF71: dout  = 8'b00000000; // 3953 :   0 - 0x0
      12'hF72: dout  = 8'b00000000; // 3954 :   0 - 0x0
      12'hF73: dout  = 8'b00000000; // 3955 :   0 - 0x0
      12'hF74: dout  = 8'b00000000; // 3956 :   0 - 0x0
      12'hF75: dout  = 8'b00000000; // 3957 :   0 - 0x0
      12'hF76: dout  = 8'b00000000; // 3958 :   0 - 0x0
      12'hF77: dout  = 8'b00000000; // 3959 :   0 - 0x0
      12'hF78: dout  = 8'b00000000; // 3960 :   0 - 0x0 -- Background 0xef
      12'hF79: dout  = 8'b00000000; // 3961 :   0 - 0x0
      12'hF7A: dout  = 8'b00000000; // 3962 :   0 - 0x0
      12'hF7B: dout  = 8'b00000000; // 3963 :   0 - 0x0
      12'hF7C: dout  = 8'b00000000; // 3964 :   0 - 0x0
      12'hF7D: dout  = 8'b00000000; // 3965 :   0 - 0x0
      12'hF7E: dout  = 8'b00000000; // 3966 :   0 - 0x0
      12'hF7F: dout  = 8'b00000000; // 3967 :   0 - 0x0
      12'hF80: dout  = 8'b00000000; // 3968 :   0 - 0x0 -- Background 0xf0
      12'hF81: dout  = 8'b00000000; // 3969 :   0 - 0x0
      12'hF82: dout  = 8'b00000000; // 3970 :   0 - 0x0
      12'hF83: dout  = 8'b00000000; // 3971 :   0 - 0x0
      12'hF84: dout  = 8'b00000000; // 3972 :   0 - 0x0
      12'hF85: dout  = 8'b00000000; // 3973 :   0 - 0x0
      12'hF86: dout  = 8'b00000000; // 3974 :   0 - 0x0
      12'hF87: dout  = 8'b00000000; // 3975 :   0 - 0x0
      12'hF88: dout  = 8'b00000000; // 3976 :   0 - 0x0 -- Background 0xf1
      12'hF89: dout  = 8'b00000000; // 3977 :   0 - 0x0
      12'hF8A: dout  = 8'b00000000; // 3978 :   0 - 0x0
      12'hF8B: dout  = 8'b00000000; // 3979 :   0 - 0x0
      12'hF8C: dout  = 8'b00000000; // 3980 :   0 - 0x0
      12'hF8D: dout  = 8'b00000000; // 3981 :   0 - 0x0
      12'hF8E: dout  = 8'b00000000; // 3982 :   0 - 0x0
      12'hF8F: dout  = 8'b00000000; // 3983 :   0 - 0x0
      12'hF90: dout  = 8'b00000000; // 3984 :   0 - 0x0 -- Background 0xf2
      12'hF91: dout  = 8'b00000000; // 3985 :   0 - 0x0
      12'hF92: dout  = 8'b00000000; // 3986 :   0 - 0x0
      12'hF93: dout  = 8'b00000000; // 3987 :   0 - 0x0
      12'hF94: dout  = 8'b00000000; // 3988 :   0 - 0x0
      12'hF95: dout  = 8'b00000000; // 3989 :   0 - 0x0
      12'hF96: dout  = 8'b00000000; // 3990 :   0 - 0x0
      12'hF97: dout  = 8'b00000000; // 3991 :   0 - 0x0
      12'hF98: dout  = 8'b00000000; // 3992 :   0 - 0x0 -- Background 0xf3
      12'hF99: dout  = 8'b00000000; // 3993 :   0 - 0x0
      12'hF9A: dout  = 8'b00000000; // 3994 :   0 - 0x0
      12'hF9B: dout  = 8'b00000000; // 3995 :   0 - 0x0
      12'hF9C: dout  = 8'b00000000; // 3996 :   0 - 0x0
      12'hF9D: dout  = 8'b00000000; // 3997 :   0 - 0x0
      12'hF9E: dout  = 8'b00000000; // 3998 :   0 - 0x0
      12'hF9F: dout  = 8'b00000000; // 3999 :   0 - 0x0
      12'hFA0: dout  = 8'b00000000; // 4000 :   0 - 0x0 -- Background 0xf4
      12'hFA1: dout  = 8'b00000000; // 4001 :   0 - 0x0
      12'hFA2: dout  = 8'b00000000; // 4002 :   0 - 0x0
      12'hFA3: dout  = 8'b00000000; // 4003 :   0 - 0x0
      12'hFA4: dout  = 8'b00000000; // 4004 :   0 - 0x0
      12'hFA5: dout  = 8'b00000000; // 4005 :   0 - 0x0
      12'hFA6: dout  = 8'b00000000; // 4006 :   0 - 0x0
      12'hFA7: dout  = 8'b00000000; // 4007 :   0 - 0x0
      12'hFA8: dout  = 8'b00000000; // 4008 :   0 - 0x0 -- Background 0xf5
      12'hFA9: dout  = 8'b00000000; // 4009 :   0 - 0x0
      12'hFAA: dout  = 8'b00000000; // 4010 :   0 - 0x0
      12'hFAB: dout  = 8'b00000000; // 4011 :   0 - 0x0
      12'hFAC: dout  = 8'b00000000; // 4012 :   0 - 0x0
      12'hFAD: dout  = 8'b00000000; // 4013 :   0 - 0x0
      12'hFAE: dout  = 8'b00000000; // 4014 :   0 - 0x0
      12'hFAF: dout  = 8'b00000000; // 4015 :   0 - 0x0
      12'hFB0: dout  = 8'b00000000; // 4016 :   0 - 0x0 -- Background 0xf6
      12'hFB1: dout  = 8'b00000000; // 4017 :   0 - 0x0
      12'hFB2: dout  = 8'b00000000; // 4018 :   0 - 0x0
      12'hFB3: dout  = 8'b00000000; // 4019 :   0 - 0x0
      12'hFB4: dout  = 8'b00000000; // 4020 :   0 - 0x0
      12'hFB5: dout  = 8'b00000000; // 4021 :   0 - 0x0
      12'hFB6: dout  = 8'b00000000; // 4022 :   0 - 0x0
      12'hFB7: dout  = 8'b00000000; // 4023 :   0 - 0x0
      12'hFB8: dout  = 8'b00000000; // 4024 :   0 - 0x0 -- Background 0xf7
      12'hFB9: dout  = 8'b00000000; // 4025 :   0 - 0x0
      12'hFBA: dout  = 8'b00000000; // 4026 :   0 - 0x0
      12'hFBB: dout  = 8'b00000000; // 4027 :   0 - 0x0
      12'hFBC: dout  = 8'b00000000; // 4028 :   0 - 0x0
      12'hFBD: dout  = 8'b00000000; // 4029 :   0 - 0x0
      12'hFBE: dout  = 8'b00000000; // 4030 :   0 - 0x0
      12'hFBF: dout  = 8'b00000000; // 4031 :   0 - 0x0
      12'hFC0: dout  = 8'b00000000; // 4032 :   0 - 0x0 -- Background 0xf8
      12'hFC1: dout  = 8'b00000000; // 4033 :   0 - 0x0
      12'hFC2: dout  = 8'b00000000; // 4034 :   0 - 0x0
      12'hFC3: dout  = 8'b00000000; // 4035 :   0 - 0x0
      12'hFC4: dout  = 8'b00000000; // 4036 :   0 - 0x0
      12'hFC5: dout  = 8'b00000000; // 4037 :   0 - 0x0
      12'hFC6: dout  = 8'b00000000; // 4038 :   0 - 0x0
      12'hFC7: dout  = 8'b00000000; // 4039 :   0 - 0x0
      12'hFC8: dout  = 8'b00000000; // 4040 :   0 - 0x0 -- Background 0xf9
      12'hFC9: dout  = 8'b00000000; // 4041 :   0 - 0x0
      12'hFCA: dout  = 8'b00000000; // 4042 :   0 - 0x0
      12'hFCB: dout  = 8'b00000000; // 4043 :   0 - 0x0
      12'hFCC: dout  = 8'b00000000; // 4044 :   0 - 0x0
      12'hFCD: dout  = 8'b00000000; // 4045 :   0 - 0x0
      12'hFCE: dout  = 8'b00000000; // 4046 :   0 - 0x0
      12'hFCF: dout  = 8'b00000000; // 4047 :   0 - 0x0
      12'hFD0: dout  = 8'b00000000; // 4048 :   0 - 0x0 -- Background 0xfa
      12'hFD1: dout  = 8'b00000000; // 4049 :   0 - 0x0
      12'hFD2: dout  = 8'b00000000; // 4050 :   0 - 0x0
      12'hFD3: dout  = 8'b00000000; // 4051 :   0 - 0x0
      12'hFD4: dout  = 8'b00000000; // 4052 :   0 - 0x0
      12'hFD5: dout  = 8'b00000000; // 4053 :   0 - 0x0
      12'hFD6: dout  = 8'b00000000; // 4054 :   0 - 0x0
      12'hFD7: dout  = 8'b00000000; // 4055 :   0 - 0x0
      12'hFD8: dout  = 8'b00000000; // 4056 :   0 - 0x0 -- Background 0xfb
      12'hFD9: dout  = 8'b00000000; // 4057 :   0 - 0x0
      12'hFDA: dout  = 8'b00000000; // 4058 :   0 - 0x0
      12'hFDB: dout  = 8'b00000000; // 4059 :   0 - 0x0
      12'hFDC: dout  = 8'b00000000; // 4060 :   0 - 0x0
      12'hFDD: dout  = 8'b00000000; // 4061 :   0 - 0x0
      12'hFDE: dout  = 8'b00000000; // 4062 :   0 - 0x0
      12'hFDF: dout  = 8'b00000000; // 4063 :   0 - 0x0
      12'hFE0: dout  = 8'b00000000; // 4064 :   0 - 0x0 -- Background 0xfc
      12'hFE1: dout  = 8'b00000000; // 4065 :   0 - 0x0
      12'hFE2: dout  = 8'b00000000; // 4066 :   0 - 0x0
      12'hFE3: dout  = 8'b00000000; // 4067 :   0 - 0x0
      12'hFE4: dout  = 8'b00000000; // 4068 :   0 - 0x0
      12'hFE5: dout  = 8'b00000000; // 4069 :   0 - 0x0
      12'hFE6: dout  = 8'b00000000; // 4070 :   0 - 0x0
      12'hFE7: dout  = 8'b00000000; // 4071 :   0 - 0x0
      12'hFE8: dout  = 8'b00000000; // 4072 :   0 - 0x0 -- Background 0xfd
      12'hFE9: dout  = 8'b00000000; // 4073 :   0 - 0x0
      12'hFEA: dout  = 8'b00000000; // 4074 :   0 - 0x0
      12'hFEB: dout  = 8'b00000000; // 4075 :   0 - 0x0
      12'hFEC: dout  = 8'b00000000; // 4076 :   0 - 0x0
      12'hFED: dout  = 8'b00000000; // 4077 :   0 - 0x0
      12'hFEE: dout  = 8'b00000000; // 4078 :   0 - 0x0
      12'hFEF: dout  = 8'b00000000; // 4079 :   0 - 0x0
      12'hFF0: dout  = 8'b00000000; // 4080 :   0 - 0x0 -- Background 0xfe
      12'hFF1: dout  = 8'b00000000; // 4081 :   0 - 0x0
      12'hFF2: dout  = 8'b00000000; // 4082 :   0 - 0x0
      12'hFF3: dout  = 8'b00000000; // 4083 :   0 - 0x0
      12'hFF4: dout  = 8'b00000000; // 4084 :   0 - 0x0
      12'hFF5: dout  = 8'b00000000; // 4085 :   0 - 0x0
      12'hFF6: dout  = 8'b00000000; // 4086 :   0 - 0x0
      12'hFF7: dout  = 8'b00000000; // 4087 :   0 - 0x0
      12'hFF8: dout  = 8'b00000000; // 4088 :   0 - 0x0 -- Background 0xff
      12'hFF9: dout  = 8'b00000000; // 4089 :   0 - 0x0
      12'hFFA: dout  = 8'b00000000; // 4090 :   0 - 0x0
      12'hFFB: dout  = 8'b00000000; // 4091 :   0 - 0x0
      12'hFFC: dout  = 8'b00000000; // 4092 :   0 - 0x0
      12'hFFD: dout  = 8'b00000000; // 4093 :   0 - 0x0
      12'hFFE: dout  = 8'b00000000; // 4094 :   0 - 0x0
      12'hFFF: dout  = 8'b00000000; // 4095 :   0 - 0x0
    endcase
  end

endmodule
