------- ROM creada automaticamente por ppm2rom -----------
------- Felipe Machado -----------------------------------
------- Area de Tecnologia Electronica -------------------
------- Universidad Rey Juan Carlos ----------------------
------- https://github.com/felipe-m ----------------------
----------------------------------------------------------
--------Datos de la imagen -------------------------------
--- Fichero original    : monster_16x16_rojo.ppm 
--- Filas    : 16 
--- Columnas : 16 
----------------------------------------------------------
--------Codificacion de la memoria------------------------
--- Palabras de 3 bits
--- De cada palabra hay 1 bit para cada color : "RGB" 8 colores



------ Puertos -------------------------------------------
-- Entradas ----------------------------------------------
--    clk  :  senal de reloj
--    addr :  direccion de la memoria
-- Salidas  ----------------------------------------------
--    dout :  dato de 3 bits de la direccion addr (un ciclo despues)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;
entity ROM_RGB_3b_monster_16x16_rojo is
  port (
    clk  : in  std_logic;   -- reloj
    addr : in  std_logic_vector(8-1 downto 0);
    dout : out std_logic_vector(3-1 downto 0) 
  );
end ROM_RGB_3b_monster_16x16_rojo;


architecture BEHAVIORAL of ROM_RGB_3b_monster_16x16_rojo is
  signal addr_int  : natural range 0 to 2**8-1;
  type memostruct is array (natural range<>) of std_logic_vector(3-1 downto 0);
  constant filaimg : memostruct := (
     --"RGB"
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "100",
       "100",
       "100",
       "100",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "000",
       "000",
       "000",
       "000",
       "000",
       "100",
       "111",
       "111",
       "100",
       "100",
       "100",
       "100",
       "111",
       "111",
       "100",
       "100",
       "100",
       "000",
       "000",
       "000",
       "000",
       "111",
       "111",
       "111",
       "111",
       "100",
       "100",
       "111",
       "111",
       "111",
       "111",
       "100",
       "100",
       "000",
       "000",
       "000",
       "000",
       "001",
       "001",
       "111",
       "111",
       "100",
       "100",
       "001",
       "001",
       "111",
       "111",
       "100",
       "100",
       "000",
       "000",
       "000",
       "100",
       "001",
       "001",
       "111",
       "111",
       "100",
       "100",
       "001",
       "001",
       "111",
       "111",
       "100",
       "100",
       "100",
       "000",
       "000",
       "100",
       "100",
       "111",
       "111",
       "100",
       "100",
       "100",
       "100",
       "111",
       "111",
       "100",
       "100",
       "100",
       "100",
       "000",
       "000",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "000",
       "000",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "000",
       "000",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "000",
       "000",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "100",
       "000",
       "000",
       "100",
       "100",
       "000",
       "100",
       "100",
       "100",
       "000",
       "000",
       "100",
       "100",
       "100",
       "000",
       "100",
       "100",
       "000",
       "000",
       "100",
       "000",
       "000",
       "000",
       "100",
       "100",
       "000",
       "000",
       "100",
       "100",
       "000",
       "000",
       "000",
       "100",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000",
       "000"
        );

begin

  addr_int <= TO_INTEGER(unsigned(addr));

  P_ROM: process (clk)
  begin
    if clk'event and clk='1' then
      dout <= filaimg(addr_int);
    end if;
  end process;

end BEHAVIORAL;

