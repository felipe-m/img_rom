--- Autcmatically generated VHDL ROM from a NES memory file----
---   NAME TABLE
-- https://wiki.nesdev.com/w/index.php/PPU_nametables
--- Only the first Name Table: 1KiB


---  Original memory dump file name: pacman_ntable_start.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory with clock ------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_NTABLE_PACMAN_START is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(10-1 downto 0);  --1024 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_NTABLE_PACMAN_START;

architecture BEHAVIORAL of ROM_NTABLE_PACMAN_START is
  signal addr_int  : natural range 0 to 2**10-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
     ------- Name Table 0---------
    "00100000", --    0 -  0x0  :   32 - 0x20 -- line 0x0
    "00100000", --    1 -  0x1  :   32 - 0x20
    "00100000", --    2 -  0x2  :   32 - 0x20
    "00100000", --    3 -  0x3  :   32 - 0x20
    "00100000", --    4 -  0x4  :   32 - 0x20
    "00100000", --    5 -  0x5  :   32 - 0x20
    "00100000", --    6 -  0x6  :   32 - 0x20
    "00100000", --    7 -  0x7  :   32 - 0x20
    "00100000", --    8 -  0x8  :   32 - 0x20
    "00100000", --    9 -  0x9  :   32 - 0x20
    "00100000", --   10 -  0xa  :   32 - 0x20
    "00100000", --   11 -  0xb  :   32 - 0x20
    "00100000", --   12 -  0xc  :   32 - 0x20
    "00100000", --   13 -  0xd  :   32 - 0x20
    "00100000", --   14 -  0xe  :   32 - 0x20
    "00100000", --   15 -  0xf  :   32 - 0x20
    "00100000", --   16 - 0x10  :   32 - 0x20
    "00100000", --   17 - 0x11  :   32 - 0x20
    "00100000", --   18 - 0x12  :   32 - 0x20
    "00100000", --   19 - 0x13  :   32 - 0x20
    "00100000", --   20 - 0x14  :   32 - 0x20
    "00100000", --   21 - 0x15  :   32 - 0x20
    "00100000", --   22 - 0x16  :   32 - 0x20
    "00100000", --   23 - 0x17  :   32 - 0x20
    "00100000", --   24 - 0x18  :   32 - 0x20
    "00100000", --   25 - 0x19  :   32 - 0x20
    "00100000", --   26 - 0x1a  :   32 - 0x20
    "00100000", --   27 - 0x1b  :   32 - 0x20
    "00100000", --   28 - 0x1c  :   32 - 0x20
    "00100000", --   29 - 0x1d  :   32 - 0x20
    "00100000", --   30 - 0x1e  :   32 - 0x20
    "00100000", --   31 - 0x1f  :   32 - 0x20
    "00100000", --   32 - 0x20  :   32 - 0x20 -- line 0x1
    "00100000", --   33 - 0x21  :   32 - 0x20
    "00100000", --   34 - 0x22  :   32 - 0x20
    "00100000", --   35 - 0x23  :   32 - 0x20
    "00100000", --   36 - 0x24  :   32 - 0x20
    "00100000", --   37 - 0x25  :   32 - 0x20
    "00100000", --   38 - 0x26  :   32 - 0x20
    "00100000", --   39 - 0x27  :   32 - 0x20
    "00100000", --   40 - 0x28  :   32 - 0x20
    "00100000", --   41 - 0x29  :   32 - 0x20
    "00100000", --   42 - 0x2a  :   32 - 0x20
    "00100000", --   43 - 0x2b  :   32 - 0x20
    "00100000", --   44 - 0x2c  :   32 - 0x20
    "00100000", --   45 - 0x2d  :   32 - 0x20
    "00100000", --   46 - 0x2e  :   32 - 0x20
    "00100000", --   47 - 0x2f  :   32 - 0x20
    "00100000", --   48 - 0x30  :   32 - 0x20
    "00100000", --   49 - 0x31  :   32 - 0x20
    "00100000", --   50 - 0x32  :   32 - 0x20
    "00100000", --   51 - 0x33  :   32 - 0x20
    "00100000", --   52 - 0x34  :   32 - 0x20
    "00100000", --   53 - 0x35  :   32 - 0x20
    "00100000", --   54 - 0x36  :   32 - 0x20
    "00100000", --   55 - 0x37  :   32 - 0x20
    "00100000", --   56 - 0x38  :   32 - 0x20
    "00100000", --   57 - 0x39  :   32 - 0x20
    "00100000", --   58 - 0x3a  :   32 - 0x20
    "00100000", --   59 - 0x3b  :   32 - 0x20
    "00100000", --   60 - 0x3c  :   32 - 0x20
    "00100000", --   61 - 0x3d  :   32 - 0x20
    "00100000", --   62 - 0x3e  :   32 - 0x20
    "00100000", --   63 - 0x3f  :   32 - 0x20
    "00100000", --   64 - 0x40  :   32 - 0x20 -- line 0x2
    "00100000", --   65 - 0x41  :   32 - 0x20
    "00100000", --   66 - 0x42  :   32 - 0x20
    "00100000", --   67 - 0x43  :   32 - 0x20
    "00100000", --   68 - 0x44  :   32 - 0x20
    "00100000", --   69 - 0x45  :   32 - 0x20
    "00100000", --   70 - 0x46  :   32 - 0x20
    "00100000", --   71 - 0x47  :   32 - 0x20
    "00100000", --   72 - 0x48  :   32 - 0x20
    "00100000", --   73 - 0x49  :   32 - 0x20
    "00100000", --   74 - 0x4a  :   32 - 0x20
    "00100000", --   75 - 0x4b  :   32 - 0x20
    "00100000", --   76 - 0x4c  :   32 - 0x20
    "00100000", --   77 - 0x4d  :   32 - 0x20
    "00100000", --   78 - 0x4e  :   32 - 0x20
    "00100000", --   79 - 0x4f  :   32 - 0x20
    "00100000", --   80 - 0x50  :   32 - 0x20
    "00100000", --   81 - 0x51  :   32 - 0x20
    "00100000", --   82 - 0x52  :   32 - 0x20
    "00100000", --   83 - 0x53  :   32 - 0x20
    "00100000", --   84 - 0x54  :   32 - 0x20
    "00100000", --   85 - 0x55  :   32 - 0x20
    "00100000", --   86 - 0x56  :   32 - 0x20
    "00100000", --   87 - 0x57  :   32 - 0x20
    "00100000", --   88 - 0x58  :   32 - 0x20
    "00100000", --   89 - 0x59  :   32 - 0x20
    "00100000", --   90 - 0x5a  :   32 - 0x20
    "00100000", --   91 - 0x5b  :   32 - 0x20
    "00100000", --   92 - 0x5c  :   32 - 0x20
    "00100000", --   93 - 0x5d  :   32 - 0x20
    "00100000", --   94 - 0x5e  :   32 - 0x20
    "00100000", --   95 - 0x5f  :   32 - 0x20
    "00100000", --   96 - 0x60  :   32 - 0x20 -- line 0x3
    "00100000", --   97 - 0x61  :   32 - 0x20
    "00100000", --   98 - 0x62  :   32 - 0x20
    "00100000", --   99 - 0x63  :   32 - 0x20
    "00100000", --  100 - 0x64  :   32 - 0x20
    "10110000", --  101 - 0x65  :  176 - 0xb0
    "10110011", --  102 - 0x66  :  179 - 0xb3
    "10110010", --  103 - 0x67  :  178 - 0xb2
    "00100000", --  104 - 0x68  :   32 - 0x20
    "00100000", --  105 - 0x69  :   32 - 0x20
    "00100000", --  106 - 0x6a  :   32 - 0x20
    "00100000", --  107 - 0x6b  :   32 - 0x20
    "10110100", --  108 - 0x6c  :  180 - 0xb4
    "10110101", --  109 - 0x6d  :  181 - 0xb5
    "10110110", --  110 - 0x6e  :  182 - 0xb6
    "10110111", --  111 - 0x6f  :  183 - 0xb7
    "10111000", --  112 - 0x70  :  184 - 0xb8
    "10111001", --  113 - 0x71  :  185 - 0xb9
    "10111010", --  114 - 0x72  :  186 - 0xba
    "10111011", --  115 - 0x73  :  187 - 0xbb
    "00100000", --  116 - 0x74  :   32 - 0x20
    "00100000", --  117 - 0x75  :   32 - 0x20
    "00100000", --  118 - 0x76  :   32 - 0x20
    "10110001", --  119 - 0x77  :  177 - 0xb1
    "10110011", --  120 - 0x78  :  179 - 0xb3
    "10110010", --  121 - 0x79  :  178 - 0xb2
    "00100000", --  122 - 0x7a  :   32 - 0x20
    "00100000", --  123 - 0x7b  :   32 - 0x20
    "00100000", --  124 - 0x7c  :   32 - 0x20
    "00100000", --  125 - 0x7d  :   32 - 0x20
    "00100000", --  126 - 0x7e  :   32 - 0x20
    "00100000", --  127 - 0x7f  :   32 - 0x20
    "00100000", --  128 - 0x80  :   32 - 0x20 -- line 0x4
    "00100000", --  129 - 0x81  :   32 - 0x20
    "00100000", --  130 - 0x82  :   32 - 0x20
    "00100000", --  131 - 0x83  :   32 - 0x20
    "00100000", --  132 - 0x84  :   32 - 0x20
    "00100000", --  133 - 0x85  :   32 - 0x20
    "00100000", --  134 - 0x86  :   32 - 0x20
    "00100000", --  135 - 0x87  :   32 - 0x20
    "00110101", --  136 - 0x88  :   53 - 0x35
    "00110000", --  137 - 0x89  :   48 - 0x30
    "00100000", --  138 - 0x8a  :   32 - 0x20
    "00100000", --  139 - 0x8b  :   32 - 0x20
    "00100000", --  140 - 0x8c  :   32 - 0x20
    "00100000", --  141 - 0x8d  :   32 - 0x20
    "00110001", --  142 - 0x8e  :   49 - 0x31
    "00110000", --  143 - 0x8f  :   48 - 0x30
    "00110000", --  144 - 0x90  :   48 - 0x30
    "00110000", --  145 - 0x91  :   48 - 0x30
    "00110000", --  146 - 0x92  :   48 - 0x30
    "00100000", --  147 - 0x93  :   32 - 0x20
    "00100000", --  148 - 0x94  :   32 - 0x20
    "00100000", --  149 - 0x95  :   32 - 0x20
    "00100000", --  150 - 0x96  :   32 - 0x20
    "00100000", --  151 - 0x97  :   32 - 0x20
    "00100000", --  152 - 0x98  :   32 - 0x20
    "00100000", --  153 - 0x99  :   32 - 0x20
    "00110000", --  154 - 0x9a  :   48 - 0x30
    "00110000", --  155 - 0x9b  :   48 - 0x30
    "00100000", --  156 - 0x9c  :   32 - 0x20
    "00100000", --  157 - 0x9d  :   32 - 0x20
    "00100000", --  158 - 0x9e  :   32 - 0x20
    "00100000", --  159 - 0x9f  :   32 - 0x20
    "00100000", --  160 - 0xa0  :   32 - 0x20 -- line 0x5
    "00100000", --  161 - 0xa1  :   32 - 0x20
    "00100000", --  162 - 0xa2  :   32 - 0x20
    "00100000", --  163 - 0xa3  :   32 - 0x20
    "00100000", --  164 - 0xa4  :   32 - 0x20
    "00100000", --  165 - 0xa5  :   32 - 0x20
    "00100000", --  166 - 0xa6  :   32 - 0x20
    "00100000", --  167 - 0xa7  :   32 - 0x20
    "00100000", --  168 - 0xa8  :   32 - 0x20
    "00100000", --  169 - 0xa9  :   32 - 0x20
    "00100000", --  170 - 0xaa  :   32 - 0x20
    "00100000", --  171 - 0xab  :   32 - 0x20
    "00100000", --  172 - 0xac  :   32 - 0x20
    "00100000", --  173 - 0xad  :   32 - 0x20
    "00100000", --  174 - 0xae  :   32 - 0x20
    "00100000", --  175 - 0xaf  :   32 - 0x20
    "00100000", --  176 - 0xb0  :   32 - 0x20
    "00100000", --  177 - 0xb1  :   32 - 0x20
    "00100000", --  178 - 0xb2  :   32 - 0x20
    "00100000", --  179 - 0xb3  :   32 - 0x20
    "00100000", --  180 - 0xb4  :   32 - 0x20
    "00100000", --  181 - 0xb5  :   32 - 0x20
    "00100000", --  182 - 0xb6  :   32 - 0x20
    "00100000", --  183 - 0xb7  :   32 - 0x20
    "00100000", --  184 - 0xb8  :   32 - 0x20
    "00100000", --  185 - 0xb9  :   32 - 0x20
    "00100000", --  186 - 0xba  :   32 - 0x20
    "00100000", --  187 - 0xbb  :   32 - 0x20
    "00100000", --  188 - 0xbc  :   32 - 0x20
    "00100000", --  189 - 0xbd  :   32 - 0x20
    "00100000", --  190 - 0xbe  :   32 - 0x20
    "00100000", --  191 - 0xbf  :   32 - 0x20
    "00100000", --  192 - 0xc0  :   32 - 0x20 -- line 0x6
    "00100000", --  193 - 0xc1  :   32 - 0x20
    "00100000", --  194 - 0xc2  :   32 - 0x20
    "00100000", --  195 - 0xc3  :   32 - 0x20
    "00100000", --  196 - 0xc4  :   32 - 0x20
    "00100000", --  197 - 0xc5  :   32 - 0x20
    "00100000", --  198 - 0xc6  :   32 - 0x20
    "00100000", --  199 - 0xc7  :   32 - 0x20
    "00100000", --  200 - 0xc8  :   32 - 0x20
    "00100000", --  201 - 0xc9  :   32 - 0x20
    "00100000", --  202 - 0xca  :   32 - 0x20
    "00100000", --  203 - 0xcb  :   32 - 0x20
    "00100000", --  204 - 0xcc  :   32 - 0x20
    "00100000", --  205 - 0xcd  :   32 - 0x20
    "00100000", --  206 - 0xce  :   32 - 0x20
    "00100000", --  207 - 0xcf  :   32 - 0x20
    "00100000", --  208 - 0xd0  :   32 - 0x20
    "00100000", --  209 - 0xd1  :   32 - 0x20
    "00100000", --  210 - 0xd2  :   32 - 0x20
    "00100000", --  211 - 0xd3  :   32 - 0x20
    "00100000", --  212 - 0xd4  :   32 - 0x20
    "00100000", --  213 - 0xd5  :   32 - 0x20
    "00100000", --  214 - 0xd6  :   32 - 0x20
    "00100000", --  215 - 0xd7  :   32 - 0x20
    "00100000", --  216 - 0xd8  :   32 - 0x20
    "00100000", --  217 - 0xd9  :   32 - 0x20
    "00100000", --  218 - 0xda  :   32 - 0x20
    "00100000", --  219 - 0xdb  :   32 - 0x20
    "00100000", --  220 - 0xdc  :   32 - 0x20
    "00100000", --  221 - 0xdd  :   32 - 0x20
    "00100000", --  222 - 0xde  :   32 - 0x20
    "00100000", --  223 - 0xdf  :   32 - 0x20
    "00100000", --  224 - 0xe0  :   32 - 0x20 -- line 0x7
    "00100000", --  225 - 0xe1  :   32 - 0x20
    "00100000", --  226 - 0xe2  :   32 - 0x20
    "00100000", --  227 - 0xe3  :   32 - 0x20
    "00100000", --  228 - 0xe4  :   32 - 0x20
    "11100100", --  229 - 0xe5  :  228 - 0xe4
    "11101000", --  230 - 0xe6  :  232 - 0xe8
    "11101000", --  231 - 0xe7  :  232 - 0xe8
    "11101000", --  232 - 0xe8  :  232 - 0xe8
    "11101000", --  233 - 0xe9  :  232 - 0xe8
    "11101000", --  234 - 0xea  :  232 - 0xe8
    "11101000", --  235 - 0xeb  :  232 - 0xe8
    "11101000", --  236 - 0xec  :  232 - 0xe8
    "11101000", --  237 - 0xed  :  232 - 0xe8
    "11101000", --  238 - 0xee  :  232 - 0xe8
    "11101000", --  239 - 0xef  :  232 - 0xe8
    "11101000", --  240 - 0xf0  :  232 - 0xe8
    "11101000", --  241 - 0xf1  :  232 - 0xe8
    "11101000", --  242 - 0xf2  :  232 - 0xe8
    "11101000", --  243 - 0xf3  :  232 - 0xe8
    "11101000", --  244 - 0xf4  :  232 - 0xe8
    "11101000", --  245 - 0xf5  :  232 - 0xe8
    "11101000", --  246 - 0xf6  :  232 - 0xe8
    "11101000", --  247 - 0xf7  :  232 - 0xe8
    "11101000", --  248 - 0xf8  :  232 - 0xe8
    "11101000", --  249 - 0xf9  :  232 - 0xe8
    "11101000", --  250 - 0xfa  :  232 - 0xe8
    "11100101", --  251 - 0xfb  :  229 - 0xe5
    "00100000", --  252 - 0xfc  :   32 - 0x20
    "00100000", --  253 - 0xfd  :   32 - 0x20
    "00100000", --  254 - 0xfe  :   32 - 0x20
    "00100000", --  255 - 0xff  :   32 - 0x20
    "00100000", --  256 - 0x100  :   32 - 0x20 -- line 0x8
    "00100000", --  257 - 0x101  :   32 - 0x20
    "00100000", --  258 - 0x102  :   32 - 0x20
    "00100000", --  259 - 0x103  :   32 - 0x20
    "00100000", --  260 - 0x104  :   32 - 0x20
    "11101011", --  261 - 0x105  :  235 - 0xeb
    "10001000", --  262 - 0x106  :  136 - 0x88
    "10000000", --  263 - 0x107  :  128 - 0x80
    "10000001", --  264 - 0x108  :  129 - 0x81
    "10000010", --  265 - 0x109  :  130 - 0x82
    "10000011", --  266 - 0x10a  :  131 - 0x83
    "10000100", --  267 - 0x10b  :  132 - 0x84
    "10000101", --  268 - 0x10c  :  133 - 0x85
    "10000110", --  269 - 0x10d  :  134 - 0x86
    "10000111", --  270 - 0x10e  :  135 - 0x87
    "10001000", --  271 - 0x10f  :  136 - 0x88
    "10001000", --  272 - 0x110  :  136 - 0x88
    "10001001", --  273 - 0x111  :  137 - 0x89
    "10001010", --  274 - 0x112  :  138 - 0x8a
    "10001011", --  275 - 0x113  :  139 - 0x8b
    "10001100", --  276 - 0x114  :  140 - 0x8c
    "10001101", --  277 - 0x115  :  141 - 0x8d
    "10001110", --  278 - 0x116  :  142 - 0x8e
    "10001111", --  279 - 0x117  :  143 - 0x8f
    "10010000", --  280 - 0x118  :  144 - 0x90
    "10010001", --  281 - 0x119  :  145 - 0x91
    "10100011", --  282 - 0x11a  :  163 - 0xa3
    "11101001", --  283 - 0x11b  :  233 - 0xe9
    "00100000", --  284 - 0x11c  :   32 - 0x20
    "00100000", --  285 - 0x11d  :   32 - 0x20
    "00100000", --  286 - 0x11e  :   32 - 0x20
    "00100000", --  287 - 0x11f  :   32 - 0x20
    "00100000", --  288 - 0x120  :   32 - 0x20 -- line 0x9
    "00100000", --  289 - 0x121  :   32 - 0x20
    "00100000", --  290 - 0x122  :   32 - 0x20
    "00100000", --  291 - 0x123  :   32 - 0x20
    "00100000", --  292 - 0x124  :   32 - 0x20
    "11101011", --  293 - 0x125  :  235 - 0xeb
    "10001000", --  294 - 0x126  :  136 - 0x88
    "10010010", --  295 - 0x127  :  146 - 0x92
    "10010011", --  296 - 0x128  :  147 - 0x93
    "10010100", --  297 - 0x129  :  148 - 0x94
    "10010101", --  298 - 0x12a  :  149 - 0x95
    "10010110", --  299 - 0x12b  :  150 - 0x96
    "10010111", --  300 - 0x12c  :  151 - 0x97
    "10011000", --  301 - 0x12d  :  152 - 0x98
    "10011001", --  302 - 0x12e  :  153 - 0x99
    "10011010", --  303 - 0x12f  :  154 - 0x9a
    "10011011", --  304 - 0x130  :  155 - 0x9b
    "10011100", --  305 - 0x131  :  156 - 0x9c
    "10011101", --  306 - 0x132  :  157 - 0x9d
    "10011110", --  307 - 0x133  :  158 - 0x9e
    "10011111", --  308 - 0x134  :  159 - 0x9f
    "10100000", --  309 - 0x135  :  160 - 0xa0
    "10100001", --  310 - 0x136  :  161 - 0xa1
    "10100010", --  311 - 0x137  :  162 - 0xa2
    "10100011", --  312 - 0x138  :  163 - 0xa3
    "10100100", --  313 - 0x139  :  164 - 0xa4
    "10100011", --  314 - 0x13a  :  163 - 0xa3
    "11101001", --  315 - 0x13b  :  233 - 0xe9
    "00100000", --  316 - 0x13c  :   32 - 0x20
    "00100000", --  317 - 0x13d  :   32 - 0x20
    "00100000", --  318 - 0x13e  :   32 - 0x20
    "00100000", --  319 - 0x13f  :   32 - 0x20
    "00100000", --  320 - 0x140  :   32 - 0x20 -- line 0xa
    "00100000", --  321 - 0x141  :   32 - 0x20
    "00100000", --  322 - 0x142  :   32 - 0x20
    "00100000", --  323 - 0x143  :   32 - 0x20
    "00100000", --  324 - 0x144  :   32 - 0x20
    "11101011", --  325 - 0x145  :  235 - 0xeb
    "10001000", --  326 - 0x146  :  136 - 0x88
    "10010010", --  327 - 0x147  :  146 - 0x92
    "10100101", --  328 - 0x148  :  165 - 0xa5
    "10100110", --  329 - 0x149  :  166 - 0xa6
    "10100111", --  330 - 0x14a  :  167 - 0xa7
    "10101000", --  331 - 0x14b  :  168 - 0xa8
    "10101001", --  332 - 0x14c  :  169 - 0xa9
    "10101010", --  333 - 0x14d  :  170 - 0xaa
    "10101011", --  334 - 0x14e  :  171 - 0xab
    "10101100", --  335 - 0x14f  :  172 - 0xac
    "10101101", --  336 - 0x150  :  173 - 0xad
    "10101110", --  337 - 0x151  :  174 - 0xae
    "10100011", --  338 - 0x152  :  163 - 0xa3
    "10101111", --  339 - 0x153  :  175 - 0xaf
    "11010000", --  340 - 0x154  :  208 - 0xd0
    "11010001", --  341 - 0x155  :  209 - 0xd1
    "11010010", --  342 - 0x156  :  210 - 0xd2
    "10100011", --  343 - 0x157  :  163 - 0xa3
    "11010011", --  344 - 0x158  :  211 - 0xd3
    "10100100", --  345 - 0x159  :  164 - 0xa4
    "10100011", --  346 - 0x15a  :  163 - 0xa3
    "11101001", --  347 - 0x15b  :  233 - 0xe9
    "00100000", --  348 - 0x15c  :   32 - 0x20
    "00100000", --  349 - 0x15d  :   32 - 0x20
    "00100000", --  350 - 0x15e  :   32 - 0x20
    "00100000", --  351 - 0x15f  :   32 - 0x20
    "00100000", --  352 - 0x160  :   32 - 0x20 -- line 0xb
    "00100000", --  353 - 0x161  :   32 - 0x20
    "00100000", --  354 - 0x162  :   32 - 0x20
    "00100000", --  355 - 0x163  :   32 - 0x20
    "00100000", --  356 - 0x164  :   32 - 0x20
    "11101011", --  357 - 0x165  :  235 - 0xeb
    "10001000", --  358 - 0x166  :  136 - 0x88
    "11010100", --  359 - 0x167  :  212 - 0xd4
    "11010101", --  360 - 0x168  :  213 - 0xd5
    "11010110", --  361 - 0x169  :  214 - 0xd6
    "11010111", --  362 - 0x16a  :  215 - 0xd7
    "11011000", --  363 - 0x16b  :  216 - 0xd8
    "11011001", --  364 - 0x16c  :  217 - 0xd9
    "11011010", --  365 - 0x16d  :  218 - 0xda
    "11011011", --  366 - 0x16e  :  219 - 0xdb
    "10001000", --  367 - 0x16f  :  136 - 0x88
    "10001000", --  368 - 0x170  :  136 - 0x88
    "11011100", --  369 - 0x171  :  220 - 0xdc
    "11010111", --  370 - 0x172  :  215 - 0xd7
    "11011101", --  371 - 0x173  :  221 - 0xdd
    "11011110", --  372 - 0x174  :  222 - 0xde
    "11011111", --  373 - 0x175  :  223 - 0xdf
    "11100000", --  374 - 0x176  :  224 - 0xe0
    "11100001", --  375 - 0x177  :  225 - 0xe1
    "11100010", --  376 - 0x178  :  226 - 0xe2
    "11100011", --  377 - 0x179  :  227 - 0xe3
    "10100011", --  378 - 0x17a  :  163 - 0xa3
    "11101001", --  379 - 0x17b  :  233 - 0xe9
    "00100000", --  380 - 0x17c  :   32 - 0x20
    "00100000", --  381 - 0x17d  :   32 - 0x20
    "00100000", --  382 - 0x17e  :   32 - 0x20
    "00100000", --  383 - 0x17f  :   32 - 0x20
    "00100000", --  384 - 0x180  :   32 - 0x20 -- line 0xc
    "00100000", --  385 - 0x181  :   32 - 0x20
    "00100000", --  386 - 0x182  :   32 - 0x20
    "00100000", --  387 - 0x183  :   32 - 0x20
    "00100000", --  388 - 0x184  :   32 - 0x20
    "11100111", --  389 - 0x185  :  231 - 0xe7
    "11101010", --  390 - 0x186  :  234 - 0xea
    "11101010", --  391 - 0x187  :  234 - 0xea
    "11101010", --  392 - 0x188  :  234 - 0xea
    "11101010", --  393 - 0x189  :  234 - 0xea
    "11101010", --  394 - 0x18a  :  234 - 0xea
    "11101010", --  395 - 0x18b  :  234 - 0xea
    "11101010", --  396 - 0x18c  :  234 - 0xea
    "11101010", --  397 - 0x18d  :  234 - 0xea
    "11101010", --  398 - 0x18e  :  234 - 0xea
    "11101010", --  399 - 0x18f  :  234 - 0xea
    "11101010", --  400 - 0x190  :  234 - 0xea
    "11101010", --  401 - 0x191  :  234 - 0xea
    "11101010", --  402 - 0x192  :  234 - 0xea
    "11101010", --  403 - 0x193  :  234 - 0xea
    "11101010", --  404 - 0x194  :  234 - 0xea
    "11101010", --  405 - 0x195  :  234 - 0xea
    "11101010", --  406 - 0x196  :  234 - 0xea
    "11101010", --  407 - 0x197  :  234 - 0xea
    "11101010", --  408 - 0x198  :  234 - 0xea
    "11101010", --  409 - 0x199  :  234 - 0xea
    "11101010", --  410 - 0x19a  :  234 - 0xea
    "11100110", --  411 - 0x19b  :  230 - 0xe6
    "00100000", --  412 - 0x19c  :   32 - 0x20
    "00100000", --  413 - 0x19d  :   32 - 0x20
    "00100000", --  414 - 0x19e  :   32 - 0x20
    "00100000", --  415 - 0x19f  :   32 - 0x20
    "00100000", --  416 - 0x1a0  :   32 - 0x20 -- line 0xd
    "00100000", --  417 - 0x1a1  :   32 - 0x20
    "00100000", --  418 - 0x1a2  :   32 - 0x20
    "00100000", --  419 - 0x1a3  :   32 - 0x20
    "00100000", --  420 - 0x1a4  :   32 - 0x20
    "00100000", --  421 - 0x1a5  :   32 - 0x20
    "00100000", --  422 - 0x1a6  :   32 - 0x20
    "00100000", --  423 - 0x1a7  :   32 - 0x20
    "00100000", --  424 - 0x1a8  :   32 - 0x20
    "00100000", --  425 - 0x1a9  :   32 - 0x20
    "00100000", --  426 - 0x1aa  :   32 - 0x20
    "00100000", --  427 - 0x1ab  :   32 - 0x20
    "00100000", --  428 - 0x1ac  :   32 - 0x20
    "00100000", --  429 - 0x1ad  :   32 - 0x20
    "00100000", --  430 - 0x1ae  :   32 - 0x20
    "00100000", --  431 - 0x1af  :   32 - 0x20
    "00100000", --  432 - 0x1b0  :   32 - 0x20
    "00100000", --  433 - 0x1b1  :   32 - 0x20
    "00100000", --  434 - 0x1b2  :   32 - 0x20
    "00100000", --  435 - 0x1b3  :   32 - 0x20
    "00100000", --  436 - 0x1b4  :   32 - 0x20
    "00100000", --  437 - 0x1b5  :   32 - 0x20
    "00100000", --  438 - 0x1b6  :   32 - 0x20
    "00100000", --  439 - 0x1b7  :   32 - 0x20
    "00100000", --  440 - 0x1b8  :   32 - 0x20
    "00100000", --  441 - 0x1b9  :   32 - 0x20
    "00100000", --  442 - 0x1ba  :   32 - 0x20
    "00100000", --  443 - 0x1bb  :   32 - 0x20
    "00100000", --  444 - 0x1bc  :   32 - 0x20
    "00100000", --  445 - 0x1bd  :   32 - 0x20
    "00100000", --  446 - 0x1be  :   32 - 0x20
    "00100000", --  447 - 0x1bf  :   32 - 0x20
    "00100000", --  448 - 0x1c0  :   32 - 0x20 -- line 0xe
    "00100000", --  449 - 0x1c1  :   32 - 0x20
    "00100000", --  450 - 0x1c2  :   32 - 0x20
    "00100000", --  451 - 0x1c3  :   32 - 0x20
    "00100000", --  452 - 0x1c4  :   32 - 0x20
    "00100000", --  453 - 0x1c5  :   32 - 0x20
    "00100000", --  454 - 0x1c6  :   32 - 0x20
    "00100000", --  455 - 0x1c7  :   32 - 0x20
    "00100000", --  456 - 0x1c8  :   32 - 0x20
    "00100000", --  457 - 0x1c9  :   32 - 0x20
    "00100000", --  458 - 0x1ca  :   32 - 0x20
    "00100000", --  459 - 0x1cb  :   32 - 0x20
    "00100000", --  460 - 0x1cc  :   32 - 0x20
    "00100000", --  461 - 0x1cd  :   32 - 0x20
    "00100000", --  462 - 0x1ce  :   32 - 0x20
    "00100000", --  463 - 0x1cf  :   32 - 0x20
    "00100000", --  464 - 0x1d0  :   32 - 0x20
    "00100000", --  465 - 0x1d1  :   32 - 0x20
    "00100000", --  466 - 0x1d2  :   32 - 0x20
    "00100000", --  467 - 0x1d3  :   32 - 0x20
    "00100000", --  468 - 0x1d4  :   32 - 0x20
    "00100000", --  469 - 0x1d5  :   32 - 0x20
    "00100000", --  470 - 0x1d6  :   32 - 0x20
    "00100000", --  471 - 0x1d7  :   32 - 0x20
    "00100000", --  472 - 0x1d8  :   32 - 0x20
    "00100000", --  473 - 0x1d9  :   32 - 0x20
    "00100000", --  474 - 0x1da  :   32 - 0x20
    "00100000", --  475 - 0x1db  :   32 - 0x20
    "00100000", --  476 - 0x1dc  :   32 - 0x20
    "00100000", --  477 - 0x1dd  :   32 - 0x20
    "00100000", --  478 - 0x1de  :   32 - 0x20
    "00100000", --  479 - 0x1df  :   32 - 0x20
    "00100000", --  480 - 0x1e0  :   32 - 0x20 -- line 0xf
    "00100000", --  481 - 0x1e1  :   32 - 0x20
    "00100000", --  482 - 0x1e2  :   32 - 0x20
    "00100000", --  483 - 0x1e3  :   32 - 0x20
    "00100000", --  484 - 0x1e4  :   32 - 0x20
    "00100000", --  485 - 0x1e5  :   32 - 0x20
    "00100000", --  486 - 0x1e6  :   32 - 0x20
    "00100000", --  487 - 0x1e7  :   32 - 0x20
    "00100000", --  488 - 0x1e8  :   32 - 0x20
    "00100000", --  489 - 0x1e9  :   32 - 0x20
    "00100000", --  490 - 0x1ea  :   32 - 0x20
    "00100000", --  491 - 0x1eb  :   32 - 0x20
    "00100000", --  492 - 0x1ec  :   32 - 0x20
    "00100000", --  493 - 0x1ed  :   32 - 0x20
    "00100000", --  494 - 0x1ee  :   32 - 0x20
    "00100000", --  495 - 0x1ef  :   32 - 0x20
    "00100000", --  496 - 0x1f0  :   32 - 0x20
    "00100000", --  497 - 0x1f1  :   32 - 0x20
    "00100000", --  498 - 0x1f2  :   32 - 0x20
    "00100000", --  499 - 0x1f3  :   32 - 0x20
    "00100000", --  500 - 0x1f4  :   32 - 0x20
    "00100000", --  501 - 0x1f5  :   32 - 0x20
    "00100000", --  502 - 0x1f6  :   32 - 0x20
    "00100000", --  503 - 0x1f7  :   32 - 0x20
    "00100000", --  504 - 0x1f8  :   32 - 0x20
    "00100000", --  505 - 0x1f9  :   32 - 0x20
    "00100000", --  506 - 0x1fa  :   32 - 0x20
    "00100000", --  507 - 0x1fb  :   32 - 0x20
    "00100000", --  508 - 0x1fc  :   32 - 0x20
    "00100000", --  509 - 0x1fd  :   32 - 0x20
    "00100000", --  510 - 0x1fe  :   32 - 0x20
    "00100000", --  511 - 0x1ff  :   32 - 0x20
    "00100000", --  512 - 0x200  :   32 - 0x20 -- line 0x10
    "00100000", --  513 - 0x201  :   32 - 0x20
    "00100000", --  514 - 0x202  :   32 - 0x20
    "00100000", --  515 - 0x203  :   32 - 0x20
    "00100000", --  516 - 0x204  :   32 - 0x20
    "00100000", --  517 - 0x205  :   32 - 0x20
    "00100000", --  518 - 0x206  :   32 - 0x20
    "00100000", --  519 - 0x207  :   32 - 0x20
    "00100000", --  520 - 0x208  :   32 - 0x20
    "00100000", --  521 - 0x209  :   32 - 0x20
    "01011100", --  522 - 0x20a  :   92 - 0x5c
    "00100000", --  523 - 0x20b  :   32 - 0x20
    "00110001", --  524 - 0x20c  :   49 - 0x31
    "00100000", --  525 - 0x20d  :   32 - 0x20
    "01010000", --  526 - 0x20e  :   80 - 0x50
    "01001100", --  527 - 0x20f  :   76 - 0x4c
    "01000001", --  528 - 0x210  :   65 - 0x41
    "01011001", --  529 - 0x211  :   89 - 0x59
    "01000101", --  530 - 0x212  :   69 - 0x45
    "01010010", --  531 - 0x213  :   82 - 0x52
    "00100000", --  532 - 0x214  :   32 - 0x20
    "00100000", --  533 - 0x215  :   32 - 0x20
    "00100000", --  534 - 0x216  :   32 - 0x20
    "00100000", --  535 - 0x217  :   32 - 0x20
    "00100000", --  536 - 0x218  :   32 - 0x20
    "00100000", --  537 - 0x219  :   32 - 0x20
    "00100000", --  538 - 0x21a  :   32 - 0x20
    "00100000", --  539 - 0x21b  :   32 - 0x20
    "00100000", --  540 - 0x21c  :   32 - 0x20
    "00100000", --  541 - 0x21d  :   32 - 0x20
    "00100000", --  542 - 0x21e  :   32 - 0x20
    "00100000", --  543 - 0x21f  :   32 - 0x20
    "00100000", --  544 - 0x220  :   32 - 0x20 -- line 0x11
    "00100000", --  545 - 0x221  :   32 - 0x20
    "00100000", --  546 - 0x222  :   32 - 0x20
    "00100000", --  547 - 0x223  :   32 - 0x20
    "00100000", --  548 - 0x224  :   32 - 0x20
    "00100000", --  549 - 0x225  :   32 - 0x20
    "00100000", --  550 - 0x226  :   32 - 0x20
    "00100000", --  551 - 0x227  :   32 - 0x20
    "00100000", --  552 - 0x228  :   32 - 0x20
    "00100000", --  553 - 0x229  :   32 - 0x20
    "00100000", --  554 - 0x22a  :   32 - 0x20
    "00100000", --  555 - 0x22b  :   32 - 0x20
    "00100000", --  556 - 0x22c  :   32 - 0x20
    "00100000", --  557 - 0x22d  :   32 - 0x20
    "00100000", --  558 - 0x22e  :   32 - 0x20
    "00100000", --  559 - 0x22f  :   32 - 0x20
    "00100000", --  560 - 0x230  :   32 - 0x20
    "00100000", --  561 - 0x231  :   32 - 0x20
    "00100000", --  562 - 0x232  :   32 - 0x20
    "00100000", --  563 - 0x233  :   32 - 0x20
    "00100000", --  564 - 0x234  :   32 - 0x20
    "00100000", --  565 - 0x235  :   32 - 0x20
    "00100000", --  566 - 0x236  :   32 - 0x20
    "00100000", --  567 - 0x237  :   32 - 0x20
    "00100000", --  568 - 0x238  :   32 - 0x20
    "00100000", --  569 - 0x239  :   32 - 0x20
    "00100000", --  570 - 0x23a  :   32 - 0x20
    "00100000", --  571 - 0x23b  :   32 - 0x20
    "00100000", --  572 - 0x23c  :   32 - 0x20
    "00100000", --  573 - 0x23d  :   32 - 0x20
    "00100000", --  574 - 0x23e  :   32 - 0x20
    "00100000", --  575 - 0x23f  :   32 - 0x20
    "00100000", --  576 - 0x240  :   32 - 0x20 -- line 0x12
    "00100000", --  577 - 0x241  :   32 - 0x20
    "00100000", --  578 - 0x242  :   32 - 0x20
    "00100000", --  579 - 0x243  :   32 - 0x20
    "00100000", --  580 - 0x244  :   32 - 0x20
    "00100000", --  581 - 0x245  :   32 - 0x20
    "00100000", --  582 - 0x246  :   32 - 0x20
    "00100000", --  583 - 0x247  :   32 - 0x20
    "00100000", --  584 - 0x248  :   32 - 0x20
    "00100000", --  585 - 0x249  :   32 - 0x20
    "00100000", --  586 - 0x24a  :   32 - 0x20
    "00100000", --  587 - 0x24b  :   32 - 0x20
    "00110010", --  588 - 0x24c  :   50 - 0x32
    "00100000", --  589 - 0x24d  :   32 - 0x20
    "01010000", --  590 - 0x24e  :   80 - 0x50
    "01001100", --  591 - 0x24f  :   76 - 0x4c
    "01000001", --  592 - 0x250  :   65 - 0x41
    "01011001", --  593 - 0x251  :   89 - 0x59
    "01000101", --  594 - 0x252  :   69 - 0x45
    "01010010", --  595 - 0x253  :   82 - 0x52
    "01010011", --  596 - 0x254  :   83 - 0x53
    "00100000", --  597 - 0x255  :   32 - 0x20
    "00100000", --  598 - 0x256  :   32 - 0x20
    "00100000", --  599 - 0x257  :   32 - 0x20
    "00100000", --  600 - 0x258  :   32 - 0x20
    "00100000", --  601 - 0x259  :   32 - 0x20
    "00100000", --  602 - 0x25a  :   32 - 0x20
    "00100000", --  603 - 0x25b  :   32 - 0x20
    "00100000", --  604 - 0x25c  :   32 - 0x20
    "00100000", --  605 - 0x25d  :   32 - 0x20
    "00100000", --  606 - 0x25e  :   32 - 0x20
    "00100000", --  607 - 0x25f  :   32 - 0x20
    "00100000", --  608 - 0x260  :   32 - 0x20 -- line 0x13
    "00100000", --  609 - 0x261  :   32 - 0x20
    "00100000", --  610 - 0x262  :   32 - 0x20
    "00100000", --  611 - 0x263  :   32 - 0x20
    "00100000", --  612 - 0x264  :   32 - 0x20
    "00100000", --  613 - 0x265  :   32 - 0x20
    "00100000", --  614 - 0x266  :   32 - 0x20
    "00100000", --  615 - 0x267  :   32 - 0x20
    "00100000", --  616 - 0x268  :   32 - 0x20
    "00100000", --  617 - 0x269  :   32 - 0x20
    "00100000", --  618 - 0x26a  :   32 - 0x20
    "00100000", --  619 - 0x26b  :   32 - 0x20
    "00100000", --  620 - 0x26c  :   32 - 0x20
    "00100000", --  621 - 0x26d  :   32 - 0x20
    "00100000", --  622 - 0x26e  :   32 - 0x20
    "00100000", --  623 - 0x26f  :   32 - 0x20
    "00100000", --  624 - 0x270  :   32 - 0x20
    "00100000", --  625 - 0x271  :   32 - 0x20
    "00100000", --  626 - 0x272  :   32 - 0x20
    "00100000", --  627 - 0x273  :   32 - 0x20
    "00100000", --  628 - 0x274  :   32 - 0x20
    "00100000", --  629 - 0x275  :   32 - 0x20
    "00100000", --  630 - 0x276  :   32 - 0x20
    "00100000", --  631 - 0x277  :   32 - 0x20
    "00100000", --  632 - 0x278  :   32 - 0x20
    "00100000", --  633 - 0x279  :   32 - 0x20
    "00100000", --  634 - 0x27a  :   32 - 0x20
    "00100000", --  635 - 0x27b  :   32 - 0x20
    "00100000", --  636 - 0x27c  :   32 - 0x20
    "00100000", --  637 - 0x27d  :   32 - 0x20
    "00100000", --  638 - 0x27e  :   32 - 0x20
    "00100000", --  639 - 0x27f  :   32 - 0x20
    "00100000", --  640 - 0x280  :   32 - 0x20 -- line 0x14
    "00100000", --  641 - 0x281  :   32 - 0x20
    "00100000", --  642 - 0x282  :   32 - 0x20
    "00100000", --  643 - 0x283  :   32 - 0x20
    "00100000", --  644 - 0x284  :   32 - 0x20
    "00100000", --  645 - 0x285  :   32 - 0x20
    "00100000", --  646 - 0x286  :   32 - 0x20
    "00100000", --  647 - 0x287  :   32 - 0x20
    "00100000", --  648 - 0x288  :   32 - 0x20
    "00100000", --  649 - 0x289  :   32 - 0x20
    "00100000", --  650 - 0x28a  :   32 - 0x20
    "00100000", --  651 - 0x28b  :   32 - 0x20
    "00100000", --  652 - 0x28c  :   32 - 0x20
    "00100000", --  653 - 0x28d  :   32 - 0x20
    "00100000", --  654 - 0x28e  :   32 - 0x20
    "00100000", --  655 - 0x28f  :   32 - 0x20
    "00100000", --  656 - 0x290  :   32 - 0x20
    "00100000", --  657 - 0x291  :   32 - 0x20
    "00100000", --  658 - 0x292  :   32 - 0x20
    "00100000", --  659 - 0x293  :   32 - 0x20
    "00100000", --  660 - 0x294  :   32 - 0x20
    "00100000", --  661 - 0x295  :   32 - 0x20
    "00100000", --  662 - 0x296  :   32 - 0x20
    "00100000", --  663 - 0x297  :   32 - 0x20
    "00100000", --  664 - 0x298  :   32 - 0x20
    "00100000", --  665 - 0x299  :   32 - 0x20
    "00100000", --  666 - 0x29a  :   32 - 0x20
    "00100000", --  667 - 0x29b  :   32 - 0x20
    "00100000", --  668 - 0x29c  :   32 - 0x20
    "00100000", --  669 - 0x29d  :   32 - 0x20
    "00100000", --  670 - 0x29e  :   32 - 0x20
    "00100000", --  671 - 0x29f  :   32 - 0x20
    "00100000", --  672 - 0x2a0  :   32 - 0x20 -- line 0x15
    "00100000", --  673 - 0x2a1  :   32 - 0x20
    "01010100", --  674 - 0x2a2  :   84 - 0x54
    "01001101", --  675 - 0x2a3  :   77 - 0x4d
    "00100000", --  676 - 0x2a4  :   32 - 0x20
    "01000001", --  677 - 0x2a5  :   65 - 0x41
    "01001110", --  678 - 0x2a6  :   78 - 0x4e
    "01000100", --  679 - 0x2a7  :   68 - 0x44
    "00100000", --  680 - 0x2a8  :   32 - 0x20
    "01011101", --  681 - 0x2a9  :   93 - 0x5d
    "00100000", --  682 - 0x2aa  :   32 - 0x20
    "00110001", --  683 - 0x2ab  :   49 - 0x31
    "00111001", --  684 - 0x2ac  :   57 - 0x39
    "00111000", --  685 - 0x2ad  :   56 - 0x38
    "00110000", --  686 - 0x2ae  :   48 - 0x30
    "00100000", --  687 - 0x2af  :   32 - 0x20
    "00110001", --  688 - 0x2b0  :   49 - 0x31
    "00111001", --  689 - 0x2b1  :   57 - 0x39
    "00111000", --  690 - 0x2b2  :   56 - 0x38
    "00110100", --  691 - 0x2b3  :   52 - 0x34
    "00100000", --  692 - 0x2b4  :   32 - 0x20
    "01001110", --  693 - 0x2b5  :   78 - 0x4e
    "01000001", --  694 - 0x2b6  :   65 - 0x41
    "01001101", --  695 - 0x2b7  :   77 - 0x4d
    "01000011", --  696 - 0x2b8  :   67 - 0x43
    "01001111", --  697 - 0x2b9  :   79 - 0x4f
    "00100000", --  698 - 0x2ba  :   32 - 0x20
    "01001100", --  699 - 0x2bb  :   76 - 0x4c
    "01010100", --  700 - 0x2bc  :   84 - 0x54
    "01000100", --  701 - 0x2bd  :   68 - 0x44
    "01011011", --  702 - 0x2be  :   91 - 0x5b
    "00100000", --  703 - 0x2bf  :   32 - 0x20
    "00100000", --  704 - 0x2c0  :   32 - 0x20 -- line 0x16
    "00100000", --  705 - 0x2c1  :   32 - 0x20
    "00100000", --  706 - 0x2c2  :   32 - 0x20
    "00100000", --  707 - 0x2c3  :   32 - 0x20
    "00100000", --  708 - 0x2c4  :   32 - 0x20
    "00100000", --  709 - 0x2c5  :   32 - 0x20
    "00100000", --  710 - 0x2c6  :   32 - 0x20
    "00100000", --  711 - 0x2c7  :   32 - 0x20
    "00100000", --  712 - 0x2c8  :   32 - 0x20
    "00100000", --  713 - 0x2c9  :   32 - 0x20
    "00100000", --  714 - 0x2ca  :   32 - 0x20
    "00100000", --  715 - 0x2cb  :   32 - 0x20
    "00100000", --  716 - 0x2cc  :   32 - 0x20
    "00100000", --  717 - 0x2cd  :   32 - 0x20
    "00100000", --  718 - 0x2ce  :   32 - 0x20
    "00100000", --  719 - 0x2cf  :   32 - 0x20
    "00100000", --  720 - 0x2d0  :   32 - 0x20
    "00100000", --  721 - 0x2d1  :   32 - 0x20
    "00100000", --  722 - 0x2d2  :   32 - 0x20
    "00100000", --  723 - 0x2d3  :   32 - 0x20
    "00100000", --  724 - 0x2d4  :   32 - 0x20
    "00100000", --  725 - 0x2d5  :   32 - 0x20
    "00100000", --  726 - 0x2d6  :   32 - 0x20
    "00100000", --  727 - 0x2d7  :   32 - 0x20
    "00100000", --  728 - 0x2d8  :   32 - 0x20
    "00100000", --  729 - 0x2d9  :   32 - 0x20
    "00100000", --  730 - 0x2da  :   32 - 0x20
    "00100000", --  731 - 0x2db  :   32 - 0x20
    "00100000", --  732 - 0x2dc  :   32 - 0x20
    "00100000", --  733 - 0x2dd  :   32 - 0x20
    "00100000", --  734 - 0x2de  :   32 - 0x20
    "00100000", --  735 - 0x2df  :   32 - 0x20
    "00100000", --  736 - 0x2e0  :   32 - 0x20 -- line 0x17
    "00100000", --  737 - 0x2e1  :   32 - 0x20
    "00100000", --  738 - 0x2e2  :   32 - 0x20
    "00100000", --  739 - 0x2e3  :   32 - 0x20
    "00100000", --  740 - 0x2e4  :   32 - 0x20
    "00100000", --  741 - 0x2e5  :   32 - 0x20
    "00100000", --  742 - 0x2e6  :   32 - 0x20
    "00100000", --  743 - 0x2e7  :   32 - 0x20
    "00100000", --  744 - 0x2e8  :   32 - 0x20
    "00100000", --  745 - 0x2e9  :   32 - 0x20
    "00100000", --  746 - 0x2ea  :   32 - 0x20
    "00100000", --  747 - 0x2eb  :   32 - 0x20
    "00100000", --  748 - 0x2ec  :   32 - 0x20
    "01010100", --  749 - 0x2ed  :   84 - 0x54
    "01000101", --  750 - 0x2ee  :   69 - 0x45
    "01001110", --  751 - 0x2ef  :   78 - 0x4e
    "01000111", --  752 - 0x2f0  :   71 - 0x47
    "01000101", --  753 - 0x2f1  :   69 - 0x45
    "01001110", --  754 - 0x2f2  :   78 - 0x4e
    "00100000", --  755 - 0x2f3  :   32 - 0x20
    "00100000", --  756 - 0x2f4  :   32 - 0x20
    "00100000", --  757 - 0x2f5  :   32 - 0x20
    "00100000", --  758 - 0x2f6  :   32 - 0x20
    "00100000", --  759 - 0x2f7  :   32 - 0x20
    "00100000", --  760 - 0x2f8  :   32 - 0x20
    "00100000", --  761 - 0x2f9  :   32 - 0x20
    "00100000", --  762 - 0x2fa  :   32 - 0x20
    "00100000", --  763 - 0x2fb  :   32 - 0x20
    "00100000", --  764 - 0x2fc  :   32 - 0x20
    "00100000", --  765 - 0x2fd  :   32 - 0x20
    "00100000", --  766 - 0x2fe  :   32 - 0x20
    "00100000", --  767 - 0x2ff  :   32 - 0x20
    "00100000", --  768 - 0x300  :   32 - 0x20 -- line 0x18
    "00100000", --  769 - 0x301  :   32 - 0x20
    "00100000", --  770 - 0x302  :   32 - 0x20
    "00100000", --  771 - 0x303  :   32 - 0x20
    "00100000", --  772 - 0x304  :   32 - 0x20
    "00100000", --  773 - 0x305  :   32 - 0x20
    "00100000", --  774 - 0x306  :   32 - 0x20
    "00100000", --  775 - 0x307  :   32 - 0x20
    "00100000", --  776 - 0x308  :   32 - 0x20
    "00100000", --  777 - 0x309  :   32 - 0x20
    "00100000", --  778 - 0x30a  :   32 - 0x20
    "00100000", --  779 - 0x30b  :   32 - 0x20
    "00100000", --  780 - 0x30c  :   32 - 0x20
    "00100000", --  781 - 0x30d  :   32 - 0x20
    "00100000", --  782 - 0x30e  :   32 - 0x20
    "00100000", --  783 - 0x30f  :   32 - 0x20
    "00100000", --  784 - 0x310  :   32 - 0x20
    "00100000", --  785 - 0x311  :   32 - 0x20
    "00100000", --  786 - 0x312  :   32 - 0x20
    "00100000", --  787 - 0x313  :   32 - 0x20
    "00100000", --  788 - 0x314  :   32 - 0x20
    "00100000", --  789 - 0x315  :   32 - 0x20
    "00100000", --  790 - 0x316  :   32 - 0x20
    "00100000", --  791 - 0x317  :   32 - 0x20
    "00100000", --  792 - 0x318  :   32 - 0x20
    "00100000", --  793 - 0x319  :   32 - 0x20
    "00100000", --  794 - 0x31a  :   32 - 0x20
    "00100000", --  795 - 0x31b  :   32 - 0x20
    "00100000", --  796 - 0x31c  :   32 - 0x20
    "00100000", --  797 - 0x31d  :   32 - 0x20
    "00100000", --  798 - 0x31e  :   32 - 0x20
    "00100000", --  799 - 0x31f  :   32 - 0x20
    "00100000", --  800 - 0x320  :   32 - 0x20 -- line 0x19
    "00100000", --  801 - 0x321  :   32 - 0x20
    "00100000", --  802 - 0x322  :   32 - 0x20
    "00100000", --  803 - 0x323  :   32 - 0x20
    "00100000", --  804 - 0x324  :   32 - 0x20
    "00100000", --  805 - 0x325  :   32 - 0x20
    "00100000", --  806 - 0x326  :   32 - 0x20
    "00100000", --  807 - 0x327  :   32 - 0x20
    "00100000", --  808 - 0x328  :   32 - 0x20
    "00100000", --  809 - 0x329  :   32 - 0x20
    "00100000", --  810 - 0x32a  :   32 - 0x20
    "00100000", --  811 - 0x32b  :   32 - 0x20
    "00100000", --  812 - 0x32c  :   32 - 0x20
    "00100000", --  813 - 0x32d  :   32 - 0x20
    "00100000", --  814 - 0x32e  :   32 - 0x20
    "00100000", --  815 - 0x32f  :   32 - 0x20
    "00100000", --  816 - 0x330  :   32 - 0x20
    "00100000", --  817 - 0x331  :   32 - 0x20
    "00100000", --  818 - 0x332  :   32 - 0x20
    "00100000", --  819 - 0x333  :   32 - 0x20
    "00100000", --  820 - 0x334  :   32 - 0x20
    "00100000", --  821 - 0x335  :   32 - 0x20
    "00100000", --  822 - 0x336  :   32 - 0x20
    "00100000", --  823 - 0x337  :   32 - 0x20
    "00100000", --  824 - 0x338  :   32 - 0x20
    "00100000", --  825 - 0x339  :   32 - 0x20
    "00100000", --  826 - 0x33a  :   32 - 0x20
    "00100000", --  827 - 0x33b  :   32 - 0x20
    "00100000", --  828 - 0x33c  :   32 - 0x20
    "00100000", --  829 - 0x33d  :   32 - 0x20
    "00100000", --  830 - 0x33e  :   32 - 0x20
    "00100000", --  831 - 0x33f  :   32 - 0x20
    "00100000", --  832 - 0x340  :   32 - 0x20 -- line 0x1a
    "00100000", --  833 - 0x341  :   32 - 0x20
    "00100000", --  834 - 0x342  :   32 - 0x20
    "00100000", --  835 - 0x343  :   32 - 0x20
    "00100000", --  836 - 0x344  :   32 - 0x20
    "00100000", --  837 - 0x345  :   32 - 0x20
    "00100000", --  838 - 0x346  :   32 - 0x20
    "00100000", --  839 - 0x347  :   32 - 0x20
    "00100000", --  840 - 0x348  :   32 - 0x20
    "00100000", --  841 - 0x349  :   32 - 0x20
    "00100000", --  842 - 0x34a  :   32 - 0x20
    "00100000", --  843 - 0x34b  :   32 - 0x20
    "00100000", --  844 - 0x34c  :   32 - 0x20
    "00100000", --  845 - 0x34d  :   32 - 0x20
    "00100000", --  846 - 0x34e  :   32 - 0x20
    "00100000", --  847 - 0x34f  :   32 - 0x20
    "00100000", --  848 - 0x350  :   32 - 0x20
    "00100000", --  849 - 0x351  :   32 - 0x20
    "00100000", --  850 - 0x352  :   32 - 0x20
    "00100000", --  851 - 0x353  :   32 - 0x20
    "00100000", --  852 - 0x354  :   32 - 0x20
    "00100000", --  853 - 0x355  :   32 - 0x20
    "00100000", --  854 - 0x356  :   32 - 0x20
    "00100000", --  855 - 0x357  :   32 - 0x20
    "00100000", --  856 - 0x358  :   32 - 0x20
    "00100000", --  857 - 0x359  :   32 - 0x20
    "00100000", --  858 - 0x35a  :   32 - 0x20
    "00100000", --  859 - 0x35b  :   32 - 0x20
    "00100000", --  860 - 0x35c  :   32 - 0x20
    "00100000", --  861 - 0x35d  :   32 - 0x20
    "00100000", --  862 - 0x35e  :   32 - 0x20
    "00100000", --  863 - 0x35f  :   32 - 0x20
    "00100000", --  864 - 0x360  :   32 - 0x20 -- line 0x1b
    "00100000", --  865 - 0x361  :   32 - 0x20
    "00100000", --  866 - 0x362  :   32 - 0x20
    "00100000", --  867 - 0x363  :   32 - 0x20
    "00100000", --  868 - 0x364  :   32 - 0x20
    "00100000", --  869 - 0x365  :   32 - 0x20
    "00100000", --  870 - 0x366  :   32 - 0x20
    "00100000", --  871 - 0x367  :   32 - 0x20
    "00100000", --  872 - 0x368  :   32 - 0x20
    "00100000", --  873 - 0x369  :   32 - 0x20
    "00100000", --  874 - 0x36a  :   32 - 0x20
    "00100000", --  875 - 0x36b  :   32 - 0x20
    "00100000", --  876 - 0x36c  :   32 - 0x20
    "00100000", --  877 - 0x36d  :   32 - 0x20
    "00100000", --  878 - 0x36e  :   32 - 0x20
    "00100000", --  879 - 0x36f  :   32 - 0x20
    "00100000", --  880 - 0x370  :   32 - 0x20
    "00100000", --  881 - 0x371  :   32 - 0x20
    "00100000", --  882 - 0x372  :   32 - 0x20
    "00100000", --  883 - 0x373  :   32 - 0x20
    "00100000", --  884 - 0x374  :   32 - 0x20
    "00100000", --  885 - 0x375  :   32 - 0x20
    "00100000", --  886 - 0x376  :   32 - 0x20
    "00100000", --  887 - 0x377  :   32 - 0x20
    "00100000", --  888 - 0x378  :   32 - 0x20
    "00100000", --  889 - 0x379  :   32 - 0x20
    "00100000", --  890 - 0x37a  :   32 - 0x20
    "00100000", --  891 - 0x37b  :   32 - 0x20
    "00100000", --  892 - 0x37c  :   32 - 0x20
    "00100000", --  893 - 0x37d  :   32 - 0x20
    "00100000", --  894 - 0x37e  :   32 - 0x20
    "00100000", --  895 - 0x37f  :   32 - 0x20
    "00100000", --  896 - 0x380  :   32 - 0x20 -- line 0x1c
    "00100000", --  897 - 0x381  :   32 - 0x20
    "00100000", --  898 - 0x382  :   32 - 0x20
    "00100000", --  899 - 0x383  :   32 - 0x20
    "00100000", --  900 - 0x384  :   32 - 0x20
    "00100000", --  901 - 0x385  :   32 - 0x20
    "00100000", --  902 - 0x386  :   32 - 0x20
    "00100000", --  903 - 0x387  :   32 - 0x20
    "00100000", --  904 - 0x388  :   32 - 0x20
    "00100000", --  905 - 0x389  :   32 - 0x20
    "00100000", --  906 - 0x38a  :   32 - 0x20
    "00100000", --  907 - 0x38b  :   32 - 0x20
    "00100000", --  908 - 0x38c  :   32 - 0x20
    "00100000", --  909 - 0x38d  :   32 - 0x20
    "00100000", --  910 - 0x38e  :   32 - 0x20
    "00100000", --  911 - 0x38f  :   32 - 0x20
    "00100000", --  912 - 0x390  :   32 - 0x20
    "00100000", --  913 - 0x391  :   32 - 0x20
    "00100000", --  914 - 0x392  :   32 - 0x20
    "00100000", --  915 - 0x393  :   32 - 0x20
    "00100000", --  916 - 0x394  :   32 - 0x20
    "00100000", --  917 - 0x395  :   32 - 0x20
    "00100000", --  918 - 0x396  :   32 - 0x20
    "00100000", --  919 - 0x397  :   32 - 0x20
    "00100000", --  920 - 0x398  :   32 - 0x20
    "00100000", --  921 - 0x399  :   32 - 0x20
    "00100000", --  922 - 0x39a  :   32 - 0x20
    "00100000", --  923 - 0x39b  :   32 - 0x20
    "00100000", --  924 - 0x39c  :   32 - 0x20
    "00100000", --  925 - 0x39d  :   32 - 0x20
    "00100000", --  926 - 0x39e  :   32 - 0x20
    "00100000", --  927 - 0x39f  :   32 - 0x20
    "00100000", --  928 - 0x3a0  :   32 - 0x20 -- line 0x1d
    "00100000", --  929 - 0x3a1  :   32 - 0x20
    "00100000", --  930 - 0x3a2  :   32 - 0x20
    "00100000", --  931 - 0x3a3  :   32 - 0x20
    "00100000", --  932 - 0x3a4  :   32 - 0x20
    "00100000", --  933 - 0x3a5  :   32 - 0x20
    "00100000", --  934 - 0x3a6  :   32 - 0x20
    "00100000", --  935 - 0x3a7  :   32 - 0x20
    "00100000", --  936 - 0x3a8  :   32 - 0x20
    "00100000", --  937 - 0x3a9  :   32 - 0x20
    "00100000", --  938 - 0x3aa  :   32 - 0x20
    "00100000", --  939 - 0x3ab  :   32 - 0x20
    "00100000", --  940 - 0x3ac  :   32 - 0x20
    "00100000", --  941 - 0x3ad  :   32 - 0x20
    "00100000", --  942 - 0x3ae  :   32 - 0x20
    "00100000", --  943 - 0x3af  :   32 - 0x20
    "00100000", --  944 - 0x3b0  :   32 - 0x20
    "00100000", --  945 - 0x3b1  :   32 - 0x20
    "00100000", --  946 - 0x3b2  :   32 - 0x20
    "00100000", --  947 - 0x3b3  :   32 - 0x20
    "00100000", --  948 - 0x3b4  :   32 - 0x20
    "00100000", --  949 - 0x3b5  :   32 - 0x20
    "00100000", --  950 - 0x3b6  :   32 - 0x20
    "00100000", --  951 - 0x3b7  :   32 - 0x20
    "00100000", --  952 - 0x3b8  :   32 - 0x20
    "00100000", --  953 - 0x3b9  :   32 - 0x20
    "00100000", --  954 - 0x3ba  :   32 - 0x20
    "00100000", --  955 - 0x3bb  :   32 - 0x20
    "00100000", --  956 - 0x3bc  :   32 - 0x20
    "00100000", --  957 - 0x3bd  :   32 - 0x20
    "00100000", --  958 - 0x3be  :   32 - 0x20
    "00100000", --  959 - 0x3bf  :   32 - 0x20
        ---- Attribute Table 0----
    "00000000", --  960 - 0x3c0  :    0 - 0x0
    "00000000", --  961 - 0x3c1  :    0 - 0x0
    "00000000", --  962 - 0x3c2  :    0 - 0x0
    "00000000", --  963 - 0x3c3  :    0 - 0x0
    "00000000", --  964 - 0x3c4  :    0 - 0x0
    "00000000", --  965 - 0x3c5  :    0 - 0x0
    "00000000", --  966 - 0x3c6  :    0 - 0x0
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "10000000", --  968 - 0x3c8  :  128 - 0x80
    "10100000", --  969 - 0x3c9  :  160 - 0xa0
    "10100000", --  970 - 0x3ca  :  160 - 0xa0
    "10100000", --  971 - 0x3cb  :  160 - 0xa0
    "10100000", --  972 - 0x3cc  :  160 - 0xa0
    "10100000", --  973 - 0x3cd  :  160 - 0xa0
    "10100000", --  974 - 0x3ce  :  160 - 0xa0
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "00000000", --  976 - 0x3d0  :    0 - 0x0
    "01100110", --  977 - 0x3d1  :  102 - 0x66
    "01010101", --  978 - 0x3d2  :   85 - 0x55
    "01010101", --  979 - 0x3d3  :   85 - 0x55
    "01010101", --  980 - 0x3d4  :   85 - 0x55
    "01010101", --  981 - 0x3d5  :   85 - 0x55
    "11011101", --  982 - 0x3d6  :  221 - 0xdd
    "00000000", --  983 - 0x3d7  :    0 - 0x0
    "00001000", --  984 - 0x3d8  :    8 - 0x8
    "00001010", --  985 - 0x3d9  :   10 - 0xa
    "00001010", --  986 - 0x3da  :   10 - 0xa
    "00001010", --  987 - 0x3db  :   10 - 0xa
    "00001010", --  988 - 0x3dc  :   10 - 0xa
    "00001010", --  989 - 0x3dd  :   10 - 0xa
    "00001010", --  990 - 0x3de  :   10 - 0xa
    "00000000", --  991 - 0x3df  :    0 - 0x0
    "00000000", --  992 - 0x3e0  :    0 - 0x0
    "00000000", --  993 - 0x3e1  :    0 - 0x0
    "00000000", --  994 - 0x3e2  :    0 - 0x0
    "00000000", --  995 - 0x3e3  :    0 - 0x0
    "00000000", --  996 - 0x3e4  :    0 - 0x0
    "00000000", --  997 - 0x3e5  :    0 - 0x0
    "00000000", --  998 - 0x3e6  :    0 - 0x0
    "00000000", --  999 - 0x3e7  :    0 - 0x0
    "11110000", -- 1000 - 0x3e8  :  240 - 0xf0
    "11110000", -- 1001 - 0x3e9  :  240 - 0xf0
    "11110000", -- 1002 - 0x3ea  :  240 - 0xf0
    "11110000", -- 1003 - 0x3eb  :  240 - 0xf0
    "11110000", -- 1004 - 0x3ec  :  240 - 0xf0
    "11110000", -- 1005 - 0x3ed  :  240 - 0xf0
    "11110000", -- 1006 - 0x3ee  :  240 - 0xf0
    "11110000", -- 1007 - 0x3ef  :  240 - 0xf0
    "00000000", -- 1008 - 0x3f0  :    0 - 0x0
    "00000000", -- 1009 - 0x3f1  :    0 - 0x0
    "00000000", -- 1010 - 0x3f2  :    0 - 0x0
    "00000000", -- 1011 - 0x3f3  :    0 - 0x0
    "00000000", -- 1012 - 0x3f4  :    0 - 0x0
    "00000000", -- 1013 - 0x3f5  :    0 - 0x0
    "00000000", -- 1014 - 0x3f6  :    0 - 0x0
    "00000000", -- 1015 - 0x3f7  :    0 - 0x0
    "00000000", -- 1016 - 0x3f8  :    0 - 0x0
    "00000000", -- 1017 - 0x3f9  :    0 - 0x0
    "00000000", -- 1018 - 0x3fa  :    0 - 0x0
    "00000000", -- 1019 - 0x3fb  :    0 - 0x0
    "00000000", -- 1020 - 0x3fc  :    0 - 0x0
    "00000000", -- 1021 - 0x3fd  :    0 - 0x0
    "00000000", -- 1022 - 0x3fe  :    0 - 0x0
    "00000000"  -- 1023 - 0x3ff  :    0 - 0x0
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
