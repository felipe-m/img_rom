//- Autcmatically generated verilog ROM from a NES memory file----
//-   PATTERN TABLE WITH ONLY ONE COLOR PLANE
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


//-  Original memory dump file name: smario_traspas_patron.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_PTABLE_SPRILO_color1
  (
     //input     clk,   // clock
     input      [12-1:0] addr,  //4096 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                              //  address:   value 
                              //    dec  : dec - hex
          // Sprite pattern Table
      12'h0: dout  = 8'b00000000; //    0 :   0 - 0x0 -- Sprite 0x0
      12'h1: dout  = 8'b00000000; //    1 :   0 - 0x0
      12'h2: dout  = 8'b00000000; //    2 :   0 - 0x0
      12'h3: dout  = 8'b00000000; //    3 :   0 - 0x0
      12'h4: dout  = 8'b00011111; //    4 :  31 - 0x1f
      12'h5: dout  = 8'b00111111; //    5 :  63 - 0x3f
      12'h6: dout  = 8'b00111111; //    6 :  63 - 0x3f
      12'h7: dout  = 8'b01111111; //    7 : 127 - 0x7f
      12'h8: dout  = 8'b00000000; //    8 :   0 - 0x0 -- Sprite 0x1
      12'h9: dout  = 8'b00100000; //    9 :  32 - 0x20
      12'hA: dout  = 8'b01100000; //   10 :  96 - 0x60
      12'hB: dout  = 8'b00000000; //   11 :   0 - 0x0
      12'hC: dout  = 8'b11110000; //   12 : 240 - 0xf0
      12'hD: dout  = 8'b11111100; //   13 : 252 - 0xfc
      12'hE: dout  = 8'b11111110; //   14 : 254 - 0xfe
      12'hF: dout  = 8'b11111110; //   15 : 254 - 0xfe
      12'h10: dout  = 8'b01111111; //   16 : 127 - 0x7f -- Sprite 0x2
      12'h11: dout  = 8'b01111111; //   17 : 127 - 0x7f
      12'h12: dout  = 8'b00011111; //   18 :  31 - 0x1f
      12'h13: dout  = 8'b00000111; //   19 :   7 - 0x7
      12'h14: dout  = 8'b00000000; //   20 :   0 - 0x0
      12'h15: dout  = 8'b00011110; //   21 :  30 - 0x1e
      12'h16: dout  = 8'b00111111; //   22 :  63 - 0x3f
      12'h17: dout  = 8'b01111111; //   23 : 127 - 0x7f
      12'h18: dout  = 8'b11111100; //   24 : 252 - 0xfc -- Sprite 0x3
      12'h19: dout  = 8'b11111100; //   25 : 252 - 0xfc
      12'h1A: dout  = 8'b11111000; //   26 : 248 - 0xf8
      12'h1B: dout  = 8'b11000000; //   27 : 192 - 0xc0
      12'h1C: dout  = 8'b11000010; //   28 : 194 - 0xc2
      12'h1D: dout  = 8'b01100111; //   29 : 103 - 0x67
      12'h1E: dout  = 8'b00101111; //   30 :  47 - 0x2f
      12'h1F: dout  = 8'b00110111; //   31 :  55 - 0x37
      12'h20: dout  = 8'b01111111; //   32 : 127 - 0x7f -- Sprite 0x4
      12'h21: dout  = 8'b01111110; //   33 : 126 - 0x7e
      12'h22: dout  = 8'b11111100; //   34 : 252 - 0xfc
      12'h23: dout  = 8'b11110000; //   35 : 240 - 0xf0
      12'h24: dout  = 8'b11111000; //   36 : 248 - 0xf8
      12'h25: dout  = 8'b11111000; //   37 : 248 - 0xf8
      12'h26: dout  = 8'b11110000; //   38 : 240 - 0xf0
      12'h27: dout  = 8'b01110000; //   39 : 112 - 0x70
      12'h28: dout  = 8'b00110111; //   40 :  55 - 0x37 -- Sprite 0x5
      12'h29: dout  = 8'b00110110; //   41 :  54 - 0x36
      12'h2A: dout  = 8'b01011100; //   42 :  92 - 0x5c
      12'h2B: dout  = 8'b00000000; //   43 :   0 - 0x0
      12'h2C: dout  = 8'b00000000; //   44 :   0 - 0x0
      12'h2D: dout  = 8'b00000001; //   45 :   1 - 0x1
      12'h2E: dout  = 8'b00000011; //   46 :   3 - 0x3
      12'h2F: dout  = 8'b00011111; //   47 :  31 - 0x1f
      12'h30: dout  = 8'b00001000; //   48 :   8 - 0x8 -- Sprite 0x6
      12'h31: dout  = 8'b00100100; //   49 :  36 - 0x24
      12'h32: dout  = 8'b11100011; //   50 : 227 - 0xe3
      12'h33: dout  = 8'b11110000; //   51 : 240 - 0xf0
      12'h34: dout  = 8'b11111000; //   52 : 248 - 0xf8
      12'h35: dout  = 8'b01110000; //   53 : 112 - 0x70
      12'h36: dout  = 8'b01110000; //   54 : 112 - 0x70
      12'h37: dout  = 8'b00111000; //   55 :  56 - 0x38
      12'h38: dout  = 8'b00011111; //   56 :  31 - 0x1f -- Sprite 0x7
      12'h39: dout  = 8'b00011111; //   57 :  31 - 0x1f
      12'h3A: dout  = 8'b00011111; //   58 :  31 - 0x1f
      12'h3B: dout  = 8'b00011111; //   59 :  31 - 0x1f
      12'h3C: dout  = 8'b00000000; //   60 :   0 - 0x0
      12'h3D: dout  = 8'b00000000; //   61 :   0 - 0x0
      12'h3E: dout  = 8'b00000000; //   62 :   0 - 0x0
      12'h3F: dout  = 8'b00000000; //   63 :   0 - 0x0
      12'h40: dout  = 8'b00000000; //   64 :   0 - 0x0 -- Sprite 0x8
      12'h41: dout  = 8'b00000000; //   65 :   0 - 0x0
      12'h42: dout  = 8'b00000000; //   66 :   0 - 0x0
      12'h43: dout  = 8'b00000000; //   67 :   0 - 0x0
      12'h44: dout  = 8'b00000000; //   68 :   0 - 0x0
      12'h45: dout  = 8'b00000000; //   69 :   0 - 0x0
      12'h46: dout  = 8'b00001111; //   70 :  15 - 0xf
      12'h47: dout  = 8'b00011111; //   71 :  31 - 0x1f
      12'h48: dout  = 8'b00000000; //   72 :   0 - 0x0 -- Sprite 0x9
      12'h49: dout  = 8'b00000000; //   73 :   0 - 0x0
      12'h4A: dout  = 8'b00000000; //   74 :   0 - 0x0
      12'h4B: dout  = 8'b00010000; //   75 :  16 - 0x10
      12'h4C: dout  = 8'b00110000; //   76 :  48 - 0x30
      12'h4D: dout  = 8'b00000000; //   77 :   0 - 0x0
      12'h4E: dout  = 8'b11111000; //   78 : 248 - 0xf8
      12'h4F: dout  = 8'b11111110; //   79 : 254 - 0xfe
      12'h50: dout  = 8'b00011111; //   80 :  31 - 0x1f -- Sprite 0xa
      12'h51: dout  = 8'b00111111; //   81 :  63 - 0x3f
      12'h52: dout  = 8'b00111111; //   82 :  63 - 0x3f
      12'h53: dout  = 8'b00011111; //   83 :  31 - 0x1f
      12'h54: dout  = 8'b00000111; //   84 :   7 - 0x7
      12'h55: dout  = 8'b00001000; //   85 :   8 - 0x8
      12'h56: dout  = 8'b00010111; //   86 :  23 - 0x17
      12'h57: dout  = 8'b00010111; //   87 :  23 - 0x17
      12'h58: dout  = 8'b11111111; //   88 : 255 - 0xff -- Sprite 0xb
      12'h59: dout  = 8'b11111111; //   89 : 255 - 0xff
      12'h5A: dout  = 8'b11111110; //   90 : 254 - 0xfe
      12'h5B: dout  = 8'b11111110; //   91 : 254 - 0xfe
      12'h5C: dout  = 8'b11111100; //   92 : 252 - 0xfc
      12'h5D: dout  = 8'b11100000; //   93 : 224 - 0xe0
      12'h5E: dout  = 8'b01000000; //   94 :  64 - 0x40
      12'h5F: dout  = 8'b10100000; //   95 : 160 - 0xa0
      12'h60: dout  = 8'b00110111; //   96 :  55 - 0x37 -- Sprite 0xc
      12'h61: dout  = 8'b00100111; //   97 :  39 - 0x27
      12'h62: dout  = 8'b00100011; //   98 :  35 - 0x23
      12'h63: dout  = 8'b00000011; //   99 :   3 - 0x3
      12'h64: dout  = 8'b00000001; //  100 :   1 - 0x1
      12'h65: dout  = 8'b00000000; //  101 :   0 - 0x0
      12'h66: dout  = 8'b00000000; //  102 :   0 - 0x0
      12'h67: dout  = 8'b00000000; //  103 :   0 - 0x0
      12'h68: dout  = 8'b11001100; //  104 : 204 - 0xcc -- Sprite 0xd
      12'h69: dout  = 8'b11111111; //  105 : 255 - 0xff
      12'h6A: dout  = 8'b11111111; //  106 : 255 - 0xff
      12'h6B: dout  = 8'b11111111; //  107 : 255 - 0xff
      12'h6C: dout  = 8'b11111111; //  108 : 255 - 0xff
      12'h6D: dout  = 8'b01110000; //  109 : 112 - 0x70
      12'h6E: dout  = 8'b00000000; //  110 :   0 - 0x0
      12'h6F: dout  = 8'b00001000; //  111 :   8 - 0x8
      12'h70: dout  = 8'b11110000; //  112 : 240 - 0xf0 -- Sprite 0xe
      12'h71: dout  = 8'b11110000; //  113 : 240 - 0xf0
      12'h72: dout  = 8'b11110000; //  114 : 240 - 0xf0
      12'h73: dout  = 8'b11110000; //  115 : 240 - 0xf0
      12'h74: dout  = 8'b11110000; //  116 : 240 - 0xf0
      12'h75: dout  = 8'b11000000; //  117 : 192 - 0xc0
      12'h76: dout  = 8'b10000000; //  118 : 128 - 0x80
      12'h77: dout  = 8'b00000000; //  119 :   0 - 0x0
      12'h78: dout  = 8'b00010000; //  120 :  16 - 0x10 -- Sprite 0xf
      12'h79: dout  = 8'b01100000; //  121 :  96 - 0x60
      12'h7A: dout  = 8'b10000000; //  122 : 128 - 0x80
      12'h7B: dout  = 8'b00000000; //  123 :   0 - 0x0
      12'h7C: dout  = 8'b01111000; //  124 : 120 - 0x78
      12'h7D: dout  = 8'b01111000; //  125 : 120 - 0x78
      12'h7E: dout  = 8'b01111110; //  126 : 126 - 0x7e
      12'h7F: dout  = 8'b01111110; //  127 : 126 - 0x7e
      12'h80: dout  = 8'b00000000; //  128 :   0 - 0x0 -- Sprite 0x10
      12'h81: dout  = 8'b00000000; //  129 :   0 - 0x0
      12'h82: dout  = 8'b00000000; //  130 :   0 - 0x0
      12'h83: dout  = 8'b00000000; //  131 :   0 - 0x0
      12'h84: dout  = 8'b00000000; //  132 :   0 - 0x0
      12'h85: dout  = 8'b00011111; //  133 :  31 - 0x1f
      12'h86: dout  = 8'b00111111; //  134 :  63 - 0x3f
      12'h87: dout  = 8'b00111111; //  135 :  63 - 0x3f
      12'h88: dout  = 8'b00000000; //  136 :   0 - 0x0 -- Sprite 0x11
      12'h89: dout  = 8'b00000000; //  137 :   0 - 0x0
      12'h8A: dout  = 8'b00100000; //  138 :  32 - 0x20
      12'h8B: dout  = 8'b01100000; //  139 :  96 - 0x60
      12'h8C: dout  = 8'b00000000; //  140 :   0 - 0x0
      12'h8D: dout  = 8'b11110000; //  141 : 240 - 0xf0
      12'h8E: dout  = 8'b11111100; //  142 : 252 - 0xfc
      12'h8F: dout  = 8'b11111110; //  143 : 254 - 0xfe
      12'h90: dout  = 8'b01111111; //  144 : 127 - 0x7f -- Sprite 0x12
      12'h91: dout  = 8'b01111111; //  145 : 127 - 0x7f
      12'h92: dout  = 8'b00111111; //  146 :  63 - 0x3f
      12'h93: dout  = 8'b00011111; //  147 :  31 - 0x1f
      12'h94: dout  = 8'b00000000; //  148 :   0 - 0x0
      12'h95: dout  = 8'b00010110; //  149 :  22 - 0x16
      12'h96: dout  = 8'b00101111; //  150 :  47 - 0x2f
      12'h97: dout  = 8'b00101111; //  151 :  47 - 0x2f
      12'h98: dout  = 8'b11111110; //  152 : 254 - 0xfe -- Sprite 0x13
      12'h99: dout  = 8'b11111100; //  153 : 252 - 0xfc
      12'h9A: dout  = 8'b11111100; //  154 : 252 - 0xfc
      12'h9B: dout  = 8'b11111000; //  155 : 248 - 0xf8
      12'h9C: dout  = 8'b11000000; //  156 : 192 - 0xc0
      12'h9D: dout  = 8'b01100000; //  157 :  96 - 0x60
      12'h9E: dout  = 8'b00100000; //  158 :  32 - 0x20
      12'h9F: dout  = 8'b00110000; //  159 :  48 - 0x30
      12'hA0: dout  = 8'b00101111; //  160 :  47 - 0x2f -- Sprite 0x14
      12'hA1: dout  = 8'b00101111; //  161 :  47 - 0x2f
      12'hA2: dout  = 8'b00101111; //  162 :  47 - 0x2f
      12'hA3: dout  = 8'b00001111; //  163 :  15 - 0xf
      12'hA4: dout  = 8'b00000111; //  164 :   7 - 0x7
      12'hA5: dout  = 8'b00000011; //  165 :   3 - 0x3
      12'hA6: dout  = 8'b00000000; //  166 :   0 - 0x0
      12'hA7: dout  = 8'b00000000; //  167 :   0 - 0x0
      12'hA8: dout  = 8'b00010000; //  168 :  16 - 0x10 -- Sprite 0x15
      12'hA9: dout  = 8'b11110000; //  169 : 240 - 0xf0
      12'hAA: dout  = 8'b11110000; //  170 : 240 - 0xf0
      12'hAB: dout  = 8'b11110000; //  171 : 240 - 0xf0
      12'hAC: dout  = 8'b11110000; //  172 : 240 - 0xf0
      12'hAD: dout  = 8'b11100000; //  173 : 224 - 0xe0
      12'hAE: dout  = 8'b11000000; //  174 : 192 - 0xc0
      12'hAF: dout  = 8'b11100000; //  175 : 224 - 0xe0
      12'hB0: dout  = 8'b00000001; //  176 :   1 - 0x1 -- Sprite 0x16
      12'hB1: dout  = 8'b00000011; //  177 :   3 - 0x3
      12'hB2: dout  = 8'b00000001; //  178 :   1 - 0x1
      12'hB3: dout  = 8'b00000100; //  179 :   4 - 0x4
      12'hB4: dout  = 8'b00000111; //  180 :   7 - 0x7
      12'hB5: dout  = 8'b00001111; //  181 :  15 - 0xf
      12'hB6: dout  = 8'b00001111; //  182 :  15 - 0xf
      12'hB7: dout  = 8'b00000011; //  183 :   3 - 0x3
      12'hB8: dout  = 8'b11111000; //  184 : 248 - 0xf8 -- Sprite 0x17
      12'hB9: dout  = 8'b11110000; //  185 : 240 - 0xf0
      12'hBA: dout  = 8'b11100000; //  186 : 224 - 0xe0
      12'hBB: dout  = 8'b01110000; //  187 : 112 - 0x70
      12'hBC: dout  = 8'b10110000; //  188 : 176 - 0xb0
      12'hBD: dout  = 8'b10000000; //  189 : 128 - 0x80
      12'hBE: dout  = 8'b11100000; //  190 : 224 - 0xe0
      12'hBF: dout  = 8'b11100000; //  191 : 224 - 0xe0
      12'hC0: dout  = 8'b00000000; //  192 :   0 - 0x0 -- Sprite 0x18
      12'hC1: dout  = 8'b00110000; //  193 :  48 - 0x30
      12'hC2: dout  = 8'b01110000; //  194 : 112 - 0x70
      12'hC3: dout  = 8'b01111111; //  195 : 127 - 0x7f
      12'hC4: dout  = 8'b11111111; //  196 : 255 - 0xff
      12'hC5: dout  = 8'b11111111; //  197 : 255 - 0xff
      12'hC6: dout  = 8'b11110111; //  198 : 247 - 0xf7
      12'hC7: dout  = 8'b11110011; //  199 : 243 - 0xf3
      12'hC8: dout  = 8'b00000000; //  200 :   0 - 0x0 -- Sprite 0x19
      12'hC9: dout  = 8'b00011000; //  201 :  24 - 0x18
      12'hCA: dout  = 8'b00010000; //  202 :  16 - 0x10
      12'hCB: dout  = 8'b00000000; //  203 :   0 - 0x0
      12'hCC: dout  = 8'b11111000; //  204 : 248 - 0xf8
      12'hCD: dout  = 8'b11111000; //  205 : 248 - 0xf8
      12'hCE: dout  = 8'b11111110; //  206 : 254 - 0xfe
      12'hCF: dout  = 8'b11111111; //  207 : 255 - 0xff
      12'hD0: dout  = 8'b11100111; //  208 : 231 - 0xe7 -- Sprite 0x1a
      12'hD1: dout  = 8'b00001111; //  209 :  15 - 0xf
      12'hD2: dout  = 8'b00001111; //  210 :  15 - 0xf
      12'hD3: dout  = 8'b00011111; //  211 :  31 - 0x1f
      12'hD4: dout  = 8'b00011111; //  212 :  31 - 0x1f
      12'hD5: dout  = 8'b00011111; //  213 :  31 - 0x1f
      12'hD6: dout  = 8'b00001111; //  214 :  15 - 0xf
      12'hD7: dout  = 8'b00000111; //  215 :   7 - 0x7
      12'hD8: dout  = 8'b11111111; //  216 : 255 - 0xff -- Sprite 0x1b
      12'hD9: dout  = 8'b11111110; //  217 : 254 - 0xfe
      12'hDA: dout  = 8'b11111100; //  218 : 252 - 0xfc
      12'hDB: dout  = 8'b11000110; //  219 : 198 - 0xc6
      12'hDC: dout  = 8'b10001110; //  220 : 142 - 0x8e
      12'hDD: dout  = 8'b11101110; //  221 : 238 - 0xee
      12'hDE: dout  = 8'b11111111; //  222 : 255 - 0xff
      12'hDF: dout  = 8'b11111111; //  223 : 255 - 0xff
      12'hE0: dout  = 8'b00000011; //  224 :   3 - 0x3 -- Sprite 0x1c
      12'hE1: dout  = 8'b00000000; //  225 :   0 - 0x0
      12'hE2: dout  = 8'b00000000; //  226 :   0 - 0x0
      12'hE3: dout  = 8'b00001110; //  227 :  14 - 0xe
      12'hE4: dout  = 8'b00000111; //  228 :   7 - 0x7
      12'hE5: dout  = 8'b00111111; //  229 :  63 - 0x3f
      12'hE6: dout  = 8'b00111111; //  230 :  63 - 0x3f
      12'hE7: dout  = 8'b00111111; //  231 :  63 - 0x3f
      12'hE8: dout  = 8'b11111111; //  232 : 255 - 0xff -- Sprite 0x1d
      12'hE9: dout  = 8'b01111111; //  233 : 127 - 0x7f
      12'hEA: dout  = 8'b00111111; //  234 :  63 - 0x3f
      12'hEB: dout  = 8'b00001110; //  235 :  14 - 0xe
      12'hEC: dout  = 8'b11000000; //  236 : 192 - 0xc0
      12'hED: dout  = 8'b11000000; //  237 : 192 - 0xc0
      12'hEE: dout  = 8'b11100000; //  238 : 224 - 0xe0
      12'hEF: dout  = 8'b11100000; //  239 : 224 - 0xe0
      12'hF0: dout  = 8'b00000000; //  240 :   0 - 0x0 -- Sprite 0x1e
      12'hF1: dout  = 8'b10000000; //  241 : 128 - 0x80
      12'hF2: dout  = 8'b11001000; //  242 : 200 - 0xc8
      12'hF3: dout  = 8'b11111110; //  243 : 254 - 0xfe
      12'hF4: dout  = 8'b01111111; //  244 : 127 - 0x7f
      12'hF5: dout  = 8'b00111111; //  245 :  63 - 0x3f
      12'hF6: dout  = 8'b00011110; //  246 :  30 - 0x1e
      12'hF7: dout  = 8'b00001110; //  247 :  14 - 0xe
      12'hF8: dout  = 8'b11100000; //  248 : 224 - 0xe0 -- Sprite 0x1f
      12'hF9: dout  = 8'b00000000; //  249 :   0 - 0x0
      12'hFA: dout  = 8'b00000000; //  250 :   0 - 0x0
      12'hFB: dout  = 8'b00000000; //  251 :   0 - 0x0
      12'hFC: dout  = 8'b00000000; //  252 :   0 - 0x0
      12'hFD: dout  = 8'b00000000; //  253 :   0 - 0x0
      12'hFE: dout  = 8'b00000000; //  254 :   0 - 0x0
      12'hFF: dout  = 8'b00000000; //  255 :   0 - 0x0
      12'h100: dout  = 8'b00000000; //  256 :   0 - 0x0 -- Sprite 0x20
      12'h101: dout  = 8'b00000000; //  257 :   0 - 0x0
      12'h102: dout  = 8'b00000000; //  258 :   0 - 0x0
      12'h103: dout  = 8'b00000000; //  259 :   0 - 0x0
      12'h104: dout  = 8'b00000000; //  260 :   0 - 0x0
      12'h105: dout  = 8'b00000000; //  261 :   0 - 0x0
      12'h106: dout  = 8'b00011111; //  262 :  31 - 0x1f
      12'h107: dout  = 8'b00111111; //  263 :  63 - 0x3f
      12'h108: dout  = 8'b00001110; //  264 :  14 - 0xe -- Sprite 0x21
      12'h109: dout  = 8'b00011111; //  265 :  31 - 0x1f
      12'h10A: dout  = 8'b00011111; //  266 :  31 - 0x1f
      12'h10B: dout  = 8'b00011111; //  267 :  31 - 0x1f
      12'h10C: dout  = 8'b00011111; //  268 :  31 - 0x1f
      12'h10D: dout  = 8'b00000011; //  269 :   3 - 0x3
      12'h10E: dout  = 8'b11111111; //  270 : 255 - 0xff
      12'h10F: dout  = 8'b11111111; //  271 : 255 - 0xff
      12'h110: dout  = 8'b00111111; //  272 :  63 - 0x3f -- Sprite 0x22
      12'h111: dout  = 8'b00111111; //  273 :  63 - 0x3f
      12'h112: dout  = 8'b01111111; //  274 : 127 - 0x7f
      12'h113: dout  = 8'b01111111; //  275 : 127 - 0x7f
      12'h114: dout  = 8'b00011111; //  276 :  31 - 0x1f
      12'h115: dout  = 8'b00000000; //  277 :   0 - 0x0
      12'h116: dout  = 8'b01111110; //  278 : 126 - 0x7e
      12'h117: dout  = 8'b11111111; //  279 : 255 - 0xff
      12'h118: dout  = 8'b11111111; //  280 : 255 - 0xff -- Sprite 0x23
      12'h119: dout  = 8'b11111111; //  281 : 255 - 0xff
      12'h11A: dout  = 8'b11111110; //  282 : 254 - 0xfe
      12'h11B: dout  = 8'b11111110; //  283 : 254 - 0xfe
      12'h11C: dout  = 8'b11111110; //  284 : 254 - 0xfe
      12'h11D: dout  = 8'b11011110; //  285 : 222 - 0xde
      12'h11E: dout  = 8'b01011100; //  286 :  92 - 0x5c
      12'h11F: dout  = 8'b01101100; //  287 : 108 - 0x6c
      12'h120: dout  = 8'b11111111; //  288 : 255 - 0xff -- Sprite 0x24
      12'h121: dout  = 8'b11111111; //  289 : 255 - 0xff
      12'h122: dout  = 8'b11111110; //  290 : 254 - 0xfe
      12'h123: dout  = 8'b11111100; //  291 : 252 - 0xfc
      12'h124: dout  = 8'b11111000; //  292 : 248 - 0xf8
      12'h125: dout  = 8'b10110000; //  293 : 176 - 0xb0
      12'h126: dout  = 8'b01100000; //  294 :  96 - 0x60
      12'h127: dout  = 8'b00000000; //  295 :   0 - 0x0
      12'h128: dout  = 8'b00101000; //  296 :  40 - 0x28 -- Sprite 0x25
      12'h129: dout  = 8'b00110000; //  297 :  48 - 0x30
      12'h12A: dout  = 8'b00011000; //  298 :  24 - 0x18
      12'h12B: dout  = 8'b01000000; //  299 :  64 - 0x40
      12'h12C: dout  = 8'b00000000; //  300 :   0 - 0x0
      12'h12D: dout  = 8'b00000001; //  301 :   1 - 0x1
      12'h12E: dout  = 8'b00000011; //  302 :   3 - 0x3
      12'h12F: dout  = 8'b00001111; //  303 :  15 - 0xf
      12'h130: dout  = 8'b00010000; //  304 :  16 - 0x10 -- Sprite 0x26
      12'h131: dout  = 8'b11101100; //  305 : 236 - 0xec
      12'h132: dout  = 8'b11100011; //  306 : 227 - 0xe3
      12'h133: dout  = 8'b11100000; //  307 : 224 - 0xe0
      12'h134: dout  = 8'b11100000; //  308 : 224 - 0xe0
      12'h135: dout  = 8'b11100000; //  309 : 224 - 0xe0
      12'h136: dout  = 8'b11000000; //  310 : 192 - 0xc0
      12'h137: dout  = 8'b10000000; //  311 : 128 - 0x80
      12'h138: dout  = 8'b00001111; //  312 :  15 - 0xf -- Sprite 0x27
      12'h139: dout  = 8'b00001111; //  313 :  15 - 0xf
      12'h13A: dout  = 8'b00001111; //  314 :  15 - 0xf
      12'h13B: dout  = 8'b00001111; //  315 :  15 - 0xf
      12'h13C: dout  = 8'b00000000; //  316 :   0 - 0x0
      12'h13D: dout  = 8'b00000000; //  317 :   0 - 0x0
      12'h13E: dout  = 8'b00000000; //  318 :   0 - 0x0
      12'h13F: dout  = 8'b00000000; //  319 :   0 - 0x0
      12'h140: dout  = 8'b00011111; //  320 :  31 - 0x1f -- Sprite 0x28
      12'h141: dout  = 8'b00111111; //  321 :  63 - 0x3f
      12'h142: dout  = 8'b00111111; //  322 :  63 - 0x3f
      12'h143: dout  = 8'b00011111; //  323 :  31 - 0x1f
      12'h144: dout  = 8'b00000111; //  324 :   7 - 0x7
      12'h145: dout  = 8'b00001001; //  325 :   9 - 0x9
      12'h146: dout  = 8'b00010011; //  326 :  19 - 0x13
      12'h147: dout  = 8'b00010111; //  327 :  23 - 0x17
      12'h148: dout  = 8'b11111111; //  328 : 255 - 0xff -- Sprite 0x29
      12'h149: dout  = 8'b11111111; //  329 : 255 - 0xff
      12'h14A: dout  = 8'b11111110; //  330 : 254 - 0xfe
      12'h14B: dout  = 8'b11111111; //  331 : 255 - 0xff
      12'h14C: dout  = 8'b11111110; //  332 : 254 - 0xfe
      12'h14D: dout  = 8'b11111100; //  333 : 252 - 0xfc
      12'h14E: dout  = 8'b11111000; //  334 : 248 - 0xf8
      12'h14F: dout  = 8'b11100000; //  335 : 224 - 0xe0
      12'h150: dout  = 8'b00010111; //  336 :  23 - 0x17 -- Sprite 0x2a
      12'h151: dout  = 8'b00010111; //  337 :  23 - 0x17
      12'h152: dout  = 8'b00000011; //  338 :   3 - 0x3
      12'h153: dout  = 8'b00000000; //  339 :   0 - 0x0
      12'h154: dout  = 8'b00000000; //  340 :   0 - 0x0
      12'h155: dout  = 8'b00000000; //  341 :   0 - 0x0
      12'h156: dout  = 8'b00000000; //  342 :   0 - 0x0
      12'h157: dout  = 8'b00000000; //  343 :   0 - 0x0
      12'h158: dout  = 8'b11010000; //  344 : 208 - 0xd0 -- Sprite 0x2b
      12'h159: dout  = 8'b10010000; //  345 : 144 - 0x90
      12'h15A: dout  = 8'b00011000; //  346 :  24 - 0x18
      12'h15B: dout  = 8'b00001000; //  347 :   8 - 0x8
      12'h15C: dout  = 8'b01000000; //  348 :  64 - 0x40
      12'h15D: dout  = 8'b00000000; //  349 :   0 - 0x0
      12'h15E: dout  = 8'b00000000; //  350 :   0 - 0x0
      12'h15F: dout  = 8'b00000000; //  351 :   0 - 0x0
      12'h160: dout  = 8'b00110000; //  352 :  48 - 0x30 -- Sprite 0x2c
      12'h161: dout  = 8'b11110000; //  353 : 240 - 0xf0
      12'h162: dout  = 8'b11110000; //  354 : 240 - 0xf0
      12'h163: dout  = 8'b11110001; //  355 : 241 - 0xf1
      12'h164: dout  = 8'b11110110; //  356 : 246 - 0xf6
      12'h165: dout  = 8'b11000110; //  357 : 198 - 0xc6
      12'h166: dout  = 8'b10000100; //  358 : 132 - 0x84
      12'h167: dout  = 8'b00000000; //  359 :   0 - 0x0
      12'h168: dout  = 8'b00000000; //  360 :   0 - 0x0 -- Sprite 0x2d
      12'h169: dout  = 8'b00000000; //  361 :   0 - 0x0
      12'h16A: dout  = 8'b00000000; //  362 :   0 - 0x0
      12'h16B: dout  = 8'b00000000; //  363 :   0 - 0x0
      12'h16C: dout  = 8'b00000000; //  364 :   0 - 0x0
      12'h16D: dout  = 8'b00000000; //  365 :   0 - 0x0
      12'h16E: dout  = 8'b00000000; //  366 :   0 - 0x0
      12'h16F: dout  = 8'b00000000; //  367 :   0 - 0x0
      12'h170: dout  = 8'b00011111; //  368 :  31 - 0x1f -- Sprite 0x2e
      12'h171: dout  = 8'b00011111; //  369 :  31 - 0x1f
      12'h172: dout  = 8'b00111111; //  370 :  63 - 0x3f
      12'h173: dout  = 8'b00111110; //  371 :  62 - 0x3e
      12'h174: dout  = 8'b01111100; //  372 : 124 - 0x7c
      12'h175: dout  = 8'b01111000; //  373 : 120 - 0x78
      12'h176: dout  = 8'b11110000; //  374 : 240 - 0xf0
      12'h177: dout  = 8'b11100000; //  375 : 224 - 0xe0
      12'h178: dout  = 8'b10110000; //  376 : 176 - 0xb0 -- Sprite 0x2f
      12'h179: dout  = 8'b10010000; //  377 : 144 - 0x90
      12'h17A: dout  = 8'b00011000; //  378 :  24 - 0x18
      12'h17B: dout  = 8'b00001000; //  379 :   8 - 0x8
      12'h17C: dout  = 8'b01000000; //  380 :  64 - 0x40
      12'h17D: dout  = 8'b00000000; //  381 :   0 - 0x0
      12'h17E: dout  = 8'b00000000; //  382 :   0 - 0x0
      12'h17F: dout  = 8'b00000000; //  383 :   0 - 0x0
      12'h180: dout  = 8'b11000000; //  384 : 192 - 0xc0 -- Sprite 0x30
      12'h181: dout  = 8'b11100000; //  385 : 224 - 0xe0
      12'h182: dout  = 8'b11111100; //  386 : 252 - 0xfc
      12'h183: dout  = 8'b11111110; //  387 : 254 - 0xfe
      12'h184: dout  = 8'b11111111; //  388 : 255 - 0xff
      12'h185: dout  = 8'b01111111; //  389 : 127 - 0x7f
      12'h186: dout  = 8'b00000011; //  390 :   3 - 0x3
      12'h187: dout  = 8'b00000000; //  391 :   0 - 0x0
      12'h188: dout  = 8'b00000000; //  392 :   0 - 0x0 -- Sprite 0x31
      12'h189: dout  = 8'b00000000; //  393 :   0 - 0x0
      12'h18A: dout  = 8'b00010000; //  394 :  16 - 0x10
      12'h18B: dout  = 8'b00111000; //  395 :  56 - 0x38
      12'h18C: dout  = 8'b00111110; //  396 :  62 - 0x3e
      12'h18D: dout  = 8'b00111100; //  397 :  60 - 0x3c
      12'h18E: dout  = 8'b00111000; //  398 :  56 - 0x38
      12'h18F: dout  = 8'b00011000; //  399 :  24 - 0x18
      12'h190: dout  = 8'b00000000; //  400 :   0 - 0x0 -- Sprite 0x32
      12'h191: dout  = 8'b00000000; //  401 :   0 - 0x0
      12'h192: dout  = 8'b00000000; //  402 :   0 - 0x0
      12'h193: dout  = 8'b00000111; //  403 :   7 - 0x7
      12'h194: dout  = 8'b00001111; //  404 :  15 - 0xf
      12'h195: dout  = 8'b00001111; //  405 :  15 - 0xf
      12'h196: dout  = 8'b00001111; //  406 :  15 - 0xf
      12'h197: dout  = 8'b00000011; //  407 :   3 - 0x3
      12'h198: dout  = 8'b00000000; //  408 :   0 - 0x0 -- Sprite 0x33
      12'h199: dout  = 8'b00000000; //  409 :   0 - 0x0
      12'h19A: dout  = 8'b00000000; //  410 :   0 - 0x0
      12'h19B: dout  = 8'b11110000; //  411 : 240 - 0xf0
      12'h19C: dout  = 8'b11111100; //  412 : 252 - 0xfc
      12'h19D: dout  = 8'b11111110; //  413 : 254 - 0xfe
      12'h19E: dout  = 8'b11111100; //  414 : 252 - 0xfc
      12'h19F: dout  = 8'b11111000; //  415 : 248 - 0xf8
      12'h1A0: dout  = 8'b00000111; //  416 :   7 - 0x7 -- Sprite 0x34
      12'h1A1: dout  = 8'b00001111; //  417 :  15 - 0xf
      12'h1A2: dout  = 8'b00011011; //  418 :  27 - 0x1b
      12'h1A3: dout  = 8'b00011000; //  419 :  24 - 0x18
      12'h1A4: dout  = 8'b00010000; //  420 :  16 - 0x10
      12'h1A5: dout  = 8'b00110000; //  421 :  48 - 0x30
      12'h1A6: dout  = 8'b00100001; //  422 :  33 - 0x21
      12'h1A7: dout  = 8'b00000001; //  423 :   1 - 0x1
      12'h1A8: dout  = 8'b10101000; //  424 : 168 - 0xa8 -- Sprite 0x35
      12'h1A9: dout  = 8'b11111100; //  425 : 252 - 0xfc
      12'h1AA: dout  = 8'b11111000; //  426 : 248 - 0xf8
      12'h1AB: dout  = 8'b00000000; //  427 :   0 - 0x0
      12'h1AC: dout  = 8'b00000000; //  428 :   0 - 0x0
      12'h1AD: dout  = 8'b00000000; //  429 :   0 - 0x0
      12'h1AE: dout  = 8'b11000000; //  430 : 192 - 0xc0
      12'h1AF: dout  = 8'b11100000; //  431 : 224 - 0xe0
      12'h1B0: dout  = 8'b00000000; //  432 :   0 - 0x0 -- Sprite 0x36
      12'h1B1: dout  = 8'b00000000; //  433 :   0 - 0x0
      12'h1B2: dout  = 8'b00001111; //  434 :  15 - 0xf
      12'h1B3: dout  = 8'b00011111; //  435 :  31 - 0x1f
      12'h1B4: dout  = 8'b00011111; //  436 :  31 - 0x1f
      12'h1B5: dout  = 8'b00011111; //  437 :  31 - 0x1f
      12'h1B6: dout  = 8'b00000111; //  438 :   7 - 0x7
      12'h1B7: dout  = 8'b00111100; //  439 :  60 - 0x3c
      12'h1B8: dout  = 8'b00000000; //  440 :   0 - 0x0 -- Sprite 0x37
      12'h1B9: dout  = 8'b00000000; //  441 :   0 - 0x0
      12'h1BA: dout  = 8'b11100000; //  442 : 224 - 0xe0
      12'h1BB: dout  = 8'b11111000; //  443 : 248 - 0xf8
      12'h1BC: dout  = 8'b11111100; //  444 : 252 - 0xfc
      12'h1BD: dout  = 8'b11111000; //  445 : 248 - 0xf8
      12'h1BE: dout  = 8'b11110000; //  446 : 240 - 0xf0
      12'h1BF: dout  = 8'b11000000; //  447 : 192 - 0xc0
      12'h1C0: dout  = 8'b11111100; //  448 : 252 - 0xfc -- Sprite 0x38
      12'h1C1: dout  = 8'b11101101; //  449 : 237 - 0xed
      12'h1C2: dout  = 8'b11000000; //  450 : 192 - 0xc0
      12'h1C3: dout  = 8'b00000000; //  451 :   0 - 0x0
      12'h1C4: dout  = 8'b00000000; //  452 :   0 - 0x0
      12'h1C5: dout  = 8'b01100000; //  453 :  96 - 0x60
      12'h1C6: dout  = 8'b01110000; //  454 : 112 - 0x70
      12'h1C7: dout  = 8'b00111000; //  455 :  56 - 0x38
      12'h1C8: dout  = 8'b01111110; //  456 : 126 - 0x7e -- Sprite 0x39
      12'h1C9: dout  = 8'b00011110; //  457 :  30 - 0x1e
      12'h1CA: dout  = 8'b00000100; //  458 :   4 - 0x4
      12'h1CB: dout  = 8'b00001100; //  459 :  12 - 0xc
      12'h1CC: dout  = 8'b00001100; //  460 :  12 - 0xc
      12'h1CD: dout  = 8'b00001100; //  461 :  12 - 0xc
      12'h1CE: dout  = 8'b00000000; //  462 :   0 - 0x0
      12'h1CF: dout  = 8'b00000000; //  463 :   0 - 0x0
      12'h1D0: dout  = 8'b00000000; //  464 :   0 - 0x0 -- Sprite 0x3a
      12'h1D1: dout  = 8'b00000000; //  465 :   0 - 0x0
      12'h1D2: dout  = 8'b00001111; //  466 :  15 - 0xf
      12'h1D3: dout  = 8'b00011111; //  467 :  31 - 0x1f
      12'h1D4: dout  = 8'b00011111; //  468 :  31 - 0x1f
      12'h1D5: dout  = 8'b00011111; //  469 :  31 - 0x1f
      12'h1D6: dout  = 8'b00000111; //  470 :   7 - 0x7
      12'h1D7: dout  = 8'b00001101; //  471 :  13 - 0xd
      12'h1D8: dout  = 8'b00011110; //  472 :  30 - 0x1e -- Sprite 0x3b
      12'h1D9: dout  = 8'b00011100; //  473 :  28 - 0x1c
      12'h1DA: dout  = 8'b00011110; //  474 :  30 - 0x1e
      12'h1DB: dout  = 8'b00001111; //  475 :  15 - 0xf
      12'h1DC: dout  = 8'b00000111; //  476 :   7 - 0x7
      12'h1DD: dout  = 8'b00000000; //  477 :   0 - 0x0
      12'h1DE: dout  = 8'b00000111; //  478 :   7 - 0x7
      12'h1DF: dout  = 8'b00000111; //  479 :   7 - 0x7
      12'h1E0: dout  = 8'b01100000; //  480 :  96 - 0x60 -- Sprite 0x3c
      12'h1E1: dout  = 8'b10010000; //  481 : 144 - 0x90
      12'h1E2: dout  = 8'b00000000; //  482 :   0 - 0x0
      12'h1E3: dout  = 8'b10000000; //  483 : 128 - 0x80
      12'h1E4: dout  = 8'b00000000; //  484 :   0 - 0x0
      12'h1E5: dout  = 8'b11100000; //  485 : 224 - 0xe0
      12'h1E6: dout  = 8'b11110000; //  486 : 240 - 0xf0
      12'h1E7: dout  = 8'b10000000; //  487 : 128 - 0x80
      12'h1E8: dout  = 8'b00000000; //  488 :   0 - 0x0 -- Sprite 0x3d
      12'h1E9: dout  = 8'b00010000; //  489 :  16 - 0x10
      12'h1EA: dout  = 8'b00111111; //  490 :  63 - 0x3f
      12'h1EB: dout  = 8'b01111111; //  491 : 127 - 0x7f
      12'h1EC: dout  = 8'b01111111; //  492 : 127 - 0x7f
      12'h1ED: dout  = 8'b00111111; //  493 :  63 - 0x3f
      12'h1EE: dout  = 8'b00000011; //  494 :   3 - 0x3
      12'h1EF: dout  = 8'b00001111; //  495 :  15 - 0xf
      12'h1F0: dout  = 8'b00000000; //  496 :   0 - 0x0 -- Sprite 0x3e
      12'h1F1: dout  = 8'b00000000; //  497 :   0 - 0x0
      12'h1F2: dout  = 8'b11100000; //  498 : 224 - 0xe0
      12'h1F3: dout  = 8'b11111000; //  499 : 248 - 0xf8
      12'h1F4: dout  = 8'b11111100; //  500 : 252 - 0xfc
      12'h1F5: dout  = 8'b11111000; //  501 : 248 - 0xf8
      12'h1F6: dout  = 8'b10110000; //  502 : 176 - 0xb0
      12'h1F7: dout  = 8'b00111000; //  503 :  56 - 0x38
      12'h1F8: dout  = 8'b00011111; //  504 :  31 - 0x1f -- Sprite 0x3f
      12'h1F9: dout  = 8'b00000111; //  505 :   7 - 0x7
      12'h1FA: dout  = 8'b00000000; //  506 :   0 - 0x0
      12'h1FB: dout  = 8'b00001110; //  507 :  14 - 0xe
      12'h1FC: dout  = 8'b00001111; //  508 :  15 - 0xf
      12'h1FD: dout  = 8'b01010011; //  509 :  83 - 0x53
      12'h1FE: dout  = 8'b01111100; //  510 : 124 - 0x7c
      12'h1FF: dout  = 8'b00111100; //  511 :  60 - 0x3c
      12'h200: dout  = 8'b11111000; //  512 : 248 - 0xf8 -- Sprite 0x40
      12'h201: dout  = 8'b11111000; //  513 : 248 - 0xf8
      12'h202: dout  = 8'b11110000; //  514 : 240 - 0xf0
      12'h203: dout  = 8'b00000000; //  515 :   0 - 0x0
      12'h204: dout  = 8'b00000000; //  516 :   0 - 0x0
      12'h205: dout  = 8'b10000000; //  517 : 128 - 0x80
      12'h206: dout  = 8'b00000000; //  518 :   0 - 0x0
      12'h207: dout  = 8'b00000000; //  519 :   0 - 0x0
      12'h208: dout  = 8'b00000111; //  520 :   7 - 0x7 -- Sprite 0x41
      12'h209: dout  = 8'b00000111; //  521 :   7 - 0x7
      12'h20A: dout  = 8'b00000011; //  522 :   3 - 0x3
      12'h20B: dout  = 8'b11110111; //  523 : 247 - 0xf7
      12'h20C: dout  = 8'b11111111; //  524 : 255 - 0xff
      12'h20D: dout  = 8'b11111111; //  525 : 255 - 0xff
      12'h20E: dout  = 8'b11111110; //  526 : 254 - 0xfe
      12'h20F: dout  = 8'b11111100; //  527 : 252 - 0xfc
      12'h210: dout  = 8'b00111110; //  528 :  62 - 0x3e -- Sprite 0x42
      12'h211: dout  = 8'b01111111; //  529 : 127 - 0x7f
      12'h212: dout  = 8'b11111111; //  530 : 255 - 0xff
      12'h213: dout  = 8'b11100010; //  531 : 226 - 0xe2
      12'h214: dout  = 8'b01010000; //  532 :  80 - 0x50
      12'h215: dout  = 8'b00111000; //  533 :  56 - 0x38
      12'h216: dout  = 8'b01110000; //  534 : 112 - 0x70
      12'h217: dout  = 8'b01000000; //  535 :  64 - 0x40
      12'h218: dout  = 8'b11101000; //  536 : 232 - 0xe8 -- Sprite 0x43
      12'h219: dout  = 8'b01110001; //  537 : 113 - 0x71
      12'h21A: dout  = 8'b00000001; //  538 :   1 - 0x1
      12'h21B: dout  = 8'b01001011; //  539 :  75 - 0x4b
      12'h21C: dout  = 8'b00000011; //  540 :   3 - 0x3
      12'h21D: dout  = 8'b00000011; //  541 :   3 - 0x3
      12'h21E: dout  = 8'b00000000; //  542 :   0 - 0x0
      12'h21F: dout  = 8'b00000000; //  543 :   0 - 0x0
      12'h220: dout  = 8'b00000101; //  544 :   5 - 0x5 -- Sprite 0x44
      12'h221: dout  = 8'b00000011; //  545 :   3 - 0x3
      12'h222: dout  = 8'b00000001; //  546 :   1 - 0x1
      12'h223: dout  = 8'b00110000; //  547 :  48 - 0x30
      12'h224: dout  = 8'b00110000; //  548 :  48 - 0x30
      12'h225: dout  = 8'b00110000; //  549 :  48 - 0x30
      12'h226: dout  = 8'b00100110; //  550 :  38 - 0x26
      12'h227: dout  = 8'b00000100; //  551 :   4 - 0x4
      12'h228: dout  = 8'b11111110; //  552 : 254 - 0xfe -- Sprite 0x45
      12'h229: dout  = 8'b11111100; //  553 : 252 - 0xfc
      12'h22A: dout  = 8'b11100000; //  554 : 224 - 0xe0
      12'h22B: dout  = 8'b00000000; //  555 :   0 - 0x0
      12'h22C: dout  = 8'b00000000; //  556 :   0 - 0x0
      12'h22D: dout  = 8'b00000000; //  557 :   0 - 0x0
      12'h22E: dout  = 8'b00000000; //  558 :   0 - 0x0
      12'h22F: dout  = 8'b00000000; //  559 :   0 - 0x0
      12'h230: dout  = 8'b00000101; //  560 :   5 - 0x5 -- Sprite 0x46
      12'h231: dout  = 8'b00000011; //  561 :   3 - 0x3
      12'h232: dout  = 8'b00000001; //  562 :   1 - 0x1
      12'h233: dout  = 8'b00010000; //  563 :  16 - 0x10
      12'h234: dout  = 8'b00110000; //  564 :  48 - 0x30
      12'h235: dout  = 8'b00001100; //  565 :  12 - 0xc
      12'h236: dout  = 8'b00011100; //  566 :  28 - 0x1c
      12'h237: dout  = 8'b00011000; //  567 :  24 - 0x18
      12'h238: dout  = 8'b11000000; //  568 : 192 - 0xc0 -- Sprite 0x47
      12'h239: dout  = 8'b11100000; //  569 : 224 - 0xe0
      12'h23A: dout  = 8'b11110000; //  570 : 240 - 0xf0
      12'h23B: dout  = 8'b01111000; //  571 : 120 - 0x78
      12'h23C: dout  = 8'b00011000; //  572 :  24 - 0x18
      12'h23D: dout  = 8'b00001000; //  573 :   8 - 0x8
      12'h23E: dout  = 8'b00000000; //  574 :   0 - 0x0
      12'h23F: dout  = 8'b00000000; //  575 :   0 - 0x0
      12'h240: dout  = 8'b00000111; //  576 :   7 - 0x7 -- Sprite 0x48
      12'h241: dout  = 8'b00001111; //  577 :  15 - 0xf
      12'h242: dout  = 8'b00111110; //  578 :  62 - 0x3e
      12'h243: dout  = 8'b01111100; //  579 : 124 - 0x7c
      12'h244: dout  = 8'b00110000; //  580 :  48 - 0x30
      12'h245: dout  = 8'b00001100; //  581 :  12 - 0xc
      12'h246: dout  = 8'b00011100; //  582 :  28 - 0x1c
      12'h247: dout  = 8'b00011000; //  583 :  24 - 0x18
      12'h248: dout  = 8'b01100000; //  584 :  96 - 0x60 -- Sprite 0x49
      12'h249: dout  = 8'b01100000; //  585 :  96 - 0x60
      12'h24A: dout  = 8'b01100000; //  586 :  96 - 0x60
      12'h24B: dout  = 8'b10000000; //  587 : 128 - 0x80
      12'h24C: dout  = 8'b00000000; //  588 :   0 - 0x0
      12'h24D: dout  = 8'b00000000; //  589 :   0 - 0x0
      12'h24E: dout  = 8'b00000000; //  590 :   0 - 0x0
      12'h24F: dout  = 8'b00000000; //  591 :   0 - 0x0
      12'h250: dout  = 8'b01110011; //  592 : 115 - 0x73 -- Sprite 0x4a
      12'h251: dout  = 8'b11110011; //  593 : 243 - 0xf3
      12'h252: dout  = 8'b11110000; //  594 : 240 - 0xf0
      12'h253: dout  = 8'b11110100; //  595 : 244 - 0xf4
      12'h254: dout  = 8'b11110000; //  596 : 240 - 0xf0
      12'h255: dout  = 8'b11110000; //  597 : 240 - 0xf0
      12'h256: dout  = 8'b01110000; //  598 : 112 - 0x70
      12'h257: dout  = 8'b01100000; //  599 :  96 - 0x60
      12'h258: dout  = 8'b00000000; //  600 :   0 - 0x0 -- Sprite 0x4b
      12'h259: dout  = 8'b00000000; //  601 :   0 - 0x0
      12'h25A: dout  = 8'b00000000; //  602 :   0 - 0x0
      12'h25B: dout  = 8'b00000000; //  603 :   0 - 0x0
      12'h25C: dout  = 8'b00111100; //  604 :  60 - 0x3c
      12'h25D: dout  = 8'b00111100; //  605 :  60 - 0x3c
      12'h25E: dout  = 8'b11111100; //  606 : 252 - 0xfc
      12'h25F: dout  = 8'b11111100; //  607 : 252 - 0xfc
      12'h260: dout  = 8'b01111111; //  608 : 127 - 0x7f -- Sprite 0x4c
      12'h261: dout  = 8'b01111111; //  609 : 127 - 0x7f
      12'h262: dout  = 8'b00011111; //  610 :  31 - 0x1f
      12'h263: dout  = 8'b00000111; //  611 :   7 - 0x7
      12'h264: dout  = 8'b00001011; //  612 :  11 - 0xb
      12'h265: dout  = 8'b00011011; //  613 :  27 - 0x1b
      12'h266: dout  = 8'b00111011; //  614 :  59 - 0x3b
      12'h267: dout  = 8'b01111011; //  615 : 123 - 0x7b
      12'h268: dout  = 8'b11111100; //  616 : 252 - 0xfc -- Sprite 0x4d
      12'h269: dout  = 8'b11111100; //  617 : 252 - 0xfc
      12'h26A: dout  = 8'b11111000; //  618 : 248 - 0xf8
      12'h26B: dout  = 8'b11100000; //  619 : 224 - 0xe0
      12'h26C: dout  = 8'b11010000; //  620 : 208 - 0xd0
      12'h26D: dout  = 8'b11011000; //  621 : 216 - 0xd8
      12'h26E: dout  = 8'b11011100; //  622 : 220 - 0xdc
      12'h26F: dout  = 8'b11011110; //  623 : 222 - 0xde
      12'h270: dout  = 8'b11000100; //  624 : 196 - 0xc4 -- Sprite 0x4e
      12'h271: dout  = 8'b11100000; //  625 : 224 - 0xe0
      12'h272: dout  = 8'b11100000; //  626 : 224 - 0xe0
      12'h273: dout  = 8'b01000000; //  627 :  64 - 0x40
      12'h274: dout  = 8'b00000000; //  628 :   0 - 0x0
      12'h275: dout  = 8'b00111100; //  629 :  60 - 0x3c
      12'h276: dout  = 8'b00111100; //  630 :  60 - 0x3c
      12'h277: dout  = 8'b01111100; //  631 : 124 - 0x7c
      12'h278: dout  = 8'b00011101; //  632 :  29 - 0x1d -- Sprite 0x4f
      12'h279: dout  = 8'b00111100; //  633 :  60 - 0x3c
      12'h27A: dout  = 8'b00111010; //  634 :  58 - 0x3a
      12'h27B: dout  = 8'b00111000; //  635 :  56 - 0x38
      12'h27C: dout  = 8'b00110000; //  636 :  48 - 0x30
      12'h27D: dout  = 8'b00000000; //  637 :   0 - 0x0
      12'h27E: dout  = 8'b00011100; //  638 :  28 - 0x1c
      12'h27F: dout  = 8'b00111100; //  639 :  60 - 0x3c
      12'h280: dout  = 8'b00100010; //  640 :  34 - 0x22 -- Sprite 0x50
      12'h281: dout  = 8'b01010101; //  641 :  85 - 0x55
      12'h282: dout  = 8'b01010101; //  642 :  85 - 0x55
      12'h283: dout  = 8'b01010101; //  643 :  85 - 0x55
      12'h284: dout  = 8'b01010101; //  644 :  85 - 0x55
      12'h285: dout  = 8'b01010101; //  645 :  85 - 0x55
      12'h286: dout  = 8'b01110111; //  646 : 119 - 0x77
      12'h287: dout  = 8'b00100010; //  647 :  34 - 0x22
      12'h288: dout  = 8'b00000000; //  648 :   0 - 0x0 -- Sprite 0x51
      12'h289: dout  = 8'b00000000; //  649 :   0 - 0x0
      12'h28A: dout  = 8'b00000000; //  650 :   0 - 0x0
      12'h28B: dout  = 8'b00000000; //  651 :   0 - 0x0
      12'h28C: dout  = 8'b00000000; //  652 :   0 - 0x0
      12'h28D: dout  = 8'b00000000; //  653 :   0 - 0x0
      12'h28E: dout  = 8'b00000000; //  654 :   0 - 0x0
      12'h28F: dout  = 8'b00000000; //  655 :   0 - 0x0
      12'h290: dout  = 8'b00000000; //  656 :   0 - 0x0 -- Sprite 0x52
      12'h291: dout  = 8'b00000000; //  657 :   0 - 0x0
      12'h292: dout  = 8'b11001111; //  658 : 207 - 0xcf
      12'h293: dout  = 8'b00000111; //  659 :   7 - 0x7
      12'h294: dout  = 8'b01111111; //  660 : 127 - 0x7f
      12'h295: dout  = 8'b00000000; //  661 :   0 - 0x0
      12'h296: dout  = 8'b00000000; //  662 :   0 - 0x0
      12'h297: dout  = 8'b00000000; //  663 :   0 - 0x0
      12'h298: dout  = 8'b00000000; //  664 :   0 - 0x0 -- Sprite 0x53
      12'h299: dout  = 8'b00000000; //  665 :   0 - 0x0
      12'h29A: dout  = 8'b00111100; //  666 :  60 - 0x3c
      12'h29B: dout  = 8'b11111100; //  667 : 252 - 0xfc
      12'h29C: dout  = 8'b11111110; //  668 : 254 - 0xfe
      12'h29D: dout  = 8'b11100000; //  669 : 224 - 0xe0
      12'h29E: dout  = 8'b00000000; //  670 :   0 - 0x0
      12'h29F: dout  = 8'b00000000; //  671 :   0 - 0x0
      12'h2A0: dout  = 8'b01000000; //  672 :  64 - 0x40 -- Sprite 0x54
      12'h2A1: dout  = 8'b11100000; //  673 : 224 - 0xe0
      12'h2A2: dout  = 8'b01000000; //  674 :  64 - 0x40
      12'h2A3: dout  = 8'b00111111; //  675 :  63 - 0x3f
      12'h2A4: dout  = 8'b00111110; //  676 :  62 - 0x3e
      12'h2A5: dout  = 8'b00111110; //  677 :  62 - 0x3e
      12'h2A6: dout  = 8'b00110000; //  678 :  48 - 0x30
      12'h2A7: dout  = 8'b00111000; //  679 :  56 - 0x38
      12'h2A8: dout  = 8'b00000000; //  680 :   0 - 0x0 -- Sprite 0x55
      12'h2A9: dout  = 8'b00000000; //  681 :   0 - 0x0
      12'h2AA: dout  = 8'b00000000; //  682 :   0 - 0x0
      12'h2AB: dout  = 8'b11111000; //  683 : 248 - 0xf8
      12'h2AC: dout  = 8'b11111000; //  684 : 248 - 0xf8
      12'h2AD: dout  = 8'b11111000; //  685 : 248 - 0xf8
      12'h2AE: dout  = 8'b00011000; //  686 :  24 - 0x18
      12'h2AF: dout  = 8'b00111000; //  687 :  56 - 0x38
      12'h2B0: dout  = 8'b00111100; //  688 :  60 - 0x3c -- Sprite 0x56
      12'h2B1: dout  = 8'b00111001; //  689 :  57 - 0x39
      12'h2B2: dout  = 8'b00111011; //  690 :  59 - 0x3b
      12'h2B3: dout  = 8'b00111111; //  691 :  63 - 0x3f
      12'h2B4: dout  = 8'b00000000; //  692 :   0 - 0x0
      12'h2B5: dout  = 8'b00000000; //  693 :   0 - 0x0
      12'h2B6: dout  = 8'b00000000; //  694 :   0 - 0x0
      12'h2B7: dout  = 8'b00000000; //  695 :   0 - 0x0
      12'h2B8: dout  = 8'b01111000; //  696 : 120 - 0x78 -- Sprite 0x57
      12'h2B9: dout  = 8'b00111000; //  697 :  56 - 0x38
      12'h2BA: dout  = 8'b10111000; //  698 : 184 - 0xb8
      12'h2BB: dout  = 8'b11111000; //  699 : 248 - 0xf8
      12'h2BC: dout  = 8'b00000000; //  700 :   0 - 0x0
      12'h2BD: dout  = 8'b00000000; //  701 :   0 - 0x0
      12'h2BE: dout  = 8'b00000000; //  702 :   0 - 0x0
      12'h2BF: dout  = 8'b00000000; //  703 :   0 - 0x0
      12'h2C0: dout  = 8'b00111111; //  704 :  63 - 0x3f -- Sprite 0x58
      12'h2C1: dout  = 8'b00111111; //  705 :  63 - 0x3f
      12'h2C2: dout  = 8'b00001111; //  706 :  15 - 0xf
      12'h2C3: dout  = 8'b01110111; //  707 : 119 - 0x77
      12'h2C4: dout  = 8'b01110111; //  708 : 119 - 0x77
      12'h2C5: dout  = 8'b11110111; //  709 : 247 - 0xf7
      12'h2C6: dout  = 8'b11110111; //  710 : 247 - 0xf7
      12'h2C7: dout  = 8'b11110111; //  711 : 247 - 0xf7
      12'h2C8: dout  = 8'b11111111; //  712 : 255 - 0xff -- Sprite 0x59
      12'h2C9: dout  = 8'b11111110; //  713 : 254 - 0xfe
      12'h2CA: dout  = 8'b11111110; //  714 : 254 - 0xfe
      12'h2CB: dout  = 8'b11111110; //  715 : 254 - 0xfe
      12'h2CC: dout  = 8'b11111010; //  716 : 250 - 0xfa
      12'h2CD: dout  = 8'b11111010; //  717 : 250 - 0xfa
      12'h2CE: dout  = 8'b11110011; //  718 : 243 - 0xf3
      12'h2CF: dout  = 8'b11100111; //  719 : 231 - 0xe7
      12'h2D0: dout  = 8'b11110000; //  720 : 240 - 0xf0 -- Sprite 0x5a
      12'h2D1: dout  = 8'b11111000; //  721 : 248 - 0xf8
      12'h2D2: dout  = 8'b11111100; //  722 : 252 - 0xfc
      12'h2D3: dout  = 8'b01111100; //  723 : 124 - 0x7c
      12'h2D4: dout  = 8'b01111000; //  724 : 120 - 0x78
      12'h2D5: dout  = 8'b00111000; //  725 :  56 - 0x38
      12'h2D6: dout  = 8'b00111100; //  726 :  60 - 0x3c
      12'h2D7: dout  = 8'b11111100; //  727 : 252 - 0xfc
      12'h2D8: dout  = 8'b11111111; //  728 : 255 - 0xff -- Sprite 0x5b
      12'h2D9: dout  = 8'b00000000; //  729 :   0 - 0x0
      12'h2DA: dout  = 8'b11000011; //  730 : 195 - 0xc3
      12'h2DB: dout  = 8'b10000001; //  731 : 129 - 0x81
      12'h2DC: dout  = 8'b10000001; //  732 : 129 - 0x81
      12'h2DD: dout  = 8'b11000011; //  733 : 195 - 0xc3
      12'h2DE: dout  = 8'b11111111; //  734 : 255 - 0xff
      12'h2DF: dout  = 8'b00000000; //  735 :   0 - 0x0
      12'h2E0: dout  = 8'b00000000; //  736 :   0 - 0x0 -- Sprite 0x5c
      12'h2E1: dout  = 8'b00000000; //  737 :   0 - 0x0
      12'h2E2: dout  = 8'b00000000; //  738 :   0 - 0x0
      12'h2E3: dout  = 8'b00000000; //  739 :   0 - 0x0
      12'h2E4: dout  = 8'b00000000; //  740 :   0 - 0x0
      12'h2E5: dout  = 8'b00000000; //  741 :   0 - 0x0
      12'h2E6: dout  = 8'b00000000; //  742 :   0 - 0x0
      12'h2E7: dout  = 8'b00000000; //  743 :   0 - 0x0
      12'h2E8: dout  = 8'b00000000; //  744 :   0 - 0x0 -- Sprite 0x5d
      12'h2E9: dout  = 8'b00001011; //  745 :  11 - 0xb
      12'h2EA: dout  = 8'b00011111; //  746 :  31 - 0x1f
      12'h2EB: dout  = 8'b00011111; //  747 :  31 - 0x1f
      12'h2EC: dout  = 8'b00011110; //  748 :  30 - 0x1e
      12'h2ED: dout  = 8'b00111110; //  749 :  62 - 0x3e
      12'h2EE: dout  = 8'b00001100; //  750 :  12 - 0xc
      12'h2EF: dout  = 8'b00000100; //  751 :   4 - 0x4
      12'h2F0: dout  = 8'b00000000; //  752 :   0 - 0x0 -- Sprite 0x5e
      12'h2F1: dout  = 8'b00000000; //  753 :   0 - 0x0
      12'h2F2: dout  = 8'b00000000; //  754 :   0 - 0x0
      12'h2F3: dout  = 8'b00000000; //  755 :   0 - 0x0
      12'h2F4: dout  = 8'b00000000; //  756 :   0 - 0x0
      12'h2F5: dout  = 8'b00000000; //  757 :   0 - 0x0
      12'h2F6: dout  = 8'b00000000; //  758 :   0 - 0x0
      12'h2F7: dout  = 8'b00000000; //  759 :   0 - 0x0
      12'h2F8: dout  = 8'b00000011; //  760 :   3 - 0x3 -- Sprite 0x5f
      12'h2F9: dout  = 8'b00001111; //  761 :  15 - 0xf
      12'h2FA: dout  = 8'b00001111; //  762 :  15 - 0xf
      12'h2FB: dout  = 8'b00001111; //  763 :  15 - 0xf
      12'h2FC: dout  = 8'b00001111; //  764 :  15 - 0xf
      12'h2FD: dout  = 8'b00000000; //  765 :   0 - 0x0
      12'h2FE: dout  = 8'b00000000; //  766 :   0 - 0x0
      12'h2FF: dout  = 8'b00000000; //  767 :   0 - 0x0
      12'h300: dout  = 8'b00000000; //  768 :   0 - 0x0 -- Sprite 0x60
      12'h301: dout  = 8'b00011000; //  769 :  24 - 0x18
      12'h302: dout  = 8'b00111100; //  770 :  60 - 0x3c
      12'h303: dout  = 8'b01111110; //  771 : 126 - 0x7e
      12'h304: dout  = 8'b01110110; //  772 : 118 - 0x76
      12'h305: dout  = 8'b11111011; //  773 : 251 - 0xfb
      12'h306: dout  = 8'b11111011; //  774 : 251 - 0xfb
      12'h307: dout  = 8'b11111011; //  775 : 251 - 0xfb
      12'h308: dout  = 8'b00000000; //  776 :   0 - 0x0 -- Sprite 0x61
      12'h309: dout  = 8'b00010000; //  777 :  16 - 0x10
      12'h30A: dout  = 8'b00010000; //  778 :  16 - 0x10
      12'h30B: dout  = 8'b00100000; //  779 :  32 - 0x20
      12'h30C: dout  = 8'b00100000; //  780 :  32 - 0x20
      12'h30D: dout  = 8'b00100000; //  781 :  32 - 0x20
      12'h30E: dout  = 8'b00100000; //  782 :  32 - 0x20
      12'h30F: dout  = 8'b00100000; //  783 :  32 - 0x20
      12'h310: dout  = 8'b00000000; //  784 :   0 - 0x0 -- Sprite 0x62
      12'h311: dout  = 8'b00001000; //  785 :   8 - 0x8
      12'h312: dout  = 8'b00001000; //  786 :   8 - 0x8
      12'h313: dout  = 8'b00001000; //  787 :   8 - 0x8
      12'h314: dout  = 8'b00001000; //  788 :   8 - 0x8
      12'h315: dout  = 8'b00001000; //  789 :   8 - 0x8
      12'h316: dout  = 8'b00001000; //  790 :   8 - 0x8
      12'h317: dout  = 8'b00001000; //  791 :   8 - 0x8
      12'h318: dout  = 8'b00000000; //  792 :   0 - 0x0 -- Sprite 0x63
      12'h319: dout  = 8'b00010000; //  793 :  16 - 0x10
      12'h31A: dout  = 8'b00010000; //  794 :  16 - 0x10
      12'h31B: dout  = 8'b00111000; //  795 :  56 - 0x38
      12'h31C: dout  = 8'b00111000; //  796 :  56 - 0x38
      12'h31D: dout  = 8'b00111000; //  797 :  56 - 0x38
      12'h31E: dout  = 8'b00111000; //  798 :  56 - 0x38
      12'h31F: dout  = 8'b00111000; //  799 :  56 - 0x38
      12'h320: dout  = 8'b00000000; //  800 :   0 - 0x0 -- Sprite 0x64
      12'h321: dout  = 8'b00011000; //  801 :  24 - 0x18
      12'h322: dout  = 8'b00111100; //  802 :  60 - 0x3c
      12'h323: dout  = 8'b00001110; //  803 :  14 - 0xe
      12'h324: dout  = 8'b00001110; //  804 :  14 - 0xe
      12'h325: dout  = 8'b00000100; //  805 :   4 - 0x4
      12'h326: dout  = 8'b00000000; //  806 :   0 - 0x0
      12'h327: dout  = 8'b00000000; //  807 :   0 - 0x0
      12'h328: dout  = 8'b00000000; //  808 :   0 - 0x0 -- Sprite 0x65
      12'h329: dout  = 8'b00000000; //  809 :   0 - 0x0
      12'h32A: dout  = 8'b00000100; //  810 :   4 - 0x4
      12'h32B: dout  = 8'b00000110; //  811 :   6 - 0x6
      12'h32C: dout  = 8'b00011110; //  812 :  30 - 0x1e
      12'h32D: dout  = 8'b00111100; //  813 :  60 - 0x3c
      12'h32E: dout  = 8'b00011000; //  814 :  24 - 0x18
      12'h32F: dout  = 8'b00000000; //  815 :   0 - 0x0
      12'h330: dout  = 8'b00000000; //  816 :   0 - 0x0 -- Sprite 0x66
      12'h331: dout  = 8'b00000000; //  817 :   0 - 0x0
      12'h332: dout  = 8'b00000001; //  818 :   1 - 0x1
      12'h333: dout  = 8'b00001010; //  819 :  10 - 0xa
      12'h334: dout  = 8'b00010111; //  820 :  23 - 0x17
      12'h335: dout  = 8'b00001111; //  821 :  15 - 0xf
      12'h336: dout  = 8'b00101111; //  822 :  47 - 0x2f
      12'h337: dout  = 8'b00011111; //  823 :  31 - 0x1f
      12'h338: dout  = 8'b00000000; //  824 :   0 - 0x0 -- Sprite 0x67
      12'h339: dout  = 8'b00000000; //  825 :   0 - 0x0
      12'h33A: dout  = 8'b00000000; //  826 :   0 - 0x0
      12'h33B: dout  = 8'b00000000; //  827 :   0 - 0x0
      12'h33C: dout  = 8'b00000101; //  828 :   5 - 0x5
      12'h33D: dout  = 8'b00000111; //  829 :   7 - 0x7
      12'h33E: dout  = 8'b00001111; //  830 :  15 - 0xf
      12'h33F: dout  = 8'b00000111; //  831 :   7 - 0x7
      12'h340: dout  = 8'b00000000; //  832 :   0 - 0x0 -- Sprite 0x68
      12'h341: dout  = 8'b00000000; //  833 :   0 - 0x0
      12'h342: dout  = 8'b00000000; //  834 :   0 - 0x0
      12'h343: dout  = 8'b00000000; //  835 :   0 - 0x0
      12'h344: dout  = 8'b00000000; //  836 :   0 - 0x0
      12'h345: dout  = 8'b00000000; //  837 :   0 - 0x0
      12'h346: dout  = 8'b00000001; //  838 :   1 - 0x1
      12'h347: dout  = 8'b00000011; //  839 :   3 - 0x3
      12'h348: dout  = 8'b00000000; //  840 :   0 - 0x0 -- Sprite 0x69
      12'h349: dout  = 8'b01100000; //  841 :  96 - 0x60
      12'h34A: dout  = 8'b11110000; //  842 : 240 - 0xf0
      12'h34B: dout  = 8'b11111000; //  843 : 248 - 0xf8
      12'h34C: dout  = 8'b01111100; //  844 : 124 - 0x7c
      12'h34D: dout  = 8'b00111110; //  845 :  62 - 0x3e
      12'h34E: dout  = 8'b01111110; //  846 : 126 - 0x7e
      12'h34F: dout  = 8'b01111111; //  847 : 127 - 0x7f
      12'h350: dout  = 8'b00111111; //  848 :  63 - 0x3f -- Sprite 0x6a
      12'h351: dout  = 8'b01011111; //  849 :  95 - 0x5f
      12'h352: dout  = 8'b01111111; //  850 : 127 - 0x7f
      12'h353: dout  = 8'b00111110; //  851 :  62 - 0x3e
      12'h354: dout  = 8'b00001110; //  852 :  14 - 0xe
      12'h355: dout  = 8'b00001010; //  853 :  10 - 0xa
      12'h356: dout  = 8'b01010001; //  854 :  81 - 0x51
      12'h357: dout  = 8'b00100000; //  855 :  32 - 0x20
      12'h358: dout  = 8'b00000000; //  856 :   0 - 0x0 -- Sprite 0x6b
      12'h359: dout  = 8'b00000000; //  857 :   0 - 0x0
      12'h35A: dout  = 8'b00000000; //  858 :   0 - 0x0
      12'h35B: dout  = 8'b00000000; //  859 :   0 - 0x0
      12'h35C: dout  = 8'b00000000; //  860 :   0 - 0x0
      12'h35D: dout  = 8'b00000000; //  861 :   0 - 0x0
      12'h35E: dout  = 8'b00001110; //  862 :  14 - 0xe
      12'h35F: dout  = 8'b00011111; //  863 :  31 - 0x1f
      12'h360: dout  = 8'b00111111; //  864 :  63 - 0x3f -- Sprite 0x6c
      12'h361: dout  = 8'b01111111; //  865 : 127 - 0x7f
      12'h362: dout  = 8'b01111111; //  866 : 127 - 0x7f
      12'h363: dout  = 8'b11111110; //  867 : 254 - 0xfe
      12'h364: dout  = 8'b11101100; //  868 : 236 - 0xec
      12'h365: dout  = 8'b11001010; //  869 : 202 - 0xca
      12'h366: dout  = 8'b01010001; //  870 :  81 - 0x51
      12'h367: dout  = 8'b00100000; //  871 :  32 - 0x20
      12'h368: dout  = 8'b00000000; //  872 :   0 - 0x0 -- Sprite 0x6d
      12'h369: dout  = 8'b01000000; //  873 :  64 - 0x40
      12'h36A: dout  = 8'b01100011; //  874 :  99 - 0x63
      12'h36B: dout  = 8'b01110111; //  875 : 119 - 0x77
      12'h36C: dout  = 8'b01111100; //  876 : 124 - 0x7c
      12'h36D: dout  = 8'b00111000; //  877 :  56 - 0x38
      12'h36E: dout  = 8'b11111000; //  878 : 248 - 0xf8
      12'h36F: dout  = 8'b11100100; //  879 : 228 - 0xe4
      12'h370: dout  = 8'b00000000; //  880 :   0 - 0x0 -- Sprite 0x6e
      12'h371: dout  = 8'b00000000; //  881 :   0 - 0x0
      12'h372: dout  = 8'b00000011; //  882 :   3 - 0x3
      12'h373: dout  = 8'b00000111; //  883 :   7 - 0x7
      12'h374: dout  = 8'b00001100; //  884 :  12 - 0xc
      12'h375: dout  = 8'b00011000; //  885 :  24 - 0x18
      12'h376: dout  = 8'b11111000; //  886 : 248 - 0xf8
      12'h377: dout  = 8'b11100100; //  887 : 228 - 0xe4
      12'h378: dout  = 8'b00000011; //  888 :   3 - 0x3 -- Sprite 0x6f
      12'h379: dout  = 8'b01000100; //  889 :  68 - 0x44
      12'h37A: dout  = 8'b00101000; //  890 :  40 - 0x28
      12'h37B: dout  = 8'b00010000; //  891 :  16 - 0x10
      12'h37C: dout  = 8'b00001000; //  892 :   8 - 0x8
      12'h37D: dout  = 8'b00000100; //  893 :   4 - 0x4
      12'h37E: dout  = 8'b00000011; //  894 :   3 - 0x3
      12'h37F: dout  = 8'b00000100; //  895 :   4 - 0x4
      12'h380: dout  = 8'b00000011; //  896 :   3 - 0x3 -- Sprite 0x70
      12'h381: dout  = 8'b00000111; //  897 :   7 - 0x7
      12'h382: dout  = 8'b00001111; //  898 :  15 - 0xf
      12'h383: dout  = 8'b00011111; //  899 :  31 - 0x1f
      12'h384: dout  = 8'b00100111; //  900 :  39 - 0x27
      12'h385: dout  = 8'b01111011; //  901 : 123 - 0x7b
      12'h386: dout  = 8'b01111000; //  902 : 120 - 0x78
      12'h387: dout  = 8'b11111011; //  903 : 251 - 0xfb
      12'h388: dout  = 8'b11000000; //  904 : 192 - 0xc0 -- Sprite 0x71
      12'h389: dout  = 8'b11100000; //  905 : 224 - 0xe0
      12'h38A: dout  = 8'b11110000; //  906 : 240 - 0xf0
      12'h38B: dout  = 8'b11111000; //  907 : 248 - 0xf8
      12'h38C: dout  = 8'b11100100; //  908 : 228 - 0xe4
      12'h38D: dout  = 8'b11011110; //  909 : 222 - 0xde
      12'h38E: dout  = 8'b00011110; //  910 :  30 - 0x1e
      12'h38F: dout  = 8'b11011111; //  911 : 223 - 0xdf
      12'h390: dout  = 8'b11111111; //  912 : 255 - 0xff -- Sprite 0x72
      12'h391: dout  = 8'b11111111; //  913 : 255 - 0xff
      12'h392: dout  = 8'b01111111; //  914 : 127 - 0x7f
      12'h393: dout  = 8'b00001111; //  915 :  15 - 0xf
      12'h394: dout  = 8'b00001111; //  916 :  15 - 0xf
      12'h395: dout  = 8'b00000111; //  917 :   7 - 0x7
      12'h396: dout  = 8'b00000011; //  918 :   3 - 0x3
      12'h397: dout  = 8'b00000000; //  919 :   0 - 0x0
      12'h398: dout  = 8'b11111111; //  920 : 255 - 0xff -- Sprite 0x73
      12'h399: dout  = 8'b11111111; //  921 : 255 - 0xff
      12'h39A: dout  = 8'b11111110; //  922 : 254 - 0xfe
      12'h39B: dout  = 8'b11110000; //  923 : 240 - 0xf0
      12'h39C: dout  = 8'b11110000; //  924 : 240 - 0xf0
      12'h39D: dout  = 8'b11000000; //  925 : 192 - 0xc0
      12'h39E: dout  = 8'b10000000; //  926 : 128 - 0x80
      12'h39F: dout  = 8'b00000000; //  927 :   0 - 0x0
      12'h3A0: dout  = 8'b00000000; //  928 :   0 - 0x0 -- Sprite 0x74
      12'h3A1: dout  = 8'b00000000; //  929 :   0 - 0x0
      12'h3A2: dout  = 8'b00011000; //  930 :  24 - 0x18
      12'h3A3: dout  = 8'b00100100; //  931 :  36 - 0x24
      12'h3A4: dout  = 8'b00100100; //  932 :  36 - 0x24
      12'h3A5: dout  = 8'b00011000; //  933 :  24 - 0x18
      12'h3A6: dout  = 8'b00000000; //  934 :   0 - 0x0
      12'h3A7: dout  = 8'b00000000; //  935 :   0 - 0x0
      12'h3A8: dout  = 8'b00111100; //  936 :  60 - 0x3c -- Sprite 0x75
      12'h3A9: dout  = 8'b01111110; //  937 : 126 - 0x7e
      12'h3AA: dout  = 8'b11111111; //  938 : 255 - 0xff
      12'h3AB: dout  = 8'b11111111; //  939 : 255 - 0xff
      12'h3AC: dout  = 8'b11111111; //  940 : 255 - 0xff
      12'h3AD: dout  = 8'b11111111; //  941 : 255 - 0xff
      12'h3AE: dout  = 8'b01111110; //  942 : 126 - 0x7e
      12'h3AF: dout  = 8'b00111100; //  943 :  60 - 0x3c
      12'h3B0: dout  = 8'b00000011; //  944 :   3 - 0x3 -- Sprite 0x76
      12'h3B1: dout  = 8'b00000111; //  945 :   7 - 0x7
      12'h3B2: dout  = 8'b00001111; //  946 :  15 - 0xf
      12'h3B3: dout  = 8'b00011111; //  947 :  31 - 0x1f
      12'h3B4: dout  = 8'b00111111; //  948 :  63 - 0x3f
      12'h3B5: dout  = 8'b01100011; //  949 :  99 - 0x63
      12'h3B6: dout  = 8'b01000001; //  950 :  65 - 0x41
      12'h3B7: dout  = 8'b11000001; //  951 : 193 - 0xc1
      12'h3B8: dout  = 8'b11000000; //  952 : 192 - 0xc0 -- Sprite 0x77
      12'h3B9: dout  = 8'b10000000; //  953 : 128 - 0x80
      12'h3BA: dout  = 8'b00000000; //  954 :   0 - 0x0
      12'h3BB: dout  = 8'b00000000; //  955 :   0 - 0x0
      12'h3BC: dout  = 8'b10001100; //  956 : 140 - 0x8c
      12'h3BD: dout  = 8'b11111110; //  957 : 254 - 0xfe
      12'h3BE: dout  = 8'b11111110; //  958 : 254 - 0xfe
      12'h3BF: dout  = 8'b11110011; //  959 : 243 - 0xf3
      12'h3C0: dout  = 8'b11000001; //  960 : 193 - 0xc1 -- Sprite 0x78
      12'h3C1: dout  = 8'b11100011; //  961 : 227 - 0xe3
      12'h3C2: dout  = 8'b11111111; //  962 : 255 - 0xff
      12'h3C3: dout  = 8'b01000111; //  963 :  71 - 0x47
      12'h3C4: dout  = 8'b00001111; //  964 :  15 - 0xf
      12'h3C5: dout  = 8'b00001111; //  965 :  15 - 0xf
      12'h3C6: dout  = 8'b00001111; //  966 :  15 - 0xf
      12'h3C7: dout  = 8'b00000111; //  967 :   7 - 0x7
      12'h3C8: dout  = 8'b11110001; //  968 : 241 - 0xf1 -- Sprite 0x79
      12'h3C9: dout  = 8'b11111001; //  969 : 249 - 0xf9
      12'h3CA: dout  = 8'b11111111; //  970 : 255 - 0xff
      12'h3CB: dout  = 8'b11100010; //  971 : 226 - 0xe2
      12'h3CC: dout  = 8'b11110000; //  972 : 240 - 0xf0
      12'h3CD: dout  = 8'b11110000; //  973 : 240 - 0xf0
      12'h3CE: dout  = 8'b11110000; //  974 : 240 - 0xf0
      12'h3CF: dout  = 8'b11100000; //  975 : 224 - 0xe0
      12'h3D0: dout  = 8'b00010110; //  976 :  22 - 0x16 -- Sprite 0x7a
      12'h3D1: dout  = 8'b00011111; //  977 :  31 - 0x1f
      12'h3D2: dout  = 8'b00000000; //  978 :   0 - 0x0
      12'h3D3: dout  = 8'b00000000; //  979 :   0 - 0x0
      12'h3D4: dout  = 8'b00000101; //  980 :   5 - 0x5
      12'h3D5: dout  = 8'b00001101; //  981 :  13 - 0xd
      12'h3D6: dout  = 8'b00111111; //  982 :  63 - 0x3f
      12'h3D7: dout  = 8'b00011111; //  983 :  31 - 0x1f
      12'h3D8: dout  = 8'b10000000; //  984 : 128 - 0x80 -- Sprite 0x7b
      12'h3D9: dout  = 8'b10000000; //  985 : 128 - 0x80
      12'h3DA: dout  = 8'b00000000; //  986 :   0 - 0x0
      12'h3DB: dout  = 8'b00000000; //  987 :   0 - 0x0
      12'h3DC: dout  = 8'b00000000; //  988 :   0 - 0x0
      12'h3DD: dout  = 8'b10100000; //  989 : 160 - 0xa0
      12'h3DE: dout  = 8'b10100000; //  990 : 160 - 0xa0
      12'h3DF: dout  = 8'b11100000; //  991 : 224 - 0xe0
      12'h3E0: dout  = 8'b00000000; //  992 :   0 - 0x0 -- Sprite 0x7c
      12'h3E1: dout  = 8'b00000100; //  993 :   4 - 0x4
      12'h3E2: dout  = 8'b01001110; //  994 :  78 - 0x4e
      12'h3E3: dout  = 8'b10001100; //  995 : 140 - 0x8c
      12'h3E4: dout  = 8'b00001100; //  996 :  12 - 0xc
      12'h3E5: dout  = 8'b01111111; //  997 : 127 - 0x7f
      12'h3E6: dout  = 8'b11111111; //  998 : 255 - 0xff
      12'h3E7: dout  = 8'b11111111; //  999 : 255 - 0xff
      12'h3E8: dout  = 8'b00000000; // 1000 :   0 - 0x0 -- Sprite 0x7d
      12'h3E9: dout  = 8'b00000000; // 1001 :   0 - 0x0
      12'h3EA: dout  = 8'b00000000; // 1002 :   0 - 0x0
      12'h3EB: dout  = 8'b00000000; // 1003 :   0 - 0x0
      12'h3EC: dout  = 8'b00000000; // 1004 :   0 - 0x0
      12'h3ED: dout  = 8'b00000000; // 1005 :   0 - 0x0
      12'h3EE: dout  = 8'b00000001; // 1006 :   1 - 0x1
      12'h3EF: dout  = 8'b00000001; // 1007 :   1 - 0x1
      12'h3F0: dout  = 8'b11111111; // 1008 : 255 - 0xff -- Sprite 0x7e
      12'h3F1: dout  = 8'b01111111; // 1009 : 127 - 0x7f
      12'h3F2: dout  = 8'b00111111; // 1010 :  63 - 0x3f
      12'h3F3: dout  = 8'b00011111; // 1011 :  31 - 0x1f
      12'h3F4: dout  = 8'b00001111; // 1012 :  15 - 0xf
      12'h3F5: dout  = 8'b00000111; // 1013 :   7 - 0x7
      12'h3F6: dout  = 8'b00000011; // 1014 :   3 - 0x3
      12'h3F7: dout  = 8'b00000001; // 1015 :   1 - 0x1
      12'h3F8: dout  = 8'b11111111; // 1016 : 255 - 0xff -- Sprite 0x7f
      12'h3F9: dout  = 8'b10000011; // 1017 : 131 - 0x83
      12'h3FA: dout  = 8'b00101001; // 1018 :  41 - 0x29
      12'h3FB: dout  = 8'b01101101; // 1019 : 109 - 0x6d
      12'h3FC: dout  = 8'b01000101; // 1020 :  69 - 0x45
      12'h3FD: dout  = 8'b00010001; // 1021 :  17 - 0x11
      12'h3FE: dout  = 8'b00000001; // 1022 :   1 - 0x1
      12'h3FF: dout  = 8'b11000111; // 1023 : 199 - 0xc7
      12'h400: dout  = 8'b00001000; // 1024 :   8 - 0x8 -- Sprite 0x80
      12'h401: dout  = 8'b00001000; // 1025 :   8 - 0x8
      12'h402: dout  = 8'b00000010; // 1026 :   2 - 0x2
      12'h403: dout  = 8'b00011111; // 1027 :  31 - 0x1f
      12'h404: dout  = 8'b00100010; // 1028 :  34 - 0x22
      12'h405: dout  = 8'b00000010; // 1029 :   2 - 0x2
      12'h406: dout  = 8'b00000010; // 1030 :   2 - 0x2
      12'h407: dout  = 8'b00000000; // 1031 :   0 - 0x0
      12'h408: dout  = 8'b00001000; // 1032 :   8 - 0x8 -- Sprite 0x81
      12'h409: dout  = 8'b00001000; // 1033 :   8 - 0x8
      12'h40A: dout  = 8'b00001000; // 1034 :   8 - 0x8
      12'h40B: dout  = 8'b00001000; // 1035 :   8 - 0x8
      12'h40C: dout  = 8'b00001000; // 1036 :   8 - 0x8
      12'h40D: dout  = 8'b00001000; // 1037 :   8 - 0x8
      12'h40E: dout  = 8'b00001000; // 1038 :   8 - 0x8
      12'h40F: dout  = 8'b00001000; // 1039 :   8 - 0x8
      12'h410: dout  = 8'b00010000; // 1040 :  16 - 0x10 -- Sprite 0x82
      12'h411: dout  = 8'b00011110; // 1041 :  30 - 0x1e
      12'h412: dout  = 8'b00010000; // 1042 :  16 - 0x10
      12'h413: dout  = 8'b01010000; // 1043 :  80 - 0x50
      12'h414: dout  = 8'b00010000; // 1044 :  16 - 0x10
      12'h415: dout  = 8'b00001000; // 1045 :   8 - 0x8
      12'h416: dout  = 8'b00000000; // 1046 :   0 - 0x0
      12'h417: dout  = 8'b00000000; // 1047 :   0 - 0x0
      12'h418: dout  = 8'b00000000; // 1048 :   0 - 0x0 -- Sprite 0x83
      12'h419: dout  = 8'b00000000; // 1049 :   0 - 0x0
      12'h41A: dout  = 8'b00000000; // 1050 :   0 - 0x0
      12'h41B: dout  = 8'b11111110; // 1051 : 254 - 0xfe
      12'h41C: dout  = 8'b00000000; // 1052 :   0 - 0x0
      12'h41D: dout  = 8'b00000000; // 1053 :   0 - 0x0
      12'h41E: dout  = 8'b00000000; // 1054 :   0 - 0x0
      12'h41F: dout  = 8'b00000000; // 1055 :   0 - 0x0
      12'h420: dout  = 8'b00011100; // 1056 :  28 - 0x1c -- Sprite 0x84
      12'h421: dout  = 8'b00101010; // 1057 :  42 - 0x2a
      12'h422: dout  = 8'b01110111; // 1058 : 119 - 0x77
      12'h423: dout  = 8'b11101110; // 1059 : 238 - 0xee
      12'h424: dout  = 8'b11011101; // 1060 : 221 - 0xdd
      12'h425: dout  = 8'b10101010; // 1061 : 170 - 0xaa
      12'h426: dout  = 8'b01110100; // 1062 : 116 - 0x74
      12'h427: dout  = 8'b00101000; // 1063 :  40 - 0x28
      12'h428: dout  = 8'b11111111; // 1064 : 255 - 0xff -- Sprite 0x85
      12'h429: dout  = 8'b11111110; // 1065 : 254 - 0xfe
      12'h42A: dout  = 8'b11111110; // 1066 : 254 - 0xfe
      12'h42B: dout  = 8'b00000000; // 1067 :   0 - 0x0
      12'h42C: dout  = 8'b11101111; // 1068 : 239 - 0xef
      12'h42D: dout  = 8'b11101111; // 1069 : 239 - 0xef
      12'h42E: dout  = 8'b11101111; // 1070 : 239 - 0xef
      12'h42F: dout  = 8'b00000000; // 1071 :   0 - 0x0
      12'h430: dout  = 8'b11111110; // 1072 : 254 - 0xfe -- Sprite 0x86
      12'h431: dout  = 8'b11111110; // 1073 : 254 - 0xfe
      12'h432: dout  = 8'b11111110; // 1074 : 254 - 0xfe
      12'h433: dout  = 8'b00000000; // 1075 :   0 - 0x0
      12'h434: dout  = 8'b11101111; // 1076 : 239 - 0xef
      12'h435: dout  = 8'b11101111; // 1077 : 239 - 0xef
      12'h436: dout  = 8'b11101111; // 1078 : 239 - 0xef
      12'h437: dout  = 8'b00000000; // 1079 :   0 - 0x0
      12'h438: dout  = 8'b00000000; // 1080 :   0 - 0x0 -- Sprite 0x87
      12'h439: dout  = 8'b01111111; // 1081 : 127 - 0x7f
      12'h43A: dout  = 8'b01011111; // 1082 :  95 - 0x5f
      12'h43B: dout  = 8'b01111111; // 1083 : 127 - 0x7f
      12'h43C: dout  = 8'b01111111; // 1084 : 127 - 0x7f
      12'h43D: dout  = 8'b01111111; // 1085 : 127 - 0x7f
      12'h43E: dout  = 8'b01111111; // 1086 : 127 - 0x7f
      12'h43F: dout  = 8'b01111111; // 1087 : 127 - 0x7f
      12'h440: dout  = 8'b10111000; // 1088 : 184 - 0xb8 -- Sprite 0x88
      12'h441: dout  = 8'b10011110; // 1089 : 158 - 0x9e
      12'h442: dout  = 8'b10000000; // 1090 : 128 - 0x80
      12'h443: dout  = 8'b11000000; // 1091 : 192 - 0xc0
      12'h444: dout  = 8'b11100000; // 1092 : 224 - 0xe0
      12'h445: dout  = 8'b11110000; // 1093 : 240 - 0xf0
      12'h446: dout  = 8'b11111000; // 1094 : 248 - 0xf8
      12'h447: dout  = 8'b01111100; // 1095 : 124 - 0x7c
      12'h448: dout  = 8'b00000000; // 1096 :   0 - 0x0 -- Sprite 0x89
      12'h449: dout  = 8'b00100011; // 1097 :  35 - 0x23
      12'h44A: dout  = 8'b01010111; // 1098 :  87 - 0x57
      12'h44B: dout  = 8'b01001111; // 1099 :  79 - 0x4f
      12'h44C: dout  = 8'b01010111; // 1100 :  87 - 0x57
      12'h44D: dout  = 8'b00100111; // 1101 :  39 - 0x27
      12'h44E: dout  = 8'b11000011; // 1102 : 195 - 0xc3
      12'h44F: dout  = 8'b00100001; // 1103 :  33 - 0x21
      12'h450: dout  = 8'b00000000; // 1104 :   0 - 0x0 -- Sprite 0x8a
      12'h451: dout  = 8'b00110000; // 1105 :  48 - 0x30
      12'h452: dout  = 8'b01110000; // 1106 : 112 - 0x70
      12'h453: dout  = 8'b01110000; // 1107 : 112 - 0x70
      12'h454: dout  = 8'b11110000; // 1108 : 240 - 0xf0
      12'h455: dout  = 8'b11100000; // 1109 : 224 - 0xe0
      12'h456: dout  = 8'b11000000; // 1110 : 192 - 0xc0
      12'h457: dout  = 8'b00000000; // 1111 :   0 - 0x0
      12'h458: dout  = 8'b00010011; // 1112 :  19 - 0x13 -- Sprite 0x8b
      12'h459: dout  = 8'b00001111; // 1113 :  15 - 0xf
      12'h45A: dout  = 8'b00011110; // 1114 :  30 - 0x1e
      12'h45B: dout  = 8'b11110000; // 1115 : 240 - 0xf0
      12'h45C: dout  = 8'b11111100; // 1116 : 252 - 0xfc
      12'h45D: dout  = 8'b11111000; // 1117 : 248 - 0xf8
      12'h45E: dout  = 8'b11110000; // 1118 : 240 - 0xf0
      12'h45F: dout  = 8'b11100000; // 1119 : 224 - 0xe0
      12'h460: dout  = 8'b10111110; // 1120 : 190 - 0xbe -- Sprite 0x8c
      12'h461: dout  = 8'b10010000; // 1121 : 144 - 0x90
      12'h462: dout  = 8'b10000000; // 1122 : 128 - 0x80
      12'h463: dout  = 8'b11000000; // 1123 : 192 - 0xc0
      12'h464: dout  = 8'b11000000; // 1124 : 192 - 0xc0
      12'h465: dout  = 8'b10000000; // 1125 : 128 - 0x80
      12'h466: dout  = 8'b00000000; // 1126 :   0 - 0x0
      12'h467: dout  = 8'b00000000; // 1127 :   0 - 0x0
      12'h468: dout  = 8'b00000001; // 1128 :   1 - 0x1 -- Sprite 0x8d
      12'h469: dout  = 8'b00000001; // 1129 :   1 - 0x1
      12'h46A: dout  = 8'b00000011; // 1130 :   3 - 0x3
      12'h46B: dout  = 8'b00000011; // 1131 :   3 - 0x3
      12'h46C: dout  = 8'b00000111; // 1132 :   7 - 0x7
      12'h46D: dout  = 8'b01111111; // 1133 : 127 - 0x7f
      12'h46E: dout  = 8'b01111101; // 1134 : 125 - 0x7d
      12'h46F: dout  = 8'b00111101; // 1135 :  61 - 0x3d
      12'h470: dout  = 8'b00000110; // 1136 :   6 - 0x6 -- Sprite 0x8e
      12'h471: dout  = 8'b00000100; // 1137 :   4 - 0x4
      12'h472: dout  = 8'b00110000; // 1138 :  48 - 0x30
      12'h473: dout  = 8'b00100011; // 1139 :  35 - 0x23
      12'h474: dout  = 8'b00000110; // 1140 :   6 - 0x6
      12'h475: dout  = 8'b01100100; // 1141 : 100 - 0x64
      12'h476: dout  = 8'b01100000; // 1142 :  96 - 0x60
      12'h477: dout  = 8'b00000000; // 1143 :   0 - 0x0
      12'h478: dout  = 8'b00000000; // 1144 :   0 - 0x0 -- Sprite 0x8f
      12'h479: dout  = 8'b01100000; // 1145 :  96 - 0x60
      12'h47A: dout  = 8'b01100000; // 1146 :  96 - 0x60
      12'h47B: dout  = 8'b00000000; // 1147 :   0 - 0x0
      12'h47C: dout  = 8'b00100000; // 1148 :  32 - 0x20
      12'h47D: dout  = 8'b00110000; // 1149 :  48 - 0x30
      12'h47E: dout  = 8'b00000100; // 1150 :   4 - 0x4
      12'h47F: dout  = 8'b00000110; // 1151 :   6 - 0x6
      12'h480: dout  = 8'b00000000; // 1152 :   0 - 0x0 -- Sprite 0x90
      12'h481: dout  = 8'b00000001; // 1153 :   1 - 0x1
      12'h482: dout  = 8'b00000001; // 1154 :   1 - 0x1
      12'h483: dout  = 8'b00000000; // 1155 :   0 - 0x0
      12'h484: dout  = 8'b00000000; // 1156 :   0 - 0x0
      12'h485: dout  = 8'b00000000; // 1157 :   0 - 0x0
      12'h486: dout  = 8'b00000000; // 1158 :   0 - 0x0
      12'h487: dout  = 8'b00000000; // 1159 :   0 - 0x0
      12'h488: dout  = 8'b11111110; // 1160 : 254 - 0xfe -- Sprite 0x91
      12'h489: dout  = 8'b11111111; // 1161 : 255 - 0xff
      12'h48A: dout  = 8'b11111111; // 1162 : 255 - 0xff
      12'h48B: dout  = 8'b01000000; // 1163 :  64 - 0x40
      12'h48C: dout  = 8'b00000001; // 1164 :   1 - 0x1
      12'h48D: dout  = 8'b00000011; // 1165 :   3 - 0x3
      12'h48E: dout  = 8'b00000011; // 1166 :   3 - 0x3
      12'h48F: dout  = 8'b00000011; // 1167 :   3 - 0x3
      12'h490: dout  = 8'b00000001; // 1168 :   1 - 0x1 -- Sprite 0x92
      12'h491: dout  = 8'b00000001; // 1169 :   1 - 0x1
      12'h492: dout  = 8'b00000000; // 1170 :   0 - 0x0
      12'h493: dout  = 8'b00000000; // 1171 :   0 - 0x0
      12'h494: dout  = 8'b00000000; // 1172 :   0 - 0x0
      12'h495: dout  = 8'b00000000; // 1173 :   0 - 0x0
      12'h496: dout  = 8'b00000000; // 1174 :   0 - 0x0
      12'h497: dout  = 8'b00000000; // 1175 :   0 - 0x0
      12'h498: dout  = 8'b11100000; // 1176 : 224 - 0xe0 -- Sprite 0x93
      12'h499: dout  = 8'b11111110; // 1177 : 254 - 0xfe
      12'h49A: dout  = 8'b11111111; // 1178 : 255 - 0xff
      12'h49B: dout  = 8'b01111111; // 1179 : 127 - 0x7f
      12'h49C: dout  = 8'b00000011; // 1180 :   3 - 0x3
      12'h49D: dout  = 8'b00000010; // 1181 :   2 - 0x2
      12'h49E: dout  = 8'b00000000; // 1182 :   0 - 0x0
      12'h49F: dout  = 8'b00000000; // 1183 :   0 - 0x0
      12'h4A0: dout  = 8'b00000001; // 1184 :   1 - 0x1 -- Sprite 0x94
      12'h4A1: dout  = 8'b00001101; // 1185 :  13 - 0xd
      12'h4A2: dout  = 8'b00001000; // 1186 :   8 - 0x8
      12'h4A3: dout  = 8'b00000000; // 1187 :   0 - 0x0
      12'h4A4: dout  = 8'b00110110; // 1188 :  54 - 0x36
      12'h4A5: dout  = 8'b00101100; // 1189 :  44 - 0x2c
      12'h4A6: dout  = 8'b00001000; // 1190 :   8 - 0x8
      12'h4A7: dout  = 8'b01100000; // 1191 :  96 - 0x60
      12'h4A8: dout  = 8'b01100000; // 1192 :  96 - 0x60 -- Sprite 0x95
      12'h4A9: dout  = 8'b00000000; // 1193 :   0 - 0x0
      12'h4AA: dout  = 8'b00100000; // 1194 :  32 - 0x20
      12'h4AB: dout  = 8'b00110000; // 1195 :  48 - 0x30
      12'h4AC: dout  = 8'b00000000; // 1196 :   0 - 0x0
      12'h4AD: dout  = 8'b00001000; // 1197 :   8 - 0x8
      12'h4AE: dout  = 8'b00001101; // 1198 :  13 - 0xd
      12'h4AF: dout  = 8'b00000001; // 1199 :   1 - 0x1
      12'h4B0: dout  = 8'b00000001; // 1200 :   1 - 0x1 -- Sprite 0x96
      12'h4B1: dout  = 8'b00000001; // 1201 :   1 - 0x1
      12'h4B2: dout  = 8'b00000011; // 1202 :   3 - 0x3
      12'h4B3: dout  = 8'b01000011; // 1203 :  67 - 0x43
      12'h4B4: dout  = 8'b01100111; // 1204 : 103 - 0x67
      12'h4B5: dout  = 8'b01110111; // 1205 : 119 - 0x77
      12'h4B6: dout  = 8'b01111011; // 1206 : 123 - 0x7b
      12'h4B7: dout  = 8'b01111000; // 1207 : 120 - 0x78
      12'h4B8: dout  = 8'b00000000; // 1208 :   0 - 0x0 -- Sprite 0x97
      12'h4B9: dout  = 8'b00000000; // 1209 :   0 - 0x0
      12'h4BA: dout  = 8'b10000000; // 1210 : 128 - 0x80
      12'h4BB: dout  = 8'b10000100; // 1211 : 132 - 0x84
      12'h4BC: dout  = 8'b11001100; // 1212 : 204 - 0xcc
      12'h4BD: dout  = 8'b11011100; // 1213 : 220 - 0xdc
      12'h4BE: dout  = 8'b10111100; // 1214 : 188 - 0xbc
      12'h4BF: dout  = 8'b00111100; // 1215 :  60 - 0x3c
      12'h4C0: dout  = 8'b00110011; // 1216 :  51 - 0x33 -- Sprite 0x98
      12'h4C1: dout  = 8'b00000111; // 1217 :   7 - 0x7
      12'h4C2: dout  = 8'b00000111; // 1218 :   7 - 0x7
      12'h4C3: dout  = 8'b11100011; // 1219 : 227 - 0xe3
      12'h4C4: dout  = 8'b00111000; // 1220 :  56 - 0x38
      12'h4C5: dout  = 8'b00111111; // 1221 :  63 - 0x3f
      12'h4C6: dout  = 8'b00011100; // 1222 :  28 - 0x1c
      12'h4C7: dout  = 8'b00001100; // 1223 :  12 - 0xc
      12'h4C8: dout  = 8'b10011000; // 1224 : 152 - 0x98 -- Sprite 0x99
      12'h4C9: dout  = 8'b11000111; // 1225 : 199 - 0xc7
      12'h4CA: dout  = 8'b11001000; // 1226 : 200 - 0xc8
      12'h4CB: dout  = 8'b10010010; // 1227 : 146 - 0x92
      12'h4CC: dout  = 8'b00110000; // 1228 :  48 - 0x30
      12'h4CD: dout  = 8'b11111000; // 1229 : 248 - 0xf8
      12'h4CE: dout  = 8'b01110000; // 1230 : 112 - 0x70
      12'h4CF: dout  = 8'b01100000; // 1231 :  96 - 0x60
      12'h4D0: dout  = 8'b00000000; // 1232 :   0 - 0x0 -- Sprite 0x9a
      12'h4D1: dout  = 8'b00000001; // 1233 :   1 - 0x1
      12'h4D2: dout  = 8'b00000001; // 1234 :   1 - 0x1
      12'h4D3: dout  = 8'b00000011; // 1235 :   3 - 0x3
      12'h4D4: dout  = 8'b01000011; // 1236 :  67 - 0x43
      12'h4D5: dout  = 8'b01100111; // 1237 : 103 - 0x67
      12'h4D6: dout  = 8'b01110111; // 1238 : 119 - 0x77
      12'h4D7: dout  = 8'b01111011; // 1239 : 123 - 0x7b
      12'h4D8: dout  = 8'b00000000; // 1240 :   0 - 0x0 -- Sprite 0x9b
      12'h4D9: dout  = 8'b00000000; // 1241 :   0 - 0x0
      12'h4DA: dout  = 8'b00000000; // 1242 :   0 - 0x0
      12'h4DB: dout  = 8'b10000000; // 1243 : 128 - 0x80
      12'h4DC: dout  = 8'b10000100; // 1244 : 132 - 0x84
      12'h4DD: dout  = 8'b11001100; // 1245 : 204 - 0xcc
      12'h4DE: dout  = 8'b11011100; // 1246 : 220 - 0xdc
      12'h4DF: dout  = 8'b10111100; // 1247 : 188 - 0xbc
      12'h4E0: dout  = 8'b01111000; // 1248 : 120 - 0x78 -- Sprite 0x9c
      12'h4E1: dout  = 8'b00110011; // 1249 :  51 - 0x33
      12'h4E2: dout  = 8'b00000111; // 1250 :   7 - 0x7
      12'h4E3: dout  = 8'b00000111; // 1251 :   7 - 0x7
      12'h4E4: dout  = 8'b11100011; // 1252 : 227 - 0xe3
      12'h4E5: dout  = 8'b00111000; // 1253 :  56 - 0x38
      12'h4E6: dout  = 8'b01111111; // 1254 : 127 - 0x7f
      12'h4E7: dout  = 8'b11110000; // 1255 : 240 - 0xf0
      12'h4E8: dout  = 8'b00111100; // 1256 :  60 - 0x3c -- Sprite 0x9d
      12'h4E9: dout  = 8'b10011000; // 1257 : 152 - 0x98
      12'h4EA: dout  = 8'b11000111; // 1258 : 199 - 0xc7
      12'h4EB: dout  = 8'b11001000; // 1259 : 200 - 0xc8
      12'h4EC: dout  = 8'b10010010; // 1260 : 146 - 0x92
      12'h4ED: dout  = 8'b00110000; // 1261 :  48 - 0x30
      12'h4EE: dout  = 8'b11111000; // 1262 : 248 - 0xf8
      12'h4EF: dout  = 8'b00111100; // 1263 :  60 - 0x3c
      12'h4F0: dout  = 8'b00000000; // 1264 :   0 - 0x0 -- Sprite 0x9e
      12'h4F1: dout  = 8'b00010000; // 1265 :  16 - 0x10
      12'h4F2: dout  = 8'b01111111; // 1266 : 127 - 0x7f
      12'h4F3: dout  = 8'b01111111; // 1267 : 127 - 0x7f
      12'h4F4: dout  = 8'b01111111; // 1268 : 127 - 0x7f
      12'h4F5: dout  = 8'b00011111; // 1269 :  31 - 0x1f
      12'h4F6: dout  = 8'b00001111; // 1270 :  15 - 0xf
      12'h4F7: dout  = 8'b00001111; // 1271 :  15 - 0xf
      12'h4F8: dout  = 8'b00000011; // 1272 :   3 - 0x3 -- Sprite 0x9f
      12'h4F9: dout  = 8'b00110011; // 1273 :  51 - 0x33
      12'h4FA: dout  = 8'b00111001; // 1274 :  57 - 0x39
      12'h4FB: dout  = 8'b00111010; // 1275 :  58 - 0x3a
      12'h4FC: dout  = 8'b00111000; // 1276 :  56 - 0x38
      12'h4FD: dout  = 8'b00011000; // 1277 :  24 - 0x18
      12'h4FE: dout  = 8'b00000000; // 1278 :   0 - 0x0
      12'h4FF: dout  = 8'b00000000; // 1279 :   0 - 0x0
      12'h500: dout  = 8'b00010000; // 1280 :  16 - 0x10 -- Sprite 0xa0
      12'h501: dout  = 8'b00111000; // 1281 :  56 - 0x38
      12'h502: dout  = 8'b00111100; // 1282 :  60 - 0x3c
      12'h503: dout  = 8'b01110100; // 1283 : 116 - 0x74
      12'h504: dout  = 8'b01110110; // 1284 : 118 - 0x76
      12'h505: dout  = 8'b01110110; // 1285 : 118 - 0x76
      12'h506: dout  = 8'b01111110; // 1286 : 126 - 0x7e
      12'h507: dout  = 8'b01111101; // 1287 : 125 - 0x7d
      12'h508: dout  = 8'b00000000; // 1288 :   0 - 0x0 -- Sprite 0xa1
      12'h509: dout  = 8'b00000000; // 1289 :   0 - 0x0
      12'h50A: dout  = 8'b00010001; // 1290 :  17 - 0x11
      12'h50B: dout  = 8'b00001010; // 1291 :  10 - 0xa
      12'h50C: dout  = 8'b00110100; // 1292 :  52 - 0x34
      12'h50D: dout  = 8'b00101010; // 1293 :  42 - 0x2a
      12'h50E: dout  = 8'b01010001; // 1294 :  81 - 0x51
      12'h50F: dout  = 8'b00100000; // 1295 :  32 - 0x20
      12'h510: dout  = 8'b01111111; // 1296 : 127 - 0x7f -- Sprite 0xa2
      12'h511: dout  = 8'b01100111; // 1297 : 103 - 0x67
      12'h512: dout  = 8'b01100011; // 1298 :  99 - 0x63
      12'h513: dout  = 8'b01110000; // 1299 : 112 - 0x70
      12'h514: dout  = 8'b00111000; // 1300 :  56 - 0x38
      12'h515: dout  = 8'b00111110; // 1301 :  62 - 0x3e
      12'h516: dout  = 8'b01111100; // 1302 : 124 - 0x7c
      12'h517: dout  = 8'b10111000; // 1303 : 184 - 0xb8
      12'h518: dout  = 8'b01010001; // 1304 :  81 - 0x51 -- Sprite 0xa3
      12'h519: dout  = 8'b00001010; // 1305 :  10 - 0xa
      12'h51A: dout  = 8'b00000100; // 1306 :   4 - 0x4
      12'h51B: dout  = 8'b11101010; // 1307 : 234 - 0xea
      12'h51C: dout  = 8'b01111001; // 1308 : 121 - 0x79
      12'h51D: dout  = 8'b01111111; // 1309 : 127 - 0x7f
      12'h51E: dout  = 8'b01110000; // 1310 : 112 - 0x70
      12'h51F: dout  = 8'b00111001; // 1311 :  57 - 0x39
      12'h520: dout  = 8'b01011000; // 1312 :  88 - 0x58 -- Sprite 0xa4
      12'h521: dout  = 8'b00111000; // 1313 :  56 - 0x38
      12'h522: dout  = 8'b00010000; // 1314 :  16 - 0x10
      12'h523: dout  = 8'b00110000; // 1315 :  48 - 0x30
      12'h524: dout  = 8'b11110000; // 1316 : 240 - 0xf0
      12'h525: dout  = 8'b11110000; // 1317 : 240 - 0xf0
      12'h526: dout  = 8'b11100000; // 1318 : 224 - 0xe0
      12'h527: dout  = 8'b11000000; // 1319 : 192 - 0xc0
      12'h528: dout  = 8'b00000000; // 1320 :   0 - 0x0 -- Sprite 0xa5
      12'h529: dout  = 8'b00001000; // 1321 :   8 - 0x8
      12'h52A: dout  = 8'b00011100; // 1322 :  28 - 0x1c
      12'h52B: dout  = 8'b00111100; // 1323 :  60 - 0x3c
      12'h52C: dout  = 8'b01111010; // 1324 : 122 - 0x7a
      12'h52D: dout  = 8'b01111010; // 1325 : 122 - 0x7a
      12'h52E: dout  = 8'b01111010; // 1326 : 122 - 0x7a
      12'h52F: dout  = 8'b01111110; // 1327 : 126 - 0x7e
      12'h530: dout  = 8'b00000000; // 1328 :   0 - 0x0 -- Sprite 0xa6
      12'h531: dout  = 8'b00000000; // 1329 :   0 - 0x0
      12'h532: dout  = 8'b00000000; // 1330 :   0 - 0x0
      12'h533: dout  = 8'b00010001; // 1331 :  17 - 0x11
      12'h534: dout  = 8'b00001010; // 1332 :  10 - 0xa
      12'h535: dout  = 8'b00110100; // 1333 :  52 - 0x34
      12'h536: dout  = 8'b00101010; // 1334 :  42 - 0x2a
      12'h537: dout  = 8'b01010001; // 1335 :  81 - 0x51
      12'h538: dout  = 8'b01111111; // 1336 : 127 - 0x7f -- Sprite 0xa7
      12'h539: dout  = 8'b01111101; // 1337 : 125 - 0x7d
      12'h53A: dout  = 8'b00111111; // 1338 :  63 - 0x3f
      12'h53B: dout  = 8'b00110111; // 1339 :  55 - 0x37
      12'h53C: dout  = 8'b00110011; // 1340 :  51 - 0x33
      12'h53D: dout  = 8'b00111011; // 1341 :  59 - 0x3b
      12'h53E: dout  = 8'b00111010; // 1342 :  58 - 0x3a
      12'h53F: dout  = 8'b01111000; // 1343 : 120 - 0x78
      12'h540: dout  = 8'b00100000; // 1344 :  32 - 0x20 -- Sprite 0xa8
      12'h541: dout  = 8'b01010001; // 1345 :  81 - 0x51
      12'h542: dout  = 8'b00001010; // 1346 :  10 - 0xa
      12'h543: dout  = 8'b00000100; // 1347 :   4 - 0x4
      12'h544: dout  = 8'b11101010; // 1348 : 234 - 0xea
      12'h545: dout  = 8'b00111001; // 1349 :  57 - 0x39
      12'h546: dout  = 8'b01111111; // 1350 : 127 - 0x7f
      12'h547: dout  = 8'b11110000; // 1351 : 240 - 0xf0
      12'h548: dout  = 8'b10111100; // 1352 : 188 - 0xbc -- Sprite 0xa9
      12'h549: dout  = 8'b01011000; // 1353 :  88 - 0x58
      12'h54A: dout  = 8'b00111000; // 1354 :  56 - 0x38
      12'h54B: dout  = 8'b00010000; // 1355 :  16 - 0x10
      12'h54C: dout  = 8'b00110000; // 1356 :  48 - 0x30
      12'h54D: dout  = 8'b11111000; // 1357 : 248 - 0xf8
      12'h54E: dout  = 8'b11111100; // 1358 : 252 - 0xfc
      12'h54F: dout  = 8'b00111110; // 1359 :  62 - 0x3e
      12'h550: dout  = 8'b00000000; // 1360 :   0 - 0x0 -- Sprite 0xaa
      12'h551: dout  = 8'b00000000; // 1361 :   0 - 0x0
      12'h552: dout  = 8'b00000000; // 1362 :   0 - 0x0
      12'h553: dout  = 8'b00000110; // 1363 :   6 - 0x6
      12'h554: dout  = 8'b00001110; // 1364 :  14 - 0xe
      12'h555: dout  = 8'b00001100; // 1365 :  12 - 0xc
      12'h556: dout  = 8'b00000000; // 1366 :   0 - 0x0
      12'h557: dout  = 8'b00000000; // 1367 :   0 - 0x0
      12'h558: dout  = 8'b00000000; // 1368 :   0 - 0x0 -- Sprite 0xab
      12'h559: dout  = 8'b00000000; // 1369 :   0 - 0x0
      12'h55A: dout  = 8'b00000000; // 1370 :   0 - 0x0
      12'h55B: dout  = 8'b00000000; // 1371 :   0 - 0x0
      12'h55C: dout  = 8'b00000000; // 1372 :   0 - 0x0
      12'h55D: dout  = 8'b00000000; // 1373 :   0 - 0x0
      12'h55E: dout  = 8'b00001111; // 1374 :  15 - 0xf
      12'h55F: dout  = 8'b00011000; // 1375 :  24 - 0x18
      12'h560: dout  = 8'b00000000; // 1376 :   0 - 0x0 -- Sprite 0xac
      12'h561: dout  = 8'b00000000; // 1377 :   0 - 0x0
      12'h562: dout  = 8'b00000000; // 1378 :   0 - 0x0
      12'h563: dout  = 8'b00000000; // 1379 :   0 - 0x0
      12'h564: dout  = 8'b11111000; // 1380 : 248 - 0xf8
      12'h565: dout  = 8'b00111110; // 1381 :  62 - 0x3e
      12'h566: dout  = 8'b00111011; // 1382 :  59 - 0x3b
      12'h567: dout  = 8'b00011000; // 1383 :  24 - 0x18
      12'h568: dout  = 8'b00010000; // 1384 :  16 - 0x10 -- Sprite 0xad
      12'h569: dout  = 8'b00010100; // 1385 :  20 - 0x14
      12'h56A: dout  = 8'b00010000; // 1386 :  16 - 0x10
      12'h56B: dout  = 8'b00010000; // 1387 :  16 - 0x10
      12'h56C: dout  = 8'b00111000; // 1388 :  56 - 0x38
      12'h56D: dout  = 8'b01111000; // 1389 : 120 - 0x78
      12'h56E: dout  = 8'b11111000; // 1390 : 248 - 0xf8
      12'h56F: dout  = 8'b00110000; // 1391 :  48 - 0x30
      12'h570: dout  = 8'b00000000; // 1392 :   0 - 0x0 -- Sprite 0xae
      12'h571: dout  = 8'b00000000; // 1393 :   0 - 0x0
      12'h572: dout  = 8'b00000000; // 1394 :   0 - 0x0
      12'h573: dout  = 8'b00000000; // 1395 :   0 - 0x0
      12'h574: dout  = 8'b00000110; // 1396 :   6 - 0x6
      12'h575: dout  = 8'b00001110; // 1397 :  14 - 0xe
      12'h576: dout  = 8'b00001100; // 1398 :  12 - 0xc
      12'h577: dout  = 8'b00000000; // 1399 :   0 - 0x0
      12'h578: dout  = 8'b00000000; // 1400 :   0 - 0x0 -- Sprite 0xaf
      12'h579: dout  = 8'b00000000; // 1401 :   0 - 0x0
      12'h57A: dout  = 8'b00000000; // 1402 :   0 - 0x0
      12'h57B: dout  = 8'b00000000; // 1403 :   0 - 0x0
      12'h57C: dout  = 8'b00000000; // 1404 :   0 - 0x0
      12'h57D: dout  = 8'b00000000; // 1405 :   0 - 0x0
      12'h57E: dout  = 8'b00000000; // 1406 :   0 - 0x0
      12'h57F: dout  = 8'b00001111; // 1407 :  15 - 0xf
      12'h580: dout  = 8'b00000000; // 1408 :   0 - 0x0 -- Sprite 0xb0
      12'h581: dout  = 8'b00000000; // 1409 :   0 - 0x0
      12'h582: dout  = 8'b00000000; // 1410 :   0 - 0x0
      12'h583: dout  = 8'b00000000; // 1411 :   0 - 0x0
      12'h584: dout  = 8'b00000000; // 1412 :   0 - 0x0
      12'h585: dout  = 8'b11111000; // 1413 : 248 - 0xf8
      12'h586: dout  = 8'b01111110; // 1414 : 126 - 0x7e
      12'h587: dout  = 8'b11110011; // 1415 : 243 - 0xf3
      12'h588: dout  = 8'b00011000; // 1416 :  24 - 0x18 -- Sprite 0xb1
      12'h589: dout  = 8'b00010000; // 1417 :  16 - 0x10
      12'h58A: dout  = 8'b00010100; // 1418 :  20 - 0x14
      12'h58B: dout  = 8'b00010000; // 1419 :  16 - 0x10
      12'h58C: dout  = 8'b00010000; // 1420 :  16 - 0x10
      12'h58D: dout  = 8'b00111000; // 1421 :  56 - 0x38
      12'h58E: dout  = 8'b01111100; // 1422 : 124 - 0x7c
      12'h58F: dout  = 8'b11011110; // 1423 : 222 - 0xde
      12'h590: dout  = 8'b00000000; // 1424 :   0 - 0x0 -- Sprite 0xb2
      12'h591: dout  = 8'b00001101; // 1425 :  13 - 0xd
      12'h592: dout  = 8'b00011110; // 1426 :  30 - 0x1e
      12'h593: dout  = 8'b00011110; // 1427 :  30 - 0x1e
      12'h594: dout  = 8'b00011110; // 1428 :  30 - 0x1e
      12'h595: dout  = 8'b00011111; // 1429 :  31 - 0x1f
      12'h596: dout  = 8'b00001111; // 1430 :  15 - 0xf
      12'h597: dout  = 8'b00000111; // 1431 :   7 - 0x7
      12'h598: dout  = 8'b01111000; // 1432 : 120 - 0x78 -- Sprite 0xb3
      12'h599: dout  = 8'b11110000; // 1433 : 240 - 0xf0
      12'h59A: dout  = 8'b00000000; // 1434 :   0 - 0x0
      12'h59B: dout  = 8'b00011010; // 1435 :  26 - 0x1a
      12'h59C: dout  = 8'b00111111; // 1436 :  63 - 0x3f
      12'h59D: dout  = 8'b00110101; // 1437 :  53 - 0x35
      12'h59E: dout  = 8'b00110101; // 1438 :  53 - 0x35
      12'h59F: dout  = 8'b00111111; // 1439 :  63 - 0x3f
      12'h5A0: dout  = 8'b00000000; // 1440 :   0 - 0x0 -- Sprite 0xb4
      12'h5A1: dout  = 8'b00000000; // 1441 :   0 - 0x0
      12'h5A2: dout  = 8'b10000000; // 1442 : 128 - 0x80
      12'h5A3: dout  = 8'b11100000; // 1443 : 224 - 0xe0
      12'h5A4: dout  = 8'b11100000; // 1444 : 224 - 0xe0
      12'h5A5: dout  = 8'b01110000; // 1445 : 112 - 0x70
      12'h5A6: dout  = 8'b01110011; // 1446 : 115 - 0x73
      12'h5A7: dout  = 8'b00100001; // 1447 :  33 - 0x21
      12'h5A8: dout  = 8'b00011010; // 1448 :  26 - 0x1a -- Sprite 0xb5
      12'h5A9: dout  = 8'b00000111; // 1449 :   7 - 0x7
      12'h5AA: dout  = 8'b00001100; // 1450 :  12 - 0xc
      12'h5AB: dout  = 8'b00011000; // 1451 :  24 - 0x18
      12'h5AC: dout  = 8'b01111000; // 1452 : 120 - 0x78
      12'h5AD: dout  = 8'b11111110; // 1453 : 254 - 0xfe
      12'h5AE: dout  = 8'b11111100; // 1454 : 252 - 0xfc
      12'h5AF: dout  = 8'b11110000; // 1455 : 240 - 0xf0
      12'h5B0: dout  = 8'b00000000; // 1456 :   0 - 0x0 -- Sprite 0xb6
      12'h5B1: dout  = 8'b00000001; // 1457 :   1 - 0x1
      12'h5B2: dout  = 8'b00000010; // 1458 :   2 - 0x2
      12'h5B3: dout  = 8'b00000000; // 1459 :   0 - 0x0
      12'h5B4: dout  = 8'b00111000; // 1460 :  56 - 0x38
      12'h5B5: dout  = 8'b01111100; // 1461 : 124 - 0x7c
      12'h5B6: dout  = 8'b01111110; // 1462 : 126 - 0x7e
      12'h5B7: dout  = 8'b00111111; // 1463 :  63 - 0x3f
      12'h5B8: dout  = 8'b00111111; // 1464 :  63 - 0x3f -- Sprite 0xb7
      12'h5B9: dout  = 8'b01000000; // 1465 :  64 - 0x40
      12'h5BA: dout  = 8'b01100000; // 1466 :  96 - 0x60
      12'h5BB: dout  = 8'b01100000; // 1467 :  96 - 0x60
      12'h5BC: dout  = 8'b00100000; // 1468 :  32 - 0x20
      12'h5BD: dout  = 8'b00110000; // 1469 :  48 - 0x30
      12'h5BE: dout  = 8'b00010011; // 1470 :  19 - 0x13
      12'h5BF: dout  = 8'b00000001; // 1471 :   1 - 0x1
      12'h5C0: dout  = 8'b11000000; // 1472 : 192 - 0xc0 -- Sprite 0xb8
      12'h5C1: dout  = 8'b11100000; // 1473 : 224 - 0xe0
      12'h5C2: dout  = 8'b00110000; // 1474 :  48 - 0x30
      12'h5C3: dout  = 8'b11010000; // 1475 : 208 - 0xd0
      12'h5C4: dout  = 8'b11010000; // 1476 : 208 - 0xd0
      12'h5C5: dout  = 8'b11010000; // 1477 : 208 - 0xd0
      12'h5C6: dout  = 8'b11010000; // 1478 : 208 - 0xd0
      12'h5C7: dout  = 8'b00000000; // 1479 :   0 - 0x0
      12'h5C8: dout  = 8'b00000111; // 1480 :   7 - 0x7 -- Sprite 0xb9
      12'h5C9: dout  = 8'b00001111; // 1481 :  15 - 0xf
      12'h5CA: dout  = 8'b00000010; // 1482 :   2 - 0x2
      12'h5CB: dout  = 8'b00011101; // 1483 :  29 - 0x1d
      12'h5CC: dout  = 8'b00011111; // 1484 :  31 - 0x1f
      12'h5CD: dout  = 8'b00011010; // 1485 :  26 - 0x1a
      12'h5CE: dout  = 8'b00011010; // 1486 :  26 - 0x1a
      12'h5CF: dout  = 8'b00000010; // 1487 :   2 - 0x2
      12'h5D0: dout  = 8'b00111000; // 1488 :  56 - 0x38 -- Sprite 0xba
      12'h5D1: dout  = 8'b01111100; // 1489 : 124 - 0x7c
      12'h5D2: dout  = 8'b11111100; // 1490 : 252 - 0xfc
      12'h5D3: dout  = 8'b11111100; // 1491 : 252 - 0xfc
      12'h5D4: dout  = 8'b11111100; // 1492 : 252 - 0xfc
      12'h5D5: dout  = 8'b11111110; // 1493 : 254 - 0xfe
      12'h5D6: dout  = 8'b10111110; // 1494 : 190 - 0xbe
      12'h5D7: dout  = 8'b10111110; // 1495 : 190 - 0xbe
      12'h5D8: dout  = 8'b00011100; // 1496 :  28 - 0x1c -- Sprite 0xbb
      12'h5D9: dout  = 8'b00111110; // 1497 :  62 - 0x3e
      12'h5DA: dout  = 8'b00111111; // 1498 :  63 - 0x3f
      12'h5DB: dout  = 8'b00111111; // 1499 :  63 - 0x3f
      12'h5DC: dout  = 8'b00111111; // 1500 :  63 - 0x3f
      12'h5DD: dout  = 8'b01111111; // 1501 : 127 - 0x7f
      12'h5DE: dout  = 8'b01111101; // 1502 : 125 - 0x7d
      12'h5DF: dout  = 8'b01111101; // 1503 : 125 - 0x7d
      12'h5E0: dout  = 8'b01111101; // 1504 : 125 - 0x7d -- Sprite 0xbc
      12'h5E1: dout  = 8'b01111111; // 1505 : 127 - 0x7f
      12'h5E2: dout  = 8'b01011111; // 1506 :  95 - 0x5f
      12'h5E3: dout  = 8'b00111011; // 1507 :  59 - 0x3b
      12'h5E4: dout  = 8'b00111100; // 1508 :  60 - 0x3c
      12'h5E5: dout  = 8'b00111111; // 1509 :  63 - 0x3f
      12'h5E6: dout  = 8'b00011110; // 1510 :  30 - 0x1e
      12'h5E7: dout  = 8'b00000000; // 1511 :   0 - 0x0
      12'h5E8: dout  = 8'b00011100; // 1512 :  28 - 0x1c -- Sprite 0xbd
      12'h5E9: dout  = 8'b00111110; // 1513 :  62 - 0x3e
      12'h5EA: dout  = 8'b00111111; // 1514 :  63 - 0x3f
      12'h5EB: dout  = 8'b00011111; // 1515 :  31 - 0x1f
      12'h5EC: dout  = 8'b00111111; // 1516 :  63 - 0x3f
      12'h5ED: dout  = 8'b01111111; // 1517 : 127 - 0x7f
      12'h5EE: dout  = 8'b01111101; // 1518 : 125 - 0x7d
      12'h5EF: dout  = 8'b01111101; // 1519 : 125 - 0x7d
      12'h5F0: dout  = 8'b00000000; // 1520 :   0 - 0x0 -- Sprite 0xbe
      12'h5F1: dout  = 8'b00000000; // 1521 :   0 - 0x0
      12'h5F2: dout  = 8'b00000000; // 1522 :   0 - 0x0
      12'h5F3: dout  = 8'b01100000; // 1523 :  96 - 0x60
      12'h5F4: dout  = 8'b01100010; // 1524 :  98 - 0x62
      12'h5F5: dout  = 8'b01100101; // 1525 : 101 - 0x65
      12'h5F6: dout  = 8'b00111111; // 1526 :  63 - 0x3f
      12'h5F7: dout  = 8'b00011111; // 1527 :  31 - 0x1f
      12'h5F8: dout  = 8'b01110000; // 1528 : 112 - 0x70 -- Sprite 0xbf
      12'h5F9: dout  = 8'b00111100; // 1529 :  60 - 0x3c
      12'h5FA: dout  = 8'b00111100; // 1530 :  60 - 0x3c
      12'h5FB: dout  = 8'b00011000; // 1531 :  24 - 0x18
      12'h5FC: dout  = 8'b00000000; // 1532 :   0 - 0x0
      12'h5FD: dout  = 8'b00000000; // 1533 :   0 - 0x0
      12'h5FE: dout  = 8'b00000010; // 1534 :   2 - 0x2
      12'h5FF: dout  = 8'b00000111; // 1535 :   7 - 0x7
      12'h600: dout  = 8'b11001111; // 1536 : 207 - 0xcf -- Sprite 0xc0
      12'h601: dout  = 8'b01111010; // 1537 : 122 - 0x7a
      12'h602: dout  = 8'b01011010; // 1538 :  90 - 0x5a
      12'h603: dout  = 8'b00010000; // 1539 :  16 - 0x10
      12'h604: dout  = 8'b00000000; // 1540 :   0 - 0x0
      12'h605: dout  = 8'b00000000; // 1541 :   0 - 0x0
      12'h606: dout  = 8'b11000000; // 1542 : 192 - 0xc0
      12'h607: dout  = 8'b10000000; // 1543 : 128 - 0x80
      12'h608: dout  = 8'b10000101; // 1544 : 133 - 0x85 -- Sprite 0xc1
      12'h609: dout  = 8'b10000100; // 1545 : 132 - 0x84
      12'h60A: dout  = 8'b10000110; // 1546 : 134 - 0x86
      12'h60B: dout  = 8'b11000110; // 1547 : 198 - 0xc6
      12'h60C: dout  = 8'b11100111; // 1548 : 231 - 0xe7
      12'h60D: dout  = 8'b01110011; // 1549 : 115 - 0x73
      12'h60E: dout  = 8'b01110011; // 1550 : 115 - 0x73
      12'h60F: dout  = 8'b11100001; // 1551 : 225 - 0xe1
      12'h610: dout  = 8'b10000000; // 1552 : 128 - 0x80 -- Sprite 0xc2
      12'h611: dout  = 8'b01001110; // 1553 :  78 - 0x4e
      12'h612: dout  = 8'b01110111; // 1554 : 119 - 0x77
      12'h613: dout  = 8'b11110011; // 1555 : 243 - 0xf3
      12'h614: dout  = 8'b11111011; // 1556 : 251 - 0xfb
      12'h615: dout  = 8'b11111001; // 1557 : 249 - 0xf9
      12'h616: dout  = 8'b11111010; // 1558 : 250 - 0xfa
      12'h617: dout  = 8'b01111000; // 1559 : 120 - 0x78
      12'h618: dout  = 8'b00010001; // 1560 :  17 - 0x11 -- Sprite 0xc3
      12'h619: dout  = 8'b00111001; // 1561 :  57 - 0x39
      12'h61A: dout  = 8'b01111101; // 1562 : 125 - 0x7d
      12'h61B: dout  = 8'b00111001; // 1563 :  57 - 0x39
      12'h61C: dout  = 8'b00000000; // 1564 :   0 - 0x0
      12'h61D: dout  = 8'b00000000; // 1565 :   0 - 0x0
      12'h61E: dout  = 8'b11100000; // 1566 : 224 - 0xe0
      12'h61F: dout  = 8'b11100111; // 1567 : 231 - 0xe7
      12'h620: dout  = 8'b00000000; // 1568 :   0 - 0x0 -- Sprite 0xc4
      12'h621: dout  = 8'b00000000; // 1569 :   0 - 0x0
      12'h622: dout  = 8'b00000111; // 1570 :   7 - 0x7
      12'h623: dout  = 8'b00000111; // 1571 :   7 - 0x7
      12'h624: dout  = 8'b00010110; // 1572 :  22 - 0x16
      12'h625: dout  = 8'b00010000; // 1573 :  16 - 0x10
      12'h626: dout  = 8'b00000000; // 1574 :   0 - 0x0
      12'h627: dout  = 8'b00111000; // 1575 :  56 - 0x38
      12'h628: dout  = 8'b11001111; // 1576 : 207 - 0xcf -- Sprite 0xc5
      12'h629: dout  = 8'b00011111; // 1577 :  31 - 0x1f
      12'h62A: dout  = 8'b00010111; // 1578 :  23 - 0x17
      12'h62B: dout  = 8'b00010000; // 1579 :  16 - 0x10
      12'h62C: dout  = 8'b00110011; // 1580 :  51 - 0x33
      12'h62D: dout  = 8'b00110000; // 1581 :  48 - 0x30
      12'h62E: dout  = 8'b00110000; // 1582 :  48 - 0x30
      12'h62F: dout  = 8'b00100000; // 1583 :  32 - 0x20
      12'h630: dout  = 8'b00111000; // 1584 :  56 - 0x38 -- Sprite 0xc6
      12'h631: dout  = 8'b00110000; // 1585 :  48 - 0x30
      12'h632: dout  = 8'b01000000; // 1586 :  64 - 0x40
      12'h633: dout  = 8'b11000111; // 1587 : 199 - 0xc7
      12'h634: dout  = 8'b00000111; // 1588 :   7 - 0x7
      12'h635: dout  = 8'b01100110; // 1589 : 102 - 0x66
      12'h636: dout  = 8'b11100000; // 1590 : 224 - 0xe0
      12'h637: dout  = 8'b01101100; // 1591 : 108 - 0x6c
      12'h638: dout  = 8'b01100000; // 1592 :  96 - 0x60 -- Sprite 0xc7
      12'h639: dout  = 8'b11000000; // 1593 : 192 - 0xc0
      12'h63A: dout  = 8'b10000000; // 1594 : 128 - 0x80
      12'h63B: dout  = 8'b00000100; // 1595 :   4 - 0x4
      12'h63C: dout  = 8'b10011110; // 1596 : 158 - 0x9e
      12'h63D: dout  = 8'b11111111; // 1597 : 255 - 0xff
      12'h63E: dout  = 8'b11110000; // 1598 : 240 - 0xf0
      12'h63F: dout  = 8'b11111000; // 1599 : 248 - 0xf8
      12'h640: dout  = 8'b00100100; // 1600 :  36 - 0x24 -- Sprite 0xc8
      12'h641: dout  = 8'b00000001; // 1601 :   1 - 0x1
      12'h642: dout  = 8'b00000111; // 1602 :   7 - 0x7
      12'h643: dout  = 8'b11111110; // 1603 : 254 - 0xfe
      12'h644: dout  = 8'b11111111; // 1604 : 255 - 0xff
      12'h645: dout  = 8'b01111111; // 1605 : 127 - 0x7f
      12'h646: dout  = 8'b00111111; // 1606 :  63 - 0x3f
      12'h647: dout  = 8'b01111111; // 1607 : 127 - 0x7f
      12'h648: dout  = 8'b11001111; // 1608 : 207 - 0xcf -- Sprite 0xc9
      12'h649: dout  = 8'b01111010; // 1609 : 122 - 0x7a
      12'h64A: dout  = 8'b00001010; // 1610 :  10 - 0xa
      12'h64B: dout  = 8'b11111110; // 1611 : 254 - 0xfe
      12'h64C: dout  = 8'b11111100; // 1612 : 252 - 0xfc
      12'h64D: dout  = 8'b00000000; // 1613 :   0 - 0x0
      12'h64E: dout  = 8'b00000000; // 1614 :   0 - 0x0
      12'h64F: dout  = 8'b00000000; // 1615 :   0 - 0x0
      12'h650: dout  = 8'b10000101; // 1616 : 133 - 0x85 -- Sprite 0xca
      12'h651: dout  = 8'b10000110; // 1617 : 134 - 0x86
      12'h652: dout  = 8'b10000011; // 1618 : 131 - 0x83
      12'h653: dout  = 8'b11000011; // 1619 : 195 - 0xc3
      12'h654: dout  = 8'b11100001; // 1620 : 225 - 0xe1
      12'h655: dout  = 8'b01110000; // 1621 : 112 - 0x70
      12'h656: dout  = 8'b01110000; // 1622 : 112 - 0x70
      12'h657: dout  = 8'b11100000; // 1623 : 224 - 0xe0
      12'h658: dout  = 8'b01100000; // 1624 :  96 - 0x60 -- Sprite 0xcb
      12'h659: dout  = 8'b11000000; // 1625 : 192 - 0xc0
      12'h65A: dout  = 8'b10000000; // 1626 : 128 - 0x80
      12'h65B: dout  = 8'b00000000; // 1627 :   0 - 0x0
      12'h65C: dout  = 8'b10011000; // 1628 : 152 - 0x98
      12'h65D: dout  = 8'b11111100; // 1629 : 252 - 0xfc
      12'h65E: dout  = 8'b11111110; // 1630 : 254 - 0xfe
      12'h65F: dout  = 8'b11111111; // 1631 : 255 - 0xff
      12'h660: dout  = 8'b00100100; // 1632 :  36 - 0x24 -- Sprite 0xcc
      12'h661: dout  = 8'b00000000; // 1633 :   0 - 0x0
      12'h662: dout  = 8'b00000111; // 1634 :   7 - 0x7
      12'h663: dout  = 8'b11111110; // 1635 : 254 - 0xfe
      12'h664: dout  = 8'b11111111; // 1636 : 255 - 0xff
      12'h665: dout  = 8'b01111111; // 1637 : 127 - 0x7f
      12'h666: dout  = 8'b11111111; // 1638 : 255 - 0xff
      12'h667: dout  = 8'b00000011; // 1639 :   3 - 0x3
      12'h668: dout  = 8'b00000011; // 1640 :   3 - 0x3 -- Sprite 0xcd
      12'h669: dout  = 8'b00001111; // 1641 :  15 - 0xf
      12'h66A: dout  = 8'b00100011; // 1642 :  35 - 0x23
      12'h66B: dout  = 8'b01100010; // 1643 :  98 - 0x62
      12'h66C: dout  = 8'b01100100; // 1644 : 100 - 0x64
      12'h66D: dout  = 8'b00111100; // 1645 :  60 - 0x3c
      12'h66E: dout  = 8'b00011100; // 1646 :  28 - 0x1c
      12'h66F: dout  = 8'b00011110; // 1647 :  30 - 0x1e
      12'h670: dout  = 8'b00011111; // 1648 :  31 - 0x1f -- Sprite 0xce
      12'h671: dout  = 8'b00111101; // 1649 :  61 - 0x3d
      12'h672: dout  = 8'b01101101; // 1650 : 109 - 0x6d
      12'h673: dout  = 8'b01001111; // 1651 :  79 - 0x4f
      12'h674: dout  = 8'b11101110; // 1652 : 238 - 0xee
      12'h675: dout  = 8'b11110011; // 1653 : 243 - 0xf3
      12'h676: dout  = 8'b00100000; // 1654 :  32 - 0x20
      12'h677: dout  = 8'b00000011; // 1655 :   3 - 0x3
      12'h678: dout  = 8'b00000111; // 1656 :   7 - 0x7 -- Sprite 0xcf
      12'h679: dout  = 8'b00000111; // 1657 :   7 - 0x7
      12'h67A: dout  = 8'b00011111; // 1658 :  31 - 0x1f
      12'h67B: dout  = 8'b00111111; // 1659 :  63 - 0x3f
      12'h67C: dout  = 8'b00001111; // 1660 :  15 - 0xf
      12'h67D: dout  = 8'b01000111; // 1661 :  71 - 0x47
      12'h67E: dout  = 8'b00000011; // 1662 :   3 - 0x3
      12'h67F: dout  = 8'b00000000; // 1663 :   0 - 0x0
      12'h680: dout  = 8'b00000000; // 1664 :   0 - 0x0 -- Sprite 0xd0
      12'h681: dout  = 8'b00000000; // 1665 :   0 - 0x0
      12'h682: dout  = 8'b00000011; // 1666 :   3 - 0x3
      12'h683: dout  = 8'b00000111; // 1667 :   7 - 0x7
      12'h684: dout  = 8'b00001111; // 1668 :  15 - 0xf
      12'h685: dout  = 8'b00001111; // 1669 :  15 - 0xf
      12'h686: dout  = 8'b00011111; // 1670 :  31 - 0x1f
      12'h687: dout  = 8'b00011111; // 1671 :  31 - 0x1f
      12'h688: dout  = 8'b00000000; // 1672 :   0 - 0x0 -- Sprite 0xd1
      12'h689: dout  = 8'b00100011; // 1673 :  35 - 0x23
      12'h68A: dout  = 8'b01010111; // 1674 :  87 - 0x57
      12'h68B: dout  = 8'b01001111; // 1675 :  79 - 0x4f
      12'h68C: dout  = 8'b01010111; // 1676 :  87 - 0x57
      12'h68D: dout  = 8'b00101111; // 1677 :  47 - 0x2f
      12'h68E: dout  = 8'b11011111; // 1678 : 223 - 0xdf
      12'h68F: dout  = 8'b00100001; // 1679 :  33 - 0x21
      12'h690: dout  = 8'b00000000; // 1680 :   0 - 0x0 -- Sprite 0xd2
      12'h691: dout  = 8'b00000000; // 1681 :   0 - 0x0
      12'h692: dout  = 8'b00000000; // 1682 :   0 - 0x0
      12'h693: dout  = 8'b00000000; // 1683 :   0 - 0x0
      12'h694: dout  = 8'b10000000; // 1684 : 128 - 0x80
      12'h695: dout  = 8'b10000000; // 1685 : 128 - 0x80
      12'h696: dout  = 8'b00000000; // 1686 :   0 - 0x0
      12'h697: dout  = 8'b00000000; // 1687 :   0 - 0x0
      12'h698: dout  = 8'b00100011; // 1688 :  35 - 0x23 -- Sprite 0xd3
      12'h699: dout  = 8'b00001111; // 1689 :  15 - 0xf
      12'h69A: dout  = 8'b00011110; // 1690 :  30 - 0x1e
      12'h69B: dout  = 8'b11110000; // 1691 : 240 - 0xf0
      12'h69C: dout  = 8'b00011100; // 1692 :  28 - 0x1c
      12'h69D: dout  = 8'b00111111; // 1693 :  63 - 0x3f
      12'h69E: dout  = 8'b00011111; // 1694 :  31 - 0x1f
      12'h69F: dout  = 8'b00011110; // 1695 :  30 - 0x1e
      12'h6A0: dout  = 8'b00000000; // 1696 :   0 - 0x0 -- Sprite 0xd4
      12'h6A1: dout  = 8'b10000000; // 1697 : 128 - 0x80
      12'h6A2: dout  = 8'b00011000; // 1698 :  24 - 0x18
      12'h6A3: dout  = 8'b00110000; // 1699 :  48 - 0x30
      12'h6A4: dout  = 8'b00110100; // 1700 :  52 - 0x34
      12'h6A5: dout  = 8'b11111110; // 1701 : 254 - 0xfe
      12'h6A6: dout  = 8'b11111110; // 1702 : 254 - 0xfe
      12'h6A7: dout  = 8'b11111110; // 1703 : 254 - 0xfe
      12'h6A8: dout  = 8'b00000000; // 1704 :   0 - 0x0 -- Sprite 0xd5
      12'h6A9: dout  = 8'b00000000; // 1705 :   0 - 0x0
      12'h6AA: dout  = 8'b00000001; // 1706 :   1 - 0x1
      12'h6AB: dout  = 8'b00000100; // 1707 :   4 - 0x4
      12'h6AC: dout  = 8'b00000110; // 1708 :   6 - 0x6
      12'h6AD: dout  = 8'b00000110; // 1709 :   6 - 0x6
      12'h6AE: dout  = 8'b00000111; // 1710 :   7 - 0x7
      12'h6AF: dout  = 8'b00000111; // 1711 :   7 - 0x7
      12'h6B0: dout  = 8'b00001111; // 1712 :  15 - 0xf -- Sprite 0xd6
      12'h6B1: dout  = 8'b00111111; // 1713 :  63 - 0x3f
      12'h6B2: dout  = 8'b01111111; // 1714 : 127 - 0x7f
      12'h6B3: dout  = 8'b11111000; // 1715 : 248 - 0xf8
      12'h6B4: dout  = 8'b11111000; // 1716 : 248 - 0xf8
      12'h6B5: dout  = 8'b01111111; // 1717 : 127 - 0x7f
      12'h6B6: dout  = 8'b00111111; // 1718 :  63 - 0x3f
      12'h6B7: dout  = 8'b00001111; // 1719 :  15 - 0xf
      12'h6B8: dout  = 8'b00011111; // 1720 :  31 - 0x1f -- Sprite 0xd7
      12'h6B9: dout  = 8'b00011111; // 1721 :  31 - 0x1f
      12'h6BA: dout  = 8'b00011111; // 1722 :  31 - 0x1f
      12'h6BB: dout  = 8'b00001011; // 1723 :  11 - 0xb
      12'h6BC: dout  = 8'b00000001; // 1724 :   1 - 0x1
      12'h6BD: dout  = 8'b00000001; // 1725 :   1 - 0x1
      12'h6BE: dout  = 8'b00000000; // 1726 :   0 - 0x0
      12'h6BF: dout  = 8'b00000000; // 1727 :   0 - 0x0
      12'h6C0: dout  = 8'b00000011; // 1728 :   3 - 0x3 -- Sprite 0xd8
      12'h6C1: dout  = 8'b00011111; // 1729 :  31 - 0x1f
      12'h6C2: dout  = 8'b00111111; // 1730 :  63 - 0x3f
      12'h6C3: dout  = 8'b00111111; // 1731 :  63 - 0x3f
      12'h6C4: dout  = 8'b01111000; // 1732 : 120 - 0x78
      12'h6C5: dout  = 8'b00000000; // 1733 :   0 - 0x0
      12'h6C6: dout  = 8'b00000011; // 1734 :   3 - 0x3
      12'h6C7: dout  = 8'b11111111; // 1735 : 255 - 0xff
      12'h6C8: dout  = 8'b00000000; // 1736 :   0 - 0x0 -- Sprite 0xd9
      12'h6C9: dout  = 8'b00000000; // 1737 :   0 - 0x0
      12'h6CA: dout  = 8'b00000000; // 1738 :   0 - 0x0
      12'h6CB: dout  = 8'b00000000; // 1739 :   0 - 0x0
      12'h6CC: dout  = 8'b00000000; // 1740 :   0 - 0x0
      12'h6CD: dout  = 8'b00000000; // 1741 :   0 - 0x0
      12'h6CE: dout  = 8'b00000000; // 1742 :   0 - 0x0
      12'h6CF: dout  = 8'b00000000; // 1743 :   0 - 0x0
      12'h6D0: dout  = 8'b00100011; // 1744 :  35 - 0x23 -- Sprite 0xda
      12'h6D1: dout  = 8'b00100111; // 1745 :  39 - 0x27
      12'h6D2: dout  = 8'b00011111; // 1746 :  31 - 0x1f
      12'h6D3: dout  = 8'b00000111; // 1747 :   7 - 0x7
      12'h6D4: dout  = 8'b00001111; // 1748 :  15 - 0xf
      12'h6D5: dout  = 8'b00011111; // 1749 :  31 - 0x1f
      12'h6D6: dout  = 8'b01111111; // 1750 : 127 - 0x7f
      12'h6D7: dout  = 8'b00111111; // 1751 :  63 - 0x3f
      12'h6D8: dout  = 8'b11100000; // 1752 : 224 - 0xe0 -- Sprite 0xdb
      12'h6D9: dout  = 8'b10000000; // 1753 : 128 - 0x80
      12'h6DA: dout  = 8'b10000000; // 1754 : 128 - 0x80
      12'h6DB: dout  = 8'b01000000; // 1755 :  64 - 0x40
      12'h6DC: dout  = 8'b11100000; // 1756 : 224 - 0xe0
      12'h6DD: dout  = 8'b11100000; // 1757 : 224 - 0xe0
      12'h6DE: dout  = 8'b11100000; // 1758 : 224 - 0xe0
      12'h6DF: dout  = 8'b11000000; // 1759 : 192 - 0xc0
      12'h6E0: dout  = 8'b00000011; // 1760 :   3 - 0x3 -- Sprite 0xdc
      12'h6E1: dout  = 8'b00000111; // 1761 :   7 - 0x7
      12'h6E2: dout  = 8'b00001111; // 1762 :  15 - 0xf
      12'h6E3: dout  = 8'b00011111; // 1763 :  31 - 0x1f
      12'h6E4: dout  = 8'b00111111; // 1764 :  63 - 0x3f
      12'h6E5: dout  = 8'b01111111; // 1765 : 127 - 0x7f
      12'h6E6: dout  = 8'b11111111; // 1766 : 255 - 0xff
      12'h6E7: dout  = 8'b00011111; // 1767 :  31 - 0x1f
      12'h6E8: dout  = 8'b00011111; // 1768 :  31 - 0x1f -- Sprite 0xdd
      12'h6E9: dout  = 8'b00010000; // 1769 :  16 - 0x10
      12'h6EA: dout  = 8'b00001100; // 1770 :  12 - 0xc
      12'h6EB: dout  = 8'b00010010; // 1771 :  18 - 0x12
      12'h6EC: dout  = 8'b00010010; // 1772 :  18 - 0x12
      12'h6ED: dout  = 8'b00101100; // 1773 :  44 - 0x2c
      12'h6EE: dout  = 8'b00111111; // 1774 :  63 - 0x3f
      12'h6EF: dout  = 8'b00111111; // 1775 :  63 - 0x3f
      12'h6F0: dout  = 8'b00110111; // 1776 :  55 - 0x37 -- Sprite 0xde
      12'h6F1: dout  = 8'b00110110; // 1777 :  54 - 0x36
      12'h6F2: dout  = 8'b00110110; // 1778 :  54 - 0x36
      12'h6F3: dout  = 8'b00110110; // 1779 :  54 - 0x36
      12'h6F4: dout  = 8'b00010110; // 1780 :  22 - 0x16
      12'h6F5: dout  = 8'b00010110; // 1781 :  22 - 0x16
      12'h6F6: dout  = 8'b00010010; // 1782 :  18 - 0x12
      12'h6F7: dout  = 8'b00000010; // 1783 :   2 - 0x2
      12'h6F8: dout  = 8'b00010000; // 1784 :  16 - 0x10 -- Sprite 0xdf
      12'h6F9: dout  = 8'b01111110; // 1785 : 126 - 0x7e
      12'h6FA: dout  = 8'b11111111; // 1786 : 255 - 0xff
      12'h6FB: dout  = 8'b11111111; // 1787 : 255 - 0xff
      12'h6FC: dout  = 8'b11110110; // 1788 : 246 - 0xf6
      12'h6FD: dout  = 8'b01110110; // 1789 : 118 - 0x76
      12'h6FE: dout  = 8'b00111010; // 1790 :  58 - 0x3a
      12'h6FF: dout  = 8'b00011010; // 1791 :  26 - 0x1a
      12'h700: dout  = 8'b00000000; // 1792 :   0 - 0x0 -- Sprite 0xe0
      12'h701: dout  = 8'b00000000; // 1793 :   0 - 0x0
      12'h702: dout  = 8'b00111000; // 1794 :  56 - 0x38
      12'h703: dout  = 8'b00000100; // 1795 :   4 - 0x4
      12'h704: dout  = 8'b00000000; // 1796 :   0 - 0x0
      12'h705: dout  = 8'b00000000; // 1797 :   0 - 0x0
      12'h706: dout  = 8'b00000000; // 1798 :   0 - 0x0
      12'h707: dout  = 8'b00000000; // 1799 :   0 - 0x0
      12'h708: dout  = 8'b00000000; // 1800 :   0 - 0x0 -- Sprite 0xe1
      12'h709: dout  = 8'b00000000; // 1801 :   0 - 0x0
      12'h70A: dout  = 8'b00000000; // 1802 :   0 - 0x0
      12'h70B: dout  = 8'b00111000; // 1803 :  56 - 0x38
      12'h70C: dout  = 8'b01000000; // 1804 :  64 - 0x40
      12'h70D: dout  = 8'b00000000; // 1805 :   0 - 0x0
      12'h70E: dout  = 8'b00000000; // 1806 :   0 - 0x0
      12'h70F: dout  = 8'b00000000; // 1807 :   0 - 0x0
      12'h710: dout  = 8'b11111100; // 1808 : 252 - 0xfc -- Sprite 0xe2
      12'h711: dout  = 8'b10100000; // 1809 : 160 - 0xa0
      12'h712: dout  = 8'b10000000; // 1810 : 128 - 0x80
      12'h713: dout  = 8'b10000000; // 1811 : 128 - 0x80
      12'h714: dout  = 8'b00000000; // 1812 :   0 - 0x0
      12'h715: dout  = 8'b00000000; // 1813 :   0 - 0x0
      12'h716: dout  = 8'b00000000; // 1814 :   0 - 0x0
      12'h717: dout  = 8'b00000000; // 1815 :   0 - 0x0
      12'h718: dout  = 8'b00000111; // 1816 :   7 - 0x7 -- Sprite 0xe3
      12'h719: dout  = 8'b00100111; // 1817 :  39 - 0x27
      12'h71A: dout  = 8'b01010111; // 1818 :  87 - 0x57
      12'h71B: dout  = 8'b01001111; // 1819 :  79 - 0x4f
      12'h71C: dout  = 8'b01010111; // 1820 :  87 - 0x57
      12'h71D: dout  = 8'b00100111; // 1821 :  39 - 0x27
      12'h71E: dout  = 8'b11000001; // 1822 : 193 - 0xc1
      12'h71F: dout  = 8'b00100001; // 1823 :  33 - 0x21
      12'h720: dout  = 8'b00011101; // 1824 :  29 - 0x1d -- Sprite 0xe4
      12'h721: dout  = 8'b00001111; // 1825 :  15 - 0xf
      12'h722: dout  = 8'b00001111; // 1826 :  15 - 0xf
      12'h723: dout  = 8'b00011111; // 1827 :  31 - 0x1f
      12'h724: dout  = 8'b00011111; // 1828 :  31 - 0x1f
      12'h725: dout  = 8'b00011110; // 1829 :  30 - 0x1e
      12'h726: dout  = 8'b00111000; // 1830 :  56 - 0x38
      12'h727: dout  = 8'b00110000; // 1831 :  48 - 0x30
      12'h728: dout  = 8'b00000000; // 1832 :   0 - 0x0 -- Sprite 0xe5
      12'h729: dout  = 8'b00000000; // 1833 :   0 - 0x0
      12'h72A: dout  = 8'b00111000; // 1834 :  56 - 0x38
      12'h72B: dout  = 8'b00010000; // 1835 :  16 - 0x10
      12'h72C: dout  = 8'b01001100; // 1836 :  76 - 0x4c
      12'h72D: dout  = 8'b00011000; // 1837 :  24 - 0x18
      12'h72E: dout  = 8'b10000110; // 1838 : 134 - 0x86
      12'h72F: dout  = 8'b00100100; // 1839 :  36 - 0x24
      12'h730: dout  = 8'b00000000; // 1840 :   0 - 0x0 -- Sprite 0xe6
      12'h731: dout  = 8'b01000010; // 1841 :  66 - 0x42
      12'h732: dout  = 8'b00001010; // 1842 :  10 - 0xa
      12'h733: dout  = 8'b01000000; // 1843 :  64 - 0x40
      12'h734: dout  = 8'b00010000; // 1844 :  16 - 0x10
      12'h735: dout  = 8'b00000010; // 1845 :   2 - 0x2
      12'h736: dout  = 8'b00001000; // 1846 :   8 - 0x8
      12'h737: dout  = 8'b00000010; // 1847 :   2 - 0x2
      12'h738: dout  = 8'b00000000; // 1848 :   0 - 0x0 -- Sprite 0xe7
      12'h739: dout  = 8'b00000000; // 1849 :   0 - 0x0
      12'h73A: dout  = 8'b10000000; // 1850 : 128 - 0x80
      12'h73B: dout  = 8'b01000000; // 1851 :  64 - 0x40
      12'h73C: dout  = 8'b00001000; // 1852 :   8 - 0x8
      12'h73D: dout  = 8'b00001100; // 1853 :  12 - 0xc
      12'h73E: dout  = 8'b00001010; // 1854 :  10 - 0xa
      12'h73F: dout  = 8'b10000100; // 1855 : 132 - 0x84
      12'h740: dout  = 8'b00000000; // 1856 :   0 - 0x0 -- Sprite 0xe8
      12'h741: dout  = 8'b00000000; // 1857 :   0 - 0x0
      12'h742: dout  = 8'b11001111; // 1858 : 207 - 0xcf
      12'h743: dout  = 8'b00100000; // 1859 :  32 - 0x20
      12'h744: dout  = 8'b00100000; // 1860 :  32 - 0x20
      12'h745: dout  = 8'b00100000; // 1861 :  32 - 0x20
      12'h746: dout  = 8'b00100110; // 1862 :  38 - 0x26
      12'h747: dout  = 8'b00101110; // 1863 :  46 - 0x2e
      12'h748: dout  = 8'b11100000; // 1864 : 224 - 0xe0 -- Sprite 0xe9
      12'h749: dout  = 8'b11100000; // 1865 : 224 - 0xe0
      12'h74A: dout  = 8'b11000000; // 1866 : 192 - 0xc0
      12'h74B: dout  = 8'b00000000; // 1867 :   0 - 0x0
      12'h74C: dout  = 8'b00000000; // 1868 :   0 - 0x0
      12'h74D: dout  = 8'b00000000; // 1869 :   0 - 0x0
      12'h74E: dout  = 8'b00000000; // 1870 :   0 - 0x0
      12'h74F: dout  = 8'b00000000; // 1871 :   0 - 0x0
      12'h750: dout  = 8'b00101111; // 1872 :  47 - 0x2f -- Sprite 0xea
      12'h751: dout  = 8'b00100011; // 1873 :  35 - 0x23
      12'h752: dout  = 8'b00100001; // 1874 :  33 - 0x21
      12'h753: dout  = 8'b00100000; // 1875 :  32 - 0x20
      12'h754: dout  = 8'b00100000; // 1876 :  32 - 0x20
      12'h755: dout  = 8'b00000000; // 1877 :   0 - 0x0
      12'h756: dout  = 8'b00000000; // 1878 :   0 - 0x0
      12'h757: dout  = 8'b00000000; // 1879 :   0 - 0x0
      12'h758: dout  = 8'b11000001; // 1880 : 193 - 0xc1 -- Sprite 0xeb
      12'h759: dout  = 8'b10110001; // 1881 : 177 - 0xb1
      12'h75A: dout  = 8'b01011001; // 1882 :  89 - 0x59
      12'h75B: dout  = 8'b01101101; // 1883 : 109 - 0x6d
      12'h75C: dout  = 8'b00110101; // 1884 :  53 - 0x35
      12'h75D: dout  = 8'b00111011; // 1885 :  59 - 0x3b
      12'h75E: dout  = 8'b00011111; // 1886 :  31 - 0x1f
      12'h75F: dout  = 8'b00000011; // 1887 :   3 - 0x3
      12'h760: dout  = 8'b00000000; // 1888 :   0 - 0x0 -- Sprite 0xec
      12'h761: dout  = 8'b00000010; // 1889 :   2 - 0x2
      12'h762: dout  = 8'b00000000; // 1890 :   0 - 0x0
      12'h763: dout  = 8'b00001000; // 1891 :   8 - 0x8
      12'h764: dout  = 8'b00000010; // 1892 :   2 - 0x2
      12'h765: dout  = 8'b00000000; // 1893 :   0 - 0x0
      12'h766: dout  = 8'b00101000; // 1894 :  40 - 0x28
      12'h767: dout  = 8'b00000000; // 1895 :   0 - 0x0
      12'h768: dout  = 8'b00000100; // 1896 :   4 - 0x4 -- Sprite 0xed
      12'h769: dout  = 8'b00010000; // 1897 :  16 - 0x10
      12'h76A: dout  = 8'b00000010; // 1898 :   2 - 0x2
      12'h76B: dout  = 8'b00010000; // 1899 :  16 - 0x10
      12'h76C: dout  = 8'b00000100; // 1900 :   4 - 0x4
      12'h76D: dout  = 8'b00000000; // 1901 :   0 - 0x0
      12'h76E: dout  = 8'b00001010; // 1902 :  10 - 0xa
      12'h76F: dout  = 8'b00000000; // 1903 :   0 - 0x0
      12'h770: dout  = 8'b11000001; // 1904 : 193 - 0xc1 -- Sprite 0xee
      12'h771: dout  = 8'b10110001; // 1905 : 177 - 0xb1
      12'h772: dout  = 8'b01011001; // 1906 :  89 - 0x59
      12'h773: dout  = 8'b01101101; // 1907 : 109 - 0x6d
      12'h774: dout  = 8'b00110101; // 1908 :  53 - 0x35
      12'h775: dout  = 8'b00111011; // 1909 :  59 - 0x3b
      12'h776: dout  = 8'b00011111; // 1910 :  31 - 0x1f
      12'h777: dout  = 8'b00000011; // 1911 :   3 - 0x3
      12'h778: dout  = 8'b00000000; // 1912 :   0 - 0x0 -- Sprite 0xef
      12'h779: dout  = 8'b00001111; // 1913 :  15 - 0xf
      12'h77A: dout  = 8'b00011111; // 1914 :  31 - 0x1f
      12'h77B: dout  = 8'b11111111; // 1915 : 255 - 0xff
      12'h77C: dout  = 8'b11111100; // 1916 : 252 - 0xfc
      12'h77D: dout  = 8'b01100011; // 1917 :  99 - 0x63
      12'h77E: dout  = 8'b00011111; // 1918 :  31 - 0x1f
      12'h77F: dout  = 8'b00000011; // 1919 :   3 - 0x3
      12'h780: dout  = 8'b00000000; // 1920 :   0 - 0x0 -- Sprite 0xf0
      12'h781: dout  = 8'b00000000; // 1921 :   0 - 0x0
      12'h782: dout  = 8'b11111110; // 1922 : 254 - 0xfe
      12'h783: dout  = 8'b11000110; // 1923 : 198 - 0xc6
      12'h784: dout  = 8'b11000110; // 1924 : 198 - 0xc6
      12'h785: dout  = 8'b11111110; // 1925 : 254 - 0xfe
      12'h786: dout  = 8'b00000000; // 1926 :   0 - 0x0
      12'h787: dout  = 8'b00000000; // 1927 :   0 - 0x0
      12'h788: dout  = 8'b00000000; // 1928 :   0 - 0x0 -- Sprite 0xf1
      12'h789: dout  = 8'b00000000; // 1929 :   0 - 0x0
      12'h78A: dout  = 8'b00000110; // 1930 :   6 - 0x6
      12'h78B: dout  = 8'b00000110; // 1931 :   6 - 0x6
      12'h78C: dout  = 8'b00001100; // 1932 :  12 - 0xc
      12'h78D: dout  = 8'b00011000; // 1933 :  24 - 0x18
      12'h78E: dout  = 8'b01110000; // 1934 : 112 - 0x70
      12'h78F: dout  = 8'b01100000; // 1935 :  96 - 0x60
      12'h790: dout  = 8'b00000000; // 1936 :   0 - 0x0 -- Sprite 0xf2
      12'h791: dout  = 8'b00000000; // 1937 :   0 - 0x0
      12'h792: dout  = 8'b00000110; // 1938 :   6 - 0x6
      12'h793: dout  = 8'b00000110; // 1939 :   6 - 0x6
      12'h794: dout  = 8'b00000100; // 1940 :   4 - 0x4
      12'h795: dout  = 8'b00000100; // 1941 :   4 - 0x4
      12'h796: dout  = 8'b00001000; // 1942 :   8 - 0x8
      12'h797: dout  = 8'b00001000; // 1943 :   8 - 0x8
      12'h798: dout  = 8'b00001000; // 1944 :   8 - 0x8 -- Sprite 0xf3
      12'h799: dout  = 8'b00010000; // 1945 :  16 - 0x10
      12'h79A: dout  = 8'b00110000; // 1946 :  48 - 0x30
      12'h79B: dout  = 8'b00110000; // 1947 :  48 - 0x30
      12'h79C: dout  = 8'b00110000; // 1948 :  48 - 0x30
      12'h79D: dout  = 8'b00110000; // 1949 :  48 - 0x30
      12'h79E: dout  = 8'b00010000; // 1950 :  16 - 0x10
      12'h79F: dout  = 8'b00001000; // 1951 :   8 - 0x8
      12'h7A0: dout  = 8'b00000000; // 1952 :   0 - 0x0 -- Sprite 0xf4
      12'h7A1: dout  = 8'b00000000; // 1953 :   0 - 0x0
      12'h7A2: dout  = 8'b00000001; // 1954 :   1 - 0x1
      12'h7A3: dout  = 8'b00000011; // 1955 :   3 - 0x3
      12'h7A4: dout  = 8'b00000001; // 1956 :   1 - 0x1
      12'h7A5: dout  = 8'b00000000; // 1957 :   0 - 0x0
      12'h7A6: dout  = 8'b00000000; // 1958 :   0 - 0x0
      12'h7A7: dout  = 8'b00000000; // 1959 :   0 - 0x0
      12'h7A8: dout  = 8'b00000011; // 1960 :   3 - 0x3 -- Sprite 0xf5
      12'h7A9: dout  = 8'b00001110; // 1961 :  14 - 0xe
      12'h7AA: dout  = 8'b11111000; // 1962 : 248 - 0xf8
      12'h7AB: dout  = 8'b00000000; // 1963 :   0 - 0x0
      12'h7AC: dout  = 8'b00000000; // 1964 :   0 - 0x0
      12'h7AD: dout  = 8'b00000000; // 1965 :   0 - 0x0
      12'h7AE: dout  = 8'b00000000; // 1966 :   0 - 0x0
      12'h7AF: dout  = 8'b00000000; // 1967 :   0 - 0x0
      12'h7B0: dout  = 8'b00100010; // 1968 :  34 - 0x22 -- Sprite 0xf6
      12'h7B1: dout  = 8'b01100101; // 1969 : 101 - 0x65
      12'h7B2: dout  = 8'b00100101; // 1970 :  37 - 0x25
      12'h7B3: dout  = 8'b00100101; // 1971 :  37 - 0x25
      12'h7B4: dout  = 8'b00100101; // 1972 :  37 - 0x25
      12'h7B5: dout  = 8'b00100101; // 1973 :  37 - 0x25
      12'h7B6: dout  = 8'b01110111; // 1974 : 119 - 0x77
      12'h7B7: dout  = 8'b01110010; // 1975 : 114 - 0x72
      12'h7B8: dout  = 8'b01100010; // 1976 :  98 - 0x62 -- Sprite 0xf7
      12'h7B9: dout  = 8'b10010101; // 1977 : 149 - 0x95
      12'h7BA: dout  = 8'b00010101; // 1978 :  21 - 0x15
      12'h7BB: dout  = 8'b00100101; // 1979 :  37 - 0x25
      12'h7BC: dout  = 8'b01000101; // 1980 :  69 - 0x45
      12'h7BD: dout  = 8'b10000101; // 1981 : 133 - 0x85
      12'h7BE: dout  = 8'b11110111; // 1982 : 247 - 0xf7
      12'h7BF: dout  = 8'b11110010; // 1983 : 242 - 0xf2
      12'h7C0: dout  = 8'b10100010; // 1984 : 162 - 0xa2 -- Sprite 0xf8
      12'h7C1: dout  = 8'b10100101; // 1985 : 165 - 0xa5
      12'h7C2: dout  = 8'b10100101; // 1986 : 165 - 0xa5
      12'h7C3: dout  = 8'b10100101; // 1987 : 165 - 0xa5
      12'h7C4: dout  = 8'b11110101; // 1988 : 245 - 0xf5
      12'h7C5: dout  = 8'b11110101; // 1989 : 245 - 0xf5
      12'h7C6: dout  = 8'b00100111; // 1990 :  39 - 0x27
      12'h7C7: dout  = 8'b00100010; // 1991 :  34 - 0x22
      12'h7C8: dout  = 8'b11110010; // 1992 : 242 - 0xf2 -- Sprite 0xf9
      12'h7C9: dout  = 8'b10000101; // 1993 : 133 - 0x85
      12'h7CA: dout  = 8'b10000101; // 1994 : 133 - 0x85
      12'h7CB: dout  = 8'b11100101; // 1995 : 229 - 0xe5
      12'h7CC: dout  = 8'b00010101; // 1996 :  21 - 0x15
      12'h7CD: dout  = 8'b00010101; // 1997 :  21 - 0x15
      12'h7CE: dout  = 8'b11110111; // 1998 : 247 - 0xf7
      12'h7CF: dout  = 8'b11100010; // 1999 : 226 - 0xe2
      12'h7D0: dout  = 8'b01100010; // 2000 :  98 - 0x62 -- Sprite 0xfa
      12'h7D1: dout  = 8'b10010101; // 2001 : 149 - 0x95
      12'h7D2: dout  = 8'b01010101; // 2002 :  85 - 0x55
      12'h7D3: dout  = 8'b01100101; // 2003 : 101 - 0x65
      12'h7D4: dout  = 8'b10110101; // 2004 : 181 - 0xb5
      12'h7D5: dout  = 8'b10010101; // 2005 : 149 - 0x95
      12'h7D6: dout  = 8'b10010111; // 2006 : 151 - 0x97
      12'h7D7: dout  = 8'b01100010; // 2007 :  98 - 0x62
      12'h7D8: dout  = 8'b00100000; // 2008 :  32 - 0x20 -- Sprite 0xfb
      12'h7D9: dout  = 8'b01010000; // 2009 :  80 - 0x50
      12'h7DA: dout  = 8'b01010000; // 2010 :  80 - 0x50
      12'h7DB: dout  = 8'b01010000; // 2011 :  80 - 0x50
      12'h7DC: dout  = 8'b01010000; // 2012 :  80 - 0x50
      12'h7DD: dout  = 8'b01010000; // 2013 :  80 - 0x50
      12'h7DE: dout  = 8'b01110000; // 2014 : 112 - 0x70
      12'h7DF: dout  = 8'b00100000; // 2015 :  32 - 0x20
      12'h7E0: dout  = 8'b00000000; // 2016 :   0 - 0x0 -- Sprite 0xfc
      12'h7E1: dout  = 8'b00000000; // 2017 :   0 - 0x0
      12'h7E2: dout  = 8'b00000000; // 2018 :   0 - 0x0
      12'h7E3: dout  = 8'b00000000; // 2019 :   0 - 0x0
      12'h7E4: dout  = 8'b00000000; // 2020 :   0 - 0x0
      12'h7E5: dout  = 8'b00000000; // 2021 :   0 - 0x0
      12'h7E6: dout  = 8'b00000000; // 2022 :   0 - 0x0
      12'h7E7: dout  = 8'b00000000; // 2023 :   0 - 0x0
      12'h7E8: dout  = 8'b01100110; // 2024 : 102 - 0x66 -- Sprite 0xfd
      12'h7E9: dout  = 8'b11100110; // 2025 : 230 - 0xe6
      12'h7EA: dout  = 8'b01100110; // 2026 : 102 - 0x66
      12'h7EB: dout  = 8'b01100110; // 2027 : 102 - 0x66
      12'h7EC: dout  = 8'b01100110; // 2028 : 102 - 0x66
      12'h7ED: dout  = 8'b01100111; // 2029 : 103 - 0x67
      12'h7EE: dout  = 8'b11110011; // 2030 : 243 - 0xf3
      12'h7EF: dout  = 8'b00000000; // 2031 :   0 - 0x0
      12'h7F0: dout  = 8'b01011110; // 2032 :  94 - 0x5e -- Sprite 0xfe
      12'h7F1: dout  = 8'b01011001; // 2033 :  89 - 0x59
      12'h7F2: dout  = 8'b01011001; // 2034 :  89 - 0x59
      12'h7F3: dout  = 8'b01011001; // 2035 :  89 - 0x59
      12'h7F4: dout  = 8'b01011110; // 2036 :  94 - 0x5e
      12'h7F5: dout  = 8'b11011000; // 2037 : 216 - 0xd8
      12'h7F6: dout  = 8'b10011000; // 2038 : 152 - 0x98
      12'h7F7: dout  = 8'b00000000; // 2039 :   0 - 0x0
      12'h7F8: dout  = 8'b00000000; // 2040 :   0 - 0x0 -- Sprite 0xff
      12'h7F9: dout  = 8'b00000000; // 2041 :   0 - 0x0
      12'h7FA: dout  = 8'b00000000; // 2042 :   0 - 0x0
      12'h7FB: dout  = 8'b00000000; // 2043 :   0 - 0x0
      12'h7FC: dout  = 8'b00000000; // 2044 :   0 - 0x0
      12'h7FD: dout  = 8'b00000100; // 2045 :   4 - 0x4
      12'h7FE: dout  = 8'b00001000; // 2046 :   8 - 0x8
      12'h7FF: dout  = 8'b00000000; // 2047 :   0 - 0x0
          // Background pattern Table
      12'h800: dout  = 8'b00000000; // 2048 :   0 - 0x0 -- Background 0x0
      12'h801: dout  = 8'b00000000; // 2049 :   0 - 0x0
      12'h802: dout  = 8'b00000000; // 2050 :   0 - 0x0
      12'h803: dout  = 8'b00000000; // 2051 :   0 - 0x0
      12'h804: dout  = 8'b00000000; // 2052 :   0 - 0x0
      12'h805: dout  = 8'b00000000; // 2053 :   0 - 0x0
      12'h806: dout  = 8'b00000000; // 2054 :   0 - 0x0
      12'h807: dout  = 8'b00000000; // 2055 :   0 - 0x0
      12'h808: dout  = 8'b00000000; // 2056 :   0 - 0x0 -- Background 0x1
      12'h809: dout  = 8'b00000000; // 2057 :   0 - 0x0
      12'h80A: dout  = 8'b00000000; // 2058 :   0 - 0x0
      12'h80B: dout  = 8'b00000000; // 2059 :   0 - 0x0
      12'h80C: dout  = 8'b00000000; // 2060 :   0 - 0x0
      12'h80D: dout  = 8'b00000000; // 2061 :   0 - 0x0
      12'h80E: dout  = 8'b00000000; // 2062 :   0 - 0x0
      12'h80F: dout  = 8'b00000000; // 2063 :   0 - 0x0
      12'h810: dout  = 8'b00000000; // 2064 :   0 - 0x0 -- Background 0x2
      12'h811: dout  = 8'b00000000; // 2065 :   0 - 0x0
      12'h812: dout  = 8'b00000000; // 2066 :   0 - 0x0
      12'h813: dout  = 8'b00000000; // 2067 :   0 - 0x0
      12'h814: dout  = 8'b00000000; // 2068 :   0 - 0x0
      12'h815: dout  = 8'b00000000; // 2069 :   0 - 0x0
      12'h816: dout  = 8'b00000000; // 2070 :   0 - 0x0
      12'h817: dout  = 8'b00000000; // 2071 :   0 - 0x0
      12'h818: dout  = 8'b00000000; // 2072 :   0 - 0x0 -- Background 0x3
      12'h819: dout  = 8'b00000000; // 2073 :   0 - 0x0
      12'h81A: dout  = 8'b00000000; // 2074 :   0 - 0x0
      12'h81B: dout  = 8'b00000000; // 2075 :   0 - 0x0
      12'h81C: dout  = 8'b00000000; // 2076 :   0 - 0x0
      12'h81D: dout  = 8'b00000000; // 2077 :   0 - 0x0
      12'h81E: dout  = 8'b00000000; // 2078 :   0 - 0x0
      12'h81F: dout  = 8'b00000000; // 2079 :   0 - 0x0
      12'h820: dout  = 8'b00000000; // 2080 :   0 - 0x0 -- Background 0x4
      12'h821: dout  = 8'b00000000; // 2081 :   0 - 0x0
      12'h822: dout  = 8'b00000000; // 2082 :   0 - 0x0
      12'h823: dout  = 8'b00000000; // 2083 :   0 - 0x0
      12'h824: dout  = 8'b00000000; // 2084 :   0 - 0x0
      12'h825: dout  = 8'b00000000; // 2085 :   0 - 0x0
      12'h826: dout  = 8'b00000000; // 2086 :   0 - 0x0
      12'h827: dout  = 8'b00000000; // 2087 :   0 - 0x0
      12'h828: dout  = 8'b00000000; // 2088 :   0 - 0x0 -- Background 0x5
      12'h829: dout  = 8'b00000000; // 2089 :   0 - 0x0
      12'h82A: dout  = 8'b00000000; // 2090 :   0 - 0x0
      12'h82B: dout  = 8'b00000000; // 2091 :   0 - 0x0
      12'h82C: dout  = 8'b00000000; // 2092 :   0 - 0x0
      12'h82D: dout  = 8'b00000000; // 2093 :   0 - 0x0
      12'h82E: dout  = 8'b00000000; // 2094 :   0 - 0x0
      12'h82F: dout  = 8'b00000000; // 2095 :   0 - 0x0
      12'h830: dout  = 8'b00000000; // 2096 :   0 - 0x0 -- Background 0x6
      12'h831: dout  = 8'b00000000; // 2097 :   0 - 0x0
      12'h832: dout  = 8'b00000000; // 2098 :   0 - 0x0
      12'h833: dout  = 8'b00000000; // 2099 :   0 - 0x0
      12'h834: dout  = 8'b00000000; // 2100 :   0 - 0x0
      12'h835: dout  = 8'b00000000; // 2101 :   0 - 0x0
      12'h836: dout  = 8'b00000000; // 2102 :   0 - 0x0
      12'h837: dout  = 8'b00000000; // 2103 :   0 - 0x0
      12'h838: dout  = 8'b00000000; // 2104 :   0 - 0x0 -- Background 0x7
      12'h839: dout  = 8'b00000000; // 2105 :   0 - 0x0
      12'h83A: dout  = 8'b00000000; // 2106 :   0 - 0x0
      12'h83B: dout  = 8'b00000000; // 2107 :   0 - 0x0
      12'h83C: dout  = 8'b00000000; // 2108 :   0 - 0x0
      12'h83D: dout  = 8'b00000000; // 2109 :   0 - 0x0
      12'h83E: dout  = 8'b00000000; // 2110 :   0 - 0x0
      12'h83F: dout  = 8'b00000000; // 2111 :   0 - 0x0
      12'h840: dout  = 8'b00000000; // 2112 :   0 - 0x0 -- Background 0x8
      12'h841: dout  = 8'b00000000; // 2113 :   0 - 0x0
      12'h842: dout  = 8'b00000000; // 2114 :   0 - 0x0
      12'h843: dout  = 8'b00000000; // 2115 :   0 - 0x0
      12'h844: dout  = 8'b00000000; // 2116 :   0 - 0x0
      12'h845: dout  = 8'b00000000; // 2117 :   0 - 0x0
      12'h846: dout  = 8'b00000000; // 2118 :   0 - 0x0
      12'h847: dout  = 8'b00000000; // 2119 :   0 - 0x0
      12'h848: dout  = 8'b00000000; // 2120 :   0 - 0x0 -- Background 0x9
      12'h849: dout  = 8'b00000000; // 2121 :   0 - 0x0
      12'h84A: dout  = 8'b00000000; // 2122 :   0 - 0x0
      12'h84B: dout  = 8'b00000000; // 2123 :   0 - 0x0
      12'h84C: dout  = 8'b00000000; // 2124 :   0 - 0x0
      12'h84D: dout  = 8'b00000000; // 2125 :   0 - 0x0
      12'h84E: dout  = 8'b00000000; // 2126 :   0 - 0x0
      12'h84F: dout  = 8'b00000000; // 2127 :   0 - 0x0
      12'h850: dout  = 8'b00000000; // 2128 :   0 - 0x0 -- Background 0xa
      12'h851: dout  = 8'b00000000; // 2129 :   0 - 0x0
      12'h852: dout  = 8'b00000000; // 2130 :   0 - 0x0
      12'h853: dout  = 8'b00000000; // 2131 :   0 - 0x0
      12'h854: dout  = 8'b00000000; // 2132 :   0 - 0x0
      12'h855: dout  = 8'b00000000; // 2133 :   0 - 0x0
      12'h856: dout  = 8'b00000000; // 2134 :   0 - 0x0
      12'h857: dout  = 8'b00000000; // 2135 :   0 - 0x0
      12'h858: dout  = 8'b00000000; // 2136 :   0 - 0x0 -- Background 0xb
      12'h859: dout  = 8'b00000000; // 2137 :   0 - 0x0
      12'h85A: dout  = 8'b00000000; // 2138 :   0 - 0x0
      12'h85B: dout  = 8'b00000000; // 2139 :   0 - 0x0
      12'h85C: dout  = 8'b00000000; // 2140 :   0 - 0x0
      12'h85D: dout  = 8'b00000000; // 2141 :   0 - 0x0
      12'h85E: dout  = 8'b00000000; // 2142 :   0 - 0x0
      12'h85F: dout  = 8'b00000000; // 2143 :   0 - 0x0
      12'h860: dout  = 8'b00000000; // 2144 :   0 - 0x0 -- Background 0xc
      12'h861: dout  = 8'b00000000; // 2145 :   0 - 0x0
      12'h862: dout  = 8'b00000000; // 2146 :   0 - 0x0
      12'h863: dout  = 8'b00000000; // 2147 :   0 - 0x0
      12'h864: dout  = 8'b00000000; // 2148 :   0 - 0x0
      12'h865: dout  = 8'b00000000; // 2149 :   0 - 0x0
      12'h866: dout  = 8'b00000000; // 2150 :   0 - 0x0
      12'h867: dout  = 8'b00000000; // 2151 :   0 - 0x0
      12'h868: dout  = 8'b00000000; // 2152 :   0 - 0x0 -- Background 0xd
      12'h869: dout  = 8'b00000000; // 2153 :   0 - 0x0
      12'h86A: dout  = 8'b00000000; // 2154 :   0 - 0x0
      12'h86B: dout  = 8'b00000000; // 2155 :   0 - 0x0
      12'h86C: dout  = 8'b00000000; // 2156 :   0 - 0x0
      12'h86D: dout  = 8'b00000000; // 2157 :   0 - 0x0
      12'h86E: dout  = 8'b00000000; // 2158 :   0 - 0x0
      12'h86F: dout  = 8'b00000000; // 2159 :   0 - 0x0
      12'h870: dout  = 8'b00000000; // 2160 :   0 - 0x0 -- Background 0xe
      12'h871: dout  = 8'b00000000; // 2161 :   0 - 0x0
      12'h872: dout  = 8'b00000000; // 2162 :   0 - 0x0
      12'h873: dout  = 8'b00000000; // 2163 :   0 - 0x0
      12'h874: dout  = 8'b00000000; // 2164 :   0 - 0x0
      12'h875: dout  = 8'b00000000; // 2165 :   0 - 0x0
      12'h876: dout  = 8'b00000000; // 2166 :   0 - 0x0
      12'h877: dout  = 8'b00000000; // 2167 :   0 - 0x0
      12'h878: dout  = 8'b00000000; // 2168 :   0 - 0x0 -- Background 0xf
      12'h879: dout  = 8'b00000000; // 2169 :   0 - 0x0
      12'h87A: dout  = 8'b00000000; // 2170 :   0 - 0x0
      12'h87B: dout  = 8'b00000000; // 2171 :   0 - 0x0
      12'h87C: dout  = 8'b00000000; // 2172 :   0 - 0x0
      12'h87D: dout  = 8'b00000000; // 2173 :   0 - 0x0
      12'h87E: dout  = 8'b00000000; // 2174 :   0 - 0x0
      12'h87F: dout  = 8'b00000000; // 2175 :   0 - 0x0
      12'h880: dout  = 8'b00000000; // 2176 :   0 - 0x0 -- Background 0x10
      12'h881: dout  = 8'b00000000; // 2177 :   0 - 0x0
      12'h882: dout  = 8'b00000000; // 2178 :   0 - 0x0
      12'h883: dout  = 8'b00000000; // 2179 :   0 - 0x0
      12'h884: dout  = 8'b00000000; // 2180 :   0 - 0x0
      12'h885: dout  = 8'b00000000; // 2181 :   0 - 0x0
      12'h886: dout  = 8'b00000000; // 2182 :   0 - 0x0
      12'h887: dout  = 8'b00000000; // 2183 :   0 - 0x0
      12'h888: dout  = 8'b00000000; // 2184 :   0 - 0x0 -- Background 0x11
      12'h889: dout  = 8'b00000000; // 2185 :   0 - 0x0
      12'h88A: dout  = 8'b00000000; // 2186 :   0 - 0x0
      12'h88B: dout  = 8'b00000000; // 2187 :   0 - 0x0
      12'h88C: dout  = 8'b00000000; // 2188 :   0 - 0x0
      12'h88D: dout  = 8'b00000000; // 2189 :   0 - 0x0
      12'h88E: dout  = 8'b00000000; // 2190 :   0 - 0x0
      12'h88F: dout  = 8'b00000000; // 2191 :   0 - 0x0
      12'h890: dout  = 8'b00000000; // 2192 :   0 - 0x0 -- Background 0x12
      12'h891: dout  = 8'b00000000; // 2193 :   0 - 0x0
      12'h892: dout  = 8'b00000000; // 2194 :   0 - 0x0
      12'h893: dout  = 8'b00000000; // 2195 :   0 - 0x0
      12'h894: dout  = 8'b00000000; // 2196 :   0 - 0x0
      12'h895: dout  = 8'b00000000; // 2197 :   0 - 0x0
      12'h896: dout  = 8'b00000000; // 2198 :   0 - 0x0
      12'h897: dout  = 8'b00000000; // 2199 :   0 - 0x0
      12'h898: dout  = 8'b00000000; // 2200 :   0 - 0x0 -- Background 0x13
      12'h899: dout  = 8'b00000000; // 2201 :   0 - 0x0
      12'h89A: dout  = 8'b00000000; // 2202 :   0 - 0x0
      12'h89B: dout  = 8'b00000000; // 2203 :   0 - 0x0
      12'h89C: dout  = 8'b00000000; // 2204 :   0 - 0x0
      12'h89D: dout  = 8'b00000000; // 2205 :   0 - 0x0
      12'h89E: dout  = 8'b00000000; // 2206 :   0 - 0x0
      12'h89F: dout  = 8'b00000000; // 2207 :   0 - 0x0
      12'h8A0: dout  = 8'b00000000; // 2208 :   0 - 0x0 -- Background 0x14
      12'h8A1: dout  = 8'b00000000; // 2209 :   0 - 0x0
      12'h8A2: dout  = 8'b00000000; // 2210 :   0 - 0x0
      12'h8A3: dout  = 8'b00000000; // 2211 :   0 - 0x0
      12'h8A4: dout  = 8'b00000000; // 2212 :   0 - 0x0
      12'h8A5: dout  = 8'b00000000; // 2213 :   0 - 0x0
      12'h8A6: dout  = 8'b00000000; // 2214 :   0 - 0x0
      12'h8A7: dout  = 8'b00000000; // 2215 :   0 - 0x0
      12'h8A8: dout  = 8'b00000000; // 2216 :   0 - 0x0 -- Background 0x15
      12'h8A9: dout  = 8'b00000000; // 2217 :   0 - 0x0
      12'h8AA: dout  = 8'b00000000; // 2218 :   0 - 0x0
      12'h8AB: dout  = 8'b00000000; // 2219 :   0 - 0x0
      12'h8AC: dout  = 8'b00000000; // 2220 :   0 - 0x0
      12'h8AD: dout  = 8'b00000000; // 2221 :   0 - 0x0
      12'h8AE: dout  = 8'b00000000; // 2222 :   0 - 0x0
      12'h8AF: dout  = 8'b00000000; // 2223 :   0 - 0x0
      12'h8B0: dout  = 8'b00000000; // 2224 :   0 - 0x0 -- Background 0x16
      12'h8B1: dout  = 8'b00000000; // 2225 :   0 - 0x0
      12'h8B2: dout  = 8'b00000000; // 2226 :   0 - 0x0
      12'h8B3: dout  = 8'b00000000; // 2227 :   0 - 0x0
      12'h8B4: dout  = 8'b00000000; // 2228 :   0 - 0x0
      12'h8B5: dout  = 8'b00000000; // 2229 :   0 - 0x0
      12'h8B6: dout  = 8'b00000000; // 2230 :   0 - 0x0
      12'h8B7: dout  = 8'b00000000; // 2231 :   0 - 0x0
      12'h8B8: dout  = 8'b00000000; // 2232 :   0 - 0x0 -- Background 0x17
      12'h8B9: dout  = 8'b00000000; // 2233 :   0 - 0x0
      12'h8BA: dout  = 8'b00000000; // 2234 :   0 - 0x0
      12'h8BB: dout  = 8'b00000000; // 2235 :   0 - 0x0
      12'h8BC: dout  = 8'b00000000; // 2236 :   0 - 0x0
      12'h8BD: dout  = 8'b00000000; // 2237 :   0 - 0x0
      12'h8BE: dout  = 8'b00000000; // 2238 :   0 - 0x0
      12'h8BF: dout  = 8'b00000000; // 2239 :   0 - 0x0
      12'h8C0: dout  = 8'b00000000; // 2240 :   0 - 0x0 -- Background 0x18
      12'h8C1: dout  = 8'b00000000; // 2241 :   0 - 0x0
      12'h8C2: dout  = 8'b00000000; // 2242 :   0 - 0x0
      12'h8C3: dout  = 8'b00000000; // 2243 :   0 - 0x0
      12'h8C4: dout  = 8'b00000000; // 2244 :   0 - 0x0
      12'h8C5: dout  = 8'b00000000; // 2245 :   0 - 0x0
      12'h8C6: dout  = 8'b00000000; // 2246 :   0 - 0x0
      12'h8C7: dout  = 8'b00000000; // 2247 :   0 - 0x0
      12'h8C8: dout  = 8'b00000000; // 2248 :   0 - 0x0 -- Background 0x19
      12'h8C9: dout  = 8'b00000000; // 2249 :   0 - 0x0
      12'h8CA: dout  = 8'b00000000; // 2250 :   0 - 0x0
      12'h8CB: dout  = 8'b00000000; // 2251 :   0 - 0x0
      12'h8CC: dout  = 8'b00000000; // 2252 :   0 - 0x0
      12'h8CD: dout  = 8'b00000000; // 2253 :   0 - 0x0
      12'h8CE: dout  = 8'b00000000; // 2254 :   0 - 0x0
      12'h8CF: dout  = 8'b00000000; // 2255 :   0 - 0x0
      12'h8D0: dout  = 8'b00000000; // 2256 :   0 - 0x0 -- Background 0x1a
      12'h8D1: dout  = 8'b00000000; // 2257 :   0 - 0x0
      12'h8D2: dout  = 8'b00000000; // 2258 :   0 - 0x0
      12'h8D3: dout  = 8'b00000000; // 2259 :   0 - 0x0
      12'h8D4: dout  = 8'b00000000; // 2260 :   0 - 0x0
      12'h8D5: dout  = 8'b00000000; // 2261 :   0 - 0x0
      12'h8D6: dout  = 8'b00000000; // 2262 :   0 - 0x0
      12'h8D7: dout  = 8'b00000000; // 2263 :   0 - 0x0
      12'h8D8: dout  = 8'b00000000; // 2264 :   0 - 0x0 -- Background 0x1b
      12'h8D9: dout  = 8'b00000000; // 2265 :   0 - 0x0
      12'h8DA: dout  = 8'b00000000; // 2266 :   0 - 0x0
      12'h8DB: dout  = 8'b00000000; // 2267 :   0 - 0x0
      12'h8DC: dout  = 8'b00000000; // 2268 :   0 - 0x0
      12'h8DD: dout  = 8'b00000000; // 2269 :   0 - 0x0
      12'h8DE: dout  = 8'b00000000; // 2270 :   0 - 0x0
      12'h8DF: dout  = 8'b00000000; // 2271 :   0 - 0x0
      12'h8E0: dout  = 8'b00000000; // 2272 :   0 - 0x0 -- Background 0x1c
      12'h8E1: dout  = 8'b00000000; // 2273 :   0 - 0x0
      12'h8E2: dout  = 8'b00000000; // 2274 :   0 - 0x0
      12'h8E3: dout  = 8'b00000000; // 2275 :   0 - 0x0
      12'h8E4: dout  = 8'b00000000; // 2276 :   0 - 0x0
      12'h8E5: dout  = 8'b00000000; // 2277 :   0 - 0x0
      12'h8E6: dout  = 8'b00000000; // 2278 :   0 - 0x0
      12'h8E7: dout  = 8'b00000000; // 2279 :   0 - 0x0
      12'h8E8: dout  = 8'b00000000; // 2280 :   0 - 0x0 -- Background 0x1d
      12'h8E9: dout  = 8'b00000000; // 2281 :   0 - 0x0
      12'h8EA: dout  = 8'b00000000; // 2282 :   0 - 0x0
      12'h8EB: dout  = 8'b00000000; // 2283 :   0 - 0x0
      12'h8EC: dout  = 8'b00000000; // 2284 :   0 - 0x0
      12'h8ED: dout  = 8'b00000000; // 2285 :   0 - 0x0
      12'h8EE: dout  = 8'b00000000; // 2286 :   0 - 0x0
      12'h8EF: dout  = 8'b00000000; // 2287 :   0 - 0x0
      12'h8F0: dout  = 8'b00000000; // 2288 :   0 - 0x0 -- Background 0x1e
      12'h8F1: dout  = 8'b00000000; // 2289 :   0 - 0x0
      12'h8F2: dout  = 8'b00000000; // 2290 :   0 - 0x0
      12'h8F3: dout  = 8'b00000000; // 2291 :   0 - 0x0
      12'h8F4: dout  = 8'b00000000; // 2292 :   0 - 0x0
      12'h8F5: dout  = 8'b00000000; // 2293 :   0 - 0x0
      12'h8F6: dout  = 8'b00000000; // 2294 :   0 - 0x0
      12'h8F7: dout  = 8'b00000000; // 2295 :   0 - 0x0
      12'h8F8: dout  = 8'b00000000; // 2296 :   0 - 0x0 -- Background 0x1f
      12'h8F9: dout  = 8'b00000000; // 2297 :   0 - 0x0
      12'h8FA: dout  = 8'b00000000; // 2298 :   0 - 0x0
      12'h8FB: dout  = 8'b00000000; // 2299 :   0 - 0x0
      12'h8FC: dout  = 8'b00000000; // 2300 :   0 - 0x0
      12'h8FD: dout  = 8'b00000000; // 2301 :   0 - 0x0
      12'h8FE: dout  = 8'b00000000; // 2302 :   0 - 0x0
      12'h8FF: dout  = 8'b00000000; // 2303 :   0 - 0x0
      12'h900: dout  = 8'b00000000; // 2304 :   0 - 0x0 -- Background 0x20
      12'h901: dout  = 8'b00000000; // 2305 :   0 - 0x0
      12'h902: dout  = 8'b00000000; // 2306 :   0 - 0x0
      12'h903: dout  = 8'b00000000; // 2307 :   0 - 0x0
      12'h904: dout  = 8'b00000000; // 2308 :   0 - 0x0
      12'h905: dout  = 8'b00000000; // 2309 :   0 - 0x0
      12'h906: dout  = 8'b00000000; // 2310 :   0 - 0x0
      12'h907: dout  = 8'b00000000; // 2311 :   0 - 0x0
      12'h908: dout  = 8'b00000000; // 2312 :   0 - 0x0 -- Background 0x21
      12'h909: dout  = 8'b00000000; // 2313 :   0 - 0x0
      12'h90A: dout  = 8'b00000000; // 2314 :   0 - 0x0
      12'h90B: dout  = 8'b00000000; // 2315 :   0 - 0x0
      12'h90C: dout  = 8'b00000000; // 2316 :   0 - 0x0
      12'h90D: dout  = 8'b00000000; // 2317 :   0 - 0x0
      12'h90E: dout  = 8'b00000000; // 2318 :   0 - 0x0
      12'h90F: dout  = 8'b00000000; // 2319 :   0 - 0x0
      12'h910: dout  = 8'b00000000; // 2320 :   0 - 0x0 -- Background 0x22
      12'h911: dout  = 8'b00000000; // 2321 :   0 - 0x0
      12'h912: dout  = 8'b00000000; // 2322 :   0 - 0x0
      12'h913: dout  = 8'b00000000; // 2323 :   0 - 0x0
      12'h914: dout  = 8'b00000000; // 2324 :   0 - 0x0
      12'h915: dout  = 8'b00000000; // 2325 :   0 - 0x0
      12'h916: dout  = 8'b00000000; // 2326 :   0 - 0x0
      12'h917: dout  = 8'b00000000; // 2327 :   0 - 0x0
      12'h918: dout  = 8'b00000000; // 2328 :   0 - 0x0 -- Background 0x23
      12'h919: dout  = 8'b00000000; // 2329 :   0 - 0x0
      12'h91A: dout  = 8'b00000000; // 2330 :   0 - 0x0
      12'h91B: dout  = 8'b00000000; // 2331 :   0 - 0x0
      12'h91C: dout  = 8'b00000000; // 2332 :   0 - 0x0
      12'h91D: dout  = 8'b00000000; // 2333 :   0 - 0x0
      12'h91E: dout  = 8'b00000000; // 2334 :   0 - 0x0
      12'h91F: dout  = 8'b00000000; // 2335 :   0 - 0x0
      12'h920: dout  = 8'b00000000; // 2336 :   0 - 0x0 -- Background 0x24
      12'h921: dout  = 8'b00000000; // 2337 :   0 - 0x0
      12'h922: dout  = 8'b00000000; // 2338 :   0 - 0x0
      12'h923: dout  = 8'b00000000; // 2339 :   0 - 0x0
      12'h924: dout  = 8'b00000000; // 2340 :   0 - 0x0
      12'h925: dout  = 8'b00000000; // 2341 :   0 - 0x0
      12'h926: dout  = 8'b00000000; // 2342 :   0 - 0x0
      12'h927: dout  = 8'b00000000; // 2343 :   0 - 0x0
      12'h928: dout  = 8'b00000000; // 2344 :   0 - 0x0 -- Background 0x25
      12'h929: dout  = 8'b00000000; // 2345 :   0 - 0x0
      12'h92A: dout  = 8'b00000000; // 2346 :   0 - 0x0
      12'h92B: dout  = 8'b00000000; // 2347 :   0 - 0x0
      12'h92C: dout  = 8'b00000000; // 2348 :   0 - 0x0
      12'h92D: dout  = 8'b00000000; // 2349 :   0 - 0x0
      12'h92E: dout  = 8'b00000000; // 2350 :   0 - 0x0
      12'h92F: dout  = 8'b00000000; // 2351 :   0 - 0x0
      12'h930: dout  = 8'b11111111; // 2352 : 255 - 0xff -- Background 0x26
      12'h931: dout  = 8'b11111111; // 2353 : 255 - 0xff
      12'h932: dout  = 8'b11111111; // 2354 : 255 - 0xff
      12'h933: dout  = 8'b11111111; // 2355 : 255 - 0xff
      12'h934: dout  = 8'b11111111; // 2356 : 255 - 0xff
      12'h935: dout  = 8'b11111111; // 2357 : 255 - 0xff
      12'h936: dout  = 8'b11111111; // 2358 : 255 - 0xff
      12'h937: dout  = 8'b11111111; // 2359 : 255 - 0xff
      12'h938: dout  = 8'b11111111; // 2360 : 255 - 0xff -- Background 0x27
      12'h939: dout  = 8'b11111111; // 2361 : 255 - 0xff
      12'h93A: dout  = 8'b11111111; // 2362 : 255 - 0xff
      12'h93B: dout  = 8'b11111111; // 2363 : 255 - 0xff
      12'h93C: dout  = 8'b11111111; // 2364 : 255 - 0xff
      12'h93D: dout  = 8'b11111111; // 2365 : 255 - 0xff
      12'h93E: dout  = 8'b11111111; // 2366 : 255 - 0xff
      12'h93F: dout  = 8'b11111111; // 2367 : 255 - 0xff
      12'h940: dout  = 8'b00000000; // 2368 :   0 - 0x0 -- Background 0x28
      12'h941: dout  = 8'b00000000; // 2369 :   0 - 0x0
      12'h942: dout  = 8'b00000000; // 2370 :   0 - 0x0
      12'h943: dout  = 8'b00000000; // 2371 :   0 - 0x0
      12'h944: dout  = 8'b00000000; // 2372 :   0 - 0x0
      12'h945: dout  = 8'b00000000; // 2373 :   0 - 0x0
      12'h946: dout  = 8'b00000000; // 2374 :   0 - 0x0
      12'h947: dout  = 8'b00000000; // 2375 :   0 - 0x0
      12'h948: dout  = 8'b00000000; // 2376 :   0 - 0x0 -- Background 0x29
      12'h949: dout  = 8'b00000000; // 2377 :   0 - 0x0
      12'h94A: dout  = 8'b00000000; // 2378 :   0 - 0x0
      12'h94B: dout  = 8'b00000000; // 2379 :   0 - 0x0
      12'h94C: dout  = 8'b00000000; // 2380 :   0 - 0x0
      12'h94D: dout  = 8'b00000000; // 2381 :   0 - 0x0
      12'h94E: dout  = 8'b00000000; // 2382 :   0 - 0x0
      12'h94F: dout  = 8'b00000000; // 2383 :   0 - 0x0
      12'h950: dout  = 8'b01111111; // 2384 : 127 - 0x7f -- Background 0x2a
      12'h951: dout  = 8'b01111111; // 2385 : 127 - 0x7f
      12'h952: dout  = 8'b01111111; // 2386 : 127 - 0x7f
      12'h953: dout  = 8'b01111111; // 2387 : 127 - 0x7f
      12'h954: dout  = 8'b01111111; // 2388 : 127 - 0x7f
      12'h955: dout  = 8'b01111111; // 2389 : 127 - 0x7f
      12'h956: dout  = 8'b01111111; // 2390 : 127 - 0x7f
      12'h957: dout  = 8'b01111111; // 2391 : 127 - 0x7f
      12'h958: dout  = 8'b00000000; // 2392 :   0 - 0x0 -- Background 0x2b
      12'h959: dout  = 8'b00000000; // 2393 :   0 - 0x0
      12'h95A: dout  = 8'b00000000; // 2394 :   0 - 0x0
      12'h95B: dout  = 8'b00000000; // 2395 :   0 - 0x0
      12'h95C: dout  = 8'b00000000; // 2396 :   0 - 0x0
      12'h95D: dout  = 8'b00000000; // 2397 :   0 - 0x0
      12'h95E: dout  = 8'b00000000; // 2398 :   0 - 0x0
      12'h95F: dout  = 8'b00000000; // 2399 :   0 - 0x0
      12'h960: dout  = 8'b11111111; // 2400 : 255 - 0xff -- Background 0x2c
      12'h961: dout  = 8'b10000000; // 2401 : 128 - 0x80
      12'h962: dout  = 8'b10000000; // 2402 : 128 - 0x80
      12'h963: dout  = 8'b10000000; // 2403 : 128 - 0x80
      12'h964: dout  = 8'b10000000; // 2404 : 128 - 0x80
      12'h965: dout  = 8'b00000000; // 2405 :   0 - 0x0
      12'h966: dout  = 8'b00011100; // 2406 :  28 - 0x1c
      12'h967: dout  = 8'b00111110; // 2407 :  62 - 0x3e
      12'h968: dout  = 8'b01111111; // 2408 : 127 - 0x7f -- Background 0x2d
      12'h969: dout  = 8'b01111111; // 2409 : 127 - 0x7f
      12'h96A: dout  = 8'b01111111; // 2410 : 127 - 0x7f
      12'h96B: dout  = 8'b00111110; // 2411 :  62 - 0x3e
      12'h96C: dout  = 8'b00011100; // 2412 :  28 - 0x1c
      12'h96D: dout  = 8'b00000000; // 2413 :   0 - 0x0
      12'h96E: dout  = 8'b00000000; // 2414 :   0 - 0x0
      12'h96F: dout  = 8'b11111111; // 2415 : 255 - 0xff
      12'h970: dout  = 8'b00001000; // 2416 :   8 - 0x8 -- Background 0x2e
      12'h971: dout  = 8'b00000100; // 2417 :   4 - 0x4
      12'h972: dout  = 8'b00000100; // 2418 :   4 - 0x4
      12'h973: dout  = 8'b00000100; // 2419 :   4 - 0x4
      12'h974: dout  = 8'b00000100; // 2420 :   4 - 0x4
      12'h975: dout  = 8'b00000100; // 2421 :   4 - 0x4
      12'h976: dout  = 8'b00001000; // 2422 :   8 - 0x8
      12'h977: dout  = 8'b00000000; // 2423 :   0 - 0x0
      12'h978: dout  = 8'b00000011; // 2424 :   3 - 0x3 -- Background 0x2f
      12'h979: dout  = 8'b00000101; // 2425 :   5 - 0x5
      12'h97A: dout  = 8'b00001011; // 2426 :  11 - 0xb
      12'h97B: dout  = 8'b00001011; // 2427 :  11 - 0xb
      12'h97C: dout  = 8'b00001111; // 2428 :  15 - 0xf
      12'h97D: dout  = 8'b00001111; // 2429 :  15 - 0xf
      12'h97E: dout  = 8'b00000111; // 2430 :   7 - 0x7
      12'h97F: dout  = 8'b00000011; // 2431 :   3 - 0x3
      12'h980: dout  = 8'b00000001; // 2432 :   1 - 0x1 -- Background 0x30
      12'h981: dout  = 8'b00000011; // 2433 :   3 - 0x3
      12'h982: dout  = 8'b00000111; // 2434 :   7 - 0x7
      12'h983: dout  = 8'b00001111; // 2435 :  15 - 0xf
      12'h984: dout  = 8'b00011111; // 2436 :  31 - 0x1f
      12'h985: dout  = 8'b00111111; // 2437 :  63 - 0x3f
      12'h986: dout  = 8'b01111111; // 2438 : 127 - 0x7f
      12'h987: dout  = 8'b11111111; // 2439 : 255 - 0xff
      12'h988: dout  = 8'b00000000; // 2440 :   0 - 0x0 -- Background 0x31
      12'h989: dout  = 8'b00000000; // 2441 :   0 - 0x0
      12'h98A: dout  = 8'b00000000; // 2442 :   0 - 0x0
      12'h98B: dout  = 8'b00000000; // 2443 :   0 - 0x0
      12'h98C: dout  = 8'b00000000; // 2444 :   0 - 0x0
      12'h98D: dout  = 8'b00000111; // 2445 :   7 - 0x7
      12'h98E: dout  = 8'b00111111; // 2446 :  63 - 0x3f
      12'h98F: dout  = 8'b11111111; // 2447 : 255 - 0xff
      12'h990: dout  = 8'b00000000; // 2448 :   0 - 0x0 -- Background 0x32
      12'h991: dout  = 8'b00000000; // 2449 :   0 - 0x0
      12'h992: dout  = 8'b00000000; // 2450 :   0 - 0x0
      12'h993: dout  = 8'b00000000; // 2451 :   0 - 0x0
      12'h994: dout  = 8'b00000000; // 2452 :   0 - 0x0
      12'h995: dout  = 8'b11100000; // 2453 : 224 - 0xe0
      12'h996: dout  = 8'b11111100; // 2454 : 252 - 0xfc
      12'h997: dout  = 8'b11111111; // 2455 : 255 - 0xff
      12'h998: dout  = 8'b10000000; // 2456 : 128 - 0x80 -- Background 0x33
      12'h999: dout  = 8'b11000000; // 2457 : 192 - 0xc0
      12'h99A: dout  = 8'b11100000; // 2458 : 224 - 0xe0
      12'h99B: dout  = 8'b11110000; // 2459 : 240 - 0xf0
      12'h99C: dout  = 8'b11111000; // 2460 : 248 - 0xf8
      12'h99D: dout  = 8'b11111100; // 2461 : 252 - 0xfc
      12'h99E: dout  = 8'b11111110; // 2462 : 254 - 0xfe
      12'h99F: dout  = 8'b11111111; // 2463 : 255 - 0xff
      12'h9A0: dout  = 8'b11111111; // 2464 : 255 - 0xff -- Background 0x34
      12'h9A1: dout  = 8'b11111111; // 2465 : 255 - 0xff
      12'h9A2: dout  = 8'b11111111; // 2466 : 255 - 0xff
      12'h9A3: dout  = 8'b11111111; // 2467 : 255 - 0xff
      12'h9A4: dout  = 8'b11111111; // 2468 : 255 - 0xff
      12'h9A5: dout  = 8'b11111111; // 2469 : 255 - 0xff
      12'h9A6: dout  = 8'b11111111; // 2470 : 255 - 0xff
      12'h9A7: dout  = 8'b11111111; // 2471 : 255 - 0xff
      12'h9A8: dout  = 8'b00000111; // 2472 :   7 - 0x7 -- Background 0x35
      12'h9A9: dout  = 8'b00001000; // 2473 :   8 - 0x8
      12'h9AA: dout  = 8'b00010000; // 2474 :  16 - 0x10
      12'h9AB: dout  = 8'b00000000; // 2475 :   0 - 0x0
      12'h9AC: dout  = 8'b01100000; // 2476 :  96 - 0x60
      12'h9AD: dout  = 8'b10000000; // 2477 : 128 - 0x80
      12'h9AE: dout  = 8'b10000000; // 2478 : 128 - 0x80
      12'h9AF: dout  = 8'b01000000; // 2479 :  64 - 0x40
      12'h9B0: dout  = 8'b00000011; // 2480 :   3 - 0x3 -- Background 0x36
      12'h9B1: dout  = 8'b00000100; // 2481 :   4 - 0x4
      12'h9B2: dout  = 8'b00011000; // 2482 :  24 - 0x18
      12'h9B3: dout  = 8'b00100000; // 2483 :  32 - 0x20
      12'h9B4: dout  = 8'b00100000; // 2484 :  32 - 0x20
      12'h9B5: dout  = 8'b00100000; // 2485 :  32 - 0x20
      12'h9B6: dout  = 8'b01000110; // 2486 :  70 - 0x46
      12'h9B7: dout  = 8'b10001000; // 2487 : 136 - 0x88
      12'h9B8: dout  = 8'b11000000; // 2488 : 192 - 0xc0 -- Background 0x37
      12'h9B9: dout  = 8'b00100000; // 2489 :  32 - 0x20
      12'h9BA: dout  = 8'b00010000; // 2490 :  16 - 0x10
      12'h9BB: dout  = 8'b00010100; // 2491 :  20 - 0x14
      12'h9BC: dout  = 8'b00001010; // 2492 :  10 - 0xa
      12'h9BD: dout  = 8'b01000001; // 2493 :  65 - 0x41
      12'h9BE: dout  = 8'b00100001; // 2494 :  33 - 0x21
      12'h9BF: dout  = 8'b00000001; // 2495 :   1 - 0x1
      12'h9C0: dout  = 8'b10010000; // 2496 : 144 - 0x90 -- Background 0x38
      12'h9C1: dout  = 8'b10101000; // 2497 : 168 - 0xa8
      12'h9C2: dout  = 8'b01001000; // 2498 :  72 - 0x48
      12'h9C3: dout  = 8'b00001010; // 2499 :  10 - 0xa
      12'h9C4: dout  = 8'b00000101; // 2500 :   5 - 0x5
      12'h9C5: dout  = 8'b00000001; // 2501 :   1 - 0x1
      12'h9C6: dout  = 8'b00000001; // 2502 :   1 - 0x1
      12'h9C7: dout  = 8'b00000010; // 2503 :   2 - 0x2
      12'h9C8: dout  = 8'b00100100; // 2504 :  36 - 0x24 -- Background 0x39
      12'h9C9: dout  = 8'b00010010; // 2505 :  18 - 0x12
      12'h9CA: dout  = 8'b00001001; // 2506 :   9 - 0x9
      12'h9CB: dout  = 8'b00001000; // 2507 :   8 - 0x8
      12'h9CC: dout  = 8'b00000111; // 2508 :   7 - 0x7
      12'h9CD: dout  = 8'b00000000; // 2509 :   0 - 0x0
      12'h9CE: dout  = 8'b00000000; // 2510 :   0 - 0x0
      12'h9CF: dout  = 8'b00000000; // 2511 :   0 - 0x0
      12'h9D0: dout  = 8'b00000000; // 2512 :   0 - 0x0 -- Background 0x3a
      12'h9D1: dout  = 8'b01000000; // 2513 :  64 - 0x40
      12'h9D2: dout  = 8'b11100011; // 2514 : 227 - 0xe3
      12'h9D3: dout  = 8'b00111111; // 2515 :  63 - 0x3f
      12'h9D4: dout  = 8'b00001100; // 2516 :  12 - 0xc
      12'h9D5: dout  = 8'b10000001; // 2517 : 129 - 0x81
      12'h9D6: dout  = 8'b01100010; // 2518 :  98 - 0x62
      12'h9D7: dout  = 8'b00011100; // 2519 :  28 - 0x1c
      12'h9D8: dout  = 8'b01000000; // 2520 :  64 - 0x40 -- Background 0x3b
      12'h9D9: dout  = 8'b10000000; // 2521 : 128 - 0x80
      12'h9DA: dout  = 8'b11000010; // 2522 : 194 - 0xc2
      12'h9DB: dout  = 8'b01111100; // 2523 : 124 - 0x7c
      12'h9DC: dout  = 8'b00111000; // 2524 :  56 - 0x38
      12'h9DD: dout  = 8'b00000000; // 2525 :   0 - 0x0
      12'h9DE: dout  = 8'b11000011; // 2526 : 195 - 0xc3
      12'h9DF: dout  = 8'b00111100; // 2527 :  60 - 0x3c
      12'h9E0: dout  = 8'b00000100; // 2528 :   4 - 0x4 -- Background 0x3c
      12'h9E1: dout  = 8'b00000010; // 2529 :   2 - 0x2
      12'h9E2: dout  = 8'b00000001; // 2530 :   1 - 0x1
      12'h9E3: dout  = 8'b00000000; // 2531 :   0 - 0x0
      12'h9E4: dout  = 8'b00000110; // 2532 :   6 - 0x6
      12'h9E5: dout  = 8'b10011000; // 2533 : 152 - 0x98
      12'h9E6: dout  = 8'b01100000; // 2534 :  96 - 0x60
      12'h9E7: dout  = 8'b00000000; // 2535 :   0 - 0x0
      12'h9E8: dout  = 8'b11000000; // 2536 : 192 - 0xc0 -- Background 0x3d
      12'h9E9: dout  = 8'b11100000; // 2537 : 224 - 0xe0
      12'h9EA: dout  = 8'b11110000; // 2538 : 240 - 0xf0
      12'h9EB: dout  = 8'b11110000; // 2539 : 240 - 0xf0
      12'h9EC: dout  = 8'b11110000; // 2540 : 240 - 0xf0
      12'h9ED: dout  = 8'b11110000; // 2541 : 240 - 0xf0
      12'h9EE: dout  = 8'b11100000; // 2542 : 224 - 0xe0
      12'h9EF: dout  = 8'b11000000; // 2543 : 192 - 0xc0
      12'h9F0: dout  = 8'b00000000; // 2544 :   0 - 0x0 -- Background 0x3e
      12'h9F1: dout  = 8'b00000000; // 2545 :   0 - 0x0
      12'h9F2: dout  = 8'b00000000; // 2546 :   0 - 0x0
      12'h9F3: dout  = 8'b00000000; // 2547 :   0 - 0x0
      12'h9F4: dout  = 8'b00000000; // 2548 :   0 - 0x0
      12'h9F5: dout  = 8'b00000000; // 2549 :   0 - 0x0
      12'h9F6: dout  = 8'b00011100; // 2550 :  28 - 0x1c
      12'h9F7: dout  = 8'b00111110; // 2551 :  62 - 0x3e
      12'h9F8: dout  = 8'b01111111; // 2552 : 127 - 0x7f -- Background 0x3f
      12'h9F9: dout  = 8'b01111111; // 2553 : 127 - 0x7f
      12'h9FA: dout  = 8'b01111111; // 2554 : 127 - 0x7f
      12'h9FB: dout  = 8'b00111110; // 2555 :  62 - 0x3e
      12'h9FC: dout  = 8'b00011100; // 2556 :  28 - 0x1c
      12'h9FD: dout  = 8'b00000000; // 2557 :   0 - 0x0
      12'h9FE: dout  = 8'b00000000; // 2558 :   0 - 0x0
      12'h9FF: dout  = 8'b00000000; // 2559 :   0 - 0x0
      12'hA00: dout  = 8'b11111111; // 2560 : 255 - 0xff -- Background 0x40
      12'hA01: dout  = 8'b11111111; // 2561 : 255 - 0xff
      12'hA02: dout  = 8'b11111111; // 2562 : 255 - 0xff
      12'hA03: dout  = 8'b11111111; // 2563 : 255 - 0xff
      12'hA04: dout  = 8'b11111111; // 2564 : 255 - 0xff
      12'hA05: dout  = 8'b11111111; // 2565 : 255 - 0xff
      12'hA06: dout  = 8'b11111111; // 2566 : 255 - 0xff
      12'hA07: dout  = 8'b11111111; // 2567 : 255 - 0xff
      12'hA08: dout  = 8'b00000000; // 2568 :   0 - 0x0 -- Background 0x41
      12'hA09: dout  = 8'b00001000; // 2569 :   8 - 0x8
      12'hA0A: dout  = 8'b00011000; // 2570 :  24 - 0x18
      12'hA0B: dout  = 8'b00111000; // 2571 :  56 - 0x38
      12'hA0C: dout  = 8'b11111100; // 2572 : 252 - 0xfc
      12'hA0D: dout  = 8'b10111111; // 2573 : 191 - 0xbf
      12'hA0E: dout  = 8'b01011110; // 2574 :  94 - 0x5e
      12'hA0F: dout  = 8'b11011001; // 2575 : 217 - 0xd9
      12'hA10: dout  = 8'b10000001; // 2576 : 129 - 0x81 -- Background 0x42
      12'hA11: dout  = 8'b10000001; // 2577 : 129 - 0x81
      12'hA12: dout  = 8'b10000001; // 2578 : 129 - 0x81
      12'hA13: dout  = 8'b10000001; // 2579 : 129 - 0x81
      12'hA14: dout  = 8'b10000001; // 2580 : 129 - 0x81
      12'hA15: dout  = 8'b10000001; // 2581 : 129 - 0x81
      12'hA16: dout  = 8'b10000001; // 2582 : 129 - 0x81
      12'hA17: dout  = 8'b10000001; // 2583 : 129 - 0x81
      12'hA18: dout  = 8'b00000001; // 2584 :   1 - 0x1 -- Background 0x43
      12'hA19: dout  = 8'b00000001; // 2585 :   1 - 0x1
      12'hA1A: dout  = 8'b00000001; // 2586 :   1 - 0x1
      12'hA1B: dout  = 8'b00000001; // 2587 :   1 - 0x1
      12'hA1C: dout  = 8'b00000001; // 2588 :   1 - 0x1
      12'hA1D: dout  = 8'b00000001; // 2589 :   1 - 0x1
      12'hA1E: dout  = 8'b00000001; // 2590 :   1 - 0x1
      12'hA1F: dout  = 8'b00000001; // 2591 :   1 - 0x1
      12'hA20: dout  = 8'b00000000; // 2592 :   0 - 0x0 -- Background 0x44
      12'hA21: dout  = 8'b01111111; // 2593 : 127 - 0x7f
      12'hA22: dout  = 8'b01111111; // 2594 : 127 - 0x7f
      12'hA23: dout  = 8'b01100111; // 2595 : 103 - 0x67
      12'hA24: dout  = 8'b01100111; // 2596 : 103 - 0x67
      12'hA25: dout  = 8'b01111111; // 2597 : 127 - 0x7f
      12'hA26: dout  = 8'b01111111; // 2598 : 127 - 0x7f
      12'hA27: dout  = 8'b01111111; // 2599 : 127 - 0x7f
      12'hA28: dout  = 8'b00000000; // 2600 :   0 - 0x0 -- Background 0x45
      12'hA29: dout  = 8'b11111111; // 2601 : 255 - 0xff
      12'hA2A: dout  = 8'b11111111; // 2602 : 255 - 0xff
      12'hA2B: dout  = 8'b11111111; // 2603 : 255 - 0xff
      12'hA2C: dout  = 8'b11111111; // 2604 : 255 - 0xff
      12'hA2D: dout  = 8'b11111111; // 2605 : 255 - 0xff
      12'hA2E: dout  = 8'b11111111; // 2606 : 255 - 0xff
      12'hA2F: dout  = 8'b11111111; // 2607 : 255 - 0xff
      12'hA30: dout  = 8'b01111111; // 2608 : 127 - 0x7f -- Background 0x46
      12'hA31: dout  = 8'b01111111; // 2609 : 127 - 0x7f
      12'hA32: dout  = 8'b01111111; // 2610 : 127 - 0x7f
      12'hA33: dout  = 8'b01111111; // 2611 : 127 - 0x7f
      12'hA34: dout  = 8'b01111111; // 2612 : 127 - 0x7f
      12'hA35: dout  = 8'b01111111; // 2613 : 127 - 0x7f
      12'hA36: dout  = 8'b01111111; // 2614 : 127 - 0x7f
      12'hA37: dout  = 8'b01111111; // 2615 : 127 - 0x7f
      12'hA38: dout  = 8'b11111111; // 2616 : 255 - 0xff -- Background 0x47
      12'hA39: dout  = 8'b11111111; // 2617 : 255 - 0xff
      12'hA3A: dout  = 8'b11111111; // 2618 : 255 - 0xff
      12'hA3B: dout  = 8'b11111111; // 2619 : 255 - 0xff
      12'hA3C: dout  = 8'b11111111; // 2620 : 255 - 0xff
      12'hA3D: dout  = 8'b11111111; // 2621 : 255 - 0xff
      12'hA3E: dout  = 8'b11111111; // 2622 : 255 - 0xff
      12'hA3F: dout  = 8'b11111111; // 2623 : 255 - 0xff
      12'hA40: dout  = 8'b00000000; // 2624 :   0 - 0x0 -- Background 0x48
      12'hA41: dout  = 8'b11111111; // 2625 : 255 - 0xff
      12'hA42: dout  = 8'b11111111; // 2626 : 255 - 0xff
      12'hA43: dout  = 8'b11111111; // 2627 : 255 - 0xff
      12'hA44: dout  = 8'b11111111; // 2628 : 255 - 0xff
      12'hA45: dout  = 8'b11111111; // 2629 : 255 - 0xff
      12'hA46: dout  = 8'b11111111; // 2630 : 255 - 0xff
      12'hA47: dout  = 8'b11111111; // 2631 : 255 - 0xff
      12'hA48: dout  = 8'b00000000; // 2632 :   0 - 0x0 -- Background 0x49
      12'hA49: dout  = 8'b11111111; // 2633 : 255 - 0xff
      12'hA4A: dout  = 8'b11111111; // 2634 : 255 - 0xff
      12'hA4B: dout  = 8'b11100111; // 2635 : 231 - 0xe7
      12'hA4C: dout  = 8'b11100111; // 2636 : 231 - 0xe7
      12'hA4D: dout  = 8'b11111111; // 2637 : 255 - 0xff
      12'hA4E: dout  = 8'b11111111; // 2638 : 255 - 0xff
      12'hA4F: dout  = 8'b11111111; // 2639 : 255 - 0xff
      12'hA50: dout  = 8'b11111111; // 2640 : 255 - 0xff -- Background 0x4a
      12'hA51: dout  = 8'b11111111; // 2641 : 255 - 0xff
      12'hA52: dout  = 8'b11111111; // 2642 : 255 - 0xff
      12'hA53: dout  = 8'b11111111; // 2643 : 255 - 0xff
      12'hA54: dout  = 8'b11111111; // 2644 : 255 - 0xff
      12'hA55: dout  = 8'b11111111; // 2645 : 255 - 0xff
      12'hA56: dout  = 8'b11111111; // 2646 : 255 - 0xff
      12'hA57: dout  = 8'b11111111; // 2647 : 255 - 0xff
      12'hA58: dout  = 8'b00111111; // 2648 :  63 - 0x3f -- Background 0x4b
      12'hA59: dout  = 8'b01100000; // 2649 :  96 - 0x60
      12'hA5A: dout  = 8'b01000000; // 2650 :  64 - 0x40
      12'hA5B: dout  = 8'b11000000; // 2651 : 192 - 0xc0
      12'hA5C: dout  = 8'b10000000; // 2652 : 128 - 0x80
      12'hA5D: dout  = 8'b10000000; // 2653 : 128 - 0x80
      12'hA5E: dout  = 8'b10000000; // 2654 : 128 - 0x80
      12'hA5F: dout  = 8'b10000000; // 2655 : 128 - 0x80
      12'hA60: dout  = 8'b10000000; // 2656 : 128 - 0x80 -- Background 0x4c
      12'hA61: dout  = 8'b10000000; // 2657 : 128 - 0x80
      12'hA62: dout  = 8'b10000000; // 2658 : 128 - 0x80
      12'hA63: dout  = 8'b10000000; // 2659 : 128 - 0x80
      12'hA64: dout  = 8'b10000000; // 2660 : 128 - 0x80
      12'hA65: dout  = 8'b10000001; // 2661 : 129 - 0x81
      12'hA66: dout  = 8'b01000010; // 2662 :  66 - 0x42
      12'hA67: dout  = 8'b00111100; // 2663 :  60 - 0x3c
      12'hA68: dout  = 8'b11111111; // 2664 : 255 - 0xff -- Background 0x4d
      12'hA69: dout  = 8'b00000000; // 2665 :   0 - 0x0
      12'hA6A: dout  = 8'b00000000; // 2666 :   0 - 0x0
      12'hA6B: dout  = 8'b00000000; // 2667 :   0 - 0x0
      12'hA6C: dout  = 8'b00000000; // 2668 :   0 - 0x0
      12'hA6D: dout  = 8'b00000000; // 2669 :   0 - 0x0
      12'hA6E: dout  = 8'b00000000; // 2670 :   0 - 0x0
      12'hA6F: dout  = 8'b00000000; // 2671 :   0 - 0x0
      12'hA70: dout  = 8'b00000000; // 2672 :   0 - 0x0 -- Background 0x4e
      12'hA71: dout  = 8'b00000000; // 2673 :   0 - 0x0
      12'hA72: dout  = 8'b00000000; // 2674 :   0 - 0x0
      12'hA73: dout  = 8'b00000000; // 2675 :   0 - 0x0
      12'hA74: dout  = 8'b00000000; // 2676 :   0 - 0x0
      12'hA75: dout  = 8'b00000001; // 2677 :   1 - 0x1
      12'hA76: dout  = 8'b10000010; // 2678 : 130 - 0x82
      12'hA77: dout  = 8'b01111100; // 2679 : 124 - 0x7c
      12'hA78: dout  = 8'b00000000; // 2680 :   0 - 0x0 -- Background 0x4f
      12'hA79: dout  = 8'b00000000; // 2681 :   0 - 0x0
      12'hA7A: dout  = 8'b00000000; // 2682 :   0 - 0x0
      12'hA7B: dout  = 8'b00000000; // 2683 :   0 - 0x0
      12'hA7C: dout  = 8'b00000000; // 2684 :   0 - 0x0
      12'hA7D: dout  = 8'b00000001; // 2685 :   1 - 0x1
      12'hA7E: dout  = 8'b10000011; // 2686 : 131 - 0x83
      12'hA7F: dout  = 8'b11111111; // 2687 : 255 - 0xff
      12'hA80: dout  = 8'b11111000; // 2688 : 248 - 0xf8 -- Background 0x50
      12'hA81: dout  = 8'b00000100; // 2689 :   4 - 0x4
      12'hA82: dout  = 8'b00000010; // 2690 :   2 - 0x2
      12'hA83: dout  = 8'b00000010; // 2691 :   2 - 0x2
      12'hA84: dout  = 8'b00000001; // 2692 :   1 - 0x1
      12'hA85: dout  = 8'b00000001; // 2693 :   1 - 0x1
      12'hA86: dout  = 8'b00000001; // 2694 :   1 - 0x1
      12'hA87: dout  = 8'b00000001; // 2695 :   1 - 0x1
      12'hA88: dout  = 8'b00000001; // 2696 :   1 - 0x1 -- Background 0x51
      12'hA89: dout  = 8'b00000001; // 2697 :   1 - 0x1
      12'hA8A: dout  = 8'b00000001; // 2698 :   1 - 0x1
      12'hA8B: dout  = 8'b00000001; // 2699 :   1 - 0x1
      12'hA8C: dout  = 8'b00000001; // 2700 :   1 - 0x1
      12'hA8D: dout  = 8'b10000001; // 2701 : 129 - 0x81
      12'hA8E: dout  = 8'b01000010; // 2702 :  66 - 0x42
      12'hA8F: dout  = 8'b00111100; // 2703 :  60 - 0x3c
      12'hA90: dout  = 8'b11111111; // 2704 : 255 - 0xff -- Background 0x52
      12'hA91: dout  = 8'b11111111; // 2705 : 255 - 0xff
      12'hA92: dout  = 8'b11111111; // 2706 : 255 - 0xff
      12'hA93: dout  = 8'b11111111; // 2707 : 255 - 0xff
      12'hA94: dout  = 8'b11111111; // 2708 : 255 - 0xff
      12'hA95: dout  = 8'b11111111; // 2709 : 255 - 0xff
      12'hA96: dout  = 8'b11111111; // 2710 : 255 - 0xff
      12'hA97: dout  = 8'b11111111; // 2711 : 255 - 0xff
      12'hA98: dout  = 8'b01111111; // 2712 : 127 - 0x7f -- Background 0x53
      12'hA99: dout  = 8'b10000000; // 2713 : 128 - 0x80
      12'hA9A: dout  = 8'b10100000; // 2714 : 160 - 0xa0
      12'hA9B: dout  = 8'b10000111; // 2715 : 135 - 0x87
      12'hA9C: dout  = 8'b10001111; // 2716 : 143 - 0x8f
      12'hA9D: dout  = 8'b10001110; // 2717 : 142 - 0x8e
      12'hA9E: dout  = 8'b10001110; // 2718 : 142 - 0x8e
      12'hA9F: dout  = 8'b10000110; // 2719 : 134 - 0x86
      12'hAA0: dout  = 8'b11111110; // 2720 : 254 - 0xfe -- Background 0x54
      12'hAA1: dout  = 8'b00000001; // 2721 :   1 - 0x1
      12'hAA2: dout  = 8'b00000101; // 2722 :   5 - 0x5
      12'hAA3: dout  = 8'b11000001; // 2723 : 193 - 0xc1
      12'hAA4: dout  = 8'b11100001; // 2724 : 225 - 0xe1
      12'hAA5: dout  = 8'b01110001; // 2725 : 113 - 0x71
      12'hAA6: dout  = 8'b01110001; // 2726 : 113 - 0x71
      12'hAA7: dout  = 8'b11110001; // 2727 : 241 - 0xf1
      12'hAA8: dout  = 8'b10000001; // 2728 : 129 - 0x81 -- Background 0x55
      12'hAA9: dout  = 8'b10000001; // 2729 : 129 - 0x81
      12'hAAA: dout  = 8'b10000000; // 2730 : 128 - 0x80
      12'hAAB: dout  = 8'b10000001; // 2731 : 129 - 0x81
      12'hAAC: dout  = 8'b10000001; // 2732 : 129 - 0x81
      12'hAAD: dout  = 8'b10100000; // 2733 : 160 - 0xa0
      12'hAAE: dout  = 8'b10000000; // 2734 : 128 - 0x80
      12'hAAF: dout  = 8'b11111111; // 2735 : 255 - 0xff
      12'hAB0: dout  = 8'b11110001; // 2736 : 241 - 0xf1 -- Background 0x56
      12'hAB1: dout  = 8'b11000001; // 2737 : 193 - 0xc1
      12'hAB2: dout  = 8'b11000001; // 2738 : 193 - 0xc1
      12'hAB3: dout  = 8'b10000001; // 2739 : 129 - 0x81
      12'hAB4: dout  = 8'b11000001; // 2740 : 193 - 0xc1
      12'hAB5: dout  = 8'b11000101; // 2741 : 197 - 0xc5
      12'hAB6: dout  = 8'b00000001; // 2742 :   1 - 0x1
      12'hAB7: dout  = 8'b11111111; // 2743 : 255 - 0xff
      12'hAB8: dout  = 8'b01111111; // 2744 : 127 - 0x7f -- Background 0x57
      12'hAB9: dout  = 8'b11111111; // 2745 : 255 - 0xff
      12'hABA: dout  = 8'b11111111; // 2746 : 255 - 0xff
      12'hABB: dout  = 8'b11111111; // 2747 : 255 - 0xff
      12'hABC: dout  = 8'b11111111; // 2748 : 255 - 0xff
      12'hABD: dout  = 8'b11111111; // 2749 : 255 - 0xff
      12'hABE: dout  = 8'b11111111; // 2750 : 255 - 0xff
      12'hABF: dout  = 8'b11111111; // 2751 : 255 - 0xff
      12'hAC0: dout  = 8'b11111110; // 2752 : 254 - 0xfe -- Background 0x58
      12'hAC1: dout  = 8'b11111111; // 2753 : 255 - 0xff
      12'hAC2: dout  = 8'b11111111; // 2754 : 255 - 0xff
      12'hAC3: dout  = 8'b11111111; // 2755 : 255 - 0xff
      12'hAC4: dout  = 8'b11111111; // 2756 : 255 - 0xff
      12'hAC5: dout  = 8'b11111111; // 2757 : 255 - 0xff
      12'hAC6: dout  = 8'b11111111; // 2758 : 255 - 0xff
      12'hAC7: dout  = 8'b11111111; // 2759 : 255 - 0xff
      12'hAC8: dout  = 8'b11111111; // 2760 : 255 - 0xff -- Background 0x59
      12'hAC9: dout  = 8'b11111111; // 2761 : 255 - 0xff
      12'hACA: dout  = 8'b11111111; // 2762 : 255 - 0xff
      12'hACB: dout  = 8'b11111111; // 2763 : 255 - 0xff
      12'hACC: dout  = 8'b11111111; // 2764 : 255 - 0xff
      12'hACD: dout  = 8'b11111111; // 2765 : 255 - 0xff
      12'hACE: dout  = 8'b11111111; // 2766 : 255 - 0xff
      12'hACF: dout  = 8'b01111111; // 2767 : 127 - 0x7f
      12'hAD0: dout  = 8'b11111111; // 2768 : 255 - 0xff -- Background 0x5a
      12'hAD1: dout  = 8'b11111111; // 2769 : 255 - 0xff
      12'hAD2: dout  = 8'b11111111; // 2770 : 255 - 0xff
      12'hAD3: dout  = 8'b11111111; // 2771 : 255 - 0xff
      12'hAD4: dout  = 8'b11111111; // 2772 : 255 - 0xff
      12'hAD5: dout  = 8'b11111111; // 2773 : 255 - 0xff
      12'hAD6: dout  = 8'b11111111; // 2774 : 255 - 0xff
      12'hAD7: dout  = 8'b11111110; // 2775 : 254 - 0xfe
      12'hAD8: dout  = 8'b00000000; // 2776 :   0 - 0x0 -- Background 0x5b
      12'hAD9: dout  = 8'b00000000; // 2777 :   0 - 0x0
      12'hADA: dout  = 8'b00000000; // 2778 :   0 - 0x0
      12'hADB: dout  = 8'b00000000; // 2779 :   0 - 0x0
      12'hADC: dout  = 8'b00000000; // 2780 :   0 - 0x0
      12'hADD: dout  = 8'b00000000; // 2781 :   0 - 0x0
      12'hADE: dout  = 8'b00111000; // 2782 :  56 - 0x38
      12'hADF: dout  = 8'b01111100; // 2783 : 124 - 0x7c
      12'hAE0: dout  = 8'b11111110; // 2784 : 254 - 0xfe -- Background 0x5c
      12'hAE1: dout  = 8'b11111110; // 2785 : 254 - 0xfe
      12'hAE2: dout  = 8'b11111110; // 2786 : 254 - 0xfe
      12'hAE3: dout  = 8'b01111100; // 2787 : 124 - 0x7c
      12'hAE4: dout  = 8'b00111000; // 2788 :  56 - 0x38
      12'hAE5: dout  = 8'b00000000; // 2789 :   0 - 0x0
      12'hAE6: dout  = 8'b00000000; // 2790 :   0 - 0x0
      12'hAE7: dout  = 8'b00000000; // 2791 :   0 - 0x0
      12'hAE8: dout  = 8'b00100000; // 2792 :  32 - 0x20 -- Background 0x5d
      12'hAE9: dout  = 8'b11100111; // 2793 : 231 - 0xe7
      12'hAEA: dout  = 8'b11100111; // 2794 : 231 - 0xe7
      12'hAEB: dout  = 8'b11100111; // 2795 : 231 - 0xe7
      12'hAEC: dout  = 8'b11100111; // 2796 : 231 - 0xe7
      12'hAED: dout  = 8'b11100111; // 2797 : 231 - 0xe7
      12'hAEE: dout  = 8'b11101111; // 2798 : 239 - 0xef
      12'hAEF: dout  = 8'b00000000; // 2799 :   0 - 0x0
      12'hAF0: dout  = 8'b00000010; // 2800 :   2 - 0x2 -- Background 0x5e
      12'hAF1: dout  = 8'b01111110; // 2801 : 126 - 0x7e
      12'hAF2: dout  = 8'b01111110; // 2802 : 126 - 0x7e
      12'hAF3: dout  = 8'b01111110; // 2803 : 126 - 0x7e
      12'hAF4: dout  = 8'b01111110; // 2804 : 126 - 0x7e
      12'hAF5: dout  = 8'b01111110; // 2805 : 126 - 0x7e
      12'hAF6: dout  = 8'b11111110; // 2806 : 254 - 0xfe
      12'hAF7: dout  = 8'b00000000; // 2807 :   0 - 0x0
      12'hAF8: dout  = 8'b01111111; // 2808 : 127 - 0x7f -- Background 0x5f
      12'hAF9: dout  = 8'b01111111; // 2809 : 127 - 0x7f
      12'hAFA: dout  = 8'b01111111; // 2810 : 127 - 0x7f
      12'hAFB: dout  = 8'b01100111; // 2811 : 103 - 0x67
      12'hAFC: dout  = 8'b01100111; // 2812 : 103 - 0x67
      12'hAFD: dout  = 8'b01111111; // 2813 : 127 - 0x7f
      12'hAFE: dout  = 8'b01111111; // 2814 : 127 - 0x7f
      12'hAFF: dout  = 8'b01111111; // 2815 : 127 - 0x7f
      12'hB00: dout  = 8'b11111111; // 2816 : 255 - 0xff -- Background 0x60
      12'hB01: dout  = 8'b10000000; // 2817 : 128 - 0x80
      12'hB02: dout  = 8'b11111100; // 2818 : 252 - 0xfc
      12'hB03: dout  = 8'b10001100; // 2819 : 140 - 0x8c
      12'hB04: dout  = 8'b10001100; // 2820 : 140 - 0x8c
      12'hB05: dout  = 8'b10001100; // 2821 : 140 - 0x8c
      12'hB06: dout  = 8'b10001100; // 2822 : 140 - 0x8c
      12'hB07: dout  = 8'b10001100; // 2823 : 140 - 0x8c
      12'hB08: dout  = 8'b11111111; // 2824 : 255 - 0xff -- Background 0x61
      12'hB09: dout  = 8'b00000000; // 2825 :   0 - 0x0
      12'hB0A: dout  = 8'b00001111; // 2826 :  15 - 0xf
      12'hB0B: dout  = 8'b00001001; // 2827 :   9 - 0x9
      12'hB0C: dout  = 8'b00001001; // 2828 :   9 - 0x9
      12'hB0D: dout  = 8'b00001001; // 2829 :   9 - 0x9
      12'hB0E: dout  = 8'b00001001; // 2830 :   9 - 0x9
      12'hB0F: dout  = 8'b00001001; // 2831 :   9 - 0x9
      12'hB10: dout  = 8'b11111111; // 2832 : 255 - 0xff -- Background 0x62
      12'hB11: dout  = 8'b00000000; // 2833 :   0 - 0x0
      12'hB12: dout  = 8'b11111111; // 2834 : 255 - 0xff
      12'hB13: dout  = 8'b11111111; // 2835 : 255 - 0xff
      12'hB14: dout  = 8'b11111111; // 2836 : 255 - 0xff
      12'hB15: dout  = 8'b11111111; // 2837 : 255 - 0xff
      12'hB16: dout  = 8'b11111111; // 2838 : 255 - 0xff
      12'hB17: dout  = 8'b11111111; // 2839 : 255 - 0xff
      12'hB18: dout  = 8'b11111111; // 2840 : 255 - 0xff -- Background 0x63
      12'hB19: dout  = 8'b00000001; // 2841 :   1 - 0x1
      12'hB1A: dout  = 8'b11111111; // 2842 : 255 - 0xff
      12'hB1B: dout  = 8'b10101001; // 2843 : 169 - 0xa9
      12'hB1C: dout  = 8'b11010001; // 2844 : 209 - 0xd1
      12'hB1D: dout  = 8'b10101001; // 2845 : 169 - 0xa9
      12'hB1E: dout  = 8'b11010001; // 2846 : 209 - 0xd1
      12'hB1F: dout  = 8'b10101001; // 2847 : 169 - 0xa9
      12'hB20: dout  = 8'b10001100; // 2848 : 140 - 0x8c -- Background 0x64
      12'hB21: dout  = 8'b10001100; // 2849 : 140 - 0x8c
      12'hB22: dout  = 8'b10001100; // 2850 : 140 - 0x8c
      12'hB23: dout  = 8'b10001100; // 2851 : 140 - 0x8c
      12'hB24: dout  = 8'b10001100; // 2852 : 140 - 0x8c
      12'hB25: dout  = 8'b10001100; // 2853 : 140 - 0x8c
      12'hB26: dout  = 8'b11111111; // 2854 : 255 - 0xff
      12'hB27: dout  = 8'b00111111; // 2855 :  63 - 0x3f
      12'hB28: dout  = 8'b00001001; // 2856 :   9 - 0x9 -- Background 0x65
      12'hB29: dout  = 8'b00001001; // 2857 :   9 - 0x9
      12'hB2A: dout  = 8'b00001001; // 2858 :   9 - 0x9
      12'hB2B: dout  = 8'b00001001; // 2859 :   9 - 0x9
      12'hB2C: dout  = 8'b00001001; // 2860 :   9 - 0x9
      12'hB2D: dout  = 8'b00001001; // 2861 :   9 - 0x9
      12'hB2E: dout  = 8'b11111111; // 2862 : 255 - 0xff
      12'hB2F: dout  = 8'b11111111; // 2863 : 255 - 0xff
      12'hB30: dout  = 8'b11111111; // 2864 : 255 - 0xff -- Background 0x66
      12'hB31: dout  = 8'b11111111; // 2865 : 255 - 0xff
      12'hB32: dout  = 8'b11111111; // 2866 : 255 - 0xff
      12'hB33: dout  = 8'b11111111; // 2867 : 255 - 0xff
      12'hB34: dout  = 8'b11111111; // 2868 : 255 - 0xff
      12'hB35: dout  = 8'b11111111; // 2869 : 255 - 0xff
      12'hB36: dout  = 8'b11111111; // 2870 : 255 - 0xff
      12'hB37: dout  = 8'b11111111; // 2871 : 255 - 0xff
      12'hB38: dout  = 8'b11010001; // 2872 : 209 - 0xd1 -- Background 0x67
      12'hB39: dout  = 8'b10101001; // 2873 : 169 - 0xa9
      12'hB3A: dout  = 8'b11010001; // 2874 : 209 - 0xd1
      12'hB3B: dout  = 8'b10101001; // 2875 : 169 - 0xa9
      12'hB3C: dout  = 8'b11010001; // 2876 : 209 - 0xd1
      12'hB3D: dout  = 8'b10101001; // 2877 : 169 - 0xa9
      12'hB3E: dout  = 8'b11111111; // 2878 : 255 - 0xff
      12'hB3F: dout  = 8'b11111100; // 2879 : 252 - 0xfc
      12'hB40: dout  = 8'b00100011; // 2880 :  35 - 0x23 -- Background 0x68
      12'hB41: dout  = 8'b00100011; // 2881 :  35 - 0x23
      12'hB42: dout  = 8'b00100011; // 2882 :  35 - 0x23
      12'hB43: dout  = 8'b00100011; // 2883 :  35 - 0x23
      12'hB44: dout  = 8'b00100011; // 2884 :  35 - 0x23
      12'hB45: dout  = 8'b00100011; // 2885 :  35 - 0x23
      12'hB46: dout  = 8'b00100011; // 2886 :  35 - 0x23
      12'hB47: dout  = 8'b00100011; // 2887 :  35 - 0x23
      12'hB48: dout  = 8'b00000100; // 2888 :   4 - 0x4 -- Background 0x69
      12'hB49: dout  = 8'b00000100; // 2889 :   4 - 0x4
      12'hB4A: dout  = 8'b00000100; // 2890 :   4 - 0x4
      12'hB4B: dout  = 8'b00000100; // 2891 :   4 - 0x4
      12'hB4C: dout  = 8'b00000100; // 2892 :   4 - 0x4
      12'hB4D: dout  = 8'b00000100; // 2893 :   4 - 0x4
      12'hB4E: dout  = 8'b00000100; // 2894 :   4 - 0x4
      12'hB4F: dout  = 8'b00000100; // 2895 :   4 - 0x4
      12'hB50: dout  = 8'b01000100; // 2896 :  68 - 0x44 -- Background 0x6a
      12'hB51: dout  = 8'b10100100; // 2897 : 164 - 0xa4
      12'hB52: dout  = 8'b01000100; // 2898 :  68 - 0x44
      12'hB53: dout  = 8'b10100100; // 2899 : 164 - 0xa4
      12'hB54: dout  = 8'b01000100; // 2900 :  68 - 0x44
      12'hB55: dout  = 8'b10100100; // 2901 : 164 - 0xa4
      12'hB56: dout  = 8'b01000100; // 2902 :  68 - 0x44
      12'hB57: dout  = 8'b10100100; // 2903 : 164 - 0xa4
      12'hB58: dout  = 8'b00011111; // 2904 :  31 - 0x1f -- Background 0x6b
      12'hB59: dout  = 8'b00111111; // 2905 :  63 - 0x3f
      12'hB5A: dout  = 8'b01111111; // 2906 : 127 - 0x7f
      12'hB5B: dout  = 8'b01111111; // 2907 : 127 - 0x7f
      12'hB5C: dout  = 8'b11111111; // 2908 : 255 - 0xff
      12'hB5D: dout  = 8'b11111111; // 2909 : 255 - 0xff
      12'hB5E: dout  = 8'b11111111; // 2910 : 255 - 0xff
      12'hB5F: dout  = 8'b11111110; // 2911 : 254 - 0xfe
      12'hB60: dout  = 8'b11111111; // 2912 : 255 - 0xff -- Background 0x6c
      12'hB61: dout  = 8'b01111111; // 2913 : 127 - 0x7f
      12'hB62: dout  = 8'b01111111; // 2914 : 127 - 0x7f
      12'hB63: dout  = 8'b00111111; // 2915 :  63 - 0x3f
      12'hB64: dout  = 8'b00000000; // 2916 :   0 - 0x0
      12'hB65: dout  = 8'b00000000; // 2917 :   0 - 0x0
      12'hB66: dout  = 8'b00000001; // 2918 :   1 - 0x1
      12'hB67: dout  = 8'b00000001; // 2919 :   1 - 0x1
      12'hB68: dout  = 8'b11111111; // 2920 : 255 - 0xff -- Background 0x6d
      12'hB69: dout  = 8'b10000000; // 2921 : 128 - 0x80
      12'hB6A: dout  = 8'b10000000; // 2922 : 128 - 0x80
      12'hB6B: dout  = 8'b00000000; // 2923 :   0 - 0x0
      12'hB6C: dout  = 8'b00000000; // 2924 :   0 - 0x0
      12'hB6D: dout  = 8'b11111000; // 2925 : 248 - 0xf8
      12'hB6E: dout  = 8'b11111100; // 2926 : 252 - 0xfc
      12'hB6F: dout  = 8'b11111100; // 2927 : 252 - 0xfc
      12'hB70: dout  = 8'b11111111; // 2928 : 255 - 0xff -- Background 0x6e
      12'hB71: dout  = 8'b11111111; // 2929 : 255 - 0xff
      12'hB72: dout  = 8'b11111111; // 2930 : 255 - 0xff
      12'hB73: dout  = 8'b11111111; // 2931 : 255 - 0xff
      12'hB74: dout  = 8'b11111111; // 2932 : 255 - 0xff
      12'hB75: dout  = 8'b01111110; // 2933 : 126 - 0x7e
      12'hB76: dout  = 8'b00111100; // 2934 :  60 - 0x3c
      12'hB77: dout  = 8'b00000000; // 2935 :   0 - 0x0
      12'hB78: dout  = 8'b11111000; // 2936 : 248 - 0xf8 -- Background 0x6f
      12'hB79: dout  = 8'b00000100; // 2937 :   4 - 0x4
      12'hB7A: dout  = 8'b00000010; // 2938 :   2 - 0x2
      12'hB7B: dout  = 8'b00000010; // 2939 :   2 - 0x2
      12'hB7C: dout  = 8'b00011101; // 2940 :  29 - 0x1d
      12'hB7D: dout  = 8'b00111111; // 2941 :  63 - 0x3f
      12'hB7E: dout  = 8'b01111111; // 2942 : 127 - 0x7f
      12'hB7F: dout  = 8'b01111111; // 2943 : 127 - 0x7f
      12'hB80: dout  = 8'b11111100; // 2944 : 252 - 0xfc -- Background 0x70
      12'hB81: dout  = 8'b10000000; // 2945 : 128 - 0x80
      12'hB82: dout  = 8'b10000000; // 2946 : 128 - 0x80
      12'hB83: dout  = 8'b10000000; // 2947 : 128 - 0x80
      12'hB84: dout  = 8'b10000000; // 2948 : 128 - 0x80
      12'hB85: dout  = 8'b10000000; // 2949 : 128 - 0x80
      12'hB86: dout  = 8'b01100000; // 2950 :  96 - 0x60
      12'hB87: dout  = 8'b00011111; // 2951 :  31 - 0x1f
      12'hB88: dout  = 8'b00000011; // 2952 :   3 - 0x3 -- Background 0x71
      12'hB89: dout  = 8'b00000011; // 2953 :   3 - 0x3
      12'hB8A: dout  = 8'b00000011; // 2954 :   3 - 0x3
      12'hB8B: dout  = 8'b00000011; // 2955 :   3 - 0x3
      12'hB8C: dout  = 8'b00000001; // 2956 :   1 - 0x1
      12'hB8D: dout  = 8'b00000001; // 2957 :   1 - 0x1
      12'hB8E: dout  = 8'b00000000; // 2958 :   0 - 0x0
      12'hB8F: dout  = 8'b11111111; // 2959 : 255 - 0xff
      12'hB90: dout  = 8'b11111110; // 2960 : 254 - 0xfe -- Background 0x72
      12'hB91: dout  = 8'b11111110; // 2961 : 254 - 0xfe
      12'hB92: dout  = 8'b11111110; // 2962 : 254 - 0xfe
      12'hB93: dout  = 8'b11111110; // 2963 : 254 - 0xfe
      12'hB94: dout  = 8'b11111100; // 2964 : 252 - 0xfc
      12'hB95: dout  = 8'b11111100; // 2965 : 252 - 0xfc
      12'hB96: dout  = 8'b11111000; // 2966 : 248 - 0xf8
      12'hB97: dout  = 8'b11111111; // 2967 : 255 - 0xff
      12'hB98: dout  = 8'b00000000; // 2968 :   0 - 0x0 -- Background 0x73
      12'hB99: dout  = 8'b00000000; // 2969 :   0 - 0x0
      12'hB9A: dout  = 8'b00000000; // 2970 :   0 - 0x0
      12'hB9B: dout  = 8'b00000000; // 2971 :   0 - 0x0
      12'hB9C: dout  = 8'b00000000; // 2972 :   0 - 0x0
      12'hB9D: dout  = 8'b00000000; // 2973 :   0 - 0x0
      12'hB9E: dout  = 8'b00000000; // 2974 :   0 - 0x0
      12'hB9F: dout  = 8'b11111111; // 2975 : 255 - 0xff
      12'hBA0: dout  = 8'b01111111; // 2976 : 127 - 0x7f -- Background 0x74
      12'hBA1: dout  = 8'b00111111; // 2977 :  63 - 0x3f
      12'hBA2: dout  = 8'b00011101; // 2978 :  29 - 0x1d
      12'hBA3: dout  = 8'b00000001; // 2979 :   1 - 0x1
      12'hBA4: dout  = 8'b00000001; // 2980 :   1 - 0x1
      12'hBA5: dout  = 8'b00000001; // 2981 :   1 - 0x1
      12'hBA6: dout  = 8'b00000011; // 2982 :   3 - 0x3
      12'hBA7: dout  = 8'b11111110; // 2983 : 254 - 0xfe
      12'hBA8: dout  = 8'b10000000; // 2984 : 128 - 0x80 -- Background 0x75
      12'hBA9: dout  = 8'b10000000; // 2985 : 128 - 0x80
      12'hBAA: dout  = 8'b10000000; // 2986 : 128 - 0x80
      12'hBAB: dout  = 8'b10000000; // 2987 : 128 - 0x80
      12'hBAC: dout  = 8'b10000000; // 2988 : 128 - 0x80
      12'hBAD: dout  = 8'b10000100; // 2989 : 132 - 0x84
      12'hBAE: dout  = 8'b11001010; // 2990 : 202 - 0xca
      12'hBAF: dout  = 8'b10110001; // 2991 : 177 - 0xb1
      12'hBB0: dout  = 8'b00000001; // 2992 :   1 - 0x1 -- Background 0x76
      12'hBB1: dout  = 8'b00000001; // 2993 :   1 - 0x1
      12'hBB2: dout  = 8'b00000001; // 2994 :   1 - 0x1
      12'hBB3: dout  = 8'b00000001; // 2995 :   1 - 0x1
      12'hBB4: dout  = 8'b00000001; // 2996 :   1 - 0x1
      12'hBB5: dout  = 8'b00100001; // 2997 :  33 - 0x21
      12'hBB6: dout  = 8'b01010011; // 2998 :  83 - 0x53
      12'hBB7: dout  = 8'b10001101; // 2999 : 141 - 0x8d
      12'hBB8: dout  = 8'b00000000; // 3000 :   0 - 0x0 -- Background 0x77
      12'hBB9: dout  = 8'b00000000; // 3001 :   0 - 0x0
      12'hBBA: dout  = 8'b00000000; // 3002 :   0 - 0x0
      12'hBBB: dout  = 8'b00000000; // 3003 :   0 - 0x0
      12'hBBC: dout  = 8'b01110111; // 3004 : 119 - 0x77
      12'hBBD: dout  = 8'b11111111; // 3005 : 255 - 0xff
      12'hBBE: dout  = 8'b11111111; // 3006 : 255 - 0xff
      12'hBBF: dout  = 8'b11111111; // 3007 : 255 - 0xff
      12'hBC0: dout  = 8'b11111111; // 3008 : 255 - 0xff -- Background 0x78
      12'hBC1: dout  = 8'b11111111; // 3009 : 255 - 0xff
      12'hBC2: dout  = 8'b11111111; // 3010 : 255 - 0xff
      12'hBC3: dout  = 8'b11111111; // 3011 : 255 - 0xff
      12'hBC4: dout  = 8'b11111111; // 3012 : 255 - 0xff
      12'hBC5: dout  = 8'b11111111; // 3013 : 255 - 0xff
      12'hBC6: dout  = 8'b11111111; // 3014 : 255 - 0xff
      12'hBC7: dout  = 8'b11111111; // 3015 : 255 - 0xff
      12'hBC8: dout  = 8'b11111111; // 3016 : 255 - 0xff -- Background 0x79
      12'hBC9: dout  = 8'b11111111; // 3017 : 255 - 0xff
      12'hBCA: dout  = 8'b11111111; // 3018 : 255 - 0xff
      12'hBCB: dout  = 8'b01110111; // 3019 : 119 - 0x77
      12'hBCC: dout  = 8'b01110111; // 3020 : 119 - 0x77
      12'hBCD: dout  = 8'b01110111; // 3021 : 119 - 0x77
      12'hBCE: dout  = 8'b01110111; // 3022 : 119 - 0x77
      12'hBCF: dout  = 8'b01110111; // 3023 : 119 - 0x77
      12'hBD0: dout  = 8'b11111111; // 3024 : 255 - 0xff -- Background 0x7a
      12'hBD1: dout  = 8'b11111111; // 3025 : 255 - 0xff
      12'hBD2: dout  = 8'b11111111; // 3026 : 255 - 0xff
      12'hBD3: dout  = 8'b11100111; // 3027 : 231 - 0xe7
      12'hBD4: dout  = 8'b11100111; // 3028 : 231 - 0xe7
      12'hBD5: dout  = 8'b11111111; // 3029 : 255 - 0xff
      12'hBD6: dout  = 8'b11111111; // 3030 : 255 - 0xff
      12'hBD7: dout  = 8'b11111110; // 3031 : 254 - 0xfe
      12'hBD8: dout  = 8'b00000000; // 3032 :   0 - 0x0 -- Background 0x7b
      12'hBD9: dout  = 8'b00100001; // 3033 :  33 - 0x21
      12'hBDA: dout  = 8'b00100001; // 3034 :  33 - 0x21
      12'hBDB: dout  = 8'b01000001; // 3035 :  65 - 0x41
      12'hBDC: dout  = 8'b01000001; // 3036 :  65 - 0x41
      12'hBDD: dout  = 8'b01000001; // 3037 :  65 - 0x41
      12'hBDE: dout  = 8'b01000001; // 3038 :  65 - 0x41
      12'hBDF: dout  = 8'b01000001; // 3039 :  65 - 0x41
      12'hBE0: dout  = 8'b00000000; // 3040 :   0 - 0x0 -- Background 0x7c
      12'hBE1: dout  = 8'b10000000; // 3041 : 128 - 0x80
      12'hBE2: dout  = 8'b10000000; // 3042 : 128 - 0x80
      12'hBE3: dout  = 8'b10000000; // 3043 : 128 - 0x80
      12'hBE4: dout  = 8'b10000000; // 3044 : 128 - 0x80
      12'hBE5: dout  = 8'b10000000; // 3045 : 128 - 0x80
      12'hBE6: dout  = 8'b10000000; // 3046 : 128 - 0x80
      12'hBE7: dout  = 8'b10000000; // 3047 : 128 - 0x80
      12'hBE8: dout  = 8'b00100001; // 3048 :  33 - 0x21 -- Background 0x7d
      12'hBE9: dout  = 8'b00100001; // 3049 :  33 - 0x21
      12'hBEA: dout  = 8'b00000001; // 3050 :   1 - 0x1
      12'hBEB: dout  = 8'b00000001; // 3051 :   1 - 0x1
      12'hBEC: dout  = 8'b00000001; // 3052 :   1 - 0x1
      12'hBED: dout  = 8'b00000001; // 3053 :   1 - 0x1
      12'hBEE: dout  = 8'b00000001; // 3054 :   1 - 0x1
      12'hBEF: dout  = 8'b00000001; // 3055 :   1 - 0x1
      12'hBF0: dout  = 8'b10000000; // 3056 : 128 - 0x80 -- Background 0x7e
      12'hBF1: dout  = 8'b10000000; // 3057 : 128 - 0x80
      12'hBF2: dout  = 8'b10000000; // 3058 : 128 - 0x80
      12'hBF3: dout  = 8'b10000000; // 3059 : 128 - 0x80
      12'hBF4: dout  = 8'b10000000; // 3060 : 128 - 0x80
      12'hBF5: dout  = 8'b10000000; // 3061 : 128 - 0x80
      12'hBF6: dout  = 8'b10000000; // 3062 : 128 - 0x80
      12'hBF7: dout  = 8'b10000000; // 3063 : 128 - 0x80
      12'hBF8: dout  = 8'b00000001; // 3064 :   1 - 0x1 -- Background 0x7f
      12'hBF9: dout  = 8'b00000001; // 3065 :   1 - 0x1
      12'hBFA: dout  = 8'b00000110; // 3066 :   6 - 0x6
      12'hBFB: dout  = 8'b00001000; // 3067 :   8 - 0x8
      12'hBFC: dout  = 8'b00011000; // 3068 :  24 - 0x18
      12'hBFD: dout  = 8'b00100000; // 3069 :  32 - 0x20
      12'hBFE: dout  = 8'b00100000; // 3070 :  32 - 0x20
      12'hBFF: dout  = 8'b11000000; // 3071 : 192 - 0xc0
      12'hC00: dout  = 8'b00000100; // 3072 :   4 - 0x4 -- Background 0x80
      12'hC01: dout  = 8'b00000100; // 3073 :   4 - 0x4
      12'hC02: dout  = 8'b11000100; // 3074 : 196 - 0xc4
      12'hC03: dout  = 8'b11110100; // 3075 : 244 - 0xf4
      12'hC04: dout  = 8'b11110100; // 3076 : 244 - 0xf4
      12'hC05: dout  = 8'b00000100; // 3077 :   4 - 0x4
      12'hC06: dout  = 8'b00000100; // 3078 :   4 - 0x4
      12'hC07: dout  = 8'b00000101; // 3079 :   5 - 0x5
      12'hC08: dout  = 8'b01110000; // 3080 : 112 - 0x70 -- Background 0x81
      12'hC09: dout  = 8'b11110000; // 3081 : 240 - 0xf0
      12'hC0A: dout  = 8'b11110000; // 3082 : 240 - 0xf0
      12'hC0B: dout  = 8'b11111111; // 3083 : 255 - 0xff
      12'hC0C: dout  = 8'b11111111; // 3084 : 255 - 0xff
      12'hC0D: dout  = 8'b11110000; // 3085 : 240 - 0xf0
      12'hC0E: dout  = 8'b11110000; // 3086 : 240 - 0xf0
      12'hC0F: dout  = 8'b01110000; // 3087 : 112 - 0x70
      12'hC10: dout  = 8'b11000000; // 3088 : 192 - 0xc0 -- Background 0x82
      12'hC11: dout  = 8'b10000111; // 3089 : 135 - 0x87
      12'hC12: dout  = 8'b00011000; // 3090 :  24 - 0x18
      12'hC13: dout  = 8'b10110000; // 3091 : 176 - 0xb0
      12'hC14: dout  = 8'b11100111; // 3092 : 231 - 0xe7
      12'hC15: dout  = 8'b11100111; // 3093 : 231 - 0xe7
      12'hC16: dout  = 8'b11101111; // 3094 : 239 - 0xef
      12'hC17: dout  = 8'b11101111; // 3095 : 239 - 0xef
      12'hC18: dout  = 8'b01101111; // 3096 : 111 - 0x6f -- Background 0x83
      12'hC19: dout  = 8'b01000011; // 3097 :  67 - 0x43
      12'hC1A: dout  = 8'b01011101; // 3098 :  93 - 0x5d
      12'hC1B: dout  = 8'b00111111; // 3099 :  63 - 0x3f
      12'hC1C: dout  = 8'b00111111; // 3100 :  63 - 0x3f
      12'hC1D: dout  = 8'b01111111; // 3101 : 127 - 0x7f
      12'hC1E: dout  = 8'b01111111; // 3102 : 127 - 0x7f
      12'hC1F: dout  = 8'b11111111; // 3103 : 255 - 0xff
      12'hC20: dout  = 8'b00000011; // 3104 :   3 - 0x3 -- Background 0x84
      12'hC21: dout  = 8'b11111111; // 3105 : 255 - 0xff
      12'hC22: dout  = 8'b11110001; // 3106 : 241 - 0xf1
      12'hC23: dout  = 8'b01101110; // 3107 : 110 - 0x6e
      12'hC24: dout  = 8'b11001111; // 3108 : 207 - 0xcf
      12'hC25: dout  = 8'b11011111; // 3109 : 223 - 0xdf
      12'hC26: dout  = 8'b11111111; // 3110 : 255 - 0xff
      12'hC27: dout  = 8'b11111111; // 3111 : 255 - 0xff
      12'hC28: dout  = 8'b11111101; // 3112 : 253 - 0xfd -- Background 0x85
      12'hC29: dout  = 8'b11111011; // 3113 : 251 - 0xfb
      12'hC2A: dout  = 8'b11111011; // 3114 : 251 - 0xfb
      12'hC2B: dout  = 8'b11110111; // 3115 : 247 - 0xf7
      12'hC2C: dout  = 8'b11110111; // 3116 : 247 - 0xf7
      12'hC2D: dout  = 8'b00001111; // 3117 :  15 - 0xf
      12'hC2E: dout  = 8'b01111111; // 3118 : 127 - 0x7f
      12'hC2F: dout  = 8'b11111111; // 3119 : 255 - 0xff
      12'hC30: dout  = 8'b11111111; // 3120 : 255 - 0xff -- Background 0x86
      12'hC31: dout  = 8'b10000000; // 3121 : 128 - 0x80
      12'hC32: dout  = 8'b10000000; // 3122 : 128 - 0x80
      12'hC33: dout  = 8'b10000000; // 3123 : 128 - 0x80
      12'hC34: dout  = 8'b10000000; // 3124 : 128 - 0x80
      12'hC35: dout  = 8'b11111111; // 3125 : 255 - 0xff
      12'hC36: dout  = 8'b11111111; // 3126 : 255 - 0xff
      12'hC37: dout  = 8'b10000000; // 3127 : 128 - 0x80
      12'hC38: dout  = 8'b11111110; // 3128 : 254 - 0xfe -- Background 0x87
      12'hC39: dout  = 8'b00000011; // 3129 :   3 - 0x3
      12'hC3A: dout  = 8'b00000011; // 3130 :   3 - 0x3
      12'hC3B: dout  = 8'b00000011; // 3131 :   3 - 0x3
      12'hC3C: dout  = 8'b00000011; // 3132 :   3 - 0x3
      12'hC3D: dout  = 8'b11111111; // 3133 : 255 - 0xff
      12'hC3E: dout  = 8'b11111111; // 3134 : 255 - 0xff
      12'hC3F: dout  = 8'b00000011; // 3135 :   3 - 0x3
      12'hC40: dout  = 8'b00000000; // 3136 :   0 - 0x0 -- Background 0x88
      12'hC41: dout  = 8'b11111111; // 3137 : 255 - 0xff
      12'hC42: dout  = 8'b00000000; // 3138 :   0 - 0x0
      12'hC43: dout  = 8'b00000000; // 3139 :   0 - 0x0
      12'hC44: dout  = 8'b00000000; // 3140 :   0 - 0x0
      12'hC45: dout  = 8'b00000000; // 3141 :   0 - 0x0
      12'hC46: dout  = 8'b11111111; // 3142 : 255 - 0xff
      12'hC47: dout  = 8'b11111111; // 3143 : 255 - 0xff
      12'hC48: dout  = 8'b00100011; // 3144 :  35 - 0x23 -- Background 0x89
      12'hC49: dout  = 8'b11110011; // 3145 : 243 - 0xf3
      12'hC4A: dout  = 8'b00001011; // 3146 :  11 - 0xb
      12'hC4B: dout  = 8'b00001011; // 3147 :  11 - 0xb
      12'hC4C: dout  = 8'b00001011; // 3148 :  11 - 0xb
      12'hC4D: dout  = 8'b00000111; // 3149 :   7 - 0x7
      12'hC4E: dout  = 8'b11111111; // 3150 : 255 - 0xff
      12'hC4F: dout  = 8'b11111111; // 3151 : 255 - 0xff
      12'hC50: dout  = 8'b10000000; // 3152 : 128 - 0x80 -- Background 0x8a
      12'hC51: dout  = 8'b10000000; // 3153 : 128 - 0x80
      12'hC52: dout  = 8'b10000000; // 3154 : 128 - 0x80
      12'hC53: dout  = 8'b10000000; // 3155 : 128 - 0x80
      12'hC54: dout  = 8'b11111111; // 3156 : 255 - 0xff
      12'hC55: dout  = 8'b10000000; // 3157 : 128 - 0x80
      12'hC56: dout  = 8'b10000000; // 3158 : 128 - 0x80
      12'hC57: dout  = 8'b10000000; // 3159 : 128 - 0x80
      12'hC58: dout  = 8'b00000011; // 3160 :   3 - 0x3 -- Background 0x8b
      12'hC59: dout  = 8'b00000011; // 3161 :   3 - 0x3
      12'hC5A: dout  = 8'b00000011; // 3162 :   3 - 0x3
      12'hC5B: dout  = 8'b00000011; // 3163 :   3 - 0x3
      12'hC5C: dout  = 8'b11111111; // 3164 : 255 - 0xff
      12'hC5D: dout  = 8'b00000011; // 3165 :   3 - 0x3
      12'hC5E: dout  = 8'b00000011; // 3166 :   3 - 0x3
      12'hC5F: dout  = 8'b00000011; // 3167 :   3 - 0x3
      12'hC60: dout  = 8'b00000000; // 3168 :   0 - 0x0 -- Background 0x8c
      12'hC61: dout  = 8'b00000000; // 3169 :   0 - 0x0
      12'hC62: dout  = 8'b00000000; // 3170 :   0 - 0x0
      12'hC63: dout  = 8'b00000000; // 3171 :   0 - 0x0
      12'hC64: dout  = 8'b00000000; // 3172 :   0 - 0x0
      12'hC65: dout  = 8'b11111111; // 3173 : 255 - 0xff
      12'hC66: dout  = 8'b00000000; // 3174 :   0 - 0x0
      12'hC67: dout  = 8'b00000000; // 3175 :   0 - 0x0
      12'hC68: dout  = 8'b00000111; // 3176 :   7 - 0x7 -- Background 0x8d
      12'hC69: dout  = 8'b00000111; // 3177 :   7 - 0x7
      12'hC6A: dout  = 8'b00000011; // 3178 :   3 - 0x3
      12'hC6B: dout  = 8'b00000011; // 3179 :   3 - 0x3
      12'hC6C: dout  = 8'b00000011; // 3180 :   3 - 0x3
      12'hC6D: dout  = 8'b11111111; // 3181 : 255 - 0xff
      12'hC6E: dout  = 8'b00000011; // 3182 :   3 - 0x3
      12'hC6F: dout  = 8'b00000011; // 3183 :   3 - 0x3
      12'hC70: dout  = 8'b10000000; // 3184 : 128 - 0x80 -- Background 0x8e
      12'hC71: dout  = 8'b11111111; // 3185 : 255 - 0xff
      12'hC72: dout  = 8'b11111111; // 3186 : 255 - 0xff
      12'hC73: dout  = 8'b11111111; // 3187 : 255 - 0xff
      12'hC74: dout  = 8'b11111111; // 3188 : 255 - 0xff
      12'hC75: dout  = 8'b11111111; // 3189 : 255 - 0xff
      12'hC76: dout  = 8'b11111111; // 3190 : 255 - 0xff
      12'hC77: dout  = 8'b11111111; // 3191 : 255 - 0xff
      12'hC78: dout  = 8'b00000011; // 3192 :   3 - 0x3 -- Background 0x8f
      12'hC79: dout  = 8'b11111111; // 3193 : 255 - 0xff
      12'hC7A: dout  = 8'b11111111; // 3194 : 255 - 0xff
      12'hC7B: dout  = 8'b11111111; // 3195 : 255 - 0xff
      12'hC7C: dout  = 8'b11111111; // 3196 : 255 - 0xff
      12'hC7D: dout  = 8'b11111111; // 3197 : 255 - 0xff
      12'hC7E: dout  = 8'b11111111; // 3198 : 255 - 0xff
      12'hC7F: dout  = 8'b11111111; // 3199 : 255 - 0xff
      12'hC80: dout  = 8'b11111111; // 3200 : 255 - 0xff -- Background 0x90
      12'hC81: dout  = 8'b11111111; // 3201 : 255 - 0xff
      12'hC82: dout  = 8'b11111111; // 3202 : 255 - 0xff
      12'hC83: dout  = 8'b11111111; // 3203 : 255 - 0xff
      12'hC84: dout  = 8'b11111111; // 3204 : 255 - 0xff
      12'hC85: dout  = 8'b11111111; // 3205 : 255 - 0xff
      12'hC86: dout  = 8'b11111111; // 3206 : 255 - 0xff
      12'hC87: dout  = 8'b11111111; // 3207 : 255 - 0xff
      12'hC88: dout  = 8'b11111111; // 3208 : 255 - 0xff -- Background 0x91
      12'hC89: dout  = 8'b11111111; // 3209 : 255 - 0xff
      12'hC8A: dout  = 8'b11010101; // 3210 : 213 - 0xd5
      12'hC8B: dout  = 8'b10101010; // 3211 : 170 - 0xaa
      12'hC8C: dout  = 8'b11010101; // 3212 : 213 - 0xd5
      12'hC8D: dout  = 8'b10000000; // 3213 : 128 - 0x80
      12'hC8E: dout  = 8'b10000000; // 3214 : 128 - 0x80
      12'hC8F: dout  = 8'b11111111; // 3215 : 255 - 0xff
      12'hC90: dout  = 8'b11111111; // 3216 : 255 - 0xff -- Background 0x92
      12'hC91: dout  = 8'b11111111; // 3217 : 255 - 0xff
      12'hC92: dout  = 8'b01010111; // 3218 :  87 - 0x57
      12'hC93: dout  = 8'b10101011; // 3219 : 171 - 0xab
      12'hC94: dout  = 8'b01010111; // 3220 :  87 - 0x57
      12'hC95: dout  = 8'b00000011; // 3221 :   3 - 0x3
      12'hC96: dout  = 8'b00000011; // 3222 :   3 - 0x3
      12'hC97: dout  = 8'b11111110; // 3223 : 254 - 0xfe
      12'hC98: dout  = 8'b11111111; // 3224 : 255 - 0xff -- Background 0x93
      12'hC99: dout  = 8'b10101010; // 3225 : 170 - 0xaa
      12'hC9A: dout  = 8'b01010101; // 3226 :  85 - 0x55
      12'hC9B: dout  = 8'b10101010; // 3227 : 170 - 0xaa
      12'hC9C: dout  = 8'b00000000; // 3228 :   0 - 0x0
      12'hC9D: dout  = 8'b00000000; // 3229 :   0 - 0x0
      12'hC9E: dout  = 8'b11111111; // 3230 : 255 - 0xff
      12'hC9F: dout  = 8'b00000000; // 3231 :   0 - 0x0
      12'hCA0: dout  = 8'b11111111; // 3232 : 255 - 0xff -- Background 0x94
      12'hCA1: dout  = 8'b10101111; // 3233 : 175 - 0xaf
      12'hCA2: dout  = 8'b01010111; // 3234 :  87 - 0x57
      12'hCA3: dout  = 8'b10101011; // 3235 : 171 - 0xab
      12'hCA4: dout  = 8'b00001011; // 3236 :  11 - 0xb
      12'hCA5: dout  = 8'b00001011; // 3237 :  11 - 0xb
      12'hCA6: dout  = 8'b11110011; // 3238 : 243 - 0xf3
      12'hCA7: dout  = 8'b00100011; // 3239 :  35 - 0x23
      12'hCA8: dout  = 8'b11111111; // 3240 : 255 - 0xff -- Background 0x95
      12'hCA9: dout  = 8'b11111111; // 3241 : 255 - 0xff
      12'hCAA: dout  = 8'b11111111; // 3242 : 255 - 0xff
      12'hCAB: dout  = 8'b11111111; // 3243 : 255 - 0xff
      12'hCAC: dout  = 8'b11111111; // 3244 : 255 - 0xff
      12'hCAD: dout  = 8'b11111111; // 3245 : 255 - 0xff
      12'hCAE: dout  = 8'b11111111; // 3246 : 255 - 0xff
      12'hCAF: dout  = 8'b11111111; // 3247 : 255 - 0xff
      12'hCB0: dout  = 8'b11111111; // 3248 : 255 - 0xff -- Background 0x96
      12'hCB1: dout  = 8'b11111111; // 3249 : 255 - 0xff
      12'hCB2: dout  = 8'b11111111; // 3250 : 255 - 0xff
      12'hCB3: dout  = 8'b11111111; // 3251 : 255 - 0xff
      12'hCB4: dout  = 8'b11111111; // 3252 : 255 - 0xff
      12'hCB5: dout  = 8'b11111111; // 3253 : 255 - 0xff
      12'hCB6: dout  = 8'b11111111; // 3254 : 255 - 0xff
      12'hCB7: dout  = 8'b11111111; // 3255 : 255 - 0xff
      12'hCB8: dout  = 8'b11111111; // 3256 : 255 - 0xff -- Background 0x97
      12'hCB9: dout  = 8'b11111111; // 3257 : 255 - 0xff
      12'hCBA: dout  = 8'b11111111; // 3258 : 255 - 0xff
      12'hCBB: dout  = 8'b11111111; // 3259 : 255 - 0xff
      12'hCBC: dout  = 8'b11111111; // 3260 : 255 - 0xff
      12'hCBD: dout  = 8'b11111111; // 3261 : 255 - 0xff
      12'hCBE: dout  = 8'b11111111; // 3262 : 255 - 0xff
      12'hCBF: dout  = 8'b11111111; // 3263 : 255 - 0xff
      12'hCC0: dout  = 8'b11111111; // 3264 : 255 - 0xff -- Background 0x98
      12'hCC1: dout  = 8'b11111111; // 3265 : 255 - 0xff
      12'hCC2: dout  = 8'b11111111; // 3266 : 255 - 0xff
      12'hCC3: dout  = 8'b11111111; // 3267 : 255 - 0xff
      12'hCC4: dout  = 8'b11111111; // 3268 : 255 - 0xff
      12'hCC5: dout  = 8'b11111111; // 3269 : 255 - 0xff
      12'hCC6: dout  = 8'b11111111; // 3270 : 255 - 0xff
      12'hCC7: dout  = 8'b11111111; // 3271 : 255 - 0xff
      12'hCC8: dout  = 8'b00000000; // 3272 :   0 - 0x0 -- Background 0x99
      12'hCC9: dout  = 8'b00000000; // 3273 :   0 - 0x0
      12'hCCA: dout  = 8'b00000000; // 3274 :   0 - 0x0
      12'hCCB: dout  = 8'b00000000; // 3275 :   0 - 0x0
      12'hCCC: dout  = 8'b00000000; // 3276 :   0 - 0x0
      12'hCCD: dout  = 8'b00000000; // 3277 :   0 - 0x0
      12'hCCE: dout  = 8'b00000000; // 3278 :   0 - 0x0
      12'hCCF: dout  = 8'b00000000; // 3279 :   0 - 0x0
      12'hCD0: dout  = 8'b00000000; // 3280 :   0 - 0x0 -- Background 0x9a
      12'hCD1: dout  = 8'b00000000; // 3281 :   0 - 0x0
      12'hCD2: dout  = 8'b00000000; // 3282 :   0 - 0x0
      12'hCD3: dout  = 8'b00000000; // 3283 :   0 - 0x0
      12'hCD4: dout  = 8'b00000000; // 3284 :   0 - 0x0
      12'hCD5: dout  = 8'b00000000; // 3285 :   0 - 0x0
      12'hCD6: dout  = 8'b00000000; // 3286 :   0 - 0x0
      12'hCD7: dout  = 8'b00000000; // 3287 :   0 - 0x0
      12'hCD8: dout  = 8'b11111111; // 3288 : 255 - 0xff -- Background 0x9b
      12'hCD9: dout  = 8'b11111111; // 3289 : 255 - 0xff
      12'hCDA: dout  = 8'b11111111; // 3290 : 255 - 0xff
      12'hCDB: dout  = 8'b11111111; // 3291 : 255 - 0xff
      12'hCDC: dout  = 8'b11111111; // 3292 : 255 - 0xff
      12'hCDD: dout  = 8'b11111111; // 3293 : 255 - 0xff
      12'hCDE: dout  = 8'b11111111; // 3294 : 255 - 0xff
      12'hCDF: dout  = 8'b11111111; // 3295 : 255 - 0xff
      12'hCE0: dout  = 8'b11111111; // 3296 : 255 - 0xff -- Background 0x9c
      12'hCE1: dout  = 8'b11111111; // 3297 : 255 - 0xff
      12'hCE2: dout  = 8'b11111111; // 3298 : 255 - 0xff
      12'hCE3: dout  = 8'b11111111; // 3299 : 255 - 0xff
      12'hCE4: dout  = 8'b11111111; // 3300 : 255 - 0xff
      12'hCE5: dout  = 8'b11111111; // 3301 : 255 - 0xff
      12'hCE6: dout  = 8'b11111111; // 3302 : 255 - 0xff
      12'hCE7: dout  = 8'b11111111; // 3303 : 255 - 0xff
      12'hCE8: dout  = 8'b00000000; // 3304 :   0 - 0x0 -- Background 0x9d
      12'hCE9: dout  = 8'b11100000; // 3305 : 224 - 0xe0
      12'hCEA: dout  = 8'b11100000; // 3306 : 224 - 0xe0
      12'hCEB: dout  = 8'b11100000; // 3307 : 224 - 0xe0
      12'hCEC: dout  = 8'b11100000; // 3308 : 224 - 0xe0
      12'hCED: dout  = 8'b11100000; // 3309 : 224 - 0xe0
      12'hCEE: dout  = 8'b11100000; // 3310 : 224 - 0xe0
      12'hCEF: dout  = 8'b11100000; // 3311 : 224 - 0xe0
      12'hCF0: dout  = 8'b00000000; // 3312 :   0 - 0x0 -- Background 0x9e
      12'hCF1: dout  = 8'b00001111; // 3313 :  15 - 0xf
      12'hCF2: dout  = 8'b00001111; // 3314 :  15 - 0xf
      12'hCF3: dout  = 8'b00001111; // 3315 :  15 - 0xf
      12'hCF4: dout  = 8'b00001111; // 3316 :  15 - 0xf
      12'hCF5: dout  = 8'b00001111; // 3317 :  15 - 0xf
      12'hCF6: dout  = 8'b00001111; // 3318 :  15 - 0xf
      12'hCF7: dout  = 8'b00001111; // 3319 :  15 - 0xf
      12'hCF8: dout  = 8'b01001000; // 3320 :  72 - 0x48 -- Background 0x9f
      12'hCF9: dout  = 8'b01001000; // 3321 :  72 - 0x48
      12'hCFA: dout  = 8'b01101100; // 3322 : 108 - 0x6c
      12'hCFB: dout  = 8'b00000000; // 3323 :   0 - 0x0
      12'hCFC: dout  = 8'b00000000; // 3324 :   0 - 0x0
      12'hCFD: dout  = 8'b00000000; // 3325 :   0 - 0x0
      12'hCFE: dout  = 8'b11111110; // 3326 : 254 - 0xfe
      12'hCFF: dout  = 8'b00000000; // 3327 :   0 - 0x0
      12'hD00: dout  = 8'b00000101; // 3328 :   5 - 0x5 -- Background 0xa0
      12'hD01: dout  = 8'b00000101; // 3329 :   5 - 0x5
      12'hD02: dout  = 8'b11000101; // 3330 : 197 - 0xc5
      12'hD03: dout  = 8'b11110101; // 3331 : 245 - 0xf5
      12'hD04: dout  = 8'b11110100; // 3332 : 244 - 0xf4
      12'hD05: dout  = 8'b00000100; // 3333 :   4 - 0x4
      12'hD06: dout  = 8'b00000100; // 3334 :   4 - 0x4
      12'hD07: dout  = 8'b00000100; // 3335 :   4 - 0x4
      12'hD08: dout  = 8'b01110000; // 3336 : 112 - 0x70 -- Background 0xa1
      12'hD09: dout  = 8'b01110000; // 3337 : 112 - 0x70
      12'hD0A: dout  = 8'b01110000; // 3338 : 112 - 0x70
      12'hD0B: dout  = 8'b01111111; // 3339 : 127 - 0x7f
      12'hD0C: dout  = 8'b01111111; // 3340 : 127 - 0x7f
      12'hD0D: dout  = 8'b01110000; // 3341 : 112 - 0x70
      12'hD0E: dout  = 8'b01110000; // 3342 : 112 - 0x70
      12'hD0F: dout  = 8'b01110000; // 3343 : 112 - 0x70
      12'hD10: dout  = 8'b00000000; // 3344 :   0 - 0x0 -- Background 0xa2
      12'hD11: dout  = 8'b00000000; // 3345 :   0 - 0x0
      12'hD12: dout  = 8'b00000000; // 3346 :   0 - 0x0
      12'hD13: dout  = 8'b00000000; // 3347 :   0 - 0x0
      12'hD14: dout  = 8'b00000000; // 3348 :   0 - 0x0
      12'hD15: dout  = 8'b00000000; // 3349 :   0 - 0x0
      12'hD16: dout  = 8'b00000000; // 3350 :   0 - 0x0
      12'hD17: dout  = 8'b00000000; // 3351 :   0 - 0x0
      12'hD18: dout  = 8'b00000000; // 3352 :   0 - 0x0 -- Background 0xa3
      12'hD19: dout  = 8'b00000000; // 3353 :   0 - 0x0
      12'hD1A: dout  = 8'b00000000; // 3354 :   0 - 0x0
      12'hD1B: dout  = 8'b00000000; // 3355 :   0 - 0x0
      12'hD1C: dout  = 8'b00000000; // 3356 :   0 - 0x0
      12'hD1D: dout  = 8'b00000000; // 3357 :   0 - 0x0
      12'hD1E: dout  = 8'b00000000; // 3358 :   0 - 0x0
      12'hD1F: dout  = 8'b00000000; // 3359 :   0 - 0x0
      12'hD20: dout  = 8'b11111111; // 3360 : 255 - 0xff -- Background 0xa4
      12'hD21: dout  = 8'b11111111; // 3361 : 255 - 0xff
      12'hD22: dout  = 8'b11111111; // 3362 : 255 - 0xff
      12'hD23: dout  = 8'b11111111; // 3363 : 255 - 0xff
      12'hD24: dout  = 8'b11111111; // 3364 : 255 - 0xff
      12'hD25: dout  = 8'b11111110; // 3365 : 254 - 0xfe
      12'hD26: dout  = 8'b10111110; // 3366 : 190 - 0xbe
      12'hD27: dout  = 8'b11001110; // 3367 : 206 - 0xce
      12'hD28: dout  = 8'b00000000; // 3368 :   0 - 0x0 -- Background 0xa5
      12'hD29: dout  = 8'b00000000; // 3369 :   0 - 0x0
      12'hD2A: dout  = 8'b00000000; // 3370 :   0 - 0x0
      12'hD2B: dout  = 8'b00000000; // 3371 :   0 - 0x0
      12'hD2C: dout  = 8'b00000011; // 3372 :   3 - 0x3
      12'hD2D: dout  = 8'b00000100; // 3373 :   4 - 0x4
      12'hD2E: dout  = 8'b00000100; // 3374 :   4 - 0x4
      12'hD2F: dout  = 8'b00000100; // 3375 :   4 - 0x4
      12'hD30: dout  = 8'b00000000; // 3376 :   0 - 0x0 -- Background 0xa6
      12'hD31: dout  = 8'b00000000; // 3377 :   0 - 0x0
      12'hD32: dout  = 8'b01100000; // 3378 :  96 - 0x60
      12'hD33: dout  = 8'b00110000; // 3379 :  48 - 0x30
      12'hD34: dout  = 8'b00110000; // 3380 :  48 - 0x30
      12'hD35: dout  = 8'b10011000; // 3381 : 152 - 0x98
      12'hD36: dout  = 8'b10011000; // 3382 : 152 - 0x98
      12'hD37: dout  = 8'b10011000; // 3383 : 152 - 0x98
      12'hD38: dout  = 8'b00000100; // 3384 :   4 - 0x4 -- Background 0xa7
      12'hD39: dout  = 8'b00000100; // 3385 :   4 - 0x4
      12'hD3A: dout  = 8'b00000100; // 3386 :   4 - 0x4
      12'hD3B: dout  = 8'b00000100; // 3387 :   4 - 0x4
      12'hD3C: dout  = 8'b00000100; // 3388 :   4 - 0x4
      12'hD3D: dout  = 8'b00000011; // 3389 :   3 - 0x3
      12'hD3E: dout  = 8'b00000000; // 3390 :   0 - 0x0
      12'hD3F: dout  = 8'b00000000; // 3391 :   0 - 0x0
      12'hD40: dout  = 8'b10011000; // 3392 : 152 - 0x98 -- Background 0xa8
      12'hD41: dout  = 8'b10011000; // 3393 : 152 - 0x98
      12'hD42: dout  = 8'b10011000; // 3394 : 152 - 0x98
      12'hD43: dout  = 8'b10011000; // 3395 : 152 - 0x98
      12'hD44: dout  = 8'b10011000; // 3396 : 152 - 0x98
      12'hD45: dout  = 8'b00110000; // 3397 :  48 - 0x30
      12'hD46: dout  = 8'b00110000; // 3398 :  48 - 0x30
      12'hD47: dout  = 8'b01100000; // 3399 :  96 - 0x60
      12'hD48: dout  = 8'b00001111; // 3400 :  15 - 0xf -- Background 0xa9
      12'hD49: dout  = 8'b11101111; // 3401 : 239 - 0xef
      12'hD4A: dout  = 8'b11101111; // 3402 : 239 - 0xef
      12'hD4B: dout  = 8'b11101111; // 3403 : 239 - 0xef
      12'hD4C: dout  = 8'b11101111; // 3404 : 239 - 0xef
      12'hD4D: dout  = 8'b11101111; // 3405 : 239 - 0xef
      12'hD4E: dout  = 8'b11101111; // 3406 : 239 - 0xef
      12'hD4F: dout  = 8'b11100000; // 3407 : 224 - 0xe0
      12'hD50: dout  = 8'b11100000; // 3408 : 224 - 0xe0 -- Background 0xaa
      12'hD51: dout  = 8'b11101111; // 3409 : 239 - 0xef
      12'hD52: dout  = 8'b11101111; // 3410 : 239 - 0xef
      12'hD53: dout  = 8'b11101111; // 3411 : 239 - 0xef
      12'hD54: dout  = 8'b11101111; // 3412 : 239 - 0xef
      12'hD55: dout  = 8'b11101111; // 3413 : 239 - 0xef
      12'hD56: dout  = 8'b11101111; // 3414 : 239 - 0xef
      12'hD57: dout  = 8'b00001111; // 3415 :  15 - 0xf
      12'hD58: dout  = 8'b10000000; // 3416 : 128 - 0x80 -- Background 0xab
      12'hD59: dout  = 8'b01000000; // 3417 :  64 - 0x40
      12'hD5A: dout  = 8'b00100000; // 3418 :  32 - 0x20
      12'hD5B: dout  = 8'b00010000; // 3419 :  16 - 0x10
      12'hD5C: dout  = 8'b00001111; // 3420 :  15 - 0xf
      12'hD5D: dout  = 8'b00001111; // 3421 :  15 - 0xf
      12'hD5E: dout  = 8'b00001111; // 3422 :  15 - 0xf
      12'hD5F: dout  = 8'b00001111; // 3423 :  15 - 0xf
      12'hD60: dout  = 8'b00001111; // 3424 :  15 - 0xf -- Background 0xac
      12'hD61: dout  = 8'b00001111; // 3425 :  15 - 0xf
      12'hD62: dout  = 8'b00001111; // 3426 :  15 - 0xf
      12'hD63: dout  = 8'b00001111; // 3427 :  15 - 0xf
      12'hD64: dout  = 8'b00011111; // 3428 :  31 - 0x1f
      12'hD65: dout  = 8'b00111111; // 3429 :  63 - 0x3f
      12'hD66: dout  = 8'b01111111; // 3430 : 127 - 0x7f
      12'hD67: dout  = 8'b11111111; // 3431 : 255 - 0xff
      12'hD68: dout  = 8'b00000001; // 3432 :   1 - 0x1 -- Background 0xad
      12'hD69: dout  = 8'b00000011; // 3433 :   3 - 0x3
      12'hD6A: dout  = 8'b00000111; // 3434 :   7 - 0x7
      12'hD6B: dout  = 8'b00001111; // 3435 :  15 - 0xf
      12'hD6C: dout  = 8'b11111111; // 3436 : 255 - 0xff
      12'hD6D: dout  = 8'b11111111; // 3437 : 255 - 0xff
      12'hD6E: dout  = 8'b11111111; // 3438 : 255 - 0xff
      12'hD6F: dout  = 8'b11111111; // 3439 : 255 - 0xff
      12'hD70: dout  = 8'b11111111; // 3440 : 255 - 0xff -- Background 0xae
      12'hD71: dout  = 8'b11111111; // 3441 : 255 - 0xff
      12'hD72: dout  = 8'b11111111; // 3442 : 255 - 0xff
      12'hD73: dout  = 8'b11111111; // 3443 : 255 - 0xff
      12'hD74: dout  = 8'b11111111; // 3444 : 255 - 0xff
      12'hD75: dout  = 8'b11111111; // 3445 : 255 - 0xff
      12'hD76: dout  = 8'b11111111; // 3446 : 255 - 0xff
      12'hD77: dout  = 8'b11111111; // 3447 : 255 - 0xff
      12'hD78: dout  = 8'b00000000; // 3448 :   0 - 0x0 -- Background 0xaf
      12'hD79: dout  = 8'b00000000; // 3449 :   0 - 0x0
      12'hD7A: dout  = 8'b00000000; // 3450 :   0 - 0x0
      12'hD7B: dout  = 8'b00000000; // 3451 :   0 - 0x0
      12'hD7C: dout  = 8'b00000000; // 3452 :   0 - 0x0
      12'hD7D: dout  = 8'b00000000; // 3453 :   0 - 0x0
      12'hD7E: dout  = 8'b00000000; // 3454 :   0 - 0x0
      12'hD7F: dout  = 8'b00000000; // 3455 :   0 - 0x0
      12'hD80: dout  = 8'b00011111; // 3456 :  31 - 0x1f -- Background 0xb0
      12'hD81: dout  = 8'b00100000; // 3457 :  32 - 0x20
      12'hD82: dout  = 8'b01000000; // 3458 :  64 - 0x40
      12'hD83: dout  = 8'b01000000; // 3459 :  64 - 0x40
      12'hD84: dout  = 8'b01000000; // 3460 :  64 - 0x40
      12'hD85: dout  = 8'b10000000; // 3461 : 128 - 0x80
      12'hD86: dout  = 8'b10000010; // 3462 : 130 - 0x82
      12'hD87: dout  = 8'b10000010; // 3463 : 130 - 0x82
      12'hD88: dout  = 8'b10000010; // 3464 : 130 - 0x82 -- Background 0xb1
      12'hD89: dout  = 8'b10000000; // 3465 : 128 - 0x80
      12'hD8A: dout  = 8'b10100000; // 3466 : 160 - 0xa0
      12'hD8B: dout  = 8'b01000100; // 3467 :  68 - 0x44
      12'hD8C: dout  = 8'b01000011; // 3468 :  67 - 0x43
      12'hD8D: dout  = 8'b01000000; // 3469 :  64 - 0x40
      12'hD8E: dout  = 8'b00100001; // 3470 :  33 - 0x21
      12'hD8F: dout  = 8'b00011110; // 3471 :  30 - 0x1e
      12'hD90: dout  = 8'b11111000; // 3472 : 248 - 0xf8 -- Background 0xb2
      12'hD91: dout  = 8'b00000100; // 3473 :   4 - 0x4
      12'hD92: dout  = 8'b00000010; // 3474 :   2 - 0x2
      12'hD93: dout  = 8'b00000010; // 3475 :   2 - 0x2
      12'hD94: dout  = 8'b00000010; // 3476 :   2 - 0x2
      12'hD95: dout  = 8'b00000001; // 3477 :   1 - 0x1
      12'hD96: dout  = 8'b01000001; // 3478 :  65 - 0x41
      12'hD97: dout  = 8'b01000001; // 3479 :  65 - 0x41
      12'hD98: dout  = 8'b01000001; // 3480 :  65 - 0x41 -- Background 0xb3
      12'hD99: dout  = 8'b00000001; // 3481 :   1 - 0x1
      12'hD9A: dout  = 8'b00000101; // 3482 :   5 - 0x5
      12'hD9B: dout  = 8'b00100010; // 3483 :  34 - 0x22
      12'hD9C: dout  = 8'b11000010; // 3484 : 194 - 0xc2
      12'hD9D: dout  = 8'b00000010; // 3485 :   2 - 0x2
      12'hD9E: dout  = 8'b10000100; // 3486 : 132 - 0x84
      12'hD9F: dout  = 8'b01111000; // 3487 : 120 - 0x78
      12'hDA0: dout  = 8'b10000000; // 3488 : 128 - 0x80 -- Background 0xb4
      12'hDA1: dout  = 8'b01111111; // 3489 : 127 - 0x7f
      12'hDA2: dout  = 8'b01111111; // 3490 : 127 - 0x7f
      12'hDA3: dout  = 8'b01111111; // 3491 : 127 - 0x7f
      12'hDA4: dout  = 8'b01111111; // 3492 : 127 - 0x7f
      12'hDA5: dout  = 8'b01111111; // 3493 : 127 - 0x7f
      12'hDA6: dout  = 8'b01111111; // 3494 : 127 - 0x7f
      12'hDA7: dout  = 8'b01111111; // 3495 : 127 - 0x7f
      12'hDA8: dout  = 8'b01100001; // 3496 :  97 - 0x61 -- Background 0xb5
      12'hDA9: dout  = 8'b11011111; // 3497 : 223 - 0xdf
      12'hDAA: dout  = 8'b11011111; // 3498 : 223 - 0xdf
      12'hDAB: dout  = 8'b11011111; // 3499 : 223 - 0xdf
      12'hDAC: dout  = 8'b11011111; // 3500 : 223 - 0xdf
      12'hDAD: dout  = 8'b11111111; // 3501 : 255 - 0xff
      12'hDAE: dout  = 8'b11000001; // 3502 : 193 - 0xc1
      12'hDAF: dout  = 8'b11011111; // 3503 : 223 - 0xdf
      12'hDB0: dout  = 8'b01111111; // 3504 : 127 - 0x7f -- Background 0xb6
      12'hDB1: dout  = 8'b01111111; // 3505 : 127 - 0x7f
      12'hDB2: dout  = 8'b11111111; // 3506 : 255 - 0xff
      12'hDB3: dout  = 8'b00111111; // 3507 :  63 - 0x3f
      12'hDB4: dout  = 8'b01001111; // 3508 :  79 - 0x4f
      12'hDB5: dout  = 8'b01110001; // 3509 : 113 - 0x71
      12'hDB6: dout  = 8'b01111111; // 3510 : 127 - 0x7f
      12'hDB7: dout  = 8'b11111111; // 3511 : 255 - 0xff
      12'hDB8: dout  = 8'b11011111; // 3512 : 223 - 0xdf -- Background 0xb7
      12'hDB9: dout  = 8'b11011111; // 3513 : 223 - 0xdf
      12'hDBA: dout  = 8'b10111111; // 3514 : 191 - 0xbf
      12'hDBB: dout  = 8'b10111111; // 3515 : 191 - 0xbf
      12'hDBC: dout  = 8'b01111111; // 3516 : 127 - 0x7f
      12'hDBD: dout  = 8'b01111111; // 3517 : 127 - 0x7f
      12'hDBE: dout  = 8'b01111111; // 3518 : 127 - 0x7f
      12'hDBF: dout  = 8'b01111111; // 3519 : 127 - 0x7f
      12'hDC0: dout  = 8'b00000000; // 3520 :   0 - 0x0 -- Background 0xb8
      12'hDC1: dout  = 8'b00000000; // 3521 :   0 - 0x0
      12'hDC2: dout  = 8'b00000011; // 3522 :   3 - 0x3
      12'hDC3: dout  = 8'b00001100; // 3523 :  12 - 0xc
      12'hDC4: dout  = 8'b00010000; // 3524 :  16 - 0x10
      12'hDC5: dout  = 8'b00100000; // 3525 :  32 - 0x20
      12'hDC6: dout  = 8'b01000000; // 3526 :  64 - 0x40
      12'hDC7: dout  = 8'b01000000; // 3527 :  64 - 0x40
      12'hDC8: dout  = 8'b00000000; // 3528 :   0 - 0x0 -- Background 0xb9
      12'hDC9: dout  = 8'b00000000; // 3529 :   0 - 0x0
      12'hDCA: dout  = 8'b11000000; // 3530 : 192 - 0xc0
      12'hDCB: dout  = 8'b00110000; // 3531 :  48 - 0x30
      12'hDCC: dout  = 8'b00001000; // 3532 :   8 - 0x8
      12'hDCD: dout  = 8'b00000100; // 3533 :   4 - 0x4
      12'hDCE: dout  = 8'b00000010; // 3534 :   2 - 0x2
      12'hDCF: dout  = 8'b00000010; // 3535 :   2 - 0x2
      12'hDD0: dout  = 8'b10000000; // 3536 : 128 - 0x80 -- Background 0xba
      12'hDD1: dout  = 8'b10000000; // 3537 : 128 - 0x80
      12'hDD2: dout  = 8'b10000000; // 3538 : 128 - 0x80
      12'hDD3: dout  = 8'b10000000; // 3539 : 128 - 0x80
      12'hDD4: dout  = 8'b10000000; // 3540 : 128 - 0x80
      12'hDD5: dout  = 8'b10000000; // 3541 : 128 - 0x80
      12'hDD6: dout  = 8'b10000000; // 3542 : 128 - 0x80
      12'hDD7: dout  = 8'b10000000; // 3543 : 128 - 0x80
      12'hDD8: dout  = 8'b00000001; // 3544 :   1 - 0x1 -- Background 0xbb
      12'hDD9: dout  = 8'b00000001; // 3545 :   1 - 0x1
      12'hDDA: dout  = 8'b00000001; // 3546 :   1 - 0x1
      12'hDDB: dout  = 8'b00000001; // 3547 :   1 - 0x1
      12'hDDC: dout  = 8'b00000001; // 3548 :   1 - 0x1
      12'hDDD: dout  = 8'b00000001; // 3549 :   1 - 0x1
      12'hDDE: dout  = 8'b00000001; // 3550 :   1 - 0x1
      12'hDDF: dout  = 8'b00000001; // 3551 :   1 - 0x1
      12'hDE0: dout  = 8'b01000000; // 3552 :  64 - 0x40 -- Background 0xbc
      12'hDE1: dout  = 8'b01000000; // 3553 :  64 - 0x40
      12'hDE2: dout  = 8'b01000000; // 3554 :  64 - 0x40
      12'hDE3: dout  = 8'b00100000; // 3555 :  32 - 0x20
      12'hDE4: dout  = 8'b00110000; // 3556 :  48 - 0x30
      12'hDE5: dout  = 8'b00011100; // 3557 :  28 - 0x1c
      12'hDE6: dout  = 8'b00001111; // 3558 :  15 - 0xf
      12'hDE7: dout  = 8'b00000111; // 3559 :   7 - 0x7
      12'hDE8: dout  = 8'b00000010; // 3560 :   2 - 0x2 -- Background 0xbd
      12'hDE9: dout  = 8'b00000010; // 3561 :   2 - 0x2
      12'hDEA: dout  = 8'b00000010; // 3562 :   2 - 0x2
      12'hDEB: dout  = 8'b00000100; // 3563 :   4 - 0x4
      12'hDEC: dout  = 8'b00001100; // 3564 :  12 - 0xc
      12'hDED: dout  = 8'b00111000; // 3565 :  56 - 0x38
      12'hDEE: dout  = 8'b11110000; // 3566 : 240 - 0xf0
      12'hDEF: dout  = 8'b11110000; // 3567 : 240 - 0xf0
      12'hDF0: dout  = 8'b00001000; // 3568 :   8 - 0x8 -- Background 0xbe
      12'hDF1: dout  = 8'b00001000; // 3569 :   8 - 0x8
      12'hDF2: dout  = 8'b00001000; // 3570 :   8 - 0x8
      12'hDF3: dout  = 8'b00001000; // 3571 :   8 - 0x8
      12'hDF4: dout  = 8'b00001000; // 3572 :   8 - 0x8
      12'hDF5: dout  = 8'b00001100; // 3573 :  12 - 0xc
      12'hDF6: dout  = 8'b00000101; // 3574 :   5 - 0x5
      12'hDF7: dout  = 8'b00001010; // 3575 :  10 - 0xa
      12'hDF8: dout  = 8'b00010000; // 3576 :  16 - 0x10 -- Background 0xbf
      12'hDF9: dout  = 8'b01010000; // 3577 :  80 - 0x50
      12'hDFA: dout  = 8'b01010000; // 3578 :  80 - 0x50
      12'hDFB: dout  = 8'b01010000; // 3579 :  80 - 0x50
      12'hDFC: dout  = 8'b01010000; // 3580 :  80 - 0x50
      12'hDFD: dout  = 8'b00110000; // 3581 :  48 - 0x30
      12'hDFE: dout  = 8'b10100000; // 3582 : 160 - 0xa0
      12'hDFF: dout  = 8'b01010000; // 3583 :  80 - 0x50
      12'hE00: dout  = 8'b00000000; // 3584 :   0 - 0x0 -- Background 0xc0
      12'hE01: dout  = 8'b01000001; // 3585 :  65 - 0x41
      12'hE02: dout  = 8'b00100010; // 3586 :  34 - 0x22
      12'hE03: dout  = 8'b00100010; // 3587 :  34 - 0x22
      12'hE04: dout  = 8'b00011100; // 3588 :  28 - 0x1c
      12'hE05: dout  = 8'b00000000; // 3589 :   0 - 0x0
      12'hE06: dout  = 8'b00000000; // 3590 :   0 - 0x0
      12'hE07: dout  = 8'b00000000; // 3591 :   0 - 0x0
      12'hE08: dout  = 8'b11100011; // 3592 : 227 - 0xe3 -- Background 0xc1
      12'hE09: dout  = 8'b00010100; // 3593 :  20 - 0x14
      12'hE0A: dout  = 8'b00111110; // 3594 :  62 - 0x3e
      12'hE0B: dout  = 8'b00111110; // 3595 :  62 - 0x3e
      12'hE0C: dout  = 8'b00111110; // 3596 :  62 - 0x3e
      12'hE0D: dout  = 8'b00111110; // 3597 :  62 - 0x3e
      12'hE0E: dout  = 8'b00010100; // 3598 :  20 - 0x14
      12'hE0F: dout  = 8'b11100011; // 3599 : 227 - 0xe3
      12'hE10: dout  = 8'b11111111; // 3600 : 255 - 0xff -- Background 0xc2
      12'hE11: dout  = 8'b11111111; // 3601 : 255 - 0xff
      12'hE12: dout  = 8'b11111000; // 3602 : 248 - 0xf8
      12'hE13: dout  = 8'b11110000; // 3603 : 240 - 0xf0
      12'hE14: dout  = 8'b11110000; // 3604 : 240 - 0xf0
      12'hE15: dout  = 8'b11100000; // 3605 : 224 - 0xe0
      12'hE16: dout  = 8'b11100000; // 3606 : 224 - 0xe0
      12'hE17: dout  = 8'b11100000; // 3607 : 224 - 0xe0
      12'hE18: dout  = 8'b11111111; // 3608 : 255 - 0xff -- Background 0xc3
      12'hE19: dout  = 8'b11111111; // 3609 : 255 - 0xff
      12'hE1A: dout  = 8'b01111111; // 3610 : 127 - 0x7f
      12'hE1B: dout  = 8'b00111111; // 3611 :  63 - 0x3f
      12'hE1C: dout  = 8'b00111111; // 3612 :  63 - 0x3f
      12'hE1D: dout  = 8'b10011111; // 3613 : 159 - 0x9f
      12'hE1E: dout  = 8'b10011111; // 3614 : 159 - 0x9f
      12'hE1F: dout  = 8'b10011111; // 3615 : 159 - 0x9f
      12'hE20: dout  = 8'b11100000; // 3616 : 224 - 0xe0 -- Background 0xc4
      12'hE21: dout  = 8'b11100000; // 3617 : 224 - 0xe0
      12'hE22: dout  = 8'b11100000; // 3618 : 224 - 0xe0
      12'hE23: dout  = 8'b11100000; // 3619 : 224 - 0xe0
      12'hE24: dout  = 8'b11100000; // 3620 : 224 - 0xe0
      12'hE25: dout  = 8'b11110011; // 3621 : 243 - 0xf3
      12'hE26: dout  = 8'b11110000; // 3622 : 240 - 0xf0
      12'hE27: dout  = 8'b11111000; // 3623 : 248 - 0xf8
      12'hE28: dout  = 8'b10011111; // 3624 : 159 - 0x9f -- Background 0xc5
      12'hE29: dout  = 8'b10011111; // 3625 : 159 - 0x9f
      12'hE2A: dout  = 8'b10011111; // 3626 : 159 - 0x9f
      12'hE2B: dout  = 8'b10011111; // 3627 : 159 - 0x9f
      12'hE2C: dout  = 8'b10011111; // 3628 : 159 - 0x9f
      12'hE2D: dout  = 8'b00111111; // 3629 :  63 - 0x3f
      12'hE2E: dout  = 8'b00111111; // 3630 :  63 - 0x3f
      12'hE2F: dout  = 8'b01111111; // 3631 : 127 - 0x7f
      12'hE30: dout  = 8'b00000000; // 3632 :   0 - 0x0 -- Background 0xc6
      12'hE31: dout  = 8'b01110000; // 3633 : 112 - 0x70
      12'hE32: dout  = 8'b00011111; // 3634 :  31 - 0x1f
      12'hE33: dout  = 8'b00010000; // 3635 :  16 - 0x10
      12'hE34: dout  = 8'b01110000; // 3636 : 112 - 0x70
      12'hE35: dout  = 8'b01111111; // 3637 : 127 - 0x7f
      12'hE36: dout  = 8'b01111111; // 3638 : 127 - 0x7f
      12'hE37: dout  = 8'b01111111; // 3639 : 127 - 0x7f
      12'hE38: dout  = 8'b00000000; // 3640 :   0 - 0x0 -- Background 0xc7
      12'hE39: dout  = 8'b00000011; // 3641 :   3 - 0x3
      12'hE3A: dout  = 8'b11111000; // 3642 : 248 - 0xf8
      12'hE3B: dout  = 8'b00000000; // 3643 :   0 - 0x0
      12'hE3C: dout  = 8'b00000011; // 3644 :   3 - 0x3
      12'hE3D: dout  = 8'b11111011; // 3645 : 251 - 0xfb
      12'hE3E: dout  = 8'b11111011; // 3646 : 251 - 0xfb
      12'hE3F: dout  = 8'b11111011; // 3647 : 251 - 0xfb
      12'hE40: dout  = 8'b01111100; // 3648 : 124 - 0x7c -- Background 0xc8
      12'hE41: dout  = 8'b01111011; // 3649 : 123 - 0x7b
      12'hE42: dout  = 8'b01110110; // 3650 : 118 - 0x76
      12'hE43: dout  = 8'b01110101; // 3651 : 117 - 0x75
      12'hE44: dout  = 8'b01110101; // 3652 : 117 - 0x75
      12'hE45: dout  = 8'b01110111; // 3653 : 119 - 0x77
      12'hE46: dout  = 8'b00010111; // 3654 :  23 - 0x17
      12'hE47: dout  = 8'b01100111; // 3655 : 103 - 0x67
      12'hE48: dout  = 8'b00111011; // 3656 :  59 - 0x3b -- Background 0xc9
      12'hE49: dout  = 8'b11111011; // 3657 : 251 - 0xfb
      12'hE4A: dout  = 8'b01111011; // 3658 : 123 - 0x7b
      12'hE4B: dout  = 8'b11111011; // 3659 : 251 - 0xfb
      12'hE4C: dout  = 8'b11111011; // 3660 : 251 - 0xfb
      12'hE4D: dout  = 8'b11110011; // 3661 : 243 - 0xf3
      12'hE4E: dout  = 8'b11111000; // 3662 : 248 - 0xf8
      12'hE4F: dout  = 8'b11110011; // 3663 : 243 - 0xf3
      12'hE50: dout  = 8'b00001111; // 3664 :  15 - 0xf -- Background 0xca
      12'hE51: dout  = 8'b00001111; // 3665 :  15 - 0xf
      12'hE52: dout  = 8'b00011111; // 3666 :  31 - 0x1f
      12'hE53: dout  = 8'b00011111; // 3667 :  31 - 0x1f
      12'hE54: dout  = 8'b00111111; // 3668 :  63 - 0x3f
      12'hE55: dout  = 8'b00111100; // 3669 :  60 - 0x3c
      12'hE56: dout  = 8'b01111000; // 3670 : 120 - 0x78
      12'hE57: dout  = 8'b01111010; // 3671 : 122 - 0x7a
      12'hE58: dout  = 8'b11111000; // 3672 : 248 - 0xf8 -- Background 0xcb
      12'hE59: dout  = 8'b11111000; // 3673 : 248 - 0xf8
      12'hE5A: dout  = 8'b11111100; // 3674 : 252 - 0xfc
      12'hE5B: dout  = 8'b11111100; // 3675 : 252 - 0xfc
      12'hE5C: dout  = 8'b11111110; // 3676 : 254 - 0xfe
      12'hE5D: dout  = 8'b00111110; // 3677 :  62 - 0x3e
      12'hE5E: dout  = 8'b00011110; // 3678 :  30 - 0x1e
      12'hE5F: dout  = 8'b01011111; // 3679 :  95 - 0x5f
      12'hE60: dout  = 8'b01110110; // 3680 : 118 - 0x76 -- Background 0xcc
      12'hE61: dout  = 8'b01110110; // 3681 : 118 - 0x76
      12'hE62: dout  = 8'b01110110; // 3682 : 118 - 0x76
      12'hE63: dout  = 8'b01110000; // 3683 : 112 - 0x70
      12'hE64: dout  = 8'b01111101; // 3684 : 125 - 0x7d
      12'hE65: dout  = 8'b01111100; // 3685 : 124 - 0x7c
      12'hE66: dout  = 8'b01111111; // 3686 : 127 - 0x7f
      12'hE67: dout  = 8'b01111111; // 3687 : 127 - 0x7f
      12'hE68: dout  = 8'b01101111; // 3688 : 111 - 0x6f -- Background 0xcd
      12'hE69: dout  = 8'b01101111; // 3689 : 111 - 0x6f
      12'hE6A: dout  = 8'b01101111; // 3690 : 111 - 0x6f
      12'hE6B: dout  = 8'b00001111; // 3691 :  15 - 0xf
      12'hE6C: dout  = 8'b10111111; // 3692 : 191 - 0xbf
      12'hE6D: dout  = 8'b00111111; // 3693 :  63 - 0x3f
      12'hE6E: dout  = 8'b11111111; // 3694 : 255 - 0xff
      12'hE6F: dout  = 8'b11111111; // 3695 : 255 - 0xff
      12'hE70: dout  = 8'b00111100; // 3696 :  60 - 0x3c -- Background 0xce
      12'hE71: dout  = 8'b01111110; // 3697 : 126 - 0x7e
      12'hE72: dout  = 8'b01111110; // 3698 : 126 - 0x7e
      12'hE73: dout  = 8'b11111111; // 3699 : 255 - 0xff
      12'hE74: dout  = 8'b11111111; // 3700 : 255 - 0xff
      12'hE75: dout  = 8'b11111111; // 3701 : 255 - 0xff
      12'hE76: dout  = 8'b01000010; // 3702 :  66 - 0x42
      12'hE77: dout  = 8'b00000000; // 3703 :   0 - 0x0
      12'hE78: dout  = 8'b00000000; // 3704 :   0 - 0x0 -- Background 0xcf
      12'hE79: dout  = 8'b00000000; // 3705 :   0 - 0x0
      12'hE7A: dout  = 8'b00000000; // 3706 :   0 - 0x0
      12'hE7B: dout  = 8'b00000000; // 3707 :   0 - 0x0
      12'hE7C: dout  = 8'b00000000; // 3708 :   0 - 0x0
      12'hE7D: dout  = 8'b00000000; // 3709 :   0 - 0x0
      12'hE7E: dout  = 8'b00000000; // 3710 :   0 - 0x0
      12'hE7F: dout  = 8'b00000000; // 3711 :   0 - 0x0
      12'hE80: dout  = 8'b11110000; // 3712 : 240 - 0xf0 -- Background 0xd0
      12'hE81: dout  = 8'b11100000; // 3713 : 224 - 0xe0
      12'hE82: dout  = 8'b11100000; // 3714 : 224 - 0xe0
      12'hE83: dout  = 8'b11000000; // 3715 : 192 - 0xc0
      12'hE84: dout  = 8'b11000000; // 3716 : 192 - 0xc0
      12'hE85: dout  = 8'b10000000; // 3717 : 128 - 0x80
      12'hE86: dout  = 8'b10000000; // 3718 : 128 - 0x80
      12'hE87: dout  = 8'b10000000; // 3719 : 128 - 0x80
      12'hE88: dout  = 8'b00001111; // 3720 :  15 - 0xf -- Background 0xd1
      12'hE89: dout  = 8'b00000111; // 3721 :   7 - 0x7
      12'hE8A: dout  = 8'b00000111; // 3722 :   7 - 0x7
      12'hE8B: dout  = 8'b00000011; // 3723 :   3 - 0x3
      12'hE8C: dout  = 8'b00000011; // 3724 :   3 - 0x3
      12'hE8D: dout  = 8'b00000001; // 3725 :   1 - 0x1
      12'hE8E: dout  = 8'b00000001; // 3726 :   1 - 0x1
      12'hE8F: dout  = 8'b00000001; // 3727 :   1 - 0x1
      12'hE90: dout  = 8'b10000000; // 3728 : 128 - 0x80 -- Background 0xd2
      12'hE91: dout  = 8'b10000000; // 3729 : 128 - 0x80
      12'hE92: dout  = 8'b11000000; // 3730 : 192 - 0xc0
      12'hE93: dout  = 8'b11000000; // 3731 : 192 - 0xc0
      12'hE94: dout  = 8'b11100000; // 3732 : 224 - 0xe0
      12'hE95: dout  = 8'b11111000; // 3733 : 248 - 0xf8
      12'hE96: dout  = 8'b11111110; // 3734 : 254 - 0xfe
      12'hE97: dout  = 8'b11111111; // 3735 : 255 - 0xff
      12'hE98: dout  = 8'b11111111; // 3736 : 255 - 0xff -- Background 0xd3
      12'hE99: dout  = 8'b01111111; // 3737 : 127 - 0x7f
      12'hE9A: dout  = 8'b00011111; // 3738 :  31 - 0x1f
      12'hE9B: dout  = 8'b00000111; // 3739 :   7 - 0x7
      12'hE9C: dout  = 8'b00000011; // 3740 :   3 - 0x3
      12'hE9D: dout  = 8'b00000011; // 3741 :   3 - 0x3
      12'hE9E: dout  = 8'b00000001; // 3742 :   1 - 0x1
      12'hE9F: dout  = 8'b10000001; // 3743 : 129 - 0x81
      12'hEA0: dout  = 8'b10000000; // 3744 : 128 - 0x80 -- Background 0xd4
      12'hEA1: dout  = 8'b10000000; // 3745 : 128 - 0x80
      12'hEA2: dout  = 8'b10000000; // 3746 : 128 - 0x80
      12'hEA3: dout  = 8'b11000000; // 3747 : 192 - 0xc0
      12'hEA4: dout  = 8'b11000000; // 3748 : 192 - 0xc0
      12'hEA5: dout  = 8'b11100000; // 3749 : 224 - 0xe0
      12'hEA6: dout  = 8'b11100000; // 3750 : 224 - 0xe0
      12'hEA7: dout  = 8'b11110000; // 3751 : 240 - 0xf0
      12'hEA8: dout  = 8'b00000001; // 3752 :   1 - 0x1 -- Background 0xd5
      12'hEA9: dout  = 8'b00000001; // 3753 :   1 - 0x1
      12'hEAA: dout  = 8'b00000001; // 3754 :   1 - 0x1
      12'hEAB: dout  = 8'b00000011; // 3755 :   3 - 0x3
      12'hEAC: dout  = 8'b00000011; // 3756 :   3 - 0x3
      12'hEAD: dout  = 8'b00000111; // 3757 :   7 - 0x7
      12'hEAE: dout  = 8'b00000111; // 3758 :   7 - 0x7
      12'hEAF: dout  = 8'b00001111; // 3759 :  15 - 0xf
      12'hEB0: dout  = 8'b11111111; // 3760 : 255 - 0xff -- Background 0xd6
      12'hEB1: dout  = 8'b11111111; // 3761 : 255 - 0xff
      12'hEB2: dout  = 8'b11111111; // 3762 : 255 - 0xff
      12'hEB3: dout  = 8'b11111111; // 3763 : 255 - 0xff
      12'hEB4: dout  = 8'b11111111; // 3764 : 255 - 0xff
      12'hEB5: dout  = 8'b11111111; // 3765 : 255 - 0xff
      12'hEB6: dout  = 8'b11111111; // 3766 : 255 - 0xff
      12'hEB7: dout  = 8'b11111111; // 3767 : 255 - 0xff
      12'hEB8: dout  = 8'b11111111; // 3768 : 255 - 0xff -- Background 0xd7
      12'hEB9: dout  = 8'b11111111; // 3769 : 255 - 0xff
      12'hEBA: dout  = 8'b11111111; // 3770 : 255 - 0xff
      12'hEBB: dout  = 8'b11111111; // 3771 : 255 - 0xff
      12'hEBC: dout  = 8'b11111111; // 3772 : 255 - 0xff
      12'hEBD: dout  = 8'b11111111; // 3773 : 255 - 0xff
      12'hEBE: dout  = 8'b11111111; // 3774 : 255 - 0xff
      12'hEBF: dout  = 8'b11111111; // 3775 : 255 - 0xff
      12'hEC0: dout  = 8'b10000001; // 3776 : 129 - 0x81 -- Background 0xd8
      12'hEC1: dout  = 8'b10000001; // 3777 : 129 - 0x81
      12'hEC2: dout  = 8'b10000001; // 3778 : 129 - 0x81
      12'hEC3: dout  = 8'b10000001; // 3779 : 129 - 0x81
      12'hEC4: dout  = 8'b10000001; // 3780 : 129 - 0x81
      12'hEC5: dout  = 8'b10000001; // 3781 : 129 - 0x81
      12'hEC6: dout  = 8'b10000001; // 3782 : 129 - 0x81
      12'hEC7: dout  = 8'b10000001; // 3783 : 129 - 0x81
      12'hEC8: dout  = 8'b00000001; // 3784 :   1 - 0x1 -- Background 0xd9
      12'hEC9: dout  = 8'b00000001; // 3785 :   1 - 0x1
      12'hECA: dout  = 8'b00000001; // 3786 :   1 - 0x1
      12'hECB: dout  = 8'b00000011; // 3787 :   3 - 0x3
      12'hECC: dout  = 8'b00000011; // 3788 :   3 - 0x3
      12'hECD: dout  = 8'b00000111; // 3789 :   7 - 0x7
      12'hECE: dout  = 8'b00000111; // 3790 :   7 - 0x7
      12'hECF: dout  = 8'b00001111; // 3791 :  15 - 0xf
      12'hED0: dout  = 8'b00000001; // 3792 :   1 - 0x1 -- Background 0xda
      12'hED1: dout  = 8'b00000001; // 3793 :   1 - 0x1
      12'hED2: dout  = 8'b00000001; // 3794 :   1 - 0x1
      12'hED3: dout  = 8'b00000001; // 3795 :   1 - 0x1
      12'hED4: dout  = 8'b00000001; // 3796 :   1 - 0x1
      12'hED5: dout  = 8'b00000001; // 3797 :   1 - 0x1
      12'hED6: dout  = 8'b00000001; // 3798 :   1 - 0x1
      12'hED7: dout  = 8'b00000001; // 3799 :   1 - 0x1
      12'hED8: dout  = 8'b10000001; // 3800 : 129 - 0x81 -- Background 0xdb
      12'hED9: dout  = 8'b10000001; // 3801 : 129 - 0x81
      12'hEDA: dout  = 8'b10000001; // 3802 : 129 - 0x81
      12'hEDB: dout  = 8'b10000001; // 3803 : 129 - 0x81
      12'hEDC: dout  = 8'b10000001; // 3804 : 129 - 0x81
      12'hEDD: dout  = 8'b10000001; // 3805 : 129 - 0x81
      12'hEDE: dout  = 8'b10000001; // 3806 : 129 - 0x81
      12'hEDF: dout  = 8'b10000001; // 3807 : 129 - 0x81
      12'hEE0: dout  = 8'b11111111; // 3808 : 255 - 0xff -- Background 0xdc
      12'hEE1: dout  = 8'b00000011; // 3809 :   3 - 0x3
      12'hEE2: dout  = 8'b00000011; // 3810 :   3 - 0x3
      12'hEE3: dout  = 8'b00000011; // 3811 :   3 - 0x3
      12'hEE4: dout  = 8'b00000011; // 3812 :   3 - 0x3
      12'hEE5: dout  = 8'b00000011; // 3813 :   3 - 0x3
      12'hEE6: dout  = 8'b00000011; // 3814 :   3 - 0x3
      12'hEE7: dout  = 8'b11111111; // 3815 : 255 - 0xff
      12'hEE8: dout  = 8'b11111111; // 3816 : 255 - 0xff -- Background 0xdd
      12'hEE9: dout  = 8'b11111111; // 3817 : 255 - 0xff
      12'hEEA: dout  = 8'b11111111; // 3818 : 255 - 0xff
      12'hEEB: dout  = 8'b11111111; // 3819 : 255 - 0xff
      12'hEEC: dout  = 8'b11111111; // 3820 : 255 - 0xff
      12'hEED: dout  = 8'b11111111; // 3821 : 255 - 0xff
      12'hEEE: dout  = 8'b11111111; // 3822 : 255 - 0xff
      12'hEEF: dout  = 8'b11111111; // 3823 : 255 - 0xff
      12'hEF0: dout  = 8'b10000000; // 3824 : 128 - 0x80 -- Background 0xde
      12'hEF1: dout  = 8'b10000000; // 3825 : 128 - 0x80
      12'hEF2: dout  = 8'b10000000; // 3826 : 128 - 0x80
      12'hEF3: dout  = 8'b10000000; // 3827 : 128 - 0x80
      12'hEF4: dout  = 8'b10000000; // 3828 : 128 - 0x80
      12'hEF5: dout  = 8'b10000000; // 3829 : 128 - 0x80
      12'hEF6: dout  = 8'b10000000; // 3830 : 128 - 0x80
      12'hEF7: dout  = 8'b10000000; // 3831 : 128 - 0x80
      12'hEF8: dout  = 8'b00000001; // 3832 :   1 - 0x1 -- Background 0xdf
      12'hEF9: dout  = 8'b00000001; // 3833 :   1 - 0x1
      12'hEFA: dout  = 8'b00000001; // 3834 :   1 - 0x1
      12'hEFB: dout  = 8'b00000011; // 3835 :   3 - 0x3
      12'hEFC: dout  = 8'b00000111; // 3836 :   7 - 0x7
      12'hEFD: dout  = 8'b00000011; // 3837 :   3 - 0x3
      12'hEFE: dout  = 8'b00000001; // 3838 :   1 - 0x1
      12'hEFF: dout  = 8'b00000001; // 3839 :   1 - 0x1
      12'hF00: dout  = 8'b10000001; // 3840 : 129 - 0x81 -- Background 0xe0
      12'hF01: dout  = 8'b10000001; // 3841 : 129 - 0x81
      12'hF02: dout  = 8'b10000001; // 3842 : 129 - 0x81
      12'hF03: dout  = 8'b10000001; // 3843 : 129 - 0x81
      12'hF04: dout  = 8'b10000001; // 3844 : 129 - 0x81
      12'hF05: dout  = 8'b10000001; // 3845 : 129 - 0x81
      12'hF06: dout  = 8'b10000001; // 3846 : 129 - 0x81
      12'hF07: dout  = 8'b10000001; // 3847 : 129 - 0x81
      12'hF08: dout  = 8'b11111111; // 3848 : 255 - 0xff -- Background 0xe1
      12'hF09: dout  = 8'b11111111; // 3849 : 255 - 0xff
      12'hF0A: dout  = 8'b11111111; // 3850 : 255 - 0xff
      12'hF0B: dout  = 8'b11111111; // 3851 : 255 - 0xff
      12'hF0C: dout  = 8'b11111111; // 3852 : 255 - 0xff
      12'hF0D: dout  = 8'b11111111; // 3853 : 255 - 0xff
      12'hF0E: dout  = 8'b11111111; // 3854 : 255 - 0xff
      12'hF0F: dout  = 8'b11111111; // 3855 : 255 - 0xff
      12'hF10: dout  = 8'b11111111; // 3856 : 255 - 0xff -- Background 0xe2
      12'hF11: dout  = 8'b11111111; // 3857 : 255 - 0xff
      12'hF12: dout  = 8'b11111111; // 3858 : 255 - 0xff
      12'hF13: dout  = 8'b11111111; // 3859 : 255 - 0xff
      12'hF14: dout  = 8'b11111111; // 3860 : 255 - 0xff
      12'hF15: dout  = 8'b11111111; // 3861 : 255 - 0xff
      12'hF16: dout  = 8'b11111111; // 3862 : 255 - 0xff
      12'hF17: dout  = 8'b11111111; // 3863 : 255 - 0xff
      12'hF18: dout  = 8'b10000001; // 3864 : 129 - 0x81 -- Background 0xe3
      12'hF19: dout  = 8'b10000001; // 3865 : 129 - 0x81
      12'hF1A: dout  = 8'b10000001; // 3866 : 129 - 0x81
      12'hF1B: dout  = 8'b10000001; // 3867 : 129 - 0x81
      12'hF1C: dout  = 8'b10000001; // 3868 : 129 - 0x81
      12'hF1D: dout  = 8'b10000001; // 3869 : 129 - 0x81
      12'hF1E: dout  = 8'b10000001; // 3870 : 129 - 0x81
      12'hF1F: dout  = 8'b10000001; // 3871 : 129 - 0x81
      12'hF20: dout  = 8'b10000000; // 3872 : 128 - 0x80 -- Background 0xe4
      12'hF21: dout  = 8'b10000000; // 3873 : 128 - 0x80
      12'hF22: dout  = 8'b11000000; // 3874 : 192 - 0xc0
      12'hF23: dout  = 8'b11000000; // 3875 : 192 - 0xc0
      12'hF24: dout  = 8'b11100000; // 3876 : 224 - 0xe0
      12'hF25: dout  = 8'b11111000; // 3877 : 248 - 0xf8
      12'hF26: dout  = 8'b11111110; // 3878 : 254 - 0xfe
      12'hF27: dout  = 8'b11111111; // 3879 : 255 - 0xff
      12'hF28: dout  = 8'b11111111; // 3880 : 255 - 0xff -- Background 0xe5
      12'hF29: dout  = 8'b01111111; // 3881 : 127 - 0x7f
      12'hF2A: dout  = 8'b00011111; // 3882 :  31 - 0x1f
      12'hF2B: dout  = 8'b00000111; // 3883 :   7 - 0x7
      12'hF2C: dout  = 8'b00000011; // 3884 :   3 - 0x3
      12'hF2D: dout  = 8'b00000011; // 3885 :   3 - 0x3
      12'hF2E: dout  = 8'b00000001; // 3886 :   1 - 0x1
      12'hF2F: dout  = 8'b10000001; // 3887 : 129 - 0x81
      12'hF30: dout  = 8'b10000001; // 3888 : 129 - 0x81 -- Background 0xe6
      12'hF31: dout  = 8'b10000001; // 3889 : 129 - 0x81
      12'hF32: dout  = 8'b10000001; // 3890 : 129 - 0x81
      12'hF33: dout  = 8'b10000001; // 3891 : 129 - 0x81
      12'hF34: dout  = 8'b10000001; // 3892 : 129 - 0x81
      12'hF35: dout  = 8'b10000001; // 3893 : 129 - 0x81
      12'hF36: dout  = 8'b10000001; // 3894 : 129 - 0x81
      12'hF37: dout  = 8'b10000001; // 3895 : 129 - 0x81
      12'hF38: dout  = 8'b10000001; // 3896 : 129 - 0x81 -- Background 0xe7
      12'hF39: dout  = 8'b10000001; // 3897 : 129 - 0x81
      12'hF3A: dout  = 8'b10000001; // 3898 : 129 - 0x81
      12'hF3B: dout  = 8'b10000001; // 3899 : 129 - 0x81
      12'hF3C: dout  = 8'b10000001; // 3900 : 129 - 0x81
      12'hF3D: dout  = 8'b10000001; // 3901 : 129 - 0x81
      12'hF3E: dout  = 8'b10000001; // 3902 : 129 - 0x81
      12'hF3F: dout  = 8'b10000001; // 3903 : 129 - 0x81
      12'hF40: dout  = 8'b01111110; // 3904 : 126 - 0x7e -- Background 0xe8
      12'hF41: dout  = 8'b00111100; // 3905 :  60 - 0x3c
      12'hF42: dout  = 8'b00111100; // 3906 :  60 - 0x3c
      12'hF43: dout  = 8'b00011000; // 3907 :  24 - 0x18
      12'hF44: dout  = 8'b00011000; // 3908 :  24 - 0x18
      12'hF45: dout  = 8'b00000000; // 3909 :   0 - 0x0
      12'hF46: dout  = 8'b00000000; // 3910 :   0 - 0x0
      12'hF47: dout  = 8'b00000000; // 3911 :   0 - 0x0
      12'hF48: dout  = 8'b11110010; // 3912 : 242 - 0xf2 -- Background 0xe9
      12'hF49: dout  = 8'b11111110; // 3913 : 254 - 0xfe
      12'hF4A: dout  = 8'b11111110; // 3914 : 254 - 0xfe
      12'hF4B: dout  = 8'b11111111; // 3915 : 255 - 0xff
      12'hF4C: dout  = 8'b11111111; // 3916 : 255 - 0xff
      12'hF4D: dout  = 8'b11101111; // 3917 : 239 - 0xef
      12'hF4E: dout  = 8'b11110111; // 3918 : 247 - 0xf7
      12'hF4F: dout  = 8'b11111000; // 3919 : 248 - 0xf8
      12'hF50: dout  = 8'b10111111; // 3920 : 191 - 0xbf -- Background 0xea
      12'hF51: dout  = 8'b10111110; // 3921 : 190 - 0xbe
      12'hF52: dout  = 8'b10111101; // 3922 : 189 - 0xbd
      12'hF53: dout  = 8'b01111011; // 3923 : 123 - 0x7b
      12'hF54: dout  = 8'b01111011; // 3924 : 123 - 0x7b
      12'hF55: dout  = 8'b00000111; // 3925 :   7 - 0x7
      12'hF56: dout  = 8'b11110011; // 3926 : 243 - 0xf3
      12'hF57: dout  = 8'b11111101; // 3927 : 253 - 0xfd
      12'hF58: dout  = 8'b11111111; // 3928 : 255 - 0xff -- Background 0xeb
      12'hF59: dout  = 8'b11111111; // 3929 : 255 - 0xff
      12'hF5A: dout  = 8'b11111111; // 3930 : 255 - 0xff
      12'hF5B: dout  = 8'b01100111; // 3931 : 103 - 0x67
      12'hF5C: dout  = 8'b01011001; // 3932 :  89 - 0x59
      12'hF5D: dout  = 8'b10011110; // 3933 : 158 - 0x9e
      12'hF5E: dout  = 8'b10111111; // 3934 : 191 - 0xbf
      12'hF5F: dout  = 8'b10111111; // 3935 : 191 - 0xbf
      12'hF60: dout  = 8'b00100000; // 3936 :  32 - 0x20 -- Background 0xec
      12'hF61: dout  = 8'b11100110; // 3937 : 230 - 0xe6
      12'hF62: dout  = 8'b01010100; // 3938 :  84 - 0x54
      12'hF63: dout  = 8'b00100110; // 3939 :  38 - 0x26
      12'hF64: dout  = 8'b00100001; // 3940 :  33 - 0x21
      12'hF65: dout  = 8'b00000110; // 3941 :   6 - 0x6
      12'hF66: dout  = 8'b01010100; // 3942 :  84 - 0x54
      12'hF67: dout  = 8'b00100110; // 3943 :  38 - 0x26
      12'hF68: dout  = 8'b00100000; // 3944 :  32 - 0x20 -- Background 0xed
      12'hF69: dout  = 8'b10011010; // 3945 : 154 - 0x9a
      12'hF6A: dout  = 8'b00000001; // 3946 :   1 - 0x1
      12'hF6B: dout  = 8'b01001001; // 3947 :  73 - 0x49
      12'hF6C: dout  = 8'b00100000; // 3948 :  32 - 0x20
      12'hF6D: dout  = 8'b10100101; // 3949 : 165 - 0xa5
      12'hF6E: dout  = 8'b11001001; // 3950 : 201 - 0xc9
      12'hF6F: dout  = 8'b01000110; // 3951 :  70 - 0x46
      12'hF70: dout  = 8'b11010001; // 3952 : 209 - 0xd1 -- Background 0xee
      12'hF71: dout  = 8'b11011000; // 3953 : 216 - 0xd8
      12'hF72: dout  = 8'b11011000; // 3954 : 216 - 0xd8
      12'hF73: dout  = 8'b11011110; // 3955 : 222 - 0xde
      12'hF74: dout  = 8'b11010001; // 3956 : 209 - 0xd1
      12'hF75: dout  = 8'b11010000; // 3957 : 208 - 0xd0
      12'hF76: dout  = 8'b11011010; // 3958 : 218 - 0xda
      12'hF77: dout  = 8'b11011110; // 3959 : 222 - 0xde
      12'hF78: dout  = 8'b11011011; // 3960 : 219 - 0xdb -- Background 0xef
      12'hF79: dout  = 8'b11011001; // 3961 : 217 - 0xd9
      12'hF7A: dout  = 8'b11011011; // 3962 : 219 - 0xdb
      12'hF7B: dout  = 8'b11011100; // 3963 : 220 - 0xdc
      12'hF7C: dout  = 8'b11011011; // 3964 : 219 - 0xdb
      12'hF7D: dout  = 8'b11011111; // 3965 : 223 - 0xdf
      12'hF7E: dout  = 8'b00100000; // 3966 :  32 - 0x20
      12'hF7F: dout  = 8'b11100110; // 3967 : 230 - 0xe6
      12'hF80: dout  = 8'b11011010; // 3968 : 218 - 0xda -- Background 0xf0
      12'hF81: dout  = 8'b11011011; // 3969 : 219 - 0xdb
      12'hF82: dout  = 8'b11100000; // 3970 : 224 - 0xe0
      12'hF83: dout  = 8'b00100001; // 3971 :  33 - 0x21
      12'hF84: dout  = 8'b00000110; // 3972 :   6 - 0x6
      12'hF85: dout  = 8'b00001010; // 3973 :  10 - 0xa
      12'hF86: dout  = 8'b11010110; // 3974 : 214 - 0xd6
      12'hF87: dout  = 8'b11010111; // 3975 : 215 - 0xd7
      12'hF88: dout  = 8'b00100001; // 3976 :  33 - 0x21 -- Background 0xf1
      12'hF89: dout  = 8'b00100110; // 3977 :  38 - 0x26
      12'hF8A: dout  = 8'b00010100; // 3978 :  20 - 0x14
      12'hF8B: dout  = 8'b11010000; // 3979 : 208 - 0xd0
      12'hF8C: dout  = 8'b11101000; // 3980 : 232 - 0xe8
      12'hF8D: dout  = 8'b11010001; // 3981 : 209 - 0xd1
      12'hF8E: dout  = 8'b11010000; // 3982 : 208 - 0xd0
      12'hF8F: dout  = 8'b11010001; // 3983 : 209 - 0xd1
      12'hF90: dout  = 8'b11011110; // 3984 : 222 - 0xde -- Background 0xf2
      12'hF91: dout  = 8'b11010001; // 3985 : 209 - 0xd1
      12'hF92: dout  = 8'b11010000; // 3986 : 208 - 0xd0
      12'hF93: dout  = 8'b11010001; // 3987 : 209 - 0xd1
      12'hF94: dout  = 8'b11010000; // 3988 : 208 - 0xd0
      12'hF95: dout  = 8'b11010001; // 3989 : 209 - 0xd1
      12'hF96: dout  = 8'b00100110; // 3990 :  38 - 0x26
      12'hF97: dout  = 8'b00100001; // 3991 :  33 - 0x21
      12'hF98: dout  = 8'b01000010; // 3992 :  66 - 0x42 -- Background 0xf3
      12'hF99: dout  = 8'b11011011; // 3993 : 219 - 0xdb
      12'hF9A: dout  = 8'b11011011; // 3994 : 219 - 0xdb
      12'hF9B: dout  = 8'b01000010; // 3995 :  66 - 0x42
      12'hF9C: dout  = 8'b00100110; // 3996 :  38 - 0x26
      12'hF9D: dout  = 8'b11011011; // 3997 : 219 - 0xdb
      12'hF9E: dout  = 8'b01000010; // 3998 :  66 - 0x42
      12'hF9F: dout  = 8'b11011011; // 3999 : 219 - 0xdb
      12'hFA0: dout  = 8'b01000110; // 4000 :  70 - 0x46 -- Background 0xf4
      12'hFA1: dout  = 8'b11011011; // 4001 : 219 - 0xdb
      12'hFA2: dout  = 8'b00100001; // 4002 :  33 - 0x21
      12'hFA3: dout  = 8'b01101100; // 4003 : 108 - 0x6c
      12'hFA4: dout  = 8'b00001110; // 4004 :  14 - 0xe
      12'hFA5: dout  = 8'b11011111; // 4005 : 223 - 0xdf
      12'hFA6: dout  = 8'b11011011; // 4006 : 219 - 0xdb
      12'hFA7: dout  = 8'b11011011; // 4007 : 219 - 0xdb
      12'hFA8: dout  = 8'b11100100; // 4008 : 228 - 0xe4 -- Background 0xf5
      12'hFA9: dout  = 8'b11100101; // 4009 : 229 - 0xe5
      12'hFAA: dout  = 8'b00100110; // 4010 :  38 - 0x26
      12'hFAB: dout  = 8'b00100001; // 4011 :  33 - 0x21
      12'hFAC: dout  = 8'b10000110; // 4012 : 134 - 0x86
      12'hFAD: dout  = 8'b00010100; // 4013 :  20 - 0x14
      12'hFAE: dout  = 8'b11011011; // 4014 : 219 - 0xdb
      12'hFAF: dout  = 8'b11011011; // 4015 : 219 - 0xdb
      12'hFB0: dout  = 8'b00100110; // 4016 :  38 - 0x26 -- Background 0xf6
      12'hFB1: dout  = 8'b11011011; // 4017 : 219 - 0xdb
      12'hFB2: dout  = 8'b11100011; // 4018 : 227 - 0xe3
      12'hFB3: dout  = 8'b11011011; // 4019 : 219 - 0xdb
      12'hFB4: dout  = 8'b11100000; // 4020 : 224 - 0xe0
      12'hFB5: dout  = 8'b11011011; // 4021 : 219 - 0xdb
      12'hFB6: dout  = 8'b11011011; // 4022 : 219 - 0xdb
      12'hFB7: dout  = 8'b11100110; // 4023 : 230 - 0xe6
      12'hFB8: dout  = 8'b11011011; // 4024 : 219 - 0xdb -- Background 0xf7
      12'hFB9: dout  = 8'b01000010; // 4025 :  66 - 0x42
      12'hFBA: dout  = 8'b11011011; // 4026 : 219 - 0xdb
      12'hFBB: dout  = 8'b11011011; // 4027 : 219 - 0xdb
      12'hFBC: dout  = 8'b11011011; // 4028 : 219 - 0xdb
      12'hFBD: dout  = 8'b11010100; // 4029 : 212 - 0xd4
      12'hFBE: dout  = 8'b11011001; // 4030 : 217 - 0xd9
      12'hFBF: dout  = 8'b00100110; // 4031 :  38 - 0x26
      12'hFC0: dout  = 8'b11100111; // 4032 : 231 - 0xe7 -- Background 0xf8
      12'hFC1: dout  = 8'b00100001; // 4033 :  33 - 0x21
      12'hFC2: dout  = 8'b11000101; // 4034 : 197 - 0xc5
      12'hFC3: dout  = 8'b00010110; // 4035 :  22 - 0x16
      12'hFC4: dout  = 8'b01011111; // 4036 :  95 - 0x5f
      12'hFC5: dout  = 8'b10010101; // 4037 : 149 - 0x95
      12'hFC6: dout  = 8'b10010101; // 4038 : 149 - 0x95
      12'hFC7: dout  = 8'b10010101; // 4039 : 149 - 0x95
      12'hFC8: dout  = 8'b10010101; // 4040 : 149 - 0x95 -- Background 0xf9
      12'hFC9: dout  = 8'b10010110; // 4041 : 150 - 0x96
      12'hFCA: dout  = 8'b10010101; // 4042 : 149 - 0x95
      12'hFCB: dout  = 8'b10010101; // 4043 : 149 - 0x95
      12'hFCC: dout  = 8'b10010111; // 4044 : 151 - 0x97
      12'hFCD: dout  = 8'b10011000; // 4045 : 152 - 0x98
      12'hFCE: dout  = 8'b10010111; // 4046 : 151 - 0x97
      12'hFCF: dout  = 8'b10011000; // 4047 : 152 - 0x98
      12'hFD0: dout  = 8'b00001000; // 4048 :   8 - 0x8 -- Background 0xfa
      12'hFD1: dout  = 8'b00000101; // 4049 :   5 - 0x5
      12'hFD2: dout  = 8'b00100100; // 4050 :  36 - 0x24
      12'hFD3: dout  = 8'b00010111; // 4051 :  23 - 0x17
      12'hFD4: dout  = 8'b00010010; // 4052 :  18 - 0x12
      12'hFD5: dout  = 8'b00010111; // 4053 :  23 - 0x17
      12'hFD6: dout  = 8'b00011101; // 4054 :  29 - 0x1d
      12'hFD7: dout  = 8'b00001110; // 4055 :  14 - 0xe
      12'hFD8: dout  = 8'b00011001; // 4056 :  25 - 0x19 -- Background 0xfb
      12'hFD9: dout  = 8'b00010101; // 4057 :  21 - 0x15
      12'hFDA: dout  = 8'b00001010; // 4058 :  10 - 0xa
      12'hFDB: dout  = 8'b00100010; // 4059 :  34 - 0x22
      12'hFDC: dout  = 8'b00001110; // 4060 :  14 - 0xe
      12'hFDD: dout  = 8'b00011011; // 4061 :  27 - 0x1b
      12'hFDE: dout  = 8'b00100100; // 4062 :  36 - 0x24
      12'hFDF: dout  = 8'b00010000; // 4063 :  16 - 0x10
      12'hFE0: dout  = 8'b00011001; // 4064 :  25 - 0x19 -- Background 0xfc
      12'hFE1: dout  = 8'b00010101; // 4065 :  21 - 0x15
      12'hFE2: dout  = 8'b00001010; // 4066 :  10 - 0xa
      12'hFE3: dout  = 8'b00100010; // 4067 :  34 - 0x22
      12'hFE4: dout  = 8'b00001110; // 4068 :  14 - 0xe
      12'hFE5: dout  = 8'b00011011; // 4069 :  27 - 0x1b
      12'hFE6: dout  = 8'b00100100; // 4070 :  36 - 0x24
      12'hFE7: dout  = 8'b00010000; // 4071 :  16 - 0x10
      12'hFE8: dout  = 8'b00011001; // 4072 :  25 - 0x19 -- Background 0xfd
      12'hFE9: dout  = 8'b00101000; // 4073 :  40 - 0x28
      12'hFEA: dout  = 8'b00100010; // 4074 :  34 - 0x22
      12'hFEB: dout  = 8'b11110110; // 4075 : 246 - 0xf6
      12'hFEC: dout  = 8'b00000001; // 4076 :   1 - 0x1
      12'hFED: dout  = 8'b00000000; // 4077 :   0 - 0x0
      12'hFEE: dout  = 8'b00100011; // 4078 :  35 - 0x23
      12'hFEF: dout  = 8'b11001001; // 4079 : 201 - 0xc9
      12'hFF0: dout  = 8'b10101010; // 4080 : 170 - 0xaa -- Background 0xfe
      12'hFF1: dout  = 8'b00100011; // 4081 :  35 - 0x23
      12'hFF2: dout  = 8'b11101010; // 4082 : 234 - 0xea
      12'hFF3: dout  = 8'b00000100; // 4083 :   4 - 0x4
      12'hFF4: dout  = 8'b10011001; // 4084 : 153 - 0x99
      12'hFF5: dout  = 8'b10101010; // 4085 : 170 - 0xaa
      12'hFF6: dout  = 8'b10101010; // 4086 : 170 - 0xaa
      12'hFF7: dout  = 8'b10101010; // 4087 : 170 - 0xaa
      12'hFF8: dout  = 8'b11111111; // 4088 : 255 - 0xff -- Background 0xff
      12'hFF9: dout  = 8'b11111111; // 4089 : 255 - 0xff
      12'hFFA: dout  = 8'b11111111; // 4090 : 255 - 0xff
      12'hFFB: dout  = 8'b11111111; // 4091 : 255 - 0xff
      12'hFFC: dout  = 8'b11111111; // 4092 : 255 - 0xff
      12'hFFD: dout  = 8'b11111111; // 4093 : 255 - 0xff
      12'hFFE: dout  = 8'b11111111; // 4094 : 255 - 0xff
      12'hFFF: dout  = 8'b11111111; // 4095 : 255 - 0xff
    endcase
  end

endmodule
