---   Background Pattern table COLOR PLANE 1
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
--- Autcmatically generated VHDL ROM from a NES memory file----


---  Original memory dump file name: pacman_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_PACMAN_BG_PLN1 is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(11-1 downto 0);  --2048 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_PACMAN_BG_PLN1;

architecture BEHAVIORAL of ROM_PTABLE_PACMAN_BG_PLN1 is
  signal addr_int  : natural range 0 to 2**11-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Background pattern Table COLOR PLANE 1
    "00000000", --    0 -  0x0  :    0 - 0x0 -- Background 0x0
    "00000000", --    1 -  0x1  :    0 - 0x0
    "00000000", --    2 -  0x2  :    0 - 0x0
    "00000000", --    3 -  0x3  :    0 - 0x0
    "00000000", --    4 -  0x4  :    0 - 0x0
    "00000000", --    5 -  0x5  :    0 - 0x0
    "00000000", --    6 -  0x6  :    0 - 0x0
    "00000000", --    7 -  0x7  :    0 - 0x0
    "00000000", --    8 -  0x8  :    0 - 0x0 -- Background 0x1
    "00111000", --    9 -  0x9  :   56 - 0x38
    "01111100", --   10 -  0xa  :  124 - 0x7c
    "11111110", --   11 -  0xb  :  254 - 0xfe
    "11111110", --   12 -  0xc  :  254 - 0xfe
    "11111110", --   13 -  0xd  :  254 - 0xfe
    "01111100", --   14 -  0xe  :  124 - 0x7c
    "00111000", --   15 -  0xf  :   56 - 0x38
    "00000000", --   16 - 0x10  :    0 - 0x0 -- Background 0x2
    "00000000", --   17 - 0x11  :    0 - 0x0
    "00000000", --   18 - 0x12  :    0 - 0x0
    "00000000", --   19 - 0x13  :    0 - 0x0
    "00000000", --   20 - 0x14  :    0 - 0x0
    "00000000", --   21 - 0x15  :    0 - 0x0
    "00000000", --   22 - 0x16  :    0 - 0x0
    "00000000", --   23 - 0x17  :    0 - 0x0
    "00000000", --   24 - 0x18  :    0 - 0x0 -- Background 0x3
    "00000000", --   25 - 0x19  :    0 - 0x0
    "00000000", --   26 - 0x1a  :    0 - 0x0
    "00011000", --   27 - 0x1b  :   24 - 0x18
    "00011000", --   28 - 0x1c  :   24 - 0x18
    "00000000", --   29 - 0x1d  :    0 - 0x0
    "00000000", --   30 - 0x1e  :    0 - 0x0
    "00000000", --   31 - 0x1f  :    0 - 0x0
    "11111111", --   32 - 0x20  :  255 - 0xff -- Background 0x4
    "11111111", --   33 - 0x21  :  255 - 0xff
    "11111111", --   34 - 0x22  :  255 - 0xff
    "11111111", --   35 - 0x23  :  255 - 0xff
    "11111111", --   36 - 0x24  :  255 - 0xff
    "11111111", --   37 - 0x25  :  255 - 0xff
    "11111111", --   38 - 0x26  :  255 - 0xff
    "11111111", --   39 - 0x27  :  255 - 0xff
    "00001111", --   40 - 0x28  :   15 - 0xf -- Background 0x5
    "00001111", --   41 - 0x29  :   15 - 0xf
    "00001111", --   42 - 0x2a  :   15 - 0xf
    "00001111", --   43 - 0x2b  :   15 - 0xf
    "00001111", --   44 - 0x2c  :   15 - 0xf
    "00001111", --   45 - 0x2d  :   15 - 0xf
    "00001111", --   46 - 0x2e  :   15 - 0xf
    "00001111", --   47 - 0x2f  :   15 - 0xf
    "11110000", --   48 - 0x30  :  240 - 0xf0 -- Background 0x6
    "11110000", --   49 - 0x31  :  240 - 0xf0
    "11110000", --   50 - 0x32  :  240 - 0xf0
    "11110000", --   51 - 0x33  :  240 - 0xf0
    "11110000", --   52 - 0x34  :  240 - 0xf0
    "11110000", --   53 - 0x35  :  240 - 0xf0
    "11110000", --   54 - 0x36  :  240 - 0xf0
    "11110000", --   55 - 0x37  :  240 - 0xf0
    "00000000", --   56 - 0x38  :    0 - 0x0 -- Background 0x7
    "00000000", --   57 - 0x39  :    0 - 0x0
    "00000000", --   58 - 0x3a  :    0 - 0x0
    "00000000", --   59 - 0x3b  :    0 - 0x0
    "00000000", --   60 - 0x3c  :    0 - 0x0
    "00000000", --   61 - 0x3d  :    0 - 0x0
    "00000000", --   62 - 0x3e  :    0 - 0x0
    "00000000", --   63 - 0x3f  :    0 - 0x0
    "00000000", --   64 - 0x40  :    0 - 0x0 -- Background 0x8
    "00000000", --   65 - 0x41  :    0 - 0x0
    "00000000", --   66 - 0x42  :    0 - 0x0
    "00000000", --   67 - 0x43  :    0 - 0x0
    "00000000", --   68 - 0x44  :    0 - 0x0
    "00000000", --   69 - 0x45  :    0 - 0x0
    "00000000", --   70 - 0x46  :    0 - 0x0
    "00000000", --   71 - 0x47  :    0 - 0x0
    "00000000", --   72 - 0x48  :    0 - 0x0 -- Background 0x9
    "00000000", --   73 - 0x49  :    0 - 0x0
    "00000000", --   74 - 0x4a  :    0 - 0x0
    "00011000", --   75 - 0x4b  :   24 - 0x18
    "00011000", --   76 - 0x4c  :   24 - 0x18
    "00000000", --   77 - 0x4d  :    0 - 0x0
    "00000000", --   78 - 0x4e  :    0 - 0x0
    "00000000", --   79 - 0x4f  :    0 - 0x0
    "00000000", --   80 - 0x50  :    0 - 0x0 -- Background 0xa
    "00000000", --   81 - 0x51  :    0 - 0x0
    "00000000", --   82 - 0x52  :    0 - 0x0
    "00000000", --   83 - 0x53  :    0 - 0x0
    "00000000", --   84 - 0x54  :    0 - 0x0
    "00000000", --   85 - 0x55  :    0 - 0x0
    "00000000", --   86 - 0x56  :    0 - 0x0
    "00000000", --   87 - 0x57  :    0 - 0x0
    "00000000", --   88 - 0x58  :    0 - 0x0 -- Background 0xb
    "00000000", --   89 - 0x59  :    0 - 0x0
    "00000000", --   90 - 0x5a  :    0 - 0x0
    "00000000", --   91 - 0x5b  :    0 - 0x0
    "00000000", --   92 - 0x5c  :    0 - 0x0
    "00000000", --   93 - 0x5d  :    0 - 0x0
    "00000000", --   94 - 0x5e  :    0 - 0x0
    "00000000", --   95 - 0x5f  :    0 - 0x0
    "00000000", --   96 - 0x60  :    0 - 0x0 -- Background 0xc
    "00000000", --   97 - 0x61  :    0 - 0x0
    "00000000", --   98 - 0x62  :    0 - 0x0
    "00000000", --   99 - 0x63  :    0 - 0x0
    "00000000", --  100 - 0x64  :    0 - 0x0
    "00000000", --  101 - 0x65  :    0 - 0x0
    "00000000", --  102 - 0x66  :    0 - 0x0
    "00000000", --  103 - 0x67  :    0 - 0x0
    "00000000", --  104 - 0x68  :    0 - 0x0 -- Background 0xd
    "00000000", --  105 - 0x69  :    0 - 0x0
    "00000000", --  106 - 0x6a  :    0 - 0x0
    "00000000", --  107 - 0x6b  :    0 - 0x0
    "00000000", --  108 - 0x6c  :    0 - 0x0
    "00000000", --  109 - 0x6d  :    0 - 0x0
    "00000000", --  110 - 0x6e  :    0 - 0x0
    "00000000", --  111 - 0x6f  :    0 - 0x0
    "00000000", --  112 - 0x70  :    0 - 0x0 -- Background 0xe
    "00000000", --  113 - 0x71  :    0 - 0x0
    "00000000", --  114 - 0x72  :    0 - 0x0
    "00000000", --  115 - 0x73  :    0 - 0x0
    "00000000", --  116 - 0x74  :    0 - 0x0
    "00000000", --  117 - 0x75  :    0 - 0x0
    "00000000", --  118 - 0x76  :    0 - 0x0
    "00000000", --  119 - 0x77  :    0 - 0x0
    "00000000", --  120 - 0x78  :    0 - 0x0 -- Background 0xf
    "00000000", --  121 - 0x79  :    0 - 0x0
    "00000000", --  122 - 0x7a  :    0 - 0x0
    "00000000", --  123 - 0x7b  :    0 - 0x0
    "00000000", --  124 - 0x7c  :    0 - 0x0
    "00000000", --  125 - 0x7d  :    0 - 0x0
    "00000000", --  126 - 0x7e  :    0 - 0x0
    "00000000", --  127 - 0x7f  :    0 - 0x0
    "00000000", --  128 - 0x80  :    0 - 0x0 -- Background 0x10
    "00000000", --  129 - 0x81  :    0 - 0x0
    "00000000", --  130 - 0x82  :    0 - 0x0
    "00000000", --  131 - 0x83  :    0 - 0x0
    "00000000", --  132 - 0x84  :    0 - 0x0
    "00000000", --  133 - 0x85  :    0 - 0x0
    "00000000", --  134 - 0x86  :    0 - 0x0
    "00000000", --  135 - 0x87  :    0 - 0x0
    "00000000", --  136 - 0x88  :    0 - 0x0 -- Background 0x11
    "00000000", --  137 - 0x89  :    0 - 0x0
    "00000000", --  138 - 0x8a  :    0 - 0x0
    "00000000", --  139 - 0x8b  :    0 - 0x0
    "00000000", --  140 - 0x8c  :    0 - 0x0
    "00000000", --  141 - 0x8d  :    0 - 0x0
    "00000000", --  142 - 0x8e  :    0 - 0x0
    "00000000", --  143 - 0x8f  :    0 - 0x0
    "00000000", --  144 - 0x90  :    0 - 0x0 -- Background 0x12
    "00000000", --  145 - 0x91  :    0 - 0x0
    "00000000", --  146 - 0x92  :    0 - 0x0
    "00000000", --  147 - 0x93  :    0 - 0x0
    "00000000", --  148 - 0x94  :    0 - 0x0
    "00000000", --  149 - 0x95  :    0 - 0x0
    "00000000", --  150 - 0x96  :    0 - 0x0
    "00000000", --  151 - 0x97  :    0 - 0x0
    "00000000", --  152 - 0x98  :    0 - 0x0 -- Background 0x13
    "00000000", --  153 - 0x99  :    0 - 0x0
    "00000000", --  154 - 0x9a  :    0 - 0x0
    "00000000", --  155 - 0x9b  :    0 - 0x0
    "00000000", --  156 - 0x9c  :    0 - 0x0
    "00000000", --  157 - 0x9d  :    0 - 0x0
    "00000000", --  158 - 0x9e  :    0 - 0x0
    "00000000", --  159 - 0x9f  :    0 - 0x0
    "00000000", --  160 - 0xa0  :    0 - 0x0 -- Background 0x14
    "00000000", --  161 - 0xa1  :    0 - 0x0
    "00000000", --  162 - 0xa2  :    0 - 0x0
    "00000000", --  163 - 0xa3  :    0 - 0x0
    "00000000", --  164 - 0xa4  :    0 - 0x0
    "00000000", --  165 - 0xa5  :    0 - 0x0
    "00000000", --  166 - 0xa6  :    0 - 0x0
    "00000000", --  167 - 0xa7  :    0 - 0x0
    "00000000", --  168 - 0xa8  :    0 - 0x0 -- Background 0x15
    "00000000", --  169 - 0xa9  :    0 - 0x0
    "00000000", --  170 - 0xaa  :    0 - 0x0
    "00000000", --  171 - 0xab  :    0 - 0x0
    "00000000", --  172 - 0xac  :    0 - 0x0
    "00000000", --  173 - 0xad  :    0 - 0x0
    "00000000", --  174 - 0xae  :    0 - 0x0
    "00000000", --  175 - 0xaf  :    0 - 0x0
    "00000000", --  176 - 0xb0  :    0 - 0x0 -- Background 0x16
    "00000000", --  177 - 0xb1  :    0 - 0x0
    "00000000", --  178 - 0xb2  :    0 - 0x0
    "00000000", --  179 - 0xb3  :    0 - 0x0
    "00000000", --  180 - 0xb4  :    0 - 0x0
    "00000000", --  181 - 0xb5  :    0 - 0x0
    "00000000", --  182 - 0xb6  :    0 - 0x0
    "00000000", --  183 - 0xb7  :    0 - 0x0
    "00000000", --  184 - 0xb8  :    0 - 0x0 -- Background 0x17
    "00000000", --  185 - 0xb9  :    0 - 0x0
    "00000000", --  186 - 0xba  :    0 - 0x0
    "00000000", --  187 - 0xbb  :    0 - 0x0
    "00000000", --  188 - 0xbc  :    0 - 0x0
    "00000000", --  189 - 0xbd  :    0 - 0x0
    "00000000", --  190 - 0xbe  :    0 - 0x0
    "00000000", --  191 - 0xbf  :    0 - 0x0
    "00000000", --  192 - 0xc0  :    0 - 0x0 -- Background 0x18
    "00000000", --  193 - 0xc1  :    0 - 0x0
    "00000000", --  194 - 0xc2  :    0 - 0x0
    "00000000", --  195 - 0xc3  :    0 - 0x0
    "00000000", --  196 - 0xc4  :    0 - 0x0
    "00000000", --  197 - 0xc5  :    0 - 0x0
    "00000000", --  198 - 0xc6  :    0 - 0x0
    "00000000", --  199 - 0xc7  :    0 - 0x0
    "00000000", --  200 - 0xc8  :    0 - 0x0 -- Background 0x19
    "00000000", --  201 - 0xc9  :    0 - 0x0
    "00000000", --  202 - 0xca  :    0 - 0x0
    "00000000", --  203 - 0xcb  :    0 - 0x0
    "00000000", --  204 - 0xcc  :    0 - 0x0
    "00000000", --  205 - 0xcd  :    0 - 0x0
    "00000000", --  206 - 0xce  :    0 - 0x0
    "00000000", --  207 - 0xcf  :    0 - 0x0
    "00000000", --  208 - 0xd0  :    0 - 0x0 -- Background 0x1a
    "00000000", --  209 - 0xd1  :    0 - 0x0
    "00000000", --  210 - 0xd2  :    0 - 0x0
    "00000000", --  211 - 0xd3  :    0 - 0x0
    "00000000", --  212 - 0xd4  :    0 - 0x0
    "00000000", --  213 - 0xd5  :    0 - 0x0
    "00000000", --  214 - 0xd6  :    0 - 0x0
    "00000000", --  215 - 0xd7  :    0 - 0x0
    "00000000", --  216 - 0xd8  :    0 - 0x0 -- Background 0x1b
    "00000000", --  217 - 0xd9  :    0 - 0x0
    "00000000", --  218 - 0xda  :    0 - 0x0
    "00000000", --  219 - 0xdb  :    0 - 0x0
    "00000000", --  220 - 0xdc  :    0 - 0x0
    "00000000", --  221 - 0xdd  :    0 - 0x0
    "00000000", --  222 - 0xde  :    0 - 0x0
    "00000000", --  223 - 0xdf  :    0 - 0x0
    "00000000", --  224 - 0xe0  :    0 - 0x0 -- Background 0x1c
    "00000000", --  225 - 0xe1  :    0 - 0x0
    "00000000", --  226 - 0xe2  :    0 - 0x0
    "00000000", --  227 - 0xe3  :    0 - 0x0
    "00000000", --  228 - 0xe4  :    0 - 0x0
    "00000000", --  229 - 0xe5  :    0 - 0x0
    "00000000", --  230 - 0xe6  :    0 - 0x0
    "00000000", --  231 - 0xe7  :    0 - 0x0
    "00000000", --  232 - 0xe8  :    0 - 0x0 -- Background 0x1d
    "00000000", --  233 - 0xe9  :    0 - 0x0
    "00000000", --  234 - 0xea  :    0 - 0x0
    "00000000", --  235 - 0xeb  :    0 - 0x0
    "00000000", --  236 - 0xec  :    0 - 0x0
    "00000000", --  237 - 0xed  :    0 - 0x0
    "00000000", --  238 - 0xee  :    0 - 0x0
    "00000000", --  239 - 0xef  :    0 - 0x0
    "00000000", --  240 - 0xf0  :    0 - 0x0 -- Background 0x1e
    "00000000", --  241 - 0xf1  :    0 - 0x0
    "00000000", --  242 - 0xf2  :    0 - 0x0
    "00000000", --  243 - 0xf3  :    0 - 0x0
    "00000000", --  244 - 0xf4  :    0 - 0x0
    "00000000", --  245 - 0xf5  :    0 - 0x0
    "00000000", --  246 - 0xf6  :    0 - 0x0
    "00000000", --  247 - 0xf7  :    0 - 0x0
    "00000000", --  248 - 0xf8  :    0 - 0x0 -- Background 0x1f
    "00000000", --  249 - 0xf9  :    0 - 0x0
    "00000000", --  250 - 0xfa  :    0 - 0x0
    "00000000", --  251 - 0xfb  :    0 - 0x0
    "00000000", --  252 - 0xfc  :    0 - 0x0
    "00000000", --  253 - 0xfd  :    0 - 0x0
    "00000000", --  254 - 0xfe  :    0 - 0x0
    "00000000", --  255 - 0xff  :    0 - 0x0
    "00000000", --  256 - 0x100  :    0 - 0x0 -- Background 0x20
    "00000000", --  257 - 0x101  :    0 - 0x0
    "00000000", --  258 - 0x102  :    0 - 0x0
    "00000000", --  259 - 0x103  :    0 - 0x0
    "00000000", --  260 - 0x104  :    0 - 0x0
    "00000000", --  261 - 0x105  :    0 - 0x0
    "00000000", --  262 - 0x106  :    0 - 0x0
    "00000000", --  263 - 0x107  :    0 - 0x0
    "00001111", --  264 - 0x108  :   15 - 0xf -- Background 0x21
    "00001111", --  265 - 0x109  :   15 - 0xf
    "00001111", --  266 - 0x10a  :   15 - 0xf
    "00000111", --  267 - 0x10b  :    7 - 0x7
    "00000111", --  268 - 0x10c  :    7 - 0x7
    "00001111", --  269 - 0x10d  :   15 - 0xf
    "00001111", --  270 - 0x10e  :   15 - 0xf
    "00001111", --  271 - 0x10f  :   15 - 0xf
    "11110000", --  272 - 0x110  :  240 - 0xf0 -- Background 0x22
    "11110000", --  273 - 0x111  :  240 - 0xf0
    "11110000", --  274 - 0x112  :  240 - 0xf0
    "11100000", --  275 - 0x113  :  224 - 0xe0
    "11100000", --  276 - 0x114  :  224 - 0xe0
    "11110000", --  277 - 0x115  :  240 - 0xf0
    "11110000", --  278 - 0x116  :  240 - 0xf0
    "11110000", --  279 - 0x117  :  240 - 0xf0
    "11111111", --  280 - 0x118  :  255 - 0xff -- Background 0x23
    "11111111", --  281 - 0x119  :  255 - 0xff
    "11100001", --  282 - 0x11a  :  225 - 0xe1
    "11100001", --  283 - 0x11b  :  225 - 0xe1
    "11100001", --  284 - 0x11c  :  225 - 0xe1
    "11100001", --  285 - 0x11d  :  225 - 0xe1
    "11100001", --  286 - 0x11e  :  225 - 0xe1
    "11100001", --  287 - 0x11f  :  225 - 0xe1
    "10000111", --  288 - 0x120  :  135 - 0x87 -- Background 0x24
    "11000111", --  289 - 0x121  :  199 - 0xc7
    "11000000", --  290 - 0x122  :  192 - 0xc0
    "11000111", --  291 - 0x123  :  199 - 0xc7
    "11001111", --  292 - 0x124  :  207 - 0xcf
    "11001110", --  293 - 0x125  :  206 - 0xce
    "11001111", --  294 - 0x126  :  207 - 0xcf
    "11000111", --  295 - 0x127  :  199 - 0xc7
    "11111000", --  296 - 0x128  :  248 - 0xf8 -- Background 0x25
    "11111100", --  297 - 0x129  :  252 - 0xfc
    "00011100", --  298 - 0x12a  :   28 - 0x1c
    "11111100", --  299 - 0x12b  :  252 - 0xfc
    "11111100", --  300 - 0x12c  :  252 - 0xfc
    "00011100", --  301 - 0x12d  :   28 - 0x1c
    "11111100", --  302 - 0x12e  :  252 - 0xfc
    "11111100", --  303 - 0x12f  :  252 - 0xfc
    "11111111", --  304 - 0x130  :  255 - 0xff -- Background 0x26
    "11111111", --  305 - 0x131  :  255 - 0xff
    "11100111", --  306 - 0x132  :  231 - 0xe7
    "11100111", --  307 - 0x133  :  231 - 0xe7
    "11100111", --  308 - 0x134  :  231 - 0xe7
    "11100111", --  309 - 0x135  :  231 - 0xe7
    "11100111", --  310 - 0x136  :  231 - 0xe7
    "11100111", --  311 - 0x137  :  231 - 0xe7
    "11110000", --  312 - 0x138  :  240 - 0xf0 -- Background 0x27
    "11111001", --  313 - 0x139  :  249 - 0xf9
    "00111001", --  314 - 0x13a  :   57 - 0x39
    "00111001", --  315 - 0x13b  :   57 - 0x39
    "00111001", --  316 - 0x13c  :   57 - 0x39
    "00111001", --  317 - 0x13d  :   57 - 0x39
    "00111001", --  318 - 0x13e  :   57 - 0x39
    "00111000", --  319 - 0x13f  :   56 - 0x38
    "11111111", --  320 - 0x140  :  255 - 0xff -- Background 0x28
    "11111111", --  321 - 0x141  :  255 - 0xff
    "11000000", --  322 - 0x142  :  192 - 0xc0
    "11000000", --  323 - 0x143  :  192 - 0xc0
    "11000000", --  324 - 0x144  :  192 - 0xc0
    "11000000", --  325 - 0x145  :  192 - 0xc0
    "11111111", --  326 - 0x146  :  255 - 0xff
    "11111111", --  327 - 0x147  :  255 - 0xff
    "00011111", --  328 - 0x148  :   31 - 0x1f -- Background 0x29
    "00111111", --  329 - 0x149  :   63 - 0x3f
    "00110000", --  330 - 0x14a  :   48 - 0x30
    "00110000", --  331 - 0x14b  :   48 - 0x30
    "00110000", --  332 - 0x14c  :   48 - 0x30
    "00110000", --  333 - 0x14d  :   48 - 0x30
    "00111111", --  334 - 0x14e  :   63 - 0x3f
    "00011111", --  335 - 0x14f  :   31 - 0x1f
    "11100011", --  336 - 0x150  :  227 - 0xe3 -- Background 0x2a
    "11110011", --  337 - 0x151  :  243 - 0xf3
    "01110000", --  338 - 0x152  :  112 - 0x70
    "01110000", --  339 - 0x153  :  112 - 0x70
    "01110000", --  340 - 0x154  :  112 - 0x70
    "01110000", --  341 - 0x155  :  112 - 0x70
    "11110000", --  342 - 0x156  :  240 - 0xf0
    "11100000", --  343 - 0x157  :  224 - 0xe0
    "11111110", --  344 - 0x158  :  254 - 0xfe -- Background 0x2b
    "11111110", --  345 - 0x159  :  254 - 0xfe
    "01110000", --  346 - 0x15a  :  112 - 0x70
    "01110000", --  347 - 0x15b  :  112 - 0x70
    "01110000", --  348 - 0x15c  :  112 - 0x70
    "01110000", --  349 - 0x15d  :  112 - 0x70
    "01110000", --  350 - 0x15e  :  112 - 0x70
    "01110000", --  351 - 0x15f  :  112 - 0x70
    "00000000", --  352 - 0x160  :    0 - 0x0 -- Background 0x2c
    "00000000", --  353 - 0x161  :    0 - 0x0
    "00000000", --  354 - 0x162  :    0 - 0x0
    "00000000", --  355 - 0x163  :    0 - 0x0
    "00000000", --  356 - 0x164  :    0 - 0x0
    "00000000", --  357 - 0x165  :    0 - 0x0
    "00000000", --  358 - 0x166  :    0 - 0x0
    "00000000", --  359 - 0x167  :    0 - 0x0
    "11111111", --  360 - 0x168  :  255 - 0xff -- Background 0x2d
    "11111111", --  361 - 0x169  :  255 - 0xff
    "11111111", --  362 - 0x16a  :  255 - 0xff
    "11111111", --  363 - 0x16b  :  255 - 0xff
    "11111111", --  364 - 0x16c  :  255 - 0xff
    "11111111", --  365 - 0x16d  :  255 - 0xff
    "11111111", --  366 - 0x16e  :  255 - 0xff
    "11111111", --  367 - 0x16f  :  255 - 0xff
    "00000000", --  368 - 0x170  :    0 - 0x0 -- Background 0x2e
    "00000000", --  369 - 0x171  :    0 - 0x0
    "00000000", --  370 - 0x172  :    0 - 0x0
    "00000000", --  371 - 0x173  :    0 - 0x0
    "00000000", --  372 - 0x174  :    0 - 0x0
    "00000000", --  373 - 0x175  :    0 - 0x0
    "00000000", --  374 - 0x176  :    0 - 0x0
    "00000000", --  375 - 0x177  :    0 - 0x0
    "00000000", --  376 - 0x178  :    0 - 0x0 -- Background 0x2f
    "00000000", --  377 - 0x179  :    0 - 0x0
    "00000000", --  378 - 0x17a  :    0 - 0x0
    "00011000", --  379 - 0x17b  :   24 - 0x18
    "00011000", --  380 - 0x17c  :   24 - 0x18
    "00000000", --  381 - 0x17d  :    0 - 0x0
    "00000000", --  382 - 0x17e  :    0 - 0x0
    "00000000", --  383 - 0x17f  :    0 - 0x0
    "00000000", --  384 - 0x180  :    0 - 0x0 -- Background 0x30
    "00000000", --  385 - 0x181  :    0 - 0x0
    "00000000", --  386 - 0x182  :    0 - 0x0
    "00000000", --  387 - 0x183  :    0 - 0x0
    "00000000", --  388 - 0x184  :    0 - 0x0
    "00000000", --  389 - 0x185  :    0 - 0x0
    "00000000", --  390 - 0x186  :    0 - 0x0
    "00000000", --  391 - 0x187  :    0 - 0x0
    "00000000", --  392 - 0x188  :    0 - 0x0 -- Background 0x31
    "00000000", --  393 - 0x189  :    0 - 0x0
    "00000000", --  394 - 0x18a  :    0 - 0x0
    "00000000", --  395 - 0x18b  :    0 - 0x0
    "00000000", --  396 - 0x18c  :    0 - 0x0
    "00000000", --  397 - 0x18d  :    0 - 0x0
    "00000000", --  398 - 0x18e  :    0 - 0x0
    "00000000", --  399 - 0x18f  :    0 - 0x0
    "00000000", --  400 - 0x190  :    0 - 0x0 -- Background 0x32
    "00000000", --  401 - 0x191  :    0 - 0x0
    "00000000", --  402 - 0x192  :    0 - 0x0
    "00000000", --  403 - 0x193  :    0 - 0x0
    "00000000", --  404 - 0x194  :    0 - 0x0
    "00000000", --  405 - 0x195  :    0 - 0x0
    "00000000", --  406 - 0x196  :    0 - 0x0
    "00000000", --  407 - 0x197  :    0 - 0x0
    "00000000", --  408 - 0x198  :    0 - 0x0 -- Background 0x33
    "00000000", --  409 - 0x199  :    0 - 0x0
    "00000000", --  410 - 0x19a  :    0 - 0x0
    "00000000", --  411 - 0x19b  :    0 - 0x0
    "00000000", --  412 - 0x19c  :    0 - 0x0
    "00000000", --  413 - 0x19d  :    0 - 0x0
    "00000000", --  414 - 0x19e  :    0 - 0x0
    "00000000", --  415 - 0x19f  :    0 - 0x0
    "00000000", --  416 - 0x1a0  :    0 - 0x0 -- Background 0x34
    "00000000", --  417 - 0x1a1  :    0 - 0x0
    "00000000", --  418 - 0x1a2  :    0 - 0x0
    "00000000", --  419 - 0x1a3  :    0 - 0x0
    "00000000", --  420 - 0x1a4  :    0 - 0x0
    "00000000", --  421 - 0x1a5  :    0 - 0x0
    "00000000", --  422 - 0x1a6  :    0 - 0x0
    "00000000", --  423 - 0x1a7  :    0 - 0x0
    "00000000", --  424 - 0x1a8  :    0 - 0x0 -- Background 0x35
    "00000000", --  425 - 0x1a9  :    0 - 0x0
    "00000000", --  426 - 0x1aa  :    0 - 0x0
    "00000000", --  427 - 0x1ab  :    0 - 0x0
    "00000000", --  428 - 0x1ac  :    0 - 0x0
    "00000000", --  429 - 0x1ad  :    0 - 0x0
    "00000000", --  430 - 0x1ae  :    0 - 0x0
    "00000000", --  431 - 0x1af  :    0 - 0x0
    "00000000", --  432 - 0x1b0  :    0 - 0x0 -- Background 0x36
    "00000000", --  433 - 0x1b1  :    0 - 0x0
    "00000000", --  434 - 0x1b2  :    0 - 0x0
    "00000000", --  435 - 0x1b3  :    0 - 0x0
    "00000000", --  436 - 0x1b4  :    0 - 0x0
    "00000000", --  437 - 0x1b5  :    0 - 0x0
    "00000000", --  438 - 0x1b6  :    0 - 0x0
    "00000000", --  439 - 0x1b7  :    0 - 0x0
    "00000000", --  440 - 0x1b8  :    0 - 0x0 -- Background 0x37
    "00000000", --  441 - 0x1b9  :    0 - 0x0
    "00000000", --  442 - 0x1ba  :    0 - 0x0
    "00000000", --  443 - 0x1bb  :    0 - 0x0
    "00000000", --  444 - 0x1bc  :    0 - 0x0
    "00000000", --  445 - 0x1bd  :    0 - 0x0
    "00000000", --  446 - 0x1be  :    0 - 0x0
    "00000000", --  447 - 0x1bf  :    0 - 0x0
    "00000000", --  448 - 0x1c0  :    0 - 0x0 -- Background 0x38
    "00000000", --  449 - 0x1c1  :    0 - 0x0
    "00000000", --  450 - 0x1c2  :    0 - 0x0
    "00000000", --  451 - 0x1c3  :    0 - 0x0
    "00000000", --  452 - 0x1c4  :    0 - 0x0
    "00000000", --  453 - 0x1c5  :    0 - 0x0
    "00000000", --  454 - 0x1c6  :    0 - 0x0
    "00000000", --  455 - 0x1c7  :    0 - 0x0
    "00000000", --  456 - 0x1c8  :    0 - 0x0 -- Background 0x39
    "00000000", --  457 - 0x1c9  :    0 - 0x0
    "00000000", --  458 - 0x1ca  :    0 - 0x0
    "00000000", --  459 - 0x1cb  :    0 - 0x0
    "00000000", --  460 - 0x1cc  :    0 - 0x0
    "00000000", --  461 - 0x1cd  :    0 - 0x0
    "00000000", --  462 - 0x1ce  :    0 - 0x0
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "00000000", --  464 - 0x1d0  :    0 - 0x0 -- Background 0x3a
    "00000000", --  465 - 0x1d1  :    0 - 0x0
    "00000000", --  466 - 0x1d2  :    0 - 0x0
    "00000000", --  467 - 0x1d3  :    0 - 0x0
    "00000000", --  468 - 0x1d4  :    0 - 0x0
    "00000000", --  469 - 0x1d5  :    0 - 0x0
    "00000000", --  470 - 0x1d6  :    0 - 0x0
    "00000000", --  471 - 0x1d7  :    0 - 0x0
    "00000000", --  472 - 0x1d8  :    0 - 0x0 -- Background 0x3b
    "00000000", --  473 - 0x1d9  :    0 - 0x0
    "00000000", --  474 - 0x1da  :    0 - 0x0
    "00000000", --  475 - 0x1db  :    0 - 0x0
    "00000000", --  476 - 0x1dc  :    0 - 0x0
    "00000000", --  477 - 0x1dd  :    0 - 0x0
    "00000000", --  478 - 0x1de  :    0 - 0x0
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "00000000", --  480 - 0x1e0  :    0 - 0x0 -- Background 0x3c
    "00000111", --  481 - 0x1e1  :    7 - 0x7
    "00011111", --  482 - 0x1e2  :   31 - 0x1f
    "00111111", --  483 - 0x1e3  :   63 - 0x3f
    "00111111", --  484 - 0x1e4  :   63 - 0x3f
    "00001111", --  485 - 0x1e5  :   15 - 0xf
    "00000011", --  486 - 0x1e6  :    3 - 0x3
    "00000000", --  487 - 0x1e7  :    0 - 0x0
    "00000000", --  488 - 0x1e8  :    0 - 0x0 -- Background 0x3d
    "11000000", --  489 - 0x1e9  :  192 - 0xc0
    "11110000", --  490 - 0x1ea  :  240 - 0xf0
    "11111000", --  491 - 0x1eb  :  248 - 0xf8
    "11111000", --  492 - 0x1ec  :  248 - 0xf8
    "11111100", --  493 - 0x1ed  :  252 - 0xfc
    "11111100", --  494 - 0x1ee  :  252 - 0xfc
    "11111100", --  495 - 0x1ef  :  252 - 0xfc
    "00000000", --  496 - 0x1f0  :    0 - 0x0 -- Background 0x3e
    "00000011", --  497 - 0x1f1  :    3 - 0x3
    "00001111", --  498 - 0x1f2  :   15 - 0xf
    "00111111", --  499 - 0x1f3  :   63 - 0x3f
    "00111111", --  500 - 0x1f4  :   63 - 0x3f
    "00011111", --  501 - 0x1f5  :   31 - 0x1f
    "00000111", --  502 - 0x1f6  :    7 - 0x7
    "00000000", --  503 - 0x1f7  :    0 - 0x0
    "11111100", --  504 - 0x1f8  :  252 - 0xfc -- Background 0x3f
    "11111100", --  505 - 0x1f9  :  252 - 0xfc
    "11111100", --  506 - 0x1fa  :  252 - 0xfc
    "11111000", --  507 - 0x1fb  :  248 - 0xf8
    "11111000", --  508 - 0x1fc  :  248 - 0xf8
    "11110000", --  509 - 0x1fd  :  240 - 0xf0
    "11000000", --  510 - 0x1fe  :  192 - 0xc0
    "00000000", --  511 - 0x1ff  :    0 - 0x0
    "00000000", --  512 - 0x200  :    0 - 0x0 -- Background 0x40
    "00000000", --  513 - 0x201  :    0 - 0x0
    "00000000", --  514 - 0x202  :    0 - 0x0
    "00000000", --  515 - 0x203  :    0 - 0x0
    "00000000", --  516 - 0x204  :    0 - 0x0
    "00000000", --  517 - 0x205  :    0 - 0x0
    "00000000", --  518 - 0x206  :    0 - 0x0
    "00000000", --  519 - 0x207  :    0 - 0x0
    "00000000", --  520 - 0x208  :    0 - 0x0 -- Background 0x41
    "00000000", --  521 - 0x209  :    0 - 0x0
    "00000000", --  522 - 0x20a  :    0 - 0x0
    "00000000", --  523 - 0x20b  :    0 - 0x0
    "00000000", --  524 - 0x20c  :    0 - 0x0
    "00000000", --  525 - 0x20d  :    0 - 0x0
    "00000000", --  526 - 0x20e  :    0 - 0x0
    "00000000", --  527 - 0x20f  :    0 - 0x0
    "00000000", --  528 - 0x210  :    0 - 0x0 -- Background 0x42
    "00000000", --  529 - 0x211  :    0 - 0x0
    "00000000", --  530 - 0x212  :    0 - 0x0
    "00000000", --  531 - 0x213  :    0 - 0x0
    "00000000", --  532 - 0x214  :    0 - 0x0
    "00000000", --  533 - 0x215  :    0 - 0x0
    "00000000", --  534 - 0x216  :    0 - 0x0
    "00000000", --  535 - 0x217  :    0 - 0x0
    "00000000", --  536 - 0x218  :    0 - 0x0 -- Background 0x43
    "00000000", --  537 - 0x219  :    0 - 0x0
    "00000000", --  538 - 0x21a  :    0 - 0x0
    "00000000", --  539 - 0x21b  :    0 - 0x0
    "00000000", --  540 - 0x21c  :    0 - 0x0
    "00000000", --  541 - 0x21d  :    0 - 0x0
    "00000000", --  542 - 0x21e  :    0 - 0x0
    "00000000", --  543 - 0x21f  :    0 - 0x0
    "00000000", --  544 - 0x220  :    0 - 0x0 -- Background 0x44
    "00000000", --  545 - 0x221  :    0 - 0x0
    "00000000", --  546 - 0x222  :    0 - 0x0
    "00000000", --  547 - 0x223  :    0 - 0x0
    "00000000", --  548 - 0x224  :    0 - 0x0
    "00000000", --  549 - 0x225  :    0 - 0x0
    "00000000", --  550 - 0x226  :    0 - 0x0
    "00000000", --  551 - 0x227  :    0 - 0x0
    "00000000", --  552 - 0x228  :    0 - 0x0 -- Background 0x45
    "00000000", --  553 - 0x229  :    0 - 0x0
    "00000000", --  554 - 0x22a  :    0 - 0x0
    "00000000", --  555 - 0x22b  :    0 - 0x0
    "00000000", --  556 - 0x22c  :    0 - 0x0
    "00000000", --  557 - 0x22d  :    0 - 0x0
    "00000000", --  558 - 0x22e  :    0 - 0x0
    "00000000", --  559 - 0x22f  :    0 - 0x0
    "00000000", --  560 - 0x230  :    0 - 0x0 -- Background 0x46
    "00000000", --  561 - 0x231  :    0 - 0x0
    "00000000", --  562 - 0x232  :    0 - 0x0
    "00000000", --  563 - 0x233  :    0 - 0x0
    "00000000", --  564 - 0x234  :    0 - 0x0
    "00000000", --  565 - 0x235  :    0 - 0x0
    "00000000", --  566 - 0x236  :    0 - 0x0
    "00000000", --  567 - 0x237  :    0 - 0x0
    "00000000", --  568 - 0x238  :    0 - 0x0 -- Background 0x47
    "00000000", --  569 - 0x239  :    0 - 0x0
    "00000000", --  570 - 0x23a  :    0 - 0x0
    "00000000", --  571 - 0x23b  :    0 - 0x0
    "00000000", --  572 - 0x23c  :    0 - 0x0
    "00000000", --  573 - 0x23d  :    0 - 0x0
    "00000000", --  574 - 0x23e  :    0 - 0x0
    "00000000", --  575 - 0x23f  :    0 - 0x0
    "00000000", --  576 - 0x240  :    0 - 0x0 -- Background 0x48
    "00000000", --  577 - 0x241  :    0 - 0x0
    "00000000", --  578 - 0x242  :    0 - 0x0
    "00000000", --  579 - 0x243  :    0 - 0x0
    "00000000", --  580 - 0x244  :    0 - 0x0
    "00000000", --  581 - 0x245  :    0 - 0x0
    "00000000", --  582 - 0x246  :    0 - 0x0
    "00000000", --  583 - 0x247  :    0 - 0x0
    "00000000", --  584 - 0x248  :    0 - 0x0 -- Background 0x49
    "00000000", --  585 - 0x249  :    0 - 0x0
    "00000000", --  586 - 0x24a  :    0 - 0x0
    "00000000", --  587 - 0x24b  :    0 - 0x0
    "00000000", --  588 - 0x24c  :    0 - 0x0
    "00000000", --  589 - 0x24d  :    0 - 0x0
    "00000000", --  590 - 0x24e  :    0 - 0x0
    "00000000", --  591 - 0x24f  :    0 - 0x0
    "00000000", --  592 - 0x250  :    0 - 0x0 -- Background 0x4a
    "00000000", --  593 - 0x251  :    0 - 0x0
    "00000000", --  594 - 0x252  :    0 - 0x0
    "00000000", --  595 - 0x253  :    0 - 0x0
    "00000000", --  596 - 0x254  :    0 - 0x0
    "00000000", --  597 - 0x255  :    0 - 0x0
    "00000000", --  598 - 0x256  :    0 - 0x0
    "00000000", --  599 - 0x257  :    0 - 0x0
    "00000000", --  600 - 0x258  :    0 - 0x0 -- Background 0x4b
    "00000000", --  601 - 0x259  :    0 - 0x0
    "00000000", --  602 - 0x25a  :    0 - 0x0
    "00000000", --  603 - 0x25b  :    0 - 0x0
    "00000000", --  604 - 0x25c  :    0 - 0x0
    "00000000", --  605 - 0x25d  :    0 - 0x0
    "00000000", --  606 - 0x25e  :    0 - 0x0
    "00000000", --  607 - 0x25f  :    0 - 0x0
    "00000000", --  608 - 0x260  :    0 - 0x0 -- Background 0x4c
    "00000000", --  609 - 0x261  :    0 - 0x0
    "00000000", --  610 - 0x262  :    0 - 0x0
    "00000000", --  611 - 0x263  :    0 - 0x0
    "00000000", --  612 - 0x264  :    0 - 0x0
    "00000000", --  613 - 0x265  :    0 - 0x0
    "00000000", --  614 - 0x266  :    0 - 0x0
    "00000000", --  615 - 0x267  :    0 - 0x0
    "00000000", --  616 - 0x268  :    0 - 0x0 -- Background 0x4d
    "00000000", --  617 - 0x269  :    0 - 0x0
    "00000000", --  618 - 0x26a  :    0 - 0x0
    "00000000", --  619 - 0x26b  :    0 - 0x0
    "00000000", --  620 - 0x26c  :    0 - 0x0
    "00000000", --  621 - 0x26d  :    0 - 0x0
    "00000000", --  622 - 0x26e  :    0 - 0x0
    "00000000", --  623 - 0x26f  :    0 - 0x0
    "00000000", --  624 - 0x270  :    0 - 0x0 -- Background 0x4e
    "00000000", --  625 - 0x271  :    0 - 0x0
    "00000000", --  626 - 0x272  :    0 - 0x0
    "00000000", --  627 - 0x273  :    0 - 0x0
    "00000000", --  628 - 0x274  :    0 - 0x0
    "00000000", --  629 - 0x275  :    0 - 0x0
    "00000000", --  630 - 0x276  :    0 - 0x0
    "00000000", --  631 - 0x277  :    0 - 0x0
    "00000000", --  632 - 0x278  :    0 - 0x0 -- Background 0x4f
    "00000000", --  633 - 0x279  :    0 - 0x0
    "00000000", --  634 - 0x27a  :    0 - 0x0
    "00000000", --  635 - 0x27b  :    0 - 0x0
    "00000000", --  636 - 0x27c  :    0 - 0x0
    "00000000", --  637 - 0x27d  :    0 - 0x0
    "00000000", --  638 - 0x27e  :    0 - 0x0
    "00000000", --  639 - 0x27f  :    0 - 0x0
    "00000000", --  640 - 0x280  :    0 - 0x0 -- Background 0x50
    "00000000", --  641 - 0x281  :    0 - 0x0
    "00000000", --  642 - 0x282  :    0 - 0x0
    "00000000", --  643 - 0x283  :    0 - 0x0
    "00000000", --  644 - 0x284  :    0 - 0x0
    "00000000", --  645 - 0x285  :    0 - 0x0
    "00000000", --  646 - 0x286  :    0 - 0x0
    "00000000", --  647 - 0x287  :    0 - 0x0
    "00000000", --  648 - 0x288  :    0 - 0x0 -- Background 0x51
    "00000000", --  649 - 0x289  :    0 - 0x0
    "00000000", --  650 - 0x28a  :    0 - 0x0
    "00000000", --  651 - 0x28b  :    0 - 0x0
    "00000000", --  652 - 0x28c  :    0 - 0x0
    "00000000", --  653 - 0x28d  :    0 - 0x0
    "00000000", --  654 - 0x28e  :    0 - 0x0
    "00000000", --  655 - 0x28f  :    0 - 0x0
    "00000000", --  656 - 0x290  :    0 - 0x0 -- Background 0x52
    "00000000", --  657 - 0x291  :    0 - 0x0
    "00000000", --  658 - 0x292  :    0 - 0x0
    "00000000", --  659 - 0x293  :    0 - 0x0
    "00000000", --  660 - 0x294  :    0 - 0x0
    "00000000", --  661 - 0x295  :    0 - 0x0
    "00000000", --  662 - 0x296  :    0 - 0x0
    "00000000", --  663 - 0x297  :    0 - 0x0
    "00000000", --  664 - 0x298  :    0 - 0x0 -- Background 0x53
    "00000000", --  665 - 0x299  :    0 - 0x0
    "00000000", --  666 - 0x29a  :    0 - 0x0
    "00000000", --  667 - 0x29b  :    0 - 0x0
    "00000000", --  668 - 0x29c  :    0 - 0x0
    "00000000", --  669 - 0x29d  :    0 - 0x0
    "00000000", --  670 - 0x29e  :    0 - 0x0
    "00000000", --  671 - 0x29f  :    0 - 0x0
    "00000000", --  672 - 0x2a0  :    0 - 0x0 -- Background 0x54
    "00000000", --  673 - 0x2a1  :    0 - 0x0
    "00000000", --  674 - 0x2a2  :    0 - 0x0
    "00000000", --  675 - 0x2a3  :    0 - 0x0
    "00000000", --  676 - 0x2a4  :    0 - 0x0
    "00000000", --  677 - 0x2a5  :    0 - 0x0
    "00000000", --  678 - 0x2a6  :    0 - 0x0
    "00000000", --  679 - 0x2a7  :    0 - 0x0
    "00000000", --  680 - 0x2a8  :    0 - 0x0 -- Background 0x55
    "00000000", --  681 - 0x2a9  :    0 - 0x0
    "00000000", --  682 - 0x2aa  :    0 - 0x0
    "00000000", --  683 - 0x2ab  :    0 - 0x0
    "00000000", --  684 - 0x2ac  :    0 - 0x0
    "00000000", --  685 - 0x2ad  :    0 - 0x0
    "00000000", --  686 - 0x2ae  :    0 - 0x0
    "00000000", --  687 - 0x2af  :    0 - 0x0
    "00000000", --  688 - 0x2b0  :    0 - 0x0 -- Background 0x56
    "00000000", --  689 - 0x2b1  :    0 - 0x0
    "00000000", --  690 - 0x2b2  :    0 - 0x0
    "00000000", --  691 - 0x2b3  :    0 - 0x0
    "00000000", --  692 - 0x2b4  :    0 - 0x0
    "00000000", --  693 - 0x2b5  :    0 - 0x0
    "00000000", --  694 - 0x2b6  :    0 - 0x0
    "00000000", --  695 - 0x2b7  :    0 - 0x0
    "00000000", --  696 - 0x2b8  :    0 - 0x0 -- Background 0x57
    "00000000", --  697 - 0x2b9  :    0 - 0x0
    "00000000", --  698 - 0x2ba  :    0 - 0x0
    "00000000", --  699 - 0x2bb  :    0 - 0x0
    "00000000", --  700 - 0x2bc  :    0 - 0x0
    "00000000", --  701 - 0x2bd  :    0 - 0x0
    "00000000", --  702 - 0x2be  :    0 - 0x0
    "00000000", --  703 - 0x2bf  :    0 - 0x0
    "00000000", --  704 - 0x2c0  :    0 - 0x0 -- Background 0x58
    "00000000", --  705 - 0x2c1  :    0 - 0x0
    "00000000", --  706 - 0x2c2  :    0 - 0x0
    "00000000", --  707 - 0x2c3  :    0 - 0x0
    "00000000", --  708 - 0x2c4  :    0 - 0x0
    "00000000", --  709 - 0x2c5  :    0 - 0x0
    "00000000", --  710 - 0x2c6  :    0 - 0x0
    "00000000", --  711 - 0x2c7  :    0 - 0x0
    "00000000", --  712 - 0x2c8  :    0 - 0x0 -- Background 0x59
    "00000000", --  713 - 0x2c9  :    0 - 0x0
    "00000000", --  714 - 0x2ca  :    0 - 0x0
    "00000000", --  715 - 0x2cb  :    0 - 0x0
    "00000000", --  716 - 0x2cc  :    0 - 0x0
    "00000000", --  717 - 0x2cd  :    0 - 0x0
    "00000000", --  718 - 0x2ce  :    0 - 0x0
    "00000000", --  719 - 0x2cf  :    0 - 0x0
    "00000000", --  720 - 0x2d0  :    0 - 0x0 -- Background 0x5a
    "00000000", --  721 - 0x2d1  :    0 - 0x0
    "00000000", --  722 - 0x2d2  :    0 - 0x0
    "00000000", --  723 - 0x2d3  :    0 - 0x0
    "00000000", --  724 - 0x2d4  :    0 - 0x0
    "00000000", --  725 - 0x2d5  :    0 - 0x0
    "00000000", --  726 - 0x2d6  :    0 - 0x0
    "00000000", --  727 - 0x2d7  :    0 - 0x0
    "00000000", --  728 - 0x2d8  :    0 - 0x0 -- Background 0x5b
    "00000000", --  729 - 0x2d9  :    0 - 0x0
    "00000000", --  730 - 0x2da  :    0 - 0x0
    "00000000", --  731 - 0x2db  :    0 - 0x0
    "00000000", --  732 - 0x2dc  :    0 - 0x0
    "00000000", --  733 - 0x2dd  :    0 - 0x0
    "00000000", --  734 - 0x2de  :    0 - 0x0
    "00000000", --  735 - 0x2df  :    0 - 0x0
    "00000000", --  736 - 0x2e0  :    0 - 0x0 -- Background 0x5c
    "00000000", --  737 - 0x2e1  :    0 - 0x0
    "00000000", --  738 - 0x2e2  :    0 - 0x0
    "00000000", --  739 - 0x2e3  :    0 - 0x0
    "00000000", --  740 - 0x2e4  :    0 - 0x0
    "00000000", --  741 - 0x2e5  :    0 - 0x0
    "00000000", --  742 - 0x2e6  :    0 - 0x0
    "00000000", --  743 - 0x2e7  :    0 - 0x0
    "00000000", --  744 - 0x2e8  :    0 - 0x0 -- Background 0x5d
    "00000000", --  745 - 0x2e9  :    0 - 0x0
    "00000000", --  746 - 0x2ea  :    0 - 0x0
    "00000000", --  747 - 0x2eb  :    0 - 0x0
    "00000000", --  748 - 0x2ec  :    0 - 0x0
    "00000000", --  749 - 0x2ed  :    0 - 0x0
    "00000000", --  750 - 0x2ee  :    0 - 0x0
    "00000000", --  751 - 0x2ef  :    0 - 0x0
    "00000000", --  752 - 0x2f0  :    0 - 0x0 -- Background 0x5e
    "00000000", --  753 - 0x2f1  :    0 - 0x0
    "00010000", --  754 - 0x2f2  :   16 - 0x10
    "00010000", --  755 - 0x2f3  :   16 - 0x10
    "00010000", --  756 - 0x2f4  :   16 - 0x10
    "00010000", --  757 - 0x2f5  :   16 - 0x10
    "00000000", --  758 - 0x2f6  :    0 - 0x0
    "00000000", --  759 - 0x2f7  :    0 - 0x0
    "00000000", --  760 - 0x2f8  :    0 - 0x0 -- Background 0x5f
    "00000000", --  761 - 0x2f9  :    0 - 0x0
    "00000000", --  762 - 0x2fa  :    0 - 0x0
    "00000000", --  763 - 0x2fb  :    0 - 0x0
    "00000000", --  764 - 0x2fc  :    0 - 0x0
    "00000000", --  765 - 0x2fd  :    0 - 0x0
    "00000000", --  766 - 0x2fe  :    0 - 0x0
    "00000000", --  767 - 0x2ff  :    0 - 0x0
    "00000000", --  768 - 0x300  :    0 - 0x0 -- Background 0x60
    "00000000", --  769 - 0x301  :    0 - 0x0
    "00000000", --  770 - 0x302  :    0 - 0x0
    "00000000", --  771 - 0x303  :    0 - 0x0
    "00000000", --  772 - 0x304  :    0 - 0x0
    "00000000", --  773 - 0x305  :    0 - 0x0
    "00000000", --  774 - 0x306  :    0 - 0x0
    "00000000", --  775 - 0x307  :    0 - 0x0
    "00000000", --  776 - 0x308  :    0 - 0x0 -- Background 0x61
    "00000000", --  777 - 0x309  :    0 - 0x0
    "00000000", --  778 - 0x30a  :    0 - 0x0
    "00000000", --  779 - 0x30b  :    0 - 0x0
    "00000000", --  780 - 0x30c  :    0 - 0x0
    "00000000", --  781 - 0x30d  :    0 - 0x0
    "00000000", --  782 - 0x30e  :    0 - 0x0
    "00000000", --  783 - 0x30f  :    0 - 0x0
    "00000000", --  784 - 0x310  :    0 - 0x0 -- Background 0x62
    "00000000", --  785 - 0x311  :    0 - 0x0
    "00000000", --  786 - 0x312  :    0 - 0x0
    "00000000", --  787 - 0x313  :    0 - 0x0
    "00000000", --  788 - 0x314  :    0 - 0x0
    "00000000", --  789 - 0x315  :    0 - 0x0
    "00000000", --  790 - 0x316  :    0 - 0x0
    "00000000", --  791 - 0x317  :    0 - 0x0
    "00000000", --  792 - 0x318  :    0 - 0x0 -- Background 0x63
    "00000000", --  793 - 0x319  :    0 - 0x0
    "00000000", --  794 - 0x31a  :    0 - 0x0
    "00000000", --  795 - 0x31b  :    0 - 0x0
    "00000000", --  796 - 0x31c  :    0 - 0x0
    "00000000", --  797 - 0x31d  :    0 - 0x0
    "00000000", --  798 - 0x31e  :    0 - 0x0
    "00000000", --  799 - 0x31f  :    0 - 0x0
    "00000000", --  800 - 0x320  :    0 - 0x0 -- Background 0x64
    "00000000", --  801 - 0x321  :    0 - 0x0
    "00000000", --  802 - 0x322  :    0 - 0x0
    "00000000", --  803 - 0x323  :    0 - 0x0
    "00000000", --  804 - 0x324  :    0 - 0x0
    "00000000", --  805 - 0x325  :    0 - 0x0
    "00000000", --  806 - 0x326  :    0 - 0x0
    "00000000", --  807 - 0x327  :    0 - 0x0
    "00000000", --  808 - 0x328  :    0 - 0x0 -- Background 0x65
    "00000000", --  809 - 0x329  :    0 - 0x0
    "00000000", --  810 - 0x32a  :    0 - 0x0
    "00000000", --  811 - 0x32b  :    0 - 0x0
    "00000000", --  812 - 0x32c  :    0 - 0x0
    "00000000", --  813 - 0x32d  :    0 - 0x0
    "00000000", --  814 - 0x32e  :    0 - 0x0
    "00000000", --  815 - 0x32f  :    0 - 0x0
    "00000000", --  816 - 0x330  :    0 - 0x0 -- Background 0x66
    "00000000", --  817 - 0x331  :    0 - 0x0
    "00000000", --  818 - 0x332  :    0 - 0x0
    "00000000", --  819 - 0x333  :    0 - 0x0
    "00000000", --  820 - 0x334  :    0 - 0x0
    "00000000", --  821 - 0x335  :    0 - 0x0
    "00000000", --  822 - 0x336  :    0 - 0x0
    "00000000", --  823 - 0x337  :    0 - 0x0
    "00000000", --  824 - 0x338  :    0 - 0x0 -- Background 0x67
    "00000000", --  825 - 0x339  :    0 - 0x0
    "00000000", --  826 - 0x33a  :    0 - 0x0
    "00000000", --  827 - 0x33b  :    0 - 0x0
    "00000000", --  828 - 0x33c  :    0 - 0x0
    "00000000", --  829 - 0x33d  :    0 - 0x0
    "00000000", --  830 - 0x33e  :    0 - 0x0
    "00000000", --  831 - 0x33f  :    0 - 0x0
    "00000000", --  832 - 0x340  :    0 - 0x0 -- Background 0x68
    "00000000", --  833 - 0x341  :    0 - 0x0
    "00000000", --  834 - 0x342  :    0 - 0x0
    "00000001", --  835 - 0x343  :    1 - 0x1
    "00000001", --  836 - 0x344  :    1 - 0x1
    "00001011", --  837 - 0x345  :   11 - 0xb
    "00011100", --  838 - 0x346  :   28 - 0x1c
    "00111111", --  839 - 0x347  :   63 - 0x3f
    "00000000", --  840 - 0x348  :    0 - 0x0 -- Background 0x69
    "00000000", --  841 - 0x349  :    0 - 0x0
    "00110000", --  842 - 0x34a  :   48 - 0x30
    "01111000", --  843 - 0x34b  :  120 - 0x78
    "10000000", --  844 - 0x34c  :  128 - 0x80
    "11110000", --  845 - 0x34d  :  240 - 0xf0
    "11111000", --  846 - 0x34e  :  248 - 0xf8
    "11111100", --  847 - 0x34f  :  252 - 0xfc
    "00111111", --  848 - 0x350  :   63 - 0x3f -- Background 0x6a
    "00111111", --  849 - 0x351  :   63 - 0x3f
    "00111111", --  850 - 0x352  :   63 - 0x3f
    "00011111", --  851 - 0x353  :   31 - 0x1f
    "00011111", --  852 - 0x354  :   31 - 0x1f
    "00000111", --  853 - 0x355  :    7 - 0x7
    "00000000", --  854 - 0x356  :    0 - 0x0
    "00000000", --  855 - 0x357  :    0 - 0x0
    "11111100", --  856 - 0x358  :  252 - 0xfc -- Background 0x6b
    "11101100", --  857 - 0x359  :  236 - 0xec
    "11101100", --  858 - 0x35a  :  236 - 0xec
    "11011000", --  859 - 0x35b  :  216 - 0xd8
    "11111000", --  860 - 0x35c  :  248 - 0xf8
    "11100000", --  861 - 0x35d  :  224 - 0xe0
    "00000000", --  862 - 0x35e  :    0 - 0x0
    "00000000", --  863 - 0x35f  :    0 - 0x0
    "00000000", --  864 - 0x360  :    0 - 0x0 -- Background 0x6c
    "00000000", --  865 - 0x361  :    0 - 0x0
    "00000001", --  866 - 0x362  :    1 - 0x1
    "00011101", --  867 - 0x363  :   29 - 0x1d
    "00111110", --  868 - 0x364  :   62 - 0x3e
    "00111111", --  869 - 0x365  :   63 - 0x3f
    "00111111", --  870 - 0x366  :   63 - 0x3f
    "00111111", --  871 - 0x367  :   63 - 0x3f
    "00000000", --  872 - 0x368  :    0 - 0x0 -- Background 0x6d
    "10000000", --  873 - 0x369  :  128 - 0x80
    "00000000", --  874 - 0x36a  :    0 - 0x0
    "01110000", --  875 - 0x36b  :  112 - 0x70
    "11111000", --  876 - 0x36c  :  248 - 0xf8
    "11111100", --  877 - 0x36d  :  252 - 0xfc
    "11111100", --  878 - 0x36e  :  252 - 0xfc
    "11111100", --  879 - 0x36f  :  252 - 0xfc
    "00111111", --  880 - 0x370  :   63 - 0x3f -- Background 0x6e
    "00111111", --  881 - 0x371  :   63 - 0x3f
    "00011111", --  882 - 0x372  :   31 - 0x1f
    "00011111", --  883 - 0x373  :   31 - 0x1f
    "00001111", --  884 - 0x374  :   15 - 0xf
    "00000110", --  885 - 0x375  :    6 - 0x6
    "00000000", --  886 - 0x376  :    0 - 0x0
    "00000000", --  887 - 0x377  :    0 - 0x0
    "11101100", --  888 - 0x378  :  236 - 0xec -- Background 0x6f
    "11101100", --  889 - 0x379  :  236 - 0xec
    "11011000", --  890 - 0x37a  :  216 - 0xd8
    "11111000", --  891 - 0x37b  :  248 - 0xf8
    "11110000", --  892 - 0x37c  :  240 - 0xf0
    "11100000", --  893 - 0x37d  :  224 - 0xe0
    "00000000", --  894 - 0x37e  :    0 - 0x0
    "00000000", --  895 - 0x37f  :    0 - 0x0
    "00000000", --  896 - 0x380  :    0 - 0x0 -- Background 0x70
    "00000000", --  897 - 0x381  :    0 - 0x0
    "00000000", --  898 - 0x382  :    0 - 0x0
    "00000000", --  899 - 0x383  :    0 - 0x0
    "00000000", --  900 - 0x384  :    0 - 0x0
    "00000000", --  901 - 0x385  :    0 - 0x0
    "00000000", --  902 - 0x386  :    0 - 0x0
    "00000000", --  903 - 0x387  :    0 - 0x0
    "00000000", --  904 - 0x388  :    0 - 0x0 -- Background 0x71
    "00000000", --  905 - 0x389  :    0 - 0x0
    "00000000", --  906 - 0x38a  :    0 - 0x0
    "00000000", --  907 - 0x38b  :    0 - 0x0
    "00000000", --  908 - 0x38c  :    0 - 0x0
    "00000000", --  909 - 0x38d  :    0 - 0x0
    "00000000", --  910 - 0x38e  :    0 - 0x0
    "00000000", --  911 - 0x38f  :    0 - 0x0
    "00000000", --  912 - 0x390  :    0 - 0x0 -- Background 0x72
    "00000000", --  913 - 0x391  :    0 - 0x0
    "00000000", --  914 - 0x392  :    0 - 0x0
    "00000000", --  915 - 0x393  :    0 - 0x0
    "00000000", --  916 - 0x394  :    0 - 0x0
    "00000000", --  917 - 0x395  :    0 - 0x0
    "00000000", --  918 - 0x396  :    0 - 0x0
    "00000000", --  919 - 0x397  :    0 - 0x0
    "00000000", --  920 - 0x398  :    0 - 0x0 -- Background 0x73
    "00000000", --  921 - 0x399  :    0 - 0x0
    "00000000", --  922 - 0x39a  :    0 - 0x0
    "00000000", --  923 - 0x39b  :    0 - 0x0
    "00000000", --  924 - 0x39c  :    0 - 0x0
    "00000000", --  925 - 0x39d  :    0 - 0x0
    "00000000", --  926 - 0x39e  :    0 - 0x0
    "00000000", --  927 - 0x39f  :    0 - 0x0
    "00000000", --  928 - 0x3a0  :    0 - 0x0 -- Background 0x74
    "00000000", --  929 - 0x3a1  :    0 - 0x0
    "00000000", --  930 - 0x3a2  :    0 - 0x0
    "00000000", --  931 - 0x3a3  :    0 - 0x0
    "00010001", --  932 - 0x3a4  :   17 - 0x11
    "00010011", --  933 - 0x3a5  :   19 - 0x13
    "00011111", --  934 - 0x3a6  :   31 - 0x1f
    "00011111", --  935 - 0x3a7  :   31 - 0x1f
    "00000000", --  936 - 0x3a8  :    0 - 0x0 -- Background 0x75
    "00000000", --  937 - 0x3a9  :    0 - 0x0
    "00000000", --  938 - 0x3aa  :    0 - 0x0
    "10000000", --  939 - 0x3ab  :  128 - 0x80
    "11000100", --  940 - 0x3ac  :  196 - 0xc4
    "11100100", --  941 - 0x3ad  :  228 - 0xe4
    "11111100", --  942 - 0x3ae  :  252 - 0xfc
    "11111100", --  943 - 0x3af  :  252 - 0xfc
    "00011111", --  944 - 0x3b0  :   31 - 0x1f -- Background 0x76
    "00001110", --  945 - 0x3b1  :   14 - 0xe
    "00000110", --  946 - 0x3b2  :    6 - 0x6
    "00000010", --  947 - 0x3b3  :    2 - 0x2
    "00000000", --  948 - 0x3b4  :    0 - 0x0
    "00000000", --  949 - 0x3b5  :    0 - 0x0
    "00000000", --  950 - 0x3b6  :    0 - 0x0
    "00000000", --  951 - 0x3b7  :    0 - 0x0
    "11111100", --  952 - 0x3b8  :  252 - 0xfc -- Background 0x77
    "10111000", --  953 - 0x3b9  :  184 - 0xb8
    "10110000", --  954 - 0x3ba  :  176 - 0xb0
    "10100000", --  955 - 0x3bb  :  160 - 0xa0
    "10000000", --  956 - 0x3bc  :  128 - 0x80
    "00000000", --  957 - 0x3bd  :    0 - 0x0
    "00000000", --  958 - 0x3be  :    0 - 0x0
    "00000000", --  959 - 0x3bf  :    0 - 0x0
    "00000000", --  960 - 0x3c0  :    0 - 0x0 -- Background 0x78
    "00000000", --  961 - 0x3c1  :    0 - 0x0
    "00000000", --  962 - 0x3c2  :    0 - 0x0
    "00000001", --  963 - 0x3c3  :    1 - 0x1
    "00000011", --  964 - 0x3c4  :    3 - 0x3
    "00000110", --  965 - 0x3c5  :    6 - 0x6
    "00000110", --  966 - 0x3c6  :    6 - 0x6
    "00001111", --  967 - 0x3c7  :   15 - 0xf
    "00000000", --  968 - 0x3c8  :    0 - 0x0 -- Background 0x79
    "00011000", --  969 - 0x3c9  :   24 - 0x18
    "11110100", --  970 - 0x3ca  :  244 - 0xf4
    "11111000", --  971 - 0x3cb  :  248 - 0xf8
    "00111000", --  972 - 0x3cc  :   56 - 0x38
    "01111100", --  973 - 0x3cd  :  124 - 0x7c
    "11111100", --  974 - 0x3ce  :  252 - 0xfc
    "11111100", --  975 - 0x3cf  :  252 - 0xfc
    "00001111", --  976 - 0x3d0  :   15 - 0xf -- Background 0x7a
    "00011111", --  977 - 0x3d1  :   31 - 0x1f
    "00110000", --  978 - 0x3d2  :   48 - 0x30
    "00111000", --  979 - 0x3d3  :   56 - 0x38
    "00011101", --  980 - 0x3d4  :   29 - 0x1d
    "00000011", --  981 - 0x3d5  :    3 - 0x3
    "00000011", --  982 - 0x3d6  :    3 - 0x3
    "00000000", --  983 - 0x3d7  :    0 - 0x0
    "11111100", --  984 - 0x3d8  :  252 - 0xfc -- Background 0x7b
    "11111100", --  985 - 0x3d9  :  252 - 0xfc
    "01111100", --  986 - 0x3da  :  124 - 0x7c
    "10001110", --  987 - 0x3db  :  142 - 0x8e
    "10000110", --  988 - 0x3dc  :  134 - 0x86
    "10011100", --  989 - 0x3dd  :  156 - 0x9c
    "01111000", --  990 - 0x3de  :  120 - 0x78
    "00000000", --  991 - 0x3df  :    0 - 0x0
    "00000000", --  992 - 0x3e0  :    0 - 0x0 -- Background 0x7c
    "00000001", --  993 - 0x3e1  :    1 - 0x1
    "00000110", --  994 - 0x3e2  :    6 - 0x6
    "00000111", --  995 - 0x3e3  :    7 - 0x7
    "00000111", --  996 - 0x3e4  :    7 - 0x7
    "00000111", --  997 - 0x3e5  :    7 - 0x7
    "00000001", --  998 - 0x3e6  :    1 - 0x1
    "00000011", --  999 - 0x3e7  :    3 - 0x3
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0 -- Background 0x7d
    "11000000", -- 1001 - 0x3e9  :  192 - 0xc0
    "00110000", -- 1002 - 0x3ea  :   48 - 0x30
    "11110000", -- 1003 - 0x3eb  :  240 - 0xf0
    "11110000", -- 1004 - 0x3ec  :  240 - 0xf0
    "11110000", -- 1005 - 0x3ed  :  240 - 0xf0
    "01000000", -- 1006 - 0x3ee  :   64 - 0x40
    "01000000", -- 1007 - 0x3ef  :   64 - 0x40
    "00000001", -- 1008 - 0x3f0  :    1 - 0x1 -- Background 0x7e
    "00000000", -- 1009 - 0x3f1  :    0 - 0x0
    "00000001", -- 1010 - 0x3f2  :    1 - 0x1
    "00000011", -- 1011 - 0x3f3  :    3 - 0x3
    "00000001", -- 1012 - 0x3f4  :    1 - 0x1
    "00000000", -- 1013 - 0x3f5  :    0 - 0x0
    "00000000", -- 1014 - 0x3f6  :    0 - 0x0
    "00000000", -- 1015 - 0x3f7  :    0 - 0x0
    "01000000", -- 1016 - 0x3f8  :   64 - 0x40 -- Background 0x7f
    "01000000", -- 1017 - 0x3f9  :   64 - 0x40
    "01000000", -- 1018 - 0x3fa  :   64 - 0x40
    "01000000", -- 1019 - 0x3fb  :   64 - 0x40
    "01000000", -- 1020 - 0x3fc  :   64 - 0x40
    "10000000", -- 1021 - 0x3fd  :  128 - 0x80
    "00000000", -- 1022 - 0x3fe  :    0 - 0x0
    "00000000", -- 1023 - 0x3ff  :    0 - 0x0
    "00000000", -- 1024 - 0x400  :    0 - 0x0 -- Background 0x80
    "00000000", -- 1025 - 0x401  :    0 - 0x0
    "00000000", -- 1026 - 0x402  :    0 - 0x0
    "00000000", -- 1027 - 0x403  :    0 - 0x0
    "00000000", -- 1028 - 0x404  :    0 - 0x0
    "00011111", -- 1029 - 0x405  :   31 - 0x1f
    "00010000", -- 1030 - 0x406  :   16 - 0x10
    "00010111", -- 1031 - 0x407  :   23 - 0x17
    "00000000", -- 1032 - 0x408  :    0 - 0x0 -- Background 0x81
    "00000000", -- 1033 - 0x409  :    0 - 0x0
    "00000000", -- 1034 - 0x40a  :    0 - 0x0
    "00000000", -- 1035 - 0x40b  :    0 - 0x0
    "00000000", -- 1036 - 0x40c  :    0 - 0x0
    "11111111", -- 1037 - 0x40d  :  255 - 0xff
    "00000000", -- 1038 - 0x40e  :    0 - 0x0
    "11111111", -- 1039 - 0x40f  :  255 - 0xff
    "00000000", -- 1040 - 0x410  :    0 - 0x0 -- Background 0x82
    "00000000", -- 1041 - 0x411  :    0 - 0x0
    "00000000", -- 1042 - 0x412  :    0 - 0x0
    "00000000", -- 1043 - 0x413  :    0 - 0x0
    "00000000", -- 1044 - 0x414  :    0 - 0x0
    "10000000", -- 1045 - 0x415  :  128 - 0x80
    "00000000", -- 1046 - 0x416  :    0 - 0x0
    "11000000", -- 1047 - 0x417  :  192 - 0xc0
    "00000000", -- 1048 - 0x418  :    0 - 0x0 -- Background 0x83
    "00000000", -- 1049 - 0x419  :    0 - 0x0
    "00000000", -- 1050 - 0x41a  :    0 - 0x0
    "00000000", -- 1051 - 0x41b  :    0 - 0x0
    "00000000", -- 1052 - 0x41c  :    0 - 0x0
    "00001000", -- 1053 - 0x41d  :    8 - 0x8
    "00001000", -- 1054 - 0x41e  :    8 - 0x8
    "00010110", -- 1055 - 0x41f  :   22 - 0x16
    "00000000", -- 1056 - 0x420  :    0 - 0x0 -- Background 0x84
    "00000000", -- 1057 - 0x421  :    0 - 0x0
    "00000000", -- 1058 - 0x422  :    0 - 0x0
    "00000000", -- 1059 - 0x423  :    0 - 0x0
    "00000000", -- 1060 - 0x424  :    0 - 0x0
    "00000000", -- 1061 - 0x425  :    0 - 0x0
    "01000000", -- 1062 - 0x426  :   64 - 0x40
    "11000000", -- 1063 - 0x427  :  192 - 0xc0
    "00000000", -- 1064 - 0x428  :    0 - 0x0 -- Background 0x85
    "00000000", -- 1065 - 0x429  :    0 - 0x0
    "00000000", -- 1066 - 0x42a  :    0 - 0x0
    "00000000", -- 1067 - 0x42b  :    0 - 0x0
    "00000000", -- 1068 - 0x42c  :    0 - 0x0
    "00000001", -- 1069 - 0x42d  :    1 - 0x1
    "00000111", -- 1070 - 0x42e  :    7 - 0x7
    "00001100", -- 1071 - 0x42f  :   12 - 0xc
    "00000000", -- 1072 - 0x430  :    0 - 0x0 -- Background 0x86
    "00000000", -- 1073 - 0x431  :    0 - 0x0
    "00000000", -- 1074 - 0x432  :    0 - 0x0
    "00000000", -- 1075 - 0x433  :    0 - 0x0
    "00000000", -- 1076 - 0x434  :    0 - 0x0
    "11000000", -- 1077 - 0x435  :  192 - 0xc0
    "00111111", -- 1078 - 0x436  :   63 - 0x3f
    "11111111", -- 1079 - 0x437  :  255 - 0xff
    "00000000", -- 1080 - 0x438  :    0 - 0x0 -- Background 0x87
    "00000000", -- 1081 - 0x439  :    0 - 0x0
    "00000000", -- 1082 - 0x43a  :    0 - 0x0
    "00000000", -- 1083 - 0x43b  :    0 - 0x0
    "00000000", -- 1084 - 0x43c  :    0 - 0x0
    "00000000", -- 1085 - 0x43d  :    0 - 0x0
    "00000000", -- 1086 - 0x43e  :    0 - 0x0
    "11000000", -- 1087 - 0x43f  :  192 - 0xc0
    "00000000", -- 1088 - 0x440  :    0 - 0x0 -- Background 0x88
    "00000000", -- 1089 - 0x441  :    0 - 0x0
    "00000000", -- 1090 - 0x442  :    0 - 0x0
    "00000000", -- 1091 - 0x443  :    0 - 0x0
    "00000000", -- 1092 - 0x444  :    0 - 0x0
    "00000000", -- 1093 - 0x445  :    0 - 0x0
    "00000000", -- 1094 - 0x446  :    0 - 0x0
    "00000000", -- 1095 - 0x447  :    0 - 0x0
    "00000000", -- 1096 - 0x448  :    0 - 0x0 -- Background 0x89
    "00000000", -- 1097 - 0x449  :    0 - 0x0
    "00000000", -- 1098 - 0x44a  :    0 - 0x0
    "00000000", -- 1099 - 0x44b  :    0 - 0x0
    "00000000", -- 1100 - 0x44c  :    0 - 0x0
    "01000100", -- 1101 - 0x44d  :   68 - 0x44
    "01010110", -- 1102 - 0x44e  :   86 - 0x56
    "01011011", -- 1103 - 0x44f  :   91 - 0x5b
    "00000000", -- 1104 - 0x450  :    0 - 0x0 -- Background 0x8a
    "00000000", -- 1105 - 0x451  :    0 - 0x0
    "00000000", -- 1106 - 0x452  :    0 - 0x0
    "00000000", -- 1107 - 0x453  :    0 - 0x0
    "00000000", -- 1108 - 0x454  :    0 - 0x0
    "00000000", -- 1109 - 0x455  :    0 - 0x0
    "00000000", -- 1110 - 0x456  :    0 - 0x0
    "00000000", -- 1111 - 0x457  :    0 - 0x0
    "00000000", -- 1112 - 0x458  :    0 - 0x0 -- Background 0x8b
    "00000000", -- 1113 - 0x459  :    0 - 0x0
    "00000000", -- 1114 - 0x45a  :    0 - 0x0
    "00000000", -- 1115 - 0x45b  :    0 - 0x0
    "00000000", -- 1116 - 0x45c  :    0 - 0x0
    "00010000", -- 1117 - 0x45d  :   16 - 0x10
    "00110100", -- 1118 - 0x45e  :   52 - 0x34
    "01101101", -- 1119 - 0x45f  :  109 - 0x6d
    "00000000", -- 1120 - 0x460  :    0 - 0x0 -- Background 0x8c
    "00000000", -- 1121 - 0x461  :    0 - 0x0
    "00000000", -- 1122 - 0x462  :    0 - 0x0
    "00000000", -- 1123 - 0x463  :    0 - 0x0
    "00000000", -- 1124 - 0x464  :    0 - 0x0
    "00000000", -- 1125 - 0x465  :    0 - 0x0
    "00000000", -- 1126 - 0x466  :    0 - 0x0
    "00000000", -- 1127 - 0x467  :    0 - 0x0
    "00000000", -- 1128 - 0x468  :    0 - 0x0 -- Background 0x8d
    "00000000", -- 1129 - 0x469  :    0 - 0x0
    "00000000", -- 1130 - 0x46a  :    0 - 0x0
    "00000000", -- 1131 - 0x46b  :    0 - 0x0
    "01000000", -- 1132 - 0x46c  :   64 - 0x40
    "01001000", -- 1133 - 0x46d  :   72 - 0x48
    "10101000", -- 1134 - 0x46e  :  168 - 0xa8
    "10101100", -- 1135 - 0x46f  :  172 - 0xac
    "00000000", -- 1136 - 0x470  :    0 - 0x0 -- Background 0x8e
    "00000000", -- 1137 - 0x471  :    0 - 0x0
    "00000000", -- 1138 - 0x472  :    0 - 0x0
    "00000000", -- 1139 - 0x473  :    0 - 0x0
    "00000010", -- 1140 - 0x474  :    2 - 0x2
    "00000010", -- 1141 - 0x475  :    2 - 0x2
    "00000010", -- 1142 - 0x476  :    2 - 0x2
    "00000010", -- 1143 - 0x477  :    2 - 0x2
    "00000000", -- 1144 - 0x478  :    0 - 0x0 -- Background 0x8f
    "00000000", -- 1145 - 0x479  :    0 - 0x0
    "00000000", -- 1146 - 0x47a  :    0 - 0x0
    "00000011", -- 1147 - 0x47b  :    3 - 0x3
    "01000011", -- 1148 - 0x47c  :   67 - 0x43
    "01100010", -- 1149 - 0x47d  :   98 - 0x62
    "10110010", -- 1150 - 0x47e  :  178 - 0xb2
    "11011010", -- 1151 - 0x47f  :  218 - 0xda
    "00000000", -- 1152 - 0x480  :    0 - 0x0 -- Background 0x90
    "00000000", -- 1153 - 0x481  :    0 - 0x0
    "00000000", -- 1154 - 0x482  :    0 - 0x0
    "11111100", -- 1155 - 0x483  :  252 - 0xfc
    "11111100", -- 1156 - 0x484  :  252 - 0xfc
    "00000000", -- 1157 - 0x485  :    0 - 0x0
    "11111111", -- 1158 - 0x486  :  255 - 0xff
    "11111111", -- 1159 - 0x487  :  255 - 0xff
    "00000000", -- 1160 - 0x488  :    0 - 0x0 -- Background 0x91
    "00000000", -- 1161 - 0x489  :    0 - 0x0
    "00000000", -- 1162 - 0x48a  :    0 - 0x0
    "00000000", -- 1163 - 0x48b  :    0 - 0x0
    "00000000", -- 1164 - 0x48c  :    0 - 0x0
    "00000000", -- 1165 - 0x48d  :    0 - 0x0
    "00000000", -- 1166 - 0x48e  :    0 - 0x0
    "00000000", -- 1167 - 0x48f  :    0 - 0x0
    "00010111", -- 1168 - 0x490  :   23 - 0x17 -- Background 0x92
    "00010111", -- 1169 - 0x491  :   23 - 0x17
    "00010111", -- 1170 - 0x492  :   23 - 0x17
    "00010111", -- 1171 - 0x493  :   23 - 0x17
    "00010111", -- 1172 - 0x494  :   23 - 0x17
    "00010111", -- 1173 - 0x495  :   23 - 0x17
    "00010111", -- 1174 - 0x496  :   23 - 0x17
    "00010111", -- 1175 - 0x497  :   23 - 0x17
    "11111111", -- 1176 - 0x498  :  255 - 0xff -- Background 0x93
    "11111111", -- 1177 - 0x499  :  255 - 0xff
    "11111111", -- 1178 - 0x49a  :  255 - 0xff
    "11111111", -- 1179 - 0x49b  :  255 - 0xff
    "11111001", -- 1180 - 0x49c  :  249 - 0xf9
    "11111001", -- 1181 - 0x49d  :  249 - 0xf9
    "11111111", -- 1182 - 0x49e  :  255 - 0xff
    "11111111", -- 1183 - 0x49f  :  255 - 0xff
    "11110000", -- 1184 - 0x4a0  :  240 - 0xf0 -- Background 0x94
    "11111000", -- 1185 - 0x4a1  :  248 - 0xf8
    "11111000", -- 1186 - 0x4a2  :  248 - 0xf8
    "11111100", -- 1187 - 0x4a3  :  252 - 0xfc
    "11111100", -- 1188 - 0x4a4  :  252 - 0xfc
    "11111100", -- 1189 - 0x4a5  :  252 - 0xfc
    "01111100", -- 1190 - 0x4a6  :  124 - 0x7c
    "01111100", -- 1191 - 0x4a7  :  124 - 0x7c
    "00010111", -- 1192 - 0x4a8  :   23 - 0x17 -- Background 0x95
    "00101111", -- 1193 - 0x4a9  :   47 - 0x2f
    "00101111", -- 1194 - 0x4aa  :   47 - 0x2f
    "01011111", -- 1195 - 0x4ab  :   95 - 0x5f
    "01011111", -- 1196 - 0x4ac  :   95 - 0x5f
    "10111111", -- 1197 - 0x4ad  :  191 - 0xbf
    "10111111", -- 1198 - 0x4ae  :  191 - 0xbf
    "01111111", -- 1199 - 0x4af  :  127 - 0x7f
    "01100000", -- 1200 - 0x4b0  :   96 - 0x60 -- Background 0x96
    "01100000", -- 1201 - 0x4b1  :   96 - 0x60
    "10110000", -- 1202 - 0x4b2  :  176 - 0xb0
    "10110000", -- 1203 - 0x4b3  :  176 - 0xb0
    "11011000", -- 1204 - 0x4b4  :  216 - 0xd8
    "11011000", -- 1205 - 0x4b5  :  216 - 0xd8
    "11101100", -- 1206 - 0x4b6  :  236 - 0xec
    "11101100", -- 1207 - 0x4b7  :  236 - 0xec
    "00110011", -- 1208 - 0x4b8  :   51 - 0x33 -- Background 0x97
    "00101111", -- 1209 - 0x4b9  :   47 - 0x2f
    "01101111", -- 1210 - 0x4ba  :  111 - 0x6f
    "01011111", -- 1211 - 0x4bb  :   95 - 0x5f
    "11011111", -- 1212 - 0x4bc  :  223 - 0xdf
    "10111111", -- 1213 - 0x4bd  :  191 - 0xbf
    "10111111", -- 1214 - 0x4be  :  191 - 0xbf
    "10111111", -- 1215 - 0x4bf  :  191 - 0xbf
    "11111111", -- 1216 - 0x4c0  :  255 - 0xff -- Background 0x98
    "11111111", -- 1217 - 0x4c1  :  255 - 0xff
    "11111111", -- 1218 - 0x4c2  :  255 - 0xff
    "11111110", -- 1219 - 0x4c3  :  254 - 0xfe
    "11111001", -- 1220 - 0x4c4  :  249 - 0xf9
    "11100111", -- 1221 - 0x4c5  :  231 - 0xe7
    "11111100", -- 1222 - 0x4c6  :  252 - 0xfc
    "11110011", -- 1223 - 0x4c7  :  243 - 0xf3
    "11110000", -- 1224 - 0x4c8  :  240 - 0xf0 -- Background 0x99
    "11111000", -- 1225 - 0x4c9  :  248 - 0xf8
    "11111000", -- 1226 - 0x4ca  :  248 - 0xf8
    "01110000", -- 1227 - 0x4cb  :  112 - 0x70
    "11001100", -- 1228 - 0x4cc  :  204 - 0xcc
    "00110000", -- 1229 - 0x4cd  :   48 - 0x30
    "11000000", -- 1230 - 0x4ce  :  192 - 0xc0
    "00000000", -- 1231 - 0x4cf  :    0 - 0x0
    "00000000", -- 1232 - 0x4d0  :    0 - 0x0 -- Background 0x9a
    "00000000", -- 1233 - 0x4d1  :    0 - 0x0
    "00000000", -- 1234 - 0x4d2  :    0 - 0x0
    "00000000", -- 1235 - 0x4d3  :    0 - 0x0
    "00111111", -- 1236 - 0x4d4  :   63 - 0x3f
    "00100000", -- 1237 - 0x4d5  :   32 - 0x20
    "00101111", -- 1238 - 0x4d6  :   47 - 0x2f
    "00101111", -- 1239 - 0x4d7  :   47 - 0x2f
    "00000000", -- 1240 - 0x4d8  :    0 - 0x0 -- Background 0x9b
    "00000000", -- 1241 - 0x4d9  :    0 - 0x0
    "00000000", -- 1242 - 0x4da  :    0 - 0x0
    "00000000", -- 1243 - 0x4db  :    0 - 0x0
    "11100000", -- 1244 - 0x4dc  :  224 - 0xe0
    "00000000", -- 1245 - 0x4dd  :    0 - 0x0
    "11110000", -- 1246 - 0x4de  :  240 - 0xf0
    "11110000", -- 1247 - 0x4df  :  240 - 0xf0
    "01011101", -- 1248 - 0x4e0  :   93 - 0x5d -- Background 0x9c
    "01011110", -- 1249 - 0x4e1  :   94 - 0x5e
    "01011111", -- 1250 - 0x4e2  :   95 - 0x5f
    "01011111", -- 1251 - 0x4e3  :   95 - 0x5f
    "01011111", -- 1252 - 0x4e4  :   95 - 0x5f
    "01011111", -- 1253 - 0x4e5  :   95 - 0x5f
    "01011111", -- 1254 - 0x4e6  :   95 - 0x5f
    "01011111", -- 1255 - 0x4e7  :   95 - 0x5f
    "10000000", -- 1256 - 0x4e8  :  128 - 0x80 -- Background 0x9d
    "11000001", -- 1257 - 0x4e9  :  193 - 0xc1
    "01100011", -- 1258 - 0x4ea  :   99 - 0x63
    "10110110", -- 1259 - 0x4eb  :  182 - 0xb6
    "11011001", -- 1260 - 0x4ec  :  217 - 0xd9
    "11101011", -- 1261 - 0x4ed  :  235 - 0xeb
    "11110111", -- 1262 - 0x4ee  :  247 - 0xf7
    "11111111", -- 1263 - 0x4ef  :  255 - 0xff
    "11011101", -- 1264 - 0x4f0  :  221 - 0xdd -- Background 0x9e
    "10111101", -- 1265 - 0x4f1  :  189 - 0xbd
    "01111101", -- 1266 - 0x4f2  :  125 - 0x7d
    "11111101", -- 1267 - 0x4f3  :  253 - 0xfd
    "11111101", -- 1268 - 0x4f4  :  253 - 0xfd
    "11111101", -- 1269 - 0x4f5  :  253 - 0xfd
    "11111101", -- 1270 - 0x4f6  :  253 - 0xfd
    "11111101", -- 1271 - 0x4f7  :  253 - 0xfd
    "00000001", -- 1272 - 0x4f8  :    1 - 0x1 -- Background 0x9f
    "00000001", -- 1273 - 0x4f9  :    1 - 0x1
    "00000010", -- 1274 - 0x4fa  :    2 - 0x2
    "00000010", -- 1275 - 0x4fb  :    2 - 0x2
    "00000101", -- 1276 - 0x4fc  :    5 - 0x5
    "00000101", -- 1277 - 0x4fd  :    5 - 0x5
    "00001011", -- 1278 - 0x4fe  :   11 - 0xb
    "00001011", -- 1279 - 0x4ff  :   11 - 0xb
    "01110100", -- 1280 - 0x500  :  116 - 0x74 -- Background 0xa0
    "01110110", -- 1281 - 0x501  :  118 - 0x76
    "11111010", -- 1282 - 0x502  :  250 - 0xfa
    "11111011", -- 1283 - 0x503  :  251 - 0xfb
    "11111101", -- 1284 - 0x504  :  253 - 0xfd
    "11111101", -- 1285 - 0x505  :  253 - 0xfd
    "11111110", -- 1286 - 0x506  :  254 - 0xfe
    "11111110", -- 1287 - 0x507  :  254 - 0xfe
    "00000010", -- 1288 - 0x508  :    2 - 0x2 -- Background 0xa1
    "00000010", -- 1289 - 0x509  :    2 - 0x2
    "00000010", -- 1290 - 0x50a  :    2 - 0x2
    "00000010", -- 1291 - 0x50b  :    2 - 0x2
    "00000010", -- 1292 - 0x50c  :    2 - 0x2
    "10000010", -- 1293 - 0x50d  :  130 - 0x82
    "10000010", -- 1294 - 0x50e  :  130 - 0x82
    "11000010", -- 1295 - 0x50f  :  194 - 0xc2
    "11101010", -- 1296 - 0x510  :  234 - 0xea -- Background 0xa2
    "11110110", -- 1297 - 0x511  :  246 - 0xf6
    "11111010", -- 1298 - 0x512  :  250 - 0xfa
    "11111010", -- 1299 - 0x513  :  250 - 0xfa
    "11111100", -- 1300 - 0x514  :  252 - 0xfc
    "11111100", -- 1301 - 0x515  :  252 - 0xfc
    "11111110", -- 1302 - 0x516  :  254 - 0xfe
    "11111111", -- 1303 - 0x517  :  255 - 0xff
    "11111111", -- 1304 - 0x518  :  255 - 0xff -- Background 0xa3
    "11111111", -- 1305 - 0x519  :  255 - 0xff
    "11111111", -- 1306 - 0x51a  :  255 - 0xff
    "11111111", -- 1307 - 0x51b  :  255 - 0xff
    "11111111", -- 1308 - 0x51c  :  255 - 0xff
    "11111111", -- 1309 - 0x51d  :  255 - 0xff
    "11111111", -- 1310 - 0x51e  :  255 - 0xff
    "11111111", -- 1311 - 0x51f  :  255 - 0xff
    "01000000", -- 1312 - 0x520  :   64 - 0x40 -- Background 0xa4
    "01000000", -- 1313 - 0x521  :   64 - 0x40
    "01000000", -- 1314 - 0x522  :   64 - 0x40
    "01000000", -- 1315 - 0x523  :   64 - 0x40
    "01000000", -- 1316 - 0x524  :   64 - 0x40
    "01000000", -- 1317 - 0x525  :   64 - 0x40
    "01000000", -- 1318 - 0x526  :   64 - 0x40
    "01000000", -- 1319 - 0x527  :   64 - 0x40
    "11111000", -- 1320 - 0x528  :  248 - 0xf8 -- Background 0xa5
    "11111111", -- 1321 - 0x529  :  255 - 0xff
    "11111111", -- 1322 - 0x52a  :  255 - 0xff
    "11111000", -- 1323 - 0x52b  :  248 - 0xf8
    "11111011", -- 1324 - 0x52c  :  251 - 0xfb
    "11111010", -- 1325 - 0x52d  :  250 - 0xfa
    "11111010", -- 1326 - 0x52e  :  250 - 0xfa
    "11111010", -- 1327 - 0x52f  :  250 - 0xfa
    "11111100", -- 1328 - 0x530  :  252 - 0xfc -- Background 0xa6
    "11111010", -- 1329 - 0x531  :  250 - 0xfa
    "11110110", -- 1330 - 0x532  :  246 - 0xf6
    "00001101", -- 1331 - 0x533  :   13 - 0xd
    "11111001", -- 1332 - 0x534  :  249 - 0xf9
    "00000011", -- 1333 - 0x535  :    3 - 0x3
    "00010011", -- 1334 - 0x536  :   19 - 0x13
    "00110111", -- 1335 - 0x537  :   55 - 0x37
    "01111111", -- 1336 - 0x538  :  127 - 0x7f -- Background 0xa7
    "11111001", -- 1337 - 0x539  :  249 - 0xf9
    "11111001", -- 1338 - 0x53a  :  249 - 0xf9
    "11111111", -- 1339 - 0x53b  :  255 - 0xff
    "11111110", -- 1340 - 0x53c  :  254 - 0xfe
    "11111100", -- 1341 - 0x53d  :  252 - 0xfc
    "11111111", -- 1342 - 0x53e  :  255 - 0xff
    "11111111", -- 1343 - 0x53f  :  255 - 0xff
    "11110110", -- 1344 - 0x540  :  246 - 0xf6 -- Background 0xa8
    "11110110", -- 1345 - 0x541  :  246 - 0xf6
    "11111011", -- 1346 - 0x542  :  251 - 0xfb
    "01111011", -- 1347 - 0x543  :  123 - 0x7b
    "11111101", -- 1348 - 0x544  :  253 - 0xfd
    "11110101", -- 1349 - 0x545  :  245 - 0xf5
    "11110110", -- 1350 - 0x546  :  246 - 0xf6
    "11111010", -- 1351 - 0x547  :  250 - 0xfa
    "10111111", -- 1352 - 0x548  :  191 - 0xbf -- Background 0xa9
    "10111111", -- 1353 - 0x549  :  191 - 0xbf
    "00111111", -- 1354 - 0x54a  :   63 - 0x3f
    "00111111", -- 1355 - 0x54b  :   63 - 0x3f
    "10111111", -- 1356 - 0x54c  :  191 - 0xbf
    "10011111", -- 1357 - 0x54d  :  159 - 0x9f
    "11001111", -- 1358 - 0x54e  :  207 - 0xcf
    "11010111", -- 1359 - 0x54f  :  215 - 0xd7
    "11100100", -- 1360 - 0x550  :  228 - 0xe4 -- Background 0xaa
    "11111000", -- 1361 - 0x551  :  248 - 0xf8
    "11111111", -- 1362 - 0x552  :  255 - 0xff
    "11110011", -- 1363 - 0x553  :  243 - 0xf3
    "11111100", -- 1364 - 0x554  :  252 - 0xfc
    "11111111", -- 1365 - 0x555  :  255 - 0xff
    "11111111", -- 1366 - 0x556  :  255 - 0xff
    "11111111", -- 1367 - 0x557  :  255 - 0xff
    "00000000", -- 1368 - 0x558  :    0 - 0x0 -- Background 0xab
    "00000000", -- 1369 - 0x559  :    0 - 0x0
    "00000000", -- 1370 - 0x55a  :    0 - 0x0
    "11000000", -- 1371 - 0x55b  :  192 - 0xc0
    "11110000", -- 1372 - 0x55c  :  240 - 0xf0
    "00111100", -- 1373 - 0x55d  :   60 - 0x3c
    "11011000", -- 1374 - 0x55e  :  216 - 0xd8
    "10110110", -- 1375 - 0x55f  :  182 - 0xb6
    "00001111", -- 1376 - 0x560  :   15 - 0xf -- Background 0xac
    "00001111", -- 1377 - 0x561  :   15 - 0xf
    "00000000", -- 1378 - 0x562  :    0 - 0x0
    "00000011", -- 1379 - 0x563  :    3 - 0x3
    "00000000", -- 1380 - 0x564  :    0 - 0x0
    "00000000", -- 1381 - 0x565  :    0 - 0x0
    "00000000", -- 1382 - 0x566  :    0 - 0x0
    "00000000", -- 1383 - 0x567  :    0 - 0x0
    "11110100", -- 1384 - 0x568  :  244 - 0xf4 -- Background 0xad
    "11110100", -- 1385 - 0x569  :  244 - 0xf4
    "00000100", -- 1386 - 0x56a  :    4 - 0x4
    "11111100", -- 1387 - 0x56b  :  252 - 0xfc
    "00000000", -- 1388 - 0x56c  :    0 - 0x0
    "00000000", -- 1389 - 0x56d  :    0 - 0x0
    "00000000", -- 1390 - 0x56e  :    0 - 0x0
    "00000000", -- 1391 - 0x56f  :    0 - 0x0
    "01011111", -- 1392 - 0x570  :   95 - 0x5f -- Background 0xae
    "01011111", -- 1393 - 0x571  :   95 - 0x5f
    "01011111", -- 1394 - 0x572  :   95 - 0x5f
    "01011111", -- 1395 - 0x573  :   95 - 0x5f
    "01011111", -- 1396 - 0x574  :   95 - 0x5f
    "01011111", -- 1397 - 0x575  :   95 - 0x5f
    "01011111", -- 1398 - 0x576  :   95 - 0x5f
    "01011111", -- 1399 - 0x577  :   95 - 0x5f
    "11111101", -- 1400 - 0x578  :  253 - 0xfd -- Background 0xaf
    "11111101", -- 1401 - 0x579  :  253 - 0xfd
    "11111101", -- 1402 - 0x57a  :  253 - 0xfd
    "11111101", -- 1403 - 0x57b  :  253 - 0xfd
    "11110101", -- 1404 - 0x57c  :  245 - 0xf5
    "11110101", -- 1405 - 0x57d  :  245 - 0xf5
    "11110101", -- 1406 - 0x57e  :  245 - 0xf5
    "11110101", -- 1407 - 0x57f  :  245 - 0xf5
    "00001100", -- 1408 - 0x580  :   12 - 0xc -- Background 0xb0
    "00011100", -- 1409 - 0x581  :   28 - 0x1c
    "00001100", -- 1410 - 0x582  :   12 - 0xc
    "00001100", -- 1411 - 0x583  :   12 - 0xc
    "00001100", -- 1412 - 0x584  :   12 - 0xc
    "00001100", -- 1413 - 0x585  :   12 - 0xc
    "00111111", -- 1414 - 0x586  :   63 - 0x3f
    "00000000", -- 1415 - 0x587  :    0 - 0x0
    "00111110", -- 1416 - 0x588  :   62 - 0x3e -- Background 0xb1
    "01100011", -- 1417 - 0x589  :   99 - 0x63
    "00000111", -- 1418 - 0x58a  :    7 - 0x7
    "00011110", -- 1419 - 0x58b  :   30 - 0x1e
    "00111100", -- 1420 - 0x58c  :   60 - 0x3c
    "01110000", -- 1421 - 0x58d  :  112 - 0x70
    "01111111", -- 1422 - 0x58e  :  127 - 0x7f
    "00000000", -- 1423 - 0x58f  :    0 - 0x0
    "01111110", -- 1424 - 0x590  :  126 - 0x7e -- Background 0xb2
    "01100011", -- 1425 - 0x591  :   99 - 0x63
    "01100011", -- 1426 - 0x592  :   99 - 0x63
    "01100011", -- 1427 - 0x593  :   99 - 0x63
    "01111110", -- 1428 - 0x594  :  126 - 0x7e
    "01100000", -- 1429 - 0x595  :   96 - 0x60
    "01100000", -- 1430 - 0x596  :   96 - 0x60
    "00000000", -- 1431 - 0x597  :    0 - 0x0
    "01100011", -- 1432 - 0x598  :   99 - 0x63 -- Background 0xb3
    "01100011", -- 1433 - 0x599  :   99 - 0x63
    "01100011", -- 1434 - 0x59a  :   99 - 0x63
    "01100011", -- 1435 - 0x59b  :   99 - 0x63
    "01100011", -- 1436 - 0x59c  :   99 - 0x63
    "01100011", -- 1437 - 0x59d  :   99 - 0x63
    "00111110", -- 1438 - 0x59e  :   62 - 0x3e
    "00000000", -- 1439 - 0x59f  :    0 - 0x0
    "01100011", -- 1440 - 0x5a0  :   99 - 0x63 -- Background 0xb4
    "01100011", -- 1441 - 0x5a1  :   99 - 0x63
    "01100011", -- 1442 - 0x5a2  :   99 - 0x63
    "01111111", -- 1443 - 0x5a3  :  127 - 0x7f
    "01100011", -- 1444 - 0x5a4  :   99 - 0x63
    "01100011", -- 1445 - 0x5a5  :   99 - 0x63
    "01100011", -- 1446 - 0x5a6  :   99 - 0x63
    "00000000", -- 1447 - 0x5a7  :    0 - 0x0
    "00111111", -- 1448 - 0x5a8  :   63 - 0x3f -- Background 0xb5
    "00001100", -- 1449 - 0x5a9  :   12 - 0xc
    "00001100", -- 1450 - 0x5aa  :   12 - 0xc
    "00001100", -- 1451 - 0x5ab  :   12 - 0xc
    "00001100", -- 1452 - 0x5ac  :   12 - 0xc
    "00001100", -- 1453 - 0x5ad  :   12 - 0xc
    "00111111", -- 1454 - 0x5ae  :   63 - 0x3f
    "00000000", -- 1455 - 0x5af  :    0 - 0x0
    "00000000", -- 1456 - 0x5b0  :    0 - 0x0 -- Background 0xb6
    "00000000", -- 1457 - 0x5b1  :    0 - 0x0
    "00000000", -- 1458 - 0x5b2  :    0 - 0x0
    "01111110", -- 1459 - 0x5b3  :  126 - 0x7e
    "00000000", -- 1460 - 0x5b4  :    0 - 0x0
    "00000000", -- 1461 - 0x5b5  :    0 - 0x0
    "00000000", -- 1462 - 0x5b6  :    0 - 0x0
    "00000000", -- 1463 - 0x5b7  :    0 - 0x0
    "00111100", -- 1464 - 0x5b8  :   60 - 0x3c -- Background 0xb7
    "01100110", -- 1465 - 0x5b9  :  102 - 0x66
    "01100000", -- 1466 - 0x5ba  :   96 - 0x60
    "00111110", -- 1467 - 0x5bb  :   62 - 0x3e
    "00000011", -- 1468 - 0x5bc  :    3 - 0x3
    "01100011", -- 1469 - 0x5bd  :   99 - 0x63
    "00111110", -- 1470 - 0x5be  :   62 - 0x3e
    "00000000", -- 1471 - 0x5bf  :    0 - 0x0
    "00011110", -- 1472 - 0x5c0  :   30 - 0x1e -- Background 0xb8
    "00110011", -- 1473 - 0x5c1  :   51 - 0x33
    "01100000", -- 1474 - 0x5c2  :   96 - 0x60
    "01100000", -- 1475 - 0x5c3  :   96 - 0x60
    "01100000", -- 1476 - 0x5c4  :   96 - 0x60
    "00110011", -- 1477 - 0x5c5  :   51 - 0x33
    "00011110", -- 1478 - 0x5c6  :   30 - 0x1e
    "00000000", -- 1479 - 0x5c7  :    0 - 0x0
    "00111110", -- 1480 - 0x5c8  :   62 - 0x3e -- Background 0xb9
    "01100011", -- 1481 - 0x5c9  :   99 - 0x63
    "01100011", -- 1482 - 0x5ca  :   99 - 0x63
    "01100011", -- 1483 - 0x5cb  :   99 - 0x63
    "01100011", -- 1484 - 0x5cc  :   99 - 0x63
    "01100011", -- 1485 - 0x5cd  :   99 - 0x63
    "00111110", -- 1486 - 0x5ce  :   62 - 0x3e
    "00000000", -- 1487 - 0x5cf  :    0 - 0x0
    "01111110", -- 1488 - 0x5d0  :  126 - 0x7e -- Background 0xba
    "01100011", -- 1489 - 0x5d1  :   99 - 0x63
    "01100011", -- 1490 - 0x5d2  :   99 - 0x63
    "01100111", -- 1491 - 0x5d3  :  103 - 0x67
    "01111100", -- 1492 - 0x5d4  :  124 - 0x7c
    "01101110", -- 1493 - 0x5d5  :  110 - 0x6e
    "01100111", -- 1494 - 0x5d6  :  103 - 0x67
    "00000000", -- 1495 - 0x5d7  :    0 - 0x0
    "01111111", -- 1496 - 0x5d8  :  127 - 0x7f -- Background 0xbb
    "01100000", -- 1497 - 0x5d9  :   96 - 0x60
    "01100000", -- 1498 - 0x5da  :   96 - 0x60
    "01111110", -- 1499 - 0x5db  :  126 - 0x7e
    "01100000", -- 1500 - 0x5dc  :   96 - 0x60
    "01100000", -- 1501 - 0x5dd  :   96 - 0x60
    "01111111", -- 1502 - 0x5de  :  127 - 0x7f
    "00000000", -- 1503 - 0x5df  :    0 - 0x0
    "00000000", -- 1504 - 0x5e0  :    0 - 0x0 -- Background 0xbc
    "00000000", -- 1505 - 0x5e1  :    0 - 0x0
    "00000000", -- 1506 - 0x5e2  :    0 - 0x0
    "00000000", -- 1507 - 0x5e3  :    0 - 0x0
    "00000000", -- 1508 - 0x5e4  :    0 - 0x0
    "00000000", -- 1509 - 0x5e5  :    0 - 0x0
    "00000000", -- 1510 - 0x5e6  :    0 - 0x0
    "00000000", -- 1511 - 0x5e7  :    0 - 0x0
    "00000000", -- 1512 - 0x5e8  :    0 - 0x0 -- Background 0xbd
    "00000000", -- 1513 - 0x5e9  :    0 - 0x0
    "00000000", -- 1514 - 0x5ea  :    0 - 0x0
    "00000000", -- 1515 - 0x5eb  :    0 - 0x0
    "00000000", -- 1516 - 0x5ec  :    0 - 0x0
    "00000000", -- 1517 - 0x5ed  :    0 - 0x0
    "00000000", -- 1518 - 0x5ee  :    0 - 0x0
    "00000000", -- 1519 - 0x5ef  :    0 - 0x0
    "00000000", -- 1520 - 0x5f0  :    0 - 0x0 -- Background 0xbe
    "00000000", -- 1521 - 0x5f1  :    0 - 0x0
    "00000000", -- 1522 - 0x5f2  :    0 - 0x0
    "00000000", -- 1523 - 0x5f3  :    0 - 0x0
    "00000000", -- 1524 - 0x5f4  :    0 - 0x0
    "00000000", -- 1525 - 0x5f5  :    0 - 0x0
    "00000000", -- 1526 - 0x5f6  :    0 - 0x0
    "00000000", -- 1527 - 0x5f7  :    0 - 0x0
    "00000000", -- 1528 - 0x5f8  :    0 - 0x0 -- Background 0xbf
    "00000000", -- 1529 - 0x5f9  :    0 - 0x0
    "00000000", -- 1530 - 0x5fa  :    0 - 0x0
    "00000000", -- 1531 - 0x5fb  :    0 - 0x0
    "00000000", -- 1532 - 0x5fc  :    0 - 0x0
    "00000000", -- 1533 - 0x5fd  :    0 - 0x0
    "00000000", -- 1534 - 0x5fe  :    0 - 0x0
    "00000000", -- 1535 - 0x5ff  :    0 - 0x0
    "01100011", -- 1536 - 0x600  :   99 - 0x63 -- Background 0xc0
    "01100110", -- 1537 - 0x601  :  102 - 0x66
    "01101100", -- 1538 - 0x602  :  108 - 0x6c
    "01111000", -- 1539 - 0x603  :  120 - 0x78
    "01111100", -- 1540 - 0x604  :  124 - 0x7c
    "01100110", -- 1541 - 0x605  :  102 - 0x66
    "01100011", -- 1542 - 0x606  :   99 - 0x63
    "00000000", -- 1543 - 0x607  :    0 - 0x0
    "00111111", -- 1544 - 0x608  :   63 - 0x3f -- Background 0xc1
    "00001100", -- 1545 - 0x609  :   12 - 0xc
    "00001100", -- 1546 - 0x60a  :   12 - 0xc
    "00001100", -- 1547 - 0x60b  :   12 - 0xc
    "00001100", -- 1548 - 0x60c  :   12 - 0xc
    "00001100", -- 1549 - 0x60d  :   12 - 0xc
    "00111111", -- 1550 - 0x60e  :   63 - 0x3f
    "00000000", -- 1551 - 0x60f  :    0 - 0x0
    "01100011", -- 1552 - 0x610  :   99 - 0x63 -- Background 0xc2
    "01110111", -- 1553 - 0x611  :  119 - 0x77
    "01111111", -- 1554 - 0x612  :  127 - 0x7f
    "01111111", -- 1555 - 0x613  :  127 - 0x7f
    "01101011", -- 1556 - 0x614  :  107 - 0x6b
    "01100011", -- 1557 - 0x615  :   99 - 0x63
    "01100011", -- 1558 - 0x616  :   99 - 0x63
    "00000000", -- 1559 - 0x617  :    0 - 0x0
    "00011100", -- 1560 - 0x618  :   28 - 0x1c -- Background 0xc3
    "00110110", -- 1561 - 0x619  :   54 - 0x36
    "01100011", -- 1562 - 0x61a  :   99 - 0x63
    "01100011", -- 1563 - 0x61b  :   99 - 0x63
    "01111111", -- 1564 - 0x61c  :  127 - 0x7f
    "01100011", -- 1565 - 0x61d  :   99 - 0x63
    "01100011", -- 1566 - 0x61e  :   99 - 0x63
    "00000000", -- 1567 - 0x61f  :    0 - 0x0
    "00011111", -- 1568 - 0x620  :   31 - 0x1f -- Background 0xc4
    "00110000", -- 1569 - 0x621  :   48 - 0x30
    "01100000", -- 1570 - 0x622  :   96 - 0x60
    "01100111", -- 1571 - 0x623  :  103 - 0x67
    "01100011", -- 1572 - 0x624  :   99 - 0x63
    "00110011", -- 1573 - 0x625  :   51 - 0x33
    "00011111", -- 1574 - 0x626  :   31 - 0x1f
    "00000000", -- 1575 - 0x627  :    0 - 0x0
    "01100011", -- 1576 - 0x628  :   99 - 0x63 -- Background 0xc5
    "01100011", -- 1577 - 0x629  :   99 - 0x63
    "01100011", -- 1578 - 0x62a  :   99 - 0x63
    "01100011", -- 1579 - 0x62b  :   99 - 0x63
    "01100011", -- 1580 - 0x62c  :   99 - 0x63
    "01100011", -- 1581 - 0x62d  :   99 - 0x63
    "00111110", -- 1582 - 0x62e  :   62 - 0x3e
    "00000000", -- 1583 - 0x62f  :    0 - 0x0
    "01111110", -- 1584 - 0x630  :  126 - 0x7e -- Background 0xc6
    "01100011", -- 1585 - 0x631  :   99 - 0x63
    "01100011", -- 1586 - 0x632  :   99 - 0x63
    "01100111", -- 1587 - 0x633  :  103 - 0x67
    "01111100", -- 1588 - 0x634  :  124 - 0x7c
    "01101110", -- 1589 - 0x635  :  110 - 0x6e
    "01100111", -- 1590 - 0x636  :  103 - 0x67
    "00000000", -- 1591 - 0x637  :    0 - 0x0
    "01111111", -- 1592 - 0x638  :  127 - 0x7f -- Background 0xc7
    "01100000", -- 1593 - 0x639  :   96 - 0x60
    "01100000", -- 1594 - 0x63a  :   96 - 0x60
    "01111110", -- 1595 - 0x63b  :  126 - 0x7e
    "01100000", -- 1596 - 0x63c  :   96 - 0x60
    "01100000", -- 1597 - 0x63d  :   96 - 0x60
    "01111111", -- 1598 - 0x63e  :  127 - 0x7f
    "00000000", -- 1599 - 0x63f  :    0 - 0x0
    "00110110", -- 1600 - 0x640  :   54 - 0x36 -- Background 0xc8
    "00110110", -- 1601 - 0x641  :   54 - 0x36
    "00010010", -- 1602 - 0x642  :   18 - 0x12
    "00000000", -- 1603 - 0x643  :    0 - 0x0
    "00000000", -- 1604 - 0x644  :    0 - 0x0
    "00000000", -- 1605 - 0x645  :    0 - 0x0
    "00000000", -- 1606 - 0x646  :    0 - 0x0
    "00000000", -- 1607 - 0x647  :    0 - 0x0
    "00111110", -- 1608 - 0x648  :   62 - 0x3e -- Background 0xc9
    "01100011", -- 1609 - 0x649  :   99 - 0x63
    "01100011", -- 1610 - 0x64a  :   99 - 0x63
    "01100011", -- 1611 - 0x64b  :   99 - 0x63
    "01100011", -- 1612 - 0x64c  :   99 - 0x63
    "01100011", -- 1613 - 0x64d  :   99 - 0x63
    "00111110", -- 1614 - 0x64e  :   62 - 0x3e
    "00000000", -- 1615 - 0x64f  :    0 - 0x0
    "00111100", -- 1616 - 0x650  :   60 - 0x3c -- Background 0xca
    "01100110", -- 1617 - 0x651  :  102 - 0x66
    "01100000", -- 1618 - 0x652  :   96 - 0x60
    "00111110", -- 1619 - 0x653  :   62 - 0x3e
    "00000011", -- 1620 - 0x654  :    3 - 0x3
    "01100011", -- 1621 - 0x655  :   99 - 0x63
    "00111110", -- 1622 - 0x656  :   62 - 0x3e
    "00000000", -- 1623 - 0x657  :    0 - 0x0
    "00000000", -- 1624 - 0x658  :    0 - 0x0 -- Background 0xcb
    "00111000", -- 1625 - 0x659  :   56 - 0x38
    "01111100", -- 1626 - 0x65a  :  124 - 0x7c
    "11111110", -- 1627 - 0x65b  :  254 - 0xfe
    "11111110", -- 1628 - 0x65c  :  254 - 0xfe
    "11111110", -- 1629 - 0x65d  :  254 - 0xfe
    "01111100", -- 1630 - 0x65e  :  124 - 0x7c
    "00111000", -- 1631 - 0x65f  :   56 - 0x38
    "00000000", -- 1632 - 0x660  :    0 - 0x0 -- Background 0xcc
    "00000000", -- 1633 - 0x661  :    0 - 0x0
    "00000000", -- 1634 - 0x662  :    0 - 0x0
    "00000000", -- 1635 - 0x663  :    0 - 0x0
    "00000000", -- 1636 - 0x664  :    0 - 0x0
    "00000000", -- 1637 - 0x665  :    0 - 0x0
    "00000000", -- 1638 - 0x666  :    0 - 0x0
    "00000000", -- 1639 - 0x667  :    0 - 0x0
    "00000000", -- 1640 - 0x668  :    0 - 0x0 -- Background 0xcd
    "00000000", -- 1641 - 0x669  :    0 - 0x0
    "00000000", -- 1642 - 0x66a  :    0 - 0x0
    "00000000", -- 1643 - 0x66b  :    0 - 0x0
    "00000000", -- 1644 - 0x66c  :    0 - 0x0
    "00000000", -- 1645 - 0x66d  :    0 - 0x0
    "00000000", -- 1646 - 0x66e  :    0 - 0x0
    "00000000", -- 1647 - 0x66f  :    0 - 0x0
    "00000000", -- 1648 - 0x670  :    0 - 0x0 -- Background 0xce
    "00000000", -- 1649 - 0x671  :    0 - 0x0
    "00000000", -- 1650 - 0x672  :    0 - 0x0
    "00000000", -- 1651 - 0x673  :    0 - 0x0
    "00000000", -- 1652 - 0x674  :    0 - 0x0
    "00000000", -- 1653 - 0x675  :    0 - 0x0
    "00000000", -- 1654 - 0x676  :    0 - 0x0
    "00000000", -- 1655 - 0x677  :    0 - 0x0
    "00000000", -- 1656 - 0x678  :    0 - 0x0 -- Background 0xcf
    "00000000", -- 1657 - 0x679  :    0 - 0x0
    "00000000", -- 1658 - 0x67a  :    0 - 0x0
    "00000000", -- 1659 - 0x67b  :    0 - 0x0
    "00000000", -- 1660 - 0x67c  :    0 - 0x0
    "00000000", -- 1661 - 0x67d  :    0 - 0x0
    "00000000", -- 1662 - 0x67e  :    0 - 0x0
    "00000000", -- 1663 - 0x67f  :    0 - 0x0
    "00010111", -- 1664 - 0x680  :   23 - 0x17 -- Background 0xd0
    "00010111", -- 1665 - 0x681  :   23 - 0x17
    "00101111", -- 1666 - 0x682  :   47 - 0x2f
    "00101111", -- 1667 - 0x683  :   47 - 0x2f
    "01011111", -- 1668 - 0x684  :   95 - 0x5f
    "01011111", -- 1669 - 0x685  :   95 - 0x5f
    "00111111", -- 1670 - 0x686  :   63 - 0x3f
    "00111111", -- 1671 - 0x687  :   63 - 0x3f
    "11111111", -- 1672 - 0x688  :  255 - 0xff -- Background 0xd1
    "11001111", -- 1673 - 0x689  :  207 - 0xcf
    "11001111", -- 1674 - 0x68a  :  207 - 0xcf
    "11111011", -- 1675 - 0x68b  :  251 - 0xfb
    "11110111", -- 1676 - 0x68c  :  247 - 0xf7
    "11100111", -- 1677 - 0x68d  :  231 - 0xe7
    "11111111", -- 1678 - 0x68e  :  255 - 0xff
    "11111111", -- 1679 - 0x68f  :  255 - 0xff
    "01000010", -- 1680 - 0x690  :   66 - 0x42 -- Background 0xd2
    "01100010", -- 1681 - 0x691  :   98 - 0x62
    "10100010", -- 1682 - 0x692  :  162 - 0xa2
    "10110010", -- 1683 - 0x693  :  178 - 0xb2
    "01010010", -- 1684 - 0x694  :   82 - 0x52
    "01011010", -- 1685 - 0x695  :   90 - 0x5a
    "10101010", -- 1686 - 0x696  :  170 - 0xaa
    "10101100", -- 1687 - 0x697  :  172 - 0xac
    "11111111", -- 1688 - 0x698  :  255 - 0xff -- Background 0xd3
    "11111111", -- 1689 - 0x699  :  255 - 0xff
    "11111111", -- 1690 - 0x69a  :  255 - 0xff
    "11111111", -- 1691 - 0x69b  :  255 - 0xff
    "11111101", -- 1692 - 0x69c  :  253 - 0xfd
    "11111101", -- 1693 - 0x69d  :  253 - 0xfd
    "11111101", -- 1694 - 0x69e  :  253 - 0xfd
    "11111101", -- 1695 - 0x69f  :  253 - 0xfd
    "00000111", -- 1696 - 0x6a0  :    7 - 0x7 -- Background 0xd4
    "00000111", -- 1697 - 0x6a1  :    7 - 0x7
    "00000000", -- 1698 - 0x6a2  :    0 - 0x0
    "00000011", -- 1699 - 0x6a3  :    3 - 0x3
    "00000000", -- 1700 - 0x6a4  :    0 - 0x0
    "00000000", -- 1701 - 0x6a5  :    0 - 0x0
    "00000000", -- 1702 - 0x6a6  :    0 - 0x0
    "00000000", -- 1703 - 0x6a7  :    0 - 0x0
    "11111010", -- 1704 - 0x6a8  :  250 - 0xfa -- Background 0xd5
    "11111010", -- 1705 - 0x6a9  :  250 - 0xfa
    "00000010", -- 1706 - 0x6aa  :    2 - 0x2
    "11111110", -- 1707 - 0x6ab  :  254 - 0xfe
    "00000000", -- 1708 - 0x6ac  :    0 - 0x0
    "00000000", -- 1709 - 0x6ad  :    0 - 0x0
    "00000000", -- 1710 - 0x6ae  :    0 - 0x0
    "00000000", -- 1711 - 0x6af  :    0 - 0x0
    "00001111", -- 1712 - 0x6b0  :   15 - 0xf -- Background 0xd6
    "00001111", -- 1713 - 0x6b1  :   15 - 0xf
    "00000000", -- 1714 - 0x6b2  :    0 - 0x0
    "00000111", -- 1715 - 0x6b3  :    7 - 0x7
    "00000000", -- 1716 - 0x6b4  :    0 - 0x0
    "00000000", -- 1717 - 0x6b5  :    0 - 0x0
    "00000000", -- 1718 - 0x6b6  :    0 - 0x0
    "00000000", -- 1719 - 0x6b7  :    0 - 0x0
    "11111111", -- 1720 - 0x6b8  :  255 - 0xff -- Background 0xd7
    "11111111", -- 1721 - 0x6b9  :  255 - 0xff
    "00000000", -- 1722 - 0x6ba  :    0 - 0x0
    "11111111", -- 1723 - 0x6bb  :  255 - 0xff
    "00000000", -- 1724 - 0x6bc  :    0 - 0x0
    "00000000", -- 1725 - 0x6bd  :    0 - 0x0
    "00000000", -- 1726 - 0x6be  :    0 - 0x0
    "00000000", -- 1727 - 0x6bf  :    0 - 0x0
    "11000011", -- 1728 - 0x6c0  :  195 - 0xc3 -- Background 0xd8
    "11111111", -- 1729 - 0x6c1  :  255 - 0xff
    "00000000", -- 1730 - 0x6c2  :    0 - 0x0
    "11111111", -- 1731 - 0x6c3  :  255 - 0xff
    "00000000", -- 1732 - 0x6c4  :    0 - 0x0
    "00000000", -- 1733 - 0x6c5  :    0 - 0x0
    "00000000", -- 1734 - 0x6c6  :    0 - 0x0
    "00000000", -- 1735 - 0x6c7  :    0 - 0x0
    "01101011", -- 1736 - 0x6c8  :  107 - 0x6b -- Background 0xd9
    "10110101", -- 1737 - 0x6c9  :  181 - 0xb5
    "00110110", -- 1738 - 0x6ca  :   54 - 0x36
    "11111000", -- 1739 - 0x6cb  :  248 - 0xf8
    "00000000", -- 1740 - 0x6cc  :    0 - 0x0
    "00000000", -- 1741 - 0x6cd  :    0 - 0x0
    "00000000", -- 1742 - 0x6ce  :    0 - 0x0
    "00000000", -- 1743 - 0x6cf  :    0 - 0x0
    "11111111", -- 1744 - 0x6d0  :  255 - 0xff -- Background 0xda
    "11111111", -- 1745 - 0x6d1  :  255 - 0xff
    "01111110", -- 1746 - 0x6d2  :  126 - 0x7e
    "10000001", -- 1747 - 0x6d3  :  129 - 0x81
    "00011111", -- 1748 - 0x6d4  :   31 - 0x1f
    "00000000", -- 1749 - 0x6d5  :    0 - 0x0
    "00000000", -- 1750 - 0x6d6  :    0 - 0x0
    "00000000", -- 1751 - 0x6d7  :    0 - 0x0
    "01101100", -- 1752 - 0x6d8  :  108 - 0x6c -- Background 0xdb
    "11011000", -- 1753 - 0x6d9  :  216 - 0xd8
    "00110000", -- 1754 - 0x6da  :   48 - 0x30
    "11100000", -- 1755 - 0x6db  :  224 - 0xe0
    "10000000", -- 1756 - 0x6dc  :  128 - 0x80
    "00000000", -- 1757 - 0x6dd  :    0 - 0x0
    "00000000", -- 1758 - 0x6de  :    0 - 0x0
    "00000000", -- 1759 - 0x6df  :    0 - 0x0
    "00011111", -- 1760 - 0x6e0  :   31 - 0x1f -- Background 0xdc
    "00011111", -- 1761 - 0x6e1  :   31 - 0x1f
    "00000000", -- 1762 - 0x6e2  :    0 - 0x0
    "00000111", -- 1763 - 0x6e3  :    7 - 0x7
    "00000000", -- 1764 - 0x6e4  :    0 - 0x0
    "00000000", -- 1765 - 0x6e5  :    0 - 0x0
    "00000000", -- 1766 - 0x6e6  :    0 - 0x0
    "00000000", -- 1767 - 0x6e7  :    0 - 0x0
    "10000101", -- 1768 - 0x6e8  :  133 - 0x85 -- Background 0xdd
    "11111101", -- 1769 - 0x6e9  :  253 - 0xfd
    "00000001", -- 1770 - 0x6ea  :    1 - 0x1
    "11111111", -- 1771 - 0x6eb  :  255 - 0xff
    "00000000", -- 1772 - 0x6ec  :    0 - 0x0
    "00000000", -- 1773 - 0x6ed  :    0 - 0x0
    "00000000", -- 1774 - 0x6ee  :    0 - 0x0
    "00000000", -- 1775 - 0x6ef  :    0 - 0x0
    "01111111", -- 1776 - 0x6f0  :  127 - 0x7f -- Background 0xde
    "01111111", -- 1777 - 0x6f1  :  127 - 0x7f
    "00000000", -- 1778 - 0x6f2  :    0 - 0x0
    "01011111", -- 1779 - 0x6f3  :   95 - 0x5f
    "00000000", -- 1780 - 0x6f4  :    0 - 0x0
    "00000000", -- 1781 - 0x6f5  :    0 - 0x0
    "00000000", -- 1782 - 0x6f6  :    0 - 0x0
    "00000000", -- 1783 - 0x6f7  :    0 - 0x0
    "11111100", -- 1784 - 0x6f8  :  252 - 0xfc -- Background 0xdf
    "11111111", -- 1785 - 0x6f9  :  255 - 0xff
    "00000000", -- 1786 - 0x6fa  :    0 - 0x0
    "11111111", -- 1787 - 0x6fb  :  255 - 0xff
    "00000000", -- 1788 - 0x6fc  :    0 - 0x0
    "00000000", -- 1789 - 0x6fd  :    0 - 0x0
    "00000000", -- 1790 - 0x6fe  :    0 - 0x0
    "00000000", -- 1791 - 0x6ff  :    0 - 0x0
    "00110100", -- 1792 - 0x700  :   52 - 0x34 -- Background 0xe0
    "11110110", -- 1793 - 0x701  :  246 - 0xf6
    "00000010", -- 1794 - 0x702  :    2 - 0x2
    "11111111", -- 1795 - 0x703  :  255 - 0xff
    "00000000", -- 1796 - 0x704  :    0 - 0x0
    "00000000", -- 1797 - 0x705  :    0 - 0x0
    "00000000", -- 1798 - 0x706  :    0 - 0x0
    "00000000", -- 1799 - 0x707  :    0 - 0x0
    "11111111", -- 1800 - 0x708  :  255 - 0xff -- Background 0xe1
    "11111111", -- 1801 - 0x709  :  255 - 0xff
    "00000000", -- 1802 - 0x70a  :    0 - 0x0
    "01111111", -- 1803 - 0x70b  :  127 - 0x7f
    "00000000", -- 1804 - 0x70c  :    0 - 0x0
    "00000000", -- 1805 - 0x70d  :    0 - 0x0
    "00000000", -- 1806 - 0x70e  :    0 - 0x0
    "00000000", -- 1807 - 0x70f  :    0 - 0x0
    "11100001", -- 1808 - 0x710  :  225 - 0xe1 -- Background 0xe2
    "11111111", -- 1809 - 0x711  :  255 - 0xff
    "00000000", -- 1810 - 0x712  :    0 - 0x0
    "11111111", -- 1811 - 0x713  :  255 - 0xff
    "00000000", -- 1812 - 0x714  :    0 - 0x0
    "00000000", -- 1813 - 0x715  :    0 - 0x0
    "00000000", -- 1814 - 0x716  :    0 - 0x0
    "00000000", -- 1815 - 0x717  :    0 - 0x0
    "01000000", -- 1816 - 0x718  :   64 - 0x40 -- Background 0xe3
    "01000000", -- 1817 - 0x719  :   64 - 0x40
    "01000000", -- 1818 - 0x71a  :   64 - 0x40
    "11000000", -- 1819 - 0x71b  :  192 - 0xc0
    "00000000", -- 1820 - 0x71c  :    0 - 0x0
    "00000000", -- 1821 - 0x71d  :    0 - 0x0
    "00000000", -- 1822 - 0x71e  :    0 - 0x0
    "00000000", -- 1823 - 0x71f  :    0 - 0x0
    "00000000", -- 1824 - 0x720  :    0 - 0x0 -- Background 0xe4
    "00000000", -- 1825 - 0x721  :    0 - 0x0
    "00000000", -- 1826 - 0x722  :    0 - 0x0
    "00000000", -- 1827 - 0x723  :    0 - 0x0
    "00000111", -- 1828 - 0x724  :    7 - 0x7
    "00001111", -- 1829 - 0x725  :   15 - 0xf
    "00001111", -- 1830 - 0x726  :   15 - 0xf
    "00001111", -- 1831 - 0x727  :   15 - 0xf
    "00000000", -- 1832 - 0x728  :    0 - 0x0 -- Background 0xe5
    "00000000", -- 1833 - 0x729  :    0 - 0x0
    "00000000", -- 1834 - 0x72a  :    0 - 0x0
    "00000000", -- 1835 - 0x72b  :    0 - 0x0
    "11100000", -- 1836 - 0x72c  :  224 - 0xe0
    "11110000", -- 1837 - 0x72d  :  240 - 0xf0
    "11110000", -- 1838 - 0x72e  :  240 - 0xf0
    "11110000", -- 1839 - 0x72f  :  240 - 0xf0
    "11110000", -- 1840 - 0x730  :  240 - 0xf0 -- Background 0xe6
    "11110000", -- 1841 - 0x731  :  240 - 0xf0
    "11110000", -- 1842 - 0x732  :  240 - 0xf0
    "11100000", -- 1843 - 0x733  :  224 - 0xe0
    "00000000", -- 1844 - 0x734  :    0 - 0x0
    "00000000", -- 1845 - 0x735  :    0 - 0x0
    "00000000", -- 1846 - 0x736  :    0 - 0x0
    "00000000", -- 1847 - 0x737  :    0 - 0x0
    "00001111", -- 1848 - 0x738  :   15 - 0xf -- Background 0xe7
    "00001111", -- 1849 - 0x739  :   15 - 0xf
    "00001111", -- 1850 - 0x73a  :   15 - 0xf
    "00000111", -- 1851 - 0x73b  :    7 - 0x7
    "00000000", -- 1852 - 0x73c  :    0 - 0x0
    "00000000", -- 1853 - 0x73d  :    0 - 0x0
    "00000000", -- 1854 - 0x73e  :    0 - 0x0
    "00000000", -- 1855 - 0x73f  :    0 - 0x0
    "00000000", -- 1856 - 0x740  :    0 - 0x0 -- Background 0xe8
    "00000000", -- 1857 - 0x741  :    0 - 0x0
    "00000000", -- 1858 - 0x742  :    0 - 0x0
    "00000000", -- 1859 - 0x743  :    0 - 0x0
    "11111111", -- 1860 - 0x744  :  255 - 0xff
    "11111111", -- 1861 - 0x745  :  255 - 0xff
    "11111111", -- 1862 - 0x746  :  255 - 0xff
    "11111111", -- 1863 - 0x747  :  255 - 0xff
    "11110000", -- 1864 - 0x748  :  240 - 0xf0 -- Background 0xe9
    "11110000", -- 1865 - 0x749  :  240 - 0xf0
    "11110000", -- 1866 - 0x74a  :  240 - 0xf0
    "11110000", -- 1867 - 0x74b  :  240 - 0xf0
    "11110000", -- 1868 - 0x74c  :  240 - 0xf0
    "11110000", -- 1869 - 0x74d  :  240 - 0xf0
    "11110000", -- 1870 - 0x74e  :  240 - 0xf0
    "11110000", -- 1871 - 0x74f  :  240 - 0xf0
    "11111111", -- 1872 - 0x750  :  255 - 0xff -- Background 0xea
    "11111111", -- 1873 - 0x751  :  255 - 0xff
    "11111111", -- 1874 - 0x752  :  255 - 0xff
    "11111111", -- 1875 - 0x753  :  255 - 0xff
    "00000000", -- 1876 - 0x754  :    0 - 0x0
    "00000000", -- 1877 - 0x755  :    0 - 0x0
    "00000000", -- 1878 - 0x756  :    0 - 0x0
    "00000000", -- 1879 - 0x757  :    0 - 0x0
    "00001111", -- 1880 - 0x758  :   15 - 0xf -- Background 0xeb
    "00001111", -- 1881 - 0x759  :   15 - 0xf
    "00001111", -- 1882 - 0x75a  :   15 - 0xf
    "00001111", -- 1883 - 0x75b  :   15 - 0xf
    "00001111", -- 1884 - 0x75c  :   15 - 0xf
    "00001111", -- 1885 - 0x75d  :   15 - 0xf
    "00001111", -- 1886 - 0x75e  :   15 - 0xf
    "00001111", -- 1887 - 0x75f  :   15 - 0xf
    "00000000", -- 1888 - 0x760  :    0 - 0x0 -- Background 0xec
    "00000000", -- 1889 - 0x761  :    0 - 0x0
    "00000000", -- 1890 - 0x762  :    0 - 0x0
    "00000000", -- 1891 - 0x763  :    0 - 0x0
    "00000000", -- 1892 - 0x764  :    0 - 0x0
    "00000000", -- 1893 - 0x765  :    0 - 0x0
    "00000000", -- 1894 - 0x766  :    0 - 0x0
    "00000000", -- 1895 - 0x767  :    0 - 0x0
    "00000000", -- 1896 - 0x768  :    0 - 0x0 -- Background 0xed
    "00000000", -- 1897 - 0x769  :    0 - 0x0
    "00000000", -- 1898 - 0x76a  :    0 - 0x0
    "00000000", -- 1899 - 0x76b  :    0 - 0x0
    "00000000", -- 1900 - 0x76c  :    0 - 0x0
    "00000000", -- 1901 - 0x76d  :    0 - 0x0
    "00000000", -- 1902 - 0x76e  :    0 - 0x0
    "00000000", -- 1903 - 0x76f  :    0 - 0x0
    "00000000", -- 1904 - 0x770  :    0 - 0x0 -- Background 0xee
    "00000000", -- 1905 - 0x771  :    0 - 0x0
    "00000000", -- 1906 - 0x772  :    0 - 0x0
    "00000000", -- 1907 - 0x773  :    0 - 0x0
    "00000000", -- 1908 - 0x774  :    0 - 0x0
    "00000000", -- 1909 - 0x775  :    0 - 0x0
    "00000000", -- 1910 - 0x776  :    0 - 0x0
    "00000000", -- 1911 - 0x777  :    0 - 0x0
    "00000000", -- 1912 - 0x778  :    0 - 0x0 -- Background 0xef
    "00000000", -- 1913 - 0x779  :    0 - 0x0
    "00000000", -- 1914 - 0x77a  :    0 - 0x0
    "00000000", -- 1915 - 0x77b  :    0 - 0x0
    "00000000", -- 1916 - 0x77c  :    0 - 0x0
    "00000000", -- 1917 - 0x77d  :    0 - 0x0
    "00000000", -- 1918 - 0x77e  :    0 - 0x0
    "00000000", -- 1919 - 0x77f  :    0 - 0x0
    "11111111", -- 1920 - 0x780  :  255 - 0xff -- Background 0xf0
    "11111111", -- 1921 - 0x781  :  255 - 0xff
    "11111111", -- 1922 - 0x782  :  255 - 0xff
    "11111111", -- 1923 - 0x783  :  255 - 0xff
    "11111111", -- 1924 - 0x784  :  255 - 0xff
    "11111111", -- 1925 - 0x785  :  255 - 0xff
    "11111111", -- 1926 - 0x786  :  255 - 0xff
    "11111111", -- 1927 - 0x787  :  255 - 0xff
    "11111111", -- 1928 - 0x788  :  255 - 0xff -- Background 0xf1
    "11111111", -- 1929 - 0x789  :  255 - 0xff
    "11111111", -- 1930 - 0x78a  :  255 - 0xff
    "11111111", -- 1931 - 0x78b  :  255 - 0xff
    "11111111", -- 1932 - 0x78c  :  255 - 0xff
    "11111111", -- 1933 - 0x78d  :  255 - 0xff
    "11111111", -- 1934 - 0x78e  :  255 - 0xff
    "11111111", -- 1935 - 0x78f  :  255 - 0xff
    "11111111", -- 1936 - 0x790  :  255 - 0xff -- Background 0xf2
    "11111111", -- 1937 - 0x791  :  255 - 0xff
    "11111111", -- 1938 - 0x792  :  255 - 0xff
    "11111111", -- 1939 - 0x793  :  255 - 0xff
    "11111111", -- 1940 - 0x794  :  255 - 0xff
    "11111111", -- 1941 - 0x795  :  255 - 0xff
    "11111111", -- 1942 - 0x796  :  255 - 0xff
    "11111111", -- 1943 - 0x797  :  255 - 0xff
    "11111111", -- 1944 - 0x798  :  255 - 0xff -- Background 0xf3
    "11111111", -- 1945 - 0x799  :  255 - 0xff
    "11111111", -- 1946 - 0x79a  :  255 - 0xff
    "11111111", -- 1947 - 0x79b  :  255 - 0xff
    "11111111", -- 1948 - 0x79c  :  255 - 0xff
    "11111111", -- 1949 - 0x79d  :  255 - 0xff
    "11111111", -- 1950 - 0x79e  :  255 - 0xff
    "11111111", -- 1951 - 0x79f  :  255 - 0xff
    "11111111", -- 1952 - 0x7a0  :  255 - 0xff -- Background 0xf4
    "11111111", -- 1953 - 0x7a1  :  255 - 0xff
    "11111111", -- 1954 - 0x7a2  :  255 - 0xff
    "11111111", -- 1955 - 0x7a3  :  255 - 0xff
    "11111111", -- 1956 - 0x7a4  :  255 - 0xff
    "11111111", -- 1957 - 0x7a5  :  255 - 0xff
    "11111111", -- 1958 - 0x7a6  :  255 - 0xff
    "11111111", -- 1959 - 0x7a7  :  255 - 0xff
    "11111111", -- 1960 - 0x7a8  :  255 - 0xff -- Background 0xf5
    "11111111", -- 1961 - 0x7a9  :  255 - 0xff
    "11111111", -- 1962 - 0x7aa  :  255 - 0xff
    "11111111", -- 1963 - 0x7ab  :  255 - 0xff
    "11111111", -- 1964 - 0x7ac  :  255 - 0xff
    "11111111", -- 1965 - 0x7ad  :  255 - 0xff
    "11111111", -- 1966 - 0x7ae  :  255 - 0xff
    "11111111", -- 1967 - 0x7af  :  255 - 0xff
    "11111111", -- 1968 - 0x7b0  :  255 - 0xff -- Background 0xf6
    "11111111", -- 1969 - 0x7b1  :  255 - 0xff
    "11111111", -- 1970 - 0x7b2  :  255 - 0xff
    "11111111", -- 1971 - 0x7b3  :  255 - 0xff
    "11111111", -- 1972 - 0x7b4  :  255 - 0xff
    "11111111", -- 1973 - 0x7b5  :  255 - 0xff
    "11111111", -- 1974 - 0x7b6  :  255 - 0xff
    "11111111", -- 1975 - 0x7b7  :  255 - 0xff
    "11111111", -- 1976 - 0x7b8  :  255 - 0xff -- Background 0xf7
    "11111111", -- 1977 - 0x7b9  :  255 - 0xff
    "11111111", -- 1978 - 0x7ba  :  255 - 0xff
    "11111111", -- 1979 - 0x7bb  :  255 - 0xff
    "11111111", -- 1980 - 0x7bc  :  255 - 0xff
    "11111111", -- 1981 - 0x7bd  :  255 - 0xff
    "11111111", -- 1982 - 0x7be  :  255 - 0xff
    "11111111", -- 1983 - 0x7bf  :  255 - 0xff
    "11111111", -- 1984 - 0x7c0  :  255 - 0xff -- Background 0xf8
    "11111111", -- 1985 - 0x7c1  :  255 - 0xff
    "11111111", -- 1986 - 0x7c2  :  255 - 0xff
    "11111111", -- 1987 - 0x7c3  :  255 - 0xff
    "11111111", -- 1988 - 0x7c4  :  255 - 0xff
    "11111111", -- 1989 - 0x7c5  :  255 - 0xff
    "11111111", -- 1990 - 0x7c6  :  255 - 0xff
    "11111111", -- 1991 - 0x7c7  :  255 - 0xff
    "11111111", -- 1992 - 0x7c8  :  255 - 0xff -- Background 0xf9
    "11111111", -- 1993 - 0x7c9  :  255 - 0xff
    "11111111", -- 1994 - 0x7ca  :  255 - 0xff
    "11111111", -- 1995 - 0x7cb  :  255 - 0xff
    "11111111", -- 1996 - 0x7cc  :  255 - 0xff
    "11111111", -- 1997 - 0x7cd  :  255 - 0xff
    "11111111", -- 1998 - 0x7ce  :  255 - 0xff
    "11111111", -- 1999 - 0x7cf  :  255 - 0xff
    "11111111", -- 2000 - 0x7d0  :  255 - 0xff -- Background 0xfa
    "11111111", -- 2001 - 0x7d1  :  255 - 0xff
    "11111111", -- 2002 - 0x7d2  :  255 - 0xff
    "11111111", -- 2003 - 0x7d3  :  255 - 0xff
    "11111111", -- 2004 - 0x7d4  :  255 - 0xff
    "11111111", -- 2005 - 0x7d5  :  255 - 0xff
    "11111111", -- 2006 - 0x7d6  :  255 - 0xff
    "11111111", -- 2007 - 0x7d7  :  255 - 0xff
    "11111111", -- 2008 - 0x7d8  :  255 - 0xff -- Background 0xfb
    "11111111", -- 2009 - 0x7d9  :  255 - 0xff
    "11111111", -- 2010 - 0x7da  :  255 - 0xff
    "11111111", -- 2011 - 0x7db  :  255 - 0xff
    "11111111", -- 2012 - 0x7dc  :  255 - 0xff
    "11111111", -- 2013 - 0x7dd  :  255 - 0xff
    "11111111", -- 2014 - 0x7de  :  255 - 0xff
    "11111111", -- 2015 - 0x7df  :  255 - 0xff
    "11111111", -- 2016 - 0x7e0  :  255 - 0xff -- Background 0xfc
    "11111111", -- 2017 - 0x7e1  :  255 - 0xff
    "11111111", -- 2018 - 0x7e2  :  255 - 0xff
    "11111111", -- 2019 - 0x7e3  :  255 - 0xff
    "11111111", -- 2020 - 0x7e4  :  255 - 0xff
    "11111111", -- 2021 - 0x7e5  :  255 - 0xff
    "11111111", -- 2022 - 0x7e6  :  255 - 0xff
    "11111111", -- 2023 - 0x7e7  :  255 - 0xff
    "11111111", -- 2024 - 0x7e8  :  255 - 0xff -- Background 0xfd
    "11111111", -- 2025 - 0x7e9  :  255 - 0xff
    "11111111", -- 2026 - 0x7ea  :  255 - 0xff
    "11111111", -- 2027 - 0x7eb  :  255 - 0xff
    "11111111", -- 2028 - 0x7ec  :  255 - 0xff
    "11111111", -- 2029 - 0x7ed  :  255 - 0xff
    "11111111", -- 2030 - 0x7ee  :  255 - 0xff
    "11111111", -- 2031 - 0x7ef  :  255 - 0xff
    "11111111", -- 2032 - 0x7f0  :  255 - 0xff -- Background 0xfe
    "11111111", -- 2033 - 0x7f1  :  255 - 0xff
    "11111111", -- 2034 - 0x7f2  :  255 - 0xff
    "11111111", -- 2035 - 0x7f3  :  255 - 0xff
    "11111111", -- 2036 - 0x7f4  :  255 - 0xff
    "11111111", -- 2037 - 0x7f5  :  255 - 0xff
    "11111111", -- 2038 - 0x7f6  :  255 - 0xff
    "11111111", -- 2039 - 0x7f7  :  255 - 0xff
    "11111111", -- 2040 - 0x7f8  :  255 - 0xff -- Background 0xff
    "11111111", -- 2041 - 0x7f9  :  255 - 0xff
    "11111111", -- 2042 - 0x7fa  :  255 - 0xff
    "11111111", -- 2043 - 0x7fb  :  255 - 0xff
    "11111111", -- 2044 - 0x7fc  :  255 - 0xff
    "11111111", -- 2045 - 0x7fd  :  255 - 0xff
    "11111111", -- 2046 - 0x7fe  :  255 - 0xff
    "11111111"  -- 2047 - 0x7ff  :  255 - 0xff
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
