--- Autcmatically generated VHDL ROM from a NES memory file----
---   PATTERN TABLE WITH ONLY ONE COLOR PLANE
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


---  Original memory dump file name: pacman_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_PACMAN_color0 is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(12-1 downto 0);  --4096 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_PACMAN_color0;

architecture BEHAVIORAL of ROM_PTABLE_PACMAN_color0 is
  signal addr_int  : natural range 0 to 2**12-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Sprite pattern Table
    "00000000", --    0 -  0x0  :    0 - 0x0 -- Sprite 0x0
    "00000000", --    1 -  0x1  :    0 - 0x0
    "00000000", --    2 -  0x2  :    0 - 0x0
    "00000000", --    3 -  0x3  :    0 - 0x0
    "00000000", --    4 -  0x4  :    0 - 0x0
    "00000000", --    5 -  0x5  :    0 - 0x0
    "00000000", --    6 -  0x6  :    0 - 0x0
    "00000000", --    7 -  0x7  :    0 - 0x0
    "00000000", --    8 -  0x8  :    0 - 0x0 -- Sprite 0x1
    "00111000", --    9 -  0x9  :   56 - 0x38
    "01111100", --   10 -  0xa  :  124 - 0x7c
    "11111110", --   11 -  0xb  :  254 - 0xfe
    "11111110", --   12 -  0xc  :  254 - 0xfe
    "11111110", --   13 -  0xd  :  254 - 0xfe
    "01111100", --   14 -  0xe  :  124 - 0x7c
    "00111000", --   15 -  0xf  :   56 - 0x38
    "00000000", --   16 - 0x10  :    0 - 0x0 -- Sprite 0x2
    "00000000", --   17 - 0x11  :    0 - 0x0
    "00000000", --   18 - 0x12  :    0 - 0x0
    "00000000", --   19 - 0x13  :    0 - 0x0
    "00000000", --   20 - 0x14  :    0 - 0x0
    "00000000", --   21 - 0x15  :    0 - 0x0
    "00000000", --   22 - 0x16  :    0 - 0x0
    "00000000", --   23 - 0x17  :    0 - 0x0
    "00000000", --   24 - 0x18  :    0 - 0x0 -- Sprite 0x3
    "00000000", --   25 - 0x19  :    0 - 0x0
    "00000000", --   26 - 0x1a  :    0 - 0x0
    "00011000", --   27 - 0x1b  :   24 - 0x18
    "00011000", --   28 - 0x1c  :   24 - 0x18
    "00000000", --   29 - 0x1d  :    0 - 0x0
    "00000000", --   30 - 0x1e  :    0 - 0x0
    "00000000", --   31 - 0x1f  :    0 - 0x0
    "00000000", --   32 - 0x20  :    0 - 0x0 -- Sprite 0x4
    "00000000", --   33 - 0x21  :    0 - 0x0
    "00000000", --   34 - 0x22  :    0 - 0x0
    "00000000", --   35 - 0x23  :    0 - 0x0
    "00000000", --   36 - 0x24  :    0 - 0x0
    "00000000", --   37 - 0x25  :    0 - 0x0
    "00000000", --   38 - 0x26  :    0 - 0x0
    "00000000", --   39 - 0x27  :    0 - 0x0
    "00000000", --   40 - 0x28  :    0 - 0x0 -- Sprite 0x5
    "00000000", --   41 - 0x29  :    0 - 0x0
    "00000000", --   42 - 0x2a  :    0 - 0x0
    "00000000", --   43 - 0x2b  :    0 - 0x0
    "00000000", --   44 - 0x2c  :    0 - 0x0
    "00000000", --   45 - 0x2d  :    0 - 0x0
    "00000000", --   46 - 0x2e  :    0 - 0x0
    "00000000", --   47 - 0x2f  :    0 - 0x0
    "00000000", --   48 - 0x30  :    0 - 0x0 -- Sprite 0x6
    "00000000", --   49 - 0x31  :    0 - 0x0
    "00000000", --   50 - 0x32  :    0 - 0x0
    "00000000", --   51 - 0x33  :    0 - 0x0
    "00000000", --   52 - 0x34  :    0 - 0x0
    "00000000", --   53 - 0x35  :    0 - 0x0
    "00000000", --   54 - 0x36  :    0 - 0x0
    "00000000", --   55 - 0x37  :    0 - 0x0
    "00000000", --   56 - 0x38  :    0 - 0x0 -- Sprite 0x7
    "00000000", --   57 - 0x39  :    0 - 0x0
    "00000000", --   58 - 0x3a  :    0 - 0x0
    "00000000", --   59 - 0x3b  :    0 - 0x0
    "00000000", --   60 - 0x3c  :    0 - 0x0
    "00000000", --   61 - 0x3d  :    0 - 0x0
    "00000000", --   62 - 0x3e  :    0 - 0x0
    "00000000", --   63 - 0x3f  :    0 - 0x0
    "00000000", --   64 - 0x40  :    0 - 0x0 -- Sprite 0x8
    "00000000", --   65 - 0x41  :    0 - 0x0
    "00000000", --   66 - 0x42  :    0 - 0x0
    "00000000", --   67 - 0x43  :    0 - 0x0
    "00000000", --   68 - 0x44  :    0 - 0x0
    "00000000", --   69 - 0x45  :    0 - 0x0
    "00000000", --   70 - 0x46  :    0 - 0x0
    "00000000", --   71 - 0x47  :    0 - 0x0
    "00000000", --   72 - 0x48  :    0 - 0x0 -- Sprite 0x9
    "00000000", --   73 - 0x49  :    0 - 0x0
    "00000000", --   74 - 0x4a  :    0 - 0x0
    "00011000", --   75 - 0x4b  :   24 - 0x18
    "00011000", --   76 - 0x4c  :   24 - 0x18
    "00000000", --   77 - 0x4d  :    0 - 0x0
    "00000000", --   78 - 0x4e  :    0 - 0x0
    "00000000", --   79 - 0x4f  :    0 - 0x0
    "00000000", --   80 - 0x50  :    0 - 0x0 -- Sprite 0xa
    "00000000", --   81 - 0x51  :    0 - 0x0
    "00000000", --   82 - 0x52  :    0 - 0x0
    "00000000", --   83 - 0x53  :    0 - 0x0
    "00000000", --   84 - 0x54  :    0 - 0x0
    "00000000", --   85 - 0x55  :    0 - 0x0
    "00000000", --   86 - 0x56  :    0 - 0x0
    "00000000", --   87 - 0x57  :    0 - 0x0
    "00000000", --   88 - 0x58  :    0 - 0x0 -- Sprite 0xb
    "00000000", --   89 - 0x59  :    0 - 0x0
    "00000000", --   90 - 0x5a  :    0 - 0x0
    "00000000", --   91 - 0x5b  :    0 - 0x0
    "00000000", --   92 - 0x5c  :    0 - 0x0
    "00000000", --   93 - 0x5d  :    0 - 0x0
    "00000000", --   94 - 0x5e  :    0 - 0x0
    "00000000", --   95 - 0x5f  :    0 - 0x0
    "00000000", --   96 - 0x60  :    0 - 0x0 -- Sprite 0xc
    "00000000", --   97 - 0x61  :    0 - 0x0
    "00000000", --   98 - 0x62  :    0 - 0x0
    "00000000", --   99 - 0x63  :    0 - 0x0
    "00000000", --  100 - 0x64  :    0 - 0x0
    "00000000", --  101 - 0x65  :    0 - 0x0
    "00000000", --  102 - 0x66  :    0 - 0x0
    "00000000", --  103 - 0x67  :    0 - 0x0
    "00000000", --  104 - 0x68  :    0 - 0x0 -- Sprite 0xd
    "00000000", --  105 - 0x69  :    0 - 0x0
    "00000000", --  106 - 0x6a  :    0 - 0x0
    "00000000", --  107 - 0x6b  :    0 - 0x0
    "00000000", --  108 - 0x6c  :    0 - 0x0
    "00000000", --  109 - 0x6d  :    0 - 0x0
    "00000000", --  110 - 0x6e  :    0 - 0x0
    "00000000", --  111 - 0x6f  :    0 - 0x0
    "00000000", --  112 - 0x70  :    0 - 0x0 -- Sprite 0xe
    "00000000", --  113 - 0x71  :    0 - 0x0
    "00000000", --  114 - 0x72  :    0 - 0x0
    "00000000", --  115 - 0x73  :    0 - 0x0
    "00000000", --  116 - 0x74  :    0 - 0x0
    "00000000", --  117 - 0x75  :    0 - 0x0
    "00000000", --  118 - 0x76  :    0 - 0x0
    "00000000", --  119 - 0x77  :    0 - 0x0
    "00000000", --  120 - 0x78  :    0 - 0x0 -- Sprite 0xf
    "00000000", --  121 - 0x79  :    0 - 0x0
    "00000000", --  122 - 0x7a  :    0 - 0x0
    "00000000", --  123 - 0x7b  :    0 - 0x0
    "00000000", --  124 - 0x7c  :    0 - 0x0
    "00000000", --  125 - 0x7d  :    0 - 0x0
    "00000000", --  126 - 0x7e  :    0 - 0x0
    "00000000", --  127 - 0x7f  :    0 - 0x0
    "00000000", --  128 - 0x80  :    0 - 0x0 -- Sprite 0x10
    "00000000", --  129 - 0x81  :    0 - 0x0
    "11111111", --  130 - 0x82  :  255 - 0xff
    "00000000", --  131 - 0x83  :    0 - 0x0
    "00000000", --  132 - 0x84  :    0 - 0x0
    "11111111", --  133 - 0x85  :  255 - 0xff
    "00000000", --  134 - 0x86  :    0 - 0x0
    "00000000", --  135 - 0x87  :    0 - 0x0
    "00100100", --  136 - 0x88  :   36 - 0x24 -- Sprite 0x11
    "00100100", --  137 - 0x89  :   36 - 0x24
    "00100100", --  138 - 0x8a  :   36 - 0x24
    "00100100", --  139 - 0x8b  :   36 - 0x24
    "00100100", --  140 - 0x8c  :   36 - 0x24
    "00100100", --  141 - 0x8d  :   36 - 0x24
    "00100100", --  142 - 0x8e  :   36 - 0x24
    "00100100", --  143 - 0x8f  :   36 - 0x24
    "00100100", --  144 - 0x90  :   36 - 0x24 -- Sprite 0x12
    "00100100", --  145 - 0x91  :   36 - 0x24
    "11000011", --  146 - 0x92  :  195 - 0xc3
    "00000000", --  147 - 0x93  :    0 - 0x0
    "00000000", --  148 - 0x94  :    0 - 0x0
    "11111111", --  149 - 0x95  :  255 - 0xff
    "00000000", --  150 - 0x96  :    0 - 0x0
    "00000000", --  151 - 0x97  :    0 - 0x0
    "00000000", --  152 - 0x98  :    0 - 0x0 -- Sprite 0x13
    "00000000", --  153 - 0x99  :    0 - 0x0
    "11111111", --  154 - 0x9a  :  255 - 0xff
    "00000000", --  155 - 0x9b  :    0 - 0x0
    "00000000", --  156 - 0x9c  :    0 - 0x0
    "11000011", --  157 - 0x9d  :  195 - 0xc3
    "00100100", --  158 - 0x9e  :   36 - 0x24
    "00100100", --  159 - 0x9f  :   36 - 0x24
    "00100100", --  160 - 0xa0  :   36 - 0x24 -- Sprite 0x14
    "00100100", --  161 - 0xa1  :   36 - 0x24
    "11000100", --  162 - 0xa2  :  196 - 0xc4
    "00000100", --  163 - 0xa3  :    4 - 0x4
    "00000100", --  164 - 0xa4  :    4 - 0x4
    "11000100", --  165 - 0xa5  :  196 - 0xc4
    "00100100", --  166 - 0xa6  :   36 - 0x24
    "00100100", --  167 - 0xa7  :   36 - 0x24
    "00100100", --  168 - 0xa8  :   36 - 0x24 -- Sprite 0x15
    "00100100", --  169 - 0xa9  :   36 - 0x24
    "00100011", --  170 - 0xaa  :   35 - 0x23
    "00100000", --  171 - 0xab  :   32 - 0x20
    "00100000", --  172 - 0xac  :   32 - 0x20
    "00100011", --  173 - 0xad  :   35 - 0x23
    "00100100", --  174 - 0xae  :   36 - 0x24
    "00100100", --  175 - 0xaf  :   36 - 0x24
    "00000000", --  176 - 0xb0  :    0 - 0x0 -- Sprite 0x16
    "00000000", --  177 - 0xb1  :    0 - 0x0
    "00001111", --  178 - 0xb2  :   15 - 0xf
    "00010000", --  179 - 0xb3  :   16 - 0x10
    "11110000", --  180 - 0xb4  :  240 - 0xf0
    "00001111", --  181 - 0xb5  :   15 - 0xf
    "00000000", --  182 - 0xb6  :    0 - 0x0
    "00000000", --  183 - 0xb7  :    0 - 0x0
    "00000000", --  184 - 0xb8  :    0 - 0x0 -- Sprite 0x17
    "00000000", --  185 - 0xb9  :    0 - 0x0
    "11110000", --  186 - 0xba  :  240 - 0xf0
    "00001000", --  187 - 0xbb  :    8 - 0x8
    "00001111", --  188 - 0xbc  :   15 - 0xf
    "11110000", --  189 - 0xbd  :  240 - 0xf0
    "00000000", --  190 - 0xbe  :    0 - 0x0
    "00000000", --  191 - 0xbf  :    0 - 0x0
    "00000000", --  192 - 0xc0  :    0 - 0x0 -- Sprite 0x18
    "00000000", --  193 - 0xc1  :    0 - 0x0
    "11110000", --  194 - 0xc2  :  240 - 0xf0
    "00001000", --  195 - 0xc3  :    8 - 0x8
    "00001000", --  196 - 0xc4  :    8 - 0x8
    "11110000", --  197 - 0xc5  :  240 - 0xf0
    "00000000", --  198 - 0xc6  :    0 - 0x0
    "00000000", --  199 - 0xc7  :    0 - 0x0
    "00000000", --  200 - 0xc8  :    0 - 0x0 -- Sprite 0x19
    "00000000", --  201 - 0xc9  :    0 - 0x0
    "00001111", --  202 - 0xca  :   15 - 0xf
    "00010000", --  203 - 0xcb  :   16 - 0x10
    "00010000", --  204 - 0xcc  :   16 - 0x10
    "00001111", --  205 - 0xcd  :   15 - 0xf
    "00000000", --  206 - 0xce  :    0 - 0x0
    "00000000", --  207 - 0xcf  :    0 - 0x0
    "00100100", --  208 - 0xd0  :   36 - 0x24 -- Sprite 0x1a
    "00100100", --  209 - 0xd1  :   36 - 0x24
    "00100100", --  210 - 0xd2  :   36 - 0x24
    "00100100", --  211 - 0xd3  :   36 - 0x24
    "00011000", --  212 - 0xd4  :   24 - 0x18
    "00000000", --  213 - 0xd5  :    0 - 0x0
    "00000000", --  214 - 0xd6  :    0 - 0x0
    "00000000", --  215 - 0xd7  :    0 - 0x0
    "00000000", --  216 - 0xd8  :    0 - 0x0 -- Sprite 0x1b
    "00000000", --  217 - 0xd9  :    0 - 0x0
    "00000000", --  218 - 0xda  :    0 - 0x0
    "00011000", --  219 - 0xdb  :   24 - 0x18
    "00100100", --  220 - 0xdc  :   36 - 0x24
    "00100100", --  221 - 0xdd  :   36 - 0x24
    "00100100", --  222 - 0xde  :   36 - 0x24
    "00100100", --  223 - 0xdf  :   36 - 0x24
    "00100100", --  224 - 0xe0  :   36 - 0x24 -- Sprite 0x1c
    "00100100", --  225 - 0xe1  :   36 - 0x24
    "11000100", --  226 - 0xe2  :  196 - 0xc4
    "00000100", --  227 - 0xe3  :    4 - 0x4
    "00001000", --  228 - 0xe4  :    8 - 0x8
    "11110000", --  229 - 0xe5  :  240 - 0xf0
    "00000000", --  230 - 0xe6  :    0 - 0x0
    "00000000", --  231 - 0xe7  :    0 - 0x0
    "00000000", --  232 - 0xe8  :    0 - 0x0 -- Sprite 0x1d
    "00000000", --  233 - 0xe9  :    0 - 0x0
    "11110000", --  234 - 0xea  :  240 - 0xf0
    "00001000", --  235 - 0xeb  :    8 - 0x8
    "00000100", --  236 - 0xec  :    4 - 0x4
    "11000100", --  237 - 0xed  :  196 - 0xc4
    "00100100", --  238 - 0xee  :   36 - 0x24
    "00100100", --  239 - 0xef  :   36 - 0x24
    "00100100", --  240 - 0xf0  :   36 - 0x24 -- Sprite 0x1e
    "00100100", --  241 - 0xf1  :   36 - 0x24
    "00100011", --  242 - 0xf2  :   35 - 0x23
    "00100000", --  243 - 0xf3  :   32 - 0x20
    "00010000", --  244 - 0xf4  :   16 - 0x10
    "00001111", --  245 - 0xf5  :   15 - 0xf
    "00000000", --  246 - 0xf6  :    0 - 0x0
    "00000000", --  247 - 0xf7  :    0 - 0x0
    "00000000", --  248 - 0xf8  :    0 - 0x0 -- Sprite 0x1f
    "00000000", --  249 - 0xf9  :    0 - 0x0
    "00001111", --  250 - 0xfa  :   15 - 0xf
    "00010000", --  251 - 0xfb  :   16 - 0x10
    "00100000", --  252 - 0xfc  :   32 - 0x20
    "00100011", --  253 - 0xfd  :   35 - 0x23
    "00100100", --  254 - 0xfe  :   36 - 0x24
    "00100100", --  255 - 0xff  :   36 - 0x24
    "00000000", --  256 - 0x100  :    0 - 0x0 -- Sprite 0x20
    "00000000", --  257 - 0x101  :    0 - 0x0
    "00000000", --  258 - 0x102  :    0 - 0x0
    "00000000", --  259 - 0x103  :    0 - 0x0
    "00000000", --  260 - 0x104  :    0 - 0x0
    "00000000", --  261 - 0x105  :    0 - 0x0
    "00000000", --  262 - 0x106  :    0 - 0x0
    "00000000", --  263 - 0x107  :    0 - 0x0
    "00000000", --  264 - 0x108  :    0 - 0x0 -- Sprite 0x21
    "00000000", --  265 - 0x109  :    0 - 0x0
    "11110000", --  266 - 0x10a  :  240 - 0xf0
    "00001000", --  267 - 0x10b  :    8 - 0x8
    "00001000", --  268 - 0x10c  :    8 - 0x8
    "11110000", --  269 - 0x10d  :  240 - 0xf0
    "00000000", --  270 - 0x10e  :    0 - 0x0
    "00000000", --  271 - 0x10f  :    0 - 0x0
    "00000000", --  272 - 0x110  :    0 - 0x0 -- Sprite 0x22
    "00000000", --  273 - 0x111  :    0 - 0x0
    "00001111", --  274 - 0x112  :   15 - 0xf
    "00010000", --  275 - 0x113  :   16 - 0x10
    "00010000", --  276 - 0x114  :   16 - 0x10
    "00001111", --  277 - 0x115  :   15 - 0xf
    "00000000", --  278 - 0x116  :    0 - 0x0
    "00000000", --  279 - 0x117  :    0 - 0x0
    "11111111", --  280 - 0x118  :  255 - 0xff -- Sprite 0x23
    "11111111", --  281 - 0x119  :  255 - 0xff
    "11100001", --  282 - 0x11a  :  225 - 0xe1
    "11100001", --  283 - 0x11b  :  225 - 0xe1
    "11100001", --  284 - 0x11c  :  225 - 0xe1
    "11100001", --  285 - 0x11d  :  225 - 0xe1
    "11100001", --  286 - 0x11e  :  225 - 0xe1
    "11100001", --  287 - 0x11f  :  225 - 0xe1
    "10000111", --  288 - 0x120  :  135 - 0x87 -- Sprite 0x24
    "11000111", --  289 - 0x121  :  199 - 0xc7
    "11000000", --  290 - 0x122  :  192 - 0xc0
    "11000111", --  291 - 0x123  :  199 - 0xc7
    "11001111", --  292 - 0x124  :  207 - 0xcf
    "11001110", --  293 - 0x125  :  206 - 0xce
    "11001111", --  294 - 0x126  :  207 - 0xcf
    "11000111", --  295 - 0x127  :  199 - 0xc7
    "11111000", --  296 - 0x128  :  248 - 0xf8 -- Sprite 0x25
    "11111100", --  297 - 0x129  :  252 - 0xfc
    "00011100", --  298 - 0x12a  :   28 - 0x1c
    "11111100", --  299 - 0x12b  :  252 - 0xfc
    "11111100", --  300 - 0x12c  :  252 - 0xfc
    "00011100", --  301 - 0x12d  :   28 - 0x1c
    "11111100", --  302 - 0x12e  :  252 - 0xfc
    "11111100", --  303 - 0x12f  :  252 - 0xfc
    "11111111", --  304 - 0x130  :  255 - 0xff -- Sprite 0x26
    "11111111", --  305 - 0x131  :  255 - 0xff
    "11100111", --  306 - 0x132  :  231 - 0xe7
    "11100111", --  307 - 0x133  :  231 - 0xe7
    "11100111", --  308 - 0x134  :  231 - 0xe7
    "11100111", --  309 - 0x135  :  231 - 0xe7
    "11100111", --  310 - 0x136  :  231 - 0xe7
    "11100111", --  311 - 0x137  :  231 - 0xe7
    "11110000", --  312 - 0x138  :  240 - 0xf0 -- Sprite 0x27
    "11111001", --  313 - 0x139  :  249 - 0xf9
    "00111001", --  314 - 0x13a  :   57 - 0x39
    "00111001", --  315 - 0x13b  :   57 - 0x39
    "00111001", --  316 - 0x13c  :   57 - 0x39
    "00111001", --  317 - 0x13d  :   57 - 0x39
    "00111001", --  318 - 0x13e  :   57 - 0x39
    "00111000", --  319 - 0x13f  :   56 - 0x38
    "11111111", --  320 - 0x140  :  255 - 0xff -- Sprite 0x28
    "11111111", --  321 - 0x141  :  255 - 0xff
    "11000000", --  322 - 0x142  :  192 - 0xc0
    "11000000", --  323 - 0x143  :  192 - 0xc0
    "11000000", --  324 - 0x144  :  192 - 0xc0
    "11000000", --  325 - 0x145  :  192 - 0xc0
    "11111111", --  326 - 0x146  :  255 - 0xff
    "11111111", --  327 - 0x147  :  255 - 0xff
    "00011111", --  328 - 0x148  :   31 - 0x1f -- Sprite 0x29
    "00111111", --  329 - 0x149  :   63 - 0x3f
    "00110000", --  330 - 0x14a  :   48 - 0x30
    "00110000", --  331 - 0x14b  :   48 - 0x30
    "00110000", --  332 - 0x14c  :   48 - 0x30
    "00110000", --  333 - 0x14d  :   48 - 0x30
    "00111111", --  334 - 0x14e  :   63 - 0x3f
    "00011111", --  335 - 0x14f  :   31 - 0x1f
    "11100011", --  336 - 0x150  :  227 - 0xe3 -- Sprite 0x2a
    "11110011", --  337 - 0x151  :  243 - 0xf3
    "01110000", --  338 - 0x152  :  112 - 0x70
    "01110000", --  339 - 0x153  :  112 - 0x70
    "01110000", --  340 - 0x154  :  112 - 0x70
    "01110000", --  341 - 0x155  :  112 - 0x70
    "11110000", --  342 - 0x156  :  240 - 0xf0
    "11100000", --  343 - 0x157  :  224 - 0xe0
    "11111110", --  344 - 0x158  :  254 - 0xfe -- Sprite 0x2b
    "11111110", --  345 - 0x159  :  254 - 0xfe
    "01110000", --  346 - 0x15a  :  112 - 0x70
    "01110000", --  347 - 0x15b  :  112 - 0x70
    "01110000", --  348 - 0x15c  :  112 - 0x70
    "01110000", --  349 - 0x15d  :  112 - 0x70
    "01110000", --  350 - 0x15e  :  112 - 0x70
    "01110000", --  351 - 0x15f  :  112 - 0x70
    "00000000", --  352 - 0x160  :    0 - 0x0 -- Sprite 0x2c
    "00000000", --  353 - 0x161  :    0 - 0x0
    "00000000", --  354 - 0x162  :    0 - 0x0
    "00000000", --  355 - 0x163  :    0 - 0x0
    "11111111", --  356 - 0x164  :  255 - 0xff
    "00000000", --  357 - 0x165  :    0 - 0x0
    "00000000", --  358 - 0x166  :    0 - 0x0
    "00000000", --  359 - 0x167  :    0 - 0x0
    "00000000", --  360 - 0x168  :    0 - 0x0 -- Sprite 0x2d
    "00000000", --  361 - 0x169  :    0 - 0x0
    "00000000", --  362 - 0x16a  :    0 - 0x0
    "00000000", --  363 - 0x16b  :    0 - 0x0
    "00000000", --  364 - 0x16c  :    0 - 0x0
    "00000000", --  365 - 0x16d  :    0 - 0x0
    "00000000", --  366 - 0x16e  :    0 - 0x0
    "00000000", --  367 - 0x16f  :    0 - 0x0
    "00000000", --  368 - 0x170  :    0 - 0x0 -- Sprite 0x2e
    "00000000", --  369 - 0x171  :    0 - 0x0
    "00000000", --  370 - 0x172  :    0 - 0x0
    "00011000", --  371 - 0x173  :   24 - 0x18
    "00011000", --  372 - 0x174  :   24 - 0x18
    "00000000", --  373 - 0x175  :    0 - 0x0
    "00000000", --  374 - 0x176  :    0 - 0x0
    "00000000", --  375 - 0x177  :    0 - 0x0
    "00000000", --  376 - 0x178  :    0 - 0x0 -- Sprite 0x2f
    "00000000", --  377 - 0x179  :    0 - 0x0
    "00000000", --  378 - 0x17a  :    0 - 0x0
    "00000000", --  379 - 0x17b  :    0 - 0x0
    "00000000", --  380 - 0x17c  :    0 - 0x0
    "00000000", --  381 - 0x17d  :    0 - 0x0
    "00000000", --  382 - 0x17e  :    0 - 0x0
    "00000000", --  383 - 0x17f  :    0 - 0x0
    "00011100", --  384 - 0x180  :   28 - 0x1c -- Sprite 0x30
    "00100110", --  385 - 0x181  :   38 - 0x26
    "01100011", --  386 - 0x182  :   99 - 0x63
    "01100011", --  387 - 0x183  :   99 - 0x63
    "01100011", --  388 - 0x184  :   99 - 0x63
    "00110010", --  389 - 0x185  :   50 - 0x32
    "00011100", --  390 - 0x186  :   28 - 0x1c
    "00000000", --  391 - 0x187  :    0 - 0x0
    "00001100", --  392 - 0x188  :   12 - 0xc -- Sprite 0x31
    "00011100", --  393 - 0x189  :   28 - 0x1c
    "00001100", --  394 - 0x18a  :   12 - 0xc
    "00001100", --  395 - 0x18b  :   12 - 0xc
    "00001100", --  396 - 0x18c  :   12 - 0xc
    "00001100", --  397 - 0x18d  :   12 - 0xc
    "00111111", --  398 - 0x18e  :   63 - 0x3f
    "00000000", --  399 - 0x18f  :    0 - 0x0
    "00111110", --  400 - 0x190  :   62 - 0x3e -- Sprite 0x32
    "01100011", --  401 - 0x191  :   99 - 0x63
    "00000111", --  402 - 0x192  :    7 - 0x7
    "00011110", --  403 - 0x193  :   30 - 0x1e
    "00111100", --  404 - 0x194  :   60 - 0x3c
    "01110000", --  405 - 0x195  :  112 - 0x70
    "01111111", --  406 - 0x196  :  127 - 0x7f
    "00000000", --  407 - 0x197  :    0 - 0x0
    "00111111", --  408 - 0x198  :   63 - 0x3f -- Sprite 0x33
    "00000110", --  409 - 0x199  :    6 - 0x6
    "00001100", --  410 - 0x19a  :   12 - 0xc
    "00011110", --  411 - 0x19b  :   30 - 0x1e
    "00000011", --  412 - 0x19c  :    3 - 0x3
    "01100011", --  413 - 0x19d  :   99 - 0x63
    "00111110", --  414 - 0x19e  :   62 - 0x3e
    "00000000", --  415 - 0x19f  :    0 - 0x0
    "00001110", --  416 - 0x1a0  :   14 - 0xe -- Sprite 0x34
    "00011110", --  417 - 0x1a1  :   30 - 0x1e
    "00110110", --  418 - 0x1a2  :   54 - 0x36
    "01100110", --  419 - 0x1a3  :  102 - 0x66
    "01111111", --  420 - 0x1a4  :  127 - 0x7f
    "00000110", --  421 - 0x1a5  :    6 - 0x6
    "00000110", --  422 - 0x1a6  :    6 - 0x6
    "00000000", --  423 - 0x1a7  :    0 - 0x0
    "01111110", --  424 - 0x1a8  :  126 - 0x7e -- Sprite 0x35
    "01100000", --  425 - 0x1a9  :   96 - 0x60
    "01111110", --  426 - 0x1aa  :  126 - 0x7e
    "00000011", --  427 - 0x1ab  :    3 - 0x3
    "00000011", --  428 - 0x1ac  :    3 - 0x3
    "01100011", --  429 - 0x1ad  :   99 - 0x63
    "00111110", --  430 - 0x1ae  :   62 - 0x3e
    "00000000", --  431 - 0x1af  :    0 - 0x0
    "00011110", --  432 - 0x1b0  :   30 - 0x1e -- Sprite 0x36
    "00110000", --  433 - 0x1b1  :   48 - 0x30
    "01100000", --  434 - 0x1b2  :   96 - 0x60
    "01111110", --  435 - 0x1b3  :  126 - 0x7e
    "01100011", --  436 - 0x1b4  :   99 - 0x63
    "01100011", --  437 - 0x1b5  :   99 - 0x63
    "00111110", --  438 - 0x1b6  :   62 - 0x3e
    "00000000", --  439 - 0x1b7  :    0 - 0x0
    "01111111", --  440 - 0x1b8  :  127 - 0x7f -- Sprite 0x37
    "01100011", --  441 - 0x1b9  :   99 - 0x63
    "00000110", --  442 - 0x1ba  :    6 - 0x6
    "00001100", --  443 - 0x1bb  :   12 - 0xc
    "00011000", --  444 - 0x1bc  :   24 - 0x18
    "00011000", --  445 - 0x1bd  :   24 - 0x18
    "00011000", --  446 - 0x1be  :   24 - 0x18
    "00000000", --  447 - 0x1bf  :    0 - 0x0
    "00111100", --  448 - 0x1c0  :   60 - 0x3c -- Sprite 0x38
    "01100010", --  449 - 0x1c1  :   98 - 0x62
    "01110010", --  450 - 0x1c2  :  114 - 0x72
    "00111100", --  451 - 0x1c3  :   60 - 0x3c
    "01001111", --  452 - 0x1c4  :   79 - 0x4f
    "01000011", --  453 - 0x1c5  :   67 - 0x43
    "00111110", --  454 - 0x1c6  :   62 - 0x3e
    "00000000", --  455 - 0x1c7  :    0 - 0x0
    "00111110", --  456 - 0x1c8  :   62 - 0x3e -- Sprite 0x39
    "01100011", --  457 - 0x1c9  :   99 - 0x63
    "01100011", --  458 - 0x1ca  :   99 - 0x63
    "00111111", --  459 - 0x1cb  :   63 - 0x3f
    "00000011", --  460 - 0x1cc  :    3 - 0x3
    "00000110", --  461 - 0x1cd  :    6 - 0x6
    "00111100", --  462 - 0x1ce  :   60 - 0x3c
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "00000000", --  464 - 0x1d0  :    0 - 0x0 -- Sprite 0x3a
    "00000000", --  465 - 0x1d1  :    0 - 0x0
    "00000000", --  466 - 0x1d2  :    0 - 0x0
    "01111110", --  467 - 0x1d3  :  126 - 0x7e
    "00000000", --  468 - 0x1d4  :    0 - 0x0
    "00000000", --  469 - 0x1d5  :    0 - 0x0
    "00000000", --  470 - 0x1d6  :    0 - 0x0
    "00000000", --  471 - 0x1d7  :    0 - 0x0
    "00000000", --  472 - 0x1d8  :    0 - 0x0 -- Sprite 0x3b
    "00000010", --  473 - 0x1d9  :    2 - 0x2
    "00000100", --  474 - 0x1da  :    4 - 0x4
    "00001000", --  475 - 0x1db  :    8 - 0x8
    "00010000", --  476 - 0x1dc  :   16 - 0x10
    "00100000", --  477 - 0x1dd  :   32 - 0x20
    "00000000", --  478 - 0x1de  :    0 - 0x0
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "00000000", --  480 - 0x1e0  :    0 - 0x0 -- Sprite 0x3c
    "00000111", --  481 - 0x1e1  :    7 - 0x7
    "00011111", --  482 - 0x1e2  :   31 - 0x1f
    "00111111", --  483 - 0x1e3  :   63 - 0x3f
    "00111111", --  484 - 0x1e4  :   63 - 0x3f
    "00001111", --  485 - 0x1e5  :   15 - 0xf
    "00000011", --  486 - 0x1e6  :    3 - 0x3
    "00000000", --  487 - 0x1e7  :    0 - 0x0
    "00000000", --  488 - 0x1e8  :    0 - 0x0 -- Sprite 0x3d
    "11000000", --  489 - 0x1e9  :  192 - 0xc0
    "11110000", --  490 - 0x1ea  :  240 - 0xf0
    "11111000", --  491 - 0x1eb  :  248 - 0xf8
    "11111000", --  492 - 0x1ec  :  248 - 0xf8
    "11111100", --  493 - 0x1ed  :  252 - 0xfc
    "11111100", --  494 - 0x1ee  :  252 - 0xfc
    "11111100", --  495 - 0x1ef  :  252 - 0xfc
    "00000000", --  496 - 0x1f0  :    0 - 0x0 -- Sprite 0x3e
    "00000011", --  497 - 0x1f1  :    3 - 0x3
    "00001111", --  498 - 0x1f2  :   15 - 0xf
    "00111111", --  499 - 0x1f3  :   63 - 0x3f
    "00111111", --  500 - 0x1f4  :   63 - 0x3f
    "00011111", --  501 - 0x1f5  :   31 - 0x1f
    "00000111", --  502 - 0x1f6  :    7 - 0x7
    "00000000", --  503 - 0x1f7  :    0 - 0x0
    "11111100", --  504 - 0x1f8  :  252 - 0xfc -- Sprite 0x3f
    "11111100", --  505 - 0x1f9  :  252 - 0xfc
    "11111100", --  506 - 0x1fa  :  252 - 0xfc
    "11111000", --  507 - 0x1fb  :  248 - 0xf8
    "11111000", --  508 - 0x1fc  :  248 - 0xf8
    "11110000", --  509 - 0x1fd  :  240 - 0xf0
    "11000000", --  510 - 0x1fe  :  192 - 0xc0
    "00000000", --  511 - 0x1ff  :    0 - 0x0
    "00000000", --  512 - 0x200  :    0 - 0x0 -- Sprite 0x40
    "00000000", --  513 - 0x201  :    0 - 0x0
    "00000000", --  514 - 0x202  :    0 - 0x0
    "00000000", --  515 - 0x203  :    0 - 0x0
    "00000000", --  516 - 0x204  :    0 - 0x0
    "00000000", --  517 - 0x205  :    0 - 0x0
    "00000000", --  518 - 0x206  :    0 - 0x0
    "00000000", --  519 - 0x207  :    0 - 0x0
    "00011100", --  520 - 0x208  :   28 - 0x1c -- Sprite 0x41
    "00110110", --  521 - 0x209  :   54 - 0x36
    "01100011", --  522 - 0x20a  :   99 - 0x63
    "01100011", --  523 - 0x20b  :   99 - 0x63
    "01111111", --  524 - 0x20c  :  127 - 0x7f
    "01100011", --  525 - 0x20d  :   99 - 0x63
    "01100011", --  526 - 0x20e  :   99 - 0x63
    "00000000", --  527 - 0x20f  :    0 - 0x0
    "01111110", --  528 - 0x210  :  126 - 0x7e -- Sprite 0x42
    "01100011", --  529 - 0x211  :   99 - 0x63
    "01100011", --  530 - 0x212  :   99 - 0x63
    "01111110", --  531 - 0x213  :  126 - 0x7e
    "01100011", --  532 - 0x214  :   99 - 0x63
    "01100011", --  533 - 0x215  :   99 - 0x63
    "01111110", --  534 - 0x216  :  126 - 0x7e
    "00000000", --  535 - 0x217  :    0 - 0x0
    "00011110", --  536 - 0x218  :   30 - 0x1e -- Sprite 0x43
    "00110011", --  537 - 0x219  :   51 - 0x33
    "01100000", --  538 - 0x21a  :   96 - 0x60
    "01100000", --  539 - 0x21b  :   96 - 0x60
    "01100000", --  540 - 0x21c  :   96 - 0x60
    "00110011", --  541 - 0x21d  :   51 - 0x33
    "00011110", --  542 - 0x21e  :   30 - 0x1e
    "00000000", --  543 - 0x21f  :    0 - 0x0
    "01111100", --  544 - 0x220  :  124 - 0x7c -- Sprite 0x44
    "01100110", --  545 - 0x221  :  102 - 0x66
    "01100011", --  546 - 0x222  :   99 - 0x63
    "01100011", --  547 - 0x223  :   99 - 0x63
    "01100011", --  548 - 0x224  :   99 - 0x63
    "01100110", --  549 - 0x225  :  102 - 0x66
    "01111100", --  550 - 0x226  :  124 - 0x7c
    "00000000", --  551 - 0x227  :    0 - 0x0
    "01111111", --  552 - 0x228  :  127 - 0x7f -- Sprite 0x45
    "01100000", --  553 - 0x229  :   96 - 0x60
    "01100000", --  554 - 0x22a  :   96 - 0x60
    "01111110", --  555 - 0x22b  :  126 - 0x7e
    "01100000", --  556 - 0x22c  :   96 - 0x60
    "01100000", --  557 - 0x22d  :   96 - 0x60
    "01111111", --  558 - 0x22e  :  127 - 0x7f
    "00000000", --  559 - 0x22f  :    0 - 0x0
    "01111111", --  560 - 0x230  :  127 - 0x7f -- Sprite 0x46
    "01100000", --  561 - 0x231  :   96 - 0x60
    "01100000", --  562 - 0x232  :   96 - 0x60
    "01111110", --  563 - 0x233  :  126 - 0x7e
    "01100000", --  564 - 0x234  :   96 - 0x60
    "01100000", --  565 - 0x235  :   96 - 0x60
    "01100000", --  566 - 0x236  :   96 - 0x60
    "00000000", --  567 - 0x237  :    0 - 0x0
    "00011111", --  568 - 0x238  :   31 - 0x1f -- Sprite 0x47
    "00110000", --  569 - 0x239  :   48 - 0x30
    "01100000", --  570 - 0x23a  :   96 - 0x60
    "01100111", --  571 - 0x23b  :  103 - 0x67
    "01100011", --  572 - 0x23c  :   99 - 0x63
    "00110011", --  573 - 0x23d  :   51 - 0x33
    "00011111", --  574 - 0x23e  :   31 - 0x1f
    "00000000", --  575 - 0x23f  :    0 - 0x0
    "01100011", --  576 - 0x240  :   99 - 0x63 -- Sprite 0x48
    "01100011", --  577 - 0x241  :   99 - 0x63
    "01100011", --  578 - 0x242  :   99 - 0x63
    "01111111", --  579 - 0x243  :  127 - 0x7f
    "01100011", --  580 - 0x244  :   99 - 0x63
    "01100011", --  581 - 0x245  :   99 - 0x63
    "01100011", --  582 - 0x246  :   99 - 0x63
    "00000000", --  583 - 0x247  :    0 - 0x0
    "00111111", --  584 - 0x248  :   63 - 0x3f -- Sprite 0x49
    "00001100", --  585 - 0x249  :   12 - 0xc
    "00001100", --  586 - 0x24a  :   12 - 0xc
    "00001100", --  587 - 0x24b  :   12 - 0xc
    "00001100", --  588 - 0x24c  :   12 - 0xc
    "00001100", --  589 - 0x24d  :   12 - 0xc
    "00111111", --  590 - 0x24e  :   63 - 0x3f
    "00000000", --  591 - 0x24f  :    0 - 0x0
    "00000011", --  592 - 0x250  :    3 - 0x3 -- Sprite 0x4a
    "00000011", --  593 - 0x251  :    3 - 0x3
    "00000011", --  594 - 0x252  :    3 - 0x3
    "00000011", --  595 - 0x253  :    3 - 0x3
    "00000011", --  596 - 0x254  :    3 - 0x3
    "01100011", --  597 - 0x255  :   99 - 0x63
    "00111110", --  598 - 0x256  :   62 - 0x3e
    "00000000", --  599 - 0x257  :    0 - 0x0
    "01100011", --  600 - 0x258  :   99 - 0x63 -- Sprite 0x4b
    "01100110", --  601 - 0x259  :  102 - 0x66
    "01101100", --  602 - 0x25a  :  108 - 0x6c
    "01111000", --  603 - 0x25b  :  120 - 0x78
    "01111100", --  604 - 0x25c  :  124 - 0x7c
    "01100110", --  605 - 0x25d  :  102 - 0x66
    "01100011", --  606 - 0x25e  :   99 - 0x63
    "00000000", --  607 - 0x25f  :    0 - 0x0
    "01100000", --  608 - 0x260  :   96 - 0x60 -- Sprite 0x4c
    "01100000", --  609 - 0x261  :   96 - 0x60
    "01100000", --  610 - 0x262  :   96 - 0x60
    "01100000", --  611 - 0x263  :   96 - 0x60
    "01100000", --  612 - 0x264  :   96 - 0x60
    "01100000", --  613 - 0x265  :   96 - 0x60
    "01111111", --  614 - 0x266  :  127 - 0x7f
    "00000000", --  615 - 0x267  :    0 - 0x0
    "01100011", --  616 - 0x268  :   99 - 0x63 -- Sprite 0x4d
    "01110111", --  617 - 0x269  :  119 - 0x77
    "01111111", --  618 - 0x26a  :  127 - 0x7f
    "01111111", --  619 - 0x26b  :  127 - 0x7f
    "01101011", --  620 - 0x26c  :  107 - 0x6b
    "01100011", --  621 - 0x26d  :   99 - 0x63
    "01100011", --  622 - 0x26e  :   99 - 0x63
    "00000000", --  623 - 0x26f  :    0 - 0x0
    "01100011", --  624 - 0x270  :   99 - 0x63 -- Sprite 0x4e
    "01110011", --  625 - 0x271  :  115 - 0x73
    "01111011", --  626 - 0x272  :  123 - 0x7b
    "01111111", --  627 - 0x273  :  127 - 0x7f
    "01101111", --  628 - 0x274  :  111 - 0x6f
    "01100111", --  629 - 0x275  :  103 - 0x67
    "01100011", --  630 - 0x276  :   99 - 0x63
    "00000000", --  631 - 0x277  :    0 - 0x0
    "00111110", --  632 - 0x278  :   62 - 0x3e -- Sprite 0x4f
    "01100011", --  633 - 0x279  :   99 - 0x63
    "01100011", --  634 - 0x27a  :   99 - 0x63
    "01100011", --  635 - 0x27b  :   99 - 0x63
    "01100011", --  636 - 0x27c  :   99 - 0x63
    "01100011", --  637 - 0x27d  :   99 - 0x63
    "00111110", --  638 - 0x27e  :   62 - 0x3e
    "00000000", --  639 - 0x27f  :    0 - 0x0
    "01111110", --  640 - 0x280  :  126 - 0x7e -- Sprite 0x50
    "01100011", --  641 - 0x281  :   99 - 0x63
    "01100011", --  642 - 0x282  :   99 - 0x63
    "01100011", --  643 - 0x283  :   99 - 0x63
    "01111110", --  644 - 0x284  :  126 - 0x7e
    "01100000", --  645 - 0x285  :   96 - 0x60
    "01100000", --  646 - 0x286  :   96 - 0x60
    "00000000", --  647 - 0x287  :    0 - 0x0
    "00111110", --  648 - 0x288  :   62 - 0x3e -- Sprite 0x51
    "01100011", --  649 - 0x289  :   99 - 0x63
    "01100011", --  650 - 0x28a  :   99 - 0x63
    "01100011", --  651 - 0x28b  :   99 - 0x63
    "01101111", --  652 - 0x28c  :  111 - 0x6f
    "01100110", --  653 - 0x28d  :  102 - 0x66
    "00111101", --  654 - 0x28e  :   61 - 0x3d
    "00000000", --  655 - 0x28f  :    0 - 0x0
    "01111110", --  656 - 0x290  :  126 - 0x7e -- Sprite 0x52
    "01100011", --  657 - 0x291  :   99 - 0x63
    "01100011", --  658 - 0x292  :   99 - 0x63
    "01100111", --  659 - 0x293  :  103 - 0x67
    "01111100", --  660 - 0x294  :  124 - 0x7c
    "01101110", --  661 - 0x295  :  110 - 0x6e
    "01100111", --  662 - 0x296  :  103 - 0x67
    "00000000", --  663 - 0x297  :    0 - 0x0
    "00111100", --  664 - 0x298  :   60 - 0x3c -- Sprite 0x53
    "01100110", --  665 - 0x299  :  102 - 0x66
    "01100000", --  666 - 0x29a  :   96 - 0x60
    "00111110", --  667 - 0x29b  :   62 - 0x3e
    "00000011", --  668 - 0x29c  :    3 - 0x3
    "01100011", --  669 - 0x29d  :   99 - 0x63
    "00111110", --  670 - 0x29e  :   62 - 0x3e
    "00000000", --  671 - 0x29f  :    0 - 0x0
    "00111111", --  672 - 0x2a0  :   63 - 0x3f -- Sprite 0x54
    "00001100", --  673 - 0x2a1  :   12 - 0xc
    "00001100", --  674 - 0x2a2  :   12 - 0xc
    "00001100", --  675 - 0x2a3  :   12 - 0xc
    "00001100", --  676 - 0x2a4  :   12 - 0xc
    "00001100", --  677 - 0x2a5  :   12 - 0xc
    "00001100", --  678 - 0x2a6  :   12 - 0xc
    "00000000", --  679 - 0x2a7  :    0 - 0x0
    "01100011", --  680 - 0x2a8  :   99 - 0x63 -- Sprite 0x55
    "01100011", --  681 - 0x2a9  :   99 - 0x63
    "01100011", --  682 - 0x2aa  :   99 - 0x63
    "01100011", --  683 - 0x2ab  :   99 - 0x63
    "01100011", --  684 - 0x2ac  :   99 - 0x63
    "01100011", --  685 - 0x2ad  :   99 - 0x63
    "00111110", --  686 - 0x2ae  :   62 - 0x3e
    "00000000", --  687 - 0x2af  :    0 - 0x0
    "01100011", --  688 - 0x2b0  :   99 - 0x63 -- Sprite 0x56
    "01100011", --  689 - 0x2b1  :   99 - 0x63
    "01100011", --  690 - 0x2b2  :   99 - 0x63
    "01110111", --  691 - 0x2b3  :  119 - 0x77
    "00111110", --  692 - 0x2b4  :   62 - 0x3e
    "00011100", --  693 - 0x2b5  :   28 - 0x1c
    "00001000", --  694 - 0x2b6  :    8 - 0x8
    "00000000", --  695 - 0x2b7  :    0 - 0x0
    "01100011", --  696 - 0x2b8  :   99 - 0x63 -- Sprite 0x57
    "01100011", --  697 - 0x2b9  :   99 - 0x63
    "01101011", --  698 - 0x2ba  :  107 - 0x6b
    "01111111", --  699 - 0x2bb  :  127 - 0x7f
    "01111111", --  700 - 0x2bc  :  127 - 0x7f
    "01110111", --  701 - 0x2bd  :  119 - 0x77
    "01100011", --  702 - 0x2be  :   99 - 0x63
    "00000000", --  703 - 0x2bf  :    0 - 0x0
    "01100011", --  704 - 0x2c0  :   99 - 0x63 -- Sprite 0x58
    "01110111", --  705 - 0x2c1  :  119 - 0x77
    "00111110", --  706 - 0x2c2  :   62 - 0x3e
    "00011100", --  707 - 0x2c3  :   28 - 0x1c
    "00111110", --  708 - 0x2c4  :   62 - 0x3e
    "01110111", --  709 - 0x2c5  :  119 - 0x77
    "01100011", --  710 - 0x2c6  :   99 - 0x63
    "00000000", --  711 - 0x2c7  :    0 - 0x0
    "00110011", --  712 - 0x2c8  :   51 - 0x33 -- Sprite 0x59
    "00110011", --  713 - 0x2c9  :   51 - 0x33
    "00110011", --  714 - 0x2ca  :   51 - 0x33
    "00011110", --  715 - 0x2cb  :   30 - 0x1e
    "00001100", --  716 - 0x2cc  :   12 - 0xc
    "00001100", --  717 - 0x2cd  :   12 - 0xc
    "00001100", --  718 - 0x2ce  :   12 - 0xc
    "00000000", --  719 - 0x2cf  :    0 - 0x0
    "01111111", --  720 - 0x2d0  :  127 - 0x7f -- Sprite 0x5a
    "00000111", --  721 - 0x2d1  :    7 - 0x7
    "00001110", --  722 - 0x2d2  :   14 - 0xe
    "00011100", --  723 - 0x2d3  :   28 - 0x1c
    "00111000", --  724 - 0x2d4  :   56 - 0x38
    "01110000", --  725 - 0x2d5  :  112 - 0x70
    "01111111", --  726 - 0x2d6  :  127 - 0x7f
    "00000000", --  727 - 0x2d7  :    0 - 0x0
    "00000000", --  728 - 0x2d8  :    0 - 0x0 -- Sprite 0x5b
    "00000000", --  729 - 0x2d9  :    0 - 0x0
    "00000000", --  730 - 0x2da  :    0 - 0x0
    "00000000", --  731 - 0x2db  :    0 - 0x0
    "00000000", --  732 - 0x2dc  :    0 - 0x0
    "00110000", --  733 - 0x2dd  :   48 - 0x30
    "00110000", --  734 - 0x2de  :   48 - 0x30
    "00000000", --  735 - 0x2df  :    0 - 0x0
    "11000000", --  736 - 0x2e0  :  192 - 0xc0 -- Sprite 0x5c
    "11110000", --  737 - 0x2e1  :  240 - 0xf0
    "11111100", --  738 - 0x2e2  :  252 - 0xfc
    "11111111", --  739 - 0x2e3  :  255 - 0xff
    "11111100", --  740 - 0x2e4  :  252 - 0xfc
    "11110000", --  741 - 0x2e5  :  240 - 0xf0
    "11000000", --  742 - 0x2e6  :  192 - 0xc0
    "00000000", --  743 - 0x2e7  :    0 - 0x0
    "00111100", --  744 - 0x2e8  :   60 - 0x3c -- Sprite 0x5d
    "01000010", --  745 - 0x2e9  :   66 - 0x42
    "10011001", --  746 - 0x2ea  :  153 - 0x99
    "10100001", --  747 - 0x2eb  :  161 - 0xa1
    "10100001", --  748 - 0x2ec  :  161 - 0xa1
    "10011001", --  749 - 0x2ed  :  153 - 0x99
    "01000010", --  750 - 0x2ee  :   66 - 0x42
    "00111100", --  751 - 0x2ef  :   60 - 0x3c
    "00000000", --  752 - 0x2f0  :    0 - 0x0 -- Sprite 0x5e
    "00000000", --  753 - 0x2f1  :    0 - 0x0
    "00010000", --  754 - 0x2f2  :   16 - 0x10
    "00010000", --  755 - 0x2f3  :   16 - 0x10
    "00010000", --  756 - 0x2f4  :   16 - 0x10
    "00010000", --  757 - 0x2f5  :   16 - 0x10
    "00000000", --  758 - 0x2f6  :    0 - 0x0
    "00000000", --  759 - 0x2f7  :    0 - 0x0
    "00110110", --  760 - 0x2f8  :   54 - 0x36 -- Sprite 0x5f
    "00110110", --  761 - 0x2f9  :   54 - 0x36
    "00010010", --  762 - 0x2fa  :   18 - 0x12
    "00000000", --  763 - 0x2fb  :    0 - 0x0
    "00000000", --  764 - 0x2fc  :    0 - 0x0
    "00000000", --  765 - 0x2fd  :    0 - 0x0
    "00000000", --  766 - 0x2fe  :    0 - 0x0
    "00000000", --  767 - 0x2ff  :    0 - 0x0
    "00000000", --  768 - 0x300  :    0 - 0x0 -- Sprite 0x60
    "00000000", --  769 - 0x301  :    0 - 0x0
    "00000000", --  770 - 0x302  :    0 - 0x0
    "00000000", --  771 - 0x303  :    0 - 0x0
    "00000000", --  772 - 0x304  :    0 - 0x0
    "00000001", --  773 - 0x305  :    1 - 0x1
    "00011110", --  774 - 0x306  :   30 - 0x1e
    "00111011", --  775 - 0x307  :   59 - 0x3b
    "00000000", --  776 - 0x308  :    0 - 0x0 -- Sprite 0x61
    "00000000", --  777 - 0x309  :    0 - 0x0
    "00001100", --  778 - 0x30a  :   12 - 0xc
    "00111100", --  779 - 0x30b  :   60 - 0x3c
    "11010000", --  780 - 0x30c  :  208 - 0xd0
    "00010000", --  781 - 0x30d  :   16 - 0x10
    "00100000", --  782 - 0x30e  :   32 - 0x20
    "01000000", --  783 - 0x30f  :   64 - 0x40
    "00111110", --  784 - 0x310  :   62 - 0x3e -- Sprite 0x62
    "00101101", --  785 - 0x311  :   45 - 0x2d
    "00110101", --  786 - 0x312  :   53 - 0x35
    "00011101", --  787 - 0x313  :   29 - 0x1d
    "00000001", --  788 - 0x314  :    1 - 0x1
    "00000000", --  789 - 0x315  :    0 - 0x0
    "00000000", --  790 - 0x316  :    0 - 0x0
    "00000000", --  791 - 0x317  :    0 - 0x0
    "10110000", --  792 - 0x318  :  176 - 0xb0 -- Sprite 0x63
    "10111000", --  793 - 0x319  :  184 - 0xb8
    "11111000", --  794 - 0x31a  :  248 - 0xf8
    "01111000", --  795 - 0x31b  :  120 - 0x78
    "10011000", --  796 - 0x31c  :  152 - 0x98
    "11110000", --  797 - 0x31d  :  240 - 0xf0
    "00000000", --  798 - 0x31e  :    0 - 0x0
    "00000000", --  799 - 0x31f  :    0 - 0x0
    "00000000", --  800 - 0x320  :    0 - 0x0 -- Sprite 0x64
    "00000000", --  801 - 0x321  :    0 - 0x0
    "00000111", --  802 - 0x322  :    7 - 0x7
    "00000011", --  803 - 0x323  :    3 - 0x3
    "00001101", --  804 - 0x324  :   13 - 0xd
    "00011110", --  805 - 0x325  :   30 - 0x1e
    "00010111", --  806 - 0x326  :   23 - 0x17
    "00011101", --  807 - 0x327  :   29 - 0x1d
    "00000000", --  808 - 0x328  :    0 - 0x0 -- Sprite 0x65
    "10000000", --  809 - 0x329  :  128 - 0x80
    "01110000", --  810 - 0x32a  :  112 - 0x70
    "11100000", --  811 - 0x32b  :  224 - 0xe0
    "11011000", --  812 - 0x32c  :  216 - 0xd8
    "10111100", --  813 - 0x32d  :  188 - 0xbc
    "01110100", --  814 - 0x32e  :  116 - 0x74
    "11011100", --  815 - 0x32f  :  220 - 0xdc
    "00011111", --  816 - 0x330  :   31 - 0x1f -- Sprite 0x66
    "00001011", --  817 - 0x331  :   11 - 0xb
    "00001111", --  818 - 0x332  :   15 - 0xf
    "00000101", --  819 - 0x333  :    5 - 0x5
    "00000011", --  820 - 0x334  :    3 - 0x3
    "00000001", --  821 - 0x335  :    1 - 0x1
    "00000000", --  822 - 0x336  :    0 - 0x0
    "00000000", --  823 - 0x337  :    0 - 0x0
    "11111100", --  824 - 0x338  :  252 - 0xfc -- Sprite 0x67
    "01101000", --  825 - 0x339  :  104 - 0x68
    "11111000", --  826 - 0x33a  :  248 - 0xf8
    "10110000", --  827 - 0x33b  :  176 - 0xb0
    "11100000", --  828 - 0x33c  :  224 - 0xe0
    "10000000", --  829 - 0x33d  :  128 - 0x80
    "00000000", --  830 - 0x33e  :    0 - 0x0
    "00000000", --  831 - 0x33f  :    0 - 0x0
    "00000000", --  832 - 0x340  :    0 - 0x0 -- Sprite 0x68
    "00000000", --  833 - 0x341  :    0 - 0x0
    "00000000", --  834 - 0x342  :    0 - 0x0
    "00000000", --  835 - 0x343  :    0 - 0x0
    "00000000", --  836 - 0x344  :    0 - 0x0
    "00000000", --  837 - 0x345  :    0 - 0x0
    "00000000", --  838 - 0x346  :    0 - 0x0
    "00000000", --  839 - 0x347  :    0 - 0x0
    "00000000", --  840 - 0x348  :    0 - 0x0 -- Sprite 0x69
    "00000000", --  841 - 0x349  :    0 - 0x0
    "00000000", --  842 - 0x34a  :    0 - 0x0
    "00000000", --  843 - 0x34b  :    0 - 0x0
    "00000000", --  844 - 0x34c  :    0 - 0x0
    "00000000", --  845 - 0x34d  :    0 - 0x0
    "00000000", --  846 - 0x34e  :    0 - 0x0
    "00000000", --  847 - 0x34f  :    0 - 0x0
    "00000000", --  848 - 0x350  :    0 - 0x0 -- Sprite 0x6a
    "00000000", --  849 - 0x351  :    0 - 0x0
    "00000000", --  850 - 0x352  :    0 - 0x0
    "00000000", --  851 - 0x353  :    0 - 0x0
    "00000000", --  852 - 0x354  :    0 - 0x0
    "00000000", --  853 - 0x355  :    0 - 0x0
    "00000000", --  854 - 0x356  :    0 - 0x0
    "00000000", --  855 - 0x357  :    0 - 0x0
    "00000000", --  856 - 0x358  :    0 - 0x0 -- Sprite 0x6b
    "00000000", --  857 - 0x359  :    0 - 0x0
    "00000000", --  858 - 0x35a  :    0 - 0x0
    "00000000", --  859 - 0x35b  :    0 - 0x0
    "00000000", --  860 - 0x35c  :    0 - 0x0
    "00000000", --  861 - 0x35d  :    0 - 0x0
    "00000000", --  862 - 0x35e  :    0 - 0x0
    "00000000", --  863 - 0x35f  :    0 - 0x0
    "00000000", --  864 - 0x360  :    0 - 0x0 -- Sprite 0x6c
    "00000000", --  865 - 0x361  :    0 - 0x0
    "00000001", --  866 - 0x362  :    1 - 0x1
    "00011101", --  867 - 0x363  :   29 - 0x1d
    "00111110", --  868 - 0x364  :   62 - 0x3e
    "00111111", --  869 - 0x365  :   63 - 0x3f
    "00111111", --  870 - 0x366  :   63 - 0x3f
    "00111111", --  871 - 0x367  :   63 - 0x3f
    "00000000", --  872 - 0x368  :    0 - 0x0 -- Sprite 0x6d
    "10000000", --  873 - 0x369  :  128 - 0x80
    "00000000", --  874 - 0x36a  :    0 - 0x0
    "01110000", --  875 - 0x36b  :  112 - 0x70
    "11111000", --  876 - 0x36c  :  248 - 0xf8
    "11111100", --  877 - 0x36d  :  252 - 0xfc
    "11111100", --  878 - 0x36e  :  252 - 0xfc
    "11111100", --  879 - 0x36f  :  252 - 0xfc
    "00111111", --  880 - 0x370  :   63 - 0x3f -- Sprite 0x6e
    "00111111", --  881 - 0x371  :   63 - 0x3f
    "00011111", --  882 - 0x372  :   31 - 0x1f
    "00011111", --  883 - 0x373  :   31 - 0x1f
    "00001111", --  884 - 0x374  :   15 - 0xf
    "00000110", --  885 - 0x375  :    6 - 0x6
    "00000000", --  886 - 0x376  :    0 - 0x0
    "00000000", --  887 - 0x377  :    0 - 0x0
    "11101100", --  888 - 0x378  :  236 - 0xec -- Sprite 0x6f
    "11101100", --  889 - 0x379  :  236 - 0xec
    "11011000", --  890 - 0x37a  :  216 - 0xd8
    "11111000", --  891 - 0x37b  :  248 - 0xf8
    "11110000", --  892 - 0x37c  :  240 - 0xf0
    "11100000", --  893 - 0x37d  :  224 - 0xe0
    "00000000", --  894 - 0x37e  :    0 - 0x0
    "00000000", --  895 - 0x37f  :    0 - 0x0
    "00000000", --  896 - 0x380  :    0 - 0x0 -- Sprite 0x70
    "00000100", --  897 - 0x381  :    4 - 0x4
    "00000011", --  898 - 0x382  :    3 - 0x3
    "00000000", --  899 - 0x383  :    0 - 0x0
    "00000001", --  900 - 0x384  :    1 - 0x1
    "00000111", --  901 - 0x385  :    7 - 0x7
    "00001111", --  902 - 0x386  :   15 - 0xf
    "00001100", --  903 - 0x387  :   12 - 0xc
    "00000000", --  904 - 0x388  :    0 - 0x0 -- Sprite 0x71
    "00000000", --  905 - 0x389  :    0 - 0x0
    "11100000", --  906 - 0x38a  :  224 - 0xe0
    "10000000", --  907 - 0x38b  :  128 - 0x80
    "01000000", --  908 - 0x38c  :   64 - 0x40
    "11110000", --  909 - 0x38d  :  240 - 0xf0
    "10011000", --  910 - 0x38e  :  152 - 0x98
    "11111000", --  911 - 0x38f  :  248 - 0xf8
    "00011111", --  912 - 0x390  :   31 - 0x1f -- Sprite 0x72
    "00010011", --  913 - 0x391  :   19 - 0x13
    "00011111", --  914 - 0x392  :   31 - 0x1f
    "00001111", --  915 - 0x393  :   15 - 0xf
    "00001001", --  916 - 0x394  :    9 - 0x9
    "00000111", --  917 - 0x395  :    7 - 0x7
    "00000001", --  918 - 0x396  :    1 - 0x1
    "00000000", --  919 - 0x397  :    0 - 0x0
    "11100100", --  920 - 0x398  :  228 - 0xe4 -- Sprite 0x73
    "00111100", --  921 - 0x399  :   60 - 0x3c
    "11100100", --  922 - 0x39a  :  228 - 0xe4
    "00111000", --  923 - 0x39b  :   56 - 0x38
    "11111000", --  924 - 0x39c  :  248 - 0xf8
    "11110000", --  925 - 0x39d  :  240 - 0xf0
    "11000000", --  926 - 0x39e  :  192 - 0xc0
    "00000000", --  927 - 0x39f  :    0 - 0x0
    "00000000", --  928 - 0x3a0  :    0 - 0x0 -- Sprite 0x74
    "00000000", --  929 - 0x3a1  :    0 - 0x0
    "00000000", --  930 - 0x3a2  :    0 - 0x0
    "00000000", --  931 - 0x3a3  :    0 - 0x0
    "00000000", --  932 - 0x3a4  :    0 - 0x0
    "00000000", --  933 - 0x3a5  :    0 - 0x0
    "00000000", --  934 - 0x3a6  :    0 - 0x0
    "00000000", --  935 - 0x3a7  :    0 - 0x0
    "00000000", --  936 - 0x3a8  :    0 - 0x0 -- Sprite 0x75
    "00000000", --  937 - 0x3a9  :    0 - 0x0
    "00000000", --  938 - 0x3aa  :    0 - 0x0
    "00000000", --  939 - 0x3ab  :    0 - 0x0
    "00000000", --  940 - 0x3ac  :    0 - 0x0
    "00000000", --  941 - 0x3ad  :    0 - 0x0
    "00000000", --  942 - 0x3ae  :    0 - 0x0
    "00000000", --  943 - 0x3af  :    0 - 0x0
    "00000000", --  944 - 0x3b0  :    0 - 0x0 -- Sprite 0x76
    "00000000", --  945 - 0x3b1  :    0 - 0x0
    "00000000", --  946 - 0x3b2  :    0 - 0x0
    "00000000", --  947 - 0x3b3  :    0 - 0x0
    "00000000", --  948 - 0x3b4  :    0 - 0x0
    "00000000", --  949 - 0x3b5  :    0 - 0x0
    "00000000", --  950 - 0x3b6  :    0 - 0x0
    "00000000", --  951 - 0x3b7  :    0 - 0x0
    "00000000", --  952 - 0x3b8  :    0 - 0x0 -- Sprite 0x77
    "00000000", --  953 - 0x3b9  :    0 - 0x0
    "00000000", --  954 - 0x3ba  :    0 - 0x0
    "00000000", --  955 - 0x3bb  :    0 - 0x0
    "00000000", --  956 - 0x3bc  :    0 - 0x0
    "00000000", --  957 - 0x3bd  :    0 - 0x0
    "00000000", --  958 - 0x3be  :    0 - 0x0
    "00000000", --  959 - 0x3bf  :    0 - 0x0
    "00000000", --  960 - 0x3c0  :    0 - 0x0 -- Sprite 0x78
    "00000000", --  961 - 0x3c1  :    0 - 0x0
    "00000000", --  962 - 0x3c2  :    0 - 0x0
    "00000000", --  963 - 0x3c3  :    0 - 0x0
    "00000000", --  964 - 0x3c4  :    0 - 0x0
    "00000000", --  965 - 0x3c5  :    0 - 0x0
    "00000000", --  966 - 0x3c6  :    0 - 0x0
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "00000000", --  968 - 0x3c8  :    0 - 0x0 -- Sprite 0x79
    "00000000", --  969 - 0x3c9  :    0 - 0x0
    "00000000", --  970 - 0x3ca  :    0 - 0x0
    "00000000", --  971 - 0x3cb  :    0 - 0x0
    "00000000", --  972 - 0x3cc  :    0 - 0x0
    "00000000", --  973 - 0x3cd  :    0 - 0x0
    "00000000", --  974 - 0x3ce  :    0 - 0x0
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "00000000", --  976 - 0x3d0  :    0 - 0x0 -- Sprite 0x7a
    "00000000", --  977 - 0x3d1  :    0 - 0x0
    "00000000", --  978 - 0x3d2  :    0 - 0x0
    "00000000", --  979 - 0x3d3  :    0 - 0x0
    "00000000", --  980 - 0x3d4  :    0 - 0x0
    "00000000", --  981 - 0x3d5  :    0 - 0x0
    "00000000", --  982 - 0x3d6  :    0 - 0x0
    "00000000", --  983 - 0x3d7  :    0 - 0x0
    "00000000", --  984 - 0x3d8  :    0 - 0x0 -- Sprite 0x7b
    "00000000", --  985 - 0x3d9  :    0 - 0x0
    "00000000", --  986 - 0x3da  :    0 - 0x0
    "00000000", --  987 - 0x3db  :    0 - 0x0
    "00000000", --  988 - 0x3dc  :    0 - 0x0
    "00000000", --  989 - 0x3dd  :    0 - 0x0
    "00000000", --  990 - 0x3de  :    0 - 0x0
    "00000000", --  991 - 0x3df  :    0 - 0x0
    "00000000", --  992 - 0x3e0  :    0 - 0x0 -- Sprite 0x7c
    "00000001", --  993 - 0x3e1  :    1 - 0x1
    "00000110", --  994 - 0x3e2  :    6 - 0x6
    "00000111", --  995 - 0x3e3  :    7 - 0x7
    "00000111", --  996 - 0x3e4  :    7 - 0x7
    "00000111", --  997 - 0x3e5  :    7 - 0x7
    "00000001", --  998 - 0x3e6  :    1 - 0x1
    "00000011", --  999 - 0x3e7  :    3 - 0x3
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0 -- Sprite 0x7d
    "11000000", -- 1001 - 0x3e9  :  192 - 0xc0
    "00110000", -- 1002 - 0x3ea  :   48 - 0x30
    "11110000", -- 1003 - 0x3eb  :  240 - 0xf0
    "11110000", -- 1004 - 0x3ec  :  240 - 0xf0
    "11110000", -- 1005 - 0x3ed  :  240 - 0xf0
    "01000000", -- 1006 - 0x3ee  :   64 - 0x40
    "01000000", -- 1007 - 0x3ef  :   64 - 0x40
    "00000001", -- 1008 - 0x3f0  :    1 - 0x1 -- Sprite 0x7e
    "00000000", -- 1009 - 0x3f1  :    0 - 0x0
    "00000001", -- 1010 - 0x3f2  :    1 - 0x1
    "00000011", -- 1011 - 0x3f3  :    3 - 0x3
    "00000001", -- 1012 - 0x3f4  :    1 - 0x1
    "00000000", -- 1013 - 0x3f5  :    0 - 0x0
    "00000000", -- 1014 - 0x3f6  :    0 - 0x0
    "00000000", -- 1015 - 0x3f7  :    0 - 0x0
    "01000000", -- 1016 - 0x3f8  :   64 - 0x40 -- Sprite 0x7f
    "01000000", -- 1017 - 0x3f9  :   64 - 0x40
    "01000000", -- 1018 - 0x3fa  :   64 - 0x40
    "01000000", -- 1019 - 0x3fb  :   64 - 0x40
    "01000000", -- 1020 - 0x3fc  :   64 - 0x40
    "10000000", -- 1021 - 0x3fd  :  128 - 0x80
    "00000000", -- 1022 - 0x3fe  :    0 - 0x0
    "00000000", -- 1023 - 0x3ff  :    0 - 0x0
    "11111111", -- 1024 - 0x400  :  255 - 0xff -- Sprite 0x80
    "11111111", -- 1025 - 0x401  :  255 - 0xff
    "11111111", -- 1026 - 0x402  :  255 - 0xff
    "11111111", -- 1027 - 0x403  :  255 - 0xff
    "11000000", -- 1028 - 0x404  :  192 - 0xc0
    "11000000", -- 1029 - 0x405  :  192 - 0xc0
    "11000000", -- 1030 - 0x406  :  192 - 0xc0
    "11000111", -- 1031 - 0x407  :  199 - 0xc7
    "11111111", -- 1032 - 0x408  :  255 - 0xff -- Sprite 0x81
    "11111111", -- 1033 - 0x409  :  255 - 0xff
    "11111111", -- 1034 - 0x40a  :  255 - 0xff
    "11111111", -- 1035 - 0x40b  :  255 - 0xff
    "00000000", -- 1036 - 0x40c  :    0 - 0x0
    "00000000", -- 1037 - 0x40d  :    0 - 0x0
    "00000000", -- 1038 - 0x40e  :    0 - 0x0
    "11111111", -- 1039 - 0x40f  :  255 - 0xff
    "11111111", -- 1040 - 0x410  :  255 - 0xff -- Sprite 0x82
    "11111111", -- 1041 - 0x411  :  255 - 0xff
    "11111111", -- 1042 - 0x412  :  255 - 0xff
    "11111111", -- 1043 - 0x413  :  255 - 0xff
    "01111111", -- 1044 - 0x414  :  127 - 0x7f
    "00111111", -- 1045 - 0x415  :   63 - 0x3f
    "00011111", -- 1046 - 0x416  :   31 - 0x1f
    "11001111", -- 1047 - 0x417  :  207 - 0xcf
    "11111111", -- 1048 - 0x418  :  255 - 0xff -- Sprite 0x83
    "11111111", -- 1049 - 0x419  :  255 - 0xff
    "11111111", -- 1050 - 0x41a  :  255 - 0xff
    "11110111", -- 1051 - 0x41b  :  247 - 0xf7
    "11110111", -- 1052 - 0x41c  :  247 - 0xf7
    "11100010", -- 1053 - 0x41d  :  226 - 0xe2
    "11100000", -- 1054 - 0x41e  :  224 - 0xe0
    "11000110", -- 1055 - 0x41f  :  198 - 0xc6
    "11111111", -- 1056 - 0x420  :  255 - 0xff -- Sprite 0x84
    "11111111", -- 1057 - 0x421  :  255 - 0xff
    "11111111", -- 1058 - 0x422  :  255 - 0xff
    "11111111", -- 1059 - 0x423  :  255 - 0xff
    "10111111", -- 1060 - 0x424  :  191 - 0xbf
    "10111111", -- 1061 - 0x425  :  191 - 0xbf
    "00011111", -- 1062 - 0x426  :   31 - 0x1f
    "00011111", -- 1063 - 0x427  :   31 - 0x1f
    "11111111", -- 1064 - 0x428  :  255 - 0xff -- Sprite 0x85
    "11111111", -- 1065 - 0x429  :  255 - 0xff
    "11111111", -- 1066 - 0x42a  :  255 - 0xff
    "11111111", -- 1067 - 0x42b  :  255 - 0xff
    "11111110", -- 1068 - 0x42c  :  254 - 0xfe
    "11111000", -- 1069 - 0x42d  :  248 - 0xf8
    "11100000", -- 1070 - 0x42e  :  224 - 0xe0
    "11000000", -- 1071 - 0x42f  :  192 - 0xc0
    "11111111", -- 1072 - 0x430  :  255 - 0xff -- Sprite 0x86
    "11111111", -- 1073 - 0x431  :  255 - 0xff
    "11111111", -- 1074 - 0x432  :  255 - 0xff
    "11111111", -- 1075 - 0x433  :  255 - 0xff
    "00000111", -- 1076 - 0x434  :    7 - 0x7
    "00000000", -- 1077 - 0x435  :    0 - 0x0
    "00111111", -- 1078 - 0x436  :   63 - 0x3f
    "11111111", -- 1079 - 0x437  :  255 - 0xff
    "11111111", -- 1080 - 0x438  :  255 - 0xff -- Sprite 0x87
    "11111111", -- 1081 - 0x439  :  255 - 0xff
    "11111111", -- 1082 - 0x43a  :  255 - 0xff
    "11111111", -- 1083 - 0x43b  :  255 - 0xff
    "11111111", -- 1084 - 0x43c  :  255 - 0xff
    "11111111", -- 1085 - 0x43d  :  255 - 0xff
    "00111111", -- 1086 - 0x43e  :   63 - 0x3f
    "11001111", -- 1087 - 0x43f  :  207 - 0xcf
    "11111111", -- 1088 - 0x440  :  255 - 0xff -- Sprite 0x88
    "11111111", -- 1089 - 0x441  :  255 - 0xff
    "11111111", -- 1090 - 0x442  :  255 - 0xff
    "11111111", -- 1091 - 0x443  :  255 - 0xff
    "11111111", -- 1092 - 0x444  :  255 - 0xff
    "11111111", -- 1093 - 0x445  :  255 - 0xff
    "11111111", -- 1094 - 0x446  :  255 - 0xff
    "11111111", -- 1095 - 0x447  :  255 - 0xff
    "11111111", -- 1096 - 0x448  :  255 - 0xff -- Sprite 0x89
    "11111111", -- 1097 - 0x449  :  255 - 0xff
    "11111111", -- 1098 - 0x44a  :  255 - 0xff
    "01110111", -- 1099 - 0x44b  :  119 - 0x77
    "00010011", -- 1100 - 0x44c  :   19 - 0x13
    "00000001", -- 1101 - 0x44d  :    1 - 0x1
    "00010000", -- 1102 - 0x44e  :   16 - 0x10
    "00011000", -- 1103 - 0x44f  :   24 - 0x18
    "11111111", -- 1104 - 0x450  :  255 - 0xff -- Sprite 0x8a
    "11111111", -- 1105 - 0x451  :  255 - 0xff
    "11111111", -- 1106 - 0x452  :  255 - 0xff
    "11111111", -- 1107 - 0x453  :  255 - 0xff
    "11111111", -- 1108 - 0x454  :  255 - 0xff
    "11111111", -- 1109 - 0x455  :  255 - 0xff
    "11111111", -- 1110 - 0x456  :  255 - 0xff
    "01111111", -- 1111 - 0x457  :  127 - 0x7f
    "11111111", -- 1112 - 0x458  :  255 - 0xff -- Sprite 0x8b
    "11111111", -- 1113 - 0x459  :  255 - 0xff
    "11111111", -- 1114 - 0x45a  :  255 - 0xff
    "11110111", -- 1115 - 0x45b  :  247 - 0xf7
    "11100101", -- 1116 - 0x45c  :  229 - 0xe5
    "11000001", -- 1117 - 0x45d  :  193 - 0xc1
    "10000100", -- 1118 - 0x45e  :  132 - 0x84
    "00001100", -- 1119 - 0x45f  :   12 - 0xc
    "11111111", -- 1120 - 0x460  :  255 - 0xff -- Sprite 0x8c
    "11111111", -- 1121 - 0x461  :  255 - 0xff
    "11111111", -- 1122 - 0x462  :  255 - 0xff
    "11111111", -- 1123 - 0x463  :  255 - 0xff
    "11111111", -- 1124 - 0x464  :  255 - 0xff
    "01111111", -- 1125 - 0x465  :  127 - 0x7f
    "01111110", -- 1126 - 0x466  :  126 - 0x7e
    "01111110", -- 1127 - 0x467  :  126 - 0x7e
    "11111111", -- 1128 - 0x468  :  255 - 0xff -- Sprite 0x8d
    "11111111", -- 1129 - 0x469  :  255 - 0xff
    "10111111", -- 1130 - 0x46a  :  191 - 0xbf
    "10110111", -- 1131 - 0x46b  :  183 - 0xb7
    "00010111", -- 1132 - 0x46c  :   23 - 0x17
    "00000011", -- 1133 - 0x46d  :    3 - 0x3
    "00100011", -- 1134 - 0x46e  :   35 - 0x23
    "00100001", -- 1135 - 0x46f  :   33 - 0x21
    "11111111", -- 1136 - 0x470  :  255 - 0xff -- Sprite 0x8e
    "11111111", -- 1137 - 0x471  :  255 - 0xff
    "11111011", -- 1138 - 0x472  :  251 - 0xfb
    "11111001", -- 1139 - 0x473  :  249 - 0xf9
    "11111000", -- 1140 - 0x474  :  248 - 0xf8
    "11111000", -- 1141 - 0x475  :  248 - 0xf8
    "11111000", -- 1142 - 0x476  :  248 - 0xf8
    "11111000", -- 1143 - 0x477  :  248 - 0xf8
    "11111111", -- 1144 - 0x478  :  255 - 0xff -- Sprite 0x8f
    "11111111", -- 1145 - 0x479  :  255 - 0xff
    "01111000", -- 1146 - 0x47a  :  120 - 0x78
    "00111000", -- 1147 - 0x47b  :   56 - 0x38
    "00011000", -- 1148 - 0x47c  :   24 - 0x18
    "00001000", -- 1149 - 0x47d  :    8 - 0x8
    "10000000", -- 1150 - 0x47e  :  128 - 0x80
    "11000000", -- 1151 - 0x47f  :  192 - 0xc0
    "11111111", -- 1152 - 0x480  :  255 - 0xff -- Sprite 0x90
    "11111111", -- 1153 - 0x481  :  255 - 0xff
    "00000001", -- 1154 - 0x482  :    1 - 0x1
    "00000001", -- 1155 - 0x483  :    1 - 0x1
    "00000001", -- 1156 - 0x484  :    1 - 0x1
    "00000000", -- 1157 - 0x485  :    0 - 0x0
    "11111111", -- 1158 - 0x486  :  255 - 0xff
    "11111111", -- 1159 - 0x487  :  255 - 0xff
    "11111111", -- 1160 - 0x488  :  255 - 0xff -- Sprite 0x91
    "11111111", -- 1161 - 0x489  :  255 - 0xff
    "11111111", -- 1162 - 0x48a  :  255 - 0xff
    "11111111", -- 1163 - 0x48b  :  255 - 0xff
    "11111111", -- 1164 - 0x48c  :  255 - 0xff
    "11111111", -- 1165 - 0x48d  :  255 - 0xff
    "01111111", -- 1166 - 0x48e  :  127 - 0x7f
    "00111111", -- 1167 - 0x48f  :   63 - 0x3f
    "11000111", -- 1168 - 0x490  :  199 - 0xc7 -- Sprite 0x92
    "11000111", -- 1169 - 0x491  :  199 - 0xc7
    "11000111", -- 1170 - 0x492  :  199 - 0xc7
    "11000111", -- 1171 - 0x493  :  199 - 0xc7
    "11000111", -- 1172 - 0x494  :  199 - 0xc7
    "11000111", -- 1173 - 0x495  :  199 - 0xc7
    "11000111", -- 1174 - 0x496  :  199 - 0xc7
    "11000111", -- 1175 - 0x497  :  199 - 0xc7
    "11111111", -- 1176 - 0x498  :  255 - 0xff -- Sprite 0x93
    "11111111", -- 1177 - 0x499  :  255 - 0xff
    "11111111", -- 1178 - 0x49a  :  255 - 0xff
    "11111111", -- 1179 - 0x49b  :  255 - 0xff
    "11111001", -- 1180 - 0x49c  :  249 - 0xf9
    "11111001", -- 1181 - 0x49d  :  249 - 0xf9
    "11111111", -- 1182 - 0x49e  :  255 - 0xff
    "11111111", -- 1183 - 0x49f  :  255 - 0xff
    "11110111", -- 1184 - 0x4a0  :  247 - 0xf7 -- Sprite 0x94
    "11111011", -- 1185 - 0x4a1  :  251 - 0xfb
    "11111011", -- 1186 - 0x4a2  :  251 - 0xfb
    "11111101", -- 1187 - 0x4a3  :  253 - 0xfd
    "11111100", -- 1188 - 0x4a4  :  252 - 0xfc
    "11111100", -- 1189 - 0x4a5  :  252 - 0xfc
    "01111100", -- 1190 - 0x4a6  :  124 - 0x7c
    "01111100", -- 1191 - 0x4a7  :  124 - 0x7c
    "11000111", -- 1192 - 0x4a8  :  199 - 0xc7 -- Sprite 0x95
    "10001111", -- 1193 - 0x4a9  :  143 - 0x8f
    "10001111", -- 1194 - 0x4aa  :  143 - 0x8f
    "00011111", -- 1195 - 0x4ab  :   31 - 0x1f
    "00011111", -- 1196 - 0x4ac  :   31 - 0x1f
    "00111111", -- 1197 - 0x4ad  :   63 - 0x3f
    "00111111", -- 1198 - 0x4ae  :   63 - 0x3f
    "01111111", -- 1199 - 0x4af  :  127 - 0x7f
    "00001111", -- 1200 - 0x4b0  :   15 - 0xf -- Sprite 0x96
    "00001111", -- 1201 - 0x4b1  :   15 - 0xf
    "10000111", -- 1202 - 0x4b2  :  135 - 0x87
    "10000111", -- 1203 - 0x4b3  :  135 - 0x87
    "11000010", -- 1204 - 0x4b4  :  194 - 0xc2
    "11000010", -- 1205 - 0x4b5  :  194 - 0xc2
    "11100000", -- 1206 - 0x4b6  :  224 - 0xe0
    "11100000", -- 1207 - 0x4b7  :  224 - 0xe0
    "10000011", -- 1208 - 0x4b8  :  131 - 0x83 -- Sprite 0x97
    "10001111", -- 1209 - 0x4b9  :  143 - 0x8f
    "00001111", -- 1210 - 0x4ba  :   15 - 0xf
    "00011111", -- 1211 - 0x4bb  :   31 - 0x1f
    "00011111", -- 1212 - 0x4bc  :   31 - 0x1f
    "00111111", -- 1213 - 0x4bd  :   63 - 0x3f
    "00111111", -- 1214 - 0x4be  :   63 - 0x3f
    "00111111", -- 1215 - 0x4bf  :   63 - 0x3f
    "11111111", -- 1216 - 0x4c0  :  255 - 0xff -- Sprite 0x98
    "11111111", -- 1217 - 0x4c1  :  255 - 0xff
    "11111111", -- 1218 - 0x4c2  :  255 - 0xff
    "11111110", -- 1219 - 0x4c3  :  254 - 0xfe
    "11111001", -- 1220 - 0x4c4  :  249 - 0xf9
    "11100111", -- 1221 - 0x4c5  :  231 - 0xe7
    "11111100", -- 1222 - 0x4c6  :  252 - 0xfc
    "11110000", -- 1223 - 0x4c7  :  240 - 0xf0
    "11110111", -- 1224 - 0x4c8  :  247 - 0xf7 -- Sprite 0x99
    "11111011", -- 1225 - 0x4c9  :  251 - 0xfb
    "11111011", -- 1226 - 0x4ca  :  251 - 0xfb
    "01110011", -- 1227 - 0x4cb  :  115 - 0x73
    "11000001", -- 1228 - 0x4cc  :  193 - 0xc1
    "00000011", -- 1229 - 0x4cd  :    3 - 0x3
    "00001111", -- 1230 - 0x4ce  :   15 - 0xf
    "00111111", -- 1231 - 0x4cf  :   63 - 0x3f
    "11111111", -- 1232 - 0x4d0  :  255 - 0xff -- Sprite 0x9a
    "11111111", -- 1233 - 0x4d1  :  255 - 0xff
    "11111111", -- 1234 - 0x4d2  :  255 - 0xff
    "10000000", -- 1235 - 0x4d3  :  128 - 0x80
    "10000000", -- 1236 - 0x4d4  :  128 - 0x80
    "10000000", -- 1237 - 0x4d5  :  128 - 0x80
    "10001111", -- 1238 - 0x4d6  :  143 - 0x8f
    "10001111", -- 1239 - 0x4d7  :  143 - 0x8f
    "11111111", -- 1240 - 0x4d8  :  255 - 0xff -- Sprite 0x9b
    "11111111", -- 1241 - 0x4d9  :  255 - 0xff
    "11111111", -- 1242 - 0x4da  :  255 - 0xff
    "00001111", -- 1243 - 0x4db  :   15 - 0xf
    "00001111", -- 1244 - 0x4dc  :   15 - 0xf
    "00000111", -- 1245 - 0x4dd  :    7 - 0x7
    "11110111", -- 1246 - 0x4de  :  247 - 0xf7
    "11110001", -- 1247 - 0x4df  :  241 - 0xf1
    "00011100", -- 1248 - 0x4e0  :   28 - 0x1c -- Sprite 0x9c
    "00011110", -- 1249 - 0x4e1  :   30 - 0x1e
    "00011111", -- 1250 - 0x4e2  :   31 - 0x1f
    "00011111", -- 1251 - 0x4e3  :   31 - 0x1f
    "00011111", -- 1252 - 0x4e4  :   31 - 0x1f
    "00011111", -- 1253 - 0x4e5  :   31 - 0x1f
    "00011111", -- 1254 - 0x4e6  :   31 - 0x1f
    "00011111", -- 1255 - 0x4e7  :   31 - 0x1f
    "00111110", -- 1256 - 0x4e8  :   62 - 0x3e -- Sprite 0x9d
    "00011100", -- 1257 - 0x4e9  :   28 - 0x1c
    "00001000", -- 1258 - 0x4ea  :    8 - 0x8
    "10000000", -- 1259 - 0x4eb  :  128 - 0x80
    "11000001", -- 1260 - 0x4ec  :  193 - 0xc1
    "11100011", -- 1261 - 0x4ed  :  227 - 0xe3
    "11110111", -- 1262 - 0x4ee  :  247 - 0xf7
    "11111111", -- 1263 - 0x4ef  :  255 - 0xff
    "00011100", -- 1264 - 0x4f0  :   28 - 0x1c -- Sprite 0x9e
    "00111100", -- 1265 - 0x4f1  :   60 - 0x3c
    "01111100", -- 1266 - 0x4f2  :  124 - 0x7c
    "11111100", -- 1267 - 0x4f3  :  252 - 0xfc
    "11111100", -- 1268 - 0x4f4  :  252 - 0xfc
    "11111100", -- 1269 - 0x4f5  :  252 - 0xfc
    "11111100", -- 1270 - 0x4f6  :  252 - 0xfc
    "11111100", -- 1271 - 0x4f7  :  252 - 0xfc
    "01111100", -- 1272 - 0x4f8  :  124 - 0x7c -- Sprite 0x9f
    "01111100", -- 1273 - 0x4f9  :  124 - 0x7c
    "01111000", -- 1274 - 0x4fa  :  120 - 0x78
    "01111000", -- 1275 - 0x4fb  :  120 - 0x78
    "01110001", -- 1276 - 0x4fc  :  113 - 0x71
    "01110001", -- 1277 - 0x4fd  :  113 - 0x71
    "01100011", -- 1278 - 0x4fe  :   99 - 0x63
    "01100011", -- 1279 - 0x4ff  :   99 - 0x63
    "01110001", -- 1280 - 0x500  :  113 - 0x71 -- Sprite 0xa0
    "01110000", -- 1281 - 0x501  :  112 - 0x70
    "11111000", -- 1282 - 0x502  :  248 - 0xf8
    "11111000", -- 1283 - 0x503  :  248 - 0xf8
    "11111100", -- 1284 - 0x504  :  252 - 0xfc
    "11111100", -- 1285 - 0x505  :  252 - 0xfc
    "11111110", -- 1286 - 0x506  :  254 - 0xfe
    "11111110", -- 1287 - 0x507  :  254 - 0xfe
    "11111000", -- 1288 - 0x508  :  248 - 0xf8 -- Sprite 0xa1
    "11111000", -- 1289 - 0x509  :  248 - 0xf8
    "11111000", -- 1290 - 0x50a  :  248 - 0xf8
    "01111000", -- 1291 - 0x50b  :  120 - 0x78
    "01111000", -- 1292 - 0x50c  :  120 - 0x78
    "00111000", -- 1293 - 0x50d  :   56 - 0x38
    "00111000", -- 1294 - 0x50e  :   56 - 0x38
    "00011000", -- 1295 - 0x50f  :   24 - 0x18
    "11100000", -- 1296 - 0x510  :  224 - 0xe0 -- Sprite 0xa2
    "11110000", -- 1297 - 0x511  :  240 - 0xf0
    "11111000", -- 1298 - 0x512  :  248 - 0xf8
    "11111000", -- 1299 - 0x513  :  248 - 0xf8
    "11111100", -- 1300 - 0x514  :  252 - 0xfc
    "11111100", -- 1301 - 0x515  :  252 - 0xfc
    "11111110", -- 1302 - 0x516  :  254 - 0xfe
    "11111111", -- 1303 - 0x517  :  255 - 0xff
    "11111111", -- 1304 - 0x518  :  255 - 0xff -- Sprite 0xa3
    "11111111", -- 1305 - 0x519  :  255 - 0xff
    "11111111", -- 1306 - 0x51a  :  255 - 0xff
    "11111111", -- 1307 - 0x51b  :  255 - 0xff
    "11111111", -- 1308 - 0x51c  :  255 - 0xff
    "11111111", -- 1309 - 0x51d  :  255 - 0xff
    "11111111", -- 1310 - 0x51e  :  255 - 0xff
    "11111111", -- 1311 - 0x51f  :  255 - 0xff
    "00011111", -- 1312 - 0x520  :   31 - 0x1f -- Sprite 0xa4
    "00011111", -- 1313 - 0x521  :   31 - 0x1f
    "00011111", -- 1314 - 0x522  :   31 - 0x1f
    "00011111", -- 1315 - 0x523  :   31 - 0x1f
    "00011111", -- 1316 - 0x524  :   31 - 0x1f
    "00011111", -- 1317 - 0x525  :   31 - 0x1f
    "00011111", -- 1318 - 0x526  :   31 - 0x1f
    "00011111", -- 1319 - 0x527  :   31 - 0x1f
    "11111000", -- 1320 - 0x528  :  248 - 0xf8 -- Sprite 0xa5
    "11111111", -- 1321 - 0x529  :  255 - 0xff
    "11111111", -- 1322 - 0x52a  :  255 - 0xff
    "11111000", -- 1323 - 0x52b  :  248 - 0xf8
    "11111000", -- 1324 - 0x52c  :  248 - 0xf8
    "11111000", -- 1325 - 0x52d  :  248 - 0xf8
    "11111000", -- 1326 - 0x52e  :  248 - 0xf8
    "11111000", -- 1327 - 0x52f  :  248 - 0xf8
    "11111100", -- 1328 - 0x530  :  252 - 0xfc -- Sprite 0xa6
    "11111000", -- 1329 - 0x531  :  248 - 0xf8
    "11110000", -- 1330 - 0x532  :  240 - 0xf0
    "00000001", -- 1331 - 0x533  :    1 - 0x1
    "00000001", -- 1332 - 0x534  :    1 - 0x1
    "00000011", -- 1333 - 0x535  :    3 - 0x3
    "11000011", -- 1334 - 0x536  :  195 - 0xc3
    "10000111", -- 1335 - 0x537  :  135 - 0x87
    "01111111", -- 1336 - 0x538  :  127 - 0x7f -- Sprite 0xa7
    "11111001", -- 1337 - 0x539  :  249 - 0xf9
    "11111001", -- 1338 - 0x53a  :  249 - 0xf9
    "11111111", -- 1339 - 0x53b  :  255 - 0xff
    "11111110", -- 1340 - 0x53c  :  254 - 0xfe
    "11111100", -- 1341 - 0x53d  :  252 - 0xfc
    "11111111", -- 1342 - 0x53e  :  255 - 0xff
    "11111111", -- 1343 - 0x53f  :  255 - 0xff
    "11110000", -- 1344 - 0x540  :  240 - 0xf0 -- Sprite 0xa8
    "11110000", -- 1345 - 0x541  :  240 - 0xf0
    "11111000", -- 1346 - 0x542  :  248 - 0xf8
    "01111000", -- 1347 - 0x543  :  120 - 0x78
    "11111100", -- 1348 - 0x544  :  252 - 0xfc
    "11110100", -- 1349 - 0x545  :  244 - 0xf4
    "11110110", -- 1350 - 0x546  :  246 - 0xf6
    "11111010", -- 1351 - 0x547  :  250 - 0xfa
    "00111111", -- 1352 - 0x548  :   63 - 0x3f -- Sprite 0xa9
    "00111111", -- 1353 - 0x549  :   63 - 0x3f
    "00111111", -- 1354 - 0x54a  :   63 - 0x3f
    "00111111", -- 1355 - 0x54b  :   63 - 0x3f
    "00111111", -- 1356 - 0x54c  :   63 - 0x3f
    "00011111", -- 1357 - 0x54d  :   31 - 0x1f
    "00001111", -- 1358 - 0x54e  :   15 - 0xf
    "00000111", -- 1359 - 0x54f  :    7 - 0x7
    "11100000", -- 1360 - 0x550  :  224 - 0xe0 -- Sprite 0xaa
    "11111000", -- 1361 - 0x551  :  248 - 0xf8
    "11111111", -- 1362 - 0x552  :  255 - 0xff
    "11110011", -- 1363 - 0x553  :  243 - 0xf3
    "11111100", -- 1364 - 0x554  :  252 - 0xfc
    "11111111", -- 1365 - 0x555  :  255 - 0xff
    "11111111", -- 1366 - 0x556  :  255 - 0xff
    "11111111", -- 1367 - 0x557  :  255 - 0xff
    "11111111", -- 1368 - 0x558  :  255 - 0xff -- Sprite 0xab
    "11111111", -- 1369 - 0x559  :  255 - 0xff
    "00111111", -- 1370 - 0x55a  :   63 - 0x3f
    "11001111", -- 1371 - 0x55b  :  207 - 0xcf
    "11110011", -- 1372 - 0x55c  :  243 - 0xf3
    "00111101", -- 1373 - 0x55d  :   61 - 0x3d
    "11011000", -- 1374 - 0x55e  :  216 - 0xd8
    "10110000", -- 1375 - 0x55f  :  176 - 0xb0
    "10001111", -- 1376 - 0x560  :  143 - 0x8f -- Sprite 0xac
    "11101111", -- 1377 - 0x561  :  239 - 0xef
    "11100000", -- 1378 - 0x562  :  224 - 0xe0
    "11111000", -- 1379 - 0x563  :  248 - 0xf8
    "11111000", -- 1380 - 0x564  :  248 - 0xf8
    "11111111", -- 1381 - 0x565  :  255 - 0xff
    "11111111", -- 1382 - 0x566  :  255 - 0xff
    "11111111", -- 1383 - 0x567  :  255 - 0xff
    "11110001", -- 1384 - 0x568  :  241 - 0xf1 -- Sprite 0xad
    "11110001", -- 1385 - 0x569  :  241 - 0xf1
    "00000001", -- 1386 - 0x56a  :    1 - 0x1
    "00000001", -- 1387 - 0x56b  :    1 - 0x1
    "00000001", -- 1388 - 0x56c  :    1 - 0x1
    "11111111", -- 1389 - 0x56d  :  255 - 0xff
    "11111111", -- 1390 - 0x56e  :  255 - 0xff
    "11111111", -- 1391 - 0x56f  :  255 - 0xff
    "00011111", -- 1392 - 0x570  :   31 - 0x1f -- Sprite 0xae
    "00011111", -- 1393 - 0x571  :   31 - 0x1f
    "00011111", -- 1394 - 0x572  :   31 - 0x1f
    "00011111", -- 1395 - 0x573  :   31 - 0x1f
    "00011111", -- 1396 - 0x574  :   31 - 0x1f
    "00011111", -- 1397 - 0x575  :   31 - 0x1f
    "00011111", -- 1398 - 0x576  :   31 - 0x1f
    "00011111", -- 1399 - 0x577  :   31 - 0x1f
    "11111100", -- 1400 - 0x578  :  252 - 0xfc -- Sprite 0xaf
    "11111100", -- 1401 - 0x579  :  252 - 0xfc
    "11111100", -- 1402 - 0x57a  :  252 - 0xfc
    "11111100", -- 1403 - 0x57b  :  252 - 0xfc
    "11110100", -- 1404 - 0x57c  :  244 - 0xf4
    "11110100", -- 1405 - 0x57d  :  244 - 0xf4
    "11110100", -- 1406 - 0x57e  :  244 - 0xf4
    "11110100", -- 1407 - 0x57f  :  244 - 0xf4
    "00001100", -- 1408 - 0x580  :   12 - 0xc -- Sprite 0xb0
    "00011100", -- 1409 - 0x581  :   28 - 0x1c
    "00001100", -- 1410 - 0x582  :   12 - 0xc
    "00001100", -- 1411 - 0x583  :   12 - 0xc
    "00001100", -- 1412 - 0x584  :   12 - 0xc
    "00001100", -- 1413 - 0x585  :   12 - 0xc
    "00111111", -- 1414 - 0x586  :   63 - 0x3f
    "00000000", -- 1415 - 0x587  :    0 - 0x0
    "00111110", -- 1416 - 0x588  :   62 - 0x3e -- Sprite 0xb1
    "01100011", -- 1417 - 0x589  :   99 - 0x63
    "00000111", -- 1418 - 0x58a  :    7 - 0x7
    "00011110", -- 1419 - 0x58b  :   30 - 0x1e
    "00111100", -- 1420 - 0x58c  :   60 - 0x3c
    "01110000", -- 1421 - 0x58d  :  112 - 0x70
    "01111111", -- 1422 - 0x58e  :  127 - 0x7f
    "00000000", -- 1423 - 0x58f  :    0 - 0x0
    "01111110", -- 1424 - 0x590  :  126 - 0x7e -- Sprite 0xb2
    "01100011", -- 1425 - 0x591  :   99 - 0x63
    "01100011", -- 1426 - 0x592  :   99 - 0x63
    "01100011", -- 1427 - 0x593  :   99 - 0x63
    "01111110", -- 1428 - 0x594  :  126 - 0x7e
    "01100000", -- 1429 - 0x595  :   96 - 0x60
    "01100000", -- 1430 - 0x596  :   96 - 0x60
    "00000000", -- 1431 - 0x597  :    0 - 0x0
    "01100011", -- 1432 - 0x598  :   99 - 0x63 -- Sprite 0xb3
    "01100011", -- 1433 - 0x599  :   99 - 0x63
    "01100011", -- 1434 - 0x59a  :   99 - 0x63
    "01100011", -- 1435 - 0x59b  :   99 - 0x63
    "01100011", -- 1436 - 0x59c  :   99 - 0x63
    "01100011", -- 1437 - 0x59d  :   99 - 0x63
    "00111110", -- 1438 - 0x59e  :   62 - 0x3e
    "00000000", -- 1439 - 0x59f  :    0 - 0x0
    "01100011", -- 1440 - 0x5a0  :   99 - 0x63 -- Sprite 0xb4
    "01100011", -- 1441 - 0x5a1  :   99 - 0x63
    "01100011", -- 1442 - 0x5a2  :   99 - 0x63
    "01111111", -- 1443 - 0x5a3  :  127 - 0x7f
    "01100011", -- 1444 - 0x5a4  :   99 - 0x63
    "01100011", -- 1445 - 0x5a5  :   99 - 0x63
    "01100011", -- 1446 - 0x5a6  :   99 - 0x63
    "00000000", -- 1447 - 0x5a7  :    0 - 0x0
    "00111111", -- 1448 - 0x5a8  :   63 - 0x3f -- Sprite 0xb5
    "00001100", -- 1449 - 0x5a9  :   12 - 0xc
    "00001100", -- 1450 - 0x5aa  :   12 - 0xc
    "00001100", -- 1451 - 0x5ab  :   12 - 0xc
    "00001100", -- 1452 - 0x5ac  :   12 - 0xc
    "00001100", -- 1453 - 0x5ad  :   12 - 0xc
    "00111111", -- 1454 - 0x5ae  :   63 - 0x3f
    "00000000", -- 1455 - 0x5af  :    0 - 0x0
    "00000000", -- 1456 - 0x5b0  :    0 - 0x0 -- Sprite 0xb6
    "00000000", -- 1457 - 0x5b1  :    0 - 0x0
    "00000000", -- 1458 - 0x5b2  :    0 - 0x0
    "01111110", -- 1459 - 0x5b3  :  126 - 0x7e
    "00000000", -- 1460 - 0x5b4  :    0 - 0x0
    "00000000", -- 1461 - 0x5b5  :    0 - 0x0
    "00000000", -- 1462 - 0x5b6  :    0 - 0x0
    "00000000", -- 1463 - 0x5b7  :    0 - 0x0
    "00111100", -- 1464 - 0x5b8  :   60 - 0x3c -- Sprite 0xb7
    "01100110", -- 1465 - 0x5b9  :  102 - 0x66
    "01100000", -- 1466 - 0x5ba  :   96 - 0x60
    "00111110", -- 1467 - 0x5bb  :   62 - 0x3e
    "00000011", -- 1468 - 0x5bc  :    3 - 0x3
    "01100011", -- 1469 - 0x5bd  :   99 - 0x63
    "00111110", -- 1470 - 0x5be  :   62 - 0x3e
    "00000000", -- 1471 - 0x5bf  :    0 - 0x0
    "00011110", -- 1472 - 0x5c0  :   30 - 0x1e -- Sprite 0xb8
    "00110011", -- 1473 - 0x5c1  :   51 - 0x33
    "01100000", -- 1474 - 0x5c2  :   96 - 0x60
    "01100000", -- 1475 - 0x5c3  :   96 - 0x60
    "01100000", -- 1476 - 0x5c4  :   96 - 0x60
    "00110011", -- 1477 - 0x5c5  :   51 - 0x33
    "00011110", -- 1478 - 0x5c6  :   30 - 0x1e
    "00000000", -- 1479 - 0x5c7  :    0 - 0x0
    "00111110", -- 1480 - 0x5c8  :   62 - 0x3e -- Sprite 0xb9
    "01100011", -- 1481 - 0x5c9  :   99 - 0x63
    "01100011", -- 1482 - 0x5ca  :   99 - 0x63
    "01100011", -- 1483 - 0x5cb  :   99 - 0x63
    "01100011", -- 1484 - 0x5cc  :   99 - 0x63
    "01100011", -- 1485 - 0x5cd  :   99 - 0x63
    "00111110", -- 1486 - 0x5ce  :   62 - 0x3e
    "00000000", -- 1487 - 0x5cf  :    0 - 0x0
    "01111110", -- 1488 - 0x5d0  :  126 - 0x7e -- Sprite 0xba
    "01100011", -- 1489 - 0x5d1  :   99 - 0x63
    "01100011", -- 1490 - 0x5d2  :   99 - 0x63
    "01100111", -- 1491 - 0x5d3  :  103 - 0x67
    "01111100", -- 1492 - 0x5d4  :  124 - 0x7c
    "01101110", -- 1493 - 0x5d5  :  110 - 0x6e
    "01100111", -- 1494 - 0x5d6  :  103 - 0x67
    "00000000", -- 1495 - 0x5d7  :    0 - 0x0
    "01111111", -- 1496 - 0x5d8  :  127 - 0x7f -- Sprite 0xbb
    "01100000", -- 1497 - 0x5d9  :   96 - 0x60
    "01100000", -- 1498 - 0x5da  :   96 - 0x60
    "01111110", -- 1499 - 0x5db  :  126 - 0x7e
    "01100000", -- 1500 - 0x5dc  :   96 - 0x60
    "01100000", -- 1501 - 0x5dd  :   96 - 0x60
    "01111111", -- 1502 - 0x5de  :  127 - 0x7f
    "00000000", -- 1503 - 0x5df  :    0 - 0x0
    "00000000", -- 1504 - 0x5e0  :    0 - 0x0 -- Sprite 0xbc
    "00100010", -- 1505 - 0x5e1  :   34 - 0x22
    "01100101", -- 1506 - 0x5e2  :  101 - 0x65
    "00100101", -- 1507 - 0x5e3  :   37 - 0x25
    "00100101", -- 1508 - 0x5e4  :   37 - 0x25
    "01110010", -- 1509 - 0x5e5  :  114 - 0x72
    "00000000", -- 1510 - 0x5e6  :    0 - 0x0
    "00000000", -- 1511 - 0x5e7  :    0 - 0x0
    "00000000", -- 1512 - 0x5e8  :    0 - 0x0 -- Sprite 0xbd
    "01110010", -- 1513 - 0x5e9  :  114 - 0x72
    "01000101", -- 1514 - 0x5ea  :   69 - 0x45
    "01100101", -- 1515 - 0x5eb  :  101 - 0x65
    "00010101", -- 1516 - 0x5ec  :   21 - 0x15
    "01100010", -- 1517 - 0x5ed  :   98 - 0x62
    "00000000", -- 1518 - 0x5ee  :    0 - 0x0
    "00000000", -- 1519 - 0x5ef  :    0 - 0x0
    "00000000", -- 1520 - 0x5f0  :    0 - 0x0 -- Sprite 0xbe
    "01100111", -- 1521 - 0x5f1  :  103 - 0x67
    "01010010", -- 1522 - 0x5f2  :   82 - 0x52
    "01100010", -- 1523 - 0x5f3  :   98 - 0x62
    "01000010", -- 1524 - 0x5f4  :   66 - 0x42
    "01000010", -- 1525 - 0x5f5  :   66 - 0x42
    "00000000", -- 1526 - 0x5f6  :    0 - 0x0
    "00000000", -- 1527 - 0x5f7  :    0 - 0x0
    "00000000", -- 1528 - 0x5f8  :    0 - 0x0 -- Sprite 0xbf
    "01100000", -- 1529 - 0x5f9  :   96 - 0x60
    "10000000", -- 1530 - 0x5fa  :  128 - 0x80
    "01000000", -- 1531 - 0x5fb  :   64 - 0x40
    "00100000", -- 1532 - 0x5fc  :   32 - 0x20
    "11000110", -- 1533 - 0x5fd  :  198 - 0xc6
    "00000000", -- 1534 - 0x5fe  :    0 - 0x0
    "00000000", -- 1535 - 0x5ff  :    0 - 0x0
    "01100011", -- 1536 - 0x600  :   99 - 0x63 -- Sprite 0xc0
    "01100110", -- 1537 - 0x601  :  102 - 0x66
    "01101100", -- 1538 - 0x602  :  108 - 0x6c
    "01111000", -- 1539 - 0x603  :  120 - 0x78
    "01111100", -- 1540 - 0x604  :  124 - 0x7c
    "01100110", -- 1541 - 0x605  :  102 - 0x66
    "01100011", -- 1542 - 0x606  :   99 - 0x63
    "00000000", -- 1543 - 0x607  :    0 - 0x0
    "00111111", -- 1544 - 0x608  :   63 - 0x3f -- Sprite 0xc1
    "00001100", -- 1545 - 0x609  :   12 - 0xc
    "00001100", -- 1546 - 0x60a  :   12 - 0xc
    "00001100", -- 1547 - 0x60b  :   12 - 0xc
    "00001100", -- 1548 - 0x60c  :   12 - 0xc
    "00001100", -- 1549 - 0x60d  :   12 - 0xc
    "00111111", -- 1550 - 0x60e  :   63 - 0x3f
    "00000000", -- 1551 - 0x60f  :    0 - 0x0
    "01100011", -- 1552 - 0x610  :   99 - 0x63 -- Sprite 0xc2
    "01110111", -- 1553 - 0x611  :  119 - 0x77
    "01111111", -- 1554 - 0x612  :  127 - 0x7f
    "01111111", -- 1555 - 0x613  :  127 - 0x7f
    "01101011", -- 1556 - 0x614  :  107 - 0x6b
    "01100011", -- 1557 - 0x615  :   99 - 0x63
    "01100011", -- 1558 - 0x616  :   99 - 0x63
    "00000000", -- 1559 - 0x617  :    0 - 0x0
    "00011100", -- 1560 - 0x618  :   28 - 0x1c -- Sprite 0xc3
    "00110110", -- 1561 - 0x619  :   54 - 0x36
    "01100011", -- 1562 - 0x61a  :   99 - 0x63
    "01100011", -- 1563 - 0x61b  :   99 - 0x63
    "01111111", -- 1564 - 0x61c  :  127 - 0x7f
    "01100011", -- 1565 - 0x61d  :   99 - 0x63
    "01100011", -- 1566 - 0x61e  :   99 - 0x63
    "00000000", -- 1567 - 0x61f  :    0 - 0x0
    "00011111", -- 1568 - 0x620  :   31 - 0x1f -- Sprite 0xc4
    "00110000", -- 1569 - 0x621  :   48 - 0x30
    "01100000", -- 1570 - 0x622  :   96 - 0x60
    "01100111", -- 1571 - 0x623  :  103 - 0x67
    "01100011", -- 1572 - 0x624  :   99 - 0x63
    "00110011", -- 1573 - 0x625  :   51 - 0x33
    "00011111", -- 1574 - 0x626  :   31 - 0x1f
    "00000000", -- 1575 - 0x627  :    0 - 0x0
    "01100011", -- 1576 - 0x628  :   99 - 0x63 -- Sprite 0xc5
    "01100011", -- 1577 - 0x629  :   99 - 0x63
    "01100011", -- 1578 - 0x62a  :   99 - 0x63
    "01100011", -- 1579 - 0x62b  :   99 - 0x63
    "01100011", -- 1580 - 0x62c  :   99 - 0x63
    "01100011", -- 1581 - 0x62d  :   99 - 0x63
    "00111110", -- 1582 - 0x62e  :   62 - 0x3e
    "00000000", -- 1583 - 0x62f  :    0 - 0x0
    "01111110", -- 1584 - 0x630  :  126 - 0x7e -- Sprite 0xc6
    "01100011", -- 1585 - 0x631  :   99 - 0x63
    "01100011", -- 1586 - 0x632  :   99 - 0x63
    "01100111", -- 1587 - 0x633  :  103 - 0x67
    "01111100", -- 1588 - 0x634  :  124 - 0x7c
    "01101110", -- 1589 - 0x635  :  110 - 0x6e
    "01100111", -- 1590 - 0x636  :  103 - 0x67
    "00000000", -- 1591 - 0x637  :    0 - 0x0
    "01111111", -- 1592 - 0x638  :  127 - 0x7f -- Sprite 0xc7
    "01100000", -- 1593 - 0x639  :   96 - 0x60
    "01100000", -- 1594 - 0x63a  :   96 - 0x60
    "01111110", -- 1595 - 0x63b  :  126 - 0x7e
    "01100000", -- 1596 - 0x63c  :   96 - 0x60
    "01100000", -- 1597 - 0x63d  :   96 - 0x60
    "01111111", -- 1598 - 0x63e  :  127 - 0x7f
    "00000000", -- 1599 - 0x63f  :    0 - 0x0
    "00110110", -- 1600 - 0x640  :   54 - 0x36 -- Sprite 0xc8
    "00110110", -- 1601 - 0x641  :   54 - 0x36
    "00010010", -- 1602 - 0x642  :   18 - 0x12
    "00000000", -- 1603 - 0x643  :    0 - 0x0
    "00000000", -- 1604 - 0x644  :    0 - 0x0
    "00000000", -- 1605 - 0x645  :    0 - 0x0
    "00000000", -- 1606 - 0x646  :    0 - 0x0
    "00000000", -- 1607 - 0x647  :    0 - 0x0
    "00111110", -- 1608 - 0x648  :   62 - 0x3e -- Sprite 0xc9
    "01100011", -- 1609 - 0x649  :   99 - 0x63
    "01100011", -- 1610 - 0x64a  :   99 - 0x63
    "01100011", -- 1611 - 0x64b  :   99 - 0x63
    "01100011", -- 1612 - 0x64c  :   99 - 0x63
    "01100011", -- 1613 - 0x64d  :   99 - 0x63
    "00111110", -- 1614 - 0x64e  :   62 - 0x3e
    "00000000", -- 1615 - 0x64f  :    0 - 0x0
    "00111100", -- 1616 - 0x650  :   60 - 0x3c -- Sprite 0xca
    "01100110", -- 1617 - 0x651  :  102 - 0x66
    "01100000", -- 1618 - 0x652  :   96 - 0x60
    "00111110", -- 1619 - 0x653  :   62 - 0x3e
    "00000011", -- 1620 - 0x654  :    3 - 0x3
    "01100011", -- 1621 - 0x655  :   99 - 0x63
    "00111110", -- 1622 - 0x656  :   62 - 0x3e
    "00000000", -- 1623 - 0x657  :    0 - 0x0
    "00000000", -- 1624 - 0x658  :    0 - 0x0 -- Sprite 0xcb
    "00000000", -- 1625 - 0x659  :    0 - 0x0
    "00000000", -- 1626 - 0x65a  :    0 - 0x0
    "00000000", -- 1627 - 0x65b  :    0 - 0x0
    "00000000", -- 1628 - 0x65c  :    0 - 0x0
    "00000000", -- 1629 - 0x65d  :    0 - 0x0
    "00000000", -- 1630 - 0x65e  :    0 - 0x0
    "00000000", -- 1631 - 0x65f  :    0 - 0x0
    "00000000", -- 1632 - 0x660  :    0 - 0x0 -- Sprite 0xcc
    "00000000", -- 1633 - 0x661  :    0 - 0x0
    "00000000", -- 1634 - 0x662  :    0 - 0x0
    "00000000", -- 1635 - 0x663  :    0 - 0x0
    "00000000", -- 1636 - 0x664  :    0 - 0x0
    "00000000", -- 1637 - 0x665  :    0 - 0x0
    "00000000", -- 1638 - 0x666  :    0 - 0x0
    "00000000", -- 1639 - 0x667  :    0 - 0x0
    "00000000", -- 1640 - 0x668  :    0 - 0x0 -- Sprite 0xcd
    "00000000", -- 1641 - 0x669  :    0 - 0x0
    "00000000", -- 1642 - 0x66a  :    0 - 0x0
    "00000000", -- 1643 - 0x66b  :    0 - 0x0
    "00000000", -- 1644 - 0x66c  :    0 - 0x0
    "00000000", -- 1645 - 0x66d  :    0 - 0x0
    "00000000", -- 1646 - 0x66e  :    0 - 0x0
    "00000000", -- 1647 - 0x66f  :    0 - 0x0
    "00000000", -- 1648 - 0x670  :    0 - 0x0 -- Sprite 0xce
    "00000000", -- 1649 - 0x671  :    0 - 0x0
    "00000000", -- 1650 - 0x672  :    0 - 0x0
    "00000000", -- 1651 - 0x673  :    0 - 0x0
    "00000000", -- 1652 - 0x674  :    0 - 0x0
    "00000000", -- 1653 - 0x675  :    0 - 0x0
    "00000000", -- 1654 - 0x676  :    0 - 0x0
    "00000000", -- 1655 - 0x677  :    0 - 0x0
    "00000000", -- 1656 - 0x678  :    0 - 0x0 -- Sprite 0xcf
    "00000000", -- 1657 - 0x679  :    0 - 0x0
    "00000000", -- 1658 - 0x67a  :    0 - 0x0
    "00000000", -- 1659 - 0x67b  :    0 - 0x0
    "00000000", -- 1660 - 0x67c  :    0 - 0x0
    "00000000", -- 1661 - 0x67d  :    0 - 0x0
    "00000000", -- 1662 - 0x67e  :    0 - 0x0
    "00000000", -- 1663 - 0x67f  :    0 - 0x0
    "01000111", -- 1664 - 0x680  :   71 - 0x47 -- Sprite 0xd0
    "01000111", -- 1665 - 0x681  :   71 - 0x47
    "00001111", -- 1666 - 0x682  :   15 - 0xf
    "00001111", -- 1667 - 0x683  :   15 - 0xf
    "00011111", -- 1668 - 0x684  :   31 - 0x1f
    "00011111", -- 1669 - 0x685  :   31 - 0x1f
    "00111111", -- 1670 - 0x686  :   63 - 0x3f
    "00111111", -- 1671 - 0x687  :   63 - 0x3f
    "11111111", -- 1672 - 0x688  :  255 - 0xff -- Sprite 0xd1
    "11001111", -- 1673 - 0x689  :  207 - 0xcf
    "11001111", -- 1674 - 0x68a  :  207 - 0xcf
    "11111011", -- 1675 - 0x68b  :  251 - 0xfb
    "11110111", -- 1676 - 0x68c  :  247 - 0xf7
    "11100111", -- 1677 - 0x68d  :  231 - 0xe7
    "11111111", -- 1678 - 0x68e  :  255 - 0xff
    "11111111", -- 1679 - 0x68f  :  255 - 0xff
    "00011000", -- 1680 - 0x690  :   24 - 0x18 -- Sprite 0xd2
    "00001000", -- 1681 - 0x691  :    8 - 0x8
    "10001000", -- 1682 - 0x692  :  136 - 0x88
    "10000000", -- 1683 - 0x693  :  128 - 0x80
    "01000000", -- 1684 - 0x694  :   64 - 0x40
    "01000000", -- 1685 - 0x695  :   64 - 0x40
    "10100000", -- 1686 - 0x696  :  160 - 0xa0
    "10100000", -- 1687 - 0x697  :  160 - 0xa0
    "11111111", -- 1688 - 0x698  :  255 - 0xff -- Sprite 0xd3
    "11111111", -- 1689 - 0x699  :  255 - 0xff
    "11111111", -- 1690 - 0x69a  :  255 - 0xff
    "11111111", -- 1691 - 0x69b  :  255 - 0xff
    "11111101", -- 1692 - 0x69c  :  253 - 0xfd
    "11111101", -- 1693 - 0x69d  :  253 - 0xfd
    "11111101", -- 1694 - 0x69e  :  253 - 0xfd
    "11111101", -- 1695 - 0x69f  :  253 - 0xfd
    "11000111", -- 1696 - 0x6a0  :  199 - 0xc7 -- Sprite 0xd4
    "11110111", -- 1697 - 0x6a1  :  247 - 0xf7
    "11110000", -- 1698 - 0x6a2  :  240 - 0xf0
    "11111000", -- 1699 - 0x6a3  :  248 - 0xf8
    "11111000", -- 1700 - 0x6a4  :  248 - 0xf8
    "11111111", -- 1701 - 0x6a5  :  255 - 0xff
    "11111111", -- 1702 - 0x6a6  :  255 - 0xff
    "11111111", -- 1703 - 0x6a7  :  255 - 0xff
    "11111000", -- 1704 - 0x6a8  :  248 - 0xf8 -- Sprite 0xd5
    "11111000", -- 1705 - 0x6a9  :  248 - 0xf8
    "00000000", -- 1706 - 0x6aa  :    0 - 0x0
    "00000000", -- 1707 - 0x6ab  :    0 - 0x0
    "00000000", -- 1708 - 0x6ac  :    0 - 0x0
    "11111111", -- 1709 - 0x6ad  :  255 - 0xff
    "11111111", -- 1710 - 0x6ae  :  255 - 0xff
    "11111111", -- 1711 - 0x6af  :  255 - 0xff
    "10001111", -- 1712 - 0x6b0  :  143 - 0x8f -- Sprite 0xd6
    "11101111", -- 1713 - 0x6b1  :  239 - 0xef
    "11000000", -- 1714 - 0x6b2  :  192 - 0xc0
    "11110000", -- 1715 - 0x6b3  :  240 - 0xf0
    "11100000", -- 1716 - 0x6b4  :  224 - 0xe0
    "11111111", -- 1717 - 0x6b5  :  255 - 0xff
    "11111111", -- 1718 - 0x6b6  :  255 - 0xff
    "11111111", -- 1719 - 0x6b7  :  255 - 0xff
    "11111111", -- 1720 - 0x6b8  :  255 - 0xff -- Sprite 0xd7
    "11111111", -- 1721 - 0x6b9  :  255 - 0xff
    "00000000", -- 1722 - 0x6ba  :    0 - 0x0
    "00000000", -- 1723 - 0x6bb  :    0 - 0x0
    "00000000", -- 1724 - 0x6bc  :    0 - 0x0
    "11111111", -- 1725 - 0x6bd  :  255 - 0xff
    "11111111", -- 1726 - 0x6be  :  255 - 0xff
    "11111111", -- 1727 - 0x6bf  :  255 - 0xff
    "11000011", -- 1728 - 0x6c0  :  195 - 0xc3 -- Sprite 0xd8
    "11111111", -- 1729 - 0x6c1  :  255 - 0xff
    "00000000", -- 1730 - 0x6c2  :    0 - 0x0
    "00000000", -- 1731 - 0x6c3  :    0 - 0x0
    "00000000", -- 1732 - 0x6c4  :    0 - 0x0
    "11111111", -- 1733 - 0x6c5  :  255 - 0xff
    "11111111", -- 1734 - 0x6c6  :  255 - 0xff
    "11111111", -- 1735 - 0x6c7  :  255 - 0xff
    "00000011", -- 1736 - 0x6c8  :    3 - 0x3 -- Sprite 0xd9
    "10000001", -- 1737 - 0x6c9  :  129 - 0x81
    "00000000", -- 1738 - 0x6ca  :    0 - 0x0
    "00000000", -- 1739 - 0x6cb  :    0 - 0x0
    "00000011", -- 1740 - 0x6cc  :    3 - 0x3
    "11111111", -- 1741 - 0x6cd  :  255 - 0xff
    "11111111", -- 1742 - 0x6ce  :  255 - 0xff
    "11111111", -- 1743 - 0x6cf  :  255 - 0xff
    "11111111", -- 1744 - 0x6d0  :  255 - 0xff -- Sprite 0xda
    "11111111", -- 1745 - 0x6d1  :  255 - 0xff
    "01111110", -- 1746 - 0x6d2  :  126 - 0x7e
    "00000000", -- 1747 - 0x6d3  :    0 - 0x0
    "00000000", -- 1748 - 0x6d4  :    0 - 0x0
    "11100000", -- 1749 - 0x6d5  :  224 - 0xe0
    "11111111", -- 1750 - 0x6d6  :  255 - 0xff
    "11111111", -- 1751 - 0x6d7  :  255 - 0xff
    "01100001", -- 1752 - 0x6d8  :   97 - 0x61 -- Sprite 0xdb
    "11000011", -- 1753 - 0x6d9  :  195 - 0xc3
    "00000111", -- 1754 - 0x6da  :    7 - 0x7
    "00001111", -- 1755 - 0x6db  :   15 - 0xf
    "00011111", -- 1756 - 0x6dc  :   31 - 0x1f
    "01111111", -- 1757 - 0x6dd  :  127 - 0x7f
    "11111111", -- 1758 - 0x6de  :  255 - 0xff
    "11111111", -- 1759 - 0x6df  :  255 - 0xff
    "00011111", -- 1760 - 0x6e0  :   31 - 0x1f -- Sprite 0xdc
    "11011111", -- 1761 - 0x6e1  :  223 - 0xdf
    "11000000", -- 1762 - 0x6e2  :  192 - 0xc0
    "11110000", -- 1763 - 0x6e3  :  240 - 0xf0
    "11110000", -- 1764 - 0x6e4  :  240 - 0xf0
    "11111111", -- 1765 - 0x6e5  :  255 - 0xff
    "11111111", -- 1766 - 0x6e6  :  255 - 0xff
    "11111111", -- 1767 - 0x6e7  :  255 - 0xff
    "10000100", -- 1768 - 0x6e8  :  132 - 0x84 -- Sprite 0xdd
    "11111100", -- 1769 - 0x6e9  :  252 - 0xfc
    "00000000", -- 1770 - 0x6ea  :    0 - 0x0
    "00000000", -- 1771 - 0x6eb  :    0 - 0x0
    "00000000", -- 1772 - 0x6ec  :    0 - 0x0
    "11111111", -- 1773 - 0x6ed  :  255 - 0xff
    "11111111", -- 1774 - 0x6ee  :  255 - 0xff
    "11111111", -- 1775 - 0x6ef  :  255 - 0xff
    "01111111", -- 1776 - 0x6f0  :  127 - 0x7f -- Sprite 0xde
    "01111111", -- 1777 - 0x6f1  :  127 - 0x7f
    "00000000", -- 1778 - 0x6f2  :    0 - 0x0
    "00000000", -- 1779 - 0x6f3  :    0 - 0x0
    "00000000", -- 1780 - 0x6f4  :    0 - 0x0
    "11111111", -- 1781 - 0x6f5  :  255 - 0xff
    "11111111", -- 1782 - 0x6f6  :  255 - 0xff
    "11111111", -- 1783 - 0x6f7  :  255 - 0xff
    "11111100", -- 1784 - 0x6f8  :  252 - 0xfc -- Sprite 0xdf
    "11111111", -- 1785 - 0x6f9  :  255 - 0xff
    "00000000", -- 1786 - 0x6fa  :    0 - 0x0
    "00000000", -- 1787 - 0x6fb  :    0 - 0x0
    "00000000", -- 1788 - 0x6fc  :    0 - 0x0
    "11111111", -- 1789 - 0x6fd  :  255 - 0xff
    "11111111", -- 1790 - 0x6fe  :  255 - 0xff
    "11111111", -- 1791 - 0x6ff  :  255 - 0xff
    "00110000", -- 1792 - 0x700  :   48 - 0x30 -- Sprite 0xe0
    "11110000", -- 1793 - 0x701  :  240 - 0xf0
    "00000000", -- 1794 - 0x702  :    0 - 0x0
    "00000000", -- 1795 - 0x703  :    0 - 0x0
    "00000000", -- 1796 - 0x704  :    0 - 0x0
    "11111111", -- 1797 - 0x705  :  255 - 0xff
    "11111111", -- 1798 - 0x706  :  255 - 0xff
    "11111111", -- 1799 - 0x707  :  255 - 0xff
    "11111111", -- 1800 - 0x708  :  255 - 0xff -- Sprite 0xe1
    "11111111", -- 1801 - 0x709  :  255 - 0xff
    "00000000", -- 1802 - 0x70a  :    0 - 0x0
    "00000000", -- 1803 - 0x70b  :    0 - 0x0
    "00000000", -- 1804 - 0x70c  :    0 - 0x0
    "11111111", -- 1805 - 0x70d  :  255 - 0xff
    "11111111", -- 1806 - 0x70e  :  255 - 0xff
    "11111111", -- 1807 - 0x70f  :  255 - 0xff
    "11100001", -- 1808 - 0x710  :  225 - 0xe1 -- Sprite 0xe2
    "11111111", -- 1809 - 0x711  :  255 - 0xff
    "00000000", -- 1810 - 0x712  :    0 - 0x0
    "00000000", -- 1811 - 0x713  :    0 - 0x0
    "00000000", -- 1812 - 0x714  :    0 - 0x0
    "11111111", -- 1813 - 0x715  :  255 - 0xff
    "11111111", -- 1814 - 0x716  :  255 - 0xff
    "11111111", -- 1815 - 0x717  :  255 - 0xff
    "00011111", -- 1816 - 0x718  :   31 - 0x1f -- Sprite 0xe3
    "00011111", -- 1817 - 0x719  :   31 - 0x1f
    "00011111", -- 1818 - 0x71a  :   31 - 0x1f
    "00011111", -- 1819 - 0x71b  :   31 - 0x1f
    "00011111", -- 1820 - 0x71c  :   31 - 0x1f
    "11111111", -- 1821 - 0x71d  :  255 - 0xff
    "11111111", -- 1822 - 0x71e  :  255 - 0xff
    "11111111", -- 1823 - 0x71f  :  255 - 0xff
    "00000000", -- 1824 - 0x720  :    0 - 0x0 -- Sprite 0xe4
    "00011111", -- 1825 - 0x721  :   31 - 0x1f
    "00111111", -- 1826 - 0x722  :   63 - 0x3f
    "01111000", -- 1827 - 0x723  :  120 - 0x78
    "01110111", -- 1828 - 0x724  :  119 - 0x77
    "01101111", -- 1829 - 0x725  :  111 - 0x6f
    "01101111", -- 1830 - 0x726  :  111 - 0x6f
    "01101111", -- 1831 - 0x727  :  111 - 0x6f
    "00000000", -- 1832 - 0x728  :    0 - 0x0 -- Sprite 0xe5
    "11111000", -- 1833 - 0x729  :  248 - 0xf8
    "11111100", -- 1834 - 0x72a  :  252 - 0xfc
    "00011110", -- 1835 - 0x72b  :   30 - 0x1e
    "11101110", -- 1836 - 0x72c  :  238 - 0xee
    "11110110", -- 1837 - 0x72d  :  246 - 0xf6
    "11110110", -- 1838 - 0x72e  :  246 - 0xf6
    "11110110", -- 1839 - 0x72f  :  246 - 0xf6
    "11110110", -- 1840 - 0x730  :  246 - 0xf6 -- Sprite 0xe6
    "11110110", -- 1841 - 0x731  :  246 - 0xf6
    "11110110", -- 1842 - 0x732  :  246 - 0xf6
    "11101110", -- 1843 - 0x733  :  238 - 0xee
    "00011110", -- 1844 - 0x734  :   30 - 0x1e
    "11111100", -- 1845 - 0x735  :  252 - 0xfc
    "11111000", -- 1846 - 0x736  :  248 - 0xf8
    "00000000", -- 1847 - 0x737  :    0 - 0x0
    "01101111", -- 1848 - 0x738  :  111 - 0x6f -- Sprite 0xe7
    "01101111", -- 1849 - 0x739  :  111 - 0x6f
    "01101111", -- 1850 - 0x73a  :  111 - 0x6f
    "01110111", -- 1851 - 0x73b  :  119 - 0x77
    "01111000", -- 1852 - 0x73c  :  120 - 0x78
    "00111111", -- 1853 - 0x73d  :   63 - 0x3f
    "00011111", -- 1854 - 0x73e  :   31 - 0x1f
    "00000000", -- 1855 - 0x73f  :    0 - 0x0
    "00000000", -- 1856 - 0x740  :    0 - 0x0 -- Sprite 0xe8
    "11111111", -- 1857 - 0x741  :  255 - 0xff
    "11111111", -- 1858 - 0x742  :  255 - 0xff
    "00000000", -- 1859 - 0x743  :    0 - 0x0
    "11111111", -- 1860 - 0x744  :  255 - 0xff
    "11111111", -- 1861 - 0x745  :  255 - 0xff
    "11111111", -- 1862 - 0x746  :  255 - 0xff
    "11111111", -- 1863 - 0x747  :  255 - 0xff
    "11110110", -- 1864 - 0x748  :  246 - 0xf6 -- Sprite 0xe9
    "11110110", -- 1865 - 0x749  :  246 - 0xf6
    "11110110", -- 1866 - 0x74a  :  246 - 0xf6
    "11110110", -- 1867 - 0x74b  :  246 - 0xf6
    "11110110", -- 1868 - 0x74c  :  246 - 0xf6
    "11110110", -- 1869 - 0x74d  :  246 - 0xf6
    "11110110", -- 1870 - 0x74e  :  246 - 0xf6
    "11110110", -- 1871 - 0x74f  :  246 - 0xf6
    "11111111", -- 1872 - 0x750  :  255 - 0xff -- Sprite 0xea
    "11111111", -- 1873 - 0x751  :  255 - 0xff
    "11111111", -- 1874 - 0x752  :  255 - 0xff
    "11111111", -- 1875 - 0x753  :  255 - 0xff
    "00000000", -- 1876 - 0x754  :    0 - 0x0
    "11111111", -- 1877 - 0x755  :  255 - 0xff
    "11111111", -- 1878 - 0x756  :  255 - 0xff
    "00000000", -- 1879 - 0x757  :    0 - 0x0
    "01101111", -- 1880 - 0x758  :  111 - 0x6f -- Sprite 0xeb
    "01101111", -- 1881 - 0x759  :  111 - 0x6f
    "01101111", -- 1882 - 0x75a  :  111 - 0x6f
    "01101111", -- 1883 - 0x75b  :  111 - 0x6f
    "01101111", -- 1884 - 0x75c  :  111 - 0x6f
    "01101111", -- 1885 - 0x75d  :  111 - 0x6f
    "01101111", -- 1886 - 0x75e  :  111 - 0x6f
    "01101111", -- 1887 - 0x75f  :  111 - 0x6f
    "00000000", -- 1888 - 0x760  :    0 - 0x0 -- Sprite 0xec
    "00000000", -- 1889 - 0x761  :    0 - 0x0
    "00000000", -- 1890 - 0x762  :    0 - 0x0
    "00000000", -- 1891 - 0x763  :    0 - 0x0
    "00000000", -- 1892 - 0x764  :    0 - 0x0
    "00000000", -- 1893 - 0x765  :    0 - 0x0
    "00000000", -- 1894 - 0x766  :    0 - 0x0
    "00000000", -- 1895 - 0x767  :    0 - 0x0
    "00000000", -- 1896 - 0x768  :    0 - 0x0 -- Sprite 0xed
    "00000000", -- 1897 - 0x769  :    0 - 0x0
    "00000000", -- 1898 - 0x76a  :    0 - 0x0
    "00000000", -- 1899 - 0x76b  :    0 - 0x0
    "00000000", -- 1900 - 0x76c  :    0 - 0x0
    "00000000", -- 1901 - 0x76d  :    0 - 0x0
    "00000000", -- 1902 - 0x76e  :    0 - 0x0
    "00000000", -- 1903 - 0x76f  :    0 - 0x0
    "00000000", -- 1904 - 0x770  :    0 - 0x0 -- Sprite 0xee
    "00000000", -- 1905 - 0x771  :    0 - 0x0
    "00000000", -- 1906 - 0x772  :    0 - 0x0
    "00000000", -- 1907 - 0x773  :    0 - 0x0
    "00000000", -- 1908 - 0x774  :    0 - 0x0
    "00000000", -- 1909 - 0x775  :    0 - 0x0
    "00000000", -- 1910 - 0x776  :    0 - 0x0
    "00000000", -- 1911 - 0x777  :    0 - 0x0
    "00000000", -- 1912 - 0x778  :    0 - 0x0 -- Sprite 0xef
    "00000000", -- 1913 - 0x779  :    0 - 0x0
    "00000000", -- 1914 - 0x77a  :    0 - 0x0
    "00000000", -- 1915 - 0x77b  :    0 - 0x0
    "00000000", -- 1916 - 0x77c  :    0 - 0x0
    "00000000", -- 1917 - 0x77d  :    0 - 0x0
    "00000000", -- 1918 - 0x77e  :    0 - 0x0
    "00000000", -- 1919 - 0x77f  :    0 - 0x0
    "11111111", -- 1920 - 0x780  :  255 - 0xff -- Sprite 0xf0
    "11111111", -- 1921 - 0x781  :  255 - 0xff
    "11111111", -- 1922 - 0x782  :  255 - 0xff
    "11111111", -- 1923 - 0x783  :  255 - 0xff
    "11111111", -- 1924 - 0x784  :  255 - 0xff
    "11111111", -- 1925 - 0x785  :  255 - 0xff
    "11111111", -- 1926 - 0x786  :  255 - 0xff
    "11111111", -- 1927 - 0x787  :  255 - 0xff
    "11111111", -- 1928 - 0x788  :  255 - 0xff -- Sprite 0xf1
    "11111111", -- 1929 - 0x789  :  255 - 0xff
    "11111111", -- 1930 - 0x78a  :  255 - 0xff
    "11111111", -- 1931 - 0x78b  :  255 - 0xff
    "11111111", -- 1932 - 0x78c  :  255 - 0xff
    "11111111", -- 1933 - 0x78d  :  255 - 0xff
    "11111111", -- 1934 - 0x78e  :  255 - 0xff
    "11111111", -- 1935 - 0x78f  :  255 - 0xff
    "11111111", -- 1936 - 0x790  :  255 - 0xff -- Sprite 0xf2
    "11111111", -- 1937 - 0x791  :  255 - 0xff
    "11111111", -- 1938 - 0x792  :  255 - 0xff
    "11111111", -- 1939 - 0x793  :  255 - 0xff
    "11111111", -- 1940 - 0x794  :  255 - 0xff
    "11111111", -- 1941 - 0x795  :  255 - 0xff
    "11111111", -- 1942 - 0x796  :  255 - 0xff
    "11111111", -- 1943 - 0x797  :  255 - 0xff
    "11111111", -- 1944 - 0x798  :  255 - 0xff -- Sprite 0xf3
    "11111111", -- 1945 - 0x799  :  255 - 0xff
    "11111111", -- 1946 - 0x79a  :  255 - 0xff
    "11111111", -- 1947 - 0x79b  :  255 - 0xff
    "11111111", -- 1948 - 0x79c  :  255 - 0xff
    "11111111", -- 1949 - 0x79d  :  255 - 0xff
    "11111111", -- 1950 - 0x79e  :  255 - 0xff
    "11111111", -- 1951 - 0x79f  :  255 - 0xff
    "11111111", -- 1952 - 0x7a0  :  255 - 0xff -- Sprite 0xf4
    "11111111", -- 1953 - 0x7a1  :  255 - 0xff
    "11111111", -- 1954 - 0x7a2  :  255 - 0xff
    "11111111", -- 1955 - 0x7a3  :  255 - 0xff
    "11111111", -- 1956 - 0x7a4  :  255 - 0xff
    "11111111", -- 1957 - 0x7a5  :  255 - 0xff
    "11111111", -- 1958 - 0x7a6  :  255 - 0xff
    "11111111", -- 1959 - 0x7a7  :  255 - 0xff
    "11111111", -- 1960 - 0x7a8  :  255 - 0xff -- Sprite 0xf5
    "11111111", -- 1961 - 0x7a9  :  255 - 0xff
    "11111111", -- 1962 - 0x7aa  :  255 - 0xff
    "11111111", -- 1963 - 0x7ab  :  255 - 0xff
    "11111111", -- 1964 - 0x7ac  :  255 - 0xff
    "11111111", -- 1965 - 0x7ad  :  255 - 0xff
    "11111111", -- 1966 - 0x7ae  :  255 - 0xff
    "11111111", -- 1967 - 0x7af  :  255 - 0xff
    "11111111", -- 1968 - 0x7b0  :  255 - 0xff -- Sprite 0xf6
    "11111111", -- 1969 - 0x7b1  :  255 - 0xff
    "11111111", -- 1970 - 0x7b2  :  255 - 0xff
    "11111111", -- 1971 - 0x7b3  :  255 - 0xff
    "11111111", -- 1972 - 0x7b4  :  255 - 0xff
    "11111111", -- 1973 - 0x7b5  :  255 - 0xff
    "11111111", -- 1974 - 0x7b6  :  255 - 0xff
    "11111111", -- 1975 - 0x7b7  :  255 - 0xff
    "11111111", -- 1976 - 0x7b8  :  255 - 0xff -- Sprite 0xf7
    "11111111", -- 1977 - 0x7b9  :  255 - 0xff
    "11111111", -- 1978 - 0x7ba  :  255 - 0xff
    "11111111", -- 1979 - 0x7bb  :  255 - 0xff
    "11111111", -- 1980 - 0x7bc  :  255 - 0xff
    "11111111", -- 1981 - 0x7bd  :  255 - 0xff
    "11111111", -- 1982 - 0x7be  :  255 - 0xff
    "11111111", -- 1983 - 0x7bf  :  255 - 0xff
    "11111111", -- 1984 - 0x7c0  :  255 - 0xff -- Sprite 0xf8
    "11111111", -- 1985 - 0x7c1  :  255 - 0xff
    "11111111", -- 1986 - 0x7c2  :  255 - 0xff
    "11111111", -- 1987 - 0x7c3  :  255 - 0xff
    "11111111", -- 1988 - 0x7c4  :  255 - 0xff
    "11111111", -- 1989 - 0x7c5  :  255 - 0xff
    "11111111", -- 1990 - 0x7c6  :  255 - 0xff
    "11111111", -- 1991 - 0x7c7  :  255 - 0xff
    "11111111", -- 1992 - 0x7c8  :  255 - 0xff -- Sprite 0xf9
    "11111111", -- 1993 - 0x7c9  :  255 - 0xff
    "11111111", -- 1994 - 0x7ca  :  255 - 0xff
    "11111111", -- 1995 - 0x7cb  :  255 - 0xff
    "11111111", -- 1996 - 0x7cc  :  255 - 0xff
    "11111111", -- 1997 - 0x7cd  :  255 - 0xff
    "11111111", -- 1998 - 0x7ce  :  255 - 0xff
    "11111111", -- 1999 - 0x7cf  :  255 - 0xff
    "11111111", -- 2000 - 0x7d0  :  255 - 0xff -- Sprite 0xfa
    "11111111", -- 2001 - 0x7d1  :  255 - 0xff
    "11111111", -- 2002 - 0x7d2  :  255 - 0xff
    "11111111", -- 2003 - 0x7d3  :  255 - 0xff
    "11111111", -- 2004 - 0x7d4  :  255 - 0xff
    "11111111", -- 2005 - 0x7d5  :  255 - 0xff
    "11111111", -- 2006 - 0x7d6  :  255 - 0xff
    "11111111", -- 2007 - 0x7d7  :  255 - 0xff
    "11111111", -- 2008 - 0x7d8  :  255 - 0xff -- Sprite 0xfb
    "11111111", -- 2009 - 0x7d9  :  255 - 0xff
    "11111111", -- 2010 - 0x7da  :  255 - 0xff
    "11111111", -- 2011 - 0x7db  :  255 - 0xff
    "11111111", -- 2012 - 0x7dc  :  255 - 0xff
    "11111111", -- 2013 - 0x7dd  :  255 - 0xff
    "11111111", -- 2014 - 0x7de  :  255 - 0xff
    "11111111", -- 2015 - 0x7df  :  255 - 0xff
    "11111111", -- 2016 - 0x7e0  :  255 - 0xff -- Sprite 0xfc
    "11111111", -- 2017 - 0x7e1  :  255 - 0xff
    "11111111", -- 2018 - 0x7e2  :  255 - 0xff
    "11111111", -- 2019 - 0x7e3  :  255 - 0xff
    "11111111", -- 2020 - 0x7e4  :  255 - 0xff
    "11111111", -- 2021 - 0x7e5  :  255 - 0xff
    "11111111", -- 2022 - 0x7e6  :  255 - 0xff
    "11111111", -- 2023 - 0x7e7  :  255 - 0xff
    "11111111", -- 2024 - 0x7e8  :  255 - 0xff -- Sprite 0xfd
    "11111111", -- 2025 - 0x7e9  :  255 - 0xff
    "11111111", -- 2026 - 0x7ea  :  255 - 0xff
    "11111111", -- 2027 - 0x7eb  :  255 - 0xff
    "11111111", -- 2028 - 0x7ec  :  255 - 0xff
    "11111111", -- 2029 - 0x7ed  :  255 - 0xff
    "11111111", -- 2030 - 0x7ee  :  255 - 0xff
    "11111111", -- 2031 - 0x7ef  :  255 - 0xff
    "11111111", -- 2032 - 0x7f0  :  255 - 0xff -- Sprite 0xfe
    "11111111", -- 2033 - 0x7f1  :  255 - 0xff
    "11111111", -- 2034 - 0x7f2  :  255 - 0xff
    "11111111", -- 2035 - 0x7f3  :  255 - 0xff
    "11111111", -- 2036 - 0x7f4  :  255 - 0xff
    "11111111", -- 2037 - 0x7f5  :  255 - 0xff
    "11111111", -- 2038 - 0x7f6  :  255 - 0xff
    "11111111", -- 2039 - 0x7f7  :  255 - 0xff
    "11111111", -- 2040 - 0x7f8  :  255 - 0xff -- Sprite 0xff
    "11111111", -- 2041 - 0x7f9  :  255 - 0xff
    "11111111", -- 2042 - 0x7fa  :  255 - 0xff
    "11111111", -- 2043 - 0x7fb  :  255 - 0xff
    "11111111", -- 2044 - 0x7fc  :  255 - 0xff
    "11111111", -- 2045 - 0x7fd  :  255 - 0xff
    "11111111", -- 2046 - 0x7fe  :  255 - 0xff
    "11111111", -- 2047 - 0x7ff  :  255 - 0xff
          -- Background pattern Table
    "00000000", -- 2048 - 0x800  :    0 - 0x0 -- Background 0x0
    "00000011", -- 2049 - 0x801  :    3 - 0x3
    "00001111", -- 2050 - 0x802  :   15 - 0xf
    "00011111", -- 2051 - 0x803  :   31 - 0x1f
    "00111111", -- 2052 - 0x804  :   63 - 0x3f
    "00111111", -- 2053 - 0x805  :   63 - 0x3f
    "01111111", -- 2054 - 0x806  :  127 - 0x7f
    "01111111", -- 2055 - 0x807  :  127 - 0x7f
    "00000000", -- 2056 - 0x808  :    0 - 0x0 -- Background 0x1
    "11000000", -- 2057 - 0x809  :  192 - 0xc0
    "11110000", -- 2058 - 0x80a  :  240 - 0xf0
    "11111000", -- 2059 - 0x80b  :  248 - 0xf8
    "11111000", -- 2060 - 0x80c  :  248 - 0xf8
    "11111100", -- 2061 - 0x80d  :  252 - 0xfc
    "11111100", -- 2062 - 0x80e  :  252 - 0xfc
    "11111100", -- 2063 - 0x80f  :  252 - 0xfc
    "00000000", -- 2064 - 0x810  :    0 - 0x0 -- Background 0x2
    "00000111", -- 2065 - 0x811  :    7 - 0x7
    "00011111", -- 2066 - 0x812  :   31 - 0x1f
    "00111111", -- 2067 - 0x813  :   63 - 0x3f
    "00111111", -- 2068 - 0x814  :   63 - 0x3f
    "00001111", -- 2069 - 0x815  :   15 - 0xf
    "00000011", -- 2070 - 0x816  :    3 - 0x3
    "00000000", -- 2071 - 0x817  :    0 - 0x0
    "00000000", -- 2072 - 0x818  :    0 - 0x0 -- Background 0x3
    "00000000", -- 2073 - 0x819  :    0 - 0x0
    "00000111", -- 2074 - 0x81a  :    7 - 0x7
    "00011111", -- 2075 - 0x81b  :   31 - 0x1f
    "00111111", -- 2076 - 0x81c  :   63 - 0x3f
    "00111111", -- 2077 - 0x81d  :   63 - 0x3f
    "01111111", -- 2078 - 0x81e  :  127 - 0x7f
    "01111111", -- 2079 - 0x81f  :  127 - 0x7f
    "01111110", -- 2080 - 0x820  :  126 - 0x7e -- Background 0x4
    "01111110", -- 2081 - 0x821  :  126 - 0x7e
    "01111100", -- 2082 - 0x822  :  124 - 0x7c
    "00111100", -- 2083 - 0x823  :   60 - 0x3c
    "00111000", -- 2084 - 0x824  :   56 - 0x38
    "00011000", -- 2085 - 0x825  :   24 - 0x18
    "00000000", -- 2086 - 0x826  :    0 - 0x0
    "00000000", -- 2087 - 0x827  :    0 - 0x0
    "00000000", -- 2088 - 0x828  :    0 - 0x0 -- Background 0x5
    "11000000", -- 2089 - 0x829  :  192 - 0xc0
    "11110000", -- 2090 - 0x82a  :  240 - 0xf0
    "11111000", -- 2091 - 0x82b  :  248 - 0xf8
    "11111000", -- 2092 - 0x82c  :  248 - 0xf8
    "11111100", -- 2093 - 0x82d  :  252 - 0xfc
    "01111100", -- 2094 - 0x82e  :  124 - 0x7c
    "00111100", -- 2095 - 0x82f  :   60 - 0x3c
    "00000000", -- 2096 - 0x830  :    0 - 0x0 -- Background 0x6
    "00000111", -- 2097 - 0x831  :    7 - 0x7
    "00000111", -- 2098 - 0x832  :    7 - 0x7
    "00000011", -- 2099 - 0x833  :    3 - 0x3
    "00000001", -- 2100 - 0x834  :    1 - 0x1
    "00000000", -- 2101 - 0x835  :    0 - 0x0
    "00000000", -- 2102 - 0x836  :    0 - 0x0
    "00000000", -- 2103 - 0x837  :    0 - 0x0
    "00000000", -- 2104 - 0x838  :    0 - 0x0 -- Background 0x7
    "00000000", -- 2105 - 0x839  :    0 - 0x0
    "00000111", -- 2106 - 0x83a  :    7 - 0x7
    "00011111", -- 2107 - 0x83b  :   31 - 0x1f
    "00111111", -- 2108 - 0x83c  :   63 - 0x3f
    "00111111", -- 2109 - 0x83d  :   63 - 0x3f
    "01111110", -- 2110 - 0x83e  :  126 - 0x7e
    "01111100", -- 2111 - 0x83f  :  124 - 0x7c
    "01111000", -- 2112 - 0x840  :  120 - 0x78 -- Background 0x8
    "01110000", -- 2113 - 0x841  :  112 - 0x70
    "01100000", -- 2114 - 0x842  :   96 - 0x60
    "00000000", -- 2115 - 0x843  :    0 - 0x0
    "00000000", -- 2116 - 0x844  :    0 - 0x0
    "00000000", -- 2117 - 0x845  :    0 - 0x0
    "00000000", -- 2118 - 0x846  :    0 - 0x0
    "00000000", -- 2119 - 0x847  :    0 - 0x0
    "00000000", -- 2120 - 0x848  :    0 - 0x0 -- Background 0x9
    "00000000", -- 2121 - 0x849  :    0 - 0x0
    "00000000", -- 2122 - 0x84a  :    0 - 0x0
    "00000000", -- 2123 - 0x84b  :    0 - 0x0
    "00000000", -- 2124 - 0x84c  :    0 - 0x0
    "01000000", -- 2125 - 0x84d  :   64 - 0x40
    "11110000", -- 2126 - 0x84e  :  240 - 0xf0
    "11111000", -- 2127 - 0x84f  :  248 - 0xf8
    "11111110", -- 2128 - 0x850  :  254 - 0xfe -- Background 0xa
    "01111111", -- 2129 - 0x851  :  127 - 0x7f
    "01111111", -- 2130 - 0x852  :  127 - 0x7f
    "00111111", -- 2131 - 0x853  :   63 - 0x3f
    "00001110", -- 2132 - 0x854  :   14 - 0xe
    "00000000", -- 2133 - 0x855  :    0 - 0x0
    "00000000", -- 2134 - 0x856  :    0 - 0x0
    "00000000", -- 2135 - 0x857  :    0 - 0x0
    "00000000", -- 2136 - 0x858  :    0 - 0x0 -- Background 0xb
    "00000000", -- 2137 - 0x859  :    0 - 0x0
    "00000000", -- 2138 - 0x85a  :    0 - 0x0
    "00000000", -- 2139 - 0x85b  :    0 - 0x0
    "00000000", -- 2140 - 0x85c  :    0 - 0x0
    "00000000", -- 2141 - 0x85d  :    0 - 0x0
    "00000000", -- 2142 - 0x85e  :    0 - 0x0
    "11100000", -- 2143 - 0x85f  :  224 - 0xe0
    "11111100", -- 2144 - 0x860  :  252 - 0xfc -- Background 0xc
    "11111111", -- 2145 - 0x861  :  255 - 0xff
    "01111111", -- 2146 - 0x862  :  127 - 0x7f
    "00111111", -- 2147 - 0x863  :   63 - 0x3f
    "00001110", -- 2148 - 0x864  :   14 - 0xe
    "00000000", -- 2149 - 0x865  :    0 - 0x0
    "00000000", -- 2150 - 0x866  :    0 - 0x0
    "00000000", -- 2151 - 0x867  :    0 - 0x0
    "11110000", -- 2152 - 0x868  :  240 - 0xf0 -- Background 0xd
    "11111111", -- 2153 - 0x869  :  255 - 0xff
    "11111111", -- 2154 - 0x86a  :  255 - 0xff
    "01111111", -- 2155 - 0x86b  :  127 - 0x7f
    "00011110", -- 2156 - 0x86c  :   30 - 0x1e
    "00000000", -- 2157 - 0x86d  :    0 - 0x0
    "00000000", -- 2158 - 0x86e  :    0 - 0x0
    "00000000", -- 2159 - 0x86f  :    0 - 0x0
    "00000000", -- 2160 - 0x870  :    0 - 0x0 -- Background 0xe
    "00001111", -- 2161 - 0x871  :   15 - 0xf
    "11111111", -- 2162 - 0x872  :  255 - 0xff
    "11111111", -- 2163 - 0x873  :  255 - 0xff
    "01111111", -- 2164 - 0x874  :  127 - 0x7f
    "00011110", -- 2165 - 0x875  :   30 - 0x1e
    "00000000", -- 2166 - 0x876  :    0 - 0x0
    "00000000", -- 2167 - 0x877  :    0 - 0x0
    "00000000", -- 2168 - 0x878  :    0 - 0x0 -- Background 0xf
    "00000011", -- 2169 - 0x879  :    3 - 0x3
    "00001111", -- 2170 - 0x87a  :   15 - 0xf
    "01111111", -- 2171 - 0x87b  :  127 - 0x7f
    "11111111", -- 2172 - 0x87c  :  255 - 0xff
    "01111110", -- 2173 - 0x87d  :  126 - 0x7e
    "00011100", -- 2174 - 0x87e  :   28 - 0x1c
    "00000000", -- 2175 - 0x87f  :    0 - 0x0
    "00000000", -- 2176 - 0x880  :    0 - 0x0 -- Background 0x10
    "00000001", -- 2177 - 0x881  :    1 - 0x1
    "00000011", -- 2178 - 0x882  :    3 - 0x3
    "00001111", -- 2179 - 0x883  :   15 - 0xf
    "00011111", -- 2180 - 0x884  :   31 - 0x1f
    "01111111", -- 2181 - 0x885  :  127 - 0x7f
    "01111110", -- 2182 - 0x886  :  126 - 0x7e
    "00111100", -- 2183 - 0x887  :   60 - 0x3c
    "00000000", -- 2184 - 0x888  :    0 - 0x0 -- Background 0x11
    "00000001", -- 2185 - 0x889  :    1 - 0x1
    "00000011", -- 2186 - 0x88a  :    3 - 0x3
    "00000111", -- 2187 - 0x88b  :    7 - 0x7
    "00000111", -- 2188 - 0x88c  :    7 - 0x7
    "00001111", -- 2189 - 0x88d  :   15 - 0xf
    "00011111", -- 2190 - 0x88e  :   31 - 0x1f
    "00001110", -- 2191 - 0x88f  :   14 - 0xe
    "00000000", -- 2192 - 0x890  :    0 - 0x0 -- Background 0x12
    "00000000", -- 2193 - 0x891  :    0 - 0x0
    "00000001", -- 2194 - 0x892  :    1 - 0x1
    "00000011", -- 2195 - 0x893  :    3 - 0x3
    "00000011", -- 2196 - 0x894  :    3 - 0x3
    "00000011", -- 2197 - 0x895  :    3 - 0x3
    "00000111", -- 2198 - 0x896  :    7 - 0x7
    "00000010", -- 2199 - 0x897  :    2 - 0x2
    "00000000", -- 2200 - 0x898  :    0 - 0x0 -- Background 0x13
    "00000000", -- 2201 - 0x899  :    0 - 0x0
    "00000001", -- 2202 - 0x89a  :    1 - 0x1
    "00000001", -- 2203 - 0x89b  :    1 - 0x1
    "00000001", -- 2204 - 0x89c  :    1 - 0x1
    "00000001", -- 2205 - 0x89d  :    1 - 0x1
    "00000001", -- 2206 - 0x89e  :    1 - 0x1
    "00000001", -- 2207 - 0x89f  :    1 - 0x1
    "00000000", -- 2208 - 0x8a0  :    0 - 0x0 -- Background 0x14
    "00000000", -- 2209 - 0x8a1  :    0 - 0x0
    "00000000", -- 2210 - 0x8a2  :    0 - 0x0
    "00000000", -- 2211 - 0x8a3  :    0 - 0x0
    "00000000", -- 2212 - 0x8a4  :    0 - 0x0
    "00000000", -- 2213 - 0x8a5  :    0 - 0x0
    "00000100", -- 2214 - 0x8a6  :    4 - 0x4
    "00000010", -- 2215 - 0x8a7  :    2 - 0x2
    "00000000", -- 2216 - 0x8a8  :    0 - 0x0 -- Background 0x15
    "00000000", -- 2217 - 0x8a9  :    0 - 0x0
    "00000000", -- 2218 - 0x8aa  :    0 - 0x0
    "00000000", -- 2219 - 0x8ab  :    0 - 0x0
    "00000000", -- 2220 - 0x8ac  :    0 - 0x0
    "00000000", -- 2221 - 0x8ad  :    0 - 0x0
    "00100000", -- 2222 - 0x8ae  :   32 - 0x20
    "01001000", -- 2223 - 0x8af  :   72 - 0x48
    "00010000", -- 2224 - 0x8b0  :   16 - 0x10 -- Background 0x16
    "00001000", -- 2225 - 0x8b1  :    8 - 0x8
    "00000000", -- 2226 - 0x8b2  :    0 - 0x0
    "00110000", -- 2227 - 0x8b3  :   48 - 0x30
    "00000000", -- 2228 - 0x8b4  :    0 - 0x0
    "00001000", -- 2229 - 0x8b5  :    8 - 0x8
    "00010010", -- 2230 - 0x8b6  :   18 - 0x12
    "00000100", -- 2231 - 0x8b7  :    4 - 0x4
    "00010000", -- 2232 - 0x8b8  :   16 - 0x10 -- Background 0x17
    "00000000", -- 2233 - 0x8b9  :    0 - 0x0
    "00001100", -- 2234 - 0x8ba  :   12 - 0xc
    "00000000", -- 2235 - 0x8bb  :    0 - 0x0
    "00010000", -- 2236 - 0x8bc  :   16 - 0x10
    "00001000", -- 2237 - 0x8bd  :    8 - 0x8
    "01000000", -- 2238 - 0x8be  :   64 - 0x40
    "00100000", -- 2239 - 0x8bf  :   32 - 0x20
    "00000000", -- 2240 - 0x8c0  :    0 - 0x0 -- Background 0x18
    "00000000", -- 2241 - 0x8c1  :    0 - 0x0
    "00000011", -- 2242 - 0x8c2  :    3 - 0x3
    "00000011", -- 2243 - 0x8c3  :    3 - 0x3
    "00000001", -- 2244 - 0x8c4  :    1 - 0x1
    "00100001", -- 2245 - 0x8c5  :   33 - 0x21
    "00100001", -- 2246 - 0x8c6  :   33 - 0x21
    "01110011", -- 2247 - 0x8c7  :  115 - 0x73
    "01111111", -- 2248 - 0x8c8  :  127 - 0x7f -- Background 0x19
    "01111111", -- 2249 - 0x8c9  :  127 - 0x7f
    "01111111", -- 2250 - 0x8ca  :  127 - 0x7f
    "01111111", -- 2251 - 0x8cb  :  127 - 0x7f
    "01101110", -- 2252 - 0x8cc  :  110 - 0x6e
    "01000110", -- 2253 - 0x8cd  :   70 - 0x46
    "00000000", -- 2254 - 0x8ce  :    0 - 0x0
    "00000000", -- 2255 - 0x8cf  :    0 - 0x0
    "01111111", -- 2256 - 0x8d0  :  127 - 0x7f -- Background 0x1a
    "01111111", -- 2257 - 0x8d1  :  127 - 0x7f
    "01111111", -- 2258 - 0x8d2  :  127 - 0x7f
    "01111111", -- 2259 - 0x8d3  :  127 - 0x7f
    "01111011", -- 2260 - 0x8d4  :  123 - 0x7b
    "00110001", -- 2261 - 0x8d5  :   49 - 0x31
    "00000000", -- 2262 - 0x8d6  :    0 - 0x0
    "00000000", -- 2263 - 0x8d7  :    0 - 0x0
    "00000000", -- 2264 - 0x8d8  :    0 - 0x0 -- Background 0x1b
    "00000011", -- 2265 - 0x8d9  :    3 - 0x3
    "00001111", -- 2266 - 0x8da  :   15 - 0xf
    "00011111", -- 2267 - 0x8db  :   31 - 0x1f
    "00100111", -- 2268 - 0x8dc  :   39 - 0x27
    "00000011", -- 2269 - 0x8dd  :    3 - 0x3
    "00000011", -- 2270 - 0x8de  :    3 - 0x3
    "01000011", -- 2271 - 0x8df  :   67 - 0x43
    "00000000", -- 2272 - 0x8e0  :    0 - 0x0 -- Background 0x1c
    "11000000", -- 2273 - 0x8e1  :  192 - 0xc0
    "11110000", -- 2274 - 0x8e2  :  240 - 0xf0
    "11111000", -- 2275 - 0x8e3  :  248 - 0xf8
    "10011100", -- 2276 - 0x8e4  :  156 - 0x9c
    "00001100", -- 2277 - 0x8e5  :   12 - 0xc
    "00001100", -- 2278 - 0x8e6  :   12 - 0xc
    "00001110", -- 2279 - 0x8e7  :   14 - 0xe
    "01100111", -- 2280 - 0x8e8  :  103 - 0x67 -- Background 0x1d
    "01111111", -- 2281 - 0x8e9  :  127 - 0x7f
    "01111111", -- 2282 - 0x8ea  :  127 - 0x7f
    "01111111", -- 2283 - 0x8eb  :  127 - 0x7f
    "01101110", -- 2284 - 0x8ec  :  110 - 0x6e
    "01000110", -- 2285 - 0x8ed  :   70 - 0x46
    "00000000", -- 2286 - 0x8ee  :    0 - 0x0
    "00000000", -- 2287 - 0x8ef  :    0 - 0x0
    "01100111", -- 2288 - 0x8f0  :  103 - 0x67 -- Background 0x1e
    "01111111", -- 2289 - 0x8f1  :  127 - 0x7f
    "01111111", -- 2290 - 0x8f2  :  127 - 0x7f
    "01111111", -- 2291 - 0x8f3  :  127 - 0x7f
    "01111011", -- 2292 - 0x8f4  :  123 - 0x7b
    "00110001", -- 2293 - 0x8f5  :   49 - 0x31
    "00000000", -- 2294 - 0x8f6  :    0 - 0x0
    "00000000", -- 2295 - 0x8f7  :    0 - 0x0
    "10011110", -- 2296 - 0x8f8  :  158 - 0x9e -- Background 0x1f
    "11111110", -- 2297 - 0x8f9  :  254 - 0xfe
    "11111110", -- 2298 - 0x8fa  :  254 - 0xfe
    "11111110", -- 2299 - 0x8fb  :  254 - 0xfe
    "01110110", -- 2300 - 0x8fc  :  118 - 0x76
    "01100010", -- 2301 - 0x8fd  :   98 - 0x62
    "00000000", -- 2302 - 0x8fe  :    0 - 0x0
    "00000000", -- 2303 - 0x8ff  :    0 - 0x0
    "10011110", -- 2304 - 0x900  :  158 - 0x9e -- Background 0x20
    "11111110", -- 2305 - 0x901  :  254 - 0xfe
    "11111110", -- 2306 - 0x902  :  254 - 0xfe
    "11111110", -- 2307 - 0x903  :  254 - 0xfe
    "11011110", -- 2308 - 0x904  :  222 - 0xde
    "10001100", -- 2309 - 0x905  :  140 - 0x8c
    "00000000", -- 2310 - 0x906  :    0 - 0x0
    "00000000", -- 2311 - 0x907  :    0 - 0x0
    "00000000", -- 2312 - 0x908  :    0 - 0x0 -- Background 0x21
    "00000011", -- 2313 - 0x909  :    3 - 0x3
    "00001111", -- 2314 - 0x90a  :   15 - 0xf
    "00011111", -- 2315 - 0x90b  :   31 - 0x1f
    "00111111", -- 2316 - 0x90c  :   63 - 0x3f
    "00110011", -- 2317 - 0x90d  :   51 - 0x33
    "00100001", -- 2318 - 0x90e  :   33 - 0x21
    "01100001", -- 2319 - 0x90f  :   97 - 0x61
    "01100001", -- 2320 - 0x910  :   97 - 0x61 -- Background 0x22
    "01110011", -- 2321 - 0x911  :  115 - 0x73
    "01111111", -- 2322 - 0x912  :  127 - 0x7f
    "01111111", -- 2323 - 0x913  :  127 - 0x7f
    "01101110", -- 2324 - 0x914  :  110 - 0x6e
    "01000110", -- 2325 - 0x915  :   70 - 0x46
    "00000000", -- 2326 - 0x916  :    0 - 0x0
    "00000000", -- 2327 - 0x917  :    0 - 0x0
    "01100001", -- 2328 - 0x918  :   97 - 0x61 -- Background 0x23
    "01110011", -- 2329 - 0x919  :  115 - 0x73
    "01111111", -- 2330 - 0x91a  :  127 - 0x7f
    "01111111", -- 2331 - 0x91b  :  127 - 0x7f
    "01110111", -- 2332 - 0x91c  :  119 - 0x77
    "00100011", -- 2333 - 0x91d  :   35 - 0x23
    "00000000", -- 2334 - 0x91e  :    0 - 0x0
    "00000000", -- 2335 - 0x91f  :    0 - 0x0
    "00000000", -- 2336 - 0x920  :    0 - 0x0 -- Background 0x24
    "00000011", -- 2337 - 0x921  :    3 - 0x3
    "00001111", -- 2338 - 0x922  :   15 - 0xf
    "00011111", -- 2339 - 0x923  :   31 - 0x1f
    "00111111", -- 2340 - 0x924  :   63 - 0x3f
    "00111111", -- 2341 - 0x925  :   63 - 0x3f
    "00111111", -- 2342 - 0x926  :   63 - 0x3f
    "01111111", -- 2343 - 0x927  :  127 - 0x7f
    "01111111", -- 2344 - 0x928  :  127 - 0x7f -- Background 0x25
    "01111111", -- 2345 - 0x929  :  127 - 0x7f
    "01111111", -- 2346 - 0x92a  :  127 - 0x7f
    "01111111", -- 2347 - 0x92b  :  127 - 0x7f
    "01101110", -- 2348 - 0x92c  :  110 - 0x6e
    "01000110", -- 2349 - 0x92d  :   70 - 0x46
    "00000000", -- 2350 - 0x92e  :    0 - 0x0
    "00000000", -- 2351 - 0x92f  :    0 - 0x0
    "01111111", -- 2352 - 0x930  :  127 - 0x7f -- Background 0x26
    "01111111", -- 2353 - 0x931  :  127 - 0x7f
    "01111111", -- 2354 - 0x932  :  127 - 0x7f
    "01111111", -- 2355 - 0x933  :  127 - 0x7f
    "01111011", -- 2356 - 0x934  :  123 - 0x7b
    "00110001", -- 2357 - 0x935  :   49 - 0x31
    "00000000", -- 2358 - 0x936  :    0 - 0x0
    "00000000", -- 2359 - 0x937  :    0 - 0x0
    "00000000", -- 2360 - 0x938  :    0 - 0x0 -- Background 0x27
    "00000000", -- 2361 - 0x939  :    0 - 0x0
    "00000000", -- 2362 - 0x93a  :    0 - 0x0
    "00000000", -- 2363 - 0x93b  :    0 - 0x0
    "00000000", -- 2364 - 0x93c  :    0 - 0x0
    "00000000", -- 2365 - 0x93d  :    0 - 0x0
    "00000000", -- 2366 - 0x93e  :    0 - 0x0
    "00000000", -- 2367 - 0x93f  :    0 - 0x0
    "00000000", -- 2368 - 0x940  :    0 - 0x0 -- Background 0x28
    "00000000", -- 2369 - 0x941  :    0 - 0x0
    "00000000", -- 2370 - 0x942  :    0 - 0x0
    "00000000", -- 2371 - 0x943  :    0 - 0x0
    "00000000", -- 2372 - 0x944  :    0 - 0x0
    "00000000", -- 2373 - 0x945  :    0 - 0x0
    "00000000", -- 2374 - 0x946  :    0 - 0x0
    "00000000", -- 2375 - 0x947  :    0 - 0x0
    "00000000", -- 2376 - 0x948  :    0 - 0x0 -- Background 0x29
    "00000000", -- 2377 - 0x949  :    0 - 0x0
    "00000000", -- 2378 - 0x94a  :    0 - 0x0
    "00000000", -- 2379 - 0x94b  :    0 - 0x0
    "00000000", -- 2380 - 0x94c  :    0 - 0x0
    "00000000", -- 2381 - 0x94d  :    0 - 0x0
    "00000000", -- 2382 - 0x94e  :    0 - 0x0
    "00000000", -- 2383 - 0x94f  :    0 - 0x0
    "00000000", -- 2384 - 0x950  :    0 - 0x0 -- Background 0x2a
    "00000000", -- 2385 - 0x951  :    0 - 0x0
    "00000000", -- 2386 - 0x952  :    0 - 0x0
    "00000000", -- 2387 - 0x953  :    0 - 0x0
    "00000000", -- 2388 - 0x954  :    0 - 0x0
    "00000000", -- 2389 - 0x955  :    0 - 0x0
    "00000000", -- 2390 - 0x956  :    0 - 0x0
    "00000000", -- 2391 - 0x957  :    0 - 0x0
    "00000000", -- 2392 - 0x958  :    0 - 0x0 -- Background 0x2b
    "00000000", -- 2393 - 0x959  :    0 - 0x0
    "00000000", -- 2394 - 0x95a  :    0 - 0x0
    "00000000", -- 2395 - 0x95b  :    0 - 0x0
    "00000000", -- 2396 - 0x95c  :    0 - 0x0
    "00000000", -- 2397 - 0x95d  :    0 - 0x0
    "00000000", -- 2398 - 0x95e  :    0 - 0x0
    "00000000", -- 2399 - 0x95f  :    0 - 0x0
    "00000000", -- 2400 - 0x960  :    0 - 0x0 -- Background 0x2c
    "00000000", -- 2401 - 0x961  :    0 - 0x0
    "00000000", -- 2402 - 0x962  :    0 - 0x0
    "00000000", -- 2403 - 0x963  :    0 - 0x0
    "00000000", -- 2404 - 0x964  :    0 - 0x0
    "00000000", -- 2405 - 0x965  :    0 - 0x0
    "00000000", -- 2406 - 0x966  :    0 - 0x0
    "00000000", -- 2407 - 0x967  :    0 - 0x0
    "00000000", -- 2408 - 0x968  :    0 - 0x0 -- Background 0x2d
    "00000000", -- 2409 - 0x969  :    0 - 0x0
    "00000000", -- 2410 - 0x96a  :    0 - 0x0
    "00000000", -- 2411 - 0x96b  :    0 - 0x0
    "00000000", -- 2412 - 0x96c  :    0 - 0x0
    "00000000", -- 2413 - 0x96d  :    0 - 0x0
    "00000000", -- 2414 - 0x96e  :    0 - 0x0
    "00000000", -- 2415 - 0x96f  :    0 - 0x0
    "00000000", -- 2416 - 0x970  :    0 - 0x0 -- Background 0x2e
    "00000000", -- 2417 - 0x971  :    0 - 0x0
    "00000000", -- 2418 - 0x972  :    0 - 0x0
    "00000000", -- 2419 - 0x973  :    0 - 0x0
    "00000000", -- 2420 - 0x974  :    0 - 0x0
    "00000000", -- 2421 - 0x975  :    0 - 0x0
    "00000000", -- 2422 - 0x976  :    0 - 0x0
    "00000000", -- 2423 - 0x977  :    0 - 0x0
    "00000000", -- 2424 - 0x978  :    0 - 0x0 -- Background 0x2f
    "00000000", -- 2425 - 0x979  :    0 - 0x0
    "00000000", -- 2426 - 0x97a  :    0 - 0x0
    "00000000", -- 2427 - 0x97b  :    0 - 0x0
    "00000000", -- 2428 - 0x97c  :    0 - 0x0
    "00000000", -- 2429 - 0x97d  :    0 - 0x0
    "00000000", -- 2430 - 0x97e  :    0 - 0x0
    "00000000", -- 2431 - 0x97f  :    0 - 0x0
    "00000000", -- 2432 - 0x980  :    0 - 0x0 -- Background 0x30
    "00000000", -- 2433 - 0x981  :    0 - 0x0
    "00000000", -- 2434 - 0x982  :    0 - 0x0
    "00000000", -- 2435 - 0x983  :    0 - 0x0
    "00000000", -- 2436 - 0x984  :    0 - 0x0
    "00000000", -- 2437 - 0x985  :    0 - 0x0
    "00000000", -- 2438 - 0x986  :    0 - 0x0
    "00000000", -- 2439 - 0x987  :    0 - 0x0
    "00000000", -- 2440 - 0x988  :    0 - 0x0 -- Background 0x31
    "00000000", -- 2441 - 0x989  :    0 - 0x0
    "00000000", -- 2442 - 0x98a  :    0 - 0x0
    "00000000", -- 2443 - 0x98b  :    0 - 0x0
    "00000000", -- 2444 - 0x98c  :    0 - 0x0
    "00000000", -- 2445 - 0x98d  :    0 - 0x0
    "00000000", -- 2446 - 0x98e  :    0 - 0x0
    "00000000", -- 2447 - 0x98f  :    0 - 0x0
    "00000000", -- 2448 - 0x990  :    0 - 0x0 -- Background 0x32
    "00000000", -- 2449 - 0x991  :    0 - 0x0
    "00000000", -- 2450 - 0x992  :    0 - 0x0
    "00000000", -- 2451 - 0x993  :    0 - 0x0
    "00000000", -- 2452 - 0x994  :    0 - 0x0
    "00000000", -- 2453 - 0x995  :    0 - 0x0
    "00000000", -- 2454 - 0x996  :    0 - 0x0
    "00000000", -- 2455 - 0x997  :    0 - 0x0
    "00000000", -- 2456 - 0x998  :    0 - 0x0 -- Background 0x33
    "00000000", -- 2457 - 0x999  :    0 - 0x0
    "00000000", -- 2458 - 0x99a  :    0 - 0x0
    "00000000", -- 2459 - 0x99b  :    0 - 0x0
    "00000000", -- 2460 - 0x99c  :    0 - 0x0
    "00000000", -- 2461 - 0x99d  :    0 - 0x0
    "00000000", -- 2462 - 0x99e  :    0 - 0x0
    "00000000", -- 2463 - 0x99f  :    0 - 0x0
    "00000000", -- 2464 - 0x9a0  :    0 - 0x0 -- Background 0x34
    "00000000", -- 2465 - 0x9a1  :    0 - 0x0
    "00000000", -- 2466 - 0x9a2  :    0 - 0x0
    "00000000", -- 2467 - 0x9a3  :    0 - 0x0
    "00000000", -- 2468 - 0x9a4  :    0 - 0x0
    "00000000", -- 2469 - 0x9a5  :    0 - 0x0
    "00000000", -- 2470 - 0x9a6  :    0 - 0x0
    "00000000", -- 2471 - 0x9a7  :    0 - 0x0
    "00000000", -- 2472 - 0x9a8  :    0 - 0x0 -- Background 0x35
    "00000000", -- 2473 - 0x9a9  :    0 - 0x0
    "00000000", -- 2474 - 0x9aa  :    0 - 0x0
    "00000000", -- 2475 - 0x9ab  :    0 - 0x0
    "00000000", -- 2476 - 0x9ac  :    0 - 0x0
    "00000000", -- 2477 - 0x9ad  :    0 - 0x0
    "00000000", -- 2478 - 0x9ae  :    0 - 0x0
    "00000000", -- 2479 - 0x9af  :    0 - 0x0
    "00000000", -- 2480 - 0x9b0  :    0 - 0x0 -- Background 0x36
    "00000000", -- 2481 - 0x9b1  :    0 - 0x0
    "00000000", -- 2482 - 0x9b2  :    0 - 0x0
    "00000000", -- 2483 - 0x9b3  :    0 - 0x0
    "00000000", -- 2484 - 0x9b4  :    0 - 0x0
    "00000000", -- 2485 - 0x9b5  :    0 - 0x0
    "00000000", -- 2486 - 0x9b6  :    0 - 0x0
    "00000000", -- 2487 - 0x9b7  :    0 - 0x0
    "00000000", -- 2488 - 0x9b8  :    0 - 0x0 -- Background 0x37
    "00000000", -- 2489 - 0x9b9  :    0 - 0x0
    "00000000", -- 2490 - 0x9ba  :    0 - 0x0
    "00000000", -- 2491 - 0x9bb  :    0 - 0x0
    "00000000", -- 2492 - 0x9bc  :    0 - 0x0
    "00000000", -- 2493 - 0x9bd  :    0 - 0x0
    "00000000", -- 2494 - 0x9be  :    0 - 0x0
    "00000000", -- 2495 - 0x9bf  :    0 - 0x0
    "00000000", -- 2496 - 0x9c0  :    0 - 0x0 -- Background 0x38
    "00000000", -- 2497 - 0x9c1  :    0 - 0x0
    "00000000", -- 2498 - 0x9c2  :    0 - 0x0
    "00000000", -- 2499 - 0x9c3  :    0 - 0x0
    "00000000", -- 2500 - 0x9c4  :    0 - 0x0
    "00000000", -- 2501 - 0x9c5  :    0 - 0x0
    "00000000", -- 2502 - 0x9c6  :    0 - 0x0
    "00000000", -- 2503 - 0x9c7  :    0 - 0x0
    "00000000", -- 2504 - 0x9c8  :    0 - 0x0 -- Background 0x39
    "00000000", -- 2505 - 0x9c9  :    0 - 0x0
    "00000000", -- 2506 - 0x9ca  :    0 - 0x0
    "00000000", -- 2507 - 0x9cb  :    0 - 0x0
    "00000000", -- 2508 - 0x9cc  :    0 - 0x0
    "00000000", -- 2509 - 0x9cd  :    0 - 0x0
    "00000000", -- 2510 - 0x9ce  :    0 - 0x0
    "00000000", -- 2511 - 0x9cf  :    0 - 0x0
    "00000000", -- 2512 - 0x9d0  :    0 - 0x0 -- Background 0x3a
    "00000000", -- 2513 - 0x9d1  :    0 - 0x0
    "00000000", -- 2514 - 0x9d2  :    0 - 0x0
    "00000000", -- 2515 - 0x9d3  :    0 - 0x0
    "00000000", -- 2516 - 0x9d4  :    0 - 0x0
    "00000000", -- 2517 - 0x9d5  :    0 - 0x0
    "00000000", -- 2518 - 0x9d6  :    0 - 0x0
    "00000000", -- 2519 - 0x9d7  :    0 - 0x0
    "00000000", -- 2520 - 0x9d8  :    0 - 0x0 -- Background 0x3b
    "00000000", -- 2521 - 0x9d9  :    0 - 0x0
    "00000000", -- 2522 - 0x9da  :    0 - 0x0
    "00000000", -- 2523 - 0x9db  :    0 - 0x0
    "00000000", -- 2524 - 0x9dc  :    0 - 0x0
    "00000000", -- 2525 - 0x9dd  :    0 - 0x0
    "00000000", -- 2526 - 0x9de  :    0 - 0x0
    "00000000", -- 2527 - 0x9df  :    0 - 0x0
    "00000000", -- 2528 - 0x9e0  :    0 - 0x0 -- Background 0x3c
    "00000000", -- 2529 - 0x9e1  :    0 - 0x0
    "00000000", -- 2530 - 0x9e2  :    0 - 0x0
    "00000000", -- 2531 - 0x9e3  :    0 - 0x0
    "00000000", -- 2532 - 0x9e4  :    0 - 0x0
    "00000000", -- 2533 - 0x9e5  :    0 - 0x0
    "00000000", -- 2534 - 0x9e6  :    0 - 0x0
    "00000000", -- 2535 - 0x9e7  :    0 - 0x0
    "00000000", -- 2536 - 0x9e8  :    0 - 0x0 -- Background 0x3d
    "00000000", -- 2537 - 0x9e9  :    0 - 0x0
    "00000000", -- 2538 - 0x9ea  :    0 - 0x0
    "00000000", -- 2539 - 0x9eb  :    0 - 0x0
    "00000000", -- 2540 - 0x9ec  :    0 - 0x0
    "00000000", -- 2541 - 0x9ed  :    0 - 0x0
    "00000000", -- 2542 - 0x9ee  :    0 - 0x0
    "00000000", -- 2543 - 0x9ef  :    0 - 0x0
    "00000000", -- 2544 - 0x9f0  :    0 - 0x0 -- Background 0x3e
    "00000000", -- 2545 - 0x9f1  :    0 - 0x0
    "00000000", -- 2546 - 0x9f2  :    0 - 0x0
    "00000000", -- 2547 - 0x9f3  :    0 - 0x0
    "00000000", -- 2548 - 0x9f4  :    0 - 0x0
    "00000000", -- 2549 - 0x9f5  :    0 - 0x0
    "00000000", -- 2550 - 0x9f6  :    0 - 0x0
    "00000000", -- 2551 - 0x9f7  :    0 - 0x0
    "00000000", -- 2552 - 0x9f8  :    0 - 0x0 -- Background 0x3f
    "00000000", -- 2553 - 0x9f9  :    0 - 0x0
    "00000000", -- 2554 - 0x9fa  :    0 - 0x0
    "00000000", -- 2555 - 0x9fb  :    0 - 0x0
    "00000000", -- 2556 - 0x9fc  :    0 - 0x0
    "00000000", -- 2557 - 0x9fd  :    0 - 0x0
    "00000000", -- 2558 - 0x9fe  :    0 - 0x0
    "00000000", -- 2559 - 0x9ff  :    0 - 0x0
    "00000000", -- 2560 - 0xa00  :    0 - 0x0 -- Background 0x40
    "00000000", -- 2561 - 0xa01  :    0 - 0x0
    "00000000", -- 2562 - 0xa02  :    0 - 0x0
    "00000000", -- 2563 - 0xa03  :    0 - 0x0
    "00000000", -- 2564 - 0xa04  :    0 - 0x0
    "00000000", -- 2565 - 0xa05  :    0 - 0x0
    "00000000", -- 2566 - 0xa06  :    0 - 0x0
    "00000000", -- 2567 - 0xa07  :    0 - 0x0
    "00000000", -- 2568 - 0xa08  :    0 - 0x0 -- Background 0x41
    "00000000", -- 2569 - 0xa09  :    0 - 0x0
    "00000000", -- 2570 - 0xa0a  :    0 - 0x0
    "00000000", -- 2571 - 0xa0b  :    0 - 0x0
    "00000000", -- 2572 - 0xa0c  :    0 - 0x0
    "00000000", -- 2573 - 0xa0d  :    0 - 0x0
    "00000000", -- 2574 - 0xa0e  :    0 - 0x0
    "00000000", -- 2575 - 0xa0f  :    0 - 0x0
    "00000000", -- 2576 - 0xa10  :    0 - 0x0 -- Background 0x42
    "00000000", -- 2577 - 0xa11  :    0 - 0x0
    "00000000", -- 2578 - 0xa12  :    0 - 0x0
    "00000000", -- 2579 - 0xa13  :    0 - 0x0
    "00000000", -- 2580 - 0xa14  :    0 - 0x0
    "00000000", -- 2581 - 0xa15  :    0 - 0x0
    "00000000", -- 2582 - 0xa16  :    0 - 0x0
    "00000000", -- 2583 - 0xa17  :    0 - 0x0
    "00000000", -- 2584 - 0xa18  :    0 - 0x0 -- Background 0x43
    "00000000", -- 2585 - 0xa19  :    0 - 0x0
    "00000000", -- 2586 - 0xa1a  :    0 - 0x0
    "00000000", -- 2587 - 0xa1b  :    0 - 0x0
    "00000000", -- 2588 - 0xa1c  :    0 - 0x0
    "00000000", -- 2589 - 0xa1d  :    0 - 0x0
    "00000000", -- 2590 - 0xa1e  :    0 - 0x0
    "00000000", -- 2591 - 0xa1f  :    0 - 0x0
    "00000000", -- 2592 - 0xa20  :    0 - 0x0 -- Background 0x44
    "00000000", -- 2593 - 0xa21  :    0 - 0x0
    "00000000", -- 2594 - 0xa22  :    0 - 0x0
    "00000000", -- 2595 - 0xa23  :    0 - 0x0
    "00000000", -- 2596 - 0xa24  :    0 - 0x0
    "00000000", -- 2597 - 0xa25  :    0 - 0x0
    "00000000", -- 2598 - 0xa26  :    0 - 0x0
    "00000000", -- 2599 - 0xa27  :    0 - 0x0
    "00000000", -- 2600 - 0xa28  :    0 - 0x0 -- Background 0x45
    "00000000", -- 2601 - 0xa29  :    0 - 0x0
    "00000000", -- 2602 - 0xa2a  :    0 - 0x0
    "00000000", -- 2603 - 0xa2b  :    0 - 0x0
    "00000000", -- 2604 - 0xa2c  :    0 - 0x0
    "00000000", -- 2605 - 0xa2d  :    0 - 0x0
    "00000000", -- 2606 - 0xa2e  :    0 - 0x0
    "00000000", -- 2607 - 0xa2f  :    0 - 0x0
    "00000000", -- 2608 - 0xa30  :    0 - 0x0 -- Background 0x46
    "00000000", -- 2609 - 0xa31  :    0 - 0x0
    "00000000", -- 2610 - 0xa32  :    0 - 0x0
    "00000000", -- 2611 - 0xa33  :    0 - 0x0
    "00000000", -- 2612 - 0xa34  :    0 - 0x0
    "00000000", -- 2613 - 0xa35  :    0 - 0x0
    "00000000", -- 2614 - 0xa36  :    0 - 0x0
    "00000000", -- 2615 - 0xa37  :    0 - 0x0
    "00000000", -- 2616 - 0xa38  :    0 - 0x0 -- Background 0x47
    "00000000", -- 2617 - 0xa39  :    0 - 0x0
    "00000000", -- 2618 - 0xa3a  :    0 - 0x0
    "00000000", -- 2619 - 0xa3b  :    0 - 0x0
    "00000000", -- 2620 - 0xa3c  :    0 - 0x0
    "00000000", -- 2621 - 0xa3d  :    0 - 0x0
    "00000000", -- 2622 - 0xa3e  :    0 - 0x0
    "00000000", -- 2623 - 0xa3f  :    0 - 0x0
    "00000000", -- 2624 - 0xa40  :    0 - 0x0 -- Background 0x48
    "00000000", -- 2625 - 0xa41  :    0 - 0x0
    "00000000", -- 2626 - 0xa42  :    0 - 0x0
    "00000000", -- 2627 - 0xa43  :    0 - 0x0
    "00000000", -- 2628 - 0xa44  :    0 - 0x0
    "00000000", -- 2629 - 0xa45  :    0 - 0x0
    "00000000", -- 2630 - 0xa46  :    0 - 0x0
    "00000000", -- 2631 - 0xa47  :    0 - 0x0
    "00000000", -- 2632 - 0xa48  :    0 - 0x0 -- Background 0x49
    "00000000", -- 2633 - 0xa49  :    0 - 0x0
    "00000000", -- 2634 - 0xa4a  :    0 - 0x0
    "00000000", -- 2635 - 0xa4b  :    0 - 0x0
    "00000000", -- 2636 - 0xa4c  :    0 - 0x0
    "00000000", -- 2637 - 0xa4d  :    0 - 0x0
    "00000000", -- 2638 - 0xa4e  :    0 - 0x0
    "00000000", -- 2639 - 0xa4f  :    0 - 0x0
    "00000000", -- 2640 - 0xa50  :    0 - 0x0 -- Background 0x4a
    "00000000", -- 2641 - 0xa51  :    0 - 0x0
    "00000000", -- 2642 - 0xa52  :    0 - 0x0
    "00000000", -- 2643 - 0xa53  :    0 - 0x0
    "00000000", -- 2644 - 0xa54  :    0 - 0x0
    "00000000", -- 2645 - 0xa55  :    0 - 0x0
    "00000000", -- 2646 - 0xa56  :    0 - 0x0
    "00000000", -- 2647 - 0xa57  :    0 - 0x0
    "00000000", -- 2648 - 0xa58  :    0 - 0x0 -- Background 0x4b
    "00000000", -- 2649 - 0xa59  :    0 - 0x0
    "00000000", -- 2650 - 0xa5a  :    0 - 0x0
    "00000000", -- 2651 - 0xa5b  :    0 - 0x0
    "00000000", -- 2652 - 0xa5c  :    0 - 0x0
    "00000000", -- 2653 - 0xa5d  :    0 - 0x0
    "00000000", -- 2654 - 0xa5e  :    0 - 0x0
    "00000000", -- 2655 - 0xa5f  :    0 - 0x0
    "00000000", -- 2656 - 0xa60  :    0 - 0x0 -- Background 0x4c
    "00000000", -- 2657 - 0xa61  :    0 - 0x0
    "00000000", -- 2658 - 0xa62  :    0 - 0x0
    "00000000", -- 2659 - 0xa63  :    0 - 0x0
    "00000000", -- 2660 - 0xa64  :    0 - 0x0
    "00000000", -- 2661 - 0xa65  :    0 - 0x0
    "00000000", -- 2662 - 0xa66  :    0 - 0x0
    "00000000", -- 2663 - 0xa67  :    0 - 0x0
    "00000000", -- 2664 - 0xa68  :    0 - 0x0 -- Background 0x4d
    "00000000", -- 2665 - 0xa69  :    0 - 0x0
    "00000000", -- 2666 - 0xa6a  :    0 - 0x0
    "00000001", -- 2667 - 0xa6b  :    1 - 0x1
    "00000011", -- 2668 - 0xa6c  :    3 - 0x3
    "00000111", -- 2669 - 0xa6d  :    7 - 0x7
    "00001111", -- 2670 - 0xa6e  :   15 - 0xf
    "00011111", -- 2671 - 0xa6f  :   31 - 0x1f
    "00000000", -- 2672 - 0xa70  :    0 - 0x0 -- Background 0x4e
    "00001111", -- 2673 - 0xa71  :   15 - 0xf
    "01111111", -- 2674 - 0xa72  :  127 - 0x7f
    "11111111", -- 2675 - 0xa73  :  255 - 0xff
    "11111111", -- 2676 - 0xa74  :  255 - 0xff
    "11111111", -- 2677 - 0xa75  :  255 - 0xff
    "11111111", -- 2678 - 0xa76  :  255 - 0xff
    "11111111", -- 2679 - 0xa77  :  255 - 0xff
    "00011111", -- 2680 - 0xa78  :   31 - 0x1f -- Background 0x4f
    "00111111", -- 2681 - 0xa79  :   63 - 0x3f
    "00111111", -- 2682 - 0xa7a  :   63 - 0x3f
    "00111111", -- 2683 - 0xa7b  :   63 - 0x3f
    "01111111", -- 2684 - 0xa7c  :  127 - 0x7f
    "01111111", -- 2685 - 0xa7d  :  127 - 0x7f
    "01111111", -- 2686 - 0xa7e  :  127 - 0x7f
    "01111111", -- 2687 - 0xa7f  :  127 - 0x7f
    "11111111", -- 2688 - 0xa80  :  255 - 0xff -- Background 0x50
    "11111111", -- 2689 - 0xa81  :  255 - 0xff
    "11111111", -- 2690 - 0xa82  :  255 - 0xff
    "11111111", -- 2691 - 0xa83  :  255 - 0xff
    "11111111", -- 2692 - 0xa84  :  255 - 0xff
    "11111111", -- 2693 - 0xa85  :  255 - 0xff
    "11111111", -- 2694 - 0xa86  :  255 - 0xff
    "11111111", -- 2695 - 0xa87  :  255 - 0xff
    "11111111", -- 2696 - 0xa88  :  255 - 0xff -- Background 0x51
    "11111111", -- 2697 - 0xa89  :  255 - 0xff
    "11111111", -- 2698 - 0xa8a  :  255 - 0xff
    "11111111", -- 2699 - 0xa8b  :  255 - 0xff
    "11111111", -- 2700 - 0xa8c  :  255 - 0xff
    "11111111", -- 2701 - 0xa8d  :  255 - 0xff
    "11111111", -- 2702 - 0xa8e  :  255 - 0xff
    "11111110", -- 2703 - 0xa8f  :  254 - 0xfe
    "00000000", -- 2704 - 0xa90  :    0 - 0x0 -- Background 0x52
    "00000000", -- 2705 - 0xa91  :    0 - 0x0
    "00000000", -- 2706 - 0xa92  :    0 - 0x0
    "10000000", -- 2707 - 0xa93  :  128 - 0x80
    "11000000", -- 2708 - 0xa94  :  192 - 0xc0
    "11100000", -- 2709 - 0xa95  :  224 - 0xe0
    "11110000", -- 2710 - 0xa96  :  240 - 0xf0
    "11110000", -- 2711 - 0xa97  :  240 - 0xf0
    "11111111", -- 2712 - 0xa98  :  255 - 0xff -- Background 0x53
    "11111111", -- 2713 - 0xa99  :  255 - 0xff
    "11111110", -- 2714 - 0xa9a  :  254 - 0xfe
    "11111100", -- 2715 - 0xa9b  :  252 - 0xfc
    "11110000", -- 2716 - 0xa9c  :  240 - 0xf0
    "11100000", -- 2717 - 0xa9d  :  224 - 0xe0
    "10000000", -- 2718 - 0xa9e  :  128 - 0x80
    "00000000", -- 2719 - 0xa9f  :    0 - 0x0
    "11000000", -- 2720 - 0xaa0  :  192 - 0xc0 -- Background 0x54
    "10000000", -- 2721 - 0xaa1  :  128 - 0x80
    "00000000", -- 2722 - 0xaa2  :    0 - 0x0
    "00000000", -- 2723 - 0xaa3  :    0 - 0x0
    "00000000", -- 2724 - 0xaa4  :    0 - 0x0
    "00000000", -- 2725 - 0xaa5  :    0 - 0x0
    "00000000", -- 2726 - 0xaa6  :    0 - 0x0
    "00000000", -- 2727 - 0xaa7  :    0 - 0x0
    "00000000", -- 2728 - 0xaa8  :    0 - 0x0 -- Background 0x55
    "11110000", -- 2729 - 0xaa9  :  240 - 0xf0
    "11111110", -- 2730 - 0xaaa  :  254 - 0xfe
    "11111110", -- 2731 - 0xaab  :  254 - 0xfe
    "11111110", -- 2732 - 0xaac  :  254 - 0xfe
    "11111100", -- 2733 - 0xaad  :  252 - 0xfc
    "11111000", -- 2734 - 0xaae  :  248 - 0xf8
    "11111000", -- 2735 - 0xaaf  :  248 - 0xf8
    "11110000", -- 2736 - 0xab0  :  240 - 0xf0 -- Background 0x56
    "11100000", -- 2737 - 0xab1  :  224 - 0xe0
    "11100000", -- 2738 - 0xab2  :  224 - 0xe0
    "11000000", -- 2739 - 0xab3  :  192 - 0xc0
    "10000000", -- 2740 - 0xab4  :  128 - 0x80
    "10000000", -- 2741 - 0xab5  :  128 - 0x80
    "00000000", -- 2742 - 0xab6  :    0 - 0x0
    "00000000", -- 2743 - 0xab7  :    0 - 0x0
    "00000000", -- 2744 - 0xab8  :    0 - 0x0 -- Background 0x57
    "00000000", -- 2745 - 0xab9  :    0 - 0x0
    "00000000", -- 2746 - 0xaba  :    0 - 0x0
    "00000000", -- 2747 - 0xabb  :    0 - 0x0
    "00000000", -- 2748 - 0xabc  :    0 - 0x0
    "00000000", -- 2749 - 0xabd  :    0 - 0x0
    "00000000", -- 2750 - 0xabe  :    0 - 0x0
    "00000100", -- 2751 - 0xabf  :    4 - 0x4
    "00000110", -- 2752 - 0xac0  :    6 - 0x6 -- Background 0x58
    "00000110", -- 2753 - 0xac1  :    6 - 0x6
    "00000111", -- 2754 - 0xac2  :    7 - 0x7
    "00000111", -- 2755 - 0xac3  :    7 - 0x7
    "00000111", -- 2756 - 0xac4  :    7 - 0x7
    "00000111", -- 2757 - 0xac5  :    7 - 0x7
    "00000000", -- 2758 - 0xac6  :    0 - 0x0
    "00000000", -- 2759 - 0xac7  :    0 - 0x0
    "00000000", -- 2760 - 0xac8  :    0 - 0x0 -- Background 0x59
    "00000000", -- 2761 - 0xac9  :    0 - 0x0
    "00000000", -- 2762 - 0xaca  :    0 - 0x0
    "00000000", -- 2763 - 0xacb  :    0 - 0x0
    "00000000", -- 2764 - 0xacc  :    0 - 0x0
    "00000000", -- 2765 - 0xacd  :    0 - 0x0
    "00000000", -- 2766 - 0xace  :    0 - 0x0
    "00010000", -- 2767 - 0xacf  :   16 - 0x10
    "00011100", -- 2768 - 0xad0  :   28 - 0x1c -- Background 0x5a
    "00011110", -- 2769 - 0xad1  :   30 - 0x1e
    "00011111", -- 2770 - 0xad2  :   31 - 0x1f
    "00011111", -- 2771 - 0xad3  :   31 - 0x1f
    "00011111", -- 2772 - 0xad4  :   31 - 0x1f
    "00011111", -- 2773 - 0xad5  :   31 - 0x1f
    "00000000", -- 2774 - 0xad6  :    0 - 0x0
    "00000000", -- 2775 - 0xad7  :    0 - 0x0
    "00000000", -- 2776 - 0xad8  :    0 - 0x0 -- Background 0x5b
    "00000000", -- 2777 - 0xad9  :    0 - 0x0
    "00000000", -- 2778 - 0xada  :    0 - 0x0
    "00000000", -- 2779 - 0xadb  :    0 - 0x0
    "00000000", -- 2780 - 0xadc  :    0 - 0x0
    "00000000", -- 2781 - 0xadd  :    0 - 0x0
    "00000000", -- 2782 - 0xade  :    0 - 0x0
    "11000000", -- 2783 - 0xadf  :  192 - 0xc0
    "11110000", -- 2784 - 0xae0  :  240 - 0xf0 -- Background 0x5c
    "11111100", -- 2785 - 0xae1  :  252 - 0xfc
    "11111111", -- 2786 - 0xae2  :  255 - 0xff
    "11111111", -- 2787 - 0xae3  :  255 - 0xff
    "11111111", -- 2788 - 0xae4  :  255 - 0xff
    "11111111", -- 2789 - 0xae5  :  255 - 0xff
    "00000000", -- 2790 - 0xae6  :    0 - 0x0
    "00000000", -- 2791 - 0xae7  :    0 - 0x0
    "00000000", -- 2792 - 0xae8  :    0 - 0x0 -- Background 0x5d
    "00000000", -- 2793 - 0xae9  :    0 - 0x0
    "00000001", -- 2794 - 0xaea  :    1 - 0x1
    "00000011", -- 2795 - 0xaeb  :    3 - 0x3
    "00001111", -- 2796 - 0xaec  :   15 - 0xf
    "00001111", -- 2797 - 0xaed  :   15 - 0xf
    "00000000", -- 2798 - 0xaee  :    0 - 0x0
    "00000000", -- 2799 - 0xaef  :    0 - 0x0
    "11111100", -- 2800 - 0xaf0  :  252 - 0xfc -- Background 0x5e
    "11111100", -- 2801 - 0xaf1  :  252 - 0xfc
    "11111100", -- 2802 - 0xaf2  :  252 - 0xfc
    "11111100", -- 2803 - 0xaf3  :  252 - 0xfc
    "11111000", -- 2804 - 0xaf4  :  248 - 0xf8
    "11111100", -- 2805 - 0xaf5  :  252 - 0xfc
    "00111100", -- 2806 - 0xaf6  :   60 - 0x3c
    "00000000", -- 2807 - 0xaf7  :    0 - 0x0
    "00000100", -- 2808 - 0xaf8  :    4 - 0x4 -- Background 0x5f
    "00001100", -- 2809 - 0xaf9  :   12 - 0xc
    "00011100", -- 2810 - 0xafa  :   28 - 0x1c
    "00001100", -- 2811 - 0xafb  :   12 - 0xc
    "00011000", -- 2812 - 0xafc  :   24 - 0x18
    "00111100", -- 2813 - 0xafd  :   60 - 0x3c
    "00111100", -- 2814 - 0xafe  :   60 - 0x3c
    "00000000", -- 2815 - 0xaff  :    0 - 0x0
    "00000000", -- 2816 - 0xb00  :    0 - 0x0 -- Background 0x60
    "00000011", -- 2817 - 0xb01  :    3 - 0x3
    "00001111", -- 2818 - 0xb02  :   15 - 0xf
    "00010011", -- 2819 - 0xb03  :   19 - 0x13
    "00100001", -- 2820 - 0xb04  :   33 - 0x21
    "00100001", -- 2821 - 0xb05  :   33 - 0x21
    "00100001", -- 2822 - 0xb06  :   33 - 0x21
    "01110011", -- 2823 - 0xb07  :  115 - 0x73
    "00000000", -- 2824 - 0xb08  :    0 - 0x0 -- Background 0x61
    "11000000", -- 2825 - 0xb09  :  192 - 0xc0
    "11110000", -- 2826 - 0xb0a  :  240 - 0xf0
    "11001000", -- 2827 - 0xb0b  :  200 - 0xc8
    "10000100", -- 2828 - 0xb0c  :  132 - 0x84
    "10000100", -- 2829 - 0xb0d  :  132 - 0x84
    "10000100", -- 2830 - 0xb0e  :  132 - 0x84
    "11001110", -- 2831 - 0xb0f  :  206 - 0xce
    "10010100", -- 2832 - 0xb10  :  148 - 0x94 -- Background 0x62
    "11101010", -- 2833 - 0xb11  :  234 - 0xea
    "11011110", -- 2834 - 0xb12  :  222 - 0xde
    "11101110", -- 2835 - 0xb13  :  238 - 0xee
    "11011110", -- 2836 - 0xb14  :  222 - 0xde
    "01100110", -- 2837 - 0xb15  :  102 - 0x66
    "01000010", -- 2838 - 0xb16  :   66 - 0x42
    "00000000", -- 2839 - 0xb17  :    0 - 0x0
    "10010100", -- 2840 - 0xb18  :  148 - 0x94 -- Background 0x63
    "11101010", -- 2841 - 0xb19  :  234 - 0xea
    "11011110", -- 2842 - 0xb1a  :  222 - 0xde
    "11101110", -- 2843 - 0xb1b  :  238 - 0xee
    "11011110", -- 2844 - 0xb1c  :  222 - 0xde
    "11001110", -- 2845 - 0xb1d  :  206 - 0xce
    "10001100", -- 2846 - 0xb1e  :  140 - 0x8c
    "00000000", -- 2847 - 0xb1f  :    0 - 0x0
    "00000000", -- 2848 - 0xb20  :    0 - 0x0 -- Background 0x64
    "00000000", -- 2849 - 0xb21  :    0 - 0x0
    "00000000", -- 2850 - 0xb22  :    0 - 0x0
    "00000000", -- 2851 - 0xb23  :    0 - 0x0
    "00000000", -- 2852 - 0xb24  :    0 - 0x0
    "00000000", -- 2853 - 0xb25  :    0 - 0x0
    "00000000", -- 2854 - 0xb26  :    0 - 0x0
    "00000001", -- 2855 - 0xb27  :    1 - 0x1
    "00000000", -- 2856 - 0xb28  :    0 - 0x0 -- Background 0x65
    "00000000", -- 2857 - 0xb29  :    0 - 0x0
    "00000000", -- 2858 - 0xb2a  :    0 - 0x0
    "00000000", -- 2859 - 0xb2b  :    0 - 0x0
    "00000000", -- 2860 - 0xb2c  :    0 - 0x0
    "00110110", -- 2861 - 0xb2d  :   54 - 0x36
    "00110110", -- 2862 - 0xb2e  :   54 - 0x36
    "10010000", -- 2863 - 0xb2f  :  144 - 0x90
    "00000001", -- 2864 - 0xb30  :    1 - 0x1 -- Background 0x66
    "00000011", -- 2865 - 0xb31  :    3 - 0x3
    "00000111", -- 2866 - 0xb32  :    7 - 0x7
    "00000111", -- 2867 - 0xb33  :    7 - 0x7
    "00011111", -- 2868 - 0xb34  :   31 - 0x1f
    "00011111", -- 2869 - 0xb35  :   31 - 0x1f
    "00011100", -- 2870 - 0xb36  :   28 - 0x1c
    "00000000", -- 2871 - 0xb37  :    0 - 0x0
    "11111000", -- 2872 - 0xb38  :  248 - 0xf8 -- Background 0x67
    "11111000", -- 2873 - 0xb39  :  248 - 0xf8
    "11111000", -- 2874 - 0xb3a  :  248 - 0xf8
    "11111000", -- 2875 - 0xb3b  :  248 - 0xf8
    "11111110", -- 2876 - 0xb3c  :  254 - 0xfe
    "11111110", -- 2877 - 0xb3d  :  254 - 0xfe
    "00001110", -- 2878 - 0xb3e  :   14 - 0xe
    "00000000", -- 2879 - 0xb3f  :    0 - 0x0
    "00000111", -- 2880 - 0xb40  :    7 - 0x7 -- Background 0x68
    "00001111", -- 2881 - 0xb41  :   15 - 0xf
    "00011111", -- 2882 - 0xb42  :   31 - 0x1f
    "00011111", -- 2883 - 0xb43  :   31 - 0x1f
    "00111111", -- 2884 - 0xb44  :   63 - 0x3f
    "00111111", -- 2885 - 0xb45  :   63 - 0x3f
    "00111000", -- 2886 - 0xb46  :   56 - 0x38
    "00000000", -- 2887 - 0xb47  :    0 - 0x0
    "11111000", -- 2888 - 0xb48  :  248 - 0xf8 -- Background 0x69
    "11110000", -- 2889 - 0xb49  :  240 - 0xf0
    "11110000", -- 2890 - 0xb4a  :  240 - 0xf0
    "11100000", -- 2891 - 0xb4b  :  224 - 0xe0
    "11111000", -- 2892 - 0xb4c  :  248 - 0xf8
    "11111000", -- 2893 - 0xb4d  :  248 - 0xf8
    "00111000", -- 2894 - 0xb4e  :   56 - 0x38
    "00000000", -- 2895 - 0xb4f  :    0 - 0x0
    "00000000", -- 2896 - 0xb50  :    0 - 0x0 -- Background 0x6a
    "00011111", -- 2897 - 0xb51  :   31 - 0x1f
    "01111111", -- 2898 - 0xb52  :  127 - 0x7f
    "00111111", -- 2899 - 0xb53  :   63 - 0x3f
    "00001111", -- 2900 - 0xb54  :   15 - 0xf
    "00000111", -- 2901 - 0xb55  :    7 - 0x7
    "00000000", -- 2902 - 0xb56  :    0 - 0x0
    "00000000", -- 2903 - 0xb57  :    0 - 0x0
    "00000000", -- 2904 - 0xb58  :    0 - 0x0 -- Background 0x6b
    "00000000", -- 2905 - 0xb59  :    0 - 0x0
    "11000000", -- 2906 - 0xb5a  :  192 - 0xc0
    "11110000", -- 2907 - 0xb5b  :  240 - 0xf0
    "11111000", -- 2908 - 0xb5c  :  248 - 0xf8
    "11111000", -- 2909 - 0xb5d  :  248 - 0xf8
    "11100000", -- 2910 - 0xb5e  :  224 - 0xe0
    "00000000", -- 2911 - 0xb5f  :    0 - 0x0
    "00000000", -- 2912 - 0xb60  :    0 - 0x0 -- Background 0x6c
    "00000000", -- 2913 - 0xb61  :    0 - 0x0
    "00000000", -- 2914 - 0xb62  :    0 - 0x0
    "00000000", -- 2915 - 0xb63  :    0 - 0x0
    "00000000", -- 2916 - 0xb64  :    0 - 0x0
    "00000000", -- 2917 - 0xb65  :    0 - 0x0
    "00000000", -- 2918 - 0xb66  :    0 - 0x0
    "00000000", -- 2919 - 0xb67  :    0 - 0x0
    "00000000", -- 2920 - 0xb68  :    0 - 0x0 -- Background 0x6d
    "00000000", -- 2921 - 0xb69  :    0 - 0x0
    "00000000", -- 2922 - 0xb6a  :    0 - 0x0
    "00000000", -- 2923 - 0xb6b  :    0 - 0x0
    "00000000", -- 2924 - 0xb6c  :    0 - 0x0
    "00000000", -- 2925 - 0xb6d  :    0 - 0x0
    "00000000", -- 2926 - 0xb6e  :    0 - 0x0
    "00000000", -- 2927 - 0xb6f  :    0 - 0x0
    "00000000", -- 2928 - 0xb70  :    0 - 0x0 -- Background 0x6e
    "00000000", -- 2929 - 0xb71  :    0 - 0x0
    "00000000", -- 2930 - 0xb72  :    0 - 0x0
    "00000000", -- 2931 - 0xb73  :    0 - 0x0
    "00000000", -- 2932 - 0xb74  :    0 - 0x0
    "00000000", -- 2933 - 0xb75  :    0 - 0x0
    "00000000", -- 2934 - 0xb76  :    0 - 0x0
    "00000000", -- 2935 - 0xb77  :    0 - 0x0
    "00000000", -- 2936 - 0xb78  :    0 - 0x0 -- Background 0x6f
    "00000000", -- 2937 - 0xb79  :    0 - 0x0
    "00000000", -- 2938 - 0xb7a  :    0 - 0x0
    "00000000", -- 2939 - 0xb7b  :    0 - 0x0
    "00000000", -- 2940 - 0xb7c  :    0 - 0x0
    "00000000", -- 2941 - 0xb7d  :    0 - 0x0
    "00000000", -- 2942 - 0xb7e  :    0 - 0x0
    "00000000", -- 2943 - 0xb7f  :    0 - 0x0
    "11111111", -- 2944 - 0xb80  :  255 - 0xff -- Background 0x70
    "11111111", -- 2945 - 0xb81  :  255 - 0xff
    "11111111", -- 2946 - 0xb82  :  255 - 0xff
    "11111111", -- 2947 - 0xb83  :  255 - 0xff
    "11111111", -- 2948 - 0xb84  :  255 - 0xff
    "11111111", -- 2949 - 0xb85  :  255 - 0xff
    "11111111", -- 2950 - 0xb86  :  255 - 0xff
    "11111111", -- 2951 - 0xb87  :  255 - 0xff
    "11111111", -- 2952 - 0xb88  :  255 - 0xff -- Background 0x71
    "11111111", -- 2953 - 0xb89  :  255 - 0xff
    "11111111", -- 2954 - 0xb8a  :  255 - 0xff
    "11111111", -- 2955 - 0xb8b  :  255 - 0xff
    "11111111", -- 2956 - 0xb8c  :  255 - 0xff
    "11111111", -- 2957 - 0xb8d  :  255 - 0xff
    "11111111", -- 2958 - 0xb8e  :  255 - 0xff
    "11111111", -- 2959 - 0xb8f  :  255 - 0xff
    "11111111", -- 2960 - 0xb90  :  255 - 0xff -- Background 0x72
    "11111111", -- 2961 - 0xb91  :  255 - 0xff
    "11111111", -- 2962 - 0xb92  :  255 - 0xff
    "11111111", -- 2963 - 0xb93  :  255 - 0xff
    "11111111", -- 2964 - 0xb94  :  255 - 0xff
    "11111111", -- 2965 - 0xb95  :  255 - 0xff
    "11111111", -- 2966 - 0xb96  :  255 - 0xff
    "11111111", -- 2967 - 0xb97  :  255 - 0xff
    "11111111", -- 2968 - 0xb98  :  255 - 0xff -- Background 0x73
    "11111111", -- 2969 - 0xb99  :  255 - 0xff
    "11111111", -- 2970 - 0xb9a  :  255 - 0xff
    "11111111", -- 2971 - 0xb9b  :  255 - 0xff
    "11111111", -- 2972 - 0xb9c  :  255 - 0xff
    "11111111", -- 2973 - 0xb9d  :  255 - 0xff
    "11111111", -- 2974 - 0xb9e  :  255 - 0xff
    "11111111", -- 2975 - 0xb9f  :  255 - 0xff
    "11111111", -- 2976 - 0xba0  :  255 - 0xff -- Background 0x74
    "11111111", -- 2977 - 0xba1  :  255 - 0xff
    "11111111", -- 2978 - 0xba2  :  255 - 0xff
    "11111111", -- 2979 - 0xba3  :  255 - 0xff
    "11111111", -- 2980 - 0xba4  :  255 - 0xff
    "11111111", -- 2981 - 0xba5  :  255 - 0xff
    "11111111", -- 2982 - 0xba6  :  255 - 0xff
    "11111111", -- 2983 - 0xba7  :  255 - 0xff
    "11111111", -- 2984 - 0xba8  :  255 - 0xff -- Background 0x75
    "11111111", -- 2985 - 0xba9  :  255 - 0xff
    "11111111", -- 2986 - 0xbaa  :  255 - 0xff
    "11111111", -- 2987 - 0xbab  :  255 - 0xff
    "11111111", -- 2988 - 0xbac  :  255 - 0xff
    "11111111", -- 2989 - 0xbad  :  255 - 0xff
    "11111111", -- 2990 - 0xbae  :  255 - 0xff
    "11111111", -- 2991 - 0xbaf  :  255 - 0xff
    "11111111", -- 2992 - 0xbb0  :  255 - 0xff -- Background 0x76
    "11111111", -- 2993 - 0xbb1  :  255 - 0xff
    "11111111", -- 2994 - 0xbb2  :  255 - 0xff
    "11111111", -- 2995 - 0xbb3  :  255 - 0xff
    "11111111", -- 2996 - 0xbb4  :  255 - 0xff
    "11111111", -- 2997 - 0xbb5  :  255 - 0xff
    "11111111", -- 2998 - 0xbb6  :  255 - 0xff
    "11111111", -- 2999 - 0xbb7  :  255 - 0xff
    "11111111", -- 3000 - 0xbb8  :  255 - 0xff -- Background 0x77
    "11111111", -- 3001 - 0xbb9  :  255 - 0xff
    "11111111", -- 3002 - 0xbba  :  255 - 0xff
    "11111111", -- 3003 - 0xbbb  :  255 - 0xff
    "11111111", -- 3004 - 0xbbc  :  255 - 0xff
    "11111111", -- 3005 - 0xbbd  :  255 - 0xff
    "11111111", -- 3006 - 0xbbe  :  255 - 0xff
    "11111111", -- 3007 - 0xbbf  :  255 - 0xff
    "11111111", -- 3008 - 0xbc0  :  255 - 0xff -- Background 0x78
    "11111111", -- 3009 - 0xbc1  :  255 - 0xff
    "11111111", -- 3010 - 0xbc2  :  255 - 0xff
    "11111111", -- 3011 - 0xbc3  :  255 - 0xff
    "11111111", -- 3012 - 0xbc4  :  255 - 0xff
    "11111111", -- 3013 - 0xbc5  :  255 - 0xff
    "11111111", -- 3014 - 0xbc6  :  255 - 0xff
    "11111111", -- 3015 - 0xbc7  :  255 - 0xff
    "11111111", -- 3016 - 0xbc8  :  255 - 0xff -- Background 0x79
    "11111111", -- 3017 - 0xbc9  :  255 - 0xff
    "11111111", -- 3018 - 0xbca  :  255 - 0xff
    "11111111", -- 3019 - 0xbcb  :  255 - 0xff
    "11111111", -- 3020 - 0xbcc  :  255 - 0xff
    "11111111", -- 3021 - 0xbcd  :  255 - 0xff
    "11111111", -- 3022 - 0xbce  :  255 - 0xff
    "11111111", -- 3023 - 0xbcf  :  255 - 0xff
    "11111111", -- 3024 - 0xbd0  :  255 - 0xff -- Background 0x7a
    "11111111", -- 3025 - 0xbd1  :  255 - 0xff
    "11111111", -- 3026 - 0xbd2  :  255 - 0xff
    "11111111", -- 3027 - 0xbd3  :  255 - 0xff
    "11111111", -- 3028 - 0xbd4  :  255 - 0xff
    "11111111", -- 3029 - 0xbd5  :  255 - 0xff
    "11111111", -- 3030 - 0xbd6  :  255 - 0xff
    "11111111", -- 3031 - 0xbd7  :  255 - 0xff
    "11111111", -- 3032 - 0xbd8  :  255 - 0xff -- Background 0x7b
    "11111111", -- 3033 - 0xbd9  :  255 - 0xff
    "11111111", -- 3034 - 0xbda  :  255 - 0xff
    "11111111", -- 3035 - 0xbdb  :  255 - 0xff
    "11111111", -- 3036 - 0xbdc  :  255 - 0xff
    "11111111", -- 3037 - 0xbdd  :  255 - 0xff
    "11111111", -- 3038 - 0xbde  :  255 - 0xff
    "11111111", -- 3039 - 0xbdf  :  255 - 0xff
    "11111111", -- 3040 - 0xbe0  :  255 - 0xff -- Background 0x7c
    "11111111", -- 3041 - 0xbe1  :  255 - 0xff
    "11111111", -- 3042 - 0xbe2  :  255 - 0xff
    "11111111", -- 3043 - 0xbe3  :  255 - 0xff
    "11111111", -- 3044 - 0xbe4  :  255 - 0xff
    "11111111", -- 3045 - 0xbe5  :  255 - 0xff
    "11111111", -- 3046 - 0xbe6  :  255 - 0xff
    "11111111", -- 3047 - 0xbe7  :  255 - 0xff
    "11111111", -- 3048 - 0xbe8  :  255 - 0xff -- Background 0x7d
    "11111111", -- 3049 - 0xbe9  :  255 - 0xff
    "11111111", -- 3050 - 0xbea  :  255 - 0xff
    "11111111", -- 3051 - 0xbeb  :  255 - 0xff
    "11111111", -- 3052 - 0xbec  :  255 - 0xff
    "11111111", -- 3053 - 0xbed  :  255 - 0xff
    "11111111", -- 3054 - 0xbee  :  255 - 0xff
    "11111111", -- 3055 - 0xbef  :  255 - 0xff
    "11111111", -- 3056 - 0xbf0  :  255 - 0xff -- Background 0x7e
    "11111111", -- 3057 - 0xbf1  :  255 - 0xff
    "11111111", -- 3058 - 0xbf2  :  255 - 0xff
    "11111111", -- 3059 - 0xbf3  :  255 - 0xff
    "11111111", -- 3060 - 0xbf4  :  255 - 0xff
    "11111111", -- 3061 - 0xbf5  :  255 - 0xff
    "11111111", -- 3062 - 0xbf6  :  255 - 0xff
    "11111111", -- 3063 - 0xbf7  :  255 - 0xff
    "11111111", -- 3064 - 0xbf8  :  255 - 0xff -- Background 0x7f
    "11111111", -- 3065 - 0xbf9  :  255 - 0xff
    "11111111", -- 3066 - 0xbfa  :  255 - 0xff
    "11111111", -- 3067 - 0xbfb  :  255 - 0xff
    "11111111", -- 3068 - 0xbfc  :  255 - 0xff
    "11111111", -- 3069 - 0xbfd  :  255 - 0xff
    "11111111", -- 3070 - 0xbfe  :  255 - 0xff
    "11111111", -- 3071 - 0xbff  :  255 - 0xff
    "11111111", -- 3072 - 0xc00  :  255 - 0xff -- Background 0x80
    "11111111", -- 3073 - 0xc01  :  255 - 0xff
    "11111111", -- 3074 - 0xc02  :  255 - 0xff
    "11111111", -- 3075 - 0xc03  :  255 - 0xff
    "11111111", -- 3076 - 0xc04  :  255 - 0xff
    "11111111", -- 3077 - 0xc05  :  255 - 0xff
    "11111111", -- 3078 - 0xc06  :  255 - 0xff
    "11111111", -- 3079 - 0xc07  :  255 - 0xff
    "11111111", -- 3080 - 0xc08  :  255 - 0xff -- Background 0x81
    "11111111", -- 3081 - 0xc09  :  255 - 0xff
    "11111111", -- 3082 - 0xc0a  :  255 - 0xff
    "11111111", -- 3083 - 0xc0b  :  255 - 0xff
    "11111111", -- 3084 - 0xc0c  :  255 - 0xff
    "11111111", -- 3085 - 0xc0d  :  255 - 0xff
    "11111111", -- 3086 - 0xc0e  :  255 - 0xff
    "11111111", -- 3087 - 0xc0f  :  255 - 0xff
    "11111111", -- 3088 - 0xc10  :  255 - 0xff -- Background 0x82
    "11111111", -- 3089 - 0xc11  :  255 - 0xff
    "11111111", -- 3090 - 0xc12  :  255 - 0xff
    "11111111", -- 3091 - 0xc13  :  255 - 0xff
    "11111111", -- 3092 - 0xc14  :  255 - 0xff
    "11111111", -- 3093 - 0xc15  :  255 - 0xff
    "11111111", -- 3094 - 0xc16  :  255 - 0xff
    "11111111", -- 3095 - 0xc17  :  255 - 0xff
    "11111111", -- 3096 - 0xc18  :  255 - 0xff -- Background 0x83
    "11111111", -- 3097 - 0xc19  :  255 - 0xff
    "11111111", -- 3098 - 0xc1a  :  255 - 0xff
    "11111111", -- 3099 - 0xc1b  :  255 - 0xff
    "11111111", -- 3100 - 0xc1c  :  255 - 0xff
    "11111111", -- 3101 - 0xc1d  :  255 - 0xff
    "11111111", -- 3102 - 0xc1e  :  255 - 0xff
    "11111111", -- 3103 - 0xc1f  :  255 - 0xff
    "11111111", -- 3104 - 0xc20  :  255 - 0xff -- Background 0x84
    "11111111", -- 3105 - 0xc21  :  255 - 0xff
    "11111111", -- 3106 - 0xc22  :  255 - 0xff
    "11111111", -- 3107 - 0xc23  :  255 - 0xff
    "11111111", -- 3108 - 0xc24  :  255 - 0xff
    "11111111", -- 3109 - 0xc25  :  255 - 0xff
    "11111111", -- 3110 - 0xc26  :  255 - 0xff
    "11111111", -- 3111 - 0xc27  :  255 - 0xff
    "11111111", -- 3112 - 0xc28  :  255 - 0xff -- Background 0x85
    "11111111", -- 3113 - 0xc29  :  255 - 0xff
    "11111111", -- 3114 - 0xc2a  :  255 - 0xff
    "11111111", -- 3115 - 0xc2b  :  255 - 0xff
    "11111111", -- 3116 - 0xc2c  :  255 - 0xff
    "11111111", -- 3117 - 0xc2d  :  255 - 0xff
    "11111111", -- 3118 - 0xc2e  :  255 - 0xff
    "11111111", -- 3119 - 0xc2f  :  255 - 0xff
    "11111111", -- 3120 - 0xc30  :  255 - 0xff -- Background 0x86
    "11111111", -- 3121 - 0xc31  :  255 - 0xff
    "11111111", -- 3122 - 0xc32  :  255 - 0xff
    "11111111", -- 3123 - 0xc33  :  255 - 0xff
    "11111111", -- 3124 - 0xc34  :  255 - 0xff
    "11111111", -- 3125 - 0xc35  :  255 - 0xff
    "11111111", -- 3126 - 0xc36  :  255 - 0xff
    "11111111", -- 3127 - 0xc37  :  255 - 0xff
    "11111111", -- 3128 - 0xc38  :  255 - 0xff -- Background 0x87
    "11111111", -- 3129 - 0xc39  :  255 - 0xff
    "11111111", -- 3130 - 0xc3a  :  255 - 0xff
    "11111111", -- 3131 - 0xc3b  :  255 - 0xff
    "11111111", -- 3132 - 0xc3c  :  255 - 0xff
    "11111111", -- 3133 - 0xc3d  :  255 - 0xff
    "11111111", -- 3134 - 0xc3e  :  255 - 0xff
    "11111111", -- 3135 - 0xc3f  :  255 - 0xff
    "11111111", -- 3136 - 0xc40  :  255 - 0xff -- Background 0x88
    "11111111", -- 3137 - 0xc41  :  255 - 0xff
    "11111111", -- 3138 - 0xc42  :  255 - 0xff
    "11111111", -- 3139 - 0xc43  :  255 - 0xff
    "11111111", -- 3140 - 0xc44  :  255 - 0xff
    "11111111", -- 3141 - 0xc45  :  255 - 0xff
    "11111111", -- 3142 - 0xc46  :  255 - 0xff
    "11111111", -- 3143 - 0xc47  :  255 - 0xff
    "11111111", -- 3144 - 0xc48  :  255 - 0xff -- Background 0x89
    "11111111", -- 3145 - 0xc49  :  255 - 0xff
    "11111111", -- 3146 - 0xc4a  :  255 - 0xff
    "11111111", -- 3147 - 0xc4b  :  255 - 0xff
    "11111111", -- 3148 - 0xc4c  :  255 - 0xff
    "11111111", -- 3149 - 0xc4d  :  255 - 0xff
    "11111111", -- 3150 - 0xc4e  :  255 - 0xff
    "11111111", -- 3151 - 0xc4f  :  255 - 0xff
    "11111111", -- 3152 - 0xc50  :  255 - 0xff -- Background 0x8a
    "11111111", -- 3153 - 0xc51  :  255 - 0xff
    "11111111", -- 3154 - 0xc52  :  255 - 0xff
    "11111111", -- 3155 - 0xc53  :  255 - 0xff
    "11111111", -- 3156 - 0xc54  :  255 - 0xff
    "11111111", -- 3157 - 0xc55  :  255 - 0xff
    "11111111", -- 3158 - 0xc56  :  255 - 0xff
    "11111111", -- 3159 - 0xc57  :  255 - 0xff
    "11111111", -- 3160 - 0xc58  :  255 - 0xff -- Background 0x8b
    "11111111", -- 3161 - 0xc59  :  255 - 0xff
    "11111111", -- 3162 - 0xc5a  :  255 - 0xff
    "11111111", -- 3163 - 0xc5b  :  255 - 0xff
    "11111111", -- 3164 - 0xc5c  :  255 - 0xff
    "11111111", -- 3165 - 0xc5d  :  255 - 0xff
    "11111111", -- 3166 - 0xc5e  :  255 - 0xff
    "11111111", -- 3167 - 0xc5f  :  255 - 0xff
    "11111111", -- 3168 - 0xc60  :  255 - 0xff -- Background 0x8c
    "11111111", -- 3169 - 0xc61  :  255 - 0xff
    "11111111", -- 3170 - 0xc62  :  255 - 0xff
    "11111111", -- 3171 - 0xc63  :  255 - 0xff
    "11111111", -- 3172 - 0xc64  :  255 - 0xff
    "11111111", -- 3173 - 0xc65  :  255 - 0xff
    "11111111", -- 3174 - 0xc66  :  255 - 0xff
    "11111111", -- 3175 - 0xc67  :  255 - 0xff
    "11111111", -- 3176 - 0xc68  :  255 - 0xff -- Background 0x8d
    "11111111", -- 3177 - 0xc69  :  255 - 0xff
    "11111111", -- 3178 - 0xc6a  :  255 - 0xff
    "11111111", -- 3179 - 0xc6b  :  255 - 0xff
    "11111111", -- 3180 - 0xc6c  :  255 - 0xff
    "11111111", -- 3181 - 0xc6d  :  255 - 0xff
    "11111111", -- 3182 - 0xc6e  :  255 - 0xff
    "11111111", -- 3183 - 0xc6f  :  255 - 0xff
    "11111111", -- 3184 - 0xc70  :  255 - 0xff -- Background 0x8e
    "11111111", -- 3185 - 0xc71  :  255 - 0xff
    "11111111", -- 3186 - 0xc72  :  255 - 0xff
    "11111111", -- 3187 - 0xc73  :  255 - 0xff
    "11111111", -- 3188 - 0xc74  :  255 - 0xff
    "11111111", -- 3189 - 0xc75  :  255 - 0xff
    "11111111", -- 3190 - 0xc76  :  255 - 0xff
    "11111111", -- 3191 - 0xc77  :  255 - 0xff
    "11111111", -- 3192 - 0xc78  :  255 - 0xff -- Background 0x8f
    "11111111", -- 3193 - 0xc79  :  255 - 0xff
    "11111111", -- 3194 - 0xc7a  :  255 - 0xff
    "11111111", -- 3195 - 0xc7b  :  255 - 0xff
    "11111111", -- 3196 - 0xc7c  :  255 - 0xff
    "11111111", -- 3197 - 0xc7d  :  255 - 0xff
    "11111111", -- 3198 - 0xc7e  :  255 - 0xff
    "11111111", -- 3199 - 0xc7f  :  255 - 0xff
    "00000000", -- 3200 - 0xc80  :    0 - 0x0 -- Background 0x90
    "00000000", -- 3201 - 0xc81  :    0 - 0x0
    "00000000", -- 3202 - 0xc82  :    0 - 0x0
    "00000000", -- 3203 - 0xc83  :    0 - 0x0
    "00000000", -- 3204 - 0xc84  :    0 - 0x0
    "00000001", -- 3205 - 0xc85  :    1 - 0x1
    "00011110", -- 3206 - 0xc86  :   30 - 0x1e
    "00111011", -- 3207 - 0xc87  :   59 - 0x3b
    "00000000", -- 3208 - 0xc88  :    0 - 0x0 -- Background 0x91
    "00000000", -- 3209 - 0xc89  :    0 - 0x0
    "00001100", -- 3210 - 0xc8a  :   12 - 0xc
    "00111100", -- 3211 - 0xc8b  :   60 - 0x3c
    "11010000", -- 3212 - 0xc8c  :  208 - 0xd0
    "00010000", -- 3213 - 0xc8d  :   16 - 0x10
    "00100000", -- 3214 - 0xc8e  :   32 - 0x20
    "01000000", -- 3215 - 0xc8f  :   64 - 0x40
    "00111110", -- 3216 - 0xc90  :   62 - 0x3e -- Background 0x92
    "00101101", -- 3217 - 0xc91  :   45 - 0x2d
    "00110101", -- 3218 - 0xc92  :   53 - 0x35
    "00011101", -- 3219 - 0xc93  :   29 - 0x1d
    "00000001", -- 3220 - 0xc94  :    1 - 0x1
    "00000000", -- 3221 - 0xc95  :    0 - 0x0
    "00000000", -- 3222 - 0xc96  :    0 - 0x0
    "00000000", -- 3223 - 0xc97  :    0 - 0x0
    "10110000", -- 3224 - 0xc98  :  176 - 0xb0 -- Background 0x93
    "10111000", -- 3225 - 0xc99  :  184 - 0xb8
    "11111000", -- 3226 - 0xc9a  :  248 - 0xf8
    "01111000", -- 3227 - 0xc9b  :  120 - 0x78
    "10011000", -- 3228 - 0xc9c  :  152 - 0x98
    "11110000", -- 3229 - 0xc9d  :  240 - 0xf0
    "00000000", -- 3230 - 0xc9e  :    0 - 0x0
    "00000000", -- 3231 - 0xc9f  :    0 - 0x0
    "00000000", -- 3232 - 0xca0  :    0 - 0x0 -- Background 0x94
    "00000000", -- 3233 - 0xca1  :    0 - 0x0
    "00000111", -- 3234 - 0xca2  :    7 - 0x7
    "00000011", -- 3235 - 0xca3  :    3 - 0x3
    "00001101", -- 3236 - 0xca4  :   13 - 0xd
    "00011110", -- 3237 - 0xca5  :   30 - 0x1e
    "00010111", -- 3238 - 0xca6  :   23 - 0x17
    "00011101", -- 3239 - 0xca7  :   29 - 0x1d
    "00000000", -- 3240 - 0xca8  :    0 - 0x0 -- Background 0x95
    "10000000", -- 3241 - 0xca9  :  128 - 0x80
    "01110000", -- 3242 - 0xcaa  :  112 - 0x70
    "11100000", -- 3243 - 0xcab  :  224 - 0xe0
    "11011000", -- 3244 - 0xcac  :  216 - 0xd8
    "10111100", -- 3245 - 0xcad  :  188 - 0xbc
    "01110100", -- 3246 - 0xcae  :  116 - 0x74
    "11011100", -- 3247 - 0xcaf  :  220 - 0xdc
    "00011111", -- 3248 - 0xcb0  :   31 - 0x1f -- Background 0x96
    "00001011", -- 3249 - 0xcb1  :   11 - 0xb
    "00001111", -- 3250 - 0xcb2  :   15 - 0xf
    "00000101", -- 3251 - 0xcb3  :    5 - 0x5
    "00000011", -- 3252 - 0xcb4  :    3 - 0x3
    "00000001", -- 3253 - 0xcb5  :    1 - 0x1
    "00000000", -- 3254 - 0xcb6  :    0 - 0x0
    "00000000", -- 3255 - 0xcb7  :    0 - 0x0
    "11111100", -- 3256 - 0xcb8  :  252 - 0xfc -- Background 0x97
    "01101000", -- 3257 - 0xcb9  :  104 - 0x68
    "11111000", -- 3258 - 0xcba  :  248 - 0xf8
    "10110000", -- 3259 - 0xcbb  :  176 - 0xb0
    "11100000", -- 3260 - 0xcbc  :  224 - 0xe0
    "10000000", -- 3261 - 0xcbd  :  128 - 0x80
    "00000000", -- 3262 - 0xcbe  :    0 - 0x0
    "00000000", -- 3263 - 0xcbf  :    0 - 0x0
    "00000000", -- 3264 - 0xcc0  :    0 - 0x0 -- Background 0x98
    "00000000", -- 3265 - 0xcc1  :    0 - 0x0
    "00000000", -- 3266 - 0xcc2  :    0 - 0x0
    "00000001", -- 3267 - 0xcc3  :    1 - 0x1
    "00000001", -- 3268 - 0xcc4  :    1 - 0x1
    "00001011", -- 3269 - 0xcc5  :   11 - 0xb
    "00011100", -- 3270 - 0xcc6  :   28 - 0x1c
    "00111111", -- 3271 - 0xcc7  :   63 - 0x3f
    "00000000", -- 3272 - 0xcc8  :    0 - 0x0 -- Background 0x99
    "00000000", -- 3273 - 0xcc9  :    0 - 0x0
    "00110000", -- 3274 - 0xcca  :   48 - 0x30
    "01111000", -- 3275 - 0xccb  :  120 - 0x78
    "10000000", -- 3276 - 0xccc  :  128 - 0x80
    "11110000", -- 3277 - 0xccd  :  240 - 0xf0
    "11111000", -- 3278 - 0xcce  :  248 - 0xf8
    "11111100", -- 3279 - 0xccf  :  252 - 0xfc
    "00111111", -- 3280 - 0xcd0  :   63 - 0x3f -- Background 0x9a
    "00111111", -- 3281 - 0xcd1  :   63 - 0x3f
    "00111111", -- 3282 - 0xcd2  :   63 - 0x3f
    "00011111", -- 3283 - 0xcd3  :   31 - 0x1f
    "00011111", -- 3284 - 0xcd4  :   31 - 0x1f
    "00000111", -- 3285 - 0xcd5  :    7 - 0x7
    "00000000", -- 3286 - 0xcd6  :    0 - 0x0
    "00000000", -- 3287 - 0xcd7  :    0 - 0x0
    "11111100", -- 3288 - 0xcd8  :  252 - 0xfc -- Background 0x9b
    "11101100", -- 3289 - 0xcd9  :  236 - 0xec
    "11101100", -- 3290 - 0xcda  :  236 - 0xec
    "11011000", -- 3291 - 0xcdb  :  216 - 0xd8
    "11111000", -- 3292 - 0xcdc  :  248 - 0xf8
    "11100000", -- 3293 - 0xcdd  :  224 - 0xe0
    "00000000", -- 3294 - 0xcde  :    0 - 0x0
    "00000000", -- 3295 - 0xcdf  :    0 - 0x0
    "00000000", -- 3296 - 0xce0  :    0 - 0x0 -- Background 0x9c
    "00000000", -- 3297 - 0xce1  :    0 - 0x0
    "00000001", -- 3298 - 0xce2  :    1 - 0x1
    "00011101", -- 3299 - 0xce3  :   29 - 0x1d
    "00111110", -- 3300 - 0xce4  :   62 - 0x3e
    "00111111", -- 3301 - 0xce5  :   63 - 0x3f
    "00111111", -- 3302 - 0xce6  :   63 - 0x3f
    "00111111", -- 3303 - 0xce7  :   63 - 0x3f
    "00000000", -- 3304 - 0xce8  :    0 - 0x0 -- Background 0x9d
    "10000000", -- 3305 - 0xce9  :  128 - 0x80
    "00000000", -- 3306 - 0xcea  :    0 - 0x0
    "01110000", -- 3307 - 0xceb  :  112 - 0x70
    "11111000", -- 3308 - 0xcec  :  248 - 0xf8
    "11111100", -- 3309 - 0xced  :  252 - 0xfc
    "11111100", -- 3310 - 0xcee  :  252 - 0xfc
    "11111100", -- 3311 - 0xcef  :  252 - 0xfc
    "00111111", -- 3312 - 0xcf0  :   63 - 0x3f -- Background 0x9e
    "00111111", -- 3313 - 0xcf1  :   63 - 0x3f
    "00011111", -- 3314 - 0xcf2  :   31 - 0x1f
    "00011111", -- 3315 - 0xcf3  :   31 - 0x1f
    "00001111", -- 3316 - 0xcf4  :   15 - 0xf
    "00000110", -- 3317 - 0xcf5  :    6 - 0x6
    "00000000", -- 3318 - 0xcf6  :    0 - 0x0
    "00000000", -- 3319 - 0xcf7  :    0 - 0x0
    "11101100", -- 3320 - 0xcf8  :  236 - 0xec -- Background 0x9f
    "11101100", -- 3321 - 0xcf9  :  236 - 0xec
    "11011000", -- 3322 - 0xcfa  :  216 - 0xd8
    "11111000", -- 3323 - 0xcfb  :  248 - 0xf8
    "11110000", -- 3324 - 0xcfc  :  240 - 0xf0
    "11100000", -- 3325 - 0xcfd  :  224 - 0xe0
    "00000000", -- 3326 - 0xcfe  :    0 - 0x0
    "00000000", -- 3327 - 0xcff  :    0 - 0x0
    "00000000", -- 3328 - 0xd00  :    0 - 0x0 -- Background 0xa0
    "00000100", -- 3329 - 0xd01  :    4 - 0x4
    "00000011", -- 3330 - 0xd02  :    3 - 0x3
    "00000000", -- 3331 - 0xd03  :    0 - 0x0
    "00000001", -- 3332 - 0xd04  :    1 - 0x1
    "00000111", -- 3333 - 0xd05  :    7 - 0x7
    "00001111", -- 3334 - 0xd06  :   15 - 0xf
    "00001100", -- 3335 - 0xd07  :   12 - 0xc
    "00000000", -- 3336 - 0xd08  :    0 - 0x0 -- Background 0xa1
    "00000000", -- 3337 - 0xd09  :    0 - 0x0
    "11100000", -- 3338 - 0xd0a  :  224 - 0xe0
    "10000000", -- 3339 - 0xd0b  :  128 - 0x80
    "01000000", -- 3340 - 0xd0c  :   64 - 0x40
    "11110000", -- 3341 - 0xd0d  :  240 - 0xf0
    "10011000", -- 3342 - 0xd0e  :  152 - 0x98
    "11111000", -- 3343 - 0xd0f  :  248 - 0xf8
    "00011111", -- 3344 - 0xd10  :   31 - 0x1f -- Background 0xa2
    "00010011", -- 3345 - 0xd11  :   19 - 0x13
    "00011111", -- 3346 - 0xd12  :   31 - 0x1f
    "00001111", -- 3347 - 0xd13  :   15 - 0xf
    "00001001", -- 3348 - 0xd14  :    9 - 0x9
    "00000111", -- 3349 - 0xd15  :    7 - 0x7
    "00000001", -- 3350 - 0xd16  :    1 - 0x1
    "00000000", -- 3351 - 0xd17  :    0 - 0x0
    "11100100", -- 3352 - 0xd18  :  228 - 0xe4 -- Background 0xa3
    "00111100", -- 3353 - 0xd19  :   60 - 0x3c
    "11100100", -- 3354 - 0xd1a  :  228 - 0xe4
    "00111000", -- 3355 - 0xd1b  :   56 - 0x38
    "11111000", -- 3356 - 0xd1c  :  248 - 0xf8
    "11110000", -- 3357 - 0xd1d  :  240 - 0xf0
    "11000000", -- 3358 - 0xd1e  :  192 - 0xc0
    "00000000", -- 3359 - 0xd1f  :    0 - 0x0
    "00000000", -- 3360 - 0xd20  :    0 - 0x0 -- Background 0xa4
    "00000000", -- 3361 - 0xd21  :    0 - 0x0
    "00000000", -- 3362 - 0xd22  :    0 - 0x0
    "00000000", -- 3363 - 0xd23  :    0 - 0x0
    "00010001", -- 3364 - 0xd24  :   17 - 0x11
    "00010011", -- 3365 - 0xd25  :   19 - 0x13
    "00011111", -- 3366 - 0xd26  :   31 - 0x1f
    "00011111", -- 3367 - 0xd27  :   31 - 0x1f
    "00000000", -- 3368 - 0xd28  :    0 - 0x0 -- Background 0xa5
    "00000000", -- 3369 - 0xd29  :    0 - 0x0
    "00000000", -- 3370 - 0xd2a  :    0 - 0x0
    "10000000", -- 3371 - 0xd2b  :  128 - 0x80
    "11000100", -- 3372 - 0xd2c  :  196 - 0xc4
    "11100100", -- 3373 - 0xd2d  :  228 - 0xe4
    "11111100", -- 3374 - 0xd2e  :  252 - 0xfc
    "11111100", -- 3375 - 0xd2f  :  252 - 0xfc
    "00011111", -- 3376 - 0xd30  :   31 - 0x1f -- Background 0xa6
    "00001110", -- 3377 - 0xd31  :   14 - 0xe
    "00000110", -- 3378 - 0xd32  :    6 - 0x6
    "00000010", -- 3379 - 0xd33  :    2 - 0x2
    "00000000", -- 3380 - 0xd34  :    0 - 0x0
    "00000000", -- 3381 - 0xd35  :    0 - 0x0
    "00000000", -- 3382 - 0xd36  :    0 - 0x0
    "00000000", -- 3383 - 0xd37  :    0 - 0x0
    "11111100", -- 3384 - 0xd38  :  252 - 0xfc -- Background 0xa7
    "10111000", -- 3385 - 0xd39  :  184 - 0xb8
    "10110000", -- 3386 - 0xd3a  :  176 - 0xb0
    "10100000", -- 3387 - 0xd3b  :  160 - 0xa0
    "10000000", -- 3388 - 0xd3c  :  128 - 0x80
    "00000000", -- 3389 - 0xd3d  :    0 - 0x0
    "00000000", -- 3390 - 0xd3e  :    0 - 0x0
    "00000000", -- 3391 - 0xd3f  :    0 - 0x0
    "00000000", -- 3392 - 0xd40  :    0 - 0x0 -- Background 0xa8
    "00000000", -- 3393 - 0xd41  :    0 - 0x0
    "00000000", -- 3394 - 0xd42  :    0 - 0x0
    "00000001", -- 3395 - 0xd43  :    1 - 0x1
    "00000011", -- 3396 - 0xd44  :    3 - 0x3
    "00000110", -- 3397 - 0xd45  :    6 - 0x6
    "00000110", -- 3398 - 0xd46  :    6 - 0x6
    "00001111", -- 3399 - 0xd47  :   15 - 0xf
    "00000000", -- 3400 - 0xd48  :    0 - 0x0 -- Background 0xa9
    "00011000", -- 3401 - 0xd49  :   24 - 0x18
    "11110100", -- 3402 - 0xd4a  :  244 - 0xf4
    "11111000", -- 3403 - 0xd4b  :  248 - 0xf8
    "00111000", -- 3404 - 0xd4c  :   56 - 0x38
    "01111100", -- 3405 - 0xd4d  :  124 - 0x7c
    "11111100", -- 3406 - 0xd4e  :  252 - 0xfc
    "11111100", -- 3407 - 0xd4f  :  252 - 0xfc
    "00001111", -- 3408 - 0xd50  :   15 - 0xf -- Background 0xaa
    "00011111", -- 3409 - 0xd51  :   31 - 0x1f
    "00110000", -- 3410 - 0xd52  :   48 - 0x30
    "00111000", -- 3411 - 0xd53  :   56 - 0x38
    "00011101", -- 3412 - 0xd54  :   29 - 0x1d
    "00000011", -- 3413 - 0xd55  :    3 - 0x3
    "00000011", -- 3414 - 0xd56  :    3 - 0x3
    "00000000", -- 3415 - 0xd57  :    0 - 0x0
    "11111100", -- 3416 - 0xd58  :  252 - 0xfc -- Background 0xab
    "11111100", -- 3417 - 0xd59  :  252 - 0xfc
    "01111100", -- 3418 - 0xd5a  :  124 - 0x7c
    "10001110", -- 3419 - 0xd5b  :  142 - 0x8e
    "10000110", -- 3420 - 0xd5c  :  134 - 0x86
    "10011100", -- 3421 - 0xd5d  :  156 - 0x9c
    "01111000", -- 3422 - 0xd5e  :  120 - 0x78
    "00000000", -- 3423 - 0xd5f  :    0 - 0x0
    "00000000", -- 3424 - 0xd60  :    0 - 0x0 -- Background 0xac
    "00000001", -- 3425 - 0xd61  :    1 - 0x1
    "00000110", -- 3426 - 0xd62  :    6 - 0x6
    "00000111", -- 3427 - 0xd63  :    7 - 0x7
    "00000111", -- 3428 - 0xd64  :    7 - 0x7
    "00000111", -- 3429 - 0xd65  :    7 - 0x7
    "00000001", -- 3430 - 0xd66  :    1 - 0x1
    "00000011", -- 3431 - 0xd67  :    3 - 0x3
    "00000000", -- 3432 - 0xd68  :    0 - 0x0 -- Background 0xad
    "11000000", -- 3433 - 0xd69  :  192 - 0xc0
    "00110000", -- 3434 - 0xd6a  :   48 - 0x30
    "11110000", -- 3435 - 0xd6b  :  240 - 0xf0
    "11110000", -- 3436 - 0xd6c  :  240 - 0xf0
    "11110000", -- 3437 - 0xd6d  :  240 - 0xf0
    "01000000", -- 3438 - 0xd6e  :   64 - 0x40
    "01000000", -- 3439 - 0xd6f  :   64 - 0x40
    "00000001", -- 3440 - 0xd70  :    1 - 0x1 -- Background 0xae
    "00000000", -- 3441 - 0xd71  :    0 - 0x0
    "00000001", -- 3442 - 0xd72  :    1 - 0x1
    "00000011", -- 3443 - 0xd73  :    3 - 0x3
    "00000001", -- 3444 - 0xd74  :    1 - 0x1
    "00000000", -- 3445 - 0xd75  :    0 - 0x0
    "00000000", -- 3446 - 0xd76  :    0 - 0x0
    "00000000", -- 3447 - 0xd77  :    0 - 0x0
    "01000000", -- 3448 - 0xd78  :   64 - 0x40 -- Background 0xaf
    "01000000", -- 3449 - 0xd79  :   64 - 0x40
    "01000000", -- 3450 - 0xd7a  :   64 - 0x40
    "01000000", -- 3451 - 0xd7b  :   64 - 0x40
    "01000000", -- 3452 - 0xd7c  :   64 - 0x40
    "10000000", -- 3453 - 0xd7d  :  128 - 0x80
    "00000000", -- 3454 - 0xd7e  :    0 - 0x0
    "00000000", -- 3455 - 0xd7f  :    0 - 0x0
    "01111110", -- 3456 - 0xd80  :  126 - 0x7e -- Background 0xb0
    "01100011", -- 3457 - 0xd81  :   99 - 0x63
    "01100011", -- 3458 - 0xd82  :   99 - 0x63
    "01100011", -- 3459 - 0xd83  :   99 - 0x63
    "01111110", -- 3460 - 0xd84  :  126 - 0x7e
    "01100000", -- 3461 - 0xd85  :   96 - 0x60
    "01100000", -- 3462 - 0xd86  :   96 - 0x60
    "00000000", -- 3463 - 0xd87  :    0 - 0x0
    "01100000", -- 3464 - 0xd88  :   96 - 0x60 -- Background 0xb1
    "01100000", -- 3465 - 0xd89  :   96 - 0x60
    "01100000", -- 3466 - 0xd8a  :   96 - 0x60
    "01100000", -- 3467 - 0xd8b  :   96 - 0x60
    "01100000", -- 3468 - 0xd8c  :   96 - 0x60
    "01100000", -- 3469 - 0xd8d  :   96 - 0x60
    "01111111", -- 3470 - 0xd8e  :  127 - 0x7f
    "00000000", -- 3471 - 0xd8f  :    0 - 0x0
    "00011100", -- 3472 - 0xd90  :   28 - 0x1c -- Background 0xb2
    "00110110", -- 3473 - 0xd91  :   54 - 0x36
    "01100011", -- 3474 - 0xd92  :   99 - 0x63
    "01100011", -- 3475 - 0xd93  :   99 - 0x63
    "01111111", -- 3476 - 0xd94  :  127 - 0x7f
    "01100011", -- 3477 - 0xd95  :   99 - 0x63
    "01100011", -- 3478 - 0xd96  :   99 - 0x63
    "00000000", -- 3479 - 0xd97  :    0 - 0x0
    "00110011", -- 3480 - 0xd98  :   51 - 0x33 -- Background 0xb3
    "00110011", -- 3481 - 0xd99  :   51 - 0x33
    "00110011", -- 3482 - 0xd9a  :   51 - 0x33
    "00011110", -- 3483 - 0xd9b  :   30 - 0x1e
    "00001100", -- 3484 - 0xd9c  :   12 - 0xc
    "00001100", -- 3485 - 0xd9d  :   12 - 0xc
    "00001100", -- 3486 - 0xd9e  :   12 - 0xc
    "00000000", -- 3487 - 0xd9f  :    0 - 0x0
    "01111111", -- 3488 - 0xda0  :  127 - 0x7f -- Background 0xb4
    "01100000", -- 3489 - 0xda1  :   96 - 0x60
    "01100000", -- 3490 - 0xda2  :   96 - 0x60
    "01111110", -- 3491 - 0xda3  :  126 - 0x7e
    "01100000", -- 3492 - 0xda4  :   96 - 0x60
    "01100000", -- 3493 - 0xda5  :   96 - 0x60
    "01111111", -- 3494 - 0xda6  :  127 - 0x7f
    "00000000", -- 3495 - 0xda7  :    0 - 0x0
    "01111110", -- 3496 - 0xda8  :  126 - 0x7e -- Background 0xb5
    "01100011", -- 3497 - 0xda9  :   99 - 0x63
    "01100011", -- 3498 - 0xdaa  :   99 - 0x63
    "01100111", -- 3499 - 0xdab  :  103 - 0x67
    "01111100", -- 3500 - 0xdac  :  124 - 0x7c
    "01101110", -- 3501 - 0xdad  :  110 - 0x6e
    "01100111", -- 3502 - 0xdae  :  103 - 0x67
    "00000000", -- 3503 - 0xdaf  :    0 - 0x0
    "00111110", -- 3504 - 0xdb0  :   62 - 0x3e -- Background 0xb6
    "01100011", -- 3505 - 0xdb1  :   99 - 0x63
    "01100011", -- 3506 - 0xdb2  :   99 - 0x63
    "01100011", -- 3507 - 0xdb3  :   99 - 0x63
    "01100011", -- 3508 - 0xdb4  :   99 - 0x63
    "01100011", -- 3509 - 0xdb5  :   99 - 0x63
    "00111110", -- 3510 - 0xdb6  :   62 - 0x3e
    "00000000", -- 3511 - 0xdb7  :    0 - 0x0
    "01100011", -- 3512 - 0xdb8  :   99 - 0x63 -- Background 0xb7
    "01110011", -- 3513 - 0xdb9  :  115 - 0x73
    "01111011", -- 3514 - 0xdba  :  123 - 0x7b
    "01111111", -- 3515 - 0xdbb  :  127 - 0x7f
    "01101111", -- 3516 - 0xdbc  :  111 - 0x6f
    "01100111", -- 3517 - 0xdbd  :  103 - 0x67
    "01100011", -- 3518 - 0xdbe  :   99 - 0x63
    "00000000", -- 3519 - 0xdbf  :    0 - 0x0
    "00111111", -- 3520 - 0xdc0  :   63 - 0x3f -- Background 0xb8
    "00001100", -- 3521 - 0xdc1  :   12 - 0xc
    "00001100", -- 3522 - 0xdc2  :   12 - 0xc
    "00001100", -- 3523 - 0xdc3  :   12 - 0xc
    "00001100", -- 3524 - 0xdc4  :   12 - 0xc
    "00001100", -- 3525 - 0xdc5  :   12 - 0xc
    "00001100", -- 3526 - 0xdc6  :   12 - 0xc
    "00000000", -- 3527 - 0xdc7  :    0 - 0x0
    "01100011", -- 3528 - 0xdc8  :   99 - 0x63 -- Background 0xb9
    "01100011", -- 3529 - 0xdc9  :   99 - 0x63
    "01101011", -- 3530 - 0xdca  :  107 - 0x6b
    "01111111", -- 3531 - 0xdcb  :  127 - 0x7f
    "01111111", -- 3532 - 0xdcc  :  127 - 0x7f
    "01110111", -- 3533 - 0xdcd  :  119 - 0x77
    "01100011", -- 3534 - 0xdce  :   99 - 0x63
    "00000000", -- 3535 - 0xdcf  :    0 - 0x0
    "01111100", -- 3536 - 0xdd0  :  124 - 0x7c -- Background 0xba
    "01100110", -- 3537 - 0xdd1  :  102 - 0x66
    "01100011", -- 3538 - 0xdd2  :   99 - 0x63
    "01100011", -- 3539 - 0xdd3  :   99 - 0x63
    "01100011", -- 3540 - 0xdd4  :   99 - 0x63
    "01100110", -- 3541 - 0xdd5  :  102 - 0x66
    "01111100", -- 3542 - 0xdd6  :  124 - 0x7c
    "00000000", -- 3543 - 0xdd7  :    0 - 0x0
    "00011100", -- 3544 - 0xdd8  :   28 - 0x1c -- Background 0xbb
    "00011100", -- 3545 - 0xdd9  :   28 - 0x1c
    "00011100", -- 3546 - 0xdda  :   28 - 0x1c
    "00011000", -- 3547 - 0xddb  :   24 - 0x18
    "00011000", -- 3548 - 0xddc  :   24 - 0x18
    "00000000", -- 3549 - 0xddd  :    0 - 0x0
    "00011000", -- 3550 - 0xdde  :   24 - 0x18
    "00000000", -- 3551 - 0xddf  :    0 - 0x0
    "00011111", -- 3552 - 0xde0  :   31 - 0x1f -- Background 0xbc
    "00110000", -- 3553 - 0xde1  :   48 - 0x30
    "01100000", -- 3554 - 0xde2  :   96 - 0x60
    "01100111", -- 3555 - 0xde3  :  103 - 0x67
    "01100011", -- 3556 - 0xde4  :   99 - 0x63
    "00110011", -- 3557 - 0xde5  :   51 - 0x33
    "00011111", -- 3558 - 0xde6  :   31 - 0x1f
    "00000000", -- 3559 - 0xde7  :    0 - 0x0
    "01100011", -- 3560 - 0xde8  :   99 - 0x63 -- Background 0xbd
    "01110111", -- 3561 - 0xde9  :  119 - 0x77
    "01111111", -- 3562 - 0xdea  :  127 - 0x7f
    "01111111", -- 3563 - 0xdeb  :  127 - 0x7f
    "01101011", -- 3564 - 0xdec  :  107 - 0x6b
    "01100011", -- 3565 - 0xded  :   99 - 0x63
    "01100011", -- 3566 - 0xdee  :   99 - 0x63
    "00000000", -- 3567 - 0xdef  :    0 - 0x0
    "01100011", -- 3568 - 0xdf0  :   99 - 0x63 -- Background 0xbe
    "01100011", -- 3569 - 0xdf1  :   99 - 0x63
    "01100011", -- 3570 - 0xdf2  :   99 - 0x63
    "01110111", -- 3571 - 0xdf3  :  119 - 0x77
    "00111110", -- 3572 - 0xdf4  :   62 - 0x3e
    "00011100", -- 3573 - 0xdf5  :   28 - 0x1c
    "00001000", -- 3574 - 0xdf6  :    8 - 0x8
    "00000000", -- 3575 - 0xdf7  :    0 - 0x0
    "00000000", -- 3576 - 0xdf8  :    0 - 0x0 -- Background 0xbf
    "00000000", -- 3577 - 0xdf9  :    0 - 0x0
    "00000000", -- 3578 - 0xdfa  :    0 - 0x0
    "00000000", -- 3579 - 0xdfb  :    0 - 0x0
    "00000000", -- 3580 - 0xdfc  :    0 - 0x0
    "00000000", -- 3581 - 0xdfd  :    0 - 0x0
    "00000000", -- 3582 - 0xdfe  :    0 - 0x0
    "00000000", -- 3583 - 0xdff  :    0 - 0x0
    "00011111", -- 3584 - 0xe00  :   31 - 0x1f -- Background 0xc0
    "00110000", -- 3585 - 0xe01  :   48 - 0x30
    "01100000", -- 3586 - 0xe02  :   96 - 0x60
    "01100111", -- 3587 - 0xe03  :  103 - 0x67
    "01100011", -- 3588 - 0xe04  :   99 - 0x63
    "00110011", -- 3589 - 0xe05  :   51 - 0x33
    "00011111", -- 3590 - 0xe06  :   31 - 0x1f
    "00000000", -- 3591 - 0xe07  :    0 - 0x0
    "00011100", -- 3592 - 0xe08  :   28 - 0x1c -- Background 0xc1
    "00110110", -- 3593 - 0xe09  :   54 - 0x36
    "01100011", -- 3594 - 0xe0a  :   99 - 0x63
    "01100011", -- 3595 - 0xe0b  :   99 - 0x63
    "01111111", -- 3596 - 0xe0c  :  127 - 0x7f
    "01100011", -- 3597 - 0xe0d  :   99 - 0x63
    "01100011", -- 3598 - 0xe0e  :   99 - 0x63
    "00000000", -- 3599 - 0xe0f  :    0 - 0x0
    "01100011", -- 3600 - 0xe10  :   99 - 0x63 -- Background 0xc2
    "01110111", -- 3601 - 0xe11  :  119 - 0x77
    "01111111", -- 3602 - 0xe12  :  127 - 0x7f
    "01111111", -- 3603 - 0xe13  :  127 - 0x7f
    "01101011", -- 3604 - 0xe14  :  107 - 0x6b
    "01100011", -- 3605 - 0xe15  :   99 - 0x63
    "01100011", -- 3606 - 0xe16  :   99 - 0x63
    "00000000", -- 3607 - 0xe17  :    0 - 0x0
    "01111111", -- 3608 - 0xe18  :  127 - 0x7f -- Background 0xc3
    "01100000", -- 3609 - 0xe19  :   96 - 0x60
    "01100000", -- 3610 - 0xe1a  :   96 - 0x60
    "01111110", -- 3611 - 0xe1b  :  126 - 0x7e
    "01100000", -- 3612 - 0xe1c  :   96 - 0x60
    "01100000", -- 3613 - 0xe1d  :   96 - 0x60
    "01111111", -- 3614 - 0xe1e  :  127 - 0x7f
    "00000000", -- 3615 - 0xe1f  :    0 - 0x0
    "00111110", -- 3616 - 0xe20  :   62 - 0x3e -- Background 0xc4
    "01100011", -- 3617 - 0xe21  :   99 - 0x63
    "01100011", -- 3618 - 0xe22  :   99 - 0x63
    "01100011", -- 3619 - 0xe23  :   99 - 0x63
    "01100011", -- 3620 - 0xe24  :   99 - 0x63
    "01100011", -- 3621 - 0xe25  :   99 - 0x63
    "00111110", -- 3622 - 0xe26  :   62 - 0x3e
    "00000000", -- 3623 - 0xe27  :    0 - 0x0
    "01100011", -- 3624 - 0xe28  :   99 - 0x63 -- Background 0xc5
    "01100011", -- 3625 - 0xe29  :   99 - 0x63
    "01100011", -- 3626 - 0xe2a  :   99 - 0x63
    "01110111", -- 3627 - 0xe2b  :  119 - 0x77
    "00111110", -- 3628 - 0xe2c  :   62 - 0x3e
    "00011100", -- 3629 - 0xe2d  :   28 - 0x1c
    "00001000", -- 3630 - 0xe2e  :    8 - 0x8
    "00000000", -- 3631 - 0xe2f  :    0 - 0x0
    "01111110", -- 3632 - 0xe30  :  126 - 0x7e -- Background 0xc6
    "01100011", -- 3633 - 0xe31  :   99 - 0x63
    "01100011", -- 3634 - 0xe32  :   99 - 0x63
    "01100111", -- 3635 - 0xe33  :  103 - 0x67
    "01111100", -- 3636 - 0xe34  :  124 - 0x7c
    "01101110", -- 3637 - 0xe35  :  110 - 0x6e
    "01100111", -- 3638 - 0xe36  :  103 - 0x67
    "00000000", -- 3639 - 0xe37  :    0 - 0x0
    "00110011", -- 3640 - 0xe38  :   51 - 0x33 -- Background 0xc7
    "00110011", -- 3641 - 0xe39  :   51 - 0x33
    "00110011", -- 3642 - 0xe3a  :   51 - 0x33
    "00011110", -- 3643 - 0xe3b  :   30 - 0x1e
    "00001100", -- 3644 - 0xe3c  :   12 - 0xc
    "00001100", -- 3645 - 0xe3d  :   12 - 0xc
    "00001100", -- 3646 - 0xe3e  :   12 - 0xc
    "00000000", -- 3647 - 0xe3f  :    0 - 0x0
    "00000000", -- 3648 - 0xe40  :    0 - 0x0 -- Background 0xc8
    "00000000", -- 3649 - 0xe41  :    0 - 0x0
    "00000000", -- 3650 - 0xe42  :    0 - 0x0
    "00000000", -- 3651 - 0xe43  :    0 - 0x0
    "00000000", -- 3652 - 0xe44  :    0 - 0x0
    "00000000", -- 3653 - 0xe45  :    0 - 0x0
    "00000000", -- 3654 - 0xe46  :    0 - 0x0
    "00000000", -- 3655 - 0xe47  :    0 - 0x0
    "00000000", -- 3656 - 0xe48  :    0 - 0x0 -- Background 0xc9
    "00000000", -- 3657 - 0xe49  :    0 - 0x0
    "00000000", -- 3658 - 0xe4a  :    0 - 0x0
    "00000000", -- 3659 - 0xe4b  :    0 - 0x0
    "00000000", -- 3660 - 0xe4c  :    0 - 0x0
    "00000000", -- 3661 - 0xe4d  :    0 - 0x0
    "00000000", -- 3662 - 0xe4e  :    0 - 0x0
    "00000000", -- 3663 - 0xe4f  :    0 - 0x0
    "00000000", -- 3664 - 0xe50  :    0 - 0x0 -- Background 0xca
    "00000000", -- 3665 - 0xe51  :    0 - 0x0
    "00000000", -- 3666 - 0xe52  :    0 - 0x0
    "00000000", -- 3667 - 0xe53  :    0 - 0x0
    "00000000", -- 3668 - 0xe54  :    0 - 0x0
    "00000000", -- 3669 - 0xe55  :    0 - 0x0
    "00000000", -- 3670 - 0xe56  :    0 - 0x0
    "00000000", -- 3671 - 0xe57  :    0 - 0x0
    "00000000", -- 3672 - 0xe58  :    0 - 0x0 -- Background 0xcb
    "00000000", -- 3673 - 0xe59  :    0 - 0x0
    "00000000", -- 3674 - 0xe5a  :    0 - 0x0
    "00000000", -- 3675 - 0xe5b  :    0 - 0x0
    "00000000", -- 3676 - 0xe5c  :    0 - 0x0
    "00000000", -- 3677 - 0xe5d  :    0 - 0x0
    "00000000", -- 3678 - 0xe5e  :    0 - 0x0
    "00000000", -- 3679 - 0xe5f  :    0 - 0x0
    "00000000", -- 3680 - 0xe60  :    0 - 0x0 -- Background 0xcc
    "00000000", -- 3681 - 0xe61  :    0 - 0x0
    "00000000", -- 3682 - 0xe62  :    0 - 0x0
    "00000000", -- 3683 - 0xe63  :    0 - 0x0
    "00000000", -- 3684 - 0xe64  :    0 - 0x0
    "00000000", -- 3685 - 0xe65  :    0 - 0x0
    "00000000", -- 3686 - 0xe66  :    0 - 0x0
    "00000000", -- 3687 - 0xe67  :    0 - 0x0
    "00000000", -- 3688 - 0xe68  :    0 - 0x0 -- Background 0xcd
    "00000000", -- 3689 - 0xe69  :    0 - 0x0
    "00000000", -- 3690 - 0xe6a  :    0 - 0x0
    "00000000", -- 3691 - 0xe6b  :    0 - 0x0
    "00000000", -- 3692 - 0xe6c  :    0 - 0x0
    "00000000", -- 3693 - 0xe6d  :    0 - 0x0
    "00000000", -- 3694 - 0xe6e  :    0 - 0x0
    "00000000", -- 3695 - 0xe6f  :    0 - 0x0
    "00000000", -- 3696 - 0xe70  :    0 - 0x0 -- Background 0xce
    "00000000", -- 3697 - 0xe71  :    0 - 0x0
    "00000000", -- 3698 - 0xe72  :    0 - 0x0
    "00000000", -- 3699 - 0xe73  :    0 - 0x0
    "00000000", -- 3700 - 0xe74  :    0 - 0x0
    "00000000", -- 3701 - 0xe75  :    0 - 0x0
    "00000000", -- 3702 - 0xe76  :    0 - 0x0
    "00000000", -- 3703 - 0xe77  :    0 - 0x0
    "00000000", -- 3704 - 0xe78  :    0 - 0x0 -- Background 0xcf
    "00000000", -- 3705 - 0xe79  :    0 - 0x0
    "00000000", -- 3706 - 0xe7a  :    0 - 0x0
    "00000000", -- 3707 - 0xe7b  :    0 - 0x0
    "00000000", -- 3708 - 0xe7c  :    0 - 0x0
    "00000000", -- 3709 - 0xe7d  :    0 - 0x0
    "00000000", -- 3710 - 0xe7e  :    0 - 0x0
    "00000000", -- 3711 - 0xe7f  :    0 - 0x0
    "11111111", -- 3712 - 0xe80  :  255 - 0xff -- Background 0xd0
    "11111111", -- 3713 - 0xe81  :  255 - 0xff
    "11111111", -- 3714 - 0xe82  :  255 - 0xff
    "11111111", -- 3715 - 0xe83  :  255 - 0xff
    "11111111", -- 3716 - 0xe84  :  255 - 0xff
    "11111111", -- 3717 - 0xe85  :  255 - 0xff
    "11111111", -- 3718 - 0xe86  :  255 - 0xff
    "11111111", -- 3719 - 0xe87  :  255 - 0xff
    "11111111", -- 3720 - 0xe88  :  255 - 0xff -- Background 0xd1
    "11111111", -- 3721 - 0xe89  :  255 - 0xff
    "11111111", -- 3722 - 0xe8a  :  255 - 0xff
    "11111111", -- 3723 - 0xe8b  :  255 - 0xff
    "11111111", -- 3724 - 0xe8c  :  255 - 0xff
    "11111111", -- 3725 - 0xe8d  :  255 - 0xff
    "11111111", -- 3726 - 0xe8e  :  255 - 0xff
    "11111111", -- 3727 - 0xe8f  :  255 - 0xff
    "11111111", -- 3728 - 0xe90  :  255 - 0xff -- Background 0xd2
    "11111111", -- 3729 - 0xe91  :  255 - 0xff
    "11111111", -- 3730 - 0xe92  :  255 - 0xff
    "11111111", -- 3731 - 0xe93  :  255 - 0xff
    "11111111", -- 3732 - 0xe94  :  255 - 0xff
    "11111111", -- 3733 - 0xe95  :  255 - 0xff
    "11111111", -- 3734 - 0xe96  :  255 - 0xff
    "11111111", -- 3735 - 0xe97  :  255 - 0xff
    "11111111", -- 3736 - 0xe98  :  255 - 0xff -- Background 0xd3
    "11111111", -- 3737 - 0xe99  :  255 - 0xff
    "11111111", -- 3738 - 0xe9a  :  255 - 0xff
    "11111111", -- 3739 - 0xe9b  :  255 - 0xff
    "11111111", -- 3740 - 0xe9c  :  255 - 0xff
    "11111111", -- 3741 - 0xe9d  :  255 - 0xff
    "11111111", -- 3742 - 0xe9e  :  255 - 0xff
    "11111111", -- 3743 - 0xe9f  :  255 - 0xff
    "11111111", -- 3744 - 0xea0  :  255 - 0xff -- Background 0xd4
    "11111111", -- 3745 - 0xea1  :  255 - 0xff
    "11111111", -- 3746 - 0xea2  :  255 - 0xff
    "11111111", -- 3747 - 0xea3  :  255 - 0xff
    "11111111", -- 3748 - 0xea4  :  255 - 0xff
    "11111111", -- 3749 - 0xea5  :  255 - 0xff
    "11111111", -- 3750 - 0xea6  :  255 - 0xff
    "11111111", -- 3751 - 0xea7  :  255 - 0xff
    "11111111", -- 3752 - 0xea8  :  255 - 0xff -- Background 0xd5
    "11111111", -- 3753 - 0xea9  :  255 - 0xff
    "11111111", -- 3754 - 0xeaa  :  255 - 0xff
    "11111111", -- 3755 - 0xeab  :  255 - 0xff
    "11111111", -- 3756 - 0xeac  :  255 - 0xff
    "11111111", -- 3757 - 0xead  :  255 - 0xff
    "11111111", -- 3758 - 0xeae  :  255 - 0xff
    "11111111", -- 3759 - 0xeaf  :  255 - 0xff
    "11111111", -- 3760 - 0xeb0  :  255 - 0xff -- Background 0xd6
    "11111111", -- 3761 - 0xeb1  :  255 - 0xff
    "11111111", -- 3762 - 0xeb2  :  255 - 0xff
    "11111111", -- 3763 - 0xeb3  :  255 - 0xff
    "11111111", -- 3764 - 0xeb4  :  255 - 0xff
    "11111111", -- 3765 - 0xeb5  :  255 - 0xff
    "11111111", -- 3766 - 0xeb6  :  255 - 0xff
    "11111111", -- 3767 - 0xeb7  :  255 - 0xff
    "11111111", -- 3768 - 0xeb8  :  255 - 0xff -- Background 0xd7
    "11111111", -- 3769 - 0xeb9  :  255 - 0xff
    "11111111", -- 3770 - 0xeba  :  255 - 0xff
    "11111111", -- 3771 - 0xebb  :  255 - 0xff
    "11111111", -- 3772 - 0xebc  :  255 - 0xff
    "11111111", -- 3773 - 0xebd  :  255 - 0xff
    "11111111", -- 3774 - 0xebe  :  255 - 0xff
    "11111111", -- 3775 - 0xebf  :  255 - 0xff
    "11111111", -- 3776 - 0xec0  :  255 - 0xff -- Background 0xd8
    "11111111", -- 3777 - 0xec1  :  255 - 0xff
    "11111111", -- 3778 - 0xec2  :  255 - 0xff
    "11111111", -- 3779 - 0xec3  :  255 - 0xff
    "11111111", -- 3780 - 0xec4  :  255 - 0xff
    "11111111", -- 3781 - 0xec5  :  255 - 0xff
    "11111111", -- 3782 - 0xec6  :  255 - 0xff
    "11111111", -- 3783 - 0xec7  :  255 - 0xff
    "11111111", -- 3784 - 0xec8  :  255 - 0xff -- Background 0xd9
    "11111111", -- 3785 - 0xec9  :  255 - 0xff
    "11111111", -- 3786 - 0xeca  :  255 - 0xff
    "11111111", -- 3787 - 0xecb  :  255 - 0xff
    "11111111", -- 3788 - 0xecc  :  255 - 0xff
    "11111111", -- 3789 - 0xecd  :  255 - 0xff
    "11111111", -- 3790 - 0xece  :  255 - 0xff
    "11111111", -- 3791 - 0xecf  :  255 - 0xff
    "11111111", -- 3792 - 0xed0  :  255 - 0xff -- Background 0xda
    "11111111", -- 3793 - 0xed1  :  255 - 0xff
    "11111111", -- 3794 - 0xed2  :  255 - 0xff
    "11111111", -- 3795 - 0xed3  :  255 - 0xff
    "11111111", -- 3796 - 0xed4  :  255 - 0xff
    "11111111", -- 3797 - 0xed5  :  255 - 0xff
    "11111111", -- 3798 - 0xed6  :  255 - 0xff
    "11111111", -- 3799 - 0xed7  :  255 - 0xff
    "11111111", -- 3800 - 0xed8  :  255 - 0xff -- Background 0xdb
    "11111111", -- 3801 - 0xed9  :  255 - 0xff
    "11111111", -- 3802 - 0xeda  :  255 - 0xff
    "11111111", -- 3803 - 0xedb  :  255 - 0xff
    "11111111", -- 3804 - 0xedc  :  255 - 0xff
    "11111111", -- 3805 - 0xedd  :  255 - 0xff
    "11111111", -- 3806 - 0xede  :  255 - 0xff
    "11111111", -- 3807 - 0xedf  :  255 - 0xff
    "11111111", -- 3808 - 0xee0  :  255 - 0xff -- Background 0xdc
    "11111111", -- 3809 - 0xee1  :  255 - 0xff
    "11111111", -- 3810 - 0xee2  :  255 - 0xff
    "11111111", -- 3811 - 0xee3  :  255 - 0xff
    "11111111", -- 3812 - 0xee4  :  255 - 0xff
    "11111111", -- 3813 - 0xee5  :  255 - 0xff
    "11111111", -- 3814 - 0xee6  :  255 - 0xff
    "11111111", -- 3815 - 0xee7  :  255 - 0xff
    "11111111", -- 3816 - 0xee8  :  255 - 0xff -- Background 0xdd
    "11111111", -- 3817 - 0xee9  :  255 - 0xff
    "11111111", -- 3818 - 0xeea  :  255 - 0xff
    "11111111", -- 3819 - 0xeeb  :  255 - 0xff
    "11111111", -- 3820 - 0xeec  :  255 - 0xff
    "11111111", -- 3821 - 0xeed  :  255 - 0xff
    "11111111", -- 3822 - 0xeee  :  255 - 0xff
    "11111111", -- 3823 - 0xeef  :  255 - 0xff
    "11111111", -- 3824 - 0xef0  :  255 - 0xff -- Background 0xde
    "11111111", -- 3825 - 0xef1  :  255 - 0xff
    "11111111", -- 3826 - 0xef2  :  255 - 0xff
    "11111111", -- 3827 - 0xef3  :  255 - 0xff
    "11111111", -- 3828 - 0xef4  :  255 - 0xff
    "11111111", -- 3829 - 0xef5  :  255 - 0xff
    "11111111", -- 3830 - 0xef6  :  255 - 0xff
    "11111111", -- 3831 - 0xef7  :  255 - 0xff
    "11111111", -- 3832 - 0xef8  :  255 - 0xff -- Background 0xdf
    "11111111", -- 3833 - 0xef9  :  255 - 0xff
    "11111111", -- 3834 - 0xefa  :  255 - 0xff
    "11111111", -- 3835 - 0xefb  :  255 - 0xff
    "11111111", -- 3836 - 0xefc  :  255 - 0xff
    "11111111", -- 3837 - 0xefd  :  255 - 0xff
    "11111111", -- 3838 - 0xefe  :  255 - 0xff
    "11111111", -- 3839 - 0xeff  :  255 - 0xff
    "11111111", -- 3840 - 0xf00  :  255 - 0xff -- Background 0xe0
    "11111111", -- 3841 - 0xf01  :  255 - 0xff
    "11111111", -- 3842 - 0xf02  :  255 - 0xff
    "11111111", -- 3843 - 0xf03  :  255 - 0xff
    "11111111", -- 3844 - 0xf04  :  255 - 0xff
    "11111111", -- 3845 - 0xf05  :  255 - 0xff
    "11111111", -- 3846 - 0xf06  :  255 - 0xff
    "11111111", -- 3847 - 0xf07  :  255 - 0xff
    "11111111", -- 3848 - 0xf08  :  255 - 0xff -- Background 0xe1
    "11111111", -- 3849 - 0xf09  :  255 - 0xff
    "11111111", -- 3850 - 0xf0a  :  255 - 0xff
    "11111111", -- 3851 - 0xf0b  :  255 - 0xff
    "11111111", -- 3852 - 0xf0c  :  255 - 0xff
    "11111111", -- 3853 - 0xf0d  :  255 - 0xff
    "11111111", -- 3854 - 0xf0e  :  255 - 0xff
    "11111111", -- 3855 - 0xf0f  :  255 - 0xff
    "11111111", -- 3856 - 0xf10  :  255 - 0xff -- Background 0xe2
    "11111111", -- 3857 - 0xf11  :  255 - 0xff
    "11111111", -- 3858 - 0xf12  :  255 - 0xff
    "11111111", -- 3859 - 0xf13  :  255 - 0xff
    "11111111", -- 3860 - 0xf14  :  255 - 0xff
    "11111111", -- 3861 - 0xf15  :  255 - 0xff
    "11111111", -- 3862 - 0xf16  :  255 - 0xff
    "11111111", -- 3863 - 0xf17  :  255 - 0xff
    "11111111", -- 3864 - 0xf18  :  255 - 0xff -- Background 0xe3
    "11111111", -- 3865 - 0xf19  :  255 - 0xff
    "11111111", -- 3866 - 0xf1a  :  255 - 0xff
    "11111111", -- 3867 - 0xf1b  :  255 - 0xff
    "11111111", -- 3868 - 0xf1c  :  255 - 0xff
    "11111111", -- 3869 - 0xf1d  :  255 - 0xff
    "11111111", -- 3870 - 0xf1e  :  255 - 0xff
    "11111111", -- 3871 - 0xf1f  :  255 - 0xff
    "11111111", -- 3872 - 0xf20  :  255 - 0xff -- Background 0xe4
    "11111111", -- 3873 - 0xf21  :  255 - 0xff
    "11111111", -- 3874 - 0xf22  :  255 - 0xff
    "11111111", -- 3875 - 0xf23  :  255 - 0xff
    "11111111", -- 3876 - 0xf24  :  255 - 0xff
    "11111111", -- 3877 - 0xf25  :  255 - 0xff
    "11111111", -- 3878 - 0xf26  :  255 - 0xff
    "11111111", -- 3879 - 0xf27  :  255 - 0xff
    "11111111", -- 3880 - 0xf28  :  255 - 0xff -- Background 0xe5
    "11111111", -- 3881 - 0xf29  :  255 - 0xff
    "11111111", -- 3882 - 0xf2a  :  255 - 0xff
    "11111111", -- 3883 - 0xf2b  :  255 - 0xff
    "11111111", -- 3884 - 0xf2c  :  255 - 0xff
    "11111111", -- 3885 - 0xf2d  :  255 - 0xff
    "11111111", -- 3886 - 0xf2e  :  255 - 0xff
    "11111111", -- 3887 - 0xf2f  :  255 - 0xff
    "11111111", -- 3888 - 0xf30  :  255 - 0xff -- Background 0xe6
    "11111111", -- 3889 - 0xf31  :  255 - 0xff
    "11111111", -- 3890 - 0xf32  :  255 - 0xff
    "11111111", -- 3891 - 0xf33  :  255 - 0xff
    "11111111", -- 3892 - 0xf34  :  255 - 0xff
    "11111111", -- 3893 - 0xf35  :  255 - 0xff
    "11111111", -- 3894 - 0xf36  :  255 - 0xff
    "11111111", -- 3895 - 0xf37  :  255 - 0xff
    "11111111", -- 3896 - 0xf38  :  255 - 0xff -- Background 0xe7
    "11111111", -- 3897 - 0xf39  :  255 - 0xff
    "11111111", -- 3898 - 0xf3a  :  255 - 0xff
    "11111111", -- 3899 - 0xf3b  :  255 - 0xff
    "11111111", -- 3900 - 0xf3c  :  255 - 0xff
    "11111111", -- 3901 - 0xf3d  :  255 - 0xff
    "11111111", -- 3902 - 0xf3e  :  255 - 0xff
    "11111111", -- 3903 - 0xf3f  :  255 - 0xff
    "11111111", -- 3904 - 0xf40  :  255 - 0xff -- Background 0xe8
    "11111111", -- 3905 - 0xf41  :  255 - 0xff
    "11111111", -- 3906 - 0xf42  :  255 - 0xff
    "11111111", -- 3907 - 0xf43  :  255 - 0xff
    "11111111", -- 3908 - 0xf44  :  255 - 0xff
    "11111111", -- 3909 - 0xf45  :  255 - 0xff
    "11111111", -- 3910 - 0xf46  :  255 - 0xff
    "11111111", -- 3911 - 0xf47  :  255 - 0xff
    "11111111", -- 3912 - 0xf48  :  255 - 0xff -- Background 0xe9
    "11111111", -- 3913 - 0xf49  :  255 - 0xff
    "11111111", -- 3914 - 0xf4a  :  255 - 0xff
    "11111111", -- 3915 - 0xf4b  :  255 - 0xff
    "11111111", -- 3916 - 0xf4c  :  255 - 0xff
    "11111111", -- 3917 - 0xf4d  :  255 - 0xff
    "11111111", -- 3918 - 0xf4e  :  255 - 0xff
    "11111111", -- 3919 - 0xf4f  :  255 - 0xff
    "11111111", -- 3920 - 0xf50  :  255 - 0xff -- Background 0xea
    "11111111", -- 3921 - 0xf51  :  255 - 0xff
    "11111111", -- 3922 - 0xf52  :  255 - 0xff
    "11111111", -- 3923 - 0xf53  :  255 - 0xff
    "11111111", -- 3924 - 0xf54  :  255 - 0xff
    "11111111", -- 3925 - 0xf55  :  255 - 0xff
    "11111111", -- 3926 - 0xf56  :  255 - 0xff
    "11111111", -- 3927 - 0xf57  :  255 - 0xff
    "11111111", -- 3928 - 0xf58  :  255 - 0xff -- Background 0xeb
    "11111111", -- 3929 - 0xf59  :  255 - 0xff
    "11111111", -- 3930 - 0xf5a  :  255 - 0xff
    "11111111", -- 3931 - 0xf5b  :  255 - 0xff
    "11111111", -- 3932 - 0xf5c  :  255 - 0xff
    "11111111", -- 3933 - 0xf5d  :  255 - 0xff
    "11111111", -- 3934 - 0xf5e  :  255 - 0xff
    "11111111", -- 3935 - 0xf5f  :  255 - 0xff
    "11111111", -- 3936 - 0xf60  :  255 - 0xff -- Background 0xec
    "11111111", -- 3937 - 0xf61  :  255 - 0xff
    "11111111", -- 3938 - 0xf62  :  255 - 0xff
    "11111111", -- 3939 - 0xf63  :  255 - 0xff
    "11111111", -- 3940 - 0xf64  :  255 - 0xff
    "11111111", -- 3941 - 0xf65  :  255 - 0xff
    "11111111", -- 3942 - 0xf66  :  255 - 0xff
    "11111111", -- 3943 - 0xf67  :  255 - 0xff
    "11111111", -- 3944 - 0xf68  :  255 - 0xff -- Background 0xed
    "11111111", -- 3945 - 0xf69  :  255 - 0xff
    "11111111", -- 3946 - 0xf6a  :  255 - 0xff
    "11111111", -- 3947 - 0xf6b  :  255 - 0xff
    "11111111", -- 3948 - 0xf6c  :  255 - 0xff
    "11111111", -- 3949 - 0xf6d  :  255 - 0xff
    "11111111", -- 3950 - 0xf6e  :  255 - 0xff
    "11111111", -- 3951 - 0xf6f  :  255 - 0xff
    "11111111", -- 3952 - 0xf70  :  255 - 0xff -- Background 0xee
    "11111111", -- 3953 - 0xf71  :  255 - 0xff
    "11111111", -- 3954 - 0xf72  :  255 - 0xff
    "11111111", -- 3955 - 0xf73  :  255 - 0xff
    "11111111", -- 3956 - 0xf74  :  255 - 0xff
    "11111111", -- 3957 - 0xf75  :  255 - 0xff
    "11111111", -- 3958 - 0xf76  :  255 - 0xff
    "11111111", -- 3959 - 0xf77  :  255 - 0xff
    "11111111", -- 3960 - 0xf78  :  255 - 0xff -- Background 0xef
    "11111111", -- 3961 - 0xf79  :  255 - 0xff
    "11111111", -- 3962 - 0xf7a  :  255 - 0xff
    "11111111", -- 3963 - 0xf7b  :  255 - 0xff
    "11111111", -- 3964 - 0xf7c  :  255 - 0xff
    "11111111", -- 3965 - 0xf7d  :  255 - 0xff
    "11111111", -- 3966 - 0xf7e  :  255 - 0xff
    "11111111", -- 3967 - 0xf7f  :  255 - 0xff
    "11111111", -- 3968 - 0xf80  :  255 - 0xff -- Background 0xf0
    "11111111", -- 3969 - 0xf81  :  255 - 0xff
    "11111111", -- 3970 - 0xf82  :  255 - 0xff
    "11111111", -- 3971 - 0xf83  :  255 - 0xff
    "11111111", -- 3972 - 0xf84  :  255 - 0xff
    "11111111", -- 3973 - 0xf85  :  255 - 0xff
    "11111111", -- 3974 - 0xf86  :  255 - 0xff
    "11111111", -- 3975 - 0xf87  :  255 - 0xff
    "11111111", -- 3976 - 0xf88  :  255 - 0xff -- Background 0xf1
    "11111111", -- 3977 - 0xf89  :  255 - 0xff
    "11111111", -- 3978 - 0xf8a  :  255 - 0xff
    "11111111", -- 3979 - 0xf8b  :  255 - 0xff
    "11111111", -- 3980 - 0xf8c  :  255 - 0xff
    "11111111", -- 3981 - 0xf8d  :  255 - 0xff
    "11111111", -- 3982 - 0xf8e  :  255 - 0xff
    "11111111", -- 3983 - 0xf8f  :  255 - 0xff
    "11111111", -- 3984 - 0xf90  :  255 - 0xff -- Background 0xf2
    "11111111", -- 3985 - 0xf91  :  255 - 0xff
    "11111111", -- 3986 - 0xf92  :  255 - 0xff
    "11111111", -- 3987 - 0xf93  :  255 - 0xff
    "11111111", -- 3988 - 0xf94  :  255 - 0xff
    "11111111", -- 3989 - 0xf95  :  255 - 0xff
    "11111111", -- 3990 - 0xf96  :  255 - 0xff
    "11111111", -- 3991 - 0xf97  :  255 - 0xff
    "11111111", -- 3992 - 0xf98  :  255 - 0xff -- Background 0xf3
    "11111111", -- 3993 - 0xf99  :  255 - 0xff
    "11111111", -- 3994 - 0xf9a  :  255 - 0xff
    "11111111", -- 3995 - 0xf9b  :  255 - 0xff
    "11111111", -- 3996 - 0xf9c  :  255 - 0xff
    "11111111", -- 3997 - 0xf9d  :  255 - 0xff
    "11111111", -- 3998 - 0xf9e  :  255 - 0xff
    "11111111", -- 3999 - 0xf9f  :  255 - 0xff
    "11111111", -- 4000 - 0xfa0  :  255 - 0xff -- Background 0xf4
    "11111111", -- 4001 - 0xfa1  :  255 - 0xff
    "11111111", -- 4002 - 0xfa2  :  255 - 0xff
    "11111111", -- 4003 - 0xfa3  :  255 - 0xff
    "11111111", -- 4004 - 0xfa4  :  255 - 0xff
    "11111111", -- 4005 - 0xfa5  :  255 - 0xff
    "11111111", -- 4006 - 0xfa6  :  255 - 0xff
    "11111111", -- 4007 - 0xfa7  :  255 - 0xff
    "11111111", -- 4008 - 0xfa8  :  255 - 0xff -- Background 0xf5
    "11111111", -- 4009 - 0xfa9  :  255 - 0xff
    "11111111", -- 4010 - 0xfaa  :  255 - 0xff
    "11111111", -- 4011 - 0xfab  :  255 - 0xff
    "11111111", -- 4012 - 0xfac  :  255 - 0xff
    "11111111", -- 4013 - 0xfad  :  255 - 0xff
    "11111111", -- 4014 - 0xfae  :  255 - 0xff
    "11111111", -- 4015 - 0xfaf  :  255 - 0xff
    "11111111", -- 4016 - 0xfb0  :  255 - 0xff -- Background 0xf6
    "11111111", -- 4017 - 0xfb1  :  255 - 0xff
    "11111111", -- 4018 - 0xfb2  :  255 - 0xff
    "11111111", -- 4019 - 0xfb3  :  255 - 0xff
    "11111111", -- 4020 - 0xfb4  :  255 - 0xff
    "11111111", -- 4021 - 0xfb5  :  255 - 0xff
    "11111111", -- 4022 - 0xfb6  :  255 - 0xff
    "11111111", -- 4023 - 0xfb7  :  255 - 0xff
    "11111111", -- 4024 - 0xfb8  :  255 - 0xff -- Background 0xf7
    "11111111", -- 4025 - 0xfb9  :  255 - 0xff
    "11111111", -- 4026 - 0xfba  :  255 - 0xff
    "11111111", -- 4027 - 0xfbb  :  255 - 0xff
    "11111111", -- 4028 - 0xfbc  :  255 - 0xff
    "11111111", -- 4029 - 0xfbd  :  255 - 0xff
    "11111111", -- 4030 - 0xfbe  :  255 - 0xff
    "11111111", -- 4031 - 0xfbf  :  255 - 0xff
    "11111111", -- 4032 - 0xfc0  :  255 - 0xff -- Background 0xf8
    "11111111", -- 4033 - 0xfc1  :  255 - 0xff
    "11111111", -- 4034 - 0xfc2  :  255 - 0xff
    "11111111", -- 4035 - 0xfc3  :  255 - 0xff
    "11111111", -- 4036 - 0xfc4  :  255 - 0xff
    "11111111", -- 4037 - 0xfc5  :  255 - 0xff
    "11111111", -- 4038 - 0xfc6  :  255 - 0xff
    "11111111", -- 4039 - 0xfc7  :  255 - 0xff
    "11111111", -- 4040 - 0xfc8  :  255 - 0xff -- Background 0xf9
    "11111111", -- 4041 - 0xfc9  :  255 - 0xff
    "11111111", -- 4042 - 0xfca  :  255 - 0xff
    "11111111", -- 4043 - 0xfcb  :  255 - 0xff
    "11111111", -- 4044 - 0xfcc  :  255 - 0xff
    "11111111", -- 4045 - 0xfcd  :  255 - 0xff
    "11111111", -- 4046 - 0xfce  :  255 - 0xff
    "11111111", -- 4047 - 0xfcf  :  255 - 0xff
    "11111111", -- 4048 - 0xfd0  :  255 - 0xff -- Background 0xfa
    "11111111", -- 4049 - 0xfd1  :  255 - 0xff
    "11111111", -- 4050 - 0xfd2  :  255 - 0xff
    "11111111", -- 4051 - 0xfd3  :  255 - 0xff
    "11111111", -- 4052 - 0xfd4  :  255 - 0xff
    "11111111", -- 4053 - 0xfd5  :  255 - 0xff
    "11111111", -- 4054 - 0xfd6  :  255 - 0xff
    "11111111", -- 4055 - 0xfd7  :  255 - 0xff
    "11111111", -- 4056 - 0xfd8  :  255 - 0xff -- Background 0xfb
    "11111111", -- 4057 - 0xfd9  :  255 - 0xff
    "11111111", -- 4058 - 0xfda  :  255 - 0xff
    "11111111", -- 4059 - 0xfdb  :  255 - 0xff
    "11111111", -- 4060 - 0xfdc  :  255 - 0xff
    "11111111", -- 4061 - 0xfdd  :  255 - 0xff
    "11111111", -- 4062 - 0xfde  :  255 - 0xff
    "11111111", -- 4063 - 0xfdf  :  255 - 0xff
    "11111111", -- 4064 - 0xfe0  :  255 - 0xff -- Background 0xfc
    "11111111", -- 4065 - 0xfe1  :  255 - 0xff
    "11111111", -- 4066 - 0xfe2  :  255 - 0xff
    "11111111", -- 4067 - 0xfe3  :  255 - 0xff
    "11111111", -- 4068 - 0xfe4  :  255 - 0xff
    "11111111", -- 4069 - 0xfe5  :  255 - 0xff
    "11111111", -- 4070 - 0xfe6  :  255 - 0xff
    "11111111", -- 4071 - 0xfe7  :  255 - 0xff
    "11111111", -- 4072 - 0xfe8  :  255 - 0xff -- Background 0xfd
    "11111111", -- 4073 - 0xfe9  :  255 - 0xff
    "11111111", -- 4074 - 0xfea  :  255 - 0xff
    "11111111", -- 4075 - 0xfeb  :  255 - 0xff
    "11111111", -- 4076 - 0xfec  :  255 - 0xff
    "11111111", -- 4077 - 0xfed  :  255 - 0xff
    "11111111", -- 4078 - 0xfee  :  255 - 0xff
    "11111111", -- 4079 - 0xfef  :  255 - 0xff
    "11111111", -- 4080 - 0xff0  :  255 - 0xff -- Background 0xfe
    "11111111", -- 4081 - 0xff1  :  255 - 0xff
    "11111111", -- 4082 - 0xff2  :  255 - 0xff
    "11111111", -- 4083 - 0xff3  :  255 - 0xff
    "11111111", -- 4084 - 0xff4  :  255 - 0xff
    "11111111", -- 4085 - 0xff5  :  255 - 0xff
    "11111111", -- 4086 - 0xff6  :  255 - 0xff
    "11111111", -- 4087 - 0xff7  :  255 - 0xff
    "11111111", -- 4088 - 0xff8  :  255 - 0xff -- Background 0xff
    "11111111", -- 4089 - 0xff9  :  255 - 0xff
    "11111111", -- 4090 - 0xffa  :  255 - 0xff
    "11111111", -- 4091 - 0xffb  :  255 - 0xff
    "11111111", -- 4092 - 0xffc  :  255 - 0xff
    "11111111", -- 4093 - 0xffd  :  255 - 0xff
    "11111111", -- 4094 - 0xffe  :  255 - 0xff
    "11111111"  -- 4095 - 0xfff  :  255 - 0xff
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
