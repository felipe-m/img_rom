//-   Background Pattern table BOTH COLOR PLANES
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
//- Autcmatically generated verilog ROM from a NES memory file----


//-  Original memory dump file name: sprilo_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_PTABLE_SPRILO_BG
  (
     input     clk,   // clock
     input      [12-1:0] addr,  //4096 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Background pattern Table both color planes
      12'h0: dout <= 8'b00111110; //    0 :  62 - 0x3e -- Background 0x0
      12'h1: dout <= 8'b01111111; //    1 : 127 - 0x7f
      12'h2: dout <= 8'b01110111; //    2 : 119 - 0x77
      12'h3: dout <= 8'b01111111; //    3 : 127 - 0x7f
      12'h4: dout <= 8'b01111111; //    4 : 127 - 0x7f
      12'h5: dout <= 8'b01110111; //    5 : 119 - 0x77
      12'h6: dout <= 8'b01111111; //    6 : 127 - 0x7f
      12'h7: dout <= 8'b00111110; //    7 :  62 - 0x3e
      12'h8: dout <= 8'b11000011; //    8 : 195 - 0xc3 -- plane 1
      12'h9: dout <= 8'b10000001; //    9 : 129 - 0x81
      12'hA: dout <= 8'b10011001; //   10 : 153 - 0x99
      12'hB: dout <= 8'b10010001; //   11 : 145 - 0x91
      12'hC: dout <= 8'b10001001; //   12 : 137 - 0x89
      12'hD: dout <= 8'b10011001; //   13 : 153 - 0x99
      12'hE: dout <= 8'b10000001; //   14 : 129 - 0x81
      12'hF: dout <= 8'b11000011; //   15 : 195 - 0xc3
      12'h10: dout <= 8'b00011100; //   16 :  28 - 0x1c -- Background 0x1
      12'h11: dout <= 8'b00111100; //   17 :  60 - 0x3c
      12'h12: dout <= 8'b01111100; //   18 : 124 - 0x7c
      12'h13: dout <= 8'b00011100; //   19 :  28 - 0x1c
      12'h14: dout <= 8'b00011100; //   20 :  28 - 0x1c
      12'h15: dout <= 8'b00011100; //   21 :  28 - 0x1c
      12'h16: dout <= 8'b01111111; //   22 : 127 - 0x7f
      12'h17: dout <= 8'b01111111; //   23 : 127 - 0x7f
      12'h18: dout <= 8'b11100111; //   24 : 231 - 0xe7 -- plane 1
      12'h19: dout <= 8'b11000111; //   25 : 199 - 0xc7
      12'h1A: dout <= 8'b10000111; //   26 : 135 - 0x87
      12'h1B: dout <= 8'b11100111; //   27 : 231 - 0xe7
      12'h1C: dout <= 8'b11100111; //   28 : 231 - 0xe7
      12'h1D: dout <= 8'b11100111; //   29 : 231 - 0xe7
      12'h1E: dout <= 8'b10000001; //   30 : 129 - 0x81
      12'h1F: dout <= 8'b10000001; //   31 : 129 - 0x81
      12'h20: dout <= 8'b00111110; //   32 :  62 - 0x3e -- Background 0x2
      12'h21: dout <= 8'b01111111; //   33 : 127 - 0x7f
      12'h22: dout <= 8'b00000111; //   34 :   7 - 0x7
      12'h23: dout <= 8'b00111111; //   35 :  63 - 0x3f
      12'h24: dout <= 8'b01111111; //   36 : 127 - 0x7f
      12'h25: dout <= 8'b01110000; //   37 : 112 - 0x70
      12'h26: dout <= 8'b01111111; //   38 : 127 - 0x7f
      12'h27: dout <= 8'b01111111; //   39 : 127 - 0x7f
      12'h28: dout <= 8'b11000011; //   40 : 195 - 0xc3 -- plane 1
      12'h29: dout <= 8'b10000001; //   41 : 129 - 0x81
      12'h2A: dout <= 8'b11111001; //   42 : 249 - 0xf9
      12'h2B: dout <= 8'b11000001; //   43 : 193 - 0xc1
      12'h2C: dout <= 8'b10000001; //   44 : 129 - 0x81
      12'h2D: dout <= 8'b10011111; //   45 : 159 - 0x9f
      12'h2E: dout <= 8'b10000001; //   46 : 129 - 0x81
      12'h2F: dout <= 8'b10000001; //   47 : 129 - 0x81
      12'h30: dout <= 8'b00111110; //   48 :  62 - 0x3e -- Background 0x3
      12'h31: dout <= 8'b01111111; //   49 : 127 - 0x7f
      12'h32: dout <= 8'b00000111; //   50 :   7 - 0x7
      12'h33: dout <= 8'b00011111; //   51 :  31 - 0x1f
      12'h34: dout <= 8'b00011111; //   52 :  31 - 0x1f
      12'h35: dout <= 8'b00000111; //   53 :   7 - 0x7
      12'h36: dout <= 8'b01111111; //   54 : 127 - 0x7f
      12'h37: dout <= 8'b00111110; //   55 :  62 - 0x3e
      12'h38: dout <= 8'b11000011; //   56 : 195 - 0xc3 -- plane 1
      12'h39: dout <= 8'b10000001; //   57 : 129 - 0x81
      12'h3A: dout <= 8'b11111001; //   58 : 249 - 0xf9
      12'h3B: dout <= 8'b11100001; //   59 : 225 - 0xe1
      12'h3C: dout <= 8'b11100001; //   60 : 225 - 0xe1
      12'h3D: dout <= 8'b11111001; //   61 : 249 - 0xf9
      12'h3E: dout <= 8'b10000001; //   62 : 129 - 0x81
      12'h3F: dout <= 8'b11000011; //   63 : 195 - 0xc3
      12'h40: dout <= 8'b00110000; //   64 :  48 - 0x30 -- Background 0x4
      12'h41: dout <= 8'b01110000; //   65 : 112 - 0x70
      12'h42: dout <= 8'b01110111; //   66 : 119 - 0x77
      12'h43: dout <= 8'b01110111; //   67 : 119 - 0x77
      12'h44: dout <= 8'b01111111; //   68 : 127 - 0x7f
      12'h45: dout <= 8'b01111111; //   69 : 127 - 0x7f
      12'h46: dout <= 8'b00000111; //   70 :   7 - 0x7
      12'h47: dout <= 8'b00000111; //   71 :   7 - 0x7
      12'h48: dout <= 8'b11011111; //   72 : 223 - 0xdf -- plane 1
      12'h49: dout <= 8'b10011111; //   73 : 159 - 0x9f
      12'h4A: dout <= 8'b10011001; //   74 : 153 - 0x99
      12'h4B: dout <= 8'b10011001; //   75 : 153 - 0x99
      12'h4C: dout <= 8'b10000000; //   76 : 128 - 0x80
      12'h4D: dout <= 8'b10000000; //   77 : 128 - 0x80
      12'h4E: dout <= 8'b11111001; //   78 : 249 - 0xf9
      12'h4F: dout <= 8'b11111001; //   79 : 249 - 0xf9
      12'h50: dout <= 8'b01111111; //   80 : 127 - 0x7f -- Background 0x5
      12'h51: dout <= 8'b01111111; //   81 : 127 - 0x7f
      12'h52: dout <= 8'b01110000; //   82 : 112 - 0x70
      12'h53: dout <= 8'b01111110; //   83 : 126 - 0x7e
      12'h54: dout <= 8'b01111111; //   84 : 127 - 0x7f
      12'h55: dout <= 8'b00000111; //   85 :   7 - 0x7
      12'h56: dout <= 8'b01111111; //   86 : 127 - 0x7f
      12'h57: dout <= 8'b00111110; //   87 :  62 - 0x3e
      12'h58: dout <= 8'b10000001; //   88 : 129 - 0x81 -- plane 1
      12'h59: dout <= 8'b10000001; //   89 : 129 - 0x81
      12'h5A: dout <= 8'b10011111; //   90 : 159 - 0x9f
      12'h5B: dout <= 8'b10000011; //   91 : 131 - 0x83
      12'h5C: dout <= 8'b10000001; //   92 : 129 - 0x81
      12'h5D: dout <= 8'b11111001; //   93 : 249 - 0xf9
      12'h5E: dout <= 8'b10000001; //   94 : 129 - 0x81
      12'h5F: dout <= 8'b11000011; //   95 : 195 - 0xc3
      12'h60: dout <= 8'b00111110; //   96 :  62 - 0x3e -- Background 0x6
      12'h61: dout <= 8'b01111111; //   97 : 127 - 0x7f
      12'h62: dout <= 8'b01110000; //   98 : 112 - 0x70
      12'h63: dout <= 8'b01111110; //   99 : 126 - 0x7e
      12'h64: dout <= 8'b01111111; //  100 : 127 - 0x7f
      12'h65: dout <= 8'b01110111; //  101 : 119 - 0x77
      12'h66: dout <= 8'b01111111; //  102 : 127 - 0x7f
      12'h67: dout <= 8'b00111110; //  103 :  62 - 0x3e
      12'h68: dout <= 8'b11000011; //  104 : 195 - 0xc3 -- plane 1
      12'h69: dout <= 8'b10000001; //  105 : 129 - 0x81
      12'h6A: dout <= 8'b10011111; //  106 : 159 - 0x9f
      12'h6B: dout <= 8'b10000011; //  107 : 131 - 0x83
      12'h6C: dout <= 8'b10000001; //  108 : 129 - 0x81
      12'h6D: dout <= 8'b10011001; //  109 : 153 - 0x99
      12'h6E: dout <= 8'b10000001; //  110 : 129 - 0x81
      12'h6F: dout <= 8'b11000011; //  111 : 195 - 0xc3
      12'h70: dout <= 8'b01111111; //  112 : 127 - 0x7f -- Background 0x7
      12'h71: dout <= 8'b01111111; //  113 : 127 - 0x7f
      12'h72: dout <= 8'b00000111; //  114 :   7 - 0x7
      12'h73: dout <= 8'b00001110; //  115 :  14 - 0xe
      12'h74: dout <= 8'b00001110; //  116 :  14 - 0xe
      12'h75: dout <= 8'b00011100; //  117 :  28 - 0x1c
      12'h76: dout <= 8'b00011100; //  118 :  28 - 0x1c
      12'h77: dout <= 8'b00011100; //  119 :  28 - 0x1c
      12'h78: dout <= 8'b10000001; //  120 : 129 - 0x81 -- plane 1
      12'h79: dout <= 8'b10000001; //  121 : 129 - 0x81
      12'h7A: dout <= 8'b11111001; //  122 : 249 - 0xf9
      12'h7B: dout <= 8'b11110011; //  123 : 243 - 0xf3
      12'h7C: dout <= 8'b11110011; //  124 : 243 - 0xf3
      12'h7D: dout <= 8'b11100111; //  125 : 231 - 0xe7
      12'h7E: dout <= 8'b11100111; //  126 : 231 - 0xe7
      12'h7F: dout <= 8'b11100111; //  127 : 231 - 0xe7
      12'h80: dout <= 8'b00111110; //  128 :  62 - 0x3e -- Background 0x8
      12'h81: dout <= 8'b01111111; //  129 : 127 - 0x7f
      12'h82: dout <= 8'b01110111; //  130 : 119 - 0x77
      12'h83: dout <= 8'b00111110; //  131 :  62 - 0x3e
      12'h84: dout <= 8'b01111111; //  132 : 127 - 0x7f
      12'h85: dout <= 8'b01110111; //  133 : 119 - 0x77
      12'h86: dout <= 8'b01111111; //  134 : 127 - 0x7f
      12'h87: dout <= 8'b00111110; //  135 :  62 - 0x3e
      12'h88: dout <= 8'b11000011; //  136 : 195 - 0xc3 -- plane 1
      12'h89: dout <= 8'b10000001; //  137 : 129 - 0x81
      12'h8A: dout <= 8'b10011001; //  138 : 153 - 0x99
      12'h8B: dout <= 8'b11000011; //  139 : 195 - 0xc3
      12'h8C: dout <= 8'b10000001; //  140 : 129 - 0x81
      12'h8D: dout <= 8'b10011001; //  141 : 153 - 0x99
      12'h8E: dout <= 8'b10000001; //  142 : 129 - 0x81
      12'h8F: dout <= 8'b11000011; //  143 : 195 - 0xc3
      12'h90: dout <= 8'b00111110; //  144 :  62 - 0x3e -- Background 0x9
      12'h91: dout <= 8'b01111111; //  145 : 127 - 0x7f
      12'h92: dout <= 8'b01110111; //  146 : 119 - 0x77
      12'h93: dout <= 8'b01111111; //  147 : 127 - 0x7f
      12'h94: dout <= 8'b00111111; //  148 :  63 - 0x3f
      12'h95: dout <= 8'b00000111; //  149 :   7 - 0x7
      12'h96: dout <= 8'b01111111; //  150 : 127 - 0x7f
      12'h97: dout <= 8'b00111110; //  151 :  62 - 0x3e
      12'h98: dout <= 8'b11000011; //  152 : 195 - 0xc3 -- plane 1
      12'h99: dout <= 8'b10000001; //  153 : 129 - 0x81
      12'h9A: dout <= 8'b10011001; //  154 : 153 - 0x99
      12'h9B: dout <= 8'b10000001; //  155 : 129 - 0x81
      12'h9C: dout <= 8'b11000001; //  156 : 193 - 0xc1
      12'h9D: dout <= 8'b11111001; //  157 : 249 - 0xf9
      12'h9E: dout <= 8'b10000001; //  158 : 129 - 0x81
      12'h9F: dout <= 8'b11000011; //  159 : 195 - 0xc3
      12'hA0: dout <= 8'b00000000; //  160 :   0 - 0x0 -- Background 0xa
      12'hA1: dout <= 8'b00000000; //  161 :   0 - 0x0
      12'hA2: dout <= 8'b00000000; //  162 :   0 - 0x0
      12'hA3: dout <= 8'b00000000; //  163 :   0 - 0x0
      12'hA4: dout <= 8'b00000000; //  164 :   0 - 0x0
      12'hA5: dout <= 8'b00110000; //  165 :  48 - 0x30
      12'hA6: dout <= 8'b01111000; //  166 : 120 - 0x78
      12'hA7: dout <= 8'b00110000; //  167 :  48 - 0x30
      12'hA8: dout <= 8'b11111111; //  168 : 255 - 0xff -- plane 1
      12'hA9: dout <= 8'b11111111; //  169 : 255 - 0xff
      12'hAA: dout <= 8'b11111111; //  170 : 255 - 0xff
      12'hAB: dout <= 8'b11111111; //  171 : 255 - 0xff
      12'hAC: dout <= 8'b11111111; //  172 : 255 - 0xff
      12'hAD: dout <= 8'b11011111; //  173 : 223 - 0xdf
      12'hAE: dout <= 8'b10001111; //  174 : 143 - 0x8f
      12'hAF: dout <= 8'b11011111; //  175 : 223 - 0xdf
      12'hB0: dout <= 8'b01110000; //  176 : 112 - 0x70 -- Background 0xb
      12'hB1: dout <= 8'b11111000; //  177 : 248 - 0xf8
      12'hB2: dout <= 8'b11111000; //  178 : 248 - 0xf8
      12'hB3: dout <= 8'b11111000; //  179 : 248 - 0xf8
      12'hB4: dout <= 8'b01110000; //  180 : 112 - 0x70
      12'hB5: dout <= 8'b00000000; //  181 :   0 - 0x0
      12'hB6: dout <= 8'b01110000; //  182 : 112 - 0x70
      12'hB7: dout <= 8'b01110000; //  183 : 112 - 0x70
      12'hB8: dout <= 8'b10011111; //  184 : 159 - 0x9f -- plane 1
      12'hB9: dout <= 8'b00001111; //  185 :  15 - 0xf
      12'hBA: dout <= 8'b00001111; //  186 :  15 - 0xf
      12'hBB: dout <= 8'b00001111; //  187 :  15 - 0xf
      12'hBC: dout <= 8'b10011111; //  188 : 159 - 0x9f
      12'hBD: dout <= 8'b11111111; //  189 : 255 - 0xff
      12'hBE: dout <= 8'b10011111; //  190 : 159 - 0x9f
      12'hBF: dout <= 8'b10011111; //  191 : 159 - 0x9f
      12'hC0: dout <= 8'b01111000; //  192 : 120 - 0x78 -- Background 0xc
      12'hC1: dout <= 8'b11111100; //  193 : 252 - 0xfc
      12'hC2: dout <= 8'b00011100; //  194 :  28 - 0x1c
      12'hC3: dout <= 8'b00111000; //  195 :  56 - 0x38
      12'hC4: dout <= 8'b00110000; //  196 :  48 - 0x30
      12'hC5: dout <= 8'b00000000; //  197 :   0 - 0x0
      12'hC6: dout <= 8'b01110000; //  198 : 112 - 0x70
      12'hC7: dout <= 8'b01110000; //  199 : 112 - 0x70
      12'hC8: dout <= 8'b10001111; //  200 : 143 - 0x8f -- plane 1
      12'hC9: dout <= 8'b00100111; //  201 :  39 - 0x27
      12'hCA: dout <= 8'b11100111; //  202 : 231 - 0xe7
      12'hCB: dout <= 8'b11001111; //  203 : 207 - 0xcf
      12'hCC: dout <= 8'b11011111; //  204 : 223 - 0xdf
      12'hCD: dout <= 8'b11111111; //  205 : 255 - 0xff
      12'hCE: dout <= 8'b10011111; //  206 : 159 - 0x9f
      12'hCF: dout <= 8'b10011111; //  207 : 159 - 0x9f
      12'hD0: dout <= 8'b00111100; //  208 :  60 - 0x3c -- Background 0xd
      12'hD1: dout <= 8'b01111110; //  209 : 126 - 0x7e
      12'hD2: dout <= 8'b11011011; //  210 : 219 - 0xdb
      12'hD3: dout <= 8'b11011111; //  211 : 223 - 0xdf
      12'hD4: dout <= 8'b11000011; //  212 : 195 - 0xc3
      12'hD5: dout <= 8'b01100110; //  213 : 102 - 0x66
      12'hD6: dout <= 8'b00111100; //  214 :  60 - 0x3c
      12'hD7: dout <= 8'b00000000; //  215 :   0 - 0x0
      12'hD8: dout <= 8'b11000111; //  216 : 199 - 0xc7 -- plane 1
      12'hD9: dout <= 8'b10101011; //  217 : 171 - 0xab
      12'hDA: dout <= 8'b01101101; //  218 : 109 - 0x6d
      12'hDB: dout <= 8'b01100101; //  219 : 101 - 0x65
      12'hDC: dout <= 8'b01111101; //  220 : 125 - 0x7d
      12'hDD: dout <= 8'b10111011; //  221 : 187 - 0xbb
      12'hDE: dout <= 8'b11000111; //  222 : 199 - 0xc7
      12'hDF: dout <= 8'b11111111; //  223 : 255 - 0xff
      12'hE0: dout <= 8'b00000000; //  224 :   0 - 0x0 -- Background 0xe
      12'hE1: dout <= 8'b00000000; //  225 :   0 - 0x0
      12'hE2: dout <= 8'b00000000; //  226 :   0 - 0x0
      12'hE3: dout <= 8'b00111100; //  227 :  60 - 0x3c
      12'hE4: dout <= 8'b00111110; //  228 :  62 - 0x3e
      12'hE5: dout <= 8'b00011110; //  229 :  30 - 0x1e
      12'hE6: dout <= 8'b00000000; //  230 :   0 - 0x0
      12'hE7: dout <= 8'b00000000; //  231 :   0 - 0x0
      12'hE8: dout <= 8'b11111111; //  232 : 255 - 0xff -- plane 1
      12'hE9: dout <= 8'b11111111; //  233 : 255 - 0xff
      12'hEA: dout <= 8'b11111111; //  234 : 255 - 0xff
      12'hEB: dout <= 8'b11000011; //  235 : 195 - 0xc3
      12'hEC: dout <= 8'b11000011; //  236 : 195 - 0xc3
      12'hED: dout <= 8'b11111111; //  237 : 255 - 0xff
      12'hEE: dout <= 8'b11111111; //  238 : 255 - 0xff
      12'hEF: dout <= 8'b11111111; //  239 : 255 - 0xff
      12'hF0: dout <= 8'b11111111; //  240 : 255 - 0xff -- Background 0xf
      12'hF1: dout <= 8'b11111111; //  241 : 255 - 0xff
      12'hF2: dout <= 8'b11111111; //  242 : 255 - 0xff
      12'hF3: dout <= 8'b11111111; //  243 : 255 - 0xff
      12'hF4: dout <= 8'b11111111; //  244 : 255 - 0xff
      12'hF5: dout <= 8'b11111111; //  245 : 255 - 0xff
      12'hF6: dout <= 8'b11100000; //  246 : 224 - 0xe0
      12'hF7: dout <= 8'b11100000; //  247 : 224 - 0xe0
      12'hF8: dout <= 8'b00000001; //  248 :   1 - 0x1 -- plane 1
      12'hF9: dout <= 8'b00101001; //  249 :  41 - 0x29
      12'hFA: dout <= 8'b01010101; //  250 :  85 - 0x55
      12'hFB: dout <= 8'b00101001; //  251 :  41 - 0x29
      12'hFC: dout <= 8'b01010101; //  252 :  85 - 0x55
      12'hFD: dout <= 8'b00000001; //  253 :   1 - 0x1
      12'hFE: dout <= 8'b00111111; //  254 :  63 - 0x3f
      12'hFF: dout <= 8'b00111111; //  255 :  63 - 0x3f
      12'h100: dout <= 8'b00001110; //  256 :  14 - 0xe -- Background 0x10
      12'h101: dout <= 8'b00001110; //  257 :  14 - 0xe
      12'h102: dout <= 8'b00011100; //  258 :  28 - 0x1c
      12'h103: dout <= 8'b00011100; //  259 :  28 - 0x1c
      12'h104: dout <= 8'b00011100; //  260 :  28 - 0x1c
      12'h105: dout <= 8'b00011100; //  261 :  28 - 0x1c
      12'h106: dout <= 8'b00111000; //  262 :  56 - 0x38
      12'h107: dout <= 8'b00111000; //  263 :  56 - 0x38
      12'h108: dout <= 8'b11110011; //  264 : 243 - 0xf3 -- plane 1
      12'h109: dout <= 8'b11110011; //  265 : 243 - 0xf3
      12'h10A: dout <= 8'b11100111; //  266 : 231 - 0xe7
      12'h10B: dout <= 8'b11100111; //  267 : 231 - 0xe7
      12'h10C: dout <= 8'b11100111; //  268 : 231 - 0xe7
      12'h10D: dout <= 8'b11100111; //  269 : 231 - 0xe7
      12'h10E: dout <= 8'b11001111; //  270 : 207 - 0xcf
      12'h10F: dout <= 8'b11001111; //  271 : 207 - 0xcf
      12'h110: dout <= 8'b00011100; //  272 :  28 - 0x1c -- Background 0x11
      12'h111: dout <= 8'b00111110; //  273 :  62 - 0x3e
      12'h112: dout <= 8'b01110111; //  274 : 119 - 0x77
      12'h113: dout <= 8'b01110111; //  275 : 119 - 0x77
      12'h114: dout <= 8'b01111111; //  276 : 127 - 0x7f
      12'h115: dout <= 8'b01111111; //  277 : 127 - 0x7f
      12'h116: dout <= 8'b01110111; //  278 : 119 - 0x77
      12'h117: dout <= 8'b01110111; //  279 : 119 - 0x77
      12'h118: dout <= 8'b11100111; //  280 : 231 - 0xe7 -- plane 1
      12'h119: dout <= 8'b11000011; //  281 : 195 - 0xc3
      12'h11A: dout <= 8'b10011001; //  282 : 153 - 0x99
      12'h11B: dout <= 8'b10011001; //  283 : 153 - 0x99
      12'h11C: dout <= 8'b10000001; //  284 : 129 - 0x81
      12'h11D: dout <= 8'b10000001; //  285 : 129 - 0x81
      12'h11E: dout <= 8'b10011001; //  286 : 153 - 0x99
      12'h11F: dout <= 8'b10011001; //  287 : 153 - 0x99
      12'h120: dout <= 8'b01111110; //  288 : 126 - 0x7e -- Background 0x12
      12'h121: dout <= 8'b01110111; //  289 : 119 - 0x77
      12'h122: dout <= 8'b01110111; //  290 : 119 - 0x77
      12'h123: dout <= 8'b01111110; //  291 : 126 - 0x7e
      12'h124: dout <= 8'b01111110; //  292 : 126 - 0x7e
      12'h125: dout <= 8'b01110111; //  293 : 119 - 0x77
      12'h126: dout <= 8'b01110111; //  294 : 119 - 0x77
      12'h127: dout <= 8'b01111110; //  295 : 126 - 0x7e
      12'h128: dout <= 8'b10000011; //  296 : 131 - 0x83 -- plane 1
      12'h129: dout <= 8'b10011001; //  297 : 153 - 0x99
      12'h12A: dout <= 8'b10011001; //  298 : 153 - 0x99
      12'h12B: dout <= 8'b10000011; //  299 : 131 - 0x83
      12'h12C: dout <= 8'b10000011; //  300 : 131 - 0x83
      12'h12D: dout <= 8'b10011001; //  301 : 153 - 0x99
      12'h12E: dout <= 8'b10011001; //  302 : 153 - 0x99
      12'h12F: dout <= 8'b10000011; //  303 : 131 - 0x83
      12'h130: dout <= 8'b00111110; //  304 :  62 - 0x3e -- Background 0x13
      12'h131: dout <= 8'b01111111; //  305 : 127 - 0x7f
      12'h132: dout <= 8'b01110111; //  306 : 119 - 0x77
      12'h133: dout <= 8'b01110000; //  307 : 112 - 0x70
      12'h134: dout <= 8'b01110000; //  308 : 112 - 0x70
      12'h135: dout <= 8'b01110111; //  309 : 119 - 0x77
      12'h136: dout <= 8'b01111111; //  310 : 127 - 0x7f
      12'h137: dout <= 8'b00111110; //  311 :  62 - 0x3e
      12'h138: dout <= 8'b11000011; //  312 : 195 - 0xc3 -- plane 1
      12'h139: dout <= 8'b10000001; //  313 : 129 - 0x81
      12'h13A: dout <= 8'b10011001; //  314 : 153 - 0x99
      12'h13B: dout <= 8'b10011111; //  315 : 159 - 0x9f
      12'h13C: dout <= 8'b10011111; //  316 : 159 - 0x9f
      12'h13D: dout <= 8'b10011001; //  317 : 153 - 0x99
      12'h13E: dout <= 8'b10000001; //  318 : 129 - 0x81
      12'h13F: dout <= 8'b11000011; //  319 : 195 - 0xc3
      12'h140: dout <= 8'b01111110; //  320 : 126 - 0x7e -- Background 0x14
      12'h141: dout <= 8'b01111111; //  321 : 127 - 0x7f
      12'h142: dout <= 8'b01110111; //  322 : 119 - 0x77
      12'h143: dout <= 8'b01110111; //  323 : 119 - 0x77
      12'h144: dout <= 8'b01110111; //  324 : 119 - 0x77
      12'h145: dout <= 8'b01110111; //  325 : 119 - 0x77
      12'h146: dout <= 8'b01111111; //  326 : 127 - 0x7f
      12'h147: dout <= 8'b01111110; //  327 : 126 - 0x7e
      12'h148: dout <= 8'b10000011; //  328 : 131 - 0x83 -- plane 1
      12'h149: dout <= 8'b10000001; //  329 : 129 - 0x81
      12'h14A: dout <= 8'b10011001; //  330 : 153 - 0x99
      12'h14B: dout <= 8'b10011001; //  331 : 153 - 0x99
      12'h14C: dout <= 8'b10011001; //  332 : 153 - 0x99
      12'h14D: dout <= 8'b10011001; //  333 : 153 - 0x99
      12'h14E: dout <= 8'b10000001; //  334 : 129 - 0x81
      12'h14F: dout <= 8'b10000011; //  335 : 131 - 0x83
      12'h150: dout <= 8'b01111111; //  336 : 127 - 0x7f -- Background 0x15
      12'h151: dout <= 8'b01111111; //  337 : 127 - 0x7f
      12'h152: dout <= 8'b01110000; //  338 : 112 - 0x70
      12'h153: dout <= 8'b01111100; //  339 : 124 - 0x7c
      12'h154: dout <= 8'b01111100; //  340 : 124 - 0x7c
      12'h155: dout <= 8'b01110000; //  341 : 112 - 0x70
      12'h156: dout <= 8'b01111111; //  342 : 127 - 0x7f
      12'h157: dout <= 8'b01111111; //  343 : 127 - 0x7f
      12'h158: dout <= 8'b10000001; //  344 : 129 - 0x81 -- plane 1
      12'h159: dout <= 8'b10000001; //  345 : 129 - 0x81
      12'h15A: dout <= 8'b10011111; //  346 : 159 - 0x9f
      12'h15B: dout <= 8'b10000111; //  347 : 135 - 0x87
      12'h15C: dout <= 8'b10000111; //  348 : 135 - 0x87
      12'h15D: dout <= 8'b10011111; //  349 : 159 - 0x9f
      12'h15E: dout <= 8'b10000001; //  350 : 129 - 0x81
      12'h15F: dout <= 8'b10000001; //  351 : 129 - 0x81
      12'h160: dout <= 8'b01111111; //  352 : 127 - 0x7f -- Background 0x16
      12'h161: dout <= 8'b01111111; //  353 : 127 - 0x7f
      12'h162: dout <= 8'b01110000; //  354 : 112 - 0x70
      12'h163: dout <= 8'b01111100; //  355 : 124 - 0x7c
      12'h164: dout <= 8'b01111100; //  356 : 124 - 0x7c
      12'h165: dout <= 8'b01110000; //  357 : 112 - 0x70
      12'h166: dout <= 8'b01110000; //  358 : 112 - 0x70
      12'h167: dout <= 8'b01110000; //  359 : 112 - 0x70
      12'h168: dout <= 8'b10000001; //  360 : 129 - 0x81 -- plane 1
      12'h169: dout <= 8'b10000001; //  361 : 129 - 0x81
      12'h16A: dout <= 8'b10011111; //  362 : 159 - 0x9f
      12'h16B: dout <= 8'b10000111; //  363 : 135 - 0x87
      12'h16C: dout <= 8'b10000111; //  364 : 135 - 0x87
      12'h16D: dout <= 8'b10011111; //  365 : 159 - 0x9f
      12'h16E: dout <= 8'b10011111; //  366 : 159 - 0x9f
      12'h16F: dout <= 8'b10011111; //  367 : 159 - 0x9f
      12'h170: dout <= 8'b00111110; //  368 :  62 - 0x3e -- Background 0x17
      12'h171: dout <= 8'b01111111; //  369 : 127 - 0x7f
      12'h172: dout <= 8'b01110111; //  370 : 119 - 0x77
      12'h173: dout <= 8'b01110000; //  371 : 112 - 0x70
      12'h174: dout <= 8'b01111111; //  372 : 127 - 0x7f
      12'h175: dout <= 8'b01110111; //  373 : 119 - 0x77
      12'h176: dout <= 8'b01111111; //  374 : 127 - 0x7f
      12'h177: dout <= 8'b00111110; //  375 :  62 - 0x3e
      12'h178: dout <= 8'b11000011; //  376 : 195 - 0xc3 -- plane 1
      12'h179: dout <= 8'b10000001; //  377 : 129 - 0x81
      12'h17A: dout <= 8'b10011001; //  378 : 153 - 0x99
      12'h17B: dout <= 8'b10011111; //  379 : 159 - 0x9f
      12'h17C: dout <= 8'b10010001; //  380 : 145 - 0x91
      12'h17D: dout <= 8'b10011001; //  381 : 153 - 0x99
      12'h17E: dout <= 8'b10000001; //  382 : 129 - 0x81
      12'h17F: dout <= 8'b11000011; //  383 : 195 - 0xc3
      12'h180: dout <= 8'b01110111; //  384 : 119 - 0x77 -- Background 0x18
      12'h181: dout <= 8'b01110111; //  385 : 119 - 0x77
      12'h182: dout <= 8'b01110111; //  386 : 119 - 0x77
      12'h183: dout <= 8'b01111111; //  387 : 127 - 0x7f
      12'h184: dout <= 8'b01111111; //  388 : 127 - 0x7f
      12'h185: dout <= 8'b01110111; //  389 : 119 - 0x77
      12'h186: dout <= 8'b01110111; //  390 : 119 - 0x77
      12'h187: dout <= 8'b01110111; //  391 : 119 - 0x77
      12'h188: dout <= 8'b10011001; //  392 : 153 - 0x99 -- plane 1
      12'h189: dout <= 8'b10011001; //  393 : 153 - 0x99
      12'h18A: dout <= 8'b10011001; //  394 : 153 - 0x99
      12'h18B: dout <= 8'b10000001; //  395 : 129 - 0x81
      12'h18C: dout <= 8'b10000001; //  396 : 129 - 0x81
      12'h18D: dout <= 8'b10011001; //  397 : 153 - 0x99
      12'h18E: dout <= 8'b10011001; //  398 : 153 - 0x99
      12'h18F: dout <= 8'b10011001; //  399 : 153 - 0x99
      12'h190: dout <= 8'b00111110; //  400 :  62 - 0x3e -- Background 0x19
      12'h191: dout <= 8'b00111110; //  401 :  62 - 0x3e
      12'h192: dout <= 8'b00011100; //  402 :  28 - 0x1c
      12'h193: dout <= 8'b00011100; //  403 :  28 - 0x1c
      12'h194: dout <= 8'b00011100; //  404 :  28 - 0x1c
      12'h195: dout <= 8'b00011100; //  405 :  28 - 0x1c
      12'h196: dout <= 8'b00111110; //  406 :  62 - 0x3e
      12'h197: dout <= 8'b00111110; //  407 :  62 - 0x3e
      12'h198: dout <= 8'b11000011; //  408 : 195 - 0xc3 -- plane 1
      12'h199: dout <= 8'b11000011; //  409 : 195 - 0xc3
      12'h19A: dout <= 8'b11100111; //  410 : 231 - 0xe7
      12'h19B: dout <= 8'b11100111; //  411 : 231 - 0xe7
      12'h19C: dout <= 8'b11100111; //  412 : 231 - 0xe7
      12'h19D: dout <= 8'b11100111; //  413 : 231 - 0xe7
      12'h19E: dout <= 8'b11000011; //  414 : 195 - 0xc3
      12'h19F: dout <= 8'b11000011; //  415 : 195 - 0xc3
      12'h1A0: dout <= 8'b00000111; //  416 :   7 - 0x7 -- Background 0x1a
      12'h1A1: dout <= 8'b00000111; //  417 :   7 - 0x7
      12'h1A2: dout <= 8'b00000111; //  418 :   7 - 0x7
      12'h1A3: dout <= 8'b00000111; //  419 :   7 - 0x7
      12'h1A4: dout <= 8'b00000111; //  420 :   7 - 0x7
      12'h1A5: dout <= 8'b01110111; //  421 : 119 - 0x77
      12'h1A6: dout <= 8'b01111111; //  422 : 127 - 0x7f
      12'h1A7: dout <= 8'b00111110; //  423 :  62 - 0x3e
      12'h1A8: dout <= 8'b11111001; //  424 : 249 - 0xf9 -- plane 1
      12'h1A9: dout <= 8'b11111001; //  425 : 249 - 0xf9
      12'h1AA: dout <= 8'b11111001; //  426 : 249 - 0xf9
      12'h1AB: dout <= 8'b11111001; //  427 : 249 - 0xf9
      12'h1AC: dout <= 8'b11111001; //  428 : 249 - 0xf9
      12'h1AD: dout <= 8'b10011001; //  429 : 153 - 0x99
      12'h1AE: dout <= 8'b10000001; //  430 : 129 - 0x81
      12'h1AF: dout <= 8'b11000011; //  431 : 195 - 0xc3
      12'h1B0: dout <= 8'b01110011; //  432 : 115 - 0x73 -- Background 0x1b
      12'h1B1: dout <= 8'b01110111; //  433 : 119 - 0x77
      12'h1B2: dout <= 8'b01111110; //  434 : 126 - 0x7e
      12'h1B3: dout <= 8'b01111100; //  435 : 124 - 0x7c
      12'h1B4: dout <= 8'b01111110; //  436 : 126 - 0x7e
      12'h1B5: dout <= 8'b01110111; //  437 : 119 - 0x77
      12'h1B6: dout <= 8'b01110111; //  438 : 119 - 0x77
      12'h1B7: dout <= 8'b01110111; //  439 : 119 - 0x77
      12'h1B8: dout <= 8'b10011101; //  440 : 157 - 0x9d -- plane 1
      12'h1B9: dout <= 8'b10011001; //  441 : 153 - 0x99
      12'h1BA: dout <= 8'b10010011; //  442 : 147 - 0x93
      12'h1BB: dout <= 8'b10000111; //  443 : 135 - 0x87
      12'h1BC: dout <= 8'b10000011; //  444 : 131 - 0x83
      12'h1BD: dout <= 8'b10011001; //  445 : 153 - 0x99
      12'h1BE: dout <= 8'b10011001; //  446 : 153 - 0x99
      12'h1BF: dout <= 8'b10011001; //  447 : 153 - 0x99
      12'h1C0: dout <= 8'b01110000; //  448 : 112 - 0x70 -- Background 0x1c
      12'h1C1: dout <= 8'b01110000; //  449 : 112 - 0x70
      12'h1C2: dout <= 8'b01110000; //  450 : 112 - 0x70
      12'h1C3: dout <= 8'b01110000; //  451 : 112 - 0x70
      12'h1C4: dout <= 8'b01110000; //  452 : 112 - 0x70
      12'h1C5: dout <= 8'b01110000; //  453 : 112 - 0x70
      12'h1C6: dout <= 8'b01111111; //  454 : 127 - 0x7f
      12'h1C7: dout <= 8'b01111111; //  455 : 127 - 0x7f
      12'h1C8: dout <= 8'b10011111; //  456 : 159 - 0x9f -- plane 1
      12'h1C9: dout <= 8'b10011111; //  457 : 159 - 0x9f
      12'h1CA: dout <= 8'b10011111; //  458 : 159 - 0x9f
      12'h1CB: dout <= 8'b10011111; //  459 : 159 - 0x9f
      12'h1CC: dout <= 8'b10011111; //  460 : 159 - 0x9f
      12'h1CD: dout <= 8'b10011111; //  461 : 159 - 0x9f
      12'h1CE: dout <= 8'b10000001; //  462 : 129 - 0x81
      12'h1CF: dout <= 8'b10000001; //  463 : 129 - 0x81
      12'h1D0: dout <= 8'b11100111; //  464 : 231 - 0xe7 -- Background 0x1d
      12'h1D1: dout <= 8'b11111111; //  465 : 255 - 0xff
      12'h1D2: dout <= 8'b11111111; //  466 : 255 - 0xff
      12'h1D3: dout <= 8'b11111111; //  467 : 255 - 0xff
      12'h1D4: dout <= 8'b11111111; //  468 : 255 - 0xff
      12'h1D5: dout <= 8'b11100111; //  469 : 231 - 0xe7
      12'h1D6: dout <= 8'b11100111; //  470 : 231 - 0xe7
      12'h1D7: dout <= 8'b11100111; //  471 : 231 - 0xe7
      12'h1D8: dout <= 8'b00111001; //  472 :  57 - 0x39 -- plane 1
      12'h1D9: dout <= 8'b00010001; //  473 :  17 - 0x11
      12'h1DA: dout <= 8'b00000001; //  474 :   1 - 0x1
      12'h1DB: dout <= 8'b00000001; //  475 :   1 - 0x1
      12'h1DC: dout <= 8'b00101001; //  476 :  41 - 0x29
      12'h1DD: dout <= 8'b00111001; //  477 :  57 - 0x39
      12'h1DE: dout <= 8'b00111001; //  478 :  57 - 0x39
      12'h1DF: dout <= 8'b00111001; //  479 :  57 - 0x39
      12'h1E0: dout <= 8'b01110111; //  480 : 119 - 0x77 -- Background 0x1e
      12'h1E1: dout <= 8'b01110111; //  481 : 119 - 0x77
      12'h1E2: dout <= 8'b01111111; //  482 : 127 - 0x7f
      12'h1E3: dout <= 8'b01111111; //  483 : 127 - 0x7f
      12'h1E4: dout <= 8'b01111111; //  484 : 127 - 0x7f
      12'h1E5: dout <= 8'b01111111; //  485 : 127 - 0x7f
      12'h1E6: dout <= 8'b01110111; //  486 : 119 - 0x77
      12'h1E7: dout <= 8'b01110111; //  487 : 119 - 0x77
      12'h1E8: dout <= 8'b10011001; //  488 : 153 - 0x99 -- plane 1
      12'h1E9: dout <= 8'b10011001; //  489 : 153 - 0x99
      12'h1EA: dout <= 8'b10001001; //  490 : 137 - 0x89
      12'h1EB: dout <= 8'b10000001; //  491 : 129 - 0x81
      12'h1EC: dout <= 8'b10000001; //  492 : 129 - 0x81
      12'h1ED: dout <= 8'b10010001; //  493 : 145 - 0x91
      12'h1EE: dout <= 8'b10011001; //  494 : 153 - 0x99
      12'h1EF: dout <= 8'b10011001; //  495 : 153 - 0x99
      12'h1F0: dout <= 8'b00111100; //  496 :  60 - 0x3c -- Background 0x1f
      12'h1F1: dout <= 8'b01111110; //  497 : 126 - 0x7e
      12'h1F2: dout <= 8'b11100111; //  498 : 231 - 0xe7
      12'h1F3: dout <= 8'b11100111; //  499 : 231 - 0xe7
      12'h1F4: dout <= 8'b11100111; //  500 : 231 - 0xe7
      12'h1F5: dout <= 8'b11100111; //  501 : 231 - 0xe7
      12'h1F6: dout <= 8'b01111110; //  502 : 126 - 0x7e
      12'h1F7: dout <= 8'b00111100; //  503 :  60 - 0x3c
      12'h1F8: dout <= 8'b11000111; //  504 : 199 - 0xc7 -- plane 1
      12'h1F9: dout <= 8'b10000011; //  505 : 131 - 0x83
      12'h1FA: dout <= 8'b00111001; //  506 :  57 - 0x39
      12'h1FB: dout <= 8'b00111001; //  507 :  57 - 0x39
      12'h1FC: dout <= 8'b00111001; //  508 :  57 - 0x39
      12'h1FD: dout <= 8'b00111001; //  509 :  57 - 0x39
      12'h1FE: dout <= 8'b10000011; //  510 : 131 - 0x83
      12'h1FF: dout <= 8'b11000111; //  511 : 199 - 0xc7
      12'h200: dout <= 8'b01111110; //  512 : 126 - 0x7e -- Background 0x20
      12'h201: dout <= 8'b01111111; //  513 : 127 - 0x7f
      12'h202: dout <= 8'b01110111; //  514 : 119 - 0x77
      12'h203: dout <= 8'b01110111; //  515 : 119 - 0x77
      12'h204: dout <= 8'b01111111; //  516 : 127 - 0x7f
      12'h205: dout <= 8'b01111110; //  517 : 126 - 0x7e
      12'h206: dout <= 8'b01110000; //  518 : 112 - 0x70
      12'h207: dout <= 8'b01110000; //  519 : 112 - 0x70
      12'h208: dout <= 8'b10000011; //  520 : 131 - 0x83 -- plane 1
      12'h209: dout <= 8'b10000001; //  521 : 129 - 0x81
      12'h20A: dout <= 8'b10011001; //  522 : 153 - 0x99
      12'h20B: dout <= 8'b10011001; //  523 : 153 - 0x99
      12'h20C: dout <= 8'b10000001; //  524 : 129 - 0x81
      12'h20D: dout <= 8'b10000011; //  525 : 131 - 0x83
      12'h20E: dout <= 8'b10011111; //  526 : 159 - 0x9f
      12'h20F: dout <= 8'b10011111; //  527 : 159 - 0x9f
      12'h210: dout <= 8'b00111100; //  528 :  60 - 0x3c -- Background 0x21
      12'h211: dout <= 8'b01111110; //  529 : 126 - 0x7e
      12'h212: dout <= 8'b11100111; //  530 : 231 - 0xe7
      12'h213: dout <= 8'b11100111; //  531 : 231 - 0xe7
      12'h214: dout <= 8'b11100111; //  532 : 231 - 0xe7
      12'h215: dout <= 8'b11101110; //  533 : 238 - 0xee
      12'h216: dout <= 8'b01111111; //  534 : 127 - 0x7f
      12'h217: dout <= 8'b00111111; //  535 :  63 - 0x3f
      12'h218: dout <= 8'b11000111; //  536 : 199 - 0xc7 -- plane 1
      12'h219: dout <= 8'b10000011; //  537 : 131 - 0x83
      12'h21A: dout <= 8'b00111001; //  538 :  57 - 0x39
      12'h21B: dout <= 8'b00111001; //  539 :  57 - 0x39
      12'h21C: dout <= 8'b00111001; //  540 :  57 - 0x39
      12'h21D: dout <= 8'b00110011; //  541 :  51 - 0x33
      12'h21E: dout <= 8'b10000001; //  542 : 129 - 0x81
      12'h21F: dout <= 8'b11001001; //  543 : 201 - 0xc9
      12'h220: dout <= 8'b01111110; //  544 : 126 - 0x7e -- Background 0x22
      12'h221: dout <= 8'b01111111; //  545 : 127 - 0x7f
      12'h222: dout <= 8'b01110111; //  546 : 119 - 0x77
      12'h223: dout <= 8'b01110111; //  547 : 119 - 0x77
      12'h224: dout <= 8'b01111111; //  548 : 127 - 0x7f
      12'h225: dout <= 8'b01111110; //  549 : 126 - 0x7e
      12'h226: dout <= 8'b01110111; //  550 : 119 - 0x77
      12'h227: dout <= 8'b01110111; //  551 : 119 - 0x77
      12'h228: dout <= 8'b10000011; //  552 : 131 - 0x83 -- plane 1
      12'h229: dout <= 8'b10000001; //  553 : 129 - 0x81
      12'h22A: dout <= 8'b10011001; //  554 : 153 - 0x99
      12'h22B: dout <= 8'b10011001; //  555 : 153 - 0x99
      12'h22C: dout <= 8'b10000001; //  556 : 129 - 0x81
      12'h22D: dout <= 8'b10000011; //  557 : 131 - 0x83
      12'h22E: dout <= 8'b10011001; //  558 : 153 - 0x99
      12'h22F: dout <= 8'b10011001; //  559 : 153 - 0x99
      12'h230: dout <= 8'b00111110; //  560 :  62 - 0x3e -- Background 0x23
      12'h231: dout <= 8'b01111111; //  561 : 127 - 0x7f
      12'h232: dout <= 8'b01110000; //  562 : 112 - 0x70
      12'h233: dout <= 8'b01111110; //  563 : 126 - 0x7e
      12'h234: dout <= 8'b00111111; //  564 :  63 - 0x3f
      12'h235: dout <= 8'b00000111; //  565 :   7 - 0x7
      12'h236: dout <= 8'b01111111; //  566 : 127 - 0x7f
      12'h237: dout <= 8'b00111110; //  567 :  62 - 0x3e
      12'h238: dout <= 8'b11000011; //  568 : 195 - 0xc3 -- plane 1
      12'h239: dout <= 8'b10000001; //  569 : 129 - 0x81
      12'h23A: dout <= 8'b10011111; //  570 : 159 - 0x9f
      12'h23B: dout <= 8'b10000011; //  571 : 131 - 0x83
      12'h23C: dout <= 8'b11000001; //  572 : 193 - 0xc1
      12'h23D: dout <= 8'b11111001; //  573 : 249 - 0xf9
      12'h23E: dout <= 8'b10000001; //  574 : 129 - 0x81
      12'h23F: dout <= 8'b11000011; //  575 : 195 - 0xc3
      12'h240: dout <= 8'b01111111; //  576 : 127 - 0x7f -- Background 0x24
      12'h241: dout <= 8'b01111111; //  577 : 127 - 0x7f
      12'h242: dout <= 8'b00011100; //  578 :  28 - 0x1c
      12'h243: dout <= 8'b00011100; //  579 :  28 - 0x1c
      12'h244: dout <= 8'b00011100; //  580 :  28 - 0x1c
      12'h245: dout <= 8'b00011100; //  581 :  28 - 0x1c
      12'h246: dout <= 8'b00011100; //  582 :  28 - 0x1c
      12'h247: dout <= 8'b00011100; //  583 :  28 - 0x1c
      12'h248: dout <= 8'b10000001; //  584 : 129 - 0x81 -- plane 1
      12'h249: dout <= 8'b10000001; //  585 : 129 - 0x81
      12'h24A: dout <= 8'b11100111; //  586 : 231 - 0xe7
      12'h24B: dout <= 8'b11100111; //  587 : 231 - 0xe7
      12'h24C: dout <= 8'b11100111; //  588 : 231 - 0xe7
      12'h24D: dout <= 8'b11100111; //  589 : 231 - 0xe7
      12'h24E: dout <= 8'b11100111; //  590 : 231 - 0xe7
      12'h24F: dout <= 8'b11100111; //  591 : 231 - 0xe7
      12'h250: dout <= 8'b01110111; //  592 : 119 - 0x77 -- Background 0x25
      12'h251: dout <= 8'b01110111; //  593 : 119 - 0x77
      12'h252: dout <= 8'b01110111; //  594 : 119 - 0x77
      12'h253: dout <= 8'b01110111; //  595 : 119 - 0x77
      12'h254: dout <= 8'b01110111; //  596 : 119 - 0x77
      12'h255: dout <= 8'b01110111; //  597 : 119 - 0x77
      12'h256: dout <= 8'b01111111; //  598 : 127 - 0x7f
      12'h257: dout <= 8'b00111110; //  599 :  62 - 0x3e
      12'h258: dout <= 8'b10011001; //  600 : 153 - 0x99 -- plane 1
      12'h259: dout <= 8'b10011001; //  601 : 153 - 0x99
      12'h25A: dout <= 8'b10011001; //  602 : 153 - 0x99
      12'h25B: dout <= 8'b10011001; //  603 : 153 - 0x99
      12'h25C: dout <= 8'b10011001; //  604 : 153 - 0x99
      12'h25D: dout <= 8'b10011001; //  605 : 153 - 0x99
      12'h25E: dout <= 8'b10000001; //  606 : 129 - 0x81
      12'h25F: dout <= 8'b11000011; //  607 : 195 - 0xc3
      12'h260: dout <= 8'b01110111; //  608 : 119 - 0x77 -- Background 0x26
      12'h261: dout <= 8'b01110111; //  609 : 119 - 0x77
      12'h262: dout <= 8'b01110111; //  610 : 119 - 0x77
      12'h263: dout <= 8'b01110111; //  611 : 119 - 0x77
      12'h264: dout <= 8'b01110111; //  612 : 119 - 0x77
      12'h265: dout <= 8'b01110111; //  613 : 119 - 0x77
      12'h266: dout <= 8'b00111110; //  614 :  62 - 0x3e
      12'h267: dout <= 8'b00011100; //  615 :  28 - 0x1c
      12'h268: dout <= 8'b10011001; //  616 : 153 - 0x99 -- plane 1
      12'h269: dout <= 8'b10011001; //  617 : 153 - 0x99
      12'h26A: dout <= 8'b10011001; //  618 : 153 - 0x99
      12'h26B: dout <= 8'b10011001; //  619 : 153 - 0x99
      12'h26C: dout <= 8'b10011001; //  620 : 153 - 0x99
      12'h26D: dout <= 8'b10011001; //  621 : 153 - 0x99
      12'h26E: dout <= 8'b11000011; //  622 : 195 - 0xc3
      12'h26F: dout <= 8'b11100111; //  623 : 231 - 0xe7
      12'h270: dout <= 8'b11100111; //  624 : 231 - 0xe7 -- Background 0x27
      12'h271: dout <= 8'b11100111; //  625 : 231 - 0xe7
      12'h272: dout <= 8'b11100111; //  626 : 231 - 0xe7
      12'h273: dout <= 8'b11100111; //  627 : 231 - 0xe7
      12'h274: dout <= 8'b11110111; //  628 : 247 - 0xf7
      12'h275: dout <= 8'b11111111; //  629 : 255 - 0xff
      12'h276: dout <= 8'b11111111; //  630 : 255 - 0xff
      12'h277: dout <= 8'b01111110; //  631 : 126 - 0x7e
      12'h278: dout <= 8'b00111001; //  632 :  57 - 0x39 -- plane 1
      12'h279: dout <= 8'b00111001; //  633 :  57 - 0x39
      12'h27A: dout <= 8'b00111001; //  634 :  57 - 0x39
      12'h27B: dout <= 8'b00111001; //  635 :  57 - 0x39
      12'h27C: dout <= 8'b00101001; //  636 :  41 - 0x29
      12'h27D: dout <= 8'b00000001; //  637 :   1 - 0x1
      12'h27E: dout <= 8'b00000001; //  638 :   1 - 0x1
      12'h27F: dout <= 8'b10010011; //  639 : 147 - 0x93
      12'h280: dout <= 8'b01110111; //  640 : 119 - 0x77 -- Background 0x28
      12'h281: dout <= 8'b01110111; //  641 : 119 - 0x77
      12'h282: dout <= 8'b01110111; //  642 : 119 - 0x77
      12'h283: dout <= 8'b00111110; //  643 :  62 - 0x3e
      12'h284: dout <= 8'b00111110; //  644 :  62 - 0x3e
      12'h285: dout <= 8'b01110111; //  645 : 119 - 0x77
      12'h286: dout <= 8'b01110111; //  646 : 119 - 0x77
      12'h287: dout <= 8'b01110111; //  647 : 119 - 0x77
      12'h288: dout <= 8'b10011001; //  648 : 153 - 0x99 -- plane 1
      12'h289: dout <= 8'b10011001; //  649 : 153 - 0x99
      12'h28A: dout <= 8'b10011001; //  650 : 153 - 0x99
      12'h28B: dout <= 8'b11000011; //  651 : 195 - 0xc3
      12'h28C: dout <= 8'b11000011; //  652 : 195 - 0xc3
      12'h28D: dout <= 8'b10011001; //  653 : 153 - 0x99
      12'h28E: dout <= 8'b10011001; //  654 : 153 - 0x99
      12'h28F: dout <= 8'b10011001; //  655 : 153 - 0x99
      12'h290: dout <= 8'b01110111; //  656 : 119 - 0x77 -- Background 0x29
      12'h291: dout <= 8'b01110111; //  657 : 119 - 0x77
      12'h292: dout <= 8'b01110111; //  658 : 119 - 0x77
      12'h293: dout <= 8'b01111111; //  659 : 127 - 0x7f
      12'h294: dout <= 8'b00111110; //  660 :  62 - 0x3e
      12'h295: dout <= 8'b00011100; //  661 :  28 - 0x1c
      12'h296: dout <= 8'b00011100; //  662 :  28 - 0x1c
      12'h297: dout <= 8'b00011100; //  663 :  28 - 0x1c
      12'h298: dout <= 8'b10011001; //  664 : 153 - 0x99 -- plane 1
      12'h299: dout <= 8'b10011001; //  665 : 153 - 0x99
      12'h29A: dout <= 8'b10011001; //  666 : 153 - 0x99
      12'h29B: dout <= 8'b10000001; //  667 : 129 - 0x81
      12'h29C: dout <= 8'b11000011; //  668 : 195 - 0xc3
      12'h29D: dout <= 8'b11100111; //  669 : 231 - 0xe7
      12'h29E: dout <= 8'b11100111; //  670 : 231 - 0xe7
      12'h29F: dout <= 8'b11100111; //  671 : 231 - 0xe7
      12'h2A0: dout <= 8'b01111111; //  672 : 127 - 0x7f -- Background 0x2a
      12'h2A1: dout <= 8'b01111111; //  673 : 127 - 0x7f
      12'h2A2: dout <= 8'b00001110; //  674 :  14 - 0xe
      12'h2A3: dout <= 8'b00011100; //  675 :  28 - 0x1c
      12'h2A4: dout <= 8'b00011100; //  676 :  28 - 0x1c
      12'h2A5: dout <= 8'b00111000; //  677 :  56 - 0x38
      12'h2A6: dout <= 8'b01111111; //  678 : 127 - 0x7f
      12'h2A7: dout <= 8'b01111111; //  679 : 127 - 0x7f
      12'h2A8: dout <= 8'b10000001; //  680 : 129 - 0x81 -- plane 1
      12'h2A9: dout <= 8'b10000001; //  681 : 129 - 0x81
      12'h2AA: dout <= 8'b11110011; //  682 : 243 - 0xf3
      12'h2AB: dout <= 8'b11100111; //  683 : 231 - 0xe7
      12'h2AC: dout <= 8'b11100111; //  684 : 231 - 0xe7
      12'h2AD: dout <= 8'b11001111; //  685 : 207 - 0xcf
      12'h2AE: dout <= 8'b10000001; //  686 : 129 - 0x81
      12'h2AF: dout <= 8'b10000001; //  687 : 129 - 0x81
      12'h2B0: dout <= 8'b00111110; //  688 :  62 - 0x3e -- Background 0x2b
      12'h2B1: dout <= 8'b01100011; //  689 :  99 - 0x63
      12'h2B2: dout <= 8'b01101111; //  690 : 111 - 0x6f
      12'h2B3: dout <= 8'b01111111; //  691 : 127 - 0x7f
      12'h2B4: dout <= 8'b01111111; //  692 : 127 - 0x7f
      12'h2B5: dout <= 8'b01111110; //  693 : 126 - 0x7e
      12'h2B6: dout <= 8'b01100000; //  694 :  96 - 0x60
      12'h2B7: dout <= 8'b00111111; //  695 :  63 - 0x3f
      12'h2B8: dout <= 8'b11000011; //  696 : 195 - 0xc3 -- plane 1
      12'h2B9: dout <= 8'b10111101; //  697 : 189 - 0xbd
      12'h2BA: dout <= 8'b10110101; //  698 : 181 - 0xb5
      12'h2BB: dout <= 8'b10101001; //  699 : 169 - 0xa9
      12'h2BC: dout <= 8'b10101001; //  700 : 169 - 0xa9
      12'h2BD: dout <= 8'b10100011; //  701 : 163 - 0xa3
      12'h2BE: dout <= 8'b10111111; //  702 : 191 - 0xbf
      12'h2BF: dout <= 8'b11000001; //  703 : 193 - 0xc1
      12'h2C0: dout <= 8'b00000000; //  704 :   0 - 0x0 -- Background 0x2c
      12'h2C1: dout <= 8'b01110000; //  705 : 112 - 0x70
      12'h2C2: dout <= 8'b01111100; //  706 : 124 - 0x7c
      12'h2C3: dout <= 8'b01111111; //  707 : 127 - 0x7f
      12'h2C4: dout <= 8'b01111111; //  708 : 127 - 0x7f
      12'h2C5: dout <= 8'b01111100; //  709 : 124 - 0x7c
      12'h2C6: dout <= 8'b01110000; //  710 : 112 - 0x70
      12'h2C7: dout <= 8'b00000000; //  711 :   0 - 0x0
      12'h2C8: dout <= 8'b11111111; //  712 : 255 - 0xff -- plane 1
      12'h2C9: dout <= 8'b10011111; //  713 : 159 - 0x9f
      12'h2CA: dout <= 8'b10000111; //  714 : 135 - 0x87
      12'h2CB: dout <= 8'b10000001; //  715 : 129 - 0x81
      12'h2CC: dout <= 8'b10000001; //  716 : 129 - 0x81
      12'h2CD: dout <= 8'b10000111; //  717 : 135 - 0x87
      12'h2CE: dout <= 8'b10011111; //  718 : 159 - 0x9f
      12'h2CF: dout <= 8'b11111111; //  719 : 255 - 0xff
      12'h2D0: dout <= 8'b00000000; //  720 :   0 - 0x0 -- Background 0x2d
      12'h2D1: dout <= 8'b01110000; //  721 : 112 - 0x70
      12'h2D2: dout <= 8'b01110000; //  722 : 112 - 0x70
      12'h2D3: dout <= 8'b00000000; //  723 :   0 - 0x0
      12'h2D4: dout <= 8'b00000000; //  724 :   0 - 0x0
      12'h2D5: dout <= 8'b01110000; //  725 : 112 - 0x70
      12'h2D6: dout <= 8'b01110000; //  726 : 112 - 0x70
      12'h2D7: dout <= 8'b00000000; //  727 :   0 - 0x0
      12'h2D8: dout <= 8'b11111111; //  728 : 255 - 0xff -- plane 1
      12'h2D9: dout <= 8'b10011111; //  729 : 159 - 0x9f
      12'h2DA: dout <= 8'b10011111; //  730 : 159 - 0x9f
      12'h2DB: dout <= 8'b11111111; //  731 : 255 - 0xff
      12'h2DC: dout <= 8'b11111111; //  732 : 255 - 0xff
      12'h2DD: dout <= 8'b10011111; //  733 : 159 - 0x9f
      12'h2DE: dout <= 8'b10011111; //  734 : 159 - 0x9f
      12'h2DF: dout <= 8'b11111111; //  735 : 255 - 0xff
      12'h2E0: dout <= 8'b00000000; //  736 :   0 - 0x0 -- Background 0x2e
      12'h2E1: dout <= 8'b00000000; //  737 :   0 - 0x0
      12'h2E2: dout <= 8'b00000000; //  738 :   0 - 0x0
      12'h2E3: dout <= 8'b00000000; //  739 :   0 - 0x0
      12'h2E4: dout <= 8'b00000000; //  740 :   0 - 0x0
      12'h2E5: dout <= 8'b00000000; //  741 :   0 - 0x0
      12'h2E6: dout <= 8'b00000000; //  742 :   0 - 0x0
      12'h2E7: dout <= 8'b00000000; //  743 :   0 - 0x0
      12'h2E8: dout <= 8'b00000000; //  744 :   0 - 0x0 -- plane 1
      12'h2E9: dout <= 8'b00000000; //  745 :   0 - 0x0
      12'h2EA: dout <= 8'b00000000; //  746 :   0 - 0x0
      12'h2EB: dout <= 8'b00000000; //  747 :   0 - 0x0
      12'h2EC: dout <= 8'b00000000; //  748 :   0 - 0x0
      12'h2ED: dout <= 8'b00000000; //  749 :   0 - 0x0
      12'h2EE: dout <= 8'b00000000; //  750 :   0 - 0x0
      12'h2EF: dout <= 8'b00000000; //  751 :   0 - 0x0
      12'h2F0: dout <= 8'b00000000; //  752 :   0 - 0x0 -- Background 0x2f
      12'h2F1: dout <= 8'b00000000; //  753 :   0 - 0x0
      12'h2F2: dout <= 8'b00000000; //  754 :   0 - 0x0
      12'h2F3: dout <= 8'b00000000; //  755 :   0 - 0x0
      12'h2F4: dout <= 8'b00000000; //  756 :   0 - 0x0
      12'h2F5: dout <= 8'b00000000; //  757 :   0 - 0x0
      12'h2F6: dout <= 8'b00000000; //  758 :   0 - 0x0
      12'h2F7: dout <= 8'b00000000; //  759 :   0 - 0x0
      12'h2F8: dout <= 8'b00000000; //  760 :   0 - 0x0 -- plane 1
      12'h2F9: dout <= 8'b00000000; //  761 :   0 - 0x0
      12'h2FA: dout <= 8'b00000000; //  762 :   0 - 0x0
      12'h2FB: dout <= 8'b00000000; //  763 :   0 - 0x0
      12'h2FC: dout <= 8'b00000000; //  764 :   0 - 0x0
      12'h2FD: dout <= 8'b00000000; //  765 :   0 - 0x0
      12'h2FE: dout <= 8'b00000000; //  766 :   0 - 0x0
      12'h2FF: dout <= 8'b00000000; //  767 :   0 - 0x0
      12'h300: dout <= 8'b00000000; //  768 :   0 - 0x0 -- Background 0x30
      12'h301: dout <= 8'b00000000; //  769 :   0 - 0x0
      12'h302: dout <= 8'b00000000; //  770 :   0 - 0x0
      12'h303: dout <= 8'b00000000; //  771 :   0 - 0x0
      12'h304: dout <= 8'b00000000; //  772 :   0 - 0x0
      12'h305: dout <= 8'b00000000; //  773 :   0 - 0x0
      12'h306: dout <= 8'b00000000; //  774 :   0 - 0x0
      12'h307: dout <= 8'b00000000; //  775 :   0 - 0x0
      12'h308: dout <= 8'b00000000; //  776 :   0 - 0x0 -- plane 1
      12'h309: dout <= 8'b00000000; //  777 :   0 - 0x0
      12'h30A: dout <= 8'b00000000; //  778 :   0 - 0x0
      12'h30B: dout <= 8'b00000000; //  779 :   0 - 0x0
      12'h30C: dout <= 8'b00000000; //  780 :   0 - 0x0
      12'h30D: dout <= 8'b00000000; //  781 :   0 - 0x0
      12'h30E: dout <= 8'b00000000; //  782 :   0 - 0x0
      12'h30F: dout <= 8'b00000000; //  783 :   0 - 0x0
      12'h310: dout <= 8'b00000000; //  784 :   0 - 0x0 -- Background 0x31
      12'h311: dout <= 8'b00000000; //  785 :   0 - 0x0
      12'h312: dout <= 8'b00000000; //  786 :   0 - 0x0
      12'h313: dout <= 8'b00000000; //  787 :   0 - 0x0
      12'h314: dout <= 8'b00000000; //  788 :   0 - 0x0
      12'h315: dout <= 8'b00000000; //  789 :   0 - 0x0
      12'h316: dout <= 8'b00000000; //  790 :   0 - 0x0
      12'h317: dout <= 8'b00000000; //  791 :   0 - 0x0
      12'h318: dout <= 8'b00000000; //  792 :   0 - 0x0 -- plane 1
      12'h319: dout <= 8'b00000000; //  793 :   0 - 0x0
      12'h31A: dout <= 8'b00000000; //  794 :   0 - 0x0
      12'h31B: dout <= 8'b00000000; //  795 :   0 - 0x0
      12'h31C: dout <= 8'b00000000; //  796 :   0 - 0x0
      12'h31D: dout <= 8'b00000000; //  797 :   0 - 0x0
      12'h31E: dout <= 8'b00000000; //  798 :   0 - 0x0
      12'h31F: dout <= 8'b00000000; //  799 :   0 - 0x0
      12'h320: dout <= 8'b00000000; //  800 :   0 - 0x0 -- Background 0x32
      12'h321: dout <= 8'b00000000; //  801 :   0 - 0x0
      12'h322: dout <= 8'b00000000; //  802 :   0 - 0x0
      12'h323: dout <= 8'b00000000; //  803 :   0 - 0x0
      12'h324: dout <= 8'b00000000; //  804 :   0 - 0x0
      12'h325: dout <= 8'b00000000; //  805 :   0 - 0x0
      12'h326: dout <= 8'b00000000; //  806 :   0 - 0x0
      12'h327: dout <= 8'b00000000; //  807 :   0 - 0x0
      12'h328: dout <= 8'b00000000; //  808 :   0 - 0x0 -- plane 1
      12'h329: dout <= 8'b00000000; //  809 :   0 - 0x0
      12'h32A: dout <= 8'b00000000; //  810 :   0 - 0x0
      12'h32B: dout <= 8'b00000000; //  811 :   0 - 0x0
      12'h32C: dout <= 8'b00000000; //  812 :   0 - 0x0
      12'h32D: dout <= 8'b00000000; //  813 :   0 - 0x0
      12'h32E: dout <= 8'b00000000; //  814 :   0 - 0x0
      12'h32F: dout <= 8'b00000000; //  815 :   0 - 0x0
      12'h330: dout <= 8'b00000000; //  816 :   0 - 0x0 -- Background 0x33
      12'h331: dout <= 8'b00000000; //  817 :   0 - 0x0
      12'h332: dout <= 8'b00000000; //  818 :   0 - 0x0
      12'h333: dout <= 8'b00000000; //  819 :   0 - 0x0
      12'h334: dout <= 8'b00000000; //  820 :   0 - 0x0
      12'h335: dout <= 8'b00000000; //  821 :   0 - 0x0
      12'h336: dout <= 8'b00000000; //  822 :   0 - 0x0
      12'h337: dout <= 8'b00000000; //  823 :   0 - 0x0
      12'h338: dout <= 8'b00000000; //  824 :   0 - 0x0 -- plane 1
      12'h339: dout <= 8'b00000000; //  825 :   0 - 0x0
      12'h33A: dout <= 8'b00000000; //  826 :   0 - 0x0
      12'h33B: dout <= 8'b00000000; //  827 :   0 - 0x0
      12'h33C: dout <= 8'b00000000; //  828 :   0 - 0x0
      12'h33D: dout <= 8'b00000000; //  829 :   0 - 0x0
      12'h33E: dout <= 8'b00000000; //  830 :   0 - 0x0
      12'h33F: dout <= 8'b00000000; //  831 :   0 - 0x0
      12'h340: dout <= 8'b00000000; //  832 :   0 - 0x0 -- Background 0x34
      12'h341: dout <= 8'b00000000; //  833 :   0 - 0x0
      12'h342: dout <= 8'b00000000; //  834 :   0 - 0x0
      12'h343: dout <= 8'b00000000; //  835 :   0 - 0x0
      12'h344: dout <= 8'b00000000; //  836 :   0 - 0x0
      12'h345: dout <= 8'b00000000; //  837 :   0 - 0x0
      12'h346: dout <= 8'b00000000; //  838 :   0 - 0x0
      12'h347: dout <= 8'b00000000; //  839 :   0 - 0x0
      12'h348: dout <= 8'b00000000; //  840 :   0 - 0x0 -- plane 1
      12'h349: dout <= 8'b00000000; //  841 :   0 - 0x0
      12'h34A: dout <= 8'b00000000; //  842 :   0 - 0x0
      12'h34B: dout <= 8'b00000000; //  843 :   0 - 0x0
      12'h34C: dout <= 8'b00000000; //  844 :   0 - 0x0
      12'h34D: dout <= 8'b00000000; //  845 :   0 - 0x0
      12'h34E: dout <= 8'b00000000; //  846 :   0 - 0x0
      12'h34F: dout <= 8'b00000000; //  847 :   0 - 0x0
      12'h350: dout <= 8'b00000000; //  848 :   0 - 0x0 -- Background 0x35
      12'h351: dout <= 8'b00000000; //  849 :   0 - 0x0
      12'h352: dout <= 8'b00000000; //  850 :   0 - 0x0
      12'h353: dout <= 8'b00000000; //  851 :   0 - 0x0
      12'h354: dout <= 8'b00000000; //  852 :   0 - 0x0
      12'h355: dout <= 8'b00000000; //  853 :   0 - 0x0
      12'h356: dout <= 8'b00000000; //  854 :   0 - 0x0
      12'h357: dout <= 8'b00000000; //  855 :   0 - 0x0
      12'h358: dout <= 8'b00000000; //  856 :   0 - 0x0 -- plane 1
      12'h359: dout <= 8'b00000000; //  857 :   0 - 0x0
      12'h35A: dout <= 8'b00000000; //  858 :   0 - 0x0
      12'h35B: dout <= 8'b00000000; //  859 :   0 - 0x0
      12'h35C: dout <= 8'b00000000; //  860 :   0 - 0x0
      12'h35D: dout <= 8'b00000000; //  861 :   0 - 0x0
      12'h35E: dout <= 8'b00000000; //  862 :   0 - 0x0
      12'h35F: dout <= 8'b00000000; //  863 :   0 - 0x0
      12'h360: dout <= 8'b00000000; //  864 :   0 - 0x0 -- Background 0x36
      12'h361: dout <= 8'b00000000; //  865 :   0 - 0x0
      12'h362: dout <= 8'b00000000; //  866 :   0 - 0x0
      12'h363: dout <= 8'b00000000; //  867 :   0 - 0x0
      12'h364: dout <= 8'b00000000; //  868 :   0 - 0x0
      12'h365: dout <= 8'b00000000; //  869 :   0 - 0x0
      12'h366: dout <= 8'b00000000; //  870 :   0 - 0x0
      12'h367: dout <= 8'b00000000; //  871 :   0 - 0x0
      12'h368: dout <= 8'b00000000; //  872 :   0 - 0x0 -- plane 1
      12'h369: dout <= 8'b00000000; //  873 :   0 - 0x0
      12'h36A: dout <= 8'b00000000; //  874 :   0 - 0x0
      12'h36B: dout <= 8'b00000000; //  875 :   0 - 0x0
      12'h36C: dout <= 8'b00000000; //  876 :   0 - 0x0
      12'h36D: dout <= 8'b00000000; //  877 :   0 - 0x0
      12'h36E: dout <= 8'b00000000; //  878 :   0 - 0x0
      12'h36F: dout <= 8'b00000000; //  879 :   0 - 0x0
      12'h370: dout <= 8'b00000000; //  880 :   0 - 0x0 -- Background 0x37
      12'h371: dout <= 8'b00000000; //  881 :   0 - 0x0
      12'h372: dout <= 8'b00000000; //  882 :   0 - 0x0
      12'h373: dout <= 8'b00000000; //  883 :   0 - 0x0
      12'h374: dout <= 8'b00000000; //  884 :   0 - 0x0
      12'h375: dout <= 8'b00000000; //  885 :   0 - 0x0
      12'h376: dout <= 8'b00000000; //  886 :   0 - 0x0
      12'h377: dout <= 8'b00000000; //  887 :   0 - 0x0
      12'h378: dout <= 8'b00000000; //  888 :   0 - 0x0 -- plane 1
      12'h379: dout <= 8'b00000000; //  889 :   0 - 0x0
      12'h37A: dout <= 8'b00000000; //  890 :   0 - 0x0
      12'h37B: dout <= 8'b00000000; //  891 :   0 - 0x0
      12'h37C: dout <= 8'b00000000; //  892 :   0 - 0x0
      12'h37D: dout <= 8'b00000000; //  893 :   0 - 0x0
      12'h37E: dout <= 8'b00000000; //  894 :   0 - 0x0
      12'h37F: dout <= 8'b00000000; //  895 :   0 - 0x0
      12'h380: dout <= 8'b00000000; //  896 :   0 - 0x0 -- Background 0x38
      12'h381: dout <= 8'b00000000; //  897 :   0 - 0x0
      12'h382: dout <= 8'b00000000; //  898 :   0 - 0x0
      12'h383: dout <= 8'b00000000; //  899 :   0 - 0x0
      12'h384: dout <= 8'b00000000; //  900 :   0 - 0x0
      12'h385: dout <= 8'b00000000; //  901 :   0 - 0x0
      12'h386: dout <= 8'b00000000; //  902 :   0 - 0x0
      12'h387: dout <= 8'b00000000; //  903 :   0 - 0x0
      12'h388: dout <= 8'b00000000; //  904 :   0 - 0x0 -- plane 1
      12'h389: dout <= 8'b00000000; //  905 :   0 - 0x0
      12'h38A: dout <= 8'b00000000; //  906 :   0 - 0x0
      12'h38B: dout <= 8'b00000000; //  907 :   0 - 0x0
      12'h38C: dout <= 8'b00000000; //  908 :   0 - 0x0
      12'h38D: dout <= 8'b00000000; //  909 :   0 - 0x0
      12'h38E: dout <= 8'b00000000; //  910 :   0 - 0x0
      12'h38F: dout <= 8'b00000000; //  911 :   0 - 0x0
      12'h390: dout <= 8'b00000000; //  912 :   0 - 0x0 -- Background 0x39
      12'h391: dout <= 8'b00000000; //  913 :   0 - 0x0
      12'h392: dout <= 8'b00000000; //  914 :   0 - 0x0
      12'h393: dout <= 8'b00000000; //  915 :   0 - 0x0
      12'h394: dout <= 8'b00000000; //  916 :   0 - 0x0
      12'h395: dout <= 8'b00000000; //  917 :   0 - 0x0
      12'h396: dout <= 8'b00000000; //  918 :   0 - 0x0
      12'h397: dout <= 8'b00000000; //  919 :   0 - 0x0
      12'h398: dout <= 8'b00000000; //  920 :   0 - 0x0 -- plane 1
      12'h399: dout <= 8'b00000000; //  921 :   0 - 0x0
      12'h39A: dout <= 8'b00000000; //  922 :   0 - 0x0
      12'h39B: dout <= 8'b00000000; //  923 :   0 - 0x0
      12'h39C: dout <= 8'b00000000; //  924 :   0 - 0x0
      12'h39D: dout <= 8'b00000000; //  925 :   0 - 0x0
      12'h39E: dout <= 8'b00000000; //  926 :   0 - 0x0
      12'h39F: dout <= 8'b00000000; //  927 :   0 - 0x0
      12'h3A0: dout <= 8'b00000000; //  928 :   0 - 0x0 -- Background 0x3a
      12'h3A1: dout <= 8'b00000000; //  929 :   0 - 0x0
      12'h3A2: dout <= 8'b00000000; //  930 :   0 - 0x0
      12'h3A3: dout <= 8'b00000000; //  931 :   0 - 0x0
      12'h3A4: dout <= 8'b00000000; //  932 :   0 - 0x0
      12'h3A5: dout <= 8'b00000000; //  933 :   0 - 0x0
      12'h3A6: dout <= 8'b00000000; //  934 :   0 - 0x0
      12'h3A7: dout <= 8'b00000000; //  935 :   0 - 0x0
      12'h3A8: dout <= 8'b00000000; //  936 :   0 - 0x0 -- plane 1
      12'h3A9: dout <= 8'b00000000; //  937 :   0 - 0x0
      12'h3AA: dout <= 8'b00000000; //  938 :   0 - 0x0
      12'h3AB: dout <= 8'b00000000; //  939 :   0 - 0x0
      12'h3AC: dout <= 8'b00000000; //  940 :   0 - 0x0
      12'h3AD: dout <= 8'b00000000; //  941 :   0 - 0x0
      12'h3AE: dout <= 8'b00000000; //  942 :   0 - 0x0
      12'h3AF: dout <= 8'b00000000; //  943 :   0 - 0x0
      12'h3B0: dout <= 8'b00000000; //  944 :   0 - 0x0 -- Background 0x3b
      12'h3B1: dout <= 8'b00000000; //  945 :   0 - 0x0
      12'h3B2: dout <= 8'b00000000; //  946 :   0 - 0x0
      12'h3B3: dout <= 8'b00000000; //  947 :   0 - 0x0
      12'h3B4: dout <= 8'b00000000; //  948 :   0 - 0x0
      12'h3B5: dout <= 8'b00000000; //  949 :   0 - 0x0
      12'h3B6: dout <= 8'b00000000; //  950 :   0 - 0x0
      12'h3B7: dout <= 8'b00000000; //  951 :   0 - 0x0
      12'h3B8: dout <= 8'b00000000; //  952 :   0 - 0x0 -- plane 1
      12'h3B9: dout <= 8'b00000000; //  953 :   0 - 0x0
      12'h3BA: dout <= 8'b00000000; //  954 :   0 - 0x0
      12'h3BB: dout <= 8'b00000000; //  955 :   0 - 0x0
      12'h3BC: dout <= 8'b00000000; //  956 :   0 - 0x0
      12'h3BD: dout <= 8'b00000000; //  957 :   0 - 0x0
      12'h3BE: dout <= 8'b00000000; //  958 :   0 - 0x0
      12'h3BF: dout <= 8'b00000000; //  959 :   0 - 0x0
      12'h3C0: dout <= 8'b00000000; //  960 :   0 - 0x0 -- Background 0x3c
      12'h3C1: dout <= 8'b00000000; //  961 :   0 - 0x0
      12'h3C2: dout <= 8'b00000000; //  962 :   0 - 0x0
      12'h3C3: dout <= 8'b00000000; //  963 :   0 - 0x0
      12'h3C4: dout <= 8'b00000000; //  964 :   0 - 0x0
      12'h3C5: dout <= 8'b00000000; //  965 :   0 - 0x0
      12'h3C6: dout <= 8'b00000000; //  966 :   0 - 0x0
      12'h3C7: dout <= 8'b00000000; //  967 :   0 - 0x0
      12'h3C8: dout <= 8'b00000000; //  968 :   0 - 0x0 -- plane 1
      12'h3C9: dout <= 8'b00000000; //  969 :   0 - 0x0
      12'h3CA: dout <= 8'b00000000; //  970 :   0 - 0x0
      12'h3CB: dout <= 8'b00000000; //  971 :   0 - 0x0
      12'h3CC: dout <= 8'b00000000; //  972 :   0 - 0x0
      12'h3CD: dout <= 8'b00000000; //  973 :   0 - 0x0
      12'h3CE: dout <= 8'b00000000; //  974 :   0 - 0x0
      12'h3CF: dout <= 8'b00000000; //  975 :   0 - 0x0
      12'h3D0: dout <= 8'b00000000; //  976 :   0 - 0x0 -- Background 0x3d
      12'h3D1: dout <= 8'b00000000; //  977 :   0 - 0x0
      12'h3D2: dout <= 8'b00000000; //  978 :   0 - 0x0
      12'h3D3: dout <= 8'b00000000; //  979 :   0 - 0x0
      12'h3D4: dout <= 8'b00000000; //  980 :   0 - 0x0
      12'h3D5: dout <= 8'b00000000; //  981 :   0 - 0x0
      12'h3D6: dout <= 8'b00000000; //  982 :   0 - 0x0
      12'h3D7: dout <= 8'b00000000; //  983 :   0 - 0x0
      12'h3D8: dout <= 8'b00000000; //  984 :   0 - 0x0 -- plane 1
      12'h3D9: dout <= 8'b00000000; //  985 :   0 - 0x0
      12'h3DA: dout <= 8'b00000000; //  986 :   0 - 0x0
      12'h3DB: dout <= 8'b00000000; //  987 :   0 - 0x0
      12'h3DC: dout <= 8'b00000000; //  988 :   0 - 0x0
      12'h3DD: dout <= 8'b00000000; //  989 :   0 - 0x0
      12'h3DE: dout <= 8'b00000000; //  990 :   0 - 0x0
      12'h3DF: dout <= 8'b00000000; //  991 :   0 - 0x0
      12'h3E0: dout <= 8'b00000000; //  992 :   0 - 0x0 -- Background 0x3e
      12'h3E1: dout <= 8'b00000000; //  993 :   0 - 0x0
      12'h3E2: dout <= 8'b00000000; //  994 :   0 - 0x0
      12'h3E3: dout <= 8'b00000000; //  995 :   0 - 0x0
      12'h3E4: dout <= 8'b00000000; //  996 :   0 - 0x0
      12'h3E5: dout <= 8'b00000000; //  997 :   0 - 0x0
      12'h3E6: dout <= 8'b00000000; //  998 :   0 - 0x0
      12'h3E7: dout <= 8'b00000000; //  999 :   0 - 0x0
      12'h3E8: dout <= 8'b00000000; // 1000 :   0 - 0x0 -- plane 1
      12'h3E9: dout <= 8'b00000000; // 1001 :   0 - 0x0
      12'h3EA: dout <= 8'b00000000; // 1002 :   0 - 0x0
      12'h3EB: dout <= 8'b00000000; // 1003 :   0 - 0x0
      12'h3EC: dout <= 8'b00000000; // 1004 :   0 - 0x0
      12'h3ED: dout <= 8'b00000000; // 1005 :   0 - 0x0
      12'h3EE: dout <= 8'b00000000; // 1006 :   0 - 0x0
      12'h3EF: dout <= 8'b00000000; // 1007 :   0 - 0x0
      12'h3F0: dout <= 8'b00000000; // 1008 :   0 - 0x0 -- Background 0x3f
      12'h3F1: dout <= 8'b00000000; // 1009 :   0 - 0x0
      12'h3F2: dout <= 8'b00000000; // 1010 :   0 - 0x0
      12'h3F3: dout <= 8'b00000000; // 1011 :   0 - 0x0
      12'h3F4: dout <= 8'b00000000; // 1012 :   0 - 0x0
      12'h3F5: dout <= 8'b00000000; // 1013 :   0 - 0x0
      12'h3F6: dout <= 8'b00000000; // 1014 :   0 - 0x0
      12'h3F7: dout <= 8'b00000000; // 1015 :   0 - 0x0
      12'h3F8: dout <= 8'b00000000; // 1016 :   0 - 0x0 -- plane 1
      12'h3F9: dout <= 8'b00000000; // 1017 :   0 - 0x0
      12'h3FA: dout <= 8'b00000000; // 1018 :   0 - 0x0
      12'h3FB: dout <= 8'b00000000; // 1019 :   0 - 0x0
      12'h3FC: dout <= 8'b00000000; // 1020 :   0 - 0x0
      12'h3FD: dout <= 8'b00000000; // 1021 :   0 - 0x0
      12'h3FE: dout <= 8'b00000000; // 1022 :   0 - 0x0
      12'h3FF: dout <= 8'b00000000; // 1023 :   0 - 0x0
      12'h400: dout <= 8'b00000000; // 1024 :   0 - 0x0 -- Background 0x40
      12'h401: dout <= 8'b00000000; // 1025 :   0 - 0x0
      12'h402: dout <= 8'b00000000; // 1026 :   0 - 0x0
      12'h403: dout <= 8'b00000000; // 1027 :   0 - 0x0
      12'h404: dout <= 8'b00000000; // 1028 :   0 - 0x0
      12'h405: dout <= 8'b00000000; // 1029 :   0 - 0x0
      12'h406: dout <= 8'b00000000; // 1030 :   0 - 0x0
      12'h407: dout <= 8'b00000000; // 1031 :   0 - 0x0
      12'h408: dout <= 8'b00000000; // 1032 :   0 - 0x0 -- plane 1
      12'h409: dout <= 8'b00000000; // 1033 :   0 - 0x0
      12'h40A: dout <= 8'b00000000; // 1034 :   0 - 0x0
      12'h40B: dout <= 8'b00000000; // 1035 :   0 - 0x0
      12'h40C: dout <= 8'b00000000; // 1036 :   0 - 0x0
      12'h40D: dout <= 8'b00000000; // 1037 :   0 - 0x0
      12'h40E: dout <= 8'b00000000; // 1038 :   0 - 0x0
      12'h40F: dout <= 8'b00000000; // 1039 :   0 - 0x0
      12'h410: dout <= 8'b00000000; // 1040 :   0 - 0x0 -- Background 0x41
      12'h411: dout <= 8'b00000000; // 1041 :   0 - 0x0
      12'h412: dout <= 8'b00000000; // 1042 :   0 - 0x0
      12'h413: dout <= 8'b00000000; // 1043 :   0 - 0x0
      12'h414: dout <= 8'b00000000; // 1044 :   0 - 0x0
      12'h415: dout <= 8'b00000000; // 1045 :   0 - 0x0
      12'h416: dout <= 8'b00000000; // 1046 :   0 - 0x0
      12'h417: dout <= 8'b00000000; // 1047 :   0 - 0x0
      12'h418: dout <= 8'b00000000; // 1048 :   0 - 0x0 -- plane 1
      12'h419: dout <= 8'b00000000; // 1049 :   0 - 0x0
      12'h41A: dout <= 8'b00000000; // 1050 :   0 - 0x0
      12'h41B: dout <= 8'b00000000; // 1051 :   0 - 0x0
      12'h41C: dout <= 8'b00000000; // 1052 :   0 - 0x0
      12'h41D: dout <= 8'b00000000; // 1053 :   0 - 0x0
      12'h41E: dout <= 8'b00000000; // 1054 :   0 - 0x0
      12'h41F: dout <= 8'b00000000; // 1055 :   0 - 0x0
      12'h420: dout <= 8'b00000000; // 1056 :   0 - 0x0 -- Background 0x42
      12'h421: dout <= 8'b00000000; // 1057 :   0 - 0x0
      12'h422: dout <= 8'b00000000; // 1058 :   0 - 0x0
      12'h423: dout <= 8'b00000000; // 1059 :   0 - 0x0
      12'h424: dout <= 8'b00000000; // 1060 :   0 - 0x0
      12'h425: dout <= 8'b00000000; // 1061 :   0 - 0x0
      12'h426: dout <= 8'b00000000; // 1062 :   0 - 0x0
      12'h427: dout <= 8'b00000000; // 1063 :   0 - 0x0
      12'h428: dout <= 8'b00000000; // 1064 :   0 - 0x0 -- plane 1
      12'h429: dout <= 8'b00000000; // 1065 :   0 - 0x0
      12'h42A: dout <= 8'b00000000; // 1066 :   0 - 0x0
      12'h42B: dout <= 8'b00000000; // 1067 :   0 - 0x0
      12'h42C: dout <= 8'b00000000; // 1068 :   0 - 0x0
      12'h42D: dout <= 8'b00000000; // 1069 :   0 - 0x0
      12'h42E: dout <= 8'b00000000; // 1070 :   0 - 0x0
      12'h42F: dout <= 8'b00000000; // 1071 :   0 - 0x0
      12'h430: dout <= 8'b00000000; // 1072 :   0 - 0x0 -- Background 0x43
      12'h431: dout <= 8'b00000000; // 1073 :   0 - 0x0
      12'h432: dout <= 8'b00000000; // 1074 :   0 - 0x0
      12'h433: dout <= 8'b00000000; // 1075 :   0 - 0x0
      12'h434: dout <= 8'b00000000; // 1076 :   0 - 0x0
      12'h435: dout <= 8'b00000000; // 1077 :   0 - 0x0
      12'h436: dout <= 8'b00000000; // 1078 :   0 - 0x0
      12'h437: dout <= 8'b00000000; // 1079 :   0 - 0x0
      12'h438: dout <= 8'b00000000; // 1080 :   0 - 0x0 -- plane 1
      12'h439: dout <= 8'b00000000; // 1081 :   0 - 0x0
      12'h43A: dout <= 8'b00000000; // 1082 :   0 - 0x0
      12'h43B: dout <= 8'b00000000; // 1083 :   0 - 0x0
      12'h43C: dout <= 8'b00000000; // 1084 :   0 - 0x0
      12'h43D: dout <= 8'b00000000; // 1085 :   0 - 0x0
      12'h43E: dout <= 8'b00000000; // 1086 :   0 - 0x0
      12'h43F: dout <= 8'b00000000; // 1087 :   0 - 0x0
      12'h440: dout <= 8'b00000000; // 1088 :   0 - 0x0 -- Background 0x44
      12'h441: dout <= 8'b00000000; // 1089 :   0 - 0x0
      12'h442: dout <= 8'b00000000; // 1090 :   0 - 0x0
      12'h443: dout <= 8'b00000000; // 1091 :   0 - 0x0
      12'h444: dout <= 8'b00000000; // 1092 :   0 - 0x0
      12'h445: dout <= 8'b00000000; // 1093 :   0 - 0x0
      12'h446: dout <= 8'b00000000; // 1094 :   0 - 0x0
      12'h447: dout <= 8'b00000000; // 1095 :   0 - 0x0
      12'h448: dout <= 8'b00000000; // 1096 :   0 - 0x0 -- plane 1
      12'h449: dout <= 8'b00000000; // 1097 :   0 - 0x0
      12'h44A: dout <= 8'b00000000; // 1098 :   0 - 0x0
      12'h44B: dout <= 8'b00000000; // 1099 :   0 - 0x0
      12'h44C: dout <= 8'b00000000; // 1100 :   0 - 0x0
      12'h44D: dout <= 8'b00000000; // 1101 :   0 - 0x0
      12'h44E: dout <= 8'b00000000; // 1102 :   0 - 0x0
      12'h44F: dout <= 8'b00000000; // 1103 :   0 - 0x0
      12'h450: dout <= 8'b00000000; // 1104 :   0 - 0x0 -- Background 0x45
      12'h451: dout <= 8'b00000000; // 1105 :   0 - 0x0
      12'h452: dout <= 8'b00000000; // 1106 :   0 - 0x0
      12'h453: dout <= 8'b00000000; // 1107 :   0 - 0x0
      12'h454: dout <= 8'b00000000; // 1108 :   0 - 0x0
      12'h455: dout <= 8'b00000000; // 1109 :   0 - 0x0
      12'h456: dout <= 8'b00000000; // 1110 :   0 - 0x0
      12'h457: dout <= 8'b00000000; // 1111 :   0 - 0x0
      12'h458: dout <= 8'b00000000; // 1112 :   0 - 0x0 -- plane 1
      12'h459: dout <= 8'b00000000; // 1113 :   0 - 0x0
      12'h45A: dout <= 8'b00000000; // 1114 :   0 - 0x0
      12'h45B: dout <= 8'b00000000; // 1115 :   0 - 0x0
      12'h45C: dout <= 8'b00000000; // 1116 :   0 - 0x0
      12'h45D: dout <= 8'b00000000; // 1117 :   0 - 0x0
      12'h45E: dout <= 8'b00000000; // 1118 :   0 - 0x0
      12'h45F: dout <= 8'b00000000; // 1119 :   0 - 0x0
      12'h460: dout <= 8'b00000000; // 1120 :   0 - 0x0 -- Background 0x46
      12'h461: dout <= 8'b00000000; // 1121 :   0 - 0x0
      12'h462: dout <= 8'b00000000; // 1122 :   0 - 0x0
      12'h463: dout <= 8'b00000000; // 1123 :   0 - 0x0
      12'h464: dout <= 8'b00000000; // 1124 :   0 - 0x0
      12'h465: dout <= 8'b00000000; // 1125 :   0 - 0x0
      12'h466: dout <= 8'b00000000; // 1126 :   0 - 0x0
      12'h467: dout <= 8'b00000000; // 1127 :   0 - 0x0
      12'h468: dout <= 8'b00000000; // 1128 :   0 - 0x0 -- plane 1
      12'h469: dout <= 8'b00000000; // 1129 :   0 - 0x0
      12'h46A: dout <= 8'b00000000; // 1130 :   0 - 0x0
      12'h46B: dout <= 8'b00000000; // 1131 :   0 - 0x0
      12'h46C: dout <= 8'b00000000; // 1132 :   0 - 0x0
      12'h46D: dout <= 8'b00000000; // 1133 :   0 - 0x0
      12'h46E: dout <= 8'b00000000; // 1134 :   0 - 0x0
      12'h46F: dout <= 8'b00000000; // 1135 :   0 - 0x0
      12'h470: dout <= 8'b00000000; // 1136 :   0 - 0x0 -- Background 0x47
      12'h471: dout <= 8'b00000000; // 1137 :   0 - 0x0
      12'h472: dout <= 8'b00000000; // 1138 :   0 - 0x0
      12'h473: dout <= 8'b00000000; // 1139 :   0 - 0x0
      12'h474: dout <= 8'b00000000; // 1140 :   0 - 0x0
      12'h475: dout <= 8'b00000000; // 1141 :   0 - 0x0
      12'h476: dout <= 8'b00000000; // 1142 :   0 - 0x0
      12'h477: dout <= 8'b00000000; // 1143 :   0 - 0x0
      12'h478: dout <= 8'b00000000; // 1144 :   0 - 0x0 -- plane 1
      12'h479: dout <= 8'b00000000; // 1145 :   0 - 0x0
      12'h47A: dout <= 8'b00000000; // 1146 :   0 - 0x0
      12'h47B: dout <= 8'b00000000; // 1147 :   0 - 0x0
      12'h47C: dout <= 8'b00000000; // 1148 :   0 - 0x0
      12'h47D: dout <= 8'b00000000; // 1149 :   0 - 0x0
      12'h47E: dout <= 8'b00000000; // 1150 :   0 - 0x0
      12'h47F: dout <= 8'b00000000; // 1151 :   0 - 0x0
      12'h480: dout <= 8'b00000000; // 1152 :   0 - 0x0 -- Background 0x48
      12'h481: dout <= 8'b00000000; // 1153 :   0 - 0x0
      12'h482: dout <= 8'b00000000; // 1154 :   0 - 0x0
      12'h483: dout <= 8'b00000000; // 1155 :   0 - 0x0
      12'h484: dout <= 8'b00000000; // 1156 :   0 - 0x0
      12'h485: dout <= 8'b00000000; // 1157 :   0 - 0x0
      12'h486: dout <= 8'b00000000; // 1158 :   0 - 0x0
      12'h487: dout <= 8'b00000000; // 1159 :   0 - 0x0
      12'h488: dout <= 8'b00000000; // 1160 :   0 - 0x0 -- plane 1
      12'h489: dout <= 8'b00000000; // 1161 :   0 - 0x0
      12'h48A: dout <= 8'b00000000; // 1162 :   0 - 0x0
      12'h48B: dout <= 8'b00000000; // 1163 :   0 - 0x0
      12'h48C: dout <= 8'b00000000; // 1164 :   0 - 0x0
      12'h48D: dout <= 8'b00000000; // 1165 :   0 - 0x0
      12'h48E: dout <= 8'b00000000; // 1166 :   0 - 0x0
      12'h48F: dout <= 8'b00000000; // 1167 :   0 - 0x0
      12'h490: dout <= 8'b00000000; // 1168 :   0 - 0x0 -- Background 0x49
      12'h491: dout <= 8'b00000000; // 1169 :   0 - 0x0
      12'h492: dout <= 8'b00000000; // 1170 :   0 - 0x0
      12'h493: dout <= 8'b00000000; // 1171 :   0 - 0x0
      12'h494: dout <= 8'b00000000; // 1172 :   0 - 0x0
      12'h495: dout <= 8'b00000000; // 1173 :   0 - 0x0
      12'h496: dout <= 8'b00000000; // 1174 :   0 - 0x0
      12'h497: dout <= 8'b00000000; // 1175 :   0 - 0x0
      12'h498: dout <= 8'b00000000; // 1176 :   0 - 0x0 -- plane 1
      12'h499: dout <= 8'b00000000; // 1177 :   0 - 0x0
      12'h49A: dout <= 8'b00000000; // 1178 :   0 - 0x0
      12'h49B: dout <= 8'b00000000; // 1179 :   0 - 0x0
      12'h49C: dout <= 8'b00000000; // 1180 :   0 - 0x0
      12'h49D: dout <= 8'b00000000; // 1181 :   0 - 0x0
      12'h49E: dout <= 8'b00000000; // 1182 :   0 - 0x0
      12'h49F: dout <= 8'b00000000; // 1183 :   0 - 0x0
      12'h4A0: dout <= 8'b00000000; // 1184 :   0 - 0x0 -- Background 0x4a
      12'h4A1: dout <= 8'b00000000; // 1185 :   0 - 0x0
      12'h4A2: dout <= 8'b00000000; // 1186 :   0 - 0x0
      12'h4A3: dout <= 8'b00000000; // 1187 :   0 - 0x0
      12'h4A4: dout <= 8'b00000000; // 1188 :   0 - 0x0
      12'h4A5: dout <= 8'b00000000; // 1189 :   0 - 0x0
      12'h4A6: dout <= 8'b00000000; // 1190 :   0 - 0x0
      12'h4A7: dout <= 8'b00000000; // 1191 :   0 - 0x0
      12'h4A8: dout <= 8'b00000000; // 1192 :   0 - 0x0 -- plane 1
      12'h4A9: dout <= 8'b00000000; // 1193 :   0 - 0x0
      12'h4AA: dout <= 8'b00000000; // 1194 :   0 - 0x0
      12'h4AB: dout <= 8'b00000000; // 1195 :   0 - 0x0
      12'h4AC: dout <= 8'b00000000; // 1196 :   0 - 0x0
      12'h4AD: dout <= 8'b00000000; // 1197 :   0 - 0x0
      12'h4AE: dout <= 8'b00000000; // 1198 :   0 - 0x0
      12'h4AF: dout <= 8'b00000000; // 1199 :   0 - 0x0
      12'h4B0: dout <= 8'b00000000; // 1200 :   0 - 0x0 -- Background 0x4b
      12'h4B1: dout <= 8'b00000000; // 1201 :   0 - 0x0
      12'h4B2: dout <= 8'b00000000; // 1202 :   0 - 0x0
      12'h4B3: dout <= 8'b00000000; // 1203 :   0 - 0x0
      12'h4B4: dout <= 8'b00000000; // 1204 :   0 - 0x0
      12'h4B5: dout <= 8'b00000000; // 1205 :   0 - 0x0
      12'h4B6: dout <= 8'b00000000; // 1206 :   0 - 0x0
      12'h4B7: dout <= 8'b00000000; // 1207 :   0 - 0x0
      12'h4B8: dout <= 8'b00000000; // 1208 :   0 - 0x0 -- plane 1
      12'h4B9: dout <= 8'b00000000; // 1209 :   0 - 0x0
      12'h4BA: dout <= 8'b00000000; // 1210 :   0 - 0x0
      12'h4BB: dout <= 8'b00000000; // 1211 :   0 - 0x0
      12'h4BC: dout <= 8'b00000000; // 1212 :   0 - 0x0
      12'h4BD: dout <= 8'b00000000; // 1213 :   0 - 0x0
      12'h4BE: dout <= 8'b00000000; // 1214 :   0 - 0x0
      12'h4BF: dout <= 8'b00000000; // 1215 :   0 - 0x0
      12'h4C0: dout <= 8'b00000000; // 1216 :   0 - 0x0 -- Background 0x4c
      12'h4C1: dout <= 8'b00000000; // 1217 :   0 - 0x0
      12'h4C2: dout <= 8'b00000000; // 1218 :   0 - 0x0
      12'h4C3: dout <= 8'b00000000; // 1219 :   0 - 0x0
      12'h4C4: dout <= 8'b00000000; // 1220 :   0 - 0x0
      12'h4C5: dout <= 8'b00000000; // 1221 :   0 - 0x0
      12'h4C6: dout <= 8'b00000000; // 1222 :   0 - 0x0
      12'h4C7: dout <= 8'b00000000; // 1223 :   0 - 0x0
      12'h4C8: dout <= 8'b00000000; // 1224 :   0 - 0x0 -- plane 1
      12'h4C9: dout <= 8'b00000000; // 1225 :   0 - 0x0
      12'h4CA: dout <= 8'b00000000; // 1226 :   0 - 0x0
      12'h4CB: dout <= 8'b00000000; // 1227 :   0 - 0x0
      12'h4CC: dout <= 8'b00000000; // 1228 :   0 - 0x0
      12'h4CD: dout <= 8'b00000000; // 1229 :   0 - 0x0
      12'h4CE: dout <= 8'b00000000; // 1230 :   0 - 0x0
      12'h4CF: dout <= 8'b00000000; // 1231 :   0 - 0x0
      12'h4D0: dout <= 8'b00000000; // 1232 :   0 - 0x0 -- Background 0x4d
      12'h4D1: dout <= 8'b00000000; // 1233 :   0 - 0x0
      12'h4D2: dout <= 8'b00000000; // 1234 :   0 - 0x0
      12'h4D3: dout <= 8'b00000000; // 1235 :   0 - 0x0
      12'h4D4: dout <= 8'b00000000; // 1236 :   0 - 0x0
      12'h4D5: dout <= 8'b00000000; // 1237 :   0 - 0x0
      12'h4D6: dout <= 8'b00000000; // 1238 :   0 - 0x0
      12'h4D7: dout <= 8'b00000000; // 1239 :   0 - 0x0
      12'h4D8: dout <= 8'b00000000; // 1240 :   0 - 0x0 -- plane 1
      12'h4D9: dout <= 8'b00000000; // 1241 :   0 - 0x0
      12'h4DA: dout <= 8'b00000000; // 1242 :   0 - 0x0
      12'h4DB: dout <= 8'b00000000; // 1243 :   0 - 0x0
      12'h4DC: dout <= 8'b00000000; // 1244 :   0 - 0x0
      12'h4DD: dout <= 8'b00000000; // 1245 :   0 - 0x0
      12'h4DE: dout <= 8'b00000000; // 1246 :   0 - 0x0
      12'h4DF: dout <= 8'b00000000; // 1247 :   0 - 0x0
      12'h4E0: dout <= 8'b00000000; // 1248 :   0 - 0x0 -- Background 0x4e
      12'h4E1: dout <= 8'b00000000; // 1249 :   0 - 0x0
      12'h4E2: dout <= 8'b00000000; // 1250 :   0 - 0x0
      12'h4E3: dout <= 8'b00000000; // 1251 :   0 - 0x0
      12'h4E4: dout <= 8'b00000000; // 1252 :   0 - 0x0
      12'h4E5: dout <= 8'b00000000; // 1253 :   0 - 0x0
      12'h4E6: dout <= 8'b00000000; // 1254 :   0 - 0x0
      12'h4E7: dout <= 8'b00000000; // 1255 :   0 - 0x0
      12'h4E8: dout <= 8'b00000000; // 1256 :   0 - 0x0 -- plane 1
      12'h4E9: dout <= 8'b00000000; // 1257 :   0 - 0x0
      12'h4EA: dout <= 8'b00000000; // 1258 :   0 - 0x0
      12'h4EB: dout <= 8'b00000000; // 1259 :   0 - 0x0
      12'h4EC: dout <= 8'b00000000; // 1260 :   0 - 0x0
      12'h4ED: dout <= 8'b00000000; // 1261 :   0 - 0x0
      12'h4EE: dout <= 8'b00000000; // 1262 :   0 - 0x0
      12'h4EF: dout <= 8'b00000000; // 1263 :   0 - 0x0
      12'h4F0: dout <= 8'b00000000; // 1264 :   0 - 0x0 -- Background 0x4f
      12'h4F1: dout <= 8'b00000000; // 1265 :   0 - 0x0
      12'h4F2: dout <= 8'b00000000; // 1266 :   0 - 0x0
      12'h4F3: dout <= 8'b00000000; // 1267 :   0 - 0x0
      12'h4F4: dout <= 8'b00000000; // 1268 :   0 - 0x0
      12'h4F5: dout <= 8'b00000000; // 1269 :   0 - 0x0
      12'h4F6: dout <= 8'b00000000; // 1270 :   0 - 0x0
      12'h4F7: dout <= 8'b00000000; // 1271 :   0 - 0x0
      12'h4F8: dout <= 8'b00000000; // 1272 :   0 - 0x0 -- plane 1
      12'h4F9: dout <= 8'b00000000; // 1273 :   0 - 0x0
      12'h4FA: dout <= 8'b00000000; // 1274 :   0 - 0x0
      12'h4FB: dout <= 8'b00000000; // 1275 :   0 - 0x0
      12'h4FC: dout <= 8'b00000000; // 1276 :   0 - 0x0
      12'h4FD: dout <= 8'b00000000; // 1277 :   0 - 0x0
      12'h4FE: dout <= 8'b00000000; // 1278 :   0 - 0x0
      12'h4FF: dout <= 8'b00000000; // 1279 :   0 - 0x0
      12'h500: dout <= 8'b00000000; // 1280 :   0 - 0x0 -- Background 0x50
      12'h501: dout <= 8'b00000000; // 1281 :   0 - 0x0
      12'h502: dout <= 8'b00000000; // 1282 :   0 - 0x0
      12'h503: dout <= 8'b00000000; // 1283 :   0 - 0x0
      12'h504: dout <= 8'b00000000; // 1284 :   0 - 0x0
      12'h505: dout <= 8'b00000000; // 1285 :   0 - 0x0
      12'h506: dout <= 8'b00000000; // 1286 :   0 - 0x0
      12'h507: dout <= 8'b00000000; // 1287 :   0 - 0x0
      12'h508: dout <= 8'b00000000; // 1288 :   0 - 0x0 -- plane 1
      12'h509: dout <= 8'b00000000; // 1289 :   0 - 0x0
      12'h50A: dout <= 8'b00000000; // 1290 :   0 - 0x0
      12'h50B: dout <= 8'b00000000; // 1291 :   0 - 0x0
      12'h50C: dout <= 8'b00000000; // 1292 :   0 - 0x0
      12'h50D: dout <= 8'b00000000; // 1293 :   0 - 0x0
      12'h50E: dout <= 8'b00000000; // 1294 :   0 - 0x0
      12'h50F: dout <= 8'b00000000; // 1295 :   0 - 0x0
      12'h510: dout <= 8'b00000000; // 1296 :   0 - 0x0 -- Background 0x51
      12'h511: dout <= 8'b00000000; // 1297 :   0 - 0x0
      12'h512: dout <= 8'b00000000; // 1298 :   0 - 0x0
      12'h513: dout <= 8'b00000000; // 1299 :   0 - 0x0
      12'h514: dout <= 8'b00000000; // 1300 :   0 - 0x0
      12'h515: dout <= 8'b00000000; // 1301 :   0 - 0x0
      12'h516: dout <= 8'b00000000; // 1302 :   0 - 0x0
      12'h517: dout <= 8'b00000000; // 1303 :   0 - 0x0
      12'h518: dout <= 8'b00000000; // 1304 :   0 - 0x0 -- plane 1
      12'h519: dout <= 8'b00000000; // 1305 :   0 - 0x0
      12'h51A: dout <= 8'b00000000; // 1306 :   0 - 0x0
      12'h51B: dout <= 8'b00000000; // 1307 :   0 - 0x0
      12'h51C: dout <= 8'b00000000; // 1308 :   0 - 0x0
      12'h51D: dout <= 8'b00000000; // 1309 :   0 - 0x0
      12'h51E: dout <= 8'b00000000; // 1310 :   0 - 0x0
      12'h51F: dout <= 8'b00000000; // 1311 :   0 - 0x0
      12'h520: dout <= 8'b00000000; // 1312 :   0 - 0x0 -- Background 0x52
      12'h521: dout <= 8'b00000000; // 1313 :   0 - 0x0
      12'h522: dout <= 8'b00000000; // 1314 :   0 - 0x0
      12'h523: dout <= 8'b00000000; // 1315 :   0 - 0x0
      12'h524: dout <= 8'b00000000; // 1316 :   0 - 0x0
      12'h525: dout <= 8'b00000000; // 1317 :   0 - 0x0
      12'h526: dout <= 8'b00000000; // 1318 :   0 - 0x0
      12'h527: dout <= 8'b00000000; // 1319 :   0 - 0x0
      12'h528: dout <= 8'b00000000; // 1320 :   0 - 0x0 -- plane 1
      12'h529: dout <= 8'b00000000; // 1321 :   0 - 0x0
      12'h52A: dout <= 8'b00000000; // 1322 :   0 - 0x0
      12'h52B: dout <= 8'b00000000; // 1323 :   0 - 0x0
      12'h52C: dout <= 8'b00000000; // 1324 :   0 - 0x0
      12'h52D: dout <= 8'b00000000; // 1325 :   0 - 0x0
      12'h52E: dout <= 8'b00000000; // 1326 :   0 - 0x0
      12'h52F: dout <= 8'b00000000; // 1327 :   0 - 0x0
      12'h530: dout <= 8'b00000000; // 1328 :   0 - 0x0 -- Background 0x53
      12'h531: dout <= 8'b00000000; // 1329 :   0 - 0x0
      12'h532: dout <= 8'b00000000; // 1330 :   0 - 0x0
      12'h533: dout <= 8'b00000000; // 1331 :   0 - 0x0
      12'h534: dout <= 8'b00000000; // 1332 :   0 - 0x0
      12'h535: dout <= 8'b00000000; // 1333 :   0 - 0x0
      12'h536: dout <= 8'b00000000; // 1334 :   0 - 0x0
      12'h537: dout <= 8'b00000000; // 1335 :   0 - 0x0
      12'h538: dout <= 8'b00000000; // 1336 :   0 - 0x0 -- plane 1
      12'h539: dout <= 8'b00000000; // 1337 :   0 - 0x0
      12'h53A: dout <= 8'b00000000; // 1338 :   0 - 0x0
      12'h53B: dout <= 8'b00000000; // 1339 :   0 - 0x0
      12'h53C: dout <= 8'b00000000; // 1340 :   0 - 0x0
      12'h53D: dout <= 8'b00000000; // 1341 :   0 - 0x0
      12'h53E: dout <= 8'b00000000; // 1342 :   0 - 0x0
      12'h53F: dout <= 8'b00000000; // 1343 :   0 - 0x0
      12'h540: dout <= 8'b00000000; // 1344 :   0 - 0x0 -- Background 0x54
      12'h541: dout <= 8'b00000000; // 1345 :   0 - 0x0
      12'h542: dout <= 8'b00000000; // 1346 :   0 - 0x0
      12'h543: dout <= 8'b00000000; // 1347 :   0 - 0x0
      12'h544: dout <= 8'b00000000; // 1348 :   0 - 0x0
      12'h545: dout <= 8'b00000000; // 1349 :   0 - 0x0
      12'h546: dout <= 8'b00000000; // 1350 :   0 - 0x0
      12'h547: dout <= 8'b00000000; // 1351 :   0 - 0x0
      12'h548: dout <= 8'b00000000; // 1352 :   0 - 0x0 -- plane 1
      12'h549: dout <= 8'b00000000; // 1353 :   0 - 0x0
      12'h54A: dout <= 8'b00000000; // 1354 :   0 - 0x0
      12'h54B: dout <= 8'b00000000; // 1355 :   0 - 0x0
      12'h54C: dout <= 8'b00000000; // 1356 :   0 - 0x0
      12'h54D: dout <= 8'b00000000; // 1357 :   0 - 0x0
      12'h54E: dout <= 8'b00000000; // 1358 :   0 - 0x0
      12'h54F: dout <= 8'b00000000; // 1359 :   0 - 0x0
      12'h550: dout <= 8'b00000000; // 1360 :   0 - 0x0 -- Background 0x55
      12'h551: dout <= 8'b00000000; // 1361 :   0 - 0x0
      12'h552: dout <= 8'b00000000; // 1362 :   0 - 0x0
      12'h553: dout <= 8'b00000000; // 1363 :   0 - 0x0
      12'h554: dout <= 8'b00000000; // 1364 :   0 - 0x0
      12'h555: dout <= 8'b00000000; // 1365 :   0 - 0x0
      12'h556: dout <= 8'b00000000; // 1366 :   0 - 0x0
      12'h557: dout <= 8'b00000000; // 1367 :   0 - 0x0
      12'h558: dout <= 8'b00000000; // 1368 :   0 - 0x0 -- plane 1
      12'h559: dout <= 8'b00000000; // 1369 :   0 - 0x0
      12'h55A: dout <= 8'b00000000; // 1370 :   0 - 0x0
      12'h55B: dout <= 8'b00000000; // 1371 :   0 - 0x0
      12'h55C: dout <= 8'b00000000; // 1372 :   0 - 0x0
      12'h55D: dout <= 8'b00000000; // 1373 :   0 - 0x0
      12'h55E: dout <= 8'b00000000; // 1374 :   0 - 0x0
      12'h55F: dout <= 8'b00000000; // 1375 :   0 - 0x0
      12'h560: dout <= 8'b00000000; // 1376 :   0 - 0x0 -- Background 0x56
      12'h561: dout <= 8'b00000000; // 1377 :   0 - 0x0
      12'h562: dout <= 8'b00000000; // 1378 :   0 - 0x0
      12'h563: dout <= 8'b00000000; // 1379 :   0 - 0x0
      12'h564: dout <= 8'b00000000; // 1380 :   0 - 0x0
      12'h565: dout <= 8'b00000000; // 1381 :   0 - 0x0
      12'h566: dout <= 8'b00000000; // 1382 :   0 - 0x0
      12'h567: dout <= 8'b00000000; // 1383 :   0 - 0x0
      12'h568: dout <= 8'b00000000; // 1384 :   0 - 0x0 -- plane 1
      12'h569: dout <= 8'b00000000; // 1385 :   0 - 0x0
      12'h56A: dout <= 8'b00000000; // 1386 :   0 - 0x0
      12'h56B: dout <= 8'b00000000; // 1387 :   0 - 0x0
      12'h56C: dout <= 8'b00000000; // 1388 :   0 - 0x0
      12'h56D: dout <= 8'b00000000; // 1389 :   0 - 0x0
      12'h56E: dout <= 8'b00000000; // 1390 :   0 - 0x0
      12'h56F: dout <= 8'b00000000; // 1391 :   0 - 0x0
      12'h570: dout <= 8'b00000000; // 1392 :   0 - 0x0 -- Background 0x57
      12'h571: dout <= 8'b00000000; // 1393 :   0 - 0x0
      12'h572: dout <= 8'b00000000; // 1394 :   0 - 0x0
      12'h573: dout <= 8'b00000000; // 1395 :   0 - 0x0
      12'h574: dout <= 8'b00000000; // 1396 :   0 - 0x0
      12'h575: dout <= 8'b00000000; // 1397 :   0 - 0x0
      12'h576: dout <= 8'b00000000; // 1398 :   0 - 0x0
      12'h577: dout <= 8'b00000000; // 1399 :   0 - 0x0
      12'h578: dout <= 8'b00000000; // 1400 :   0 - 0x0 -- plane 1
      12'h579: dout <= 8'b00000000; // 1401 :   0 - 0x0
      12'h57A: dout <= 8'b00000000; // 1402 :   0 - 0x0
      12'h57B: dout <= 8'b00000000; // 1403 :   0 - 0x0
      12'h57C: dout <= 8'b00000000; // 1404 :   0 - 0x0
      12'h57D: dout <= 8'b00000000; // 1405 :   0 - 0x0
      12'h57E: dout <= 8'b00000000; // 1406 :   0 - 0x0
      12'h57F: dout <= 8'b00000000; // 1407 :   0 - 0x0
      12'h580: dout <= 8'b00000000; // 1408 :   0 - 0x0 -- Background 0x58
      12'h581: dout <= 8'b00000000; // 1409 :   0 - 0x0
      12'h582: dout <= 8'b00000000; // 1410 :   0 - 0x0
      12'h583: dout <= 8'b00000000; // 1411 :   0 - 0x0
      12'h584: dout <= 8'b00000000; // 1412 :   0 - 0x0
      12'h585: dout <= 8'b00000000; // 1413 :   0 - 0x0
      12'h586: dout <= 8'b00000000; // 1414 :   0 - 0x0
      12'h587: dout <= 8'b00000000; // 1415 :   0 - 0x0
      12'h588: dout <= 8'b00000000; // 1416 :   0 - 0x0 -- plane 1
      12'h589: dout <= 8'b00000000; // 1417 :   0 - 0x0
      12'h58A: dout <= 8'b00000000; // 1418 :   0 - 0x0
      12'h58B: dout <= 8'b00000000; // 1419 :   0 - 0x0
      12'h58C: dout <= 8'b00000000; // 1420 :   0 - 0x0
      12'h58D: dout <= 8'b00000000; // 1421 :   0 - 0x0
      12'h58E: dout <= 8'b00000000; // 1422 :   0 - 0x0
      12'h58F: dout <= 8'b00000000; // 1423 :   0 - 0x0
      12'h590: dout <= 8'b00000000; // 1424 :   0 - 0x0 -- Background 0x59
      12'h591: dout <= 8'b00000000; // 1425 :   0 - 0x0
      12'h592: dout <= 8'b00000000; // 1426 :   0 - 0x0
      12'h593: dout <= 8'b00000000; // 1427 :   0 - 0x0
      12'h594: dout <= 8'b00000000; // 1428 :   0 - 0x0
      12'h595: dout <= 8'b00000000; // 1429 :   0 - 0x0
      12'h596: dout <= 8'b00000000; // 1430 :   0 - 0x0
      12'h597: dout <= 8'b00000000; // 1431 :   0 - 0x0
      12'h598: dout <= 8'b00000000; // 1432 :   0 - 0x0 -- plane 1
      12'h599: dout <= 8'b00000000; // 1433 :   0 - 0x0
      12'h59A: dout <= 8'b00000000; // 1434 :   0 - 0x0
      12'h59B: dout <= 8'b00000000; // 1435 :   0 - 0x0
      12'h59C: dout <= 8'b00000000; // 1436 :   0 - 0x0
      12'h59D: dout <= 8'b00000000; // 1437 :   0 - 0x0
      12'h59E: dout <= 8'b00000000; // 1438 :   0 - 0x0
      12'h59F: dout <= 8'b00000000; // 1439 :   0 - 0x0
      12'h5A0: dout <= 8'b00000000; // 1440 :   0 - 0x0 -- Background 0x5a
      12'h5A1: dout <= 8'b00000000; // 1441 :   0 - 0x0
      12'h5A2: dout <= 8'b00000000; // 1442 :   0 - 0x0
      12'h5A3: dout <= 8'b00000000; // 1443 :   0 - 0x0
      12'h5A4: dout <= 8'b00000000; // 1444 :   0 - 0x0
      12'h5A5: dout <= 8'b00000000; // 1445 :   0 - 0x0
      12'h5A6: dout <= 8'b00000000; // 1446 :   0 - 0x0
      12'h5A7: dout <= 8'b00000000; // 1447 :   0 - 0x0
      12'h5A8: dout <= 8'b00000000; // 1448 :   0 - 0x0 -- plane 1
      12'h5A9: dout <= 8'b00000000; // 1449 :   0 - 0x0
      12'h5AA: dout <= 8'b00000000; // 1450 :   0 - 0x0
      12'h5AB: dout <= 8'b00000000; // 1451 :   0 - 0x0
      12'h5AC: dout <= 8'b00000000; // 1452 :   0 - 0x0
      12'h5AD: dout <= 8'b00000000; // 1453 :   0 - 0x0
      12'h5AE: dout <= 8'b00000000; // 1454 :   0 - 0x0
      12'h5AF: dout <= 8'b00000000; // 1455 :   0 - 0x0
      12'h5B0: dout <= 8'b00000000; // 1456 :   0 - 0x0 -- Background 0x5b
      12'h5B1: dout <= 8'b00000000; // 1457 :   0 - 0x0
      12'h5B2: dout <= 8'b00000000; // 1458 :   0 - 0x0
      12'h5B3: dout <= 8'b00000000; // 1459 :   0 - 0x0
      12'h5B4: dout <= 8'b00000000; // 1460 :   0 - 0x0
      12'h5B5: dout <= 8'b00000000; // 1461 :   0 - 0x0
      12'h5B6: dout <= 8'b00000000; // 1462 :   0 - 0x0
      12'h5B7: dout <= 8'b00000000; // 1463 :   0 - 0x0
      12'h5B8: dout <= 8'b00000000; // 1464 :   0 - 0x0 -- plane 1
      12'h5B9: dout <= 8'b00000000; // 1465 :   0 - 0x0
      12'h5BA: dout <= 8'b00000000; // 1466 :   0 - 0x0
      12'h5BB: dout <= 8'b00000000; // 1467 :   0 - 0x0
      12'h5BC: dout <= 8'b00000000; // 1468 :   0 - 0x0
      12'h5BD: dout <= 8'b00000000; // 1469 :   0 - 0x0
      12'h5BE: dout <= 8'b00000000; // 1470 :   0 - 0x0
      12'h5BF: dout <= 8'b00000000; // 1471 :   0 - 0x0
      12'h5C0: dout <= 8'b00000000; // 1472 :   0 - 0x0 -- Background 0x5c
      12'h5C1: dout <= 8'b00000000; // 1473 :   0 - 0x0
      12'h5C2: dout <= 8'b00000000; // 1474 :   0 - 0x0
      12'h5C3: dout <= 8'b00000000; // 1475 :   0 - 0x0
      12'h5C4: dout <= 8'b00000000; // 1476 :   0 - 0x0
      12'h5C5: dout <= 8'b00000000; // 1477 :   0 - 0x0
      12'h5C6: dout <= 8'b00000000; // 1478 :   0 - 0x0
      12'h5C7: dout <= 8'b00000000; // 1479 :   0 - 0x0
      12'h5C8: dout <= 8'b00000000; // 1480 :   0 - 0x0 -- plane 1
      12'h5C9: dout <= 8'b00000000; // 1481 :   0 - 0x0
      12'h5CA: dout <= 8'b00000000; // 1482 :   0 - 0x0
      12'h5CB: dout <= 8'b00000000; // 1483 :   0 - 0x0
      12'h5CC: dout <= 8'b00000000; // 1484 :   0 - 0x0
      12'h5CD: dout <= 8'b00000000; // 1485 :   0 - 0x0
      12'h5CE: dout <= 8'b00000000; // 1486 :   0 - 0x0
      12'h5CF: dout <= 8'b00000000; // 1487 :   0 - 0x0
      12'h5D0: dout <= 8'b00000000; // 1488 :   0 - 0x0 -- Background 0x5d
      12'h5D1: dout <= 8'b00000000; // 1489 :   0 - 0x0
      12'h5D2: dout <= 8'b00000000; // 1490 :   0 - 0x0
      12'h5D3: dout <= 8'b00000000; // 1491 :   0 - 0x0
      12'h5D4: dout <= 8'b00000000; // 1492 :   0 - 0x0
      12'h5D5: dout <= 8'b00000000; // 1493 :   0 - 0x0
      12'h5D6: dout <= 8'b00000000; // 1494 :   0 - 0x0
      12'h5D7: dout <= 8'b00000000; // 1495 :   0 - 0x0
      12'h5D8: dout <= 8'b00000000; // 1496 :   0 - 0x0 -- plane 1
      12'h5D9: dout <= 8'b00000000; // 1497 :   0 - 0x0
      12'h5DA: dout <= 8'b00000000; // 1498 :   0 - 0x0
      12'h5DB: dout <= 8'b00000000; // 1499 :   0 - 0x0
      12'h5DC: dout <= 8'b00000000; // 1500 :   0 - 0x0
      12'h5DD: dout <= 8'b00000000; // 1501 :   0 - 0x0
      12'h5DE: dout <= 8'b00000000; // 1502 :   0 - 0x0
      12'h5DF: dout <= 8'b00000000; // 1503 :   0 - 0x0
      12'h5E0: dout <= 8'b00000000; // 1504 :   0 - 0x0 -- Background 0x5e
      12'h5E1: dout <= 8'b00000000; // 1505 :   0 - 0x0
      12'h5E2: dout <= 8'b00000000; // 1506 :   0 - 0x0
      12'h5E3: dout <= 8'b00000000; // 1507 :   0 - 0x0
      12'h5E4: dout <= 8'b00000000; // 1508 :   0 - 0x0
      12'h5E5: dout <= 8'b00000000; // 1509 :   0 - 0x0
      12'h5E6: dout <= 8'b00000000; // 1510 :   0 - 0x0
      12'h5E7: dout <= 8'b00000000; // 1511 :   0 - 0x0
      12'h5E8: dout <= 8'b00000000; // 1512 :   0 - 0x0 -- plane 1
      12'h5E9: dout <= 8'b00000000; // 1513 :   0 - 0x0
      12'h5EA: dout <= 8'b00000000; // 1514 :   0 - 0x0
      12'h5EB: dout <= 8'b00000000; // 1515 :   0 - 0x0
      12'h5EC: dout <= 8'b00000000; // 1516 :   0 - 0x0
      12'h5ED: dout <= 8'b00000000; // 1517 :   0 - 0x0
      12'h5EE: dout <= 8'b00000000; // 1518 :   0 - 0x0
      12'h5EF: dout <= 8'b00000000; // 1519 :   0 - 0x0
      12'h5F0: dout <= 8'b00000000; // 1520 :   0 - 0x0 -- Background 0x5f
      12'h5F1: dout <= 8'b00000000; // 1521 :   0 - 0x0
      12'h5F2: dout <= 8'b00000000; // 1522 :   0 - 0x0
      12'h5F3: dout <= 8'b00000000; // 1523 :   0 - 0x0
      12'h5F4: dout <= 8'b00000000; // 1524 :   0 - 0x0
      12'h5F5: dout <= 8'b00000000; // 1525 :   0 - 0x0
      12'h5F6: dout <= 8'b00000000; // 1526 :   0 - 0x0
      12'h5F7: dout <= 8'b00000000; // 1527 :   0 - 0x0
      12'h5F8: dout <= 8'b00000000; // 1528 :   0 - 0x0 -- plane 1
      12'h5F9: dout <= 8'b00000000; // 1529 :   0 - 0x0
      12'h5FA: dout <= 8'b00000000; // 1530 :   0 - 0x0
      12'h5FB: dout <= 8'b00000000; // 1531 :   0 - 0x0
      12'h5FC: dout <= 8'b00000000; // 1532 :   0 - 0x0
      12'h5FD: dout <= 8'b00000000; // 1533 :   0 - 0x0
      12'h5FE: dout <= 8'b00000000; // 1534 :   0 - 0x0
      12'h5FF: dout <= 8'b00000000; // 1535 :   0 - 0x0
      12'h600: dout <= 8'b00000000; // 1536 :   0 - 0x0 -- Background 0x60
      12'h601: dout <= 8'b00000000; // 1537 :   0 - 0x0
      12'h602: dout <= 8'b00000000; // 1538 :   0 - 0x0
      12'h603: dout <= 8'b00000000; // 1539 :   0 - 0x0
      12'h604: dout <= 8'b00000000; // 1540 :   0 - 0x0
      12'h605: dout <= 8'b00000000; // 1541 :   0 - 0x0
      12'h606: dout <= 8'b00000000; // 1542 :   0 - 0x0
      12'h607: dout <= 8'b00000000; // 1543 :   0 - 0x0
      12'h608: dout <= 8'b00000000; // 1544 :   0 - 0x0 -- plane 1
      12'h609: dout <= 8'b00000000; // 1545 :   0 - 0x0
      12'h60A: dout <= 8'b00000000; // 1546 :   0 - 0x0
      12'h60B: dout <= 8'b00000000; // 1547 :   0 - 0x0
      12'h60C: dout <= 8'b00000000; // 1548 :   0 - 0x0
      12'h60D: dout <= 8'b00000000; // 1549 :   0 - 0x0
      12'h60E: dout <= 8'b00000000; // 1550 :   0 - 0x0
      12'h60F: dout <= 8'b00000000; // 1551 :   0 - 0x0
      12'h610: dout <= 8'b00000000; // 1552 :   0 - 0x0 -- Background 0x61
      12'h611: dout <= 8'b00000000; // 1553 :   0 - 0x0
      12'h612: dout <= 8'b00000000; // 1554 :   0 - 0x0
      12'h613: dout <= 8'b00000000; // 1555 :   0 - 0x0
      12'h614: dout <= 8'b00000000; // 1556 :   0 - 0x0
      12'h615: dout <= 8'b00000000; // 1557 :   0 - 0x0
      12'h616: dout <= 8'b00000000; // 1558 :   0 - 0x0
      12'h617: dout <= 8'b00000000; // 1559 :   0 - 0x0
      12'h618: dout <= 8'b00000000; // 1560 :   0 - 0x0 -- plane 1
      12'h619: dout <= 8'b00000000; // 1561 :   0 - 0x0
      12'h61A: dout <= 8'b00000000; // 1562 :   0 - 0x0
      12'h61B: dout <= 8'b00000000; // 1563 :   0 - 0x0
      12'h61C: dout <= 8'b00000000; // 1564 :   0 - 0x0
      12'h61D: dout <= 8'b00000000; // 1565 :   0 - 0x0
      12'h61E: dout <= 8'b00000000; // 1566 :   0 - 0x0
      12'h61F: dout <= 8'b00000000; // 1567 :   0 - 0x0
      12'h620: dout <= 8'b00000000; // 1568 :   0 - 0x0 -- Background 0x62
      12'h621: dout <= 8'b00000000; // 1569 :   0 - 0x0
      12'h622: dout <= 8'b00000000; // 1570 :   0 - 0x0
      12'h623: dout <= 8'b00000000; // 1571 :   0 - 0x0
      12'h624: dout <= 8'b00000000; // 1572 :   0 - 0x0
      12'h625: dout <= 8'b00000000; // 1573 :   0 - 0x0
      12'h626: dout <= 8'b00000000; // 1574 :   0 - 0x0
      12'h627: dout <= 8'b00000000; // 1575 :   0 - 0x0
      12'h628: dout <= 8'b00000000; // 1576 :   0 - 0x0 -- plane 1
      12'h629: dout <= 8'b00000000; // 1577 :   0 - 0x0
      12'h62A: dout <= 8'b00000000; // 1578 :   0 - 0x0
      12'h62B: dout <= 8'b00000000; // 1579 :   0 - 0x0
      12'h62C: dout <= 8'b00000000; // 1580 :   0 - 0x0
      12'h62D: dout <= 8'b00000000; // 1581 :   0 - 0x0
      12'h62E: dout <= 8'b00000000; // 1582 :   0 - 0x0
      12'h62F: dout <= 8'b00000000; // 1583 :   0 - 0x0
      12'h630: dout <= 8'b00000000; // 1584 :   0 - 0x0 -- Background 0x63
      12'h631: dout <= 8'b00000000; // 1585 :   0 - 0x0
      12'h632: dout <= 8'b00000000; // 1586 :   0 - 0x0
      12'h633: dout <= 8'b00000000; // 1587 :   0 - 0x0
      12'h634: dout <= 8'b00000000; // 1588 :   0 - 0x0
      12'h635: dout <= 8'b00000000; // 1589 :   0 - 0x0
      12'h636: dout <= 8'b00000000; // 1590 :   0 - 0x0
      12'h637: dout <= 8'b00000000; // 1591 :   0 - 0x0
      12'h638: dout <= 8'b00000000; // 1592 :   0 - 0x0 -- plane 1
      12'h639: dout <= 8'b00000000; // 1593 :   0 - 0x0
      12'h63A: dout <= 8'b00000000; // 1594 :   0 - 0x0
      12'h63B: dout <= 8'b00000000; // 1595 :   0 - 0x0
      12'h63C: dout <= 8'b00000000; // 1596 :   0 - 0x0
      12'h63D: dout <= 8'b00000000; // 1597 :   0 - 0x0
      12'h63E: dout <= 8'b00000000; // 1598 :   0 - 0x0
      12'h63F: dout <= 8'b00000000; // 1599 :   0 - 0x0
      12'h640: dout <= 8'b00000000; // 1600 :   0 - 0x0 -- Background 0x64
      12'h641: dout <= 8'b00000000; // 1601 :   0 - 0x0
      12'h642: dout <= 8'b00000000; // 1602 :   0 - 0x0
      12'h643: dout <= 8'b00000000; // 1603 :   0 - 0x0
      12'h644: dout <= 8'b00000000; // 1604 :   0 - 0x0
      12'h645: dout <= 8'b00000000; // 1605 :   0 - 0x0
      12'h646: dout <= 8'b00000000; // 1606 :   0 - 0x0
      12'h647: dout <= 8'b00000000; // 1607 :   0 - 0x0
      12'h648: dout <= 8'b00000000; // 1608 :   0 - 0x0 -- plane 1
      12'h649: dout <= 8'b00000000; // 1609 :   0 - 0x0
      12'h64A: dout <= 8'b00000000; // 1610 :   0 - 0x0
      12'h64B: dout <= 8'b00000000; // 1611 :   0 - 0x0
      12'h64C: dout <= 8'b00000000; // 1612 :   0 - 0x0
      12'h64D: dout <= 8'b00000000; // 1613 :   0 - 0x0
      12'h64E: dout <= 8'b00000000; // 1614 :   0 - 0x0
      12'h64F: dout <= 8'b00000000; // 1615 :   0 - 0x0
      12'h650: dout <= 8'b00000000; // 1616 :   0 - 0x0 -- Background 0x65
      12'h651: dout <= 8'b00000000; // 1617 :   0 - 0x0
      12'h652: dout <= 8'b00000000; // 1618 :   0 - 0x0
      12'h653: dout <= 8'b00000000; // 1619 :   0 - 0x0
      12'h654: dout <= 8'b00000000; // 1620 :   0 - 0x0
      12'h655: dout <= 8'b00000000; // 1621 :   0 - 0x0
      12'h656: dout <= 8'b00000000; // 1622 :   0 - 0x0
      12'h657: dout <= 8'b00000000; // 1623 :   0 - 0x0
      12'h658: dout <= 8'b00000000; // 1624 :   0 - 0x0 -- plane 1
      12'h659: dout <= 8'b00000000; // 1625 :   0 - 0x0
      12'h65A: dout <= 8'b00000000; // 1626 :   0 - 0x0
      12'h65B: dout <= 8'b00000000; // 1627 :   0 - 0x0
      12'h65C: dout <= 8'b00000000; // 1628 :   0 - 0x0
      12'h65D: dout <= 8'b00000000; // 1629 :   0 - 0x0
      12'h65E: dout <= 8'b00000000; // 1630 :   0 - 0x0
      12'h65F: dout <= 8'b00000000; // 1631 :   0 - 0x0
      12'h660: dout <= 8'b00000000; // 1632 :   0 - 0x0 -- Background 0x66
      12'h661: dout <= 8'b00000000; // 1633 :   0 - 0x0
      12'h662: dout <= 8'b00000000; // 1634 :   0 - 0x0
      12'h663: dout <= 8'b00000000; // 1635 :   0 - 0x0
      12'h664: dout <= 8'b00000000; // 1636 :   0 - 0x0
      12'h665: dout <= 8'b00000000; // 1637 :   0 - 0x0
      12'h666: dout <= 8'b00000000; // 1638 :   0 - 0x0
      12'h667: dout <= 8'b00000000; // 1639 :   0 - 0x0
      12'h668: dout <= 8'b00000000; // 1640 :   0 - 0x0 -- plane 1
      12'h669: dout <= 8'b00000000; // 1641 :   0 - 0x0
      12'h66A: dout <= 8'b00000000; // 1642 :   0 - 0x0
      12'h66B: dout <= 8'b00000000; // 1643 :   0 - 0x0
      12'h66C: dout <= 8'b00000000; // 1644 :   0 - 0x0
      12'h66D: dout <= 8'b00000000; // 1645 :   0 - 0x0
      12'h66E: dout <= 8'b00000000; // 1646 :   0 - 0x0
      12'h66F: dout <= 8'b00000000; // 1647 :   0 - 0x0
      12'h670: dout <= 8'b00000000; // 1648 :   0 - 0x0 -- Background 0x67
      12'h671: dout <= 8'b00000000; // 1649 :   0 - 0x0
      12'h672: dout <= 8'b00000000; // 1650 :   0 - 0x0
      12'h673: dout <= 8'b00000000; // 1651 :   0 - 0x0
      12'h674: dout <= 8'b00000000; // 1652 :   0 - 0x0
      12'h675: dout <= 8'b00000000; // 1653 :   0 - 0x0
      12'h676: dout <= 8'b00000000; // 1654 :   0 - 0x0
      12'h677: dout <= 8'b00000000; // 1655 :   0 - 0x0
      12'h678: dout <= 8'b00000000; // 1656 :   0 - 0x0 -- plane 1
      12'h679: dout <= 8'b00000000; // 1657 :   0 - 0x0
      12'h67A: dout <= 8'b00000000; // 1658 :   0 - 0x0
      12'h67B: dout <= 8'b00000000; // 1659 :   0 - 0x0
      12'h67C: dout <= 8'b00000000; // 1660 :   0 - 0x0
      12'h67D: dout <= 8'b00000000; // 1661 :   0 - 0x0
      12'h67E: dout <= 8'b00000000; // 1662 :   0 - 0x0
      12'h67F: dout <= 8'b00000000; // 1663 :   0 - 0x0
      12'h680: dout <= 8'b00000000; // 1664 :   0 - 0x0 -- Background 0x68
      12'h681: dout <= 8'b00000000; // 1665 :   0 - 0x0
      12'h682: dout <= 8'b00000000; // 1666 :   0 - 0x0
      12'h683: dout <= 8'b00000000; // 1667 :   0 - 0x0
      12'h684: dout <= 8'b00000000; // 1668 :   0 - 0x0
      12'h685: dout <= 8'b00000000; // 1669 :   0 - 0x0
      12'h686: dout <= 8'b00000000; // 1670 :   0 - 0x0
      12'h687: dout <= 8'b00000000; // 1671 :   0 - 0x0
      12'h688: dout <= 8'b00000000; // 1672 :   0 - 0x0 -- plane 1
      12'h689: dout <= 8'b00000000; // 1673 :   0 - 0x0
      12'h68A: dout <= 8'b00000000; // 1674 :   0 - 0x0
      12'h68B: dout <= 8'b00000000; // 1675 :   0 - 0x0
      12'h68C: dout <= 8'b00000000; // 1676 :   0 - 0x0
      12'h68D: dout <= 8'b00000000; // 1677 :   0 - 0x0
      12'h68E: dout <= 8'b00000000; // 1678 :   0 - 0x0
      12'h68F: dout <= 8'b00000000; // 1679 :   0 - 0x0
      12'h690: dout <= 8'b00000000; // 1680 :   0 - 0x0 -- Background 0x69
      12'h691: dout <= 8'b00000000; // 1681 :   0 - 0x0
      12'h692: dout <= 8'b00000000; // 1682 :   0 - 0x0
      12'h693: dout <= 8'b00000000; // 1683 :   0 - 0x0
      12'h694: dout <= 8'b00000000; // 1684 :   0 - 0x0
      12'h695: dout <= 8'b00000000; // 1685 :   0 - 0x0
      12'h696: dout <= 8'b00000000; // 1686 :   0 - 0x0
      12'h697: dout <= 8'b00000000; // 1687 :   0 - 0x0
      12'h698: dout <= 8'b00000000; // 1688 :   0 - 0x0 -- plane 1
      12'h699: dout <= 8'b00000000; // 1689 :   0 - 0x0
      12'h69A: dout <= 8'b00000000; // 1690 :   0 - 0x0
      12'h69B: dout <= 8'b00000000; // 1691 :   0 - 0x0
      12'h69C: dout <= 8'b00000000; // 1692 :   0 - 0x0
      12'h69D: dout <= 8'b00000000; // 1693 :   0 - 0x0
      12'h69E: dout <= 8'b00000000; // 1694 :   0 - 0x0
      12'h69F: dout <= 8'b00000000; // 1695 :   0 - 0x0
      12'h6A0: dout <= 8'b00000000; // 1696 :   0 - 0x0 -- Background 0x6a
      12'h6A1: dout <= 8'b00000000; // 1697 :   0 - 0x0
      12'h6A2: dout <= 8'b00000000; // 1698 :   0 - 0x0
      12'h6A3: dout <= 8'b00000000; // 1699 :   0 - 0x0
      12'h6A4: dout <= 8'b00000000; // 1700 :   0 - 0x0
      12'h6A5: dout <= 8'b00000000; // 1701 :   0 - 0x0
      12'h6A6: dout <= 8'b00000000; // 1702 :   0 - 0x0
      12'h6A7: dout <= 8'b00000000; // 1703 :   0 - 0x0
      12'h6A8: dout <= 8'b00000000; // 1704 :   0 - 0x0 -- plane 1
      12'h6A9: dout <= 8'b00000000; // 1705 :   0 - 0x0
      12'h6AA: dout <= 8'b00000000; // 1706 :   0 - 0x0
      12'h6AB: dout <= 8'b00000000; // 1707 :   0 - 0x0
      12'h6AC: dout <= 8'b00000000; // 1708 :   0 - 0x0
      12'h6AD: dout <= 8'b00000000; // 1709 :   0 - 0x0
      12'h6AE: dout <= 8'b00000000; // 1710 :   0 - 0x0
      12'h6AF: dout <= 8'b00000000; // 1711 :   0 - 0x0
      12'h6B0: dout <= 8'b00000000; // 1712 :   0 - 0x0 -- Background 0x6b
      12'h6B1: dout <= 8'b00000000; // 1713 :   0 - 0x0
      12'h6B2: dout <= 8'b00000000; // 1714 :   0 - 0x0
      12'h6B3: dout <= 8'b00000000; // 1715 :   0 - 0x0
      12'h6B4: dout <= 8'b00000000; // 1716 :   0 - 0x0
      12'h6B5: dout <= 8'b00000000; // 1717 :   0 - 0x0
      12'h6B6: dout <= 8'b00000000; // 1718 :   0 - 0x0
      12'h6B7: dout <= 8'b00000000; // 1719 :   0 - 0x0
      12'h6B8: dout <= 8'b00000000; // 1720 :   0 - 0x0 -- plane 1
      12'h6B9: dout <= 8'b00000000; // 1721 :   0 - 0x0
      12'h6BA: dout <= 8'b00000000; // 1722 :   0 - 0x0
      12'h6BB: dout <= 8'b00000000; // 1723 :   0 - 0x0
      12'h6BC: dout <= 8'b00000000; // 1724 :   0 - 0x0
      12'h6BD: dout <= 8'b00000000; // 1725 :   0 - 0x0
      12'h6BE: dout <= 8'b00000000; // 1726 :   0 - 0x0
      12'h6BF: dout <= 8'b00000000; // 1727 :   0 - 0x0
      12'h6C0: dout <= 8'b00000000; // 1728 :   0 - 0x0 -- Background 0x6c
      12'h6C1: dout <= 8'b00000000; // 1729 :   0 - 0x0
      12'h6C2: dout <= 8'b00000000; // 1730 :   0 - 0x0
      12'h6C3: dout <= 8'b00000000; // 1731 :   0 - 0x0
      12'h6C4: dout <= 8'b00000000; // 1732 :   0 - 0x0
      12'h6C5: dout <= 8'b00000000; // 1733 :   0 - 0x0
      12'h6C6: dout <= 8'b00000000; // 1734 :   0 - 0x0
      12'h6C7: dout <= 8'b00000000; // 1735 :   0 - 0x0
      12'h6C8: dout <= 8'b00000000; // 1736 :   0 - 0x0 -- plane 1
      12'h6C9: dout <= 8'b00000000; // 1737 :   0 - 0x0
      12'h6CA: dout <= 8'b00000000; // 1738 :   0 - 0x0
      12'h6CB: dout <= 8'b00000000; // 1739 :   0 - 0x0
      12'h6CC: dout <= 8'b00000000; // 1740 :   0 - 0x0
      12'h6CD: dout <= 8'b00000000; // 1741 :   0 - 0x0
      12'h6CE: dout <= 8'b00000000; // 1742 :   0 - 0x0
      12'h6CF: dout <= 8'b00000000; // 1743 :   0 - 0x0
      12'h6D0: dout <= 8'b00000000; // 1744 :   0 - 0x0 -- Background 0x6d
      12'h6D1: dout <= 8'b00000000; // 1745 :   0 - 0x0
      12'h6D2: dout <= 8'b00000000; // 1746 :   0 - 0x0
      12'h6D3: dout <= 8'b00000000; // 1747 :   0 - 0x0
      12'h6D4: dout <= 8'b00000000; // 1748 :   0 - 0x0
      12'h6D5: dout <= 8'b00000000; // 1749 :   0 - 0x0
      12'h6D6: dout <= 8'b00000000; // 1750 :   0 - 0x0
      12'h6D7: dout <= 8'b00000000; // 1751 :   0 - 0x0
      12'h6D8: dout <= 8'b00000000; // 1752 :   0 - 0x0 -- plane 1
      12'h6D9: dout <= 8'b00000000; // 1753 :   0 - 0x0
      12'h6DA: dout <= 8'b00000000; // 1754 :   0 - 0x0
      12'h6DB: dout <= 8'b00000000; // 1755 :   0 - 0x0
      12'h6DC: dout <= 8'b00000000; // 1756 :   0 - 0x0
      12'h6DD: dout <= 8'b00000000; // 1757 :   0 - 0x0
      12'h6DE: dout <= 8'b00000000; // 1758 :   0 - 0x0
      12'h6DF: dout <= 8'b00000000; // 1759 :   0 - 0x0
      12'h6E0: dout <= 8'b00000000; // 1760 :   0 - 0x0 -- Background 0x6e
      12'h6E1: dout <= 8'b00000000; // 1761 :   0 - 0x0
      12'h6E2: dout <= 8'b00000000; // 1762 :   0 - 0x0
      12'h6E3: dout <= 8'b00000000; // 1763 :   0 - 0x0
      12'h6E4: dout <= 8'b00000000; // 1764 :   0 - 0x0
      12'h6E5: dout <= 8'b00000000; // 1765 :   0 - 0x0
      12'h6E6: dout <= 8'b00000000; // 1766 :   0 - 0x0
      12'h6E7: dout <= 8'b00000000; // 1767 :   0 - 0x0
      12'h6E8: dout <= 8'b00000000; // 1768 :   0 - 0x0 -- plane 1
      12'h6E9: dout <= 8'b00000000; // 1769 :   0 - 0x0
      12'h6EA: dout <= 8'b00000000; // 1770 :   0 - 0x0
      12'h6EB: dout <= 8'b00000000; // 1771 :   0 - 0x0
      12'h6EC: dout <= 8'b00000000; // 1772 :   0 - 0x0
      12'h6ED: dout <= 8'b00000000; // 1773 :   0 - 0x0
      12'h6EE: dout <= 8'b00000000; // 1774 :   0 - 0x0
      12'h6EF: dout <= 8'b00000000; // 1775 :   0 - 0x0
      12'h6F0: dout <= 8'b00000000; // 1776 :   0 - 0x0 -- Background 0x6f
      12'h6F1: dout <= 8'b00000000; // 1777 :   0 - 0x0
      12'h6F2: dout <= 8'b00000000; // 1778 :   0 - 0x0
      12'h6F3: dout <= 8'b00000000; // 1779 :   0 - 0x0
      12'h6F4: dout <= 8'b00000000; // 1780 :   0 - 0x0
      12'h6F5: dout <= 8'b00000000; // 1781 :   0 - 0x0
      12'h6F6: dout <= 8'b00000000; // 1782 :   0 - 0x0
      12'h6F7: dout <= 8'b00000000; // 1783 :   0 - 0x0
      12'h6F8: dout <= 8'b00000000; // 1784 :   0 - 0x0 -- plane 1
      12'h6F9: dout <= 8'b00000000; // 1785 :   0 - 0x0
      12'h6FA: dout <= 8'b00000000; // 1786 :   0 - 0x0
      12'h6FB: dout <= 8'b00000000; // 1787 :   0 - 0x0
      12'h6FC: dout <= 8'b00000000; // 1788 :   0 - 0x0
      12'h6FD: dout <= 8'b00000000; // 1789 :   0 - 0x0
      12'h6FE: dout <= 8'b00000000; // 1790 :   0 - 0x0
      12'h6FF: dout <= 8'b00000000; // 1791 :   0 - 0x0
      12'h700: dout <= 8'b00000000; // 1792 :   0 - 0x0 -- Background 0x70
      12'h701: dout <= 8'b00000000; // 1793 :   0 - 0x0
      12'h702: dout <= 8'b00000000; // 1794 :   0 - 0x0
      12'h703: dout <= 8'b00000000; // 1795 :   0 - 0x0
      12'h704: dout <= 8'b00000000; // 1796 :   0 - 0x0
      12'h705: dout <= 8'b00000000; // 1797 :   0 - 0x0
      12'h706: dout <= 8'b00000000; // 1798 :   0 - 0x0
      12'h707: dout <= 8'b00000000; // 1799 :   0 - 0x0
      12'h708: dout <= 8'b00000000; // 1800 :   0 - 0x0 -- plane 1
      12'h709: dout <= 8'b00000000; // 1801 :   0 - 0x0
      12'h70A: dout <= 8'b00000000; // 1802 :   0 - 0x0
      12'h70B: dout <= 8'b00000000; // 1803 :   0 - 0x0
      12'h70C: dout <= 8'b00000000; // 1804 :   0 - 0x0
      12'h70D: dout <= 8'b00000000; // 1805 :   0 - 0x0
      12'h70E: dout <= 8'b00000000; // 1806 :   0 - 0x0
      12'h70F: dout <= 8'b00000000; // 1807 :   0 - 0x0
      12'h710: dout <= 8'b00000000; // 1808 :   0 - 0x0 -- Background 0x71
      12'h711: dout <= 8'b00000000; // 1809 :   0 - 0x0
      12'h712: dout <= 8'b00000000; // 1810 :   0 - 0x0
      12'h713: dout <= 8'b00000000; // 1811 :   0 - 0x0
      12'h714: dout <= 8'b00000000; // 1812 :   0 - 0x0
      12'h715: dout <= 8'b00000000; // 1813 :   0 - 0x0
      12'h716: dout <= 8'b00000000; // 1814 :   0 - 0x0
      12'h717: dout <= 8'b00000000; // 1815 :   0 - 0x0
      12'h718: dout <= 8'b00000000; // 1816 :   0 - 0x0 -- plane 1
      12'h719: dout <= 8'b00000000; // 1817 :   0 - 0x0
      12'h71A: dout <= 8'b00000000; // 1818 :   0 - 0x0
      12'h71B: dout <= 8'b00000000; // 1819 :   0 - 0x0
      12'h71C: dout <= 8'b00000000; // 1820 :   0 - 0x0
      12'h71D: dout <= 8'b00000000; // 1821 :   0 - 0x0
      12'h71E: dout <= 8'b00000000; // 1822 :   0 - 0x0
      12'h71F: dout <= 8'b00000000; // 1823 :   0 - 0x0
      12'h720: dout <= 8'b00000000; // 1824 :   0 - 0x0 -- Background 0x72
      12'h721: dout <= 8'b00000000; // 1825 :   0 - 0x0
      12'h722: dout <= 8'b00000000; // 1826 :   0 - 0x0
      12'h723: dout <= 8'b00000000; // 1827 :   0 - 0x0
      12'h724: dout <= 8'b00000000; // 1828 :   0 - 0x0
      12'h725: dout <= 8'b00000000; // 1829 :   0 - 0x0
      12'h726: dout <= 8'b00000000; // 1830 :   0 - 0x0
      12'h727: dout <= 8'b00000000; // 1831 :   0 - 0x0
      12'h728: dout <= 8'b00000000; // 1832 :   0 - 0x0 -- plane 1
      12'h729: dout <= 8'b00000000; // 1833 :   0 - 0x0
      12'h72A: dout <= 8'b00000000; // 1834 :   0 - 0x0
      12'h72B: dout <= 8'b00000000; // 1835 :   0 - 0x0
      12'h72C: dout <= 8'b00000000; // 1836 :   0 - 0x0
      12'h72D: dout <= 8'b00000000; // 1837 :   0 - 0x0
      12'h72E: dout <= 8'b00000000; // 1838 :   0 - 0x0
      12'h72F: dout <= 8'b00000000; // 1839 :   0 - 0x0
      12'h730: dout <= 8'b00000000; // 1840 :   0 - 0x0 -- Background 0x73
      12'h731: dout <= 8'b00000000; // 1841 :   0 - 0x0
      12'h732: dout <= 8'b00000000; // 1842 :   0 - 0x0
      12'h733: dout <= 8'b00000000; // 1843 :   0 - 0x0
      12'h734: dout <= 8'b00000000; // 1844 :   0 - 0x0
      12'h735: dout <= 8'b00000000; // 1845 :   0 - 0x0
      12'h736: dout <= 8'b00000000; // 1846 :   0 - 0x0
      12'h737: dout <= 8'b00000000; // 1847 :   0 - 0x0
      12'h738: dout <= 8'b00000000; // 1848 :   0 - 0x0 -- plane 1
      12'h739: dout <= 8'b00000000; // 1849 :   0 - 0x0
      12'h73A: dout <= 8'b00000000; // 1850 :   0 - 0x0
      12'h73B: dout <= 8'b00000000; // 1851 :   0 - 0x0
      12'h73C: dout <= 8'b00000000; // 1852 :   0 - 0x0
      12'h73D: dout <= 8'b00000000; // 1853 :   0 - 0x0
      12'h73E: dout <= 8'b00000000; // 1854 :   0 - 0x0
      12'h73F: dout <= 8'b00000000; // 1855 :   0 - 0x0
      12'h740: dout <= 8'b00000000; // 1856 :   0 - 0x0 -- Background 0x74
      12'h741: dout <= 8'b00000000; // 1857 :   0 - 0x0
      12'h742: dout <= 8'b00000000; // 1858 :   0 - 0x0
      12'h743: dout <= 8'b00000000; // 1859 :   0 - 0x0
      12'h744: dout <= 8'b00000000; // 1860 :   0 - 0x0
      12'h745: dout <= 8'b00000000; // 1861 :   0 - 0x0
      12'h746: dout <= 8'b00000000; // 1862 :   0 - 0x0
      12'h747: dout <= 8'b00000000; // 1863 :   0 - 0x0
      12'h748: dout <= 8'b00000000; // 1864 :   0 - 0x0 -- plane 1
      12'h749: dout <= 8'b00000000; // 1865 :   0 - 0x0
      12'h74A: dout <= 8'b00000000; // 1866 :   0 - 0x0
      12'h74B: dout <= 8'b00000000; // 1867 :   0 - 0x0
      12'h74C: dout <= 8'b00000000; // 1868 :   0 - 0x0
      12'h74D: dout <= 8'b00000000; // 1869 :   0 - 0x0
      12'h74E: dout <= 8'b00000000; // 1870 :   0 - 0x0
      12'h74F: dout <= 8'b00000000; // 1871 :   0 - 0x0
      12'h750: dout <= 8'b00000000; // 1872 :   0 - 0x0 -- Background 0x75
      12'h751: dout <= 8'b00000000; // 1873 :   0 - 0x0
      12'h752: dout <= 8'b00000000; // 1874 :   0 - 0x0
      12'h753: dout <= 8'b00000000; // 1875 :   0 - 0x0
      12'h754: dout <= 8'b00000000; // 1876 :   0 - 0x0
      12'h755: dout <= 8'b00000000; // 1877 :   0 - 0x0
      12'h756: dout <= 8'b00000000; // 1878 :   0 - 0x0
      12'h757: dout <= 8'b00000000; // 1879 :   0 - 0x0
      12'h758: dout <= 8'b00000000; // 1880 :   0 - 0x0 -- plane 1
      12'h759: dout <= 8'b00000000; // 1881 :   0 - 0x0
      12'h75A: dout <= 8'b00000000; // 1882 :   0 - 0x0
      12'h75B: dout <= 8'b00000000; // 1883 :   0 - 0x0
      12'h75C: dout <= 8'b00000000; // 1884 :   0 - 0x0
      12'h75D: dout <= 8'b00000000; // 1885 :   0 - 0x0
      12'h75E: dout <= 8'b00000000; // 1886 :   0 - 0x0
      12'h75F: dout <= 8'b00000000; // 1887 :   0 - 0x0
      12'h760: dout <= 8'b00000000; // 1888 :   0 - 0x0 -- Background 0x76
      12'h761: dout <= 8'b00000000; // 1889 :   0 - 0x0
      12'h762: dout <= 8'b00000000; // 1890 :   0 - 0x0
      12'h763: dout <= 8'b00000000; // 1891 :   0 - 0x0
      12'h764: dout <= 8'b00000000; // 1892 :   0 - 0x0
      12'h765: dout <= 8'b00000000; // 1893 :   0 - 0x0
      12'h766: dout <= 8'b00000000; // 1894 :   0 - 0x0
      12'h767: dout <= 8'b00000000; // 1895 :   0 - 0x0
      12'h768: dout <= 8'b00000000; // 1896 :   0 - 0x0 -- plane 1
      12'h769: dout <= 8'b00000000; // 1897 :   0 - 0x0
      12'h76A: dout <= 8'b00000000; // 1898 :   0 - 0x0
      12'h76B: dout <= 8'b00000000; // 1899 :   0 - 0x0
      12'h76C: dout <= 8'b00000000; // 1900 :   0 - 0x0
      12'h76D: dout <= 8'b00000000; // 1901 :   0 - 0x0
      12'h76E: dout <= 8'b00000000; // 1902 :   0 - 0x0
      12'h76F: dout <= 8'b00000000; // 1903 :   0 - 0x0
      12'h770: dout <= 8'b00000000; // 1904 :   0 - 0x0 -- Background 0x77
      12'h771: dout <= 8'b00000000; // 1905 :   0 - 0x0
      12'h772: dout <= 8'b00000000; // 1906 :   0 - 0x0
      12'h773: dout <= 8'b00000000; // 1907 :   0 - 0x0
      12'h774: dout <= 8'b00000000; // 1908 :   0 - 0x0
      12'h775: dout <= 8'b00000000; // 1909 :   0 - 0x0
      12'h776: dout <= 8'b00000000; // 1910 :   0 - 0x0
      12'h777: dout <= 8'b00000000; // 1911 :   0 - 0x0
      12'h778: dout <= 8'b00000000; // 1912 :   0 - 0x0 -- plane 1
      12'h779: dout <= 8'b00000000; // 1913 :   0 - 0x0
      12'h77A: dout <= 8'b00000000; // 1914 :   0 - 0x0
      12'h77B: dout <= 8'b00000000; // 1915 :   0 - 0x0
      12'h77C: dout <= 8'b00000000; // 1916 :   0 - 0x0
      12'h77D: dout <= 8'b00000000; // 1917 :   0 - 0x0
      12'h77E: dout <= 8'b00000000; // 1918 :   0 - 0x0
      12'h77F: dout <= 8'b00000000; // 1919 :   0 - 0x0
      12'h780: dout <= 8'b00000000; // 1920 :   0 - 0x0 -- Background 0x78
      12'h781: dout <= 8'b00000000; // 1921 :   0 - 0x0
      12'h782: dout <= 8'b00000000; // 1922 :   0 - 0x0
      12'h783: dout <= 8'b00000000; // 1923 :   0 - 0x0
      12'h784: dout <= 8'b00000000; // 1924 :   0 - 0x0
      12'h785: dout <= 8'b00000000; // 1925 :   0 - 0x0
      12'h786: dout <= 8'b00000000; // 1926 :   0 - 0x0
      12'h787: dout <= 8'b00000000; // 1927 :   0 - 0x0
      12'h788: dout <= 8'b00000000; // 1928 :   0 - 0x0 -- plane 1
      12'h789: dout <= 8'b00000000; // 1929 :   0 - 0x0
      12'h78A: dout <= 8'b00000000; // 1930 :   0 - 0x0
      12'h78B: dout <= 8'b00000000; // 1931 :   0 - 0x0
      12'h78C: dout <= 8'b00000000; // 1932 :   0 - 0x0
      12'h78D: dout <= 8'b00000000; // 1933 :   0 - 0x0
      12'h78E: dout <= 8'b00000000; // 1934 :   0 - 0x0
      12'h78F: dout <= 8'b00000000; // 1935 :   0 - 0x0
      12'h790: dout <= 8'b00000000; // 1936 :   0 - 0x0 -- Background 0x79
      12'h791: dout <= 8'b00000000; // 1937 :   0 - 0x0
      12'h792: dout <= 8'b00000000; // 1938 :   0 - 0x0
      12'h793: dout <= 8'b00000000; // 1939 :   0 - 0x0
      12'h794: dout <= 8'b00000000; // 1940 :   0 - 0x0
      12'h795: dout <= 8'b00000000; // 1941 :   0 - 0x0
      12'h796: dout <= 8'b00000000; // 1942 :   0 - 0x0
      12'h797: dout <= 8'b00000000; // 1943 :   0 - 0x0
      12'h798: dout <= 8'b00000000; // 1944 :   0 - 0x0 -- plane 1
      12'h799: dout <= 8'b00000000; // 1945 :   0 - 0x0
      12'h79A: dout <= 8'b00000000; // 1946 :   0 - 0x0
      12'h79B: dout <= 8'b00000000; // 1947 :   0 - 0x0
      12'h79C: dout <= 8'b00000000; // 1948 :   0 - 0x0
      12'h79D: dout <= 8'b00000000; // 1949 :   0 - 0x0
      12'h79E: dout <= 8'b00000000; // 1950 :   0 - 0x0
      12'h79F: dout <= 8'b00000000; // 1951 :   0 - 0x0
      12'h7A0: dout <= 8'b00000000; // 1952 :   0 - 0x0 -- Background 0x7a
      12'h7A1: dout <= 8'b00000000; // 1953 :   0 - 0x0
      12'h7A2: dout <= 8'b00000000; // 1954 :   0 - 0x0
      12'h7A3: dout <= 8'b00000000; // 1955 :   0 - 0x0
      12'h7A4: dout <= 8'b00000000; // 1956 :   0 - 0x0
      12'h7A5: dout <= 8'b00000000; // 1957 :   0 - 0x0
      12'h7A6: dout <= 8'b00000000; // 1958 :   0 - 0x0
      12'h7A7: dout <= 8'b00000000; // 1959 :   0 - 0x0
      12'h7A8: dout <= 8'b00000000; // 1960 :   0 - 0x0 -- plane 1
      12'h7A9: dout <= 8'b00000000; // 1961 :   0 - 0x0
      12'h7AA: dout <= 8'b00000000; // 1962 :   0 - 0x0
      12'h7AB: dout <= 8'b00000000; // 1963 :   0 - 0x0
      12'h7AC: dout <= 8'b00000000; // 1964 :   0 - 0x0
      12'h7AD: dout <= 8'b00000000; // 1965 :   0 - 0x0
      12'h7AE: dout <= 8'b00000000; // 1966 :   0 - 0x0
      12'h7AF: dout <= 8'b00000000; // 1967 :   0 - 0x0
      12'h7B0: dout <= 8'b00000000; // 1968 :   0 - 0x0 -- Background 0x7b
      12'h7B1: dout <= 8'b00000000; // 1969 :   0 - 0x0
      12'h7B2: dout <= 8'b00000000; // 1970 :   0 - 0x0
      12'h7B3: dout <= 8'b00000000; // 1971 :   0 - 0x0
      12'h7B4: dout <= 8'b00000000; // 1972 :   0 - 0x0
      12'h7B5: dout <= 8'b00000000; // 1973 :   0 - 0x0
      12'h7B6: dout <= 8'b00000000; // 1974 :   0 - 0x0
      12'h7B7: dout <= 8'b00000000; // 1975 :   0 - 0x0
      12'h7B8: dout <= 8'b00000000; // 1976 :   0 - 0x0 -- plane 1
      12'h7B9: dout <= 8'b00000000; // 1977 :   0 - 0x0
      12'h7BA: dout <= 8'b00000000; // 1978 :   0 - 0x0
      12'h7BB: dout <= 8'b00000000; // 1979 :   0 - 0x0
      12'h7BC: dout <= 8'b00000000; // 1980 :   0 - 0x0
      12'h7BD: dout <= 8'b00000000; // 1981 :   0 - 0x0
      12'h7BE: dout <= 8'b00000000; // 1982 :   0 - 0x0
      12'h7BF: dout <= 8'b00000000; // 1983 :   0 - 0x0
      12'h7C0: dout <= 8'b00000000; // 1984 :   0 - 0x0 -- Background 0x7c
      12'h7C1: dout <= 8'b00000000; // 1985 :   0 - 0x0
      12'h7C2: dout <= 8'b00000000; // 1986 :   0 - 0x0
      12'h7C3: dout <= 8'b00000000; // 1987 :   0 - 0x0
      12'h7C4: dout <= 8'b00000000; // 1988 :   0 - 0x0
      12'h7C5: dout <= 8'b00000000; // 1989 :   0 - 0x0
      12'h7C6: dout <= 8'b00000000; // 1990 :   0 - 0x0
      12'h7C7: dout <= 8'b00000000; // 1991 :   0 - 0x0
      12'h7C8: dout <= 8'b00000000; // 1992 :   0 - 0x0 -- plane 1
      12'h7C9: dout <= 8'b00000000; // 1993 :   0 - 0x0
      12'h7CA: dout <= 8'b00000000; // 1994 :   0 - 0x0
      12'h7CB: dout <= 8'b00000000; // 1995 :   0 - 0x0
      12'h7CC: dout <= 8'b00000000; // 1996 :   0 - 0x0
      12'h7CD: dout <= 8'b00000000; // 1997 :   0 - 0x0
      12'h7CE: dout <= 8'b00000000; // 1998 :   0 - 0x0
      12'h7CF: dout <= 8'b00000000; // 1999 :   0 - 0x0
      12'h7D0: dout <= 8'b00000000; // 2000 :   0 - 0x0 -- Background 0x7d
      12'h7D1: dout <= 8'b00000000; // 2001 :   0 - 0x0
      12'h7D2: dout <= 8'b00000000; // 2002 :   0 - 0x0
      12'h7D3: dout <= 8'b00000000; // 2003 :   0 - 0x0
      12'h7D4: dout <= 8'b00000000; // 2004 :   0 - 0x0
      12'h7D5: dout <= 8'b00000000; // 2005 :   0 - 0x0
      12'h7D6: dout <= 8'b00000000; // 2006 :   0 - 0x0
      12'h7D7: dout <= 8'b00000000; // 2007 :   0 - 0x0
      12'h7D8: dout <= 8'b00000000; // 2008 :   0 - 0x0 -- plane 1
      12'h7D9: dout <= 8'b00000000; // 2009 :   0 - 0x0
      12'h7DA: dout <= 8'b00000000; // 2010 :   0 - 0x0
      12'h7DB: dout <= 8'b00000000; // 2011 :   0 - 0x0
      12'h7DC: dout <= 8'b00000000; // 2012 :   0 - 0x0
      12'h7DD: dout <= 8'b00000000; // 2013 :   0 - 0x0
      12'h7DE: dout <= 8'b00000000; // 2014 :   0 - 0x0
      12'h7DF: dout <= 8'b00000000; // 2015 :   0 - 0x0
      12'h7E0: dout <= 8'b00000000; // 2016 :   0 - 0x0 -- Background 0x7e
      12'h7E1: dout <= 8'b00000000; // 2017 :   0 - 0x0
      12'h7E2: dout <= 8'b00000000; // 2018 :   0 - 0x0
      12'h7E3: dout <= 8'b00000000; // 2019 :   0 - 0x0
      12'h7E4: dout <= 8'b00000000; // 2020 :   0 - 0x0
      12'h7E5: dout <= 8'b00000000; // 2021 :   0 - 0x0
      12'h7E6: dout <= 8'b00000000; // 2022 :   0 - 0x0
      12'h7E7: dout <= 8'b00000000; // 2023 :   0 - 0x0
      12'h7E8: dout <= 8'b00000000; // 2024 :   0 - 0x0 -- plane 1
      12'h7E9: dout <= 8'b00000000; // 2025 :   0 - 0x0
      12'h7EA: dout <= 8'b00000000; // 2026 :   0 - 0x0
      12'h7EB: dout <= 8'b00000000; // 2027 :   0 - 0x0
      12'h7EC: dout <= 8'b00000000; // 2028 :   0 - 0x0
      12'h7ED: dout <= 8'b00000000; // 2029 :   0 - 0x0
      12'h7EE: dout <= 8'b00000000; // 2030 :   0 - 0x0
      12'h7EF: dout <= 8'b00000000; // 2031 :   0 - 0x0
      12'h7F0: dout <= 8'b00000000; // 2032 :   0 - 0x0 -- Background 0x7f
      12'h7F1: dout <= 8'b00000000; // 2033 :   0 - 0x0
      12'h7F2: dout <= 8'b00000000; // 2034 :   0 - 0x0
      12'h7F3: dout <= 8'b00000000; // 2035 :   0 - 0x0
      12'h7F4: dout <= 8'b00000000; // 2036 :   0 - 0x0
      12'h7F5: dout <= 8'b00000000; // 2037 :   0 - 0x0
      12'h7F6: dout <= 8'b00000000; // 2038 :   0 - 0x0
      12'h7F7: dout <= 8'b00000000; // 2039 :   0 - 0x0
      12'h7F8: dout <= 8'b00000000; // 2040 :   0 - 0x0 -- plane 1
      12'h7F9: dout <= 8'b00000000; // 2041 :   0 - 0x0
      12'h7FA: dout <= 8'b00000000; // 2042 :   0 - 0x0
      12'h7FB: dout <= 8'b00000000; // 2043 :   0 - 0x0
      12'h7FC: dout <= 8'b00000000; // 2044 :   0 - 0x0
      12'h7FD: dout <= 8'b00000000; // 2045 :   0 - 0x0
      12'h7FE: dout <= 8'b00000000; // 2046 :   0 - 0x0
      12'h7FF: dout <= 8'b00000000; // 2047 :   0 - 0x0
      12'h800: dout <= 8'b00000000; // 2048 :   0 - 0x0 -- Background 0x80
      12'h801: dout <= 8'b00000000; // 2049 :   0 - 0x0
      12'h802: dout <= 8'b00000000; // 2050 :   0 - 0x0
      12'h803: dout <= 8'b00000000; // 2051 :   0 - 0x0
      12'h804: dout <= 8'b00000000; // 2052 :   0 - 0x0
      12'h805: dout <= 8'b00000000; // 2053 :   0 - 0x0
      12'h806: dout <= 8'b00000000; // 2054 :   0 - 0x0
      12'h807: dout <= 8'b00000000; // 2055 :   0 - 0x0
      12'h808: dout <= 8'b00000000; // 2056 :   0 - 0x0 -- plane 1
      12'h809: dout <= 8'b00000000; // 2057 :   0 - 0x0
      12'h80A: dout <= 8'b00000000; // 2058 :   0 - 0x0
      12'h80B: dout <= 8'b00000000; // 2059 :   0 - 0x0
      12'h80C: dout <= 8'b00000000; // 2060 :   0 - 0x0
      12'h80D: dout <= 8'b00000000; // 2061 :   0 - 0x0
      12'h80E: dout <= 8'b00000000; // 2062 :   0 - 0x0
      12'h80F: dout <= 8'b00000000; // 2063 :   0 - 0x0
      12'h810: dout <= 8'b00000000; // 2064 :   0 - 0x0 -- Background 0x81
      12'h811: dout <= 8'b00000000; // 2065 :   0 - 0x0
      12'h812: dout <= 8'b00000000; // 2066 :   0 - 0x0
      12'h813: dout <= 8'b00000000; // 2067 :   0 - 0x0
      12'h814: dout <= 8'b00000000; // 2068 :   0 - 0x0
      12'h815: dout <= 8'b00000000; // 2069 :   0 - 0x0
      12'h816: dout <= 8'b00000000; // 2070 :   0 - 0x0
      12'h817: dout <= 8'b00000000; // 2071 :   0 - 0x0
      12'h818: dout <= 8'b00000000; // 2072 :   0 - 0x0 -- plane 1
      12'h819: dout <= 8'b00000000; // 2073 :   0 - 0x0
      12'h81A: dout <= 8'b00000000; // 2074 :   0 - 0x0
      12'h81B: dout <= 8'b00000000; // 2075 :   0 - 0x0
      12'h81C: dout <= 8'b00000000; // 2076 :   0 - 0x0
      12'h81D: dout <= 8'b00000000; // 2077 :   0 - 0x0
      12'h81E: dout <= 8'b00000000; // 2078 :   0 - 0x0
      12'h81F: dout <= 8'b00000000; // 2079 :   0 - 0x0
      12'h820: dout <= 8'b00000000; // 2080 :   0 - 0x0 -- Background 0x82
      12'h821: dout <= 8'b00000000; // 2081 :   0 - 0x0
      12'h822: dout <= 8'b00000000; // 2082 :   0 - 0x0
      12'h823: dout <= 8'b00000000; // 2083 :   0 - 0x0
      12'h824: dout <= 8'b00000000; // 2084 :   0 - 0x0
      12'h825: dout <= 8'b00000000; // 2085 :   0 - 0x0
      12'h826: dout <= 8'b00000000; // 2086 :   0 - 0x0
      12'h827: dout <= 8'b00000000; // 2087 :   0 - 0x0
      12'h828: dout <= 8'b00000000; // 2088 :   0 - 0x0 -- plane 1
      12'h829: dout <= 8'b00000000; // 2089 :   0 - 0x0
      12'h82A: dout <= 8'b00000000; // 2090 :   0 - 0x0
      12'h82B: dout <= 8'b00000000; // 2091 :   0 - 0x0
      12'h82C: dout <= 8'b00000000; // 2092 :   0 - 0x0
      12'h82D: dout <= 8'b00000000; // 2093 :   0 - 0x0
      12'h82E: dout <= 8'b00000000; // 2094 :   0 - 0x0
      12'h82F: dout <= 8'b00000000; // 2095 :   0 - 0x0
      12'h830: dout <= 8'b00000000; // 2096 :   0 - 0x0 -- Background 0x83
      12'h831: dout <= 8'b00000000; // 2097 :   0 - 0x0
      12'h832: dout <= 8'b00000000; // 2098 :   0 - 0x0
      12'h833: dout <= 8'b00000000; // 2099 :   0 - 0x0
      12'h834: dout <= 8'b00000000; // 2100 :   0 - 0x0
      12'h835: dout <= 8'b00000000; // 2101 :   0 - 0x0
      12'h836: dout <= 8'b00000000; // 2102 :   0 - 0x0
      12'h837: dout <= 8'b00000000; // 2103 :   0 - 0x0
      12'h838: dout <= 8'b00000000; // 2104 :   0 - 0x0 -- plane 1
      12'h839: dout <= 8'b00000000; // 2105 :   0 - 0x0
      12'h83A: dout <= 8'b00000000; // 2106 :   0 - 0x0
      12'h83B: dout <= 8'b00000000; // 2107 :   0 - 0x0
      12'h83C: dout <= 8'b00000000; // 2108 :   0 - 0x0
      12'h83D: dout <= 8'b00000000; // 2109 :   0 - 0x0
      12'h83E: dout <= 8'b00000000; // 2110 :   0 - 0x0
      12'h83F: dout <= 8'b00000000; // 2111 :   0 - 0x0
      12'h840: dout <= 8'b00000000; // 2112 :   0 - 0x0 -- Background 0x84
      12'h841: dout <= 8'b00000000; // 2113 :   0 - 0x0
      12'h842: dout <= 8'b00000000; // 2114 :   0 - 0x0
      12'h843: dout <= 8'b00000000; // 2115 :   0 - 0x0
      12'h844: dout <= 8'b00000000; // 2116 :   0 - 0x0
      12'h845: dout <= 8'b00000000; // 2117 :   0 - 0x0
      12'h846: dout <= 8'b00000000; // 2118 :   0 - 0x0
      12'h847: dout <= 8'b00000000; // 2119 :   0 - 0x0
      12'h848: dout <= 8'b00000000; // 2120 :   0 - 0x0 -- plane 1
      12'h849: dout <= 8'b00000000; // 2121 :   0 - 0x0
      12'h84A: dout <= 8'b00000000; // 2122 :   0 - 0x0
      12'h84B: dout <= 8'b00000000; // 2123 :   0 - 0x0
      12'h84C: dout <= 8'b00000000; // 2124 :   0 - 0x0
      12'h84D: dout <= 8'b00000000; // 2125 :   0 - 0x0
      12'h84E: dout <= 8'b00000000; // 2126 :   0 - 0x0
      12'h84F: dout <= 8'b00000000; // 2127 :   0 - 0x0
      12'h850: dout <= 8'b00000000; // 2128 :   0 - 0x0 -- Background 0x85
      12'h851: dout <= 8'b00000000; // 2129 :   0 - 0x0
      12'h852: dout <= 8'b00000000; // 2130 :   0 - 0x0
      12'h853: dout <= 8'b00000000; // 2131 :   0 - 0x0
      12'h854: dout <= 8'b00000000; // 2132 :   0 - 0x0
      12'h855: dout <= 8'b00000000; // 2133 :   0 - 0x0
      12'h856: dout <= 8'b00000000; // 2134 :   0 - 0x0
      12'h857: dout <= 8'b00000000; // 2135 :   0 - 0x0
      12'h858: dout <= 8'b00000000; // 2136 :   0 - 0x0 -- plane 1
      12'h859: dout <= 8'b00000000; // 2137 :   0 - 0x0
      12'h85A: dout <= 8'b00000000; // 2138 :   0 - 0x0
      12'h85B: dout <= 8'b00000000; // 2139 :   0 - 0x0
      12'h85C: dout <= 8'b00000000; // 2140 :   0 - 0x0
      12'h85D: dout <= 8'b00000000; // 2141 :   0 - 0x0
      12'h85E: dout <= 8'b00000000; // 2142 :   0 - 0x0
      12'h85F: dout <= 8'b00000000; // 2143 :   0 - 0x0
      12'h860: dout <= 8'b00000000; // 2144 :   0 - 0x0 -- Background 0x86
      12'h861: dout <= 8'b00000000; // 2145 :   0 - 0x0
      12'h862: dout <= 8'b00000000; // 2146 :   0 - 0x0
      12'h863: dout <= 8'b00000000; // 2147 :   0 - 0x0
      12'h864: dout <= 8'b00000000; // 2148 :   0 - 0x0
      12'h865: dout <= 8'b00000000; // 2149 :   0 - 0x0
      12'h866: dout <= 8'b00000000; // 2150 :   0 - 0x0
      12'h867: dout <= 8'b00000000; // 2151 :   0 - 0x0
      12'h868: dout <= 8'b00000000; // 2152 :   0 - 0x0 -- plane 1
      12'h869: dout <= 8'b00000000; // 2153 :   0 - 0x0
      12'h86A: dout <= 8'b00000000; // 2154 :   0 - 0x0
      12'h86B: dout <= 8'b00000000; // 2155 :   0 - 0x0
      12'h86C: dout <= 8'b00000000; // 2156 :   0 - 0x0
      12'h86D: dout <= 8'b00000000; // 2157 :   0 - 0x0
      12'h86E: dout <= 8'b00000000; // 2158 :   0 - 0x0
      12'h86F: dout <= 8'b00000000; // 2159 :   0 - 0x0
      12'h870: dout <= 8'b00000000; // 2160 :   0 - 0x0 -- Background 0x87
      12'h871: dout <= 8'b00000000; // 2161 :   0 - 0x0
      12'h872: dout <= 8'b00000000; // 2162 :   0 - 0x0
      12'h873: dout <= 8'b00000000; // 2163 :   0 - 0x0
      12'h874: dout <= 8'b00000000; // 2164 :   0 - 0x0
      12'h875: dout <= 8'b00000000; // 2165 :   0 - 0x0
      12'h876: dout <= 8'b00000000; // 2166 :   0 - 0x0
      12'h877: dout <= 8'b00000000; // 2167 :   0 - 0x0
      12'h878: dout <= 8'b00000000; // 2168 :   0 - 0x0 -- plane 1
      12'h879: dout <= 8'b00000000; // 2169 :   0 - 0x0
      12'h87A: dout <= 8'b00000000; // 2170 :   0 - 0x0
      12'h87B: dout <= 8'b00000000; // 2171 :   0 - 0x0
      12'h87C: dout <= 8'b00000000; // 2172 :   0 - 0x0
      12'h87D: dout <= 8'b00000000; // 2173 :   0 - 0x0
      12'h87E: dout <= 8'b00000000; // 2174 :   0 - 0x0
      12'h87F: dout <= 8'b00000000; // 2175 :   0 - 0x0
      12'h880: dout <= 8'b00000000; // 2176 :   0 - 0x0 -- Background 0x88
      12'h881: dout <= 8'b00000000; // 2177 :   0 - 0x0
      12'h882: dout <= 8'b00000000; // 2178 :   0 - 0x0
      12'h883: dout <= 8'b00000000; // 2179 :   0 - 0x0
      12'h884: dout <= 8'b00000000; // 2180 :   0 - 0x0
      12'h885: dout <= 8'b00000000; // 2181 :   0 - 0x0
      12'h886: dout <= 8'b00000000; // 2182 :   0 - 0x0
      12'h887: dout <= 8'b00000000; // 2183 :   0 - 0x0
      12'h888: dout <= 8'b00000000; // 2184 :   0 - 0x0 -- plane 1
      12'h889: dout <= 8'b00000000; // 2185 :   0 - 0x0
      12'h88A: dout <= 8'b00000000; // 2186 :   0 - 0x0
      12'h88B: dout <= 8'b00000000; // 2187 :   0 - 0x0
      12'h88C: dout <= 8'b00000000; // 2188 :   0 - 0x0
      12'h88D: dout <= 8'b00000000; // 2189 :   0 - 0x0
      12'h88E: dout <= 8'b00000000; // 2190 :   0 - 0x0
      12'h88F: dout <= 8'b00000000; // 2191 :   0 - 0x0
      12'h890: dout <= 8'b00000000; // 2192 :   0 - 0x0 -- Background 0x89
      12'h891: dout <= 8'b00000000; // 2193 :   0 - 0x0
      12'h892: dout <= 8'b00000000; // 2194 :   0 - 0x0
      12'h893: dout <= 8'b00000000; // 2195 :   0 - 0x0
      12'h894: dout <= 8'b00000000; // 2196 :   0 - 0x0
      12'h895: dout <= 8'b00000000; // 2197 :   0 - 0x0
      12'h896: dout <= 8'b00000000; // 2198 :   0 - 0x0
      12'h897: dout <= 8'b00000000; // 2199 :   0 - 0x0
      12'h898: dout <= 8'b00000000; // 2200 :   0 - 0x0 -- plane 1
      12'h899: dout <= 8'b00000000; // 2201 :   0 - 0x0
      12'h89A: dout <= 8'b00000000; // 2202 :   0 - 0x0
      12'h89B: dout <= 8'b00000000; // 2203 :   0 - 0x0
      12'h89C: dout <= 8'b00000000; // 2204 :   0 - 0x0
      12'h89D: dout <= 8'b00000000; // 2205 :   0 - 0x0
      12'h89E: dout <= 8'b00000000; // 2206 :   0 - 0x0
      12'h89F: dout <= 8'b00000000; // 2207 :   0 - 0x0
      12'h8A0: dout <= 8'b00000000; // 2208 :   0 - 0x0 -- Background 0x8a
      12'h8A1: dout <= 8'b00000000; // 2209 :   0 - 0x0
      12'h8A2: dout <= 8'b00000000; // 2210 :   0 - 0x0
      12'h8A3: dout <= 8'b00000000; // 2211 :   0 - 0x0
      12'h8A4: dout <= 8'b00000000; // 2212 :   0 - 0x0
      12'h8A5: dout <= 8'b00000000; // 2213 :   0 - 0x0
      12'h8A6: dout <= 8'b00000000; // 2214 :   0 - 0x0
      12'h8A7: dout <= 8'b00000000; // 2215 :   0 - 0x0
      12'h8A8: dout <= 8'b00000000; // 2216 :   0 - 0x0 -- plane 1
      12'h8A9: dout <= 8'b00000000; // 2217 :   0 - 0x0
      12'h8AA: dout <= 8'b00000000; // 2218 :   0 - 0x0
      12'h8AB: dout <= 8'b00000000; // 2219 :   0 - 0x0
      12'h8AC: dout <= 8'b00000000; // 2220 :   0 - 0x0
      12'h8AD: dout <= 8'b00000000; // 2221 :   0 - 0x0
      12'h8AE: dout <= 8'b00000000; // 2222 :   0 - 0x0
      12'h8AF: dout <= 8'b00000000; // 2223 :   0 - 0x0
      12'h8B0: dout <= 8'b00000000; // 2224 :   0 - 0x0 -- Background 0x8b
      12'h8B1: dout <= 8'b00000000; // 2225 :   0 - 0x0
      12'h8B2: dout <= 8'b00000000; // 2226 :   0 - 0x0
      12'h8B3: dout <= 8'b00000000; // 2227 :   0 - 0x0
      12'h8B4: dout <= 8'b00000000; // 2228 :   0 - 0x0
      12'h8B5: dout <= 8'b00000000; // 2229 :   0 - 0x0
      12'h8B6: dout <= 8'b00000000; // 2230 :   0 - 0x0
      12'h8B7: dout <= 8'b00000000; // 2231 :   0 - 0x0
      12'h8B8: dout <= 8'b00000000; // 2232 :   0 - 0x0 -- plane 1
      12'h8B9: dout <= 8'b00000000; // 2233 :   0 - 0x0
      12'h8BA: dout <= 8'b00000000; // 2234 :   0 - 0x0
      12'h8BB: dout <= 8'b00000000; // 2235 :   0 - 0x0
      12'h8BC: dout <= 8'b00000000; // 2236 :   0 - 0x0
      12'h8BD: dout <= 8'b00000000; // 2237 :   0 - 0x0
      12'h8BE: dout <= 8'b00000000; // 2238 :   0 - 0x0
      12'h8BF: dout <= 8'b00000000; // 2239 :   0 - 0x0
      12'h8C0: dout <= 8'b00000000; // 2240 :   0 - 0x0 -- Background 0x8c
      12'h8C1: dout <= 8'b00000000; // 2241 :   0 - 0x0
      12'h8C2: dout <= 8'b00000000; // 2242 :   0 - 0x0
      12'h8C3: dout <= 8'b00000000; // 2243 :   0 - 0x0
      12'h8C4: dout <= 8'b00000000; // 2244 :   0 - 0x0
      12'h8C5: dout <= 8'b00000000; // 2245 :   0 - 0x0
      12'h8C6: dout <= 8'b00000000; // 2246 :   0 - 0x0
      12'h8C7: dout <= 8'b00000000; // 2247 :   0 - 0x0
      12'h8C8: dout <= 8'b00000000; // 2248 :   0 - 0x0 -- plane 1
      12'h8C9: dout <= 8'b00000000; // 2249 :   0 - 0x0
      12'h8CA: dout <= 8'b00000000; // 2250 :   0 - 0x0
      12'h8CB: dout <= 8'b00000000; // 2251 :   0 - 0x0
      12'h8CC: dout <= 8'b00000000; // 2252 :   0 - 0x0
      12'h8CD: dout <= 8'b00000000; // 2253 :   0 - 0x0
      12'h8CE: dout <= 8'b00000000; // 2254 :   0 - 0x0
      12'h8CF: dout <= 8'b00000000; // 2255 :   0 - 0x0
      12'h8D0: dout <= 8'b00000000; // 2256 :   0 - 0x0 -- Background 0x8d
      12'h8D1: dout <= 8'b00000000; // 2257 :   0 - 0x0
      12'h8D2: dout <= 8'b00000000; // 2258 :   0 - 0x0
      12'h8D3: dout <= 8'b00000000; // 2259 :   0 - 0x0
      12'h8D4: dout <= 8'b00000000; // 2260 :   0 - 0x0
      12'h8D5: dout <= 8'b00000000; // 2261 :   0 - 0x0
      12'h8D6: dout <= 8'b00000000; // 2262 :   0 - 0x0
      12'h8D7: dout <= 8'b00000000; // 2263 :   0 - 0x0
      12'h8D8: dout <= 8'b00000000; // 2264 :   0 - 0x0 -- plane 1
      12'h8D9: dout <= 8'b00000000; // 2265 :   0 - 0x0
      12'h8DA: dout <= 8'b00000000; // 2266 :   0 - 0x0
      12'h8DB: dout <= 8'b00000000; // 2267 :   0 - 0x0
      12'h8DC: dout <= 8'b00000000; // 2268 :   0 - 0x0
      12'h8DD: dout <= 8'b00000000; // 2269 :   0 - 0x0
      12'h8DE: dout <= 8'b00000000; // 2270 :   0 - 0x0
      12'h8DF: dout <= 8'b00000000; // 2271 :   0 - 0x0
      12'h8E0: dout <= 8'b00000000; // 2272 :   0 - 0x0 -- Background 0x8e
      12'h8E1: dout <= 8'b00000000; // 2273 :   0 - 0x0
      12'h8E2: dout <= 8'b00000000; // 2274 :   0 - 0x0
      12'h8E3: dout <= 8'b00000000; // 2275 :   0 - 0x0
      12'h8E4: dout <= 8'b00000000; // 2276 :   0 - 0x0
      12'h8E5: dout <= 8'b00000000; // 2277 :   0 - 0x0
      12'h8E6: dout <= 8'b00000000; // 2278 :   0 - 0x0
      12'h8E7: dout <= 8'b00000000; // 2279 :   0 - 0x0
      12'h8E8: dout <= 8'b00000000; // 2280 :   0 - 0x0 -- plane 1
      12'h8E9: dout <= 8'b00000000; // 2281 :   0 - 0x0
      12'h8EA: dout <= 8'b00000000; // 2282 :   0 - 0x0
      12'h8EB: dout <= 8'b00000000; // 2283 :   0 - 0x0
      12'h8EC: dout <= 8'b00000000; // 2284 :   0 - 0x0
      12'h8ED: dout <= 8'b00000000; // 2285 :   0 - 0x0
      12'h8EE: dout <= 8'b00000000; // 2286 :   0 - 0x0
      12'h8EF: dout <= 8'b00000000; // 2287 :   0 - 0x0
      12'h8F0: dout <= 8'b00000000; // 2288 :   0 - 0x0 -- Background 0x8f
      12'h8F1: dout <= 8'b00000000; // 2289 :   0 - 0x0
      12'h8F2: dout <= 8'b00000000; // 2290 :   0 - 0x0
      12'h8F3: dout <= 8'b00000000; // 2291 :   0 - 0x0
      12'h8F4: dout <= 8'b00000000; // 2292 :   0 - 0x0
      12'h8F5: dout <= 8'b00000000; // 2293 :   0 - 0x0
      12'h8F6: dout <= 8'b00000000; // 2294 :   0 - 0x0
      12'h8F7: dout <= 8'b00000000; // 2295 :   0 - 0x0
      12'h8F8: dout <= 8'b00000000; // 2296 :   0 - 0x0 -- plane 1
      12'h8F9: dout <= 8'b00000000; // 2297 :   0 - 0x0
      12'h8FA: dout <= 8'b00000000; // 2298 :   0 - 0x0
      12'h8FB: dout <= 8'b00000000; // 2299 :   0 - 0x0
      12'h8FC: dout <= 8'b00000000; // 2300 :   0 - 0x0
      12'h8FD: dout <= 8'b00000000; // 2301 :   0 - 0x0
      12'h8FE: dout <= 8'b00000000; // 2302 :   0 - 0x0
      12'h8FF: dout <= 8'b00000000; // 2303 :   0 - 0x0
      12'h900: dout <= 8'b00000000; // 2304 :   0 - 0x0 -- Background 0x90
      12'h901: dout <= 8'b00000000; // 2305 :   0 - 0x0
      12'h902: dout <= 8'b00000000; // 2306 :   0 - 0x0
      12'h903: dout <= 8'b00000000; // 2307 :   0 - 0x0
      12'h904: dout <= 8'b00000000; // 2308 :   0 - 0x0
      12'h905: dout <= 8'b00000000; // 2309 :   0 - 0x0
      12'h906: dout <= 8'b00000000; // 2310 :   0 - 0x0
      12'h907: dout <= 8'b00000000; // 2311 :   0 - 0x0
      12'h908: dout <= 8'b00000000; // 2312 :   0 - 0x0 -- plane 1
      12'h909: dout <= 8'b00000000; // 2313 :   0 - 0x0
      12'h90A: dout <= 8'b00000000; // 2314 :   0 - 0x0
      12'h90B: dout <= 8'b00000000; // 2315 :   0 - 0x0
      12'h90C: dout <= 8'b00000000; // 2316 :   0 - 0x0
      12'h90D: dout <= 8'b00000000; // 2317 :   0 - 0x0
      12'h90E: dout <= 8'b00000000; // 2318 :   0 - 0x0
      12'h90F: dout <= 8'b00000000; // 2319 :   0 - 0x0
      12'h910: dout <= 8'b00000000; // 2320 :   0 - 0x0 -- Background 0x91
      12'h911: dout <= 8'b00000000; // 2321 :   0 - 0x0
      12'h912: dout <= 8'b00000000; // 2322 :   0 - 0x0
      12'h913: dout <= 8'b00000000; // 2323 :   0 - 0x0
      12'h914: dout <= 8'b00000000; // 2324 :   0 - 0x0
      12'h915: dout <= 8'b00000000; // 2325 :   0 - 0x0
      12'h916: dout <= 8'b00000000; // 2326 :   0 - 0x0
      12'h917: dout <= 8'b00000000; // 2327 :   0 - 0x0
      12'h918: dout <= 8'b00000000; // 2328 :   0 - 0x0 -- plane 1
      12'h919: dout <= 8'b00000000; // 2329 :   0 - 0x0
      12'h91A: dout <= 8'b00000000; // 2330 :   0 - 0x0
      12'h91B: dout <= 8'b00000000; // 2331 :   0 - 0x0
      12'h91C: dout <= 8'b00000000; // 2332 :   0 - 0x0
      12'h91D: dout <= 8'b00000000; // 2333 :   0 - 0x0
      12'h91E: dout <= 8'b00000000; // 2334 :   0 - 0x0
      12'h91F: dout <= 8'b00000000; // 2335 :   0 - 0x0
      12'h920: dout <= 8'b00000000; // 2336 :   0 - 0x0 -- Background 0x92
      12'h921: dout <= 8'b00000000; // 2337 :   0 - 0x0
      12'h922: dout <= 8'b00000000; // 2338 :   0 - 0x0
      12'h923: dout <= 8'b00000000; // 2339 :   0 - 0x0
      12'h924: dout <= 8'b00000000; // 2340 :   0 - 0x0
      12'h925: dout <= 8'b00000000; // 2341 :   0 - 0x0
      12'h926: dout <= 8'b00000000; // 2342 :   0 - 0x0
      12'h927: dout <= 8'b00000000; // 2343 :   0 - 0x0
      12'h928: dout <= 8'b00000000; // 2344 :   0 - 0x0 -- plane 1
      12'h929: dout <= 8'b00000000; // 2345 :   0 - 0x0
      12'h92A: dout <= 8'b00000000; // 2346 :   0 - 0x0
      12'h92B: dout <= 8'b00000000; // 2347 :   0 - 0x0
      12'h92C: dout <= 8'b00000000; // 2348 :   0 - 0x0
      12'h92D: dout <= 8'b00000000; // 2349 :   0 - 0x0
      12'h92E: dout <= 8'b00000000; // 2350 :   0 - 0x0
      12'h92F: dout <= 8'b00000000; // 2351 :   0 - 0x0
      12'h930: dout <= 8'b00000000; // 2352 :   0 - 0x0 -- Background 0x93
      12'h931: dout <= 8'b00000000; // 2353 :   0 - 0x0
      12'h932: dout <= 8'b00000000; // 2354 :   0 - 0x0
      12'h933: dout <= 8'b00000000; // 2355 :   0 - 0x0
      12'h934: dout <= 8'b00000000; // 2356 :   0 - 0x0
      12'h935: dout <= 8'b00000000; // 2357 :   0 - 0x0
      12'h936: dout <= 8'b00000000; // 2358 :   0 - 0x0
      12'h937: dout <= 8'b00000000; // 2359 :   0 - 0x0
      12'h938: dout <= 8'b00000000; // 2360 :   0 - 0x0 -- plane 1
      12'h939: dout <= 8'b00000000; // 2361 :   0 - 0x0
      12'h93A: dout <= 8'b00000000; // 2362 :   0 - 0x0
      12'h93B: dout <= 8'b00000000; // 2363 :   0 - 0x0
      12'h93C: dout <= 8'b00000000; // 2364 :   0 - 0x0
      12'h93D: dout <= 8'b00000000; // 2365 :   0 - 0x0
      12'h93E: dout <= 8'b00000000; // 2366 :   0 - 0x0
      12'h93F: dout <= 8'b00000000; // 2367 :   0 - 0x0
      12'h940: dout <= 8'b00000000; // 2368 :   0 - 0x0 -- Background 0x94
      12'h941: dout <= 8'b00000000; // 2369 :   0 - 0x0
      12'h942: dout <= 8'b00000000; // 2370 :   0 - 0x0
      12'h943: dout <= 8'b00000000; // 2371 :   0 - 0x0
      12'h944: dout <= 8'b00000000; // 2372 :   0 - 0x0
      12'h945: dout <= 8'b00000000; // 2373 :   0 - 0x0
      12'h946: dout <= 8'b00000000; // 2374 :   0 - 0x0
      12'h947: dout <= 8'b00000000; // 2375 :   0 - 0x0
      12'h948: dout <= 8'b00000000; // 2376 :   0 - 0x0 -- plane 1
      12'h949: dout <= 8'b00000000; // 2377 :   0 - 0x0
      12'h94A: dout <= 8'b00000000; // 2378 :   0 - 0x0
      12'h94B: dout <= 8'b00000000; // 2379 :   0 - 0x0
      12'h94C: dout <= 8'b00000000; // 2380 :   0 - 0x0
      12'h94D: dout <= 8'b00000000; // 2381 :   0 - 0x0
      12'h94E: dout <= 8'b00000000; // 2382 :   0 - 0x0
      12'h94F: dout <= 8'b00000000; // 2383 :   0 - 0x0
      12'h950: dout <= 8'b00000000; // 2384 :   0 - 0x0 -- Background 0x95
      12'h951: dout <= 8'b00000000; // 2385 :   0 - 0x0
      12'h952: dout <= 8'b00000000; // 2386 :   0 - 0x0
      12'h953: dout <= 8'b00000000; // 2387 :   0 - 0x0
      12'h954: dout <= 8'b00000000; // 2388 :   0 - 0x0
      12'h955: dout <= 8'b00000000; // 2389 :   0 - 0x0
      12'h956: dout <= 8'b00000000; // 2390 :   0 - 0x0
      12'h957: dout <= 8'b00000000; // 2391 :   0 - 0x0
      12'h958: dout <= 8'b00000000; // 2392 :   0 - 0x0 -- plane 1
      12'h959: dout <= 8'b00000000; // 2393 :   0 - 0x0
      12'h95A: dout <= 8'b00000000; // 2394 :   0 - 0x0
      12'h95B: dout <= 8'b00000000; // 2395 :   0 - 0x0
      12'h95C: dout <= 8'b00000000; // 2396 :   0 - 0x0
      12'h95D: dout <= 8'b00000000; // 2397 :   0 - 0x0
      12'h95E: dout <= 8'b00000000; // 2398 :   0 - 0x0
      12'h95F: dout <= 8'b00000000; // 2399 :   0 - 0x0
      12'h960: dout <= 8'b00000000; // 2400 :   0 - 0x0 -- Background 0x96
      12'h961: dout <= 8'b00000000; // 2401 :   0 - 0x0
      12'h962: dout <= 8'b00000000; // 2402 :   0 - 0x0
      12'h963: dout <= 8'b00000000; // 2403 :   0 - 0x0
      12'h964: dout <= 8'b00000000; // 2404 :   0 - 0x0
      12'h965: dout <= 8'b00000000; // 2405 :   0 - 0x0
      12'h966: dout <= 8'b00000000; // 2406 :   0 - 0x0
      12'h967: dout <= 8'b00000000; // 2407 :   0 - 0x0
      12'h968: dout <= 8'b00000000; // 2408 :   0 - 0x0 -- plane 1
      12'h969: dout <= 8'b00000000; // 2409 :   0 - 0x0
      12'h96A: dout <= 8'b00000000; // 2410 :   0 - 0x0
      12'h96B: dout <= 8'b00000000; // 2411 :   0 - 0x0
      12'h96C: dout <= 8'b00000000; // 2412 :   0 - 0x0
      12'h96D: dout <= 8'b00000000; // 2413 :   0 - 0x0
      12'h96E: dout <= 8'b00000000; // 2414 :   0 - 0x0
      12'h96F: dout <= 8'b00000000; // 2415 :   0 - 0x0
      12'h970: dout <= 8'b00000000; // 2416 :   0 - 0x0 -- Background 0x97
      12'h971: dout <= 8'b00000000; // 2417 :   0 - 0x0
      12'h972: dout <= 8'b00000000; // 2418 :   0 - 0x0
      12'h973: dout <= 8'b00000000; // 2419 :   0 - 0x0
      12'h974: dout <= 8'b00000000; // 2420 :   0 - 0x0
      12'h975: dout <= 8'b00000000; // 2421 :   0 - 0x0
      12'h976: dout <= 8'b00000000; // 2422 :   0 - 0x0
      12'h977: dout <= 8'b00000000; // 2423 :   0 - 0x0
      12'h978: dout <= 8'b00000000; // 2424 :   0 - 0x0 -- plane 1
      12'h979: dout <= 8'b00000000; // 2425 :   0 - 0x0
      12'h97A: dout <= 8'b00000000; // 2426 :   0 - 0x0
      12'h97B: dout <= 8'b00000000; // 2427 :   0 - 0x0
      12'h97C: dout <= 8'b00000000; // 2428 :   0 - 0x0
      12'h97D: dout <= 8'b00000000; // 2429 :   0 - 0x0
      12'h97E: dout <= 8'b00000000; // 2430 :   0 - 0x0
      12'h97F: dout <= 8'b00000000; // 2431 :   0 - 0x0
      12'h980: dout <= 8'b00000000; // 2432 :   0 - 0x0 -- Background 0x98
      12'h981: dout <= 8'b00000000; // 2433 :   0 - 0x0
      12'h982: dout <= 8'b00000000; // 2434 :   0 - 0x0
      12'h983: dout <= 8'b00000000; // 2435 :   0 - 0x0
      12'h984: dout <= 8'b00000000; // 2436 :   0 - 0x0
      12'h985: dout <= 8'b00000000; // 2437 :   0 - 0x0
      12'h986: dout <= 8'b00000000; // 2438 :   0 - 0x0
      12'h987: dout <= 8'b00000000; // 2439 :   0 - 0x0
      12'h988: dout <= 8'b00000000; // 2440 :   0 - 0x0 -- plane 1
      12'h989: dout <= 8'b00000000; // 2441 :   0 - 0x0
      12'h98A: dout <= 8'b00000000; // 2442 :   0 - 0x0
      12'h98B: dout <= 8'b00000000; // 2443 :   0 - 0x0
      12'h98C: dout <= 8'b00000000; // 2444 :   0 - 0x0
      12'h98D: dout <= 8'b00000000; // 2445 :   0 - 0x0
      12'h98E: dout <= 8'b00000000; // 2446 :   0 - 0x0
      12'h98F: dout <= 8'b00000000; // 2447 :   0 - 0x0
      12'h990: dout <= 8'b00000000; // 2448 :   0 - 0x0 -- Background 0x99
      12'h991: dout <= 8'b00000000; // 2449 :   0 - 0x0
      12'h992: dout <= 8'b00000000; // 2450 :   0 - 0x0
      12'h993: dout <= 8'b00000000; // 2451 :   0 - 0x0
      12'h994: dout <= 8'b00000000; // 2452 :   0 - 0x0
      12'h995: dout <= 8'b00000000; // 2453 :   0 - 0x0
      12'h996: dout <= 8'b00000000; // 2454 :   0 - 0x0
      12'h997: dout <= 8'b00000000; // 2455 :   0 - 0x0
      12'h998: dout <= 8'b00000000; // 2456 :   0 - 0x0 -- plane 1
      12'h999: dout <= 8'b00000000; // 2457 :   0 - 0x0
      12'h99A: dout <= 8'b00000000; // 2458 :   0 - 0x0
      12'h99B: dout <= 8'b00000000; // 2459 :   0 - 0x0
      12'h99C: dout <= 8'b00000000; // 2460 :   0 - 0x0
      12'h99D: dout <= 8'b00000000; // 2461 :   0 - 0x0
      12'h99E: dout <= 8'b00000000; // 2462 :   0 - 0x0
      12'h99F: dout <= 8'b00000000; // 2463 :   0 - 0x0
      12'h9A0: dout <= 8'b00000000; // 2464 :   0 - 0x0 -- Background 0x9a
      12'h9A1: dout <= 8'b00000000; // 2465 :   0 - 0x0
      12'h9A2: dout <= 8'b00000000; // 2466 :   0 - 0x0
      12'h9A3: dout <= 8'b00000000; // 2467 :   0 - 0x0
      12'h9A4: dout <= 8'b00000000; // 2468 :   0 - 0x0
      12'h9A5: dout <= 8'b00000000; // 2469 :   0 - 0x0
      12'h9A6: dout <= 8'b00000000; // 2470 :   0 - 0x0
      12'h9A7: dout <= 8'b00000000; // 2471 :   0 - 0x0
      12'h9A8: dout <= 8'b00000000; // 2472 :   0 - 0x0 -- plane 1
      12'h9A9: dout <= 8'b00000000; // 2473 :   0 - 0x0
      12'h9AA: dout <= 8'b00000000; // 2474 :   0 - 0x0
      12'h9AB: dout <= 8'b00000000; // 2475 :   0 - 0x0
      12'h9AC: dout <= 8'b00000000; // 2476 :   0 - 0x0
      12'h9AD: dout <= 8'b00000000; // 2477 :   0 - 0x0
      12'h9AE: dout <= 8'b00000000; // 2478 :   0 - 0x0
      12'h9AF: dout <= 8'b00000000; // 2479 :   0 - 0x0
      12'h9B0: dout <= 8'b00000000; // 2480 :   0 - 0x0 -- Background 0x9b
      12'h9B1: dout <= 8'b00000000; // 2481 :   0 - 0x0
      12'h9B2: dout <= 8'b00000000; // 2482 :   0 - 0x0
      12'h9B3: dout <= 8'b00000000; // 2483 :   0 - 0x0
      12'h9B4: dout <= 8'b00000000; // 2484 :   0 - 0x0
      12'h9B5: dout <= 8'b00000000; // 2485 :   0 - 0x0
      12'h9B6: dout <= 8'b00000000; // 2486 :   0 - 0x0
      12'h9B7: dout <= 8'b00000000; // 2487 :   0 - 0x0
      12'h9B8: dout <= 8'b00000000; // 2488 :   0 - 0x0 -- plane 1
      12'h9B9: dout <= 8'b00000000; // 2489 :   0 - 0x0
      12'h9BA: dout <= 8'b00000000; // 2490 :   0 - 0x0
      12'h9BB: dout <= 8'b00000000; // 2491 :   0 - 0x0
      12'h9BC: dout <= 8'b00000000; // 2492 :   0 - 0x0
      12'h9BD: dout <= 8'b00000000; // 2493 :   0 - 0x0
      12'h9BE: dout <= 8'b00000000; // 2494 :   0 - 0x0
      12'h9BF: dout <= 8'b00000000; // 2495 :   0 - 0x0
      12'h9C0: dout <= 8'b00000000; // 2496 :   0 - 0x0 -- Background 0x9c
      12'h9C1: dout <= 8'b00000000; // 2497 :   0 - 0x0
      12'h9C2: dout <= 8'b00000000; // 2498 :   0 - 0x0
      12'h9C3: dout <= 8'b00000000; // 2499 :   0 - 0x0
      12'h9C4: dout <= 8'b00000000; // 2500 :   0 - 0x0
      12'h9C5: dout <= 8'b00000000; // 2501 :   0 - 0x0
      12'h9C6: dout <= 8'b00000000; // 2502 :   0 - 0x0
      12'h9C7: dout <= 8'b00000000; // 2503 :   0 - 0x0
      12'h9C8: dout <= 8'b00000000; // 2504 :   0 - 0x0 -- plane 1
      12'h9C9: dout <= 8'b00000000; // 2505 :   0 - 0x0
      12'h9CA: dout <= 8'b00000000; // 2506 :   0 - 0x0
      12'h9CB: dout <= 8'b00000000; // 2507 :   0 - 0x0
      12'h9CC: dout <= 8'b00000000; // 2508 :   0 - 0x0
      12'h9CD: dout <= 8'b00000000; // 2509 :   0 - 0x0
      12'h9CE: dout <= 8'b00000000; // 2510 :   0 - 0x0
      12'h9CF: dout <= 8'b00000000; // 2511 :   0 - 0x0
      12'h9D0: dout <= 8'b00000000; // 2512 :   0 - 0x0 -- Background 0x9d
      12'h9D1: dout <= 8'b00000000; // 2513 :   0 - 0x0
      12'h9D2: dout <= 8'b00000000; // 2514 :   0 - 0x0
      12'h9D3: dout <= 8'b00000000; // 2515 :   0 - 0x0
      12'h9D4: dout <= 8'b00000000; // 2516 :   0 - 0x0
      12'h9D5: dout <= 8'b00000000; // 2517 :   0 - 0x0
      12'h9D6: dout <= 8'b00000000; // 2518 :   0 - 0x0
      12'h9D7: dout <= 8'b00000000; // 2519 :   0 - 0x0
      12'h9D8: dout <= 8'b00000000; // 2520 :   0 - 0x0 -- plane 1
      12'h9D9: dout <= 8'b00000000; // 2521 :   0 - 0x0
      12'h9DA: dout <= 8'b00000000; // 2522 :   0 - 0x0
      12'h9DB: dout <= 8'b00000000; // 2523 :   0 - 0x0
      12'h9DC: dout <= 8'b00000000; // 2524 :   0 - 0x0
      12'h9DD: dout <= 8'b00000000; // 2525 :   0 - 0x0
      12'h9DE: dout <= 8'b00000000; // 2526 :   0 - 0x0
      12'h9DF: dout <= 8'b00000000; // 2527 :   0 - 0x0
      12'h9E0: dout <= 8'b00000000; // 2528 :   0 - 0x0 -- Background 0x9e
      12'h9E1: dout <= 8'b00000000; // 2529 :   0 - 0x0
      12'h9E2: dout <= 8'b00000000; // 2530 :   0 - 0x0
      12'h9E3: dout <= 8'b00000000; // 2531 :   0 - 0x0
      12'h9E4: dout <= 8'b00000000; // 2532 :   0 - 0x0
      12'h9E5: dout <= 8'b00000000; // 2533 :   0 - 0x0
      12'h9E6: dout <= 8'b00000000; // 2534 :   0 - 0x0
      12'h9E7: dout <= 8'b00000000; // 2535 :   0 - 0x0
      12'h9E8: dout <= 8'b00000000; // 2536 :   0 - 0x0 -- plane 1
      12'h9E9: dout <= 8'b00000000; // 2537 :   0 - 0x0
      12'h9EA: dout <= 8'b00000000; // 2538 :   0 - 0x0
      12'h9EB: dout <= 8'b00000000; // 2539 :   0 - 0x0
      12'h9EC: dout <= 8'b00000000; // 2540 :   0 - 0x0
      12'h9ED: dout <= 8'b00000000; // 2541 :   0 - 0x0
      12'h9EE: dout <= 8'b00000000; // 2542 :   0 - 0x0
      12'h9EF: dout <= 8'b00000000; // 2543 :   0 - 0x0
      12'h9F0: dout <= 8'b00000000; // 2544 :   0 - 0x0 -- Background 0x9f
      12'h9F1: dout <= 8'b00000000; // 2545 :   0 - 0x0
      12'h9F2: dout <= 8'b00000000; // 2546 :   0 - 0x0
      12'h9F3: dout <= 8'b00000000; // 2547 :   0 - 0x0
      12'h9F4: dout <= 8'b00000000; // 2548 :   0 - 0x0
      12'h9F5: dout <= 8'b00000000; // 2549 :   0 - 0x0
      12'h9F6: dout <= 8'b00000000; // 2550 :   0 - 0x0
      12'h9F7: dout <= 8'b00000000; // 2551 :   0 - 0x0
      12'h9F8: dout <= 8'b00000000; // 2552 :   0 - 0x0 -- plane 1
      12'h9F9: dout <= 8'b00000000; // 2553 :   0 - 0x0
      12'h9FA: dout <= 8'b00000000; // 2554 :   0 - 0x0
      12'h9FB: dout <= 8'b00000000; // 2555 :   0 - 0x0
      12'h9FC: dout <= 8'b00000000; // 2556 :   0 - 0x0
      12'h9FD: dout <= 8'b00000000; // 2557 :   0 - 0x0
      12'h9FE: dout <= 8'b00000000; // 2558 :   0 - 0x0
      12'h9FF: dout <= 8'b00000000; // 2559 :   0 - 0x0
      12'hA00: dout <= 8'b00000000; // 2560 :   0 - 0x0 -- Background 0xa0
      12'hA01: dout <= 8'b00000000; // 2561 :   0 - 0x0
      12'hA02: dout <= 8'b00000000; // 2562 :   0 - 0x0
      12'hA03: dout <= 8'b00000000; // 2563 :   0 - 0x0
      12'hA04: dout <= 8'b00000000; // 2564 :   0 - 0x0
      12'hA05: dout <= 8'b00000000; // 2565 :   0 - 0x0
      12'hA06: dout <= 8'b00000000; // 2566 :   0 - 0x0
      12'hA07: dout <= 8'b00000000; // 2567 :   0 - 0x0
      12'hA08: dout <= 8'b00000000; // 2568 :   0 - 0x0 -- plane 1
      12'hA09: dout <= 8'b00000000; // 2569 :   0 - 0x0
      12'hA0A: dout <= 8'b00000000; // 2570 :   0 - 0x0
      12'hA0B: dout <= 8'b00000000; // 2571 :   0 - 0x0
      12'hA0C: dout <= 8'b00000000; // 2572 :   0 - 0x0
      12'hA0D: dout <= 8'b00000000; // 2573 :   0 - 0x0
      12'hA0E: dout <= 8'b00000000; // 2574 :   0 - 0x0
      12'hA0F: dout <= 8'b00000000; // 2575 :   0 - 0x0
      12'hA10: dout <= 8'b00000000; // 2576 :   0 - 0x0 -- Background 0xa1
      12'hA11: dout <= 8'b00000000; // 2577 :   0 - 0x0
      12'hA12: dout <= 8'b00000000; // 2578 :   0 - 0x0
      12'hA13: dout <= 8'b00000000; // 2579 :   0 - 0x0
      12'hA14: dout <= 8'b00000000; // 2580 :   0 - 0x0
      12'hA15: dout <= 8'b00000000; // 2581 :   0 - 0x0
      12'hA16: dout <= 8'b00000000; // 2582 :   0 - 0x0
      12'hA17: dout <= 8'b00000000; // 2583 :   0 - 0x0
      12'hA18: dout <= 8'b00000000; // 2584 :   0 - 0x0 -- plane 1
      12'hA19: dout <= 8'b00000000; // 2585 :   0 - 0x0
      12'hA1A: dout <= 8'b00000000; // 2586 :   0 - 0x0
      12'hA1B: dout <= 8'b00000000; // 2587 :   0 - 0x0
      12'hA1C: dout <= 8'b00000000; // 2588 :   0 - 0x0
      12'hA1D: dout <= 8'b00000000; // 2589 :   0 - 0x0
      12'hA1E: dout <= 8'b00000000; // 2590 :   0 - 0x0
      12'hA1F: dout <= 8'b00000000; // 2591 :   0 - 0x0
      12'hA20: dout <= 8'b00000000; // 2592 :   0 - 0x0 -- Background 0xa2
      12'hA21: dout <= 8'b00000000; // 2593 :   0 - 0x0
      12'hA22: dout <= 8'b00000000; // 2594 :   0 - 0x0
      12'hA23: dout <= 8'b00000000; // 2595 :   0 - 0x0
      12'hA24: dout <= 8'b00000000; // 2596 :   0 - 0x0
      12'hA25: dout <= 8'b00000000; // 2597 :   0 - 0x0
      12'hA26: dout <= 8'b00000000; // 2598 :   0 - 0x0
      12'hA27: dout <= 8'b00000000; // 2599 :   0 - 0x0
      12'hA28: dout <= 8'b00000000; // 2600 :   0 - 0x0 -- plane 1
      12'hA29: dout <= 8'b00000000; // 2601 :   0 - 0x0
      12'hA2A: dout <= 8'b00000000; // 2602 :   0 - 0x0
      12'hA2B: dout <= 8'b00000000; // 2603 :   0 - 0x0
      12'hA2C: dout <= 8'b00000000; // 2604 :   0 - 0x0
      12'hA2D: dout <= 8'b00000000; // 2605 :   0 - 0x0
      12'hA2E: dout <= 8'b00000000; // 2606 :   0 - 0x0
      12'hA2F: dout <= 8'b00000000; // 2607 :   0 - 0x0
      12'hA30: dout <= 8'b00000000; // 2608 :   0 - 0x0 -- Background 0xa3
      12'hA31: dout <= 8'b00000000; // 2609 :   0 - 0x0
      12'hA32: dout <= 8'b00000000; // 2610 :   0 - 0x0
      12'hA33: dout <= 8'b00000000; // 2611 :   0 - 0x0
      12'hA34: dout <= 8'b00000000; // 2612 :   0 - 0x0
      12'hA35: dout <= 8'b00000000; // 2613 :   0 - 0x0
      12'hA36: dout <= 8'b00000000; // 2614 :   0 - 0x0
      12'hA37: dout <= 8'b00000000; // 2615 :   0 - 0x0
      12'hA38: dout <= 8'b00000000; // 2616 :   0 - 0x0 -- plane 1
      12'hA39: dout <= 8'b00000000; // 2617 :   0 - 0x0
      12'hA3A: dout <= 8'b00000000; // 2618 :   0 - 0x0
      12'hA3B: dout <= 8'b00000000; // 2619 :   0 - 0x0
      12'hA3C: dout <= 8'b00000000; // 2620 :   0 - 0x0
      12'hA3D: dout <= 8'b00000000; // 2621 :   0 - 0x0
      12'hA3E: dout <= 8'b00000000; // 2622 :   0 - 0x0
      12'hA3F: dout <= 8'b00000000; // 2623 :   0 - 0x0
      12'hA40: dout <= 8'b00000000; // 2624 :   0 - 0x0 -- Background 0xa4
      12'hA41: dout <= 8'b00000000; // 2625 :   0 - 0x0
      12'hA42: dout <= 8'b00000000; // 2626 :   0 - 0x0
      12'hA43: dout <= 8'b00000000; // 2627 :   0 - 0x0
      12'hA44: dout <= 8'b00000000; // 2628 :   0 - 0x0
      12'hA45: dout <= 8'b00000000; // 2629 :   0 - 0x0
      12'hA46: dout <= 8'b00000000; // 2630 :   0 - 0x0
      12'hA47: dout <= 8'b00000000; // 2631 :   0 - 0x0
      12'hA48: dout <= 8'b00000000; // 2632 :   0 - 0x0 -- plane 1
      12'hA49: dout <= 8'b00000000; // 2633 :   0 - 0x0
      12'hA4A: dout <= 8'b00000000; // 2634 :   0 - 0x0
      12'hA4B: dout <= 8'b00000000; // 2635 :   0 - 0x0
      12'hA4C: dout <= 8'b00000000; // 2636 :   0 - 0x0
      12'hA4D: dout <= 8'b00000000; // 2637 :   0 - 0x0
      12'hA4E: dout <= 8'b00000000; // 2638 :   0 - 0x0
      12'hA4F: dout <= 8'b00000000; // 2639 :   0 - 0x0
      12'hA50: dout <= 8'b00000000; // 2640 :   0 - 0x0 -- Background 0xa5
      12'hA51: dout <= 8'b00000000; // 2641 :   0 - 0x0
      12'hA52: dout <= 8'b00000000; // 2642 :   0 - 0x0
      12'hA53: dout <= 8'b00000000; // 2643 :   0 - 0x0
      12'hA54: dout <= 8'b00000000; // 2644 :   0 - 0x0
      12'hA55: dout <= 8'b00000000; // 2645 :   0 - 0x0
      12'hA56: dout <= 8'b00000000; // 2646 :   0 - 0x0
      12'hA57: dout <= 8'b00000000; // 2647 :   0 - 0x0
      12'hA58: dout <= 8'b00000000; // 2648 :   0 - 0x0 -- plane 1
      12'hA59: dout <= 8'b00000000; // 2649 :   0 - 0x0
      12'hA5A: dout <= 8'b00000000; // 2650 :   0 - 0x0
      12'hA5B: dout <= 8'b00000000; // 2651 :   0 - 0x0
      12'hA5C: dout <= 8'b00000000; // 2652 :   0 - 0x0
      12'hA5D: dout <= 8'b00000000; // 2653 :   0 - 0x0
      12'hA5E: dout <= 8'b00000000; // 2654 :   0 - 0x0
      12'hA5F: dout <= 8'b00000000; // 2655 :   0 - 0x0
      12'hA60: dout <= 8'b00000000; // 2656 :   0 - 0x0 -- Background 0xa6
      12'hA61: dout <= 8'b00000000; // 2657 :   0 - 0x0
      12'hA62: dout <= 8'b00000000; // 2658 :   0 - 0x0
      12'hA63: dout <= 8'b00000000; // 2659 :   0 - 0x0
      12'hA64: dout <= 8'b00000000; // 2660 :   0 - 0x0
      12'hA65: dout <= 8'b00000000; // 2661 :   0 - 0x0
      12'hA66: dout <= 8'b00000000; // 2662 :   0 - 0x0
      12'hA67: dout <= 8'b00000000; // 2663 :   0 - 0x0
      12'hA68: dout <= 8'b00000000; // 2664 :   0 - 0x0 -- plane 1
      12'hA69: dout <= 8'b00000000; // 2665 :   0 - 0x0
      12'hA6A: dout <= 8'b00000000; // 2666 :   0 - 0x0
      12'hA6B: dout <= 8'b00000000; // 2667 :   0 - 0x0
      12'hA6C: dout <= 8'b00000000; // 2668 :   0 - 0x0
      12'hA6D: dout <= 8'b00000000; // 2669 :   0 - 0x0
      12'hA6E: dout <= 8'b00000000; // 2670 :   0 - 0x0
      12'hA6F: dout <= 8'b00000000; // 2671 :   0 - 0x0
      12'hA70: dout <= 8'b00000000; // 2672 :   0 - 0x0 -- Background 0xa7
      12'hA71: dout <= 8'b00000000; // 2673 :   0 - 0x0
      12'hA72: dout <= 8'b00000000; // 2674 :   0 - 0x0
      12'hA73: dout <= 8'b00000000; // 2675 :   0 - 0x0
      12'hA74: dout <= 8'b00000000; // 2676 :   0 - 0x0
      12'hA75: dout <= 8'b00000000; // 2677 :   0 - 0x0
      12'hA76: dout <= 8'b00000000; // 2678 :   0 - 0x0
      12'hA77: dout <= 8'b00000000; // 2679 :   0 - 0x0
      12'hA78: dout <= 8'b00000000; // 2680 :   0 - 0x0 -- plane 1
      12'hA79: dout <= 8'b00000000; // 2681 :   0 - 0x0
      12'hA7A: dout <= 8'b00000000; // 2682 :   0 - 0x0
      12'hA7B: dout <= 8'b00000000; // 2683 :   0 - 0x0
      12'hA7C: dout <= 8'b00000000; // 2684 :   0 - 0x0
      12'hA7D: dout <= 8'b00000000; // 2685 :   0 - 0x0
      12'hA7E: dout <= 8'b00000000; // 2686 :   0 - 0x0
      12'hA7F: dout <= 8'b00000000; // 2687 :   0 - 0x0
      12'hA80: dout <= 8'b00000000; // 2688 :   0 - 0x0 -- Background 0xa8
      12'hA81: dout <= 8'b00000000; // 2689 :   0 - 0x0
      12'hA82: dout <= 8'b00000000; // 2690 :   0 - 0x0
      12'hA83: dout <= 8'b00000000; // 2691 :   0 - 0x0
      12'hA84: dout <= 8'b00000000; // 2692 :   0 - 0x0
      12'hA85: dout <= 8'b00000000; // 2693 :   0 - 0x0
      12'hA86: dout <= 8'b00000000; // 2694 :   0 - 0x0
      12'hA87: dout <= 8'b00000000; // 2695 :   0 - 0x0
      12'hA88: dout <= 8'b00000000; // 2696 :   0 - 0x0 -- plane 1
      12'hA89: dout <= 8'b00000000; // 2697 :   0 - 0x0
      12'hA8A: dout <= 8'b00000000; // 2698 :   0 - 0x0
      12'hA8B: dout <= 8'b00000000; // 2699 :   0 - 0x0
      12'hA8C: dout <= 8'b00000000; // 2700 :   0 - 0x0
      12'hA8D: dout <= 8'b00000000; // 2701 :   0 - 0x0
      12'hA8E: dout <= 8'b00000000; // 2702 :   0 - 0x0
      12'hA8F: dout <= 8'b00000000; // 2703 :   0 - 0x0
      12'hA90: dout <= 8'b00000000; // 2704 :   0 - 0x0 -- Background 0xa9
      12'hA91: dout <= 8'b00000000; // 2705 :   0 - 0x0
      12'hA92: dout <= 8'b00000000; // 2706 :   0 - 0x0
      12'hA93: dout <= 8'b00000000; // 2707 :   0 - 0x0
      12'hA94: dout <= 8'b00000000; // 2708 :   0 - 0x0
      12'hA95: dout <= 8'b00000000; // 2709 :   0 - 0x0
      12'hA96: dout <= 8'b00000000; // 2710 :   0 - 0x0
      12'hA97: dout <= 8'b00000000; // 2711 :   0 - 0x0
      12'hA98: dout <= 8'b00000000; // 2712 :   0 - 0x0 -- plane 1
      12'hA99: dout <= 8'b00000000; // 2713 :   0 - 0x0
      12'hA9A: dout <= 8'b00000000; // 2714 :   0 - 0x0
      12'hA9B: dout <= 8'b00000000; // 2715 :   0 - 0x0
      12'hA9C: dout <= 8'b00000000; // 2716 :   0 - 0x0
      12'hA9D: dout <= 8'b00000000; // 2717 :   0 - 0x0
      12'hA9E: dout <= 8'b00000000; // 2718 :   0 - 0x0
      12'hA9F: dout <= 8'b00000000; // 2719 :   0 - 0x0
      12'hAA0: dout <= 8'b00000000; // 2720 :   0 - 0x0 -- Background 0xaa
      12'hAA1: dout <= 8'b00000000; // 2721 :   0 - 0x0
      12'hAA2: dout <= 8'b00000000; // 2722 :   0 - 0x0
      12'hAA3: dout <= 8'b00000000; // 2723 :   0 - 0x0
      12'hAA4: dout <= 8'b00000000; // 2724 :   0 - 0x0
      12'hAA5: dout <= 8'b00000000; // 2725 :   0 - 0x0
      12'hAA6: dout <= 8'b00000000; // 2726 :   0 - 0x0
      12'hAA7: dout <= 8'b00000000; // 2727 :   0 - 0x0
      12'hAA8: dout <= 8'b00000000; // 2728 :   0 - 0x0 -- plane 1
      12'hAA9: dout <= 8'b00000000; // 2729 :   0 - 0x0
      12'hAAA: dout <= 8'b00000000; // 2730 :   0 - 0x0
      12'hAAB: dout <= 8'b00000000; // 2731 :   0 - 0x0
      12'hAAC: dout <= 8'b00000000; // 2732 :   0 - 0x0
      12'hAAD: dout <= 8'b00000000; // 2733 :   0 - 0x0
      12'hAAE: dout <= 8'b00000000; // 2734 :   0 - 0x0
      12'hAAF: dout <= 8'b00000000; // 2735 :   0 - 0x0
      12'hAB0: dout <= 8'b00000000; // 2736 :   0 - 0x0 -- Background 0xab
      12'hAB1: dout <= 8'b00000000; // 2737 :   0 - 0x0
      12'hAB2: dout <= 8'b00000000; // 2738 :   0 - 0x0
      12'hAB3: dout <= 8'b00000000; // 2739 :   0 - 0x0
      12'hAB4: dout <= 8'b00000000; // 2740 :   0 - 0x0
      12'hAB5: dout <= 8'b00000000; // 2741 :   0 - 0x0
      12'hAB6: dout <= 8'b00000000; // 2742 :   0 - 0x0
      12'hAB7: dout <= 8'b00000000; // 2743 :   0 - 0x0
      12'hAB8: dout <= 8'b00000000; // 2744 :   0 - 0x0 -- plane 1
      12'hAB9: dout <= 8'b00000000; // 2745 :   0 - 0x0
      12'hABA: dout <= 8'b00000000; // 2746 :   0 - 0x0
      12'hABB: dout <= 8'b00000000; // 2747 :   0 - 0x0
      12'hABC: dout <= 8'b00000000; // 2748 :   0 - 0x0
      12'hABD: dout <= 8'b00000000; // 2749 :   0 - 0x0
      12'hABE: dout <= 8'b00000000; // 2750 :   0 - 0x0
      12'hABF: dout <= 8'b00000000; // 2751 :   0 - 0x0
      12'hAC0: dout <= 8'b00000000; // 2752 :   0 - 0x0 -- Background 0xac
      12'hAC1: dout <= 8'b00000000; // 2753 :   0 - 0x0
      12'hAC2: dout <= 8'b00000000; // 2754 :   0 - 0x0
      12'hAC3: dout <= 8'b00000000; // 2755 :   0 - 0x0
      12'hAC4: dout <= 8'b00000000; // 2756 :   0 - 0x0
      12'hAC5: dout <= 8'b00000000; // 2757 :   0 - 0x0
      12'hAC6: dout <= 8'b00000000; // 2758 :   0 - 0x0
      12'hAC7: dout <= 8'b00000000; // 2759 :   0 - 0x0
      12'hAC8: dout <= 8'b00000000; // 2760 :   0 - 0x0 -- plane 1
      12'hAC9: dout <= 8'b00000000; // 2761 :   0 - 0x0
      12'hACA: dout <= 8'b00000000; // 2762 :   0 - 0x0
      12'hACB: dout <= 8'b00000000; // 2763 :   0 - 0x0
      12'hACC: dout <= 8'b00000000; // 2764 :   0 - 0x0
      12'hACD: dout <= 8'b00000000; // 2765 :   0 - 0x0
      12'hACE: dout <= 8'b00000000; // 2766 :   0 - 0x0
      12'hACF: dout <= 8'b00000000; // 2767 :   0 - 0x0
      12'hAD0: dout <= 8'b00000000; // 2768 :   0 - 0x0 -- Background 0xad
      12'hAD1: dout <= 8'b00000000; // 2769 :   0 - 0x0
      12'hAD2: dout <= 8'b00000000; // 2770 :   0 - 0x0
      12'hAD3: dout <= 8'b00000000; // 2771 :   0 - 0x0
      12'hAD4: dout <= 8'b00000000; // 2772 :   0 - 0x0
      12'hAD5: dout <= 8'b00000000; // 2773 :   0 - 0x0
      12'hAD6: dout <= 8'b00000000; // 2774 :   0 - 0x0
      12'hAD7: dout <= 8'b00000000; // 2775 :   0 - 0x0
      12'hAD8: dout <= 8'b00000000; // 2776 :   0 - 0x0 -- plane 1
      12'hAD9: dout <= 8'b00000000; // 2777 :   0 - 0x0
      12'hADA: dout <= 8'b00000000; // 2778 :   0 - 0x0
      12'hADB: dout <= 8'b00000000; // 2779 :   0 - 0x0
      12'hADC: dout <= 8'b00000000; // 2780 :   0 - 0x0
      12'hADD: dout <= 8'b00000000; // 2781 :   0 - 0x0
      12'hADE: dout <= 8'b00000000; // 2782 :   0 - 0x0
      12'hADF: dout <= 8'b00000000; // 2783 :   0 - 0x0
      12'hAE0: dout <= 8'b00000000; // 2784 :   0 - 0x0 -- Background 0xae
      12'hAE1: dout <= 8'b00000000; // 2785 :   0 - 0x0
      12'hAE2: dout <= 8'b00000000; // 2786 :   0 - 0x0
      12'hAE3: dout <= 8'b00000000; // 2787 :   0 - 0x0
      12'hAE4: dout <= 8'b00000000; // 2788 :   0 - 0x0
      12'hAE5: dout <= 8'b00000000; // 2789 :   0 - 0x0
      12'hAE6: dout <= 8'b00000000; // 2790 :   0 - 0x0
      12'hAE7: dout <= 8'b00000000; // 2791 :   0 - 0x0
      12'hAE8: dout <= 8'b00000000; // 2792 :   0 - 0x0 -- plane 1
      12'hAE9: dout <= 8'b00000000; // 2793 :   0 - 0x0
      12'hAEA: dout <= 8'b00000000; // 2794 :   0 - 0x0
      12'hAEB: dout <= 8'b00000000; // 2795 :   0 - 0x0
      12'hAEC: dout <= 8'b00000000; // 2796 :   0 - 0x0
      12'hAED: dout <= 8'b00000000; // 2797 :   0 - 0x0
      12'hAEE: dout <= 8'b00000000; // 2798 :   0 - 0x0
      12'hAEF: dout <= 8'b00000000; // 2799 :   0 - 0x0
      12'hAF0: dout <= 8'b00000000; // 2800 :   0 - 0x0 -- Background 0xaf
      12'hAF1: dout <= 8'b00000000; // 2801 :   0 - 0x0
      12'hAF2: dout <= 8'b00000000; // 2802 :   0 - 0x0
      12'hAF3: dout <= 8'b00000000; // 2803 :   0 - 0x0
      12'hAF4: dout <= 8'b00000000; // 2804 :   0 - 0x0
      12'hAF5: dout <= 8'b00000000; // 2805 :   0 - 0x0
      12'hAF6: dout <= 8'b00000000; // 2806 :   0 - 0x0
      12'hAF7: dout <= 8'b00000000; // 2807 :   0 - 0x0
      12'hAF8: dout <= 8'b00000000; // 2808 :   0 - 0x0 -- plane 1
      12'hAF9: dout <= 8'b00000000; // 2809 :   0 - 0x0
      12'hAFA: dout <= 8'b00000000; // 2810 :   0 - 0x0
      12'hAFB: dout <= 8'b00000000; // 2811 :   0 - 0x0
      12'hAFC: dout <= 8'b00000000; // 2812 :   0 - 0x0
      12'hAFD: dout <= 8'b00000000; // 2813 :   0 - 0x0
      12'hAFE: dout <= 8'b00000000; // 2814 :   0 - 0x0
      12'hAFF: dout <= 8'b00000000; // 2815 :   0 - 0x0
      12'hB00: dout <= 8'b00000000; // 2816 :   0 - 0x0 -- Background 0xb0
      12'hB01: dout <= 8'b00000000; // 2817 :   0 - 0x0
      12'hB02: dout <= 8'b00000000; // 2818 :   0 - 0x0
      12'hB03: dout <= 8'b00000000; // 2819 :   0 - 0x0
      12'hB04: dout <= 8'b00000000; // 2820 :   0 - 0x0
      12'hB05: dout <= 8'b00000000; // 2821 :   0 - 0x0
      12'hB06: dout <= 8'b00000000; // 2822 :   0 - 0x0
      12'hB07: dout <= 8'b00000000; // 2823 :   0 - 0x0
      12'hB08: dout <= 8'b00000000; // 2824 :   0 - 0x0 -- plane 1
      12'hB09: dout <= 8'b00000000; // 2825 :   0 - 0x0
      12'hB0A: dout <= 8'b00000000; // 2826 :   0 - 0x0
      12'hB0B: dout <= 8'b00000000; // 2827 :   0 - 0x0
      12'hB0C: dout <= 8'b00000000; // 2828 :   0 - 0x0
      12'hB0D: dout <= 8'b00000000; // 2829 :   0 - 0x0
      12'hB0E: dout <= 8'b00000000; // 2830 :   0 - 0x0
      12'hB0F: dout <= 8'b00000000; // 2831 :   0 - 0x0
      12'hB10: dout <= 8'b00000000; // 2832 :   0 - 0x0 -- Background 0xb1
      12'hB11: dout <= 8'b00000000; // 2833 :   0 - 0x0
      12'hB12: dout <= 8'b00000000; // 2834 :   0 - 0x0
      12'hB13: dout <= 8'b00000000; // 2835 :   0 - 0x0
      12'hB14: dout <= 8'b00000000; // 2836 :   0 - 0x0
      12'hB15: dout <= 8'b00000000; // 2837 :   0 - 0x0
      12'hB16: dout <= 8'b00000000; // 2838 :   0 - 0x0
      12'hB17: dout <= 8'b00000000; // 2839 :   0 - 0x0
      12'hB18: dout <= 8'b00000000; // 2840 :   0 - 0x0 -- plane 1
      12'hB19: dout <= 8'b00000000; // 2841 :   0 - 0x0
      12'hB1A: dout <= 8'b00000000; // 2842 :   0 - 0x0
      12'hB1B: dout <= 8'b00000000; // 2843 :   0 - 0x0
      12'hB1C: dout <= 8'b00000000; // 2844 :   0 - 0x0
      12'hB1D: dout <= 8'b00000000; // 2845 :   0 - 0x0
      12'hB1E: dout <= 8'b00000000; // 2846 :   0 - 0x0
      12'hB1F: dout <= 8'b00000000; // 2847 :   0 - 0x0
      12'hB20: dout <= 8'b00000000; // 2848 :   0 - 0x0 -- Background 0xb2
      12'hB21: dout <= 8'b00000000; // 2849 :   0 - 0x0
      12'hB22: dout <= 8'b00000000; // 2850 :   0 - 0x0
      12'hB23: dout <= 8'b00000000; // 2851 :   0 - 0x0
      12'hB24: dout <= 8'b00000000; // 2852 :   0 - 0x0
      12'hB25: dout <= 8'b00000000; // 2853 :   0 - 0x0
      12'hB26: dout <= 8'b00000000; // 2854 :   0 - 0x0
      12'hB27: dout <= 8'b00000000; // 2855 :   0 - 0x0
      12'hB28: dout <= 8'b00000000; // 2856 :   0 - 0x0 -- plane 1
      12'hB29: dout <= 8'b00000000; // 2857 :   0 - 0x0
      12'hB2A: dout <= 8'b00000000; // 2858 :   0 - 0x0
      12'hB2B: dout <= 8'b00000000; // 2859 :   0 - 0x0
      12'hB2C: dout <= 8'b00000000; // 2860 :   0 - 0x0
      12'hB2D: dout <= 8'b00000000; // 2861 :   0 - 0x0
      12'hB2E: dout <= 8'b00000000; // 2862 :   0 - 0x0
      12'hB2F: dout <= 8'b00000000; // 2863 :   0 - 0x0
      12'hB30: dout <= 8'b00000000; // 2864 :   0 - 0x0 -- Background 0xb3
      12'hB31: dout <= 8'b00000000; // 2865 :   0 - 0x0
      12'hB32: dout <= 8'b00000000; // 2866 :   0 - 0x0
      12'hB33: dout <= 8'b00000000; // 2867 :   0 - 0x0
      12'hB34: dout <= 8'b00000000; // 2868 :   0 - 0x0
      12'hB35: dout <= 8'b00000000; // 2869 :   0 - 0x0
      12'hB36: dout <= 8'b00000000; // 2870 :   0 - 0x0
      12'hB37: dout <= 8'b00000000; // 2871 :   0 - 0x0
      12'hB38: dout <= 8'b00000000; // 2872 :   0 - 0x0 -- plane 1
      12'hB39: dout <= 8'b00000000; // 2873 :   0 - 0x0
      12'hB3A: dout <= 8'b00000000; // 2874 :   0 - 0x0
      12'hB3B: dout <= 8'b00000000; // 2875 :   0 - 0x0
      12'hB3C: dout <= 8'b00000000; // 2876 :   0 - 0x0
      12'hB3D: dout <= 8'b00000000; // 2877 :   0 - 0x0
      12'hB3E: dout <= 8'b00000000; // 2878 :   0 - 0x0
      12'hB3F: dout <= 8'b00000000; // 2879 :   0 - 0x0
      12'hB40: dout <= 8'b00000000; // 2880 :   0 - 0x0 -- Background 0xb4
      12'hB41: dout <= 8'b00000000; // 2881 :   0 - 0x0
      12'hB42: dout <= 8'b00000000; // 2882 :   0 - 0x0
      12'hB43: dout <= 8'b00000000; // 2883 :   0 - 0x0
      12'hB44: dout <= 8'b00000000; // 2884 :   0 - 0x0
      12'hB45: dout <= 8'b00000000; // 2885 :   0 - 0x0
      12'hB46: dout <= 8'b00000000; // 2886 :   0 - 0x0
      12'hB47: dout <= 8'b00000000; // 2887 :   0 - 0x0
      12'hB48: dout <= 8'b00000000; // 2888 :   0 - 0x0 -- plane 1
      12'hB49: dout <= 8'b00000000; // 2889 :   0 - 0x0
      12'hB4A: dout <= 8'b00000000; // 2890 :   0 - 0x0
      12'hB4B: dout <= 8'b00000000; // 2891 :   0 - 0x0
      12'hB4C: dout <= 8'b00000000; // 2892 :   0 - 0x0
      12'hB4D: dout <= 8'b00000000; // 2893 :   0 - 0x0
      12'hB4E: dout <= 8'b00000000; // 2894 :   0 - 0x0
      12'hB4F: dout <= 8'b00000000; // 2895 :   0 - 0x0
      12'hB50: dout <= 8'b00000000; // 2896 :   0 - 0x0 -- Background 0xb5
      12'hB51: dout <= 8'b00000000; // 2897 :   0 - 0x0
      12'hB52: dout <= 8'b00000000; // 2898 :   0 - 0x0
      12'hB53: dout <= 8'b00000000; // 2899 :   0 - 0x0
      12'hB54: dout <= 8'b00000000; // 2900 :   0 - 0x0
      12'hB55: dout <= 8'b00000000; // 2901 :   0 - 0x0
      12'hB56: dout <= 8'b00000000; // 2902 :   0 - 0x0
      12'hB57: dout <= 8'b00000000; // 2903 :   0 - 0x0
      12'hB58: dout <= 8'b00000000; // 2904 :   0 - 0x0 -- plane 1
      12'hB59: dout <= 8'b00000000; // 2905 :   0 - 0x0
      12'hB5A: dout <= 8'b00000000; // 2906 :   0 - 0x0
      12'hB5B: dout <= 8'b00000000; // 2907 :   0 - 0x0
      12'hB5C: dout <= 8'b00000000; // 2908 :   0 - 0x0
      12'hB5D: dout <= 8'b00000000; // 2909 :   0 - 0x0
      12'hB5E: dout <= 8'b00000000; // 2910 :   0 - 0x0
      12'hB5F: dout <= 8'b00000000; // 2911 :   0 - 0x0
      12'hB60: dout <= 8'b00000000; // 2912 :   0 - 0x0 -- Background 0xb6
      12'hB61: dout <= 8'b00000000; // 2913 :   0 - 0x0
      12'hB62: dout <= 8'b00000000; // 2914 :   0 - 0x0
      12'hB63: dout <= 8'b00000000; // 2915 :   0 - 0x0
      12'hB64: dout <= 8'b00000000; // 2916 :   0 - 0x0
      12'hB65: dout <= 8'b00000000; // 2917 :   0 - 0x0
      12'hB66: dout <= 8'b00000000; // 2918 :   0 - 0x0
      12'hB67: dout <= 8'b00000000; // 2919 :   0 - 0x0
      12'hB68: dout <= 8'b00000000; // 2920 :   0 - 0x0 -- plane 1
      12'hB69: dout <= 8'b00000000; // 2921 :   0 - 0x0
      12'hB6A: dout <= 8'b00000000; // 2922 :   0 - 0x0
      12'hB6B: dout <= 8'b00000000; // 2923 :   0 - 0x0
      12'hB6C: dout <= 8'b00000000; // 2924 :   0 - 0x0
      12'hB6D: dout <= 8'b00000000; // 2925 :   0 - 0x0
      12'hB6E: dout <= 8'b00000000; // 2926 :   0 - 0x0
      12'hB6F: dout <= 8'b00000000; // 2927 :   0 - 0x0
      12'hB70: dout <= 8'b00000000; // 2928 :   0 - 0x0 -- Background 0xb7
      12'hB71: dout <= 8'b00000000; // 2929 :   0 - 0x0
      12'hB72: dout <= 8'b00000000; // 2930 :   0 - 0x0
      12'hB73: dout <= 8'b00000000; // 2931 :   0 - 0x0
      12'hB74: dout <= 8'b00000000; // 2932 :   0 - 0x0
      12'hB75: dout <= 8'b00000000; // 2933 :   0 - 0x0
      12'hB76: dout <= 8'b00000000; // 2934 :   0 - 0x0
      12'hB77: dout <= 8'b00000000; // 2935 :   0 - 0x0
      12'hB78: dout <= 8'b00000000; // 2936 :   0 - 0x0 -- plane 1
      12'hB79: dout <= 8'b00000000; // 2937 :   0 - 0x0
      12'hB7A: dout <= 8'b00000000; // 2938 :   0 - 0x0
      12'hB7B: dout <= 8'b00000000; // 2939 :   0 - 0x0
      12'hB7C: dout <= 8'b00000000; // 2940 :   0 - 0x0
      12'hB7D: dout <= 8'b00000000; // 2941 :   0 - 0x0
      12'hB7E: dout <= 8'b00000000; // 2942 :   0 - 0x0
      12'hB7F: dout <= 8'b00000000; // 2943 :   0 - 0x0
      12'hB80: dout <= 8'b00000000; // 2944 :   0 - 0x0 -- Background 0xb8
      12'hB81: dout <= 8'b00000000; // 2945 :   0 - 0x0
      12'hB82: dout <= 8'b00000000; // 2946 :   0 - 0x0
      12'hB83: dout <= 8'b00000000; // 2947 :   0 - 0x0
      12'hB84: dout <= 8'b00000000; // 2948 :   0 - 0x0
      12'hB85: dout <= 8'b00000000; // 2949 :   0 - 0x0
      12'hB86: dout <= 8'b00000000; // 2950 :   0 - 0x0
      12'hB87: dout <= 8'b00000000; // 2951 :   0 - 0x0
      12'hB88: dout <= 8'b00000000; // 2952 :   0 - 0x0 -- plane 1
      12'hB89: dout <= 8'b00000000; // 2953 :   0 - 0x0
      12'hB8A: dout <= 8'b00000000; // 2954 :   0 - 0x0
      12'hB8B: dout <= 8'b00000000; // 2955 :   0 - 0x0
      12'hB8C: dout <= 8'b00000000; // 2956 :   0 - 0x0
      12'hB8D: dout <= 8'b00000000; // 2957 :   0 - 0x0
      12'hB8E: dout <= 8'b00000000; // 2958 :   0 - 0x0
      12'hB8F: dout <= 8'b00000000; // 2959 :   0 - 0x0
      12'hB90: dout <= 8'b00000000; // 2960 :   0 - 0x0 -- Background 0xb9
      12'hB91: dout <= 8'b00000000; // 2961 :   0 - 0x0
      12'hB92: dout <= 8'b00000000; // 2962 :   0 - 0x0
      12'hB93: dout <= 8'b00000000; // 2963 :   0 - 0x0
      12'hB94: dout <= 8'b00000000; // 2964 :   0 - 0x0
      12'hB95: dout <= 8'b00000000; // 2965 :   0 - 0x0
      12'hB96: dout <= 8'b00000000; // 2966 :   0 - 0x0
      12'hB97: dout <= 8'b00000000; // 2967 :   0 - 0x0
      12'hB98: dout <= 8'b00000000; // 2968 :   0 - 0x0 -- plane 1
      12'hB99: dout <= 8'b00000000; // 2969 :   0 - 0x0
      12'hB9A: dout <= 8'b00000000; // 2970 :   0 - 0x0
      12'hB9B: dout <= 8'b00000000; // 2971 :   0 - 0x0
      12'hB9C: dout <= 8'b00000000; // 2972 :   0 - 0x0
      12'hB9D: dout <= 8'b00000000; // 2973 :   0 - 0x0
      12'hB9E: dout <= 8'b00000000; // 2974 :   0 - 0x0
      12'hB9F: dout <= 8'b00000000; // 2975 :   0 - 0x0
      12'hBA0: dout <= 8'b00000000; // 2976 :   0 - 0x0 -- Background 0xba
      12'hBA1: dout <= 8'b00000000; // 2977 :   0 - 0x0
      12'hBA2: dout <= 8'b00000000; // 2978 :   0 - 0x0
      12'hBA3: dout <= 8'b00000000; // 2979 :   0 - 0x0
      12'hBA4: dout <= 8'b00000000; // 2980 :   0 - 0x0
      12'hBA5: dout <= 8'b00000000; // 2981 :   0 - 0x0
      12'hBA6: dout <= 8'b00000000; // 2982 :   0 - 0x0
      12'hBA7: dout <= 8'b00000000; // 2983 :   0 - 0x0
      12'hBA8: dout <= 8'b00000000; // 2984 :   0 - 0x0 -- plane 1
      12'hBA9: dout <= 8'b00000000; // 2985 :   0 - 0x0
      12'hBAA: dout <= 8'b00000000; // 2986 :   0 - 0x0
      12'hBAB: dout <= 8'b00000000; // 2987 :   0 - 0x0
      12'hBAC: dout <= 8'b00000000; // 2988 :   0 - 0x0
      12'hBAD: dout <= 8'b00000000; // 2989 :   0 - 0x0
      12'hBAE: dout <= 8'b00000000; // 2990 :   0 - 0x0
      12'hBAF: dout <= 8'b00000000; // 2991 :   0 - 0x0
      12'hBB0: dout <= 8'b00000000; // 2992 :   0 - 0x0 -- Background 0xbb
      12'hBB1: dout <= 8'b00000000; // 2993 :   0 - 0x0
      12'hBB2: dout <= 8'b00000000; // 2994 :   0 - 0x0
      12'hBB3: dout <= 8'b00000000; // 2995 :   0 - 0x0
      12'hBB4: dout <= 8'b00000000; // 2996 :   0 - 0x0
      12'hBB5: dout <= 8'b00000000; // 2997 :   0 - 0x0
      12'hBB6: dout <= 8'b00000000; // 2998 :   0 - 0x0
      12'hBB7: dout <= 8'b00000000; // 2999 :   0 - 0x0
      12'hBB8: dout <= 8'b00000000; // 3000 :   0 - 0x0 -- plane 1
      12'hBB9: dout <= 8'b00000000; // 3001 :   0 - 0x0
      12'hBBA: dout <= 8'b00000000; // 3002 :   0 - 0x0
      12'hBBB: dout <= 8'b00000000; // 3003 :   0 - 0x0
      12'hBBC: dout <= 8'b00000000; // 3004 :   0 - 0x0
      12'hBBD: dout <= 8'b00000000; // 3005 :   0 - 0x0
      12'hBBE: dout <= 8'b00000000; // 3006 :   0 - 0x0
      12'hBBF: dout <= 8'b00000000; // 3007 :   0 - 0x0
      12'hBC0: dout <= 8'b00000000; // 3008 :   0 - 0x0 -- Background 0xbc
      12'hBC1: dout <= 8'b00000000; // 3009 :   0 - 0x0
      12'hBC2: dout <= 8'b00000000; // 3010 :   0 - 0x0
      12'hBC3: dout <= 8'b00000000; // 3011 :   0 - 0x0
      12'hBC4: dout <= 8'b00000000; // 3012 :   0 - 0x0
      12'hBC5: dout <= 8'b00000000; // 3013 :   0 - 0x0
      12'hBC6: dout <= 8'b00000000; // 3014 :   0 - 0x0
      12'hBC7: dout <= 8'b00000000; // 3015 :   0 - 0x0
      12'hBC8: dout <= 8'b00000000; // 3016 :   0 - 0x0 -- plane 1
      12'hBC9: dout <= 8'b00000000; // 3017 :   0 - 0x0
      12'hBCA: dout <= 8'b00000000; // 3018 :   0 - 0x0
      12'hBCB: dout <= 8'b00000000; // 3019 :   0 - 0x0
      12'hBCC: dout <= 8'b00000000; // 3020 :   0 - 0x0
      12'hBCD: dout <= 8'b00000000; // 3021 :   0 - 0x0
      12'hBCE: dout <= 8'b00000000; // 3022 :   0 - 0x0
      12'hBCF: dout <= 8'b00000000; // 3023 :   0 - 0x0
      12'hBD0: dout <= 8'b00000000; // 3024 :   0 - 0x0 -- Background 0xbd
      12'hBD1: dout <= 8'b00000000; // 3025 :   0 - 0x0
      12'hBD2: dout <= 8'b00000000; // 3026 :   0 - 0x0
      12'hBD3: dout <= 8'b00000000; // 3027 :   0 - 0x0
      12'hBD4: dout <= 8'b00000000; // 3028 :   0 - 0x0
      12'hBD5: dout <= 8'b00000000; // 3029 :   0 - 0x0
      12'hBD6: dout <= 8'b00000000; // 3030 :   0 - 0x0
      12'hBD7: dout <= 8'b00000000; // 3031 :   0 - 0x0
      12'hBD8: dout <= 8'b00000000; // 3032 :   0 - 0x0 -- plane 1
      12'hBD9: dout <= 8'b00000000; // 3033 :   0 - 0x0
      12'hBDA: dout <= 8'b00000000; // 3034 :   0 - 0x0
      12'hBDB: dout <= 8'b00000000; // 3035 :   0 - 0x0
      12'hBDC: dout <= 8'b00000000; // 3036 :   0 - 0x0
      12'hBDD: dout <= 8'b00000000; // 3037 :   0 - 0x0
      12'hBDE: dout <= 8'b00000000; // 3038 :   0 - 0x0
      12'hBDF: dout <= 8'b00000000; // 3039 :   0 - 0x0
      12'hBE0: dout <= 8'b00000000; // 3040 :   0 - 0x0 -- Background 0xbe
      12'hBE1: dout <= 8'b00000000; // 3041 :   0 - 0x0
      12'hBE2: dout <= 8'b00000000; // 3042 :   0 - 0x0
      12'hBE3: dout <= 8'b00000000; // 3043 :   0 - 0x0
      12'hBE4: dout <= 8'b00000000; // 3044 :   0 - 0x0
      12'hBE5: dout <= 8'b00000000; // 3045 :   0 - 0x0
      12'hBE6: dout <= 8'b00000000; // 3046 :   0 - 0x0
      12'hBE7: dout <= 8'b00000000; // 3047 :   0 - 0x0
      12'hBE8: dout <= 8'b00000000; // 3048 :   0 - 0x0 -- plane 1
      12'hBE9: dout <= 8'b00000000; // 3049 :   0 - 0x0
      12'hBEA: dout <= 8'b00000000; // 3050 :   0 - 0x0
      12'hBEB: dout <= 8'b00000000; // 3051 :   0 - 0x0
      12'hBEC: dout <= 8'b00000000; // 3052 :   0 - 0x0
      12'hBED: dout <= 8'b00000000; // 3053 :   0 - 0x0
      12'hBEE: dout <= 8'b00000000; // 3054 :   0 - 0x0
      12'hBEF: dout <= 8'b00000000; // 3055 :   0 - 0x0
      12'hBF0: dout <= 8'b00000000; // 3056 :   0 - 0x0 -- Background 0xbf
      12'hBF1: dout <= 8'b00000000; // 3057 :   0 - 0x0
      12'hBF2: dout <= 8'b00000000; // 3058 :   0 - 0x0
      12'hBF3: dout <= 8'b00000000; // 3059 :   0 - 0x0
      12'hBF4: dout <= 8'b00000000; // 3060 :   0 - 0x0
      12'hBF5: dout <= 8'b00000000; // 3061 :   0 - 0x0
      12'hBF6: dout <= 8'b00000000; // 3062 :   0 - 0x0
      12'hBF7: dout <= 8'b00000000; // 3063 :   0 - 0x0
      12'hBF8: dout <= 8'b00000000; // 3064 :   0 - 0x0 -- plane 1
      12'hBF9: dout <= 8'b00000000; // 3065 :   0 - 0x0
      12'hBFA: dout <= 8'b00000000; // 3066 :   0 - 0x0
      12'hBFB: dout <= 8'b00000000; // 3067 :   0 - 0x0
      12'hBFC: dout <= 8'b00000000; // 3068 :   0 - 0x0
      12'hBFD: dout <= 8'b00000000; // 3069 :   0 - 0x0
      12'hBFE: dout <= 8'b00000000; // 3070 :   0 - 0x0
      12'hBFF: dout <= 8'b00000000; // 3071 :   0 - 0x0
      12'hC00: dout <= 8'b00000000; // 3072 :   0 - 0x0 -- Background 0xc0
      12'hC01: dout <= 8'b00000000; // 3073 :   0 - 0x0
      12'hC02: dout <= 8'b00000000; // 3074 :   0 - 0x0
      12'hC03: dout <= 8'b00000000; // 3075 :   0 - 0x0
      12'hC04: dout <= 8'b00000000; // 3076 :   0 - 0x0
      12'hC05: dout <= 8'b00000000; // 3077 :   0 - 0x0
      12'hC06: dout <= 8'b00000000; // 3078 :   0 - 0x0
      12'hC07: dout <= 8'b00000000; // 3079 :   0 - 0x0
      12'hC08: dout <= 8'b00000000; // 3080 :   0 - 0x0 -- plane 1
      12'hC09: dout <= 8'b00000000; // 3081 :   0 - 0x0
      12'hC0A: dout <= 8'b00000000; // 3082 :   0 - 0x0
      12'hC0B: dout <= 8'b00000000; // 3083 :   0 - 0x0
      12'hC0C: dout <= 8'b00000000; // 3084 :   0 - 0x0
      12'hC0D: dout <= 8'b00000000; // 3085 :   0 - 0x0
      12'hC0E: dout <= 8'b00000000; // 3086 :   0 - 0x0
      12'hC0F: dout <= 8'b00000000; // 3087 :   0 - 0x0
      12'hC10: dout <= 8'b00000000; // 3088 :   0 - 0x0 -- Background 0xc1
      12'hC11: dout <= 8'b00000000; // 3089 :   0 - 0x0
      12'hC12: dout <= 8'b00000000; // 3090 :   0 - 0x0
      12'hC13: dout <= 8'b00000000; // 3091 :   0 - 0x0
      12'hC14: dout <= 8'b00000000; // 3092 :   0 - 0x0
      12'hC15: dout <= 8'b00000000; // 3093 :   0 - 0x0
      12'hC16: dout <= 8'b00000000; // 3094 :   0 - 0x0
      12'hC17: dout <= 8'b00000000; // 3095 :   0 - 0x0
      12'hC18: dout <= 8'b00000000; // 3096 :   0 - 0x0 -- plane 1
      12'hC19: dout <= 8'b00000000; // 3097 :   0 - 0x0
      12'hC1A: dout <= 8'b00000000; // 3098 :   0 - 0x0
      12'hC1B: dout <= 8'b00000000; // 3099 :   0 - 0x0
      12'hC1C: dout <= 8'b00000000; // 3100 :   0 - 0x0
      12'hC1D: dout <= 8'b00000000; // 3101 :   0 - 0x0
      12'hC1E: dout <= 8'b00000000; // 3102 :   0 - 0x0
      12'hC1F: dout <= 8'b00000000; // 3103 :   0 - 0x0
      12'hC20: dout <= 8'b00000000; // 3104 :   0 - 0x0 -- Background 0xc2
      12'hC21: dout <= 8'b00000000; // 3105 :   0 - 0x0
      12'hC22: dout <= 8'b00000000; // 3106 :   0 - 0x0
      12'hC23: dout <= 8'b00000000; // 3107 :   0 - 0x0
      12'hC24: dout <= 8'b00000000; // 3108 :   0 - 0x0
      12'hC25: dout <= 8'b00000000; // 3109 :   0 - 0x0
      12'hC26: dout <= 8'b00000000; // 3110 :   0 - 0x0
      12'hC27: dout <= 8'b00000000; // 3111 :   0 - 0x0
      12'hC28: dout <= 8'b00000000; // 3112 :   0 - 0x0 -- plane 1
      12'hC29: dout <= 8'b00000000; // 3113 :   0 - 0x0
      12'hC2A: dout <= 8'b00000000; // 3114 :   0 - 0x0
      12'hC2B: dout <= 8'b00000000; // 3115 :   0 - 0x0
      12'hC2C: dout <= 8'b00000000; // 3116 :   0 - 0x0
      12'hC2D: dout <= 8'b00000000; // 3117 :   0 - 0x0
      12'hC2E: dout <= 8'b00000000; // 3118 :   0 - 0x0
      12'hC2F: dout <= 8'b00000000; // 3119 :   0 - 0x0
      12'hC30: dout <= 8'b00000000; // 3120 :   0 - 0x0 -- Background 0xc3
      12'hC31: dout <= 8'b00000000; // 3121 :   0 - 0x0
      12'hC32: dout <= 8'b00000000; // 3122 :   0 - 0x0
      12'hC33: dout <= 8'b00000000; // 3123 :   0 - 0x0
      12'hC34: dout <= 8'b00000000; // 3124 :   0 - 0x0
      12'hC35: dout <= 8'b00000000; // 3125 :   0 - 0x0
      12'hC36: dout <= 8'b00000000; // 3126 :   0 - 0x0
      12'hC37: dout <= 8'b00000000; // 3127 :   0 - 0x0
      12'hC38: dout <= 8'b00000000; // 3128 :   0 - 0x0 -- plane 1
      12'hC39: dout <= 8'b00000000; // 3129 :   0 - 0x0
      12'hC3A: dout <= 8'b00000000; // 3130 :   0 - 0x0
      12'hC3B: dout <= 8'b00000000; // 3131 :   0 - 0x0
      12'hC3C: dout <= 8'b00000000; // 3132 :   0 - 0x0
      12'hC3D: dout <= 8'b00000000; // 3133 :   0 - 0x0
      12'hC3E: dout <= 8'b00000000; // 3134 :   0 - 0x0
      12'hC3F: dout <= 8'b00000000; // 3135 :   0 - 0x0
      12'hC40: dout <= 8'b00000000; // 3136 :   0 - 0x0 -- Background 0xc4
      12'hC41: dout <= 8'b00000000; // 3137 :   0 - 0x0
      12'hC42: dout <= 8'b00000000; // 3138 :   0 - 0x0
      12'hC43: dout <= 8'b00000000; // 3139 :   0 - 0x0
      12'hC44: dout <= 8'b00000000; // 3140 :   0 - 0x0
      12'hC45: dout <= 8'b00000000; // 3141 :   0 - 0x0
      12'hC46: dout <= 8'b00000000; // 3142 :   0 - 0x0
      12'hC47: dout <= 8'b00000000; // 3143 :   0 - 0x0
      12'hC48: dout <= 8'b00000000; // 3144 :   0 - 0x0 -- plane 1
      12'hC49: dout <= 8'b00000000; // 3145 :   0 - 0x0
      12'hC4A: dout <= 8'b00000000; // 3146 :   0 - 0x0
      12'hC4B: dout <= 8'b00000000; // 3147 :   0 - 0x0
      12'hC4C: dout <= 8'b00000000; // 3148 :   0 - 0x0
      12'hC4D: dout <= 8'b00000000; // 3149 :   0 - 0x0
      12'hC4E: dout <= 8'b00000000; // 3150 :   0 - 0x0
      12'hC4F: dout <= 8'b00000000; // 3151 :   0 - 0x0
      12'hC50: dout <= 8'b00000000; // 3152 :   0 - 0x0 -- Background 0xc5
      12'hC51: dout <= 8'b00000000; // 3153 :   0 - 0x0
      12'hC52: dout <= 8'b00000000; // 3154 :   0 - 0x0
      12'hC53: dout <= 8'b00000000; // 3155 :   0 - 0x0
      12'hC54: dout <= 8'b00000000; // 3156 :   0 - 0x0
      12'hC55: dout <= 8'b00000000; // 3157 :   0 - 0x0
      12'hC56: dout <= 8'b00000000; // 3158 :   0 - 0x0
      12'hC57: dout <= 8'b00000000; // 3159 :   0 - 0x0
      12'hC58: dout <= 8'b00000000; // 3160 :   0 - 0x0 -- plane 1
      12'hC59: dout <= 8'b00000000; // 3161 :   0 - 0x0
      12'hC5A: dout <= 8'b00000000; // 3162 :   0 - 0x0
      12'hC5B: dout <= 8'b00000000; // 3163 :   0 - 0x0
      12'hC5C: dout <= 8'b00000000; // 3164 :   0 - 0x0
      12'hC5D: dout <= 8'b00000000; // 3165 :   0 - 0x0
      12'hC5E: dout <= 8'b00000000; // 3166 :   0 - 0x0
      12'hC5F: dout <= 8'b00000000; // 3167 :   0 - 0x0
      12'hC60: dout <= 8'b00000000; // 3168 :   0 - 0x0 -- Background 0xc6
      12'hC61: dout <= 8'b00000000; // 3169 :   0 - 0x0
      12'hC62: dout <= 8'b00000000; // 3170 :   0 - 0x0
      12'hC63: dout <= 8'b00000000; // 3171 :   0 - 0x0
      12'hC64: dout <= 8'b00000000; // 3172 :   0 - 0x0
      12'hC65: dout <= 8'b00000000; // 3173 :   0 - 0x0
      12'hC66: dout <= 8'b00000000; // 3174 :   0 - 0x0
      12'hC67: dout <= 8'b00000000; // 3175 :   0 - 0x0
      12'hC68: dout <= 8'b00000000; // 3176 :   0 - 0x0 -- plane 1
      12'hC69: dout <= 8'b00000000; // 3177 :   0 - 0x0
      12'hC6A: dout <= 8'b00000000; // 3178 :   0 - 0x0
      12'hC6B: dout <= 8'b00000000; // 3179 :   0 - 0x0
      12'hC6C: dout <= 8'b00000000; // 3180 :   0 - 0x0
      12'hC6D: dout <= 8'b00000000; // 3181 :   0 - 0x0
      12'hC6E: dout <= 8'b00000000; // 3182 :   0 - 0x0
      12'hC6F: dout <= 8'b00000000; // 3183 :   0 - 0x0
      12'hC70: dout <= 8'b00000000; // 3184 :   0 - 0x0 -- Background 0xc7
      12'hC71: dout <= 8'b00000000; // 3185 :   0 - 0x0
      12'hC72: dout <= 8'b00000000; // 3186 :   0 - 0x0
      12'hC73: dout <= 8'b00000000; // 3187 :   0 - 0x0
      12'hC74: dout <= 8'b00000000; // 3188 :   0 - 0x0
      12'hC75: dout <= 8'b00000000; // 3189 :   0 - 0x0
      12'hC76: dout <= 8'b00000000; // 3190 :   0 - 0x0
      12'hC77: dout <= 8'b00000000; // 3191 :   0 - 0x0
      12'hC78: dout <= 8'b00000000; // 3192 :   0 - 0x0 -- plane 1
      12'hC79: dout <= 8'b00000000; // 3193 :   0 - 0x0
      12'hC7A: dout <= 8'b00000000; // 3194 :   0 - 0x0
      12'hC7B: dout <= 8'b00000000; // 3195 :   0 - 0x0
      12'hC7C: dout <= 8'b00000000; // 3196 :   0 - 0x0
      12'hC7D: dout <= 8'b00000000; // 3197 :   0 - 0x0
      12'hC7E: dout <= 8'b00000000; // 3198 :   0 - 0x0
      12'hC7F: dout <= 8'b00000000; // 3199 :   0 - 0x0
      12'hC80: dout <= 8'b00000000; // 3200 :   0 - 0x0 -- Background 0xc8
      12'hC81: dout <= 8'b00000000; // 3201 :   0 - 0x0
      12'hC82: dout <= 8'b00000000; // 3202 :   0 - 0x0
      12'hC83: dout <= 8'b00000000; // 3203 :   0 - 0x0
      12'hC84: dout <= 8'b00000000; // 3204 :   0 - 0x0
      12'hC85: dout <= 8'b00000000; // 3205 :   0 - 0x0
      12'hC86: dout <= 8'b00000000; // 3206 :   0 - 0x0
      12'hC87: dout <= 8'b00000000; // 3207 :   0 - 0x0
      12'hC88: dout <= 8'b00000000; // 3208 :   0 - 0x0 -- plane 1
      12'hC89: dout <= 8'b00000000; // 3209 :   0 - 0x0
      12'hC8A: dout <= 8'b00000000; // 3210 :   0 - 0x0
      12'hC8B: dout <= 8'b00000000; // 3211 :   0 - 0x0
      12'hC8C: dout <= 8'b00000000; // 3212 :   0 - 0x0
      12'hC8D: dout <= 8'b00000000; // 3213 :   0 - 0x0
      12'hC8E: dout <= 8'b00000000; // 3214 :   0 - 0x0
      12'hC8F: dout <= 8'b00000000; // 3215 :   0 - 0x0
      12'hC90: dout <= 8'b00000000; // 3216 :   0 - 0x0 -- Background 0xc9
      12'hC91: dout <= 8'b00000000; // 3217 :   0 - 0x0
      12'hC92: dout <= 8'b00000000; // 3218 :   0 - 0x0
      12'hC93: dout <= 8'b00000000; // 3219 :   0 - 0x0
      12'hC94: dout <= 8'b00000000; // 3220 :   0 - 0x0
      12'hC95: dout <= 8'b00000000; // 3221 :   0 - 0x0
      12'hC96: dout <= 8'b00000000; // 3222 :   0 - 0x0
      12'hC97: dout <= 8'b00000000; // 3223 :   0 - 0x0
      12'hC98: dout <= 8'b00000000; // 3224 :   0 - 0x0 -- plane 1
      12'hC99: dout <= 8'b00000000; // 3225 :   0 - 0x0
      12'hC9A: dout <= 8'b00000000; // 3226 :   0 - 0x0
      12'hC9B: dout <= 8'b00000000; // 3227 :   0 - 0x0
      12'hC9C: dout <= 8'b00000000; // 3228 :   0 - 0x0
      12'hC9D: dout <= 8'b00000000; // 3229 :   0 - 0x0
      12'hC9E: dout <= 8'b00000000; // 3230 :   0 - 0x0
      12'hC9F: dout <= 8'b00000000; // 3231 :   0 - 0x0
      12'hCA0: dout <= 8'b00000000; // 3232 :   0 - 0x0 -- Background 0xca
      12'hCA1: dout <= 8'b00000000; // 3233 :   0 - 0x0
      12'hCA2: dout <= 8'b00000000; // 3234 :   0 - 0x0
      12'hCA3: dout <= 8'b00000000; // 3235 :   0 - 0x0
      12'hCA4: dout <= 8'b00000000; // 3236 :   0 - 0x0
      12'hCA5: dout <= 8'b00000000; // 3237 :   0 - 0x0
      12'hCA6: dout <= 8'b00000000; // 3238 :   0 - 0x0
      12'hCA7: dout <= 8'b00000000; // 3239 :   0 - 0x0
      12'hCA8: dout <= 8'b00000000; // 3240 :   0 - 0x0 -- plane 1
      12'hCA9: dout <= 8'b00000000; // 3241 :   0 - 0x0
      12'hCAA: dout <= 8'b00000000; // 3242 :   0 - 0x0
      12'hCAB: dout <= 8'b00000000; // 3243 :   0 - 0x0
      12'hCAC: dout <= 8'b00000000; // 3244 :   0 - 0x0
      12'hCAD: dout <= 8'b00000000; // 3245 :   0 - 0x0
      12'hCAE: dout <= 8'b00000000; // 3246 :   0 - 0x0
      12'hCAF: dout <= 8'b00000000; // 3247 :   0 - 0x0
      12'hCB0: dout <= 8'b00000000; // 3248 :   0 - 0x0 -- Background 0xcb
      12'hCB1: dout <= 8'b00000000; // 3249 :   0 - 0x0
      12'hCB2: dout <= 8'b00000000; // 3250 :   0 - 0x0
      12'hCB3: dout <= 8'b00000000; // 3251 :   0 - 0x0
      12'hCB4: dout <= 8'b00000000; // 3252 :   0 - 0x0
      12'hCB5: dout <= 8'b00000000; // 3253 :   0 - 0x0
      12'hCB6: dout <= 8'b00000000; // 3254 :   0 - 0x0
      12'hCB7: dout <= 8'b00000000; // 3255 :   0 - 0x0
      12'hCB8: dout <= 8'b00000000; // 3256 :   0 - 0x0 -- plane 1
      12'hCB9: dout <= 8'b00000000; // 3257 :   0 - 0x0
      12'hCBA: dout <= 8'b00000000; // 3258 :   0 - 0x0
      12'hCBB: dout <= 8'b00000000; // 3259 :   0 - 0x0
      12'hCBC: dout <= 8'b00000000; // 3260 :   0 - 0x0
      12'hCBD: dout <= 8'b00000000; // 3261 :   0 - 0x0
      12'hCBE: dout <= 8'b00000000; // 3262 :   0 - 0x0
      12'hCBF: dout <= 8'b00000000; // 3263 :   0 - 0x0
      12'hCC0: dout <= 8'b00000000; // 3264 :   0 - 0x0 -- Background 0xcc
      12'hCC1: dout <= 8'b00000000; // 3265 :   0 - 0x0
      12'hCC2: dout <= 8'b00000000; // 3266 :   0 - 0x0
      12'hCC3: dout <= 8'b00000000; // 3267 :   0 - 0x0
      12'hCC4: dout <= 8'b00000000; // 3268 :   0 - 0x0
      12'hCC5: dout <= 8'b00000000; // 3269 :   0 - 0x0
      12'hCC6: dout <= 8'b00000000; // 3270 :   0 - 0x0
      12'hCC7: dout <= 8'b00000000; // 3271 :   0 - 0x0
      12'hCC8: dout <= 8'b00000000; // 3272 :   0 - 0x0 -- plane 1
      12'hCC9: dout <= 8'b00000000; // 3273 :   0 - 0x0
      12'hCCA: dout <= 8'b00000000; // 3274 :   0 - 0x0
      12'hCCB: dout <= 8'b00000000; // 3275 :   0 - 0x0
      12'hCCC: dout <= 8'b00000000; // 3276 :   0 - 0x0
      12'hCCD: dout <= 8'b00000000; // 3277 :   0 - 0x0
      12'hCCE: dout <= 8'b00000000; // 3278 :   0 - 0x0
      12'hCCF: dout <= 8'b00000000; // 3279 :   0 - 0x0
      12'hCD0: dout <= 8'b00111111; // 3280 :  63 - 0x3f -- Background 0xcd
      12'hCD1: dout <= 8'b01111111; // 3281 : 127 - 0x7f
      12'hCD2: dout <= 8'b11111111; // 3282 : 255 - 0xff
      12'hCD3: dout <= 8'b11110000; // 3283 : 240 - 0xf0
      12'hCD4: dout <= 8'b11100000; // 3284 : 224 - 0xe0
      12'hCD5: dout <= 8'b11100011; // 3285 : 227 - 0xe3
      12'hCD6: dout <= 8'b11100111; // 3286 : 231 - 0xe7
      12'hCD7: dout <= 8'b11100111; // 3287 : 231 - 0xe7
      12'hCD8: dout <= 8'b11000000; // 3288 : 192 - 0xc0 -- plane 1
      12'hCD9: dout <= 8'b10000000; // 3289 : 128 - 0x80
      12'hCDA: dout <= 8'b00000000; // 3290 :   0 - 0x0
      12'hCDB: dout <= 8'b00001111; // 3291 :  15 - 0xf
      12'hCDC: dout <= 8'b00011111; // 3292 :  31 - 0x1f
      12'hCDD: dout <= 8'b00011100; // 3293 :  28 - 0x1c
      12'hCDE: dout <= 8'b00011000; // 3294 :  24 - 0x18
      12'hCDF: dout <= 8'b00011000; // 3295 :  24 - 0x18
      12'hCE0: dout <= 8'b11111100; // 3296 : 252 - 0xfc -- Background 0xce
      12'hCE1: dout <= 8'b11111110; // 3297 : 254 - 0xfe
      12'hCE2: dout <= 8'b11111111; // 3298 : 255 - 0xff
      12'hCE3: dout <= 8'b00001111; // 3299 :  15 - 0xf
      12'hCE4: dout <= 8'b00000111; // 3300 :   7 - 0x7
      12'hCE5: dout <= 8'b11000111; // 3301 : 199 - 0xc7
      12'hCE6: dout <= 8'b11100111; // 3302 : 231 - 0xe7
      12'hCE7: dout <= 8'b11100111; // 3303 : 231 - 0xe7
      12'hCE8: dout <= 8'b00000011; // 3304 :   3 - 0x3 -- plane 1
      12'hCE9: dout <= 8'b00000001; // 3305 :   1 - 0x1
      12'hCEA: dout <= 8'b00000000; // 3306 :   0 - 0x0
      12'hCEB: dout <= 8'b11110000; // 3307 : 240 - 0xf0
      12'hCEC: dout <= 8'b11111000; // 3308 : 248 - 0xf8
      12'hCED: dout <= 8'b00111000; // 3309 :  56 - 0x38
      12'hCEE: dout <= 8'b00011000; // 3310 :  24 - 0x18
      12'hCEF: dout <= 8'b00011000; // 3311 :  24 - 0x18
      12'hCF0: dout <= 8'b00000000; // 3312 :   0 - 0x0 -- Background 0xcf
      12'hCF1: dout <= 8'b00000000; // 3313 :   0 - 0x0
      12'hCF2: dout <= 8'b00000000; // 3314 :   0 - 0x0
      12'hCF3: dout <= 8'b00000000; // 3315 :   0 - 0x0
      12'hCF4: dout <= 8'b00000000; // 3316 :   0 - 0x0
      12'hCF5: dout <= 8'b00000000; // 3317 :   0 - 0x0
      12'hCF6: dout <= 8'b00000000; // 3318 :   0 - 0x0
      12'hCF7: dout <= 8'b00000000; // 3319 :   0 - 0x0
      12'hCF8: dout <= 8'b00000000; // 3320 :   0 - 0x0 -- plane 1
      12'hCF9: dout <= 8'b00000000; // 3321 :   0 - 0x0
      12'hCFA: dout <= 8'b00000000; // 3322 :   0 - 0x0
      12'hCFB: dout <= 8'b00000000; // 3323 :   0 - 0x0
      12'hCFC: dout <= 8'b00000000; // 3324 :   0 - 0x0
      12'hCFD: dout <= 8'b00000000; // 3325 :   0 - 0x0
      12'hCFE: dout <= 8'b00000000; // 3326 :   0 - 0x0
      12'hCFF: dout <= 8'b00000000; // 3327 :   0 - 0x0
      12'hD00: dout <= 8'b00000000; // 3328 :   0 - 0x0 -- Background 0xd0
      12'hD01: dout <= 8'b00000000; // 3329 :   0 - 0x0
      12'hD02: dout <= 8'b00000000; // 3330 :   0 - 0x0
      12'hD03: dout <= 8'b00000000; // 3331 :   0 - 0x0
      12'hD04: dout <= 8'b00000000; // 3332 :   0 - 0x0
      12'hD05: dout <= 8'b00000000; // 3333 :   0 - 0x0
      12'hD06: dout <= 8'b00000000; // 3334 :   0 - 0x0
      12'hD07: dout <= 8'b00000000; // 3335 :   0 - 0x0
      12'hD08: dout <= 8'b00000000; // 3336 :   0 - 0x0 -- plane 1
      12'hD09: dout <= 8'b00000000; // 3337 :   0 - 0x0
      12'hD0A: dout <= 8'b00000000; // 3338 :   0 - 0x0
      12'hD0B: dout <= 8'b00000000; // 3339 :   0 - 0x0
      12'hD0C: dout <= 8'b00000000; // 3340 :   0 - 0x0
      12'hD0D: dout <= 8'b00000000; // 3341 :   0 - 0x0
      12'hD0E: dout <= 8'b00000000; // 3342 :   0 - 0x0
      12'hD0F: dout <= 8'b00000000; // 3343 :   0 - 0x0
      12'hD10: dout <= 8'b00000000; // 3344 :   0 - 0x0 -- Background 0xd1
      12'hD11: dout <= 8'b00000000; // 3345 :   0 - 0x0
      12'hD12: dout <= 8'b00000000; // 3346 :   0 - 0x0
      12'hD13: dout <= 8'b00000000; // 3347 :   0 - 0x0
      12'hD14: dout <= 8'b00000000; // 3348 :   0 - 0x0
      12'hD15: dout <= 8'b00000000; // 3349 :   0 - 0x0
      12'hD16: dout <= 8'b00000000; // 3350 :   0 - 0x0
      12'hD17: dout <= 8'b00000000; // 3351 :   0 - 0x0
      12'hD18: dout <= 8'b00000000; // 3352 :   0 - 0x0 -- plane 1
      12'hD19: dout <= 8'b00000000; // 3353 :   0 - 0x0
      12'hD1A: dout <= 8'b00000000; // 3354 :   0 - 0x0
      12'hD1B: dout <= 8'b00000000; // 3355 :   0 - 0x0
      12'hD1C: dout <= 8'b00000000; // 3356 :   0 - 0x0
      12'hD1D: dout <= 8'b00000000; // 3357 :   0 - 0x0
      12'hD1E: dout <= 8'b00000000; // 3358 :   0 - 0x0
      12'hD1F: dout <= 8'b00000000; // 3359 :   0 - 0x0
      12'hD20: dout <= 8'b00000000; // 3360 :   0 - 0x0 -- Background 0xd2
      12'hD21: dout <= 8'b00000000; // 3361 :   0 - 0x0
      12'hD22: dout <= 8'b00000000; // 3362 :   0 - 0x0
      12'hD23: dout <= 8'b00000000; // 3363 :   0 - 0x0
      12'hD24: dout <= 8'b00000000; // 3364 :   0 - 0x0
      12'hD25: dout <= 8'b00000000; // 3365 :   0 - 0x0
      12'hD26: dout <= 8'b00000000; // 3366 :   0 - 0x0
      12'hD27: dout <= 8'b00000000; // 3367 :   0 - 0x0
      12'hD28: dout <= 8'b00000000; // 3368 :   0 - 0x0 -- plane 1
      12'hD29: dout <= 8'b00000000; // 3369 :   0 - 0x0
      12'hD2A: dout <= 8'b00000000; // 3370 :   0 - 0x0
      12'hD2B: dout <= 8'b00000000; // 3371 :   0 - 0x0
      12'hD2C: dout <= 8'b00000000; // 3372 :   0 - 0x0
      12'hD2D: dout <= 8'b00000000; // 3373 :   0 - 0x0
      12'hD2E: dout <= 8'b00000000; // 3374 :   0 - 0x0
      12'hD2F: dout <= 8'b00000000; // 3375 :   0 - 0x0
      12'hD30: dout <= 8'b00000000; // 3376 :   0 - 0x0 -- Background 0xd3
      12'hD31: dout <= 8'b00000000; // 3377 :   0 - 0x0
      12'hD32: dout <= 8'b00000000; // 3378 :   0 - 0x0
      12'hD33: dout <= 8'b00000000; // 3379 :   0 - 0x0
      12'hD34: dout <= 8'b00000000; // 3380 :   0 - 0x0
      12'hD35: dout <= 8'b00000000; // 3381 :   0 - 0x0
      12'hD36: dout <= 8'b00000000; // 3382 :   0 - 0x0
      12'hD37: dout <= 8'b00000000; // 3383 :   0 - 0x0
      12'hD38: dout <= 8'b00000000; // 3384 :   0 - 0x0 -- plane 1
      12'hD39: dout <= 8'b00000000; // 3385 :   0 - 0x0
      12'hD3A: dout <= 8'b00000000; // 3386 :   0 - 0x0
      12'hD3B: dout <= 8'b00000000; // 3387 :   0 - 0x0
      12'hD3C: dout <= 8'b00000000; // 3388 :   0 - 0x0
      12'hD3D: dout <= 8'b00000000; // 3389 :   0 - 0x0
      12'hD3E: dout <= 8'b00000000; // 3390 :   0 - 0x0
      12'hD3F: dout <= 8'b00000000; // 3391 :   0 - 0x0
      12'hD40: dout <= 8'b00000000; // 3392 :   0 - 0x0 -- Background 0xd4
      12'hD41: dout <= 8'b00000000; // 3393 :   0 - 0x0
      12'hD42: dout <= 8'b00000000; // 3394 :   0 - 0x0
      12'hD43: dout <= 8'b00000000; // 3395 :   0 - 0x0
      12'hD44: dout <= 8'b00000000; // 3396 :   0 - 0x0
      12'hD45: dout <= 8'b00000000; // 3397 :   0 - 0x0
      12'hD46: dout <= 8'b00000000; // 3398 :   0 - 0x0
      12'hD47: dout <= 8'b00000000; // 3399 :   0 - 0x0
      12'hD48: dout <= 8'b00000000; // 3400 :   0 - 0x0 -- plane 1
      12'hD49: dout <= 8'b00000000; // 3401 :   0 - 0x0
      12'hD4A: dout <= 8'b00000000; // 3402 :   0 - 0x0
      12'hD4B: dout <= 8'b00000000; // 3403 :   0 - 0x0
      12'hD4C: dout <= 8'b00000000; // 3404 :   0 - 0x0
      12'hD4D: dout <= 8'b00000000; // 3405 :   0 - 0x0
      12'hD4E: dout <= 8'b00000000; // 3406 :   0 - 0x0
      12'hD4F: dout <= 8'b00000000; // 3407 :   0 - 0x0
      12'hD50: dout <= 8'b00000000; // 3408 :   0 - 0x0 -- Background 0xd5
      12'hD51: dout <= 8'b00000000; // 3409 :   0 - 0x0
      12'hD52: dout <= 8'b00000000; // 3410 :   0 - 0x0
      12'hD53: dout <= 8'b00000000; // 3411 :   0 - 0x0
      12'hD54: dout <= 8'b00000000; // 3412 :   0 - 0x0
      12'hD55: dout <= 8'b00000000; // 3413 :   0 - 0x0
      12'hD56: dout <= 8'b00000000; // 3414 :   0 - 0x0
      12'hD57: dout <= 8'b00000000; // 3415 :   0 - 0x0
      12'hD58: dout <= 8'b00000000; // 3416 :   0 - 0x0 -- plane 1
      12'hD59: dout <= 8'b00000000; // 3417 :   0 - 0x0
      12'hD5A: dout <= 8'b00000000; // 3418 :   0 - 0x0
      12'hD5B: dout <= 8'b00000000; // 3419 :   0 - 0x0
      12'hD5C: dout <= 8'b00000000; // 3420 :   0 - 0x0
      12'hD5D: dout <= 8'b00000000; // 3421 :   0 - 0x0
      12'hD5E: dout <= 8'b00000000; // 3422 :   0 - 0x0
      12'hD5F: dout <= 8'b00000000; // 3423 :   0 - 0x0
      12'hD60: dout <= 8'b00000000; // 3424 :   0 - 0x0 -- Background 0xd6
      12'hD61: dout <= 8'b00000000; // 3425 :   0 - 0x0
      12'hD62: dout <= 8'b00000000; // 3426 :   0 - 0x0
      12'hD63: dout <= 8'b00000000; // 3427 :   0 - 0x0
      12'hD64: dout <= 8'b00000000; // 3428 :   0 - 0x0
      12'hD65: dout <= 8'b00000000; // 3429 :   0 - 0x0
      12'hD66: dout <= 8'b00000000; // 3430 :   0 - 0x0
      12'hD67: dout <= 8'b00000000; // 3431 :   0 - 0x0
      12'hD68: dout <= 8'b00000000; // 3432 :   0 - 0x0 -- plane 1
      12'hD69: dout <= 8'b00000000; // 3433 :   0 - 0x0
      12'hD6A: dout <= 8'b00000000; // 3434 :   0 - 0x0
      12'hD6B: dout <= 8'b00000000; // 3435 :   0 - 0x0
      12'hD6C: dout <= 8'b00000000; // 3436 :   0 - 0x0
      12'hD6D: dout <= 8'b00000000; // 3437 :   0 - 0x0
      12'hD6E: dout <= 8'b00000000; // 3438 :   0 - 0x0
      12'hD6F: dout <= 8'b00000000; // 3439 :   0 - 0x0
      12'hD70: dout <= 8'b00000000; // 3440 :   0 - 0x0 -- Background 0xd7
      12'hD71: dout <= 8'b00000000; // 3441 :   0 - 0x0
      12'hD72: dout <= 8'b00000000; // 3442 :   0 - 0x0
      12'hD73: dout <= 8'b00000000; // 3443 :   0 - 0x0
      12'hD74: dout <= 8'b00000000; // 3444 :   0 - 0x0
      12'hD75: dout <= 8'b00000000; // 3445 :   0 - 0x0
      12'hD76: dout <= 8'b00000000; // 3446 :   0 - 0x0
      12'hD77: dout <= 8'b00000000; // 3447 :   0 - 0x0
      12'hD78: dout <= 8'b00000000; // 3448 :   0 - 0x0 -- plane 1
      12'hD79: dout <= 8'b00000000; // 3449 :   0 - 0x0
      12'hD7A: dout <= 8'b00000000; // 3450 :   0 - 0x0
      12'hD7B: dout <= 8'b00000000; // 3451 :   0 - 0x0
      12'hD7C: dout <= 8'b00000000; // 3452 :   0 - 0x0
      12'hD7D: dout <= 8'b00000000; // 3453 :   0 - 0x0
      12'hD7E: dout <= 8'b00000000; // 3454 :   0 - 0x0
      12'hD7F: dout <= 8'b00000000; // 3455 :   0 - 0x0
      12'hD80: dout <= 8'b00000000; // 3456 :   0 - 0x0 -- Background 0xd8
      12'hD81: dout <= 8'b00000000; // 3457 :   0 - 0x0
      12'hD82: dout <= 8'b00000000; // 3458 :   0 - 0x0
      12'hD83: dout <= 8'b00000000; // 3459 :   0 - 0x0
      12'hD84: dout <= 8'b00000000; // 3460 :   0 - 0x0
      12'hD85: dout <= 8'b00000000; // 3461 :   0 - 0x0
      12'hD86: dout <= 8'b00000000; // 3462 :   0 - 0x0
      12'hD87: dout <= 8'b00000000; // 3463 :   0 - 0x0
      12'hD88: dout <= 8'b00000000; // 3464 :   0 - 0x0 -- plane 1
      12'hD89: dout <= 8'b00000000; // 3465 :   0 - 0x0
      12'hD8A: dout <= 8'b00000000; // 3466 :   0 - 0x0
      12'hD8B: dout <= 8'b00000000; // 3467 :   0 - 0x0
      12'hD8C: dout <= 8'b00000000; // 3468 :   0 - 0x0
      12'hD8D: dout <= 8'b00000000; // 3469 :   0 - 0x0
      12'hD8E: dout <= 8'b00000000; // 3470 :   0 - 0x0
      12'hD8F: dout <= 8'b00000000; // 3471 :   0 - 0x0
      12'hD90: dout <= 8'b00000000; // 3472 :   0 - 0x0 -- Background 0xd9
      12'hD91: dout <= 8'b00000000; // 3473 :   0 - 0x0
      12'hD92: dout <= 8'b00000000; // 3474 :   0 - 0x0
      12'hD93: dout <= 8'b00000000; // 3475 :   0 - 0x0
      12'hD94: dout <= 8'b00000000; // 3476 :   0 - 0x0
      12'hD95: dout <= 8'b00000000; // 3477 :   0 - 0x0
      12'hD96: dout <= 8'b00000000; // 3478 :   0 - 0x0
      12'hD97: dout <= 8'b00000000; // 3479 :   0 - 0x0
      12'hD98: dout <= 8'b00000000; // 3480 :   0 - 0x0 -- plane 1
      12'hD99: dout <= 8'b00000000; // 3481 :   0 - 0x0
      12'hD9A: dout <= 8'b00000000; // 3482 :   0 - 0x0
      12'hD9B: dout <= 8'b00000000; // 3483 :   0 - 0x0
      12'hD9C: dout <= 8'b00000000; // 3484 :   0 - 0x0
      12'hD9D: dout <= 8'b00000000; // 3485 :   0 - 0x0
      12'hD9E: dout <= 8'b00000000; // 3486 :   0 - 0x0
      12'hD9F: dout <= 8'b00000000; // 3487 :   0 - 0x0
      12'hDA0: dout <= 8'b00000000; // 3488 :   0 - 0x0 -- Background 0xda
      12'hDA1: dout <= 8'b00000000; // 3489 :   0 - 0x0
      12'hDA2: dout <= 8'b00000000; // 3490 :   0 - 0x0
      12'hDA3: dout <= 8'b00000000; // 3491 :   0 - 0x0
      12'hDA4: dout <= 8'b00000000; // 3492 :   0 - 0x0
      12'hDA5: dout <= 8'b00000000; // 3493 :   0 - 0x0
      12'hDA6: dout <= 8'b00000000; // 3494 :   0 - 0x0
      12'hDA7: dout <= 8'b00000000; // 3495 :   0 - 0x0
      12'hDA8: dout <= 8'b00000000; // 3496 :   0 - 0x0 -- plane 1
      12'hDA9: dout <= 8'b00000000; // 3497 :   0 - 0x0
      12'hDAA: dout <= 8'b00000000; // 3498 :   0 - 0x0
      12'hDAB: dout <= 8'b00000000; // 3499 :   0 - 0x0
      12'hDAC: dout <= 8'b00000000; // 3500 :   0 - 0x0
      12'hDAD: dout <= 8'b00000000; // 3501 :   0 - 0x0
      12'hDAE: dout <= 8'b00000000; // 3502 :   0 - 0x0
      12'hDAF: dout <= 8'b00000000; // 3503 :   0 - 0x0
      12'hDB0: dout <= 8'b00000000; // 3504 :   0 - 0x0 -- Background 0xdb
      12'hDB1: dout <= 8'b00000000; // 3505 :   0 - 0x0
      12'hDB2: dout <= 8'b00000000; // 3506 :   0 - 0x0
      12'hDB3: dout <= 8'b00000000; // 3507 :   0 - 0x0
      12'hDB4: dout <= 8'b00000000; // 3508 :   0 - 0x0
      12'hDB5: dout <= 8'b00000000; // 3509 :   0 - 0x0
      12'hDB6: dout <= 8'b00000000; // 3510 :   0 - 0x0
      12'hDB7: dout <= 8'b00000000; // 3511 :   0 - 0x0
      12'hDB8: dout <= 8'b00000000; // 3512 :   0 - 0x0 -- plane 1
      12'hDB9: dout <= 8'b00000000; // 3513 :   0 - 0x0
      12'hDBA: dout <= 8'b00000000; // 3514 :   0 - 0x0
      12'hDBB: dout <= 8'b00000000; // 3515 :   0 - 0x0
      12'hDBC: dout <= 8'b00000000; // 3516 :   0 - 0x0
      12'hDBD: dout <= 8'b00000000; // 3517 :   0 - 0x0
      12'hDBE: dout <= 8'b00000000; // 3518 :   0 - 0x0
      12'hDBF: dout <= 8'b00000000; // 3519 :   0 - 0x0
      12'hDC0: dout <= 8'b00000000; // 3520 :   0 - 0x0 -- Background 0xdc
      12'hDC1: dout <= 8'b00000000; // 3521 :   0 - 0x0
      12'hDC2: dout <= 8'b00000000; // 3522 :   0 - 0x0
      12'hDC3: dout <= 8'b00000000; // 3523 :   0 - 0x0
      12'hDC4: dout <= 8'b00000000; // 3524 :   0 - 0x0
      12'hDC5: dout <= 8'b00000000; // 3525 :   0 - 0x0
      12'hDC6: dout <= 8'b00000000; // 3526 :   0 - 0x0
      12'hDC7: dout <= 8'b00000000; // 3527 :   0 - 0x0
      12'hDC8: dout <= 8'b00000000; // 3528 :   0 - 0x0 -- plane 1
      12'hDC9: dout <= 8'b00000000; // 3529 :   0 - 0x0
      12'hDCA: dout <= 8'b00000000; // 3530 :   0 - 0x0
      12'hDCB: dout <= 8'b00000000; // 3531 :   0 - 0x0
      12'hDCC: dout <= 8'b00000000; // 3532 :   0 - 0x0
      12'hDCD: dout <= 8'b00000000; // 3533 :   0 - 0x0
      12'hDCE: dout <= 8'b00000000; // 3534 :   0 - 0x0
      12'hDCF: dout <= 8'b00000000; // 3535 :   0 - 0x0
      12'hDD0: dout <= 8'b11100111; // 3536 : 231 - 0xe7 -- Background 0xdd
      12'hDD1: dout <= 8'b11100111; // 3537 : 231 - 0xe7
      12'hDD2: dout <= 8'b11100011; // 3538 : 227 - 0xe3
      12'hDD3: dout <= 8'b11100000; // 3539 : 224 - 0xe0
      12'hDD4: dout <= 8'b11110000; // 3540 : 240 - 0xf0
      12'hDD5: dout <= 8'b11111111; // 3541 : 255 - 0xff
      12'hDD6: dout <= 8'b01111111; // 3542 : 127 - 0x7f
      12'hDD7: dout <= 8'b00111111; // 3543 :  63 - 0x3f
      12'hDD8: dout <= 8'b00011000; // 3544 :  24 - 0x18 -- plane 1
      12'hDD9: dout <= 8'b00011000; // 3545 :  24 - 0x18
      12'hDDA: dout <= 8'b00011100; // 3546 :  28 - 0x1c
      12'hDDB: dout <= 8'b00011111; // 3547 :  31 - 0x1f
      12'hDDC: dout <= 8'b00001111; // 3548 :  15 - 0xf
      12'hDDD: dout <= 8'b00000000; // 3549 :   0 - 0x0
      12'hDDE: dout <= 8'b10000000; // 3550 : 128 - 0x80
      12'hDDF: dout <= 8'b11000000; // 3551 : 192 - 0xc0
      12'hDE0: dout <= 8'b11100111; // 3552 : 231 - 0xe7 -- Background 0xde
      12'hDE1: dout <= 8'b11100111; // 3553 : 231 - 0xe7
      12'hDE2: dout <= 8'b11000111; // 3554 : 199 - 0xc7
      12'hDE3: dout <= 8'b00000111; // 3555 :   7 - 0x7
      12'hDE4: dout <= 8'b00001111; // 3556 :  15 - 0xf
      12'hDE5: dout <= 8'b11111111; // 3557 : 255 - 0xff
      12'hDE6: dout <= 8'b11111110; // 3558 : 254 - 0xfe
      12'hDE7: dout <= 8'b11111100; // 3559 : 252 - 0xfc
      12'hDE8: dout <= 8'b00011000; // 3560 :  24 - 0x18 -- plane 1
      12'hDE9: dout <= 8'b00011000; // 3561 :  24 - 0x18
      12'hDEA: dout <= 8'b00111000; // 3562 :  56 - 0x38
      12'hDEB: dout <= 8'b11111000; // 3563 : 248 - 0xf8
      12'hDEC: dout <= 8'b11110000; // 3564 : 240 - 0xf0
      12'hDED: dout <= 8'b00000000; // 3565 :   0 - 0x0
      12'hDEE: dout <= 8'b00000001; // 3566 :   1 - 0x1
      12'hDEF: dout <= 8'b00000011; // 3567 :   3 - 0x3
      12'hDF0: dout <= 8'b00000000; // 3568 :   0 - 0x0 -- Background 0xdf
      12'hDF1: dout <= 8'b00000000; // 3569 :   0 - 0x0
      12'hDF2: dout <= 8'b00000000; // 3570 :   0 - 0x0
      12'hDF3: dout <= 8'b00000000; // 3571 :   0 - 0x0
      12'hDF4: dout <= 8'b00000000; // 3572 :   0 - 0x0
      12'hDF5: dout <= 8'b00000000; // 3573 :   0 - 0x0
      12'hDF6: dout <= 8'b00000000; // 3574 :   0 - 0x0
      12'hDF7: dout <= 8'b00000000; // 3575 :   0 - 0x0
      12'hDF8: dout <= 8'b00000000; // 3576 :   0 - 0x0 -- plane 1
      12'hDF9: dout <= 8'b00000000; // 3577 :   0 - 0x0
      12'hDFA: dout <= 8'b00000000; // 3578 :   0 - 0x0
      12'hDFB: dout <= 8'b00000000; // 3579 :   0 - 0x0
      12'hDFC: dout <= 8'b00000000; // 3580 :   0 - 0x0
      12'hDFD: dout <= 8'b00000000; // 3581 :   0 - 0x0
      12'hDFE: dout <= 8'b00000000; // 3582 :   0 - 0x0
      12'hDFF: dout <= 8'b00000000; // 3583 :   0 - 0x0
      12'hE00: dout <= 8'b00000000; // 3584 :   0 - 0x0 -- Background 0xe0
      12'hE01: dout <= 8'b00000000; // 3585 :   0 - 0x0
      12'hE02: dout <= 8'b00000000; // 3586 :   0 - 0x0
      12'hE03: dout <= 8'b00000000; // 3587 :   0 - 0x0
      12'hE04: dout <= 8'b00000000; // 3588 :   0 - 0x0
      12'hE05: dout <= 8'b00000000; // 3589 :   0 - 0x0
      12'hE06: dout <= 8'b00000000; // 3590 :   0 - 0x0
      12'hE07: dout <= 8'b00000000; // 3591 :   0 - 0x0
      12'hE08: dout <= 8'b00000000; // 3592 :   0 - 0x0 -- plane 1
      12'hE09: dout <= 8'b00000000; // 3593 :   0 - 0x0
      12'hE0A: dout <= 8'b00000000; // 3594 :   0 - 0x0
      12'hE0B: dout <= 8'b00000000; // 3595 :   0 - 0x0
      12'hE0C: dout <= 8'b00000000; // 3596 :   0 - 0x0
      12'hE0D: dout <= 8'b00000000; // 3597 :   0 - 0x0
      12'hE0E: dout <= 8'b00000000; // 3598 :   0 - 0x0
      12'hE0F: dout <= 8'b00000000; // 3599 :   0 - 0x0
      12'hE10: dout <= 8'b00000000; // 3600 :   0 - 0x0 -- Background 0xe1
      12'hE11: dout <= 8'b00000000; // 3601 :   0 - 0x0
      12'hE12: dout <= 8'b00000000; // 3602 :   0 - 0x0
      12'hE13: dout <= 8'b00000000; // 3603 :   0 - 0x0
      12'hE14: dout <= 8'b00000000; // 3604 :   0 - 0x0
      12'hE15: dout <= 8'b00000000; // 3605 :   0 - 0x0
      12'hE16: dout <= 8'b00000000; // 3606 :   0 - 0x0
      12'hE17: dout <= 8'b00000000; // 3607 :   0 - 0x0
      12'hE18: dout <= 8'b00000000; // 3608 :   0 - 0x0 -- plane 1
      12'hE19: dout <= 8'b00000000; // 3609 :   0 - 0x0
      12'hE1A: dout <= 8'b00000000; // 3610 :   0 - 0x0
      12'hE1B: dout <= 8'b00000000; // 3611 :   0 - 0x0
      12'hE1C: dout <= 8'b00000000; // 3612 :   0 - 0x0
      12'hE1D: dout <= 8'b00000000; // 3613 :   0 - 0x0
      12'hE1E: dout <= 8'b00000000; // 3614 :   0 - 0x0
      12'hE1F: dout <= 8'b00000000; // 3615 :   0 - 0x0
      12'hE20: dout <= 8'b00000000; // 3616 :   0 - 0x0 -- Background 0xe2
      12'hE21: dout <= 8'b00000000; // 3617 :   0 - 0x0
      12'hE22: dout <= 8'b00000000; // 3618 :   0 - 0x0
      12'hE23: dout <= 8'b00000000; // 3619 :   0 - 0x0
      12'hE24: dout <= 8'b00000000; // 3620 :   0 - 0x0
      12'hE25: dout <= 8'b00000000; // 3621 :   0 - 0x0
      12'hE26: dout <= 8'b00000000; // 3622 :   0 - 0x0
      12'hE27: dout <= 8'b00000000; // 3623 :   0 - 0x0
      12'hE28: dout <= 8'b00000000; // 3624 :   0 - 0x0 -- plane 1
      12'hE29: dout <= 8'b00000000; // 3625 :   0 - 0x0
      12'hE2A: dout <= 8'b00000000; // 3626 :   0 - 0x0
      12'hE2B: dout <= 8'b00000000; // 3627 :   0 - 0x0
      12'hE2C: dout <= 8'b00000000; // 3628 :   0 - 0x0
      12'hE2D: dout <= 8'b00000000; // 3629 :   0 - 0x0
      12'hE2E: dout <= 8'b00000000; // 3630 :   0 - 0x0
      12'hE2F: dout <= 8'b00000000; // 3631 :   0 - 0x0
      12'hE30: dout <= 8'b00000000; // 3632 :   0 - 0x0 -- Background 0xe3
      12'hE31: dout <= 8'b00000000; // 3633 :   0 - 0x0
      12'hE32: dout <= 8'b00000000; // 3634 :   0 - 0x0
      12'hE33: dout <= 8'b00000000; // 3635 :   0 - 0x0
      12'hE34: dout <= 8'b00000000; // 3636 :   0 - 0x0
      12'hE35: dout <= 8'b00000000; // 3637 :   0 - 0x0
      12'hE36: dout <= 8'b00000000; // 3638 :   0 - 0x0
      12'hE37: dout <= 8'b00000000; // 3639 :   0 - 0x0
      12'hE38: dout <= 8'b00000000; // 3640 :   0 - 0x0 -- plane 1
      12'hE39: dout <= 8'b00000000; // 3641 :   0 - 0x0
      12'hE3A: dout <= 8'b00000000; // 3642 :   0 - 0x0
      12'hE3B: dout <= 8'b00000000; // 3643 :   0 - 0x0
      12'hE3C: dout <= 8'b00000000; // 3644 :   0 - 0x0
      12'hE3D: dout <= 8'b00000000; // 3645 :   0 - 0x0
      12'hE3E: dout <= 8'b00000000; // 3646 :   0 - 0x0
      12'hE3F: dout <= 8'b00000000; // 3647 :   0 - 0x0
      12'hE40: dout <= 8'b00000000; // 3648 :   0 - 0x0 -- Background 0xe4
      12'hE41: dout <= 8'b00000000; // 3649 :   0 - 0x0
      12'hE42: dout <= 8'b00000000; // 3650 :   0 - 0x0
      12'hE43: dout <= 8'b00000000; // 3651 :   0 - 0x0
      12'hE44: dout <= 8'b00000000; // 3652 :   0 - 0x0
      12'hE45: dout <= 8'b00000000; // 3653 :   0 - 0x0
      12'hE46: dout <= 8'b00000000; // 3654 :   0 - 0x0
      12'hE47: dout <= 8'b00000000; // 3655 :   0 - 0x0
      12'hE48: dout <= 8'b00000000; // 3656 :   0 - 0x0 -- plane 1
      12'hE49: dout <= 8'b00000000; // 3657 :   0 - 0x0
      12'hE4A: dout <= 8'b00000000; // 3658 :   0 - 0x0
      12'hE4B: dout <= 8'b00000000; // 3659 :   0 - 0x0
      12'hE4C: dout <= 8'b00000000; // 3660 :   0 - 0x0
      12'hE4D: dout <= 8'b00000000; // 3661 :   0 - 0x0
      12'hE4E: dout <= 8'b00000000; // 3662 :   0 - 0x0
      12'hE4F: dout <= 8'b00000000; // 3663 :   0 - 0x0
      12'hE50: dout <= 8'b01111111; // 3664 : 127 - 0x7f -- Background 0xe5
      12'hE51: dout <= 8'b11111111; // 3665 : 255 - 0xff
      12'hE52: dout <= 8'b11111111; // 3666 : 255 - 0xff
      12'hE53: dout <= 8'b11100000; // 3667 : 224 - 0xe0
      12'hE54: dout <= 8'b11100000; // 3668 : 224 - 0xe0
      12'hE55: dout <= 8'b11100000; // 3669 : 224 - 0xe0
      12'hE56: dout <= 8'b11100000; // 3670 : 224 - 0xe0
      12'hE57: dout <= 8'b11100001; // 3671 : 225 - 0xe1
      12'hE58: dout <= 8'b00000000; // 3672 :   0 - 0x0 -- plane 1
      12'hE59: dout <= 8'b00000000; // 3673 :   0 - 0x0
      12'hE5A: dout <= 8'b00000000; // 3674 :   0 - 0x0
      12'hE5B: dout <= 8'b00000000; // 3675 :   0 - 0x0
      12'hE5C: dout <= 8'b00000000; // 3676 :   0 - 0x0
      12'hE5D: dout <= 8'b00000000; // 3677 :   0 - 0x0
      12'hE5E: dout <= 8'b00000000; // 3678 :   0 - 0x0
      12'hE5F: dout <= 8'b00000000; // 3679 :   0 - 0x0
      12'hE60: dout <= 8'b11111110; // 3680 : 254 - 0xfe -- Background 0xe6
      12'hE61: dout <= 8'b11111111; // 3681 : 255 - 0xff
      12'hE62: dout <= 8'b11111111; // 3682 : 255 - 0xff
      12'hE63: dout <= 8'b00000111; // 3683 :   7 - 0x7
      12'hE64: dout <= 8'b00000111; // 3684 :   7 - 0x7
      12'hE65: dout <= 8'b00000111; // 3685 :   7 - 0x7
      12'hE66: dout <= 8'b00000111; // 3686 :   7 - 0x7
      12'hE67: dout <= 8'b10000111; // 3687 : 135 - 0x87
      12'hE68: dout <= 8'b00000000; // 3688 :   0 - 0x0 -- plane 1
      12'hE69: dout <= 8'b00000000; // 3689 :   0 - 0x0
      12'hE6A: dout <= 8'b00000000; // 3690 :   0 - 0x0
      12'hE6B: dout <= 8'b00000000; // 3691 :   0 - 0x0
      12'hE6C: dout <= 8'b00000000; // 3692 :   0 - 0x0
      12'hE6D: dout <= 8'b00000000; // 3693 :   0 - 0x0
      12'hE6E: dout <= 8'b00000000; // 3694 :   0 - 0x0
      12'hE6F: dout <= 8'b00000000; // 3695 :   0 - 0x0
      12'hE70: dout <= 8'b00011111; // 3696 :  31 - 0x1f -- Background 0xe7
      12'hE71: dout <= 8'b00100000; // 3697 :  32 - 0x20
      12'hE72: dout <= 8'b01000000; // 3698 :  64 - 0x40
      12'hE73: dout <= 8'b10000000; // 3699 : 128 - 0x80
      12'hE74: dout <= 8'b10000000; // 3700 : 128 - 0x80
      12'hE75: dout <= 8'b10000011; // 3701 : 131 - 0x83
      12'hE76: dout <= 8'b10000111; // 3702 : 135 - 0x87
      12'hE77: dout <= 8'b10000111; // 3703 : 135 - 0x87
      12'hE78: dout <= 8'b11100000; // 3704 : 224 - 0xe0 -- plane 1
      12'hE79: dout <= 8'b11000000; // 3705 : 192 - 0xc0
      12'hE7A: dout <= 8'b10000000; // 3706 : 128 - 0x80
      12'hE7B: dout <= 8'b00000000; // 3707 :   0 - 0x0
      12'hE7C: dout <= 8'b00000000; // 3708 :   0 - 0x0
      12'hE7D: dout <= 8'b00000000; // 3709 :   0 - 0x0
      12'hE7E: dout <= 8'b00000000; // 3710 :   0 - 0x0
      12'hE7F: dout <= 8'b00000000; // 3711 :   0 - 0x0
      12'hE80: dout <= 8'b11111000; // 3712 : 248 - 0xf8 -- Background 0xe8
      12'hE81: dout <= 8'b00000100; // 3713 :   4 - 0x4
      12'hE82: dout <= 8'b00000010; // 3714 :   2 - 0x2
      12'hE83: dout <= 8'b00000001; // 3715 :   1 - 0x1
      12'hE84: dout <= 8'b00000001; // 3716 :   1 - 0x1
      12'hE85: dout <= 8'b11000001; // 3717 : 193 - 0xc1
      12'hE86: dout <= 8'b11100001; // 3718 : 225 - 0xe1
      12'hE87: dout <= 8'b11100001; // 3719 : 225 - 0xe1
      12'hE88: dout <= 8'b00000111; // 3720 :   7 - 0x7 -- plane 1
      12'hE89: dout <= 8'b00000011; // 3721 :   3 - 0x3
      12'hE8A: dout <= 8'b00000001; // 3722 :   1 - 0x1
      12'hE8B: dout <= 8'b00000000; // 3723 :   0 - 0x0
      12'hE8C: dout <= 8'b00000000; // 3724 :   0 - 0x0
      12'hE8D: dout <= 8'b00000000; // 3725 :   0 - 0x0
      12'hE8E: dout <= 8'b00000000; // 3726 :   0 - 0x0
      12'hE8F: dout <= 8'b00000000; // 3727 :   0 - 0x0
      12'hE90: dout <= 8'b00000000; // 3728 :   0 - 0x0 -- Background 0xe9
      12'hE91: dout <= 8'b00000000; // 3729 :   0 - 0x0
      12'hE92: dout <= 8'b00001000; // 3730 :   8 - 0x8
      12'hE93: dout <= 8'b00010100; // 3731 :  20 - 0x14
      12'hE94: dout <= 8'b00000000; // 3732 :   0 - 0x0
      12'hE95: dout <= 8'b00000000; // 3733 :   0 - 0x0
      12'hE96: dout <= 8'b01000000; // 3734 :  64 - 0x40
      12'hE97: dout <= 8'b10100000; // 3735 : 160 - 0xa0
      12'hE98: dout <= 8'b11111111; // 3736 : 255 - 0xff -- plane 1
      12'hE99: dout <= 8'b11111111; // 3737 : 255 - 0xff
      12'hE9A: dout <= 8'b11111111; // 3738 : 255 - 0xff
      12'hE9B: dout <= 8'b11111111; // 3739 : 255 - 0xff
      12'hE9C: dout <= 8'b11111111; // 3740 : 255 - 0xff
      12'hE9D: dout <= 8'b11111111; // 3741 : 255 - 0xff
      12'hE9E: dout <= 8'b11111111; // 3742 : 255 - 0xff
      12'hE9F: dout <= 8'b11111111; // 3743 : 255 - 0xff
      12'hEA0: dout <= 8'b01000000; // 3744 :  64 - 0x40 -- Background 0xea
      12'hEA1: dout <= 8'b10100010; // 3745 : 162 - 0xa2
      12'hEA2: dout <= 8'b00000101; // 3746 :   5 - 0x5
      12'hEA3: dout <= 8'b00000000; // 3747 :   0 - 0x0
      12'hEA4: dout <= 8'b00000000; // 3748 :   0 - 0x0
      12'hEA5: dout <= 8'b00010000; // 3749 :  16 - 0x10
      12'hEA6: dout <= 8'b00101000; // 3750 :  40 - 0x28
      12'hEA7: dout <= 8'b00000000; // 3751 :   0 - 0x0
      12'hEA8: dout <= 8'b11111111; // 3752 : 255 - 0xff -- plane 1
      12'hEA9: dout <= 8'b11111111; // 3753 : 255 - 0xff
      12'hEAA: dout <= 8'b11111111; // 3754 : 255 - 0xff
      12'hEAB: dout <= 8'b11111111; // 3755 : 255 - 0xff
      12'hEAC: dout <= 8'b11111111; // 3756 : 255 - 0xff
      12'hEAD: dout <= 8'b11111111; // 3757 : 255 - 0xff
      12'hEAE: dout <= 8'b11111111; // 3758 : 255 - 0xff
      12'hEAF: dout <= 8'b11111111; // 3759 : 255 - 0xff
      12'hEB0: dout <= 8'b11111111; // 3760 : 255 - 0xff -- Background 0xeb
      12'hEB1: dout <= 8'b11111111; // 3761 : 255 - 0xff
      12'hEB2: dout <= 8'b11111111; // 3762 : 255 - 0xff
      12'hEB3: dout <= 8'b00000000; // 3763 :   0 - 0x0
      12'hEB4: dout <= 8'b00000000; // 3764 :   0 - 0x0
      12'hEB5: dout <= 8'b00000000; // 3765 :   0 - 0x0
      12'hEB6: dout <= 8'b00000000; // 3766 :   0 - 0x0
      12'hEB7: dout <= 8'b11111111; // 3767 : 255 - 0xff
      12'hEB8: dout <= 8'b00000000; // 3768 :   0 - 0x0 -- plane 1
      12'hEB9: dout <= 8'b00000000; // 3769 :   0 - 0x0
      12'hEBA: dout <= 8'b00000000; // 3770 :   0 - 0x0
      12'hEBB: dout <= 8'b00000000; // 3771 :   0 - 0x0
      12'hEBC: dout <= 8'b00000000; // 3772 :   0 - 0x0
      12'hEBD: dout <= 8'b00000000; // 3773 :   0 - 0x0
      12'hEBE: dout <= 8'b00000000; // 3774 :   0 - 0x0
      12'hEBF: dout <= 8'b00000000; // 3775 :   0 - 0x0
      12'hEC0: dout <= 8'b11100001; // 3776 : 225 - 0xe1 -- Background 0xec
      12'hEC1: dout <= 8'b11100001; // 3777 : 225 - 0xe1
      12'hEC2: dout <= 8'b11100001; // 3778 : 225 - 0xe1
      12'hEC3: dout <= 8'b11100001; // 3779 : 225 - 0xe1
      12'hEC4: dout <= 8'b11100001; // 3780 : 225 - 0xe1
      12'hEC5: dout <= 8'b11100001; // 3781 : 225 - 0xe1
      12'hEC6: dout <= 8'b11100001; // 3782 : 225 - 0xe1
      12'hEC7: dout <= 8'b11100001; // 3783 : 225 - 0xe1
      12'hEC8: dout <= 8'b00000000; // 3784 :   0 - 0x0 -- plane 1
      12'hEC9: dout <= 8'b00000000; // 3785 :   0 - 0x0
      12'hECA: dout <= 8'b00000000; // 3786 :   0 - 0x0
      12'hECB: dout <= 8'b00000000; // 3787 :   0 - 0x0
      12'hECC: dout <= 8'b00000000; // 3788 :   0 - 0x0
      12'hECD: dout <= 8'b00000000; // 3789 :   0 - 0x0
      12'hECE: dout <= 8'b00000000; // 3790 :   0 - 0x0
      12'hECF: dout <= 8'b00000000; // 3791 :   0 - 0x0
      12'hED0: dout <= 8'b11111111; // 3792 : 255 - 0xff -- Background 0xed
      12'hED1: dout <= 8'b11111111; // 3793 : 255 - 0xff
      12'hED2: dout <= 8'b11111111; // 3794 : 255 - 0xff
      12'hED3: dout <= 8'b00000000; // 3795 :   0 - 0x0
      12'hED4: dout <= 8'b00000000; // 3796 :   0 - 0x0
      12'hED5: dout <= 8'b11111111; // 3797 : 255 - 0xff
      12'hED6: dout <= 8'b11111111; // 3798 : 255 - 0xff
      12'hED7: dout <= 8'b11111111; // 3799 : 255 - 0xff
      12'hED8: dout <= 8'b00000000; // 3800 :   0 - 0x0 -- plane 1
      12'hED9: dout <= 8'b00000000; // 3801 :   0 - 0x0
      12'hEDA: dout <= 8'b00000000; // 3802 :   0 - 0x0
      12'hEDB: dout <= 8'b11111111; // 3803 : 255 - 0xff
      12'hEDC: dout <= 8'b11111111; // 3804 : 255 - 0xff
      12'hEDD: dout <= 8'b00000000; // 3805 :   0 - 0x0
      12'hEDE: dout <= 8'b00000000; // 3806 :   0 - 0x0
      12'hEDF: dout <= 8'b00000000; // 3807 :   0 - 0x0
      12'hEE0: dout <= 8'b11100111; // 3808 : 231 - 0xe7 -- Background 0xee
      12'hEE1: dout <= 8'b11100111; // 3809 : 231 - 0xe7
      12'hEE2: dout <= 8'b11100111; // 3810 : 231 - 0xe7
      12'hEE3: dout <= 8'b11100111; // 3811 : 231 - 0xe7
      12'hEE4: dout <= 8'b11100111; // 3812 : 231 - 0xe7
      12'hEE5: dout <= 8'b11100111; // 3813 : 231 - 0xe7
      12'hEE6: dout <= 8'b11100111; // 3814 : 231 - 0xe7
      12'hEE7: dout <= 8'b11100111; // 3815 : 231 - 0xe7
      12'hEE8: dout <= 8'b00011000; // 3816 :  24 - 0x18 -- plane 1
      12'hEE9: dout <= 8'b00011000; // 3817 :  24 - 0x18
      12'hEEA: dout <= 8'b00011000; // 3818 :  24 - 0x18
      12'hEEB: dout <= 8'b00011000; // 3819 :  24 - 0x18
      12'hEEC: dout <= 8'b00011000; // 3820 :  24 - 0x18
      12'hEED: dout <= 8'b00011000; // 3821 :  24 - 0x18
      12'hEEE: dout <= 8'b00011000; // 3822 :  24 - 0x18
      12'hEEF: dout <= 8'b00011000; // 3823 :  24 - 0x18
      12'hEF0: dout <= 8'b11111111; // 3824 : 255 - 0xff -- Background 0xef
      12'hEF1: dout <= 8'b11111111; // 3825 : 255 - 0xff
      12'hEF2: dout <= 8'b11111111; // 3826 : 255 - 0xff
      12'hEF3: dout <= 8'b11111111; // 3827 : 255 - 0xff
      12'hEF4: dout <= 8'b11111111; // 3828 : 255 - 0xff
      12'hEF5: dout <= 8'b11111111; // 3829 : 255 - 0xff
      12'hEF6: dout <= 8'b11111111; // 3830 : 255 - 0xff
      12'hEF7: dout <= 8'b11111111; // 3831 : 255 - 0xff
      12'hEF8: dout <= 8'b00110011; // 3832 :  51 - 0x33 -- plane 1
      12'hEF9: dout <= 8'b00110011; // 3833 :  51 - 0x33
      12'hEFA: dout <= 8'b11001100; // 3834 : 204 - 0xcc
      12'hEFB: dout <= 8'b11001100; // 3835 : 204 - 0xcc
      12'hEFC: dout <= 8'b00110011; // 3836 :  51 - 0x33
      12'hEFD: dout <= 8'b00110011; // 3837 :  51 - 0x33
      12'hEFE: dout <= 8'b11001100; // 3838 : 204 - 0xcc
      12'hEFF: dout <= 8'b11001100; // 3839 : 204 - 0xcc
      12'hF00: dout <= 8'b00000000; // 3840 :   0 - 0x0 -- Background 0xf0
      12'hF01: dout <= 8'b00000000; // 3841 :   0 - 0x0
      12'hF02: dout <= 8'b00000000; // 3842 :   0 - 0x0
      12'hF03: dout <= 8'b00000000; // 3843 :   0 - 0x0
      12'hF04: dout <= 8'b00000000; // 3844 :   0 - 0x0
      12'hF05: dout <= 8'b00000000; // 3845 :   0 - 0x0
      12'hF06: dout <= 8'b00000000; // 3846 :   0 - 0x0
      12'hF07: dout <= 8'b00000000; // 3847 :   0 - 0x0
      12'hF08: dout <= 8'b00000000; // 3848 :   0 - 0x0 -- plane 1
      12'hF09: dout <= 8'b00000000; // 3849 :   0 - 0x0
      12'hF0A: dout <= 8'b00000000; // 3850 :   0 - 0x0
      12'hF0B: dout <= 8'b00000000; // 3851 :   0 - 0x0
      12'hF0C: dout <= 8'b00000000; // 3852 :   0 - 0x0
      12'hF0D: dout <= 8'b00000000; // 3853 :   0 - 0x0
      12'hF0E: dout <= 8'b00000000; // 3854 :   0 - 0x0
      12'hF0F: dout <= 8'b00000000; // 3855 :   0 - 0x0
      12'hF10: dout <= 8'b00000000; // 3856 :   0 - 0x0 -- Background 0xf1
      12'hF11: dout <= 8'b00000000; // 3857 :   0 - 0x0
      12'hF12: dout <= 8'b00000000; // 3858 :   0 - 0x0
      12'hF13: dout <= 8'b00000000; // 3859 :   0 - 0x0
      12'hF14: dout <= 8'b00000000; // 3860 :   0 - 0x0
      12'hF15: dout <= 8'b00000000; // 3861 :   0 - 0x0
      12'hF16: dout <= 8'b00000000; // 3862 :   0 - 0x0
      12'hF17: dout <= 8'b00000000; // 3863 :   0 - 0x0
      12'hF18: dout <= 8'b00000000; // 3864 :   0 - 0x0 -- plane 1
      12'hF19: dout <= 8'b00000000; // 3865 :   0 - 0x0
      12'hF1A: dout <= 8'b00000000; // 3866 :   0 - 0x0
      12'hF1B: dout <= 8'b00000000; // 3867 :   0 - 0x0
      12'hF1C: dout <= 8'b00000000; // 3868 :   0 - 0x0
      12'hF1D: dout <= 8'b00000000; // 3869 :   0 - 0x0
      12'hF1E: dout <= 8'b00000000; // 3870 :   0 - 0x0
      12'hF1F: dout <= 8'b00000000; // 3871 :   0 - 0x0
      12'hF20: dout <= 8'b00000000; // 3872 :   0 - 0x0 -- Background 0xf2
      12'hF21: dout <= 8'b00000000; // 3873 :   0 - 0x0
      12'hF22: dout <= 8'b00000000; // 3874 :   0 - 0x0
      12'hF23: dout <= 8'b00000000; // 3875 :   0 - 0x0
      12'hF24: dout <= 8'b00000000; // 3876 :   0 - 0x0
      12'hF25: dout <= 8'b00000000; // 3877 :   0 - 0x0
      12'hF26: dout <= 8'b00000000; // 3878 :   0 - 0x0
      12'hF27: dout <= 8'b00000000; // 3879 :   0 - 0x0
      12'hF28: dout <= 8'b00000000; // 3880 :   0 - 0x0 -- plane 1
      12'hF29: dout <= 8'b00000000; // 3881 :   0 - 0x0
      12'hF2A: dout <= 8'b00000000; // 3882 :   0 - 0x0
      12'hF2B: dout <= 8'b00000000; // 3883 :   0 - 0x0
      12'hF2C: dout <= 8'b00000000; // 3884 :   0 - 0x0
      12'hF2D: dout <= 8'b00000000; // 3885 :   0 - 0x0
      12'hF2E: dout <= 8'b00000000; // 3886 :   0 - 0x0
      12'hF2F: dout <= 8'b00000000; // 3887 :   0 - 0x0
      12'hF30: dout <= 8'b00000000; // 3888 :   0 - 0x0 -- Background 0xf3
      12'hF31: dout <= 8'b00000000; // 3889 :   0 - 0x0
      12'hF32: dout <= 8'b00000000; // 3890 :   0 - 0x0
      12'hF33: dout <= 8'b00000000; // 3891 :   0 - 0x0
      12'hF34: dout <= 8'b00000000; // 3892 :   0 - 0x0
      12'hF35: dout <= 8'b00000000; // 3893 :   0 - 0x0
      12'hF36: dout <= 8'b00000000; // 3894 :   0 - 0x0
      12'hF37: dout <= 8'b00000000; // 3895 :   0 - 0x0
      12'hF38: dout <= 8'b00000000; // 3896 :   0 - 0x0 -- plane 1
      12'hF39: dout <= 8'b00000000; // 3897 :   0 - 0x0
      12'hF3A: dout <= 8'b00000000; // 3898 :   0 - 0x0
      12'hF3B: dout <= 8'b00000000; // 3899 :   0 - 0x0
      12'hF3C: dout <= 8'b00000000; // 3900 :   0 - 0x0
      12'hF3D: dout <= 8'b00000000; // 3901 :   0 - 0x0
      12'hF3E: dout <= 8'b00000000; // 3902 :   0 - 0x0
      12'hF3F: dout <= 8'b00000000; // 3903 :   0 - 0x0
      12'hF40: dout <= 8'b11100111; // 3904 : 231 - 0xe7 -- Background 0xf4
      12'hF41: dout <= 8'b10011001; // 3905 : 153 - 0x99
      12'hF42: dout <= 8'b10000001; // 3906 : 129 - 0x81
      12'hF43: dout <= 8'b11000011; // 3907 : 195 - 0xc3
      12'hF44: dout <= 8'b11111111; // 3908 : 255 - 0xff
      12'hF45: dout <= 8'b10111101; // 3909 : 189 - 0xbd
      12'hF46: dout <= 8'b10000001; // 3910 : 129 - 0x81
      12'hF47: dout <= 8'b11000011; // 3911 : 195 - 0xc3
      12'hF48: dout <= 8'b00100100; // 3912 :  36 - 0x24 -- plane 1
      12'hF49: dout <= 8'b00011000; // 3913 :  24 - 0x18
      12'hF4A: dout <= 8'b00000000; // 3914 :   0 - 0x0
      12'hF4B: dout <= 8'b01000010; // 3915 :  66 - 0x42
      12'hF4C: dout <= 8'b01111110; // 3916 : 126 - 0x7e
      12'hF4D: dout <= 8'b00111100; // 3917 :  60 - 0x3c
      12'hF4E: dout <= 8'b00000000; // 3918 :   0 - 0x0
      12'hF4F: dout <= 8'b00000000; // 3919 :   0 - 0x0
      12'hF50: dout <= 8'b11100001; // 3920 : 225 - 0xe1 -- Background 0xf5
      12'hF51: dout <= 8'b11100000; // 3921 : 224 - 0xe0
      12'hF52: dout <= 8'b11100000; // 3922 : 224 - 0xe0
      12'hF53: dout <= 8'b11100000; // 3923 : 224 - 0xe0
      12'hF54: dout <= 8'b11100000; // 3924 : 224 - 0xe0
      12'hF55: dout <= 8'b11111111; // 3925 : 255 - 0xff
      12'hF56: dout <= 8'b11111111; // 3926 : 255 - 0xff
      12'hF57: dout <= 8'b01111111; // 3927 : 127 - 0x7f
      12'hF58: dout <= 8'b00000000; // 3928 :   0 - 0x0 -- plane 1
      12'hF59: dout <= 8'b00000000; // 3929 :   0 - 0x0
      12'hF5A: dout <= 8'b00000000; // 3930 :   0 - 0x0
      12'hF5B: dout <= 8'b00000000; // 3931 :   0 - 0x0
      12'hF5C: dout <= 8'b00000000; // 3932 :   0 - 0x0
      12'hF5D: dout <= 8'b00000000; // 3933 :   0 - 0x0
      12'hF5E: dout <= 8'b00000000; // 3934 :   0 - 0x0
      12'hF5F: dout <= 8'b00000000; // 3935 :   0 - 0x0
      12'hF60: dout <= 8'b10000111; // 3936 : 135 - 0x87 -- Background 0xf6
      12'hF61: dout <= 8'b00000111; // 3937 :   7 - 0x7
      12'hF62: dout <= 8'b00000111; // 3938 :   7 - 0x7
      12'hF63: dout <= 8'b00000111; // 3939 :   7 - 0x7
      12'hF64: dout <= 8'b00000111; // 3940 :   7 - 0x7
      12'hF65: dout <= 8'b11111111; // 3941 : 255 - 0xff
      12'hF66: dout <= 8'b11111111; // 3942 : 255 - 0xff
      12'hF67: dout <= 8'b11111110; // 3943 : 254 - 0xfe
      12'hF68: dout <= 8'b00000000; // 3944 :   0 - 0x0 -- plane 1
      12'hF69: dout <= 8'b00000000; // 3945 :   0 - 0x0
      12'hF6A: dout <= 8'b00000000; // 3946 :   0 - 0x0
      12'hF6B: dout <= 8'b00000000; // 3947 :   0 - 0x0
      12'hF6C: dout <= 8'b00000000; // 3948 :   0 - 0x0
      12'hF6D: dout <= 8'b00000000; // 3949 :   0 - 0x0
      12'hF6E: dout <= 8'b00000000; // 3950 :   0 - 0x0
      12'hF6F: dout <= 8'b00000000; // 3951 :   0 - 0x0
      12'hF70: dout <= 8'b10000111; // 3952 : 135 - 0x87 -- Background 0xf7
      12'hF71: dout <= 8'b10000111; // 3953 : 135 - 0x87
      12'hF72: dout <= 8'b10000011; // 3954 : 131 - 0x83
      12'hF73: dout <= 8'b10000000; // 3955 : 128 - 0x80
      12'hF74: dout <= 8'b10000000; // 3956 : 128 - 0x80
      12'hF75: dout <= 8'b01000000; // 3957 :  64 - 0x40
      12'hF76: dout <= 8'b00100000; // 3958 :  32 - 0x20
      12'hF77: dout <= 8'b00011111; // 3959 :  31 - 0x1f
      12'hF78: dout <= 8'b00000000; // 3960 :   0 - 0x0 -- plane 1
      12'hF79: dout <= 8'b00000000; // 3961 :   0 - 0x0
      12'hF7A: dout <= 8'b00000000; // 3962 :   0 - 0x0
      12'hF7B: dout <= 8'b00000000; // 3963 :   0 - 0x0
      12'hF7C: dout <= 8'b00000000; // 3964 :   0 - 0x0
      12'hF7D: dout <= 8'b10000000; // 3965 : 128 - 0x80
      12'hF7E: dout <= 8'b11000000; // 3966 : 192 - 0xc0
      12'hF7F: dout <= 8'b11100000; // 3967 : 224 - 0xe0
      12'hF80: dout <= 8'b11100001; // 3968 : 225 - 0xe1 -- Background 0xf8
      12'hF81: dout <= 8'b11100001; // 3969 : 225 - 0xe1
      12'hF82: dout <= 8'b11000001; // 3970 : 193 - 0xc1
      12'hF83: dout <= 8'b00000001; // 3971 :   1 - 0x1
      12'hF84: dout <= 8'b00000001; // 3972 :   1 - 0x1
      12'hF85: dout <= 8'b00000010; // 3973 :   2 - 0x2
      12'hF86: dout <= 8'b00000100; // 3974 :   4 - 0x4
      12'hF87: dout <= 8'b11111000; // 3975 : 248 - 0xf8
      12'hF88: dout <= 8'b00000000; // 3976 :   0 - 0x0 -- plane 1
      12'hF89: dout <= 8'b00000000; // 3977 :   0 - 0x0
      12'hF8A: dout <= 8'b00000000; // 3978 :   0 - 0x0
      12'hF8B: dout <= 8'b00000000; // 3979 :   0 - 0x0
      12'hF8C: dout <= 8'b00000000; // 3980 :   0 - 0x0
      12'hF8D: dout <= 8'b00000001; // 3981 :   1 - 0x1
      12'hF8E: dout <= 8'b00000011; // 3982 :   3 - 0x3
      12'hF8F: dout <= 8'b00000111; // 3983 :   7 - 0x7
      12'hF90: dout <= 8'b00000000; // 3984 :   0 - 0x0 -- Background 0xf9
      12'hF91: dout <= 8'b00000010; // 3985 :   2 - 0x2
      12'hF92: dout <= 8'b00000101; // 3986 :   5 - 0x5
      12'hF93: dout <= 8'b00000000; // 3987 :   0 - 0x0
      12'hF94: dout <= 8'b00100000; // 3988 :  32 - 0x20
      12'hF95: dout <= 8'b01010000; // 3989 :  80 - 0x50
      12'hF96: dout <= 8'b00000000; // 3990 :   0 - 0x0
      12'hF97: dout <= 8'b00000000; // 3991 :   0 - 0x0
      12'hF98: dout <= 8'b11111111; // 3992 : 255 - 0xff -- plane 1
      12'hF99: dout <= 8'b11111111; // 3993 : 255 - 0xff
      12'hF9A: dout <= 8'b11111111; // 3994 : 255 - 0xff
      12'hF9B: dout <= 8'b11111111; // 3995 : 255 - 0xff
      12'hF9C: dout <= 8'b11111111; // 3996 : 255 - 0xff
      12'hF9D: dout <= 8'b11111111; // 3997 : 255 - 0xff
      12'hF9E: dout <= 8'b11111111; // 3998 : 255 - 0xff
      12'hF9F: dout <= 8'b11111111; // 3999 : 255 - 0xff
      12'hFA0: dout <= 8'b00000000; // 4000 :   0 - 0x0 -- Background 0xfa
      12'hFA1: dout <= 8'b00000000; // 4001 :   0 - 0x0
      12'hFA2: dout <= 8'b00000000; // 4002 :   0 - 0x0
      12'hFA3: dout <= 8'b00000000; // 4003 :   0 - 0x0
      12'hFA4: dout <= 8'b00000000; // 4004 :   0 - 0x0
      12'hFA5: dout <= 8'b00000000; // 4005 :   0 - 0x0
      12'hFA6: dout <= 8'b00000000; // 4006 :   0 - 0x0
      12'hFA7: dout <= 8'b00000000; // 4007 :   0 - 0x0
      12'hFA8: dout <= 8'b11111111; // 4008 : 255 - 0xff -- plane 1
      12'hFA9: dout <= 8'b11111111; // 4009 : 255 - 0xff
      12'hFAA: dout <= 8'b11111111; // 4010 : 255 - 0xff
      12'hFAB: dout <= 8'b11111111; // 4011 : 255 - 0xff
      12'hFAC: dout <= 8'b11111111; // 4012 : 255 - 0xff
      12'hFAD: dout <= 8'b11111111; // 4013 : 255 - 0xff
      12'hFAE: dout <= 8'b11111111; // 4014 : 255 - 0xff
      12'hFAF: dout <= 8'b11111111; // 4015 : 255 - 0xff
      12'hFB0: dout <= 8'b11111111; // 4016 : 255 - 0xff -- Background 0xfb
      12'hFB1: dout <= 8'b00000000; // 4017 :   0 - 0x0
      12'hFB2: dout <= 8'b00000000; // 4018 :   0 - 0x0
      12'hFB3: dout <= 8'b00000000; // 4019 :   0 - 0x0
      12'hFB4: dout <= 8'b00000000; // 4020 :   0 - 0x0
      12'hFB5: dout <= 8'b11111111; // 4021 : 255 - 0xff
      12'hFB6: dout <= 8'b11111111; // 4022 : 255 - 0xff
      12'hFB7: dout <= 8'b11111111; // 4023 : 255 - 0xff
      12'hFB8: dout <= 8'b00000000; // 4024 :   0 - 0x0 -- plane 1
      12'hFB9: dout <= 8'b00000000; // 4025 :   0 - 0x0
      12'hFBA: dout <= 8'b00000000; // 4026 :   0 - 0x0
      12'hFBB: dout <= 8'b00000000; // 4027 :   0 - 0x0
      12'hFBC: dout <= 8'b00000000; // 4028 :   0 - 0x0
      12'hFBD: dout <= 8'b00000000; // 4029 :   0 - 0x0
      12'hFBE: dout <= 8'b00000000; // 4030 :   0 - 0x0
      12'hFBF: dout <= 8'b00000000; // 4031 :   0 - 0x0
      12'hFC0: dout <= 8'b10000111; // 4032 : 135 - 0x87 -- Background 0xfc
      12'hFC1: dout <= 8'b10000111; // 4033 : 135 - 0x87
      12'hFC2: dout <= 8'b10000111; // 4034 : 135 - 0x87
      12'hFC3: dout <= 8'b10000111; // 4035 : 135 - 0x87
      12'hFC4: dout <= 8'b10000111; // 4036 : 135 - 0x87
      12'hFC5: dout <= 8'b10000111; // 4037 : 135 - 0x87
      12'hFC6: dout <= 8'b10000111; // 4038 : 135 - 0x87
      12'hFC7: dout <= 8'b10000111; // 4039 : 135 - 0x87
      12'hFC8: dout <= 8'b00000000; // 4040 :   0 - 0x0 -- plane 1
      12'hFC9: dout <= 8'b00000000; // 4041 :   0 - 0x0
      12'hFCA: dout <= 8'b00000000; // 4042 :   0 - 0x0
      12'hFCB: dout <= 8'b00000000; // 4043 :   0 - 0x0
      12'hFCC: dout <= 8'b00000000; // 4044 :   0 - 0x0
      12'hFCD: dout <= 8'b00000000; // 4045 :   0 - 0x0
      12'hFCE: dout <= 8'b00000000; // 4046 :   0 - 0x0
      12'hFCF: dout <= 8'b00000000; // 4047 :   0 - 0x0
      12'hFD0: dout <= 8'b11111111; // 4048 : 255 - 0xff -- Background 0xfd
      12'hFD1: dout <= 8'b11111111; // 4049 : 255 - 0xff
      12'hFD2: dout <= 8'b11111111; // 4050 : 255 - 0xff
      12'hFD3: dout <= 8'b11000011; // 4051 : 195 - 0xc3
      12'hFD4: dout <= 8'b11000011; // 4052 : 195 - 0xc3
      12'hFD5: dout <= 8'b11111111; // 4053 : 255 - 0xff
      12'hFD6: dout <= 8'b11111111; // 4054 : 255 - 0xff
      12'hFD7: dout <= 8'b11111111; // 4055 : 255 - 0xff
      12'hFD8: dout <= 8'b00000000; // 4056 :   0 - 0x0 -- plane 1
      12'hFD9: dout <= 8'b00000000; // 4057 :   0 - 0x0
      12'hFDA: dout <= 8'b00000000; // 4058 :   0 - 0x0
      12'hFDB: dout <= 8'b00111100; // 4059 :  60 - 0x3c
      12'hFDC: dout <= 8'b00111100; // 4060 :  60 - 0x3c
      12'hFDD: dout <= 8'b00000000; // 4061 :   0 - 0x0
      12'hFDE: dout <= 8'b00000000; // 4062 :   0 - 0x0
      12'hFDF: dout <= 8'b00000000; // 4063 :   0 - 0x0
      12'hFE0: dout <= 8'b11111111; // 4064 : 255 - 0xff -- Background 0xfe
      12'hFE1: dout <= 8'b11111111; // 4065 : 255 - 0xff
      12'hFE2: dout <= 8'b11100111; // 4066 : 231 - 0xe7
      12'hFE3: dout <= 8'b11100111; // 4067 : 231 - 0xe7
      12'hFE4: dout <= 8'b11100111; // 4068 : 231 - 0xe7
      12'hFE5: dout <= 8'b11100111; // 4069 : 231 - 0xe7
      12'hFE6: dout <= 8'b11111111; // 4070 : 255 - 0xff
      12'hFE7: dout <= 8'b11111111; // 4071 : 255 - 0xff
      12'hFE8: dout <= 8'b00000000; // 4072 :   0 - 0x0 -- plane 1
      12'hFE9: dout <= 8'b00000000; // 4073 :   0 - 0x0
      12'hFEA: dout <= 8'b00011000; // 4074 :  24 - 0x18
      12'hFEB: dout <= 8'b00011000; // 4075 :  24 - 0x18
      12'hFEC: dout <= 8'b00011000; // 4076 :  24 - 0x18
      12'hFED: dout <= 8'b00011000; // 4077 :  24 - 0x18
      12'hFEE: dout <= 8'b00000000; // 4078 :   0 - 0x0
      12'hFEF: dout <= 8'b00000000; // 4079 :   0 - 0x0
      12'hFF0: dout <= 8'b11111111; // 4080 : 255 - 0xff -- Background 0xff
      12'hFF1: dout <= 8'b11111111; // 4081 : 255 - 0xff
      12'hFF2: dout <= 8'b11111111; // 4082 : 255 - 0xff
      12'hFF3: dout <= 8'b11111111; // 4083 : 255 - 0xff
      12'hFF4: dout <= 8'b11111111; // 4084 : 255 - 0xff
      12'hFF5: dout <= 8'b11111111; // 4085 : 255 - 0xff
      12'hFF6: dout <= 8'b11111111; // 4086 : 255 - 0xff
      12'hFF7: dout <= 8'b11111111; // 4087 : 255 - 0xff
      12'hFF8: dout <= 8'b00000000; // 4088 :   0 - 0x0 -- plane 1
      12'hFF9: dout <= 8'b00000000; // 4089 :   0 - 0x0
      12'hFFA: dout <= 8'b00000000; // 4090 :   0 - 0x0
      12'hFFB: dout <= 8'b00000000; // 4091 :   0 - 0x0
      12'hFFC: dout <= 8'b00000000; // 4092 :   0 - 0x0
      12'hFFD: dout <= 8'b00000000; // 4093 :   0 - 0x0
      12'hFFE: dout <= 8'b00000000; // 4094 :   0 - 0x0
      12'hFFF: dout <= 8'b00000000; // 4095 :   0 - 0x0
    endcase
  end

endmodule
