//- Autcmatically generated verilog ROM from a NES memory file----
//-   PATTERN TABLE
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


//-  Original memory dump file name: pacman_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_PTABLE_PACMAN
  (
     input     clk,   // clock
     input      [13-1:0] addr,  //8192 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Pattern Table 0---------
      13'h0: dout <= 8'b00000000; //    0 :   0 - 0x0 -- Sprite 0x0
      13'h1: dout <= 8'b00000000; //    1 :   0 - 0x0
      13'h2: dout <= 8'b00000000; //    2 :   0 - 0x0
      13'h3: dout <= 8'b00000000; //    3 :   0 - 0x0
      13'h4: dout <= 8'b00000000; //    4 :   0 - 0x0
      13'h5: dout <= 8'b00000000; //    5 :   0 - 0x0
      13'h6: dout <= 8'b00000000; //    6 :   0 - 0x0
      13'h7: dout <= 8'b00000000; //    7 :   0 - 0x0
      13'h8: dout <= 8'b00000000; //    8 :   0 - 0x0
      13'h9: dout <= 8'b00000000; //    9 :   0 - 0x0
      13'hA: dout <= 8'b00000000; //   10 :   0 - 0x0
      13'hB: dout <= 8'b00000000; //   11 :   0 - 0x0
      13'hC: dout <= 8'b00000000; //   12 :   0 - 0x0
      13'hD: dout <= 8'b00000000; //   13 :   0 - 0x0
      13'hE: dout <= 8'b00000000; //   14 :   0 - 0x0
      13'hF: dout <= 8'b00000000; //   15 :   0 - 0x0
      13'h10: dout <= 8'b00000000; //   16 :   0 - 0x0 -- Sprite 0x1
      13'h11: dout <= 8'b00111000; //   17 :  56 - 0x38
      13'h12: dout <= 8'b01111100; //   18 : 124 - 0x7c
      13'h13: dout <= 8'b11111110; //   19 : 254 - 0xfe
      13'h14: dout <= 8'b11111110; //   20 : 254 - 0xfe
      13'h15: dout <= 8'b11111110; //   21 : 254 - 0xfe
      13'h16: dout <= 8'b01111100; //   22 : 124 - 0x7c
      13'h17: dout <= 8'b00111000; //   23 :  56 - 0x38
      13'h18: dout <= 8'b00000000; //   24 :   0 - 0x0
      13'h19: dout <= 8'b00111000; //   25 :  56 - 0x38
      13'h1A: dout <= 8'b01111100; //   26 : 124 - 0x7c
      13'h1B: dout <= 8'b11111110; //   27 : 254 - 0xfe
      13'h1C: dout <= 8'b11111110; //   28 : 254 - 0xfe
      13'h1D: dout <= 8'b11111110; //   29 : 254 - 0xfe
      13'h1E: dout <= 8'b01111100; //   30 : 124 - 0x7c
      13'h1F: dout <= 8'b00111000; //   31 :  56 - 0x38
      13'h20: dout <= 8'b00000000; //   32 :   0 - 0x0 -- Sprite 0x2
      13'h21: dout <= 8'b00000000; //   33 :   0 - 0x0
      13'h22: dout <= 8'b00000000; //   34 :   0 - 0x0
      13'h23: dout <= 8'b00000000; //   35 :   0 - 0x0
      13'h24: dout <= 8'b00000000; //   36 :   0 - 0x0
      13'h25: dout <= 8'b00000000; //   37 :   0 - 0x0
      13'h26: dout <= 8'b00000000; //   38 :   0 - 0x0
      13'h27: dout <= 8'b00000000; //   39 :   0 - 0x0
      13'h28: dout <= 8'b00000000; //   40 :   0 - 0x0
      13'h29: dout <= 8'b00000000; //   41 :   0 - 0x0
      13'h2A: dout <= 8'b00000000; //   42 :   0 - 0x0
      13'h2B: dout <= 8'b00000000; //   43 :   0 - 0x0
      13'h2C: dout <= 8'b00000000; //   44 :   0 - 0x0
      13'h2D: dout <= 8'b00000000; //   45 :   0 - 0x0
      13'h2E: dout <= 8'b00000000; //   46 :   0 - 0x0
      13'h2F: dout <= 8'b00000000; //   47 :   0 - 0x0
      13'h30: dout <= 8'b00000000; //   48 :   0 - 0x0 -- Sprite 0x3
      13'h31: dout <= 8'b00000000; //   49 :   0 - 0x0
      13'h32: dout <= 8'b00000000; //   50 :   0 - 0x0
      13'h33: dout <= 8'b00011000; //   51 :  24 - 0x18
      13'h34: dout <= 8'b00011000; //   52 :  24 - 0x18
      13'h35: dout <= 8'b00000000; //   53 :   0 - 0x0
      13'h36: dout <= 8'b00000000; //   54 :   0 - 0x0
      13'h37: dout <= 8'b00000000; //   55 :   0 - 0x0
      13'h38: dout <= 8'b00000000; //   56 :   0 - 0x0
      13'h39: dout <= 8'b00000000; //   57 :   0 - 0x0
      13'h3A: dout <= 8'b00000000; //   58 :   0 - 0x0
      13'h3B: dout <= 8'b00011000; //   59 :  24 - 0x18
      13'h3C: dout <= 8'b00011000; //   60 :  24 - 0x18
      13'h3D: dout <= 8'b00000000; //   61 :   0 - 0x0
      13'h3E: dout <= 8'b00000000; //   62 :   0 - 0x0
      13'h3F: dout <= 8'b00000000; //   63 :   0 - 0x0
      13'h40: dout <= 8'b00000000; //   64 :   0 - 0x0 -- Sprite 0x4
      13'h41: dout <= 8'b00000000; //   65 :   0 - 0x0
      13'h42: dout <= 8'b00000000; //   66 :   0 - 0x0
      13'h43: dout <= 8'b00000000; //   67 :   0 - 0x0
      13'h44: dout <= 8'b00000000; //   68 :   0 - 0x0
      13'h45: dout <= 8'b00000000; //   69 :   0 - 0x0
      13'h46: dout <= 8'b00000000; //   70 :   0 - 0x0
      13'h47: dout <= 8'b00000000; //   71 :   0 - 0x0
      13'h48: dout <= 8'b11111111; //   72 : 255 - 0xff
      13'h49: dout <= 8'b11111111; //   73 : 255 - 0xff
      13'h4A: dout <= 8'b11111111; //   74 : 255 - 0xff
      13'h4B: dout <= 8'b11111111; //   75 : 255 - 0xff
      13'h4C: dout <= 8'b11111111; //   76 : 255 - 0xff
      13'h4D: dout <= 8'b11111111; //   77 : 255 - 0xff
      13'h4E: dout <= 8'b11111111; //   78 : 255 - 0xff
      13'h4F: dout <= 8'b11111111; //   79 : 255 - 0xff
      13'h50: dout <= 8'b00000000; //   80 :   0 - 0x0 -- Sprite 0x5
      13'h51: dout <= 8'b00000000; //   81 :   0 - 0x0
      13'h52: dout <= 8'b00000000; //   82 :   0 - 0x0
      13'h53: dout <= 8'b00000000; //   83 :   0 - 0x0
      13'h54: dout <= 8'b00000000; //   84 :   0 - 0x0
      13'h55: dout <= 8'b00000000; //   85 :   0 - 0x0
      13'h56: dout <= 8'b00000000; //   86 :   0 - 0x0
      13'h57: dout <= 8'b00000000; //   87 :   0 - 0x0
      13'h58: dout <= 8'b00001111; //   88 :  15 - 0xf
      13'h59: dout <= 8'b00001111; //   89 :  15 - 0xf
      13'h5A: dout <= 8'b00001111; //   90 :  15 - 0xf
      13'h5B: dout <= 8'b00001111; //   91 :  15 - 0xf
      13'h5C: dout <= 8'b00001111; //   92 :  15 - 0xf
      13'h5D: dout <= 8'b00001111; //   93 :  15 - 0xf
      13'h5E: dout <= 8'b00001111; //   94 :  15 - 0xf
      13'h5F: dout <= 8'b00001111; //   95 :  15 - 0xf
      13'h60: dout <= 8'b00000000; //   96 :   0 - 0x0 -- Sprite 0x6
      13'h61: dout <= 8'b00000000; //   97 :   0 - 0x0
      13'h62: dout <= 8'b00000000; //   98 :   0 - 0x0
      13'h63: dout <= 8'b00000000; //   99 :   0 - 0x0
      13'h64: dout <= 8'b00000000; //  100 :   0 - 0x0
      13'h65: dout <= 8'b00000000; //  101 :   0 - 0x0
      13'h66: dout <= 8'b00000000; //  102 :   0 - 0x0
      13'h67: dout <= 8'b00000000; //  103 :   0 - 0x0
      13'h68: dout <= 8'b11110000; //  104 : 240 - 0xf0
      13'h69: dout <= 8'b11110000; //  105 : 240 - 0xf0
      13'h6A: dout <= 8'b11110000; //  106 : 240 - 0xf0
      13'h6B: dout <= 8'b11110000; //  107 : 240 - 0xf0
      13'h6C: dout <= 8'b11110000; //  108 : 240 - 0xf0
      13'h6D: dout <= 8'b11110000; //  109 : 240 - 0xf0
      13'h6E: dout <= 8'b11110000; //  110 : 240 - 0xf0
      13'h6F: dout <= 8'b11110000; //  111 : 240 - 0xf0
      13'h70: dout <= 8'b00000000; //  112 :   0 - 0x0 -- Sprite 0x7
      13'h71: dout <= 8'b00000000; //  113 :   0 - 0x0
      13'h72: dout <= 8'b00000000; //  114 :   0 - 0x0
      13'h73: dout <= 8'b00000000; //  115 :   0 - 0x0
      13'h74: dout <= 8'b00000000; //  116 :   0 - 0x0
      13'h75: dout <= 8'b00000000; //  117 :   0 - 0x0
      13'h76: dout <= 8'b00000000; //  118 :   0 - 0x0
      13'h77: dout <= 8'b00000000; //  119 :   0 - 0x0
      13'h78: dout <= 8'b00000000; //  120 :   0 - 0x0
      13'h79: dout <= 8'b00000000; //  121 :   0 - 0x0
      13'h7A: dout <= 8'b00000000; //  122 :   0 - 0x0
      13'h7B: dout <= 8'b00000000; //  123 :   0 - 0x0
      13'h7C: dout <= 8'b00000000; //  124 :   0 - 0x0
      13'h7D: dout <= 8'b00000000; //  125 :   0 - 0x0
      13'h7E: dout <= 8'b00000000; //  126 :   0 - 0x0
      13'h7F: dout <= 8'b00000000; //  127 :   0 - 0x0
      13'h80: dout <= 8'b00000000; //  128 :   0 - 0x0 -- Sprite 0x8
      13'h81: dout <= 8'b00000000; //  129 :   0 - 0x0
      13'h82: dout <= 8'b00000000; //  130 :   0 - 0x0
      13'h83: dout <= 8'b00000000; //  131 :   0 - 0x0
      13'h84: dout <= 8'b00000000; //  132 :   0 - 0x0
      13'h85: dout <= 8'b00000000; //  133 :   0 - 0x0
      13'h86: dout <= 8'b00000000; //  134 :   0 - 0x0
      13'h87: dout <= 8'b00000000; //  135 :   0 - 0x0
      13'h88: dout <= 8'b00000000; //  136 :   0 - 0x0
      13'h89: dout <= 8'b00000000; //  137 :   0 - 0x0
      13'h8A: dout <= 8'b00000000; //  138 :   0 - 0x0
      13'h8B: dout <= 8'b00000000; //  139 :   0 - 0x0
      13'h8C: dout <= 8'b00000000; //  140 :   0 - 0x0
      13'h8D: dout <= 8'b00000000; //  141 :   0 - 0x0
      13'h8E: dout <= 8'b00000000; //  142 :   0 - 0x0
      13'h8F: dout <= 8'b00000000; //  143 :   0 - 0x0
      13'h90: dout <= 8'b00000000; //  144 :   0 - 0x0 -- Sprite 0x9
      13'h91: dout <= 8'b00000000; //  145 :   0 - 0x0
      13'h92: dout <= 8'b00000000; //  146 :   0 - 0x0
      13'h93: dout <= 8'b00011000; //  147 :  24 - 0x18
      13'h94: dout <= 8'b00011000; //  148 :  24 - 0x18
      13'h95: dout <= 8'b00000000; //  149 :   0 - 0x0
      13'h96: dout <= 8'b00000000; //  150 :   0 - 0x0
      13'h97: dout <= 8'b00000000; //  151 :   0 - 0x0
      13'h98: dout <= 8'b00000000; //  152 :   0 - 0x0
      13'h99: dout <= 8'b00000000; //  153 :   0 - 0x0
      13'h9A: dout <= 8'b00000000; //  154 :   0 - 0x0
      13'h9B: dout <= 8'b00011000; //  155 :  24 - 0x18
      13'h9C: dout <= 8'b00011000; //  156 :  24 - 0x18
      13'h9D: dout <= 8'b00000000; //  157 :   0 - 0x0
      13'h9E: dout <= 8'b00000000; //  158 :   0 - 0x0
      13'h9F: dout <= 8'b00000000; //  159 :   0 - 0x0
      13'hA0: dout <= 8'b00000000; //  160 :   0 - 0x0 -- Sprite 0xa
      13'hA1: dout <= 8'b00000000; //  161 :   0 - 0x0
      13'hA2: dout <= 8'b00000000; //  162 :   0 - 0x0
      13'hA3: dout <= 8'b00000000; //  163 :   0 - 0x0
      13'hA4: dout <= 8'b00000000; //  164 :   0 - 0x0
      13'hA5: dout <= 8'b00000000; //  165 :   0 - 0x0
      13'hA6: dout <= 8'b00000000; //  166 :   0 - 0x0
      13'hA7: dout <= 8'b00000000; //  167 :   0 - 0x0
      13'hA8: dout <= 8'b00000000; //  168 :   0 - 0x0
      13'hA9: dout <= 8'b00000000; //  169 :   0 - 0x0
      13'hAA: dout <= 8'b00000000; //  170 :   0 - 0x0
      13'hAB: dout <= 8'b00000000; //  171 :   0 - 0x0
      13'hAC: dout <= 8'b00000000; //  172 :   0 - 0x0
      13'hAD: dout <= 8'b00000000; //  173 :   0 - 0x0
      13'hAE: dout <= 8'b00000000; //  174 :   0 - 0x0
      13'hAF: dout <= 8'b00000000; //  175 :   0 - 0x0
      13'hB0: dout <= 8'b00000000; //  176 :   0 - 0x0 -- Sprite 0xb
      13'hB1: dout <= 8'b00000000; //  177 :   0 - 0x0
      13'hB2: dout <= 8'b00000000; //  178 :   0 - 0x0
      13'hB3: dout <= 8'b00000000; //  179 :   0 - 0x0
      13'hB4: dout <= 8'b00000000; //  180 :   0 - 0x0
      13'hB5: dout <= 8'b00000000; //  181 :   0 - 0x0
      13'hB6: dout <= 8'b00000000; //  182 :   0 - 0x0
      13'hB7: dout <= 8'b00000000; //  183 :   0 - 0x0
      13'hB8: dout <= 8'b00000000; //  184 :   0 - 0x0
      13'hB9: dout <= 8'b00000000; //  185 :   0 - 0x0
      13'hBA: dout <= 8'b00000000; //  186 :   0 - 0x0
      13'hBB: dout <= 8'b00000000; //  187 :   0 - 0x0
      13'hBC: dout <= 8'b00000000; //  188 :   0 - 0x0
      13'hBD: dout <= 8'b00000000; //  189 :   0 - 0x0
      13'hBE: dout <= 8'b00000000; //  190 :   0 - 0x0
      13'hBF: dout <= 8'b00000000; //  191 :   0 - 0x0
      13'hC0: dout <= 8'b00000000; //  192 :   0 - 0x0 -- Sprite 0xc
      13'hC1: dout <= 8'b00000000; //  193 :   0 - 0x0
      13'hC2: dout <= 8'b00000000; //  194 :   0 - 0x0
      13'hC3: dout <= 8'b00000000; //  195 :   0 - 0x0
      13'hC4: dout <= 8'b00000000; //  196 :   0 - 0x0
      13'hC5: dout <= 8'b00000000; //  197 :   0 - 0x0
      13'hC6: dout <= 8'b00000000; //  198 :   0 - 0x0
      13'hC7: dout <= 8'b00000000; //  199 :   0 - 0x0
      13'hC8: dout <= 8'b00000000; //  200 :   0 - 0x0
      13'hC9: dout <= 8'b00000000; //  201 :   0 - 0x0
      13'hCA: dout <= 8'b00000000; //  202 :   0 - 0x0
      13'hCB: dout <= 8'b00000000; //  203 :   0 - 0x0
      13'hCC: dout <= 8'b00000000; //  204 :   0 - 0x0
      13'hCD: dout <= 8'b00000000; //  205 :   0 - 0x0
      13'hCE: dout <= 8'b00000000; //  206 :   0 - 0x0
      13'hCF: dout <= 8'b00000000; //  207 :   0 - 0x0
      13'hD0: dout <= 8'b00000000; //  208 :   0 - 0x0 -- Sprite 0xd
      13'hD1: dout <= 8'b00000000; //  209 :   0 - 0x0
      13'hD2: dout <= 8'b00000000; //  210 :   0 - 0x0
      13'hD3: dout <= 8'b00000000; //  211 :   0 - 0x0
      13'hD4: dout <= 8'b00000000; //  212 :   0 - 0x0
      13'hD5: dout <= 8'b00000000; //  213 :   0 - 0x0
      13'hD6: dout <= 8'b00000000; //  214 :   0 - 0x0
      13'hD7: dout <= 8'b00000000; //  215 :   0 - 0x0
      13'hD8: dout <= 8'b00000000; //  216 :   0 - 0x0
      13'hD9: dout <= 8'b00000000; //  217 :   0 - 0x0
      13'hDA: dout <= 8'b00000000; //  218 :   0 - 0x0
      13'hDB: dout <= 8'b00000000; //  219 :   0 - 0x0
      13'hDC: dout <= 8'b00000000; //  220 :   0 - 0x0
      13'hDD: dout <= 8'b00000000; //  221 :   0 - 0x0
      13'hDE: dout <= 8'b00000000; //  222 :   0 - 0x0
      13'hDF: dout <= 8'b00000000; //  223 :   0 - 0x0
      13'hE0: dout <= 8'b00000000; //  224 :   0 - 0x0 -- Sprite 0xe
      13'hE1: dout <= 8'b00000000; //  225 :   0 - 0x0
      13'hE2: dout <= 8'b00000000; //  226 :   0 - 0x0
      13'hE3: dout <= 8'b00000000; //  227 :   0 - 0x0
      13'hE4: dout <= 8'b00000000; //  228 :   0 - 0x0
      13'hE5: dout <= 8'b00000000; //  229 :   0 - 0x0
      13'hE6: dout <= 8'b00000000; //  230 :   0 - 0x0
      13'hE7: dout <= 8'b00000000; //  231 :   0 - 0x0
      13'hE8: dout <= 8'b00000000; //  232 :   0 - 0x0
      13'hE9: dout <= 8'b00000000; //  233 :   0 - 0x0
      13'hEA: dout <= 8'b00000000; //  234 :   0 - 0x0
      13'hEB: dout <= 8'b00000000; //  235 :   0 - 0x0
      13'hEC: dout <= 8'b00000000; //  236 :   0 - 0x0
      13'hED: dout <= 8'b00000000; //  237 :   0 - 0x0
      13'hEE: dout <= 8'b00000000; //  238 :   0 - 0x0
      13'hEF: dout <= 8'b00000000; //  239 :   0 - 0x0
      13'hF0: dout <= 8'b00000000; //  240 :   0 - 0x0 -- Sprite 0xf
      13'hF1: dout <= 8'b00000000; //  241 :   0 - 0x0
      13'hF2: dout <= 8'b00000000; //  242 :   0 - 0x0
      13'hF3: dout <= 8'b00000000; //  243 :   0 - 0x0
      13'hF4: dout <= 8'b00000000; //  244 :   0 - 0x0
      13'hF5: dout <= 8'b00000000; //  245 :   0 - 0x0
      13'hF6: dout <= 8'b00000000; //  246 :   0 - 0x0
      13'hF7: dout <= 8'b00000000; //  247 :   0 - 0x0
      13'hF8: dout <= 8'b00000000; //  248 :   0 - 0x0
      13'hF9: dout <= 8'b00000000; //  249 :   0 - 0x0
      13'hFA: dout <= 8'b00000000; //  250 :   0 - 0x0
      13'hFB: dout <= 8'b00000000; //  251 :   0 - 0x0
      13'hFC: dout <= 8'b00000000; //  252 :   0 - 0x0
      13'hFD: dout <= 8'b00000000; //  253 :   0 - 0x0
      13'hFE: dout <= 8'b00000000; //  254 :   0 - 0x0
      13'hFF: dout <= 8'b00000000; //  255 :   0 - 0x0
      13'h100: dout <= 8'b00000000; //  256 :   0 - 0x0 -- Sprite 0x10
      13'h101: dout <= 8'b00000000; //  257 :   0 - 0x0
      13'h102: dout <= 8'b11111111; //  258 : 255 - 0xff
      13'h103: dout <= 8'b00000000; //  259 :   0 - 0x0
      13'h104: dout <= 8'b00000000; //  260 :   0 - 0x0
      13'h105: dout <= 8'b11111111; //  261 : 255 - 0xff
      13'h106: dout <= 8'b00000000; //  262 :   0 - 0x0
      13'h107: dout <= 8'b00000000; //  263 :   0 - 0x0
      13'h108: dout <= 8'b00000000; //  264 :   0 - 0x0
      13'h109: dout <= 8'b00000000; //  265 :   0 - 0x0
      13'h10A: dout <= 8'b00000000; //  266 :   0 - 0x0
      13'h10B: dout <= 8'b00000000; //  267 :   0 - 0x0
      13'h10C: dout <= 8'b00000000; //  268 :   0 - 0x0
      13'h10D: dout <= 8'b00000000; //  269 :   0 - 0x0
      13'h10E: dout <= 8'b00000000; //  270 :   0 - 0x0
      13'h10F: dout <= 8'b00000000; //  271 :   0 - 0x0
      13'h110: dout <= 8'b00100100; //  272 :  36 - 0x24 -- Sprite 0x11
      13'h111: dout <= 8'b00100100; //  273 :  36 - 0x24
      13'h112: dout <= 8'b00100100; //  274 :  36 - 0x24
      13'h113: dout <= 8'b00100100; //  275 :  36 - 0x24
      13'h114: dout <= 8'b00100100; //  276 :  36 - 0x24
      13'h115: dout <= 8'b00100100; //  277 :  36 - 0x24
      13'h116: dout <= 8'b00100100; //  278 :  36 - 0x24
      13'h117: dout <= 8'b00100100; //  279 :  36 - 0x24
      13'h118: dout <= 8'b00000000; //  280 :   0 - 0x0
      13'h119: dout <= 8'b00000000; //  281 :   0 - 0x0
      13'h11A: dout <= 8'b00000000; //  282 :   0 - 0x0
      13'h11B: dout <= 8'b00000000; //  283 :   0 - 0x0
      13'h11C: dout <= 8'b00000000; //  284 :   0 - 0x0
      13'h11D: dout <= 8'b00000000; //  285 :   0 - 0x0
      13'h11E: dout <= 8'b00000000; //  286 :   0 - 0x0
      13'h11F: dout <= 8'b00000000; //  287 :   0 - 0x0
      13'h120: dout <= 8'b00100100; //  288 :  36 - 0x24 -- Sprite 0x12
      13'h121: dout <= 8'b00100100; //  289 :  36 - 0x24
      13'h122: dout <= 8'b11000011; //  290 : 195 - 0xc3
      13'h123: dout <= 8'b00000000; //  291 :   0 - 0x0
      13'h124: dout <= 8'b00000000; //  292 :   0 - 0x0
      13'h125: dout <= 8'b11111111; //  293 : 255 - 0xff
      13'h126: dout <= 8'b00000000; //  294 :   0 - 0x0
      13'h127: dout <= 8'b00000000; //  295 :   0 - 0x0
      13'h128: dout <= 8'b00000000; //  296 :   0 - 0x0
      13'h129: dout <= 8'b00000000; //  297 :   0 - 0x0
      13'h12A: dout <= 8'b00000000; //  298 :   0 - 0x0
      13'h12B: dout <= 8'b00000000; //  299 :   0 - 0x0
      13'h12C: dout <= 8'b00000000; //  300 :   0 - 0x0
      13'h12D: dout <= 8'b00000000; //  301 :   0 - 0x0
      13'h12E: dout <= 8'b00000000; //  302 :   0 - 0x0
      13'h12F: dout <= 8'b00000000; //  303 :   0 - 0x0
      13'h130: dout <= 8'b00000000; //  304 :   0 - 0x0 -- Sprite 0x13
      13'h131: dout <= 8'b00000000; //  305 :   0 - 0x0
      13'h132: dout <= 8'b11111111; //  306 : 255 - 0xff
      13'h133: dout <= 8'b00000000; //  307 :   0 - 0x0
      13'h134: dout <= 8'b00000000; //  308 :   0 - 0x0
      13'h135: dout <= 8'b11000011; //  309 : 195 - 0xc3
      13'h136: dout <= 8'b00100100; //  310 :  36 - 0x24
      13'h137: dout <= 8'b00100100; //  311 :  36 - 0x24
      13'h138: dout <= 8'b00000000; //  312 :   0 - 0x0
      13'h139: dout <= 8'b00000000; //  313 :   0 - 0x0
      13'h13A: dout <= 8'b00000000; //  314 :   0 - 0x0
      13'h13B: dout <= 8'b00000000; //  315 :   0 - 0x0
      13'h13C: dout <= 8'b00000000; //  316 :   0 - 0x0
      13'h13D: dout <= 8'b00000000; //  317 :   0 - 0x0
      13'h13E: dout <= 8'b00000000; //  318 :   0 - 0x0
      13'h13F: dout <= 8'b00000000; //  319 :   0 - 0x0
      13'h140: dout <= 8'b00100100; //  320 :  36 - 0x24 -- Sprite 0x14
      13'h141: dout <= 8'b00100100; //  321 :  36 - 0x24
      13'h142: dout <= 8'b11000100; //  322 : 196 - 0xc4
      13'h143: dout <= 8'b00000100; //  323 :   4 - 0x4
      13'h144: dout <= 8'b00000100; //  324 :   4 - 0x4
      13'h145: dout <= 8'b11000100; //  325 : 196 - 0xc4
      13'h146: dout <= 8'b00100100; //  326 :  36 - 0x24
      13'h147: dout <= 8'b00100100; //  327 :  36 - 0x24
      13'h148: dout <= 8'b00000000; //  328 :   0 - 0x0
      13'h149: dout <= 8'b00000000; //  329 :   0 - 0x0
      13'h14A: dout <= 8'b00000000; //  330 :   0 - 0x0
      13'h14B: dout <= 8'b00000000; //  331 :   0 - 0x0
      13'h14C: dout <= 8'b00000000; //  332 :   0 - 0x0
      13'h14D: dout <= 8'b00000000; //  333 :   0 - 0x0
      13'h14E: dout <= 8'b00000000; //  334 :   0 - 0x0
      13'h14F: dout <= 8'b00000000; //  335 :   0 - 0x0
      13'h150: dout <= 8'b00100100; //  336 :  36 - 0x24 -- Sprite 0x15
      13'h151: dout <= 8'b00100100; //  337 :  36 - 0x24
      13'h152: dout <= 8'b00100011; //  338 :  35 - 0x23
      13'h153: dout <= 8'b00100000; //  339 :  32 - 0x20
      13'h154: dout <= 8'b00100000; //  340 :  32 - 0x20
      13'h155: dout <= 8'b00100011; //  341 :  35 - 0x23
      13'h156: dout <= 8'b00100100; //  342 :  36 - 0x24
      13'h157: dout <= 8'b00100100; //  343 :  36 - 0x24
      13'h158: dout <= 8'b00000000; //  344 :   0 - 0x0
      13'h159: dout <= 8'b00000000; //  345 :   0 - 0x0
      13'h15A: dout <= 8'b00000000; //  346 :   0 - 0x0
      13'h15B: dout <= 8'b00000000; //  347 :   0 - 0x0
      13'h15C: dout <= 8'b00000000; //  348 :   0 - 0x0
      13'h15D: dout <= 8'b00000000; //  349 :   0 - 0x0
      13'h15E: dout <= 8'b00000000; //  350 :   0 - 0x0
      13'h15F: dout <= 8'b00000000; //  351 :   0 - 0x0
      13'h160: dout <= 8'b00000000; //  352 :   0 - 0x0 -- Sprite 0x16
      13'h161: dout <= 8'b00000000; //  353 :   0 - 0x0
      13'h162: dout <= 8'b00001111; //  354 :  15 - 0xf
      13'h163: dout <= 8'b00010000; //  355 :  16 - 0x10
      13'h164: dout <= 8'b11110000; //  356 : 240 - 0xf0
      13'h165: dout <= 8'b00001111; //  357 :  15 - 0xf
      13'h166: dout <= 8'b00000000; //  358 :   0 - 0x0
      13'h167: dout <= 8'b00000000; //  359 :   0 - 0x0
      13'h168: dout <= 8'b00000000; //  360 :   0 - 0x0
      13'h169: dout <= 8'b00000000; //  361 :   0 - 0x0
      13'h16A: dout <= 8'b00000000; //  362 :   0 - 0x0
      13'h16B: dout <= 8'b00000000; //  363 :   0 - 0x0
      13'h16C: dout <= 8'b00000000; //  364 :   0 - 0x0
      13'h16D: dout <= 8'b00000000; //  365 :   0 - 0x0
      13'h16E: dout <= 8'b00000000; //  366 :   0 - 0x0
      13'h16F: dout <= 8'b00000000; //  367 :   0 - 0x0
      13'h170: dout <= 8'b00000000; //  368 :   0 - 0x0 -- Sprite 0x17
      13'h171: dout <= 8'b00000000; //  369 :   0 - 0x0
      13'h172: dout <= 8'b11110000; //  370 : 240 - 0xf0
      13'h173: dout <= 8'b00001000; //  371 :   8 - 0x8
      13'h174: dout <= 8'b00001111; //  372 :  15 - 0xf
      13'h175: dout <= 8'b11110000; //  373 : 240 - 0xf0
      13'h176: dout <= 8'b00000000; //  374 :   0 - 0x0
      13'h177: dout <= 8'b00000000; //  375 :   0 - 0x0
      13'h178: dout <= 8'b00000000; //  376 :   0 - 0x0
      13'h179: dout <= 8'b00000000; //  377 :   0 - 0x0
      13'h17A: dout <= 8'b00000000; //  378 :   0 - 0x0
      13'h17B: dout <= 8'b00000000; //  379 :   0 - 0x0
      13'h17C: dout <= 8'b00000000; //  380 :   0 - 0x0
      13'h17D: dout <= 8'b00000000; //  381 :   0 - 0x0
      13'h17E: dout <= 8'b00000000; //  382 :   0 - 0x0
      13'h17F: dout <= 8'b00000000; //  383 :   0 - 0x0
      13'h180: dout <= 8'b00000000; //  384 :   0 - 0x0 -- Sprite 0x18
      13'h181: dout <= 8'b00000000; //  385 :   0 - 0x0
      13'h182: dout <= 8'b11110000; //  386 : 240 - 0xf0
      13'h183: dout <= 8'b00001000; //  387 :   8 - 0x8
      13'h184: dout <= 8'b00001000; //  388 :   8 - 0x8
      13'h185: dout <= 8'b11110000; //  389 : 240 - 0xf0
      13'h186: dout <= 8'b00000000; //  390 :   0 - 0x0
      13'h187: dout <= 8'b00000000; //  391 :   0 - 0x0
      13'h188: dout <= 8'b00000000; //  392 :   0 - 0x0
      13'h189: dout <= 8'b00000000; //  393 :   0 - 0x0
      13'h18A: dout <= 8'b00000000; //  394 :   0 - 0x0
      13'h18B: dout <= 8'b00000000; //  395 :   0 - 0x0
      13'h18C: dout <= 8'b00000000; //  396 :   0 - 0x0
      13'h18D: dout <= 8'b00000000; //  397 :   0 - 0x0
      13'h18E: dout <= 8'b00000000; //  398 :   0 - 0x0
      13'h18F: dout <= 8'b00000000; //  399 :   0 - 0x0
      13'h190: dout <= 8'b00000000; //  400 :   0 - 0x0 -- Sprite 0x19
      13'h191: dout <= 8'b00000000; //  401 :   0 - 0x0
      13'h192: dout <= 8'b00001111; //  402 :  15 - 0xf
      13'h193: dout <= 8'b00010000; //  403 :  16 - 0x10
      13'h194: dout <= 8'b00010000; //  404 :  16 - 0x10
      13'h195: dout <= 8'b00001111; //  405 :  15 - 0xf
      13'h196: dout <= 8'b00000000; //  406 :   0 - 0x0
      13'h197: dout <= 8'b00000000; //  407 :   0 - 0x0
      13'h198: dout <= 8'b00000000; //  408 :   0 - 0x0
      13'h199: dout <= 8'b00000000; //  409 :   0 - 0x0
      13'h19A: dout <= 8'b00000000; //  410 :   0 - 0x0
      13'h19B: dout <= 8'b00000000; //  411 :   0 - 0x0
      13'h19C: dout <= 8'b00000000; //  412 :   0 - 0x0
      13'h19D: dout <= 8'b00000000; //  413 :   0 - 0x0
      13'h19E: dout <= 8'b00000000; //  414 :   0 - 0x0
      13'h19F: dout <= 8'b00000000; //  415 :   0 - 0x0
      13'h1A0: dout <= 8'b00100100; //  416 :  36 - 0x24 -- Sprite 0x1a
      13'h1A1: dout <= 8'b00100100; //  417 :  36 - 0x24
      13'h1A2: dout <= 8'b00100100; //  418 :  36 - 0x24
      13'h1A3: dout <= 8'b00100100; //  419 :  36 - 0x24
      13'h1A4: dout <= 8'b00011000; //  420 :  24 - 0x18
      13'h1A5: dout <= 8'b00000000; //  421 :   0 - 0x0
      13'h1A6: dout <= 8'b00000000; //  422 :   0 - 0x0
      13'h1A7: dout <= 8'b00000000; //  423 :   0 - 0x0
      13'h1A8: dout <= 8'b00000000; //  424 :   0 - 0x0
      13'h1A9: dout <= 8'b00000000; //  425 :   0 - 0x0
      13'h1AA: dout <= 8'b00000000; //  426 :   0 - 0x0
      13'h1AB: dout <= 8'b00000000; //  427 :   0 - 0x0
      13'h1AC: dout <= 8'b00000000; //  428 :   0 - 0x0
      13'h1AD: dout <= 8'b00000000; //  429 :   0 - 0x0
      13'h1AE: dout <= 8'b00000000; //  430 :   0 - 0x0
      13'h1AF: dout <= 8'b00000000; //  431 :   0 - 0x0
      13'h1B0: dout <= 8'b00000000; //  432 :   0 - 0x0 -- Sprite 0x1b
      13'h1B1: dout <= 8'b00000000; //  433 :   0 - 0x0
      13'h1B2: dout <= 8'b00000000; //  434 :   0 - 0x0
      13'h1B3: dout <= 8'b00011000; //  435 :  24 - 0x18
      13'h1B4: dout <= 8'b00100100; //  436 :  36 - 0x24
      13'h1B5: dout <= 8'b00100100; //  437 :  36 - 0x24
      13'h1B6: dout <= 8'b00100100; //  438 :  36 - 0x24
      13'h1B7: dout <= 8'b00100100; //  439 :  36 - 0x24
      13'h1B8: dout <= 8'b00000000; //  440 :   0 - 0x0
      13'h1B9: dout <= 8'b00000000; //  441 :   0 - 0x0
      13'h1BA: dout <= 8'b00000000; //  442 :   0 - 0x0
      13'h1BB: dout <= 8'b00000000; //  443 :   0 - 0x0
      13'h1BC: dout <= 8'b00000000; //  444 :   0 - 0x0
      13'h1BD: dout <= 8'b00000000; //  445 :   0 - 0x0
      13'h1BE: dout <= 8'b00000000; //  446 :   0 - 0x0
      13'h1BF: dout <= 8'b00000000; //  447 :   0 - 0x0
      13'h1C0: dout <= 8'b00100100; //  448 :  36 - 0x24 -- Sprite 0x1c
      13'h1C1: dout <= 8'b00100100; //  449 :  36 - 0x24
      13'h1C2: dout <= 8'b11000100; //  450 : 196 - 0xc4
      13'h1C3: dout <= 8'b00000100; //  451 :   4 - 0x4
      13'h1C4: dout <= 8'b00001000; //  452 :   8 - 0x8
      13'h1C5: dout <= 8'b11110000; //  453 : 240 - 0xf0
      13'h1C6: dout <= 8'b00000000; //  454 :   0 - 0x0
      13'h1C7: dout <= 8'b00000000; //  455 :   0 - 0x0
      13'h1C8: dout <= 8'b00000000; //  456 :   0 - 0x0
      13'h1C9: dout <= 8'b00000000; //  457 :   0 - 0x0
      13'h1CA: dout <= 8'b00000000; //  458 :   0 - 0x0
      13'h1CB: dout <= 8'b00000000; //  459 :   0 - 0x0
      13'h1CC: dout <= 8'b00000000; //  460 :   0 - 0x0
      13'h1CD: dout <= 8'b00000000; //  461 :   0 - 0x0
      13'h1CE: dout <= 8'b00000000; //  462 :   0 - 0x0
      13'h1CF: dout <= 8'b00000000; //  463 :   0 - 0x0
      13'h1D0: dout <= 8'b00000000; //  464 :   0 - 0x0 -- Sprite 0x1d
      13'h1D1: dout <= 8'b00000000; //  465 :   0 - 0x0
      13'h1D2: dout <= 8'b11110000; //  466 : 240 - 0xf0
      13'h1D3: dout <= 8'b00001000; //  467 :   8 - 0x8
      13'h1D4: dout <= 8'b00000100; //  468 :   4 - 0x4
      13'h1D5: dout <= 8'b11000100; //  469 : 196 - 0xc4
      13'h1D6: dout <= 8'b00100100; //  470 :  36 - 0x24
      13'h1D7: dout <= 8'b00100100; //  471 :  36 - 0x24
      13'h1D8: dout <= 8'b00000000; //  472 :   0 - 0x0
      13'h1D9: dout <= 8'b00000000; //  473 :   0 - 0x0
      13'h1DA: dout <= 8'b00000000; //  474 :   0 - 0x0
      13'h1DB: dout <= 8'b00000000; //  475 :   0 - 0x0
      13'h1DC: dout <= 8'b00000000; //  476 :   0 - 0x0
      13'h1DD: dout <= 8'b00000000; //  477 :   0 - 0x0
      13'h1DE: dout <= 8'b00000000; //  478 :   0 - 0x0
      13'h1DF: dout <= 8'b00000000; //  479 :   0 - 0x0
      13'h1E0: dout <= 8'b00100100; //  480 :  36 - 0x24 -- Sprite 0x1e
      13'h1E1: dout <= 8'b00100100; //  481 :  36 - 0x24
      13'h1E2: dout <= 8'b00100011; //  482 :  35 - 0x23
      13'h1E3: dout <= 8'b00100000; //  483 :  32 - 0x20
      13'h1E4: dout <= 8'b00010000; //  484 :  16 - 0x10
      13'h1E5: dout <= 8'b00001111; //  485 :  15 - 0xf
      13'h1E6: dout <= 8'b00000000; //  486 :   0 - 0x0
      13'h1E7: dout <= 8'b00000000; //  487 :   0 - 0x0
      13'h1E8: dout <= 8'b00000000; //  488 :   0 - 0x0
      13'h1E9: dout <= 8'b00000000; //  489 :   0 - 0x0
      13'h1EA: dout <= 8'b00000000; //  490 :   0 - 0x0
      13'h1EB: dout <= 8'b00000000; //  491 :   0 - 0x0
      13'h1EC: dout <= 8'b00000000; //  492 :   0 - 0x0
      13'h1ED: dout <= 8'b00000000; //  493 :   0 - 0x0
      13'h1EE: dout <= 8'b00000000; //  494 :   0 - 0x0
      13'h1EF: dout <= 8'b00000000; //  495 :   0 - 0x0
      13'h1F0: dout <= 8'b00000000; //  496 :   0 - 0x0 -- Sprite 0x1f
      13'h1F1: dout <= 8'b00000000; //  497 :   0 - 0x0
      13'h1F2: dout <= 8'b00001111; //  498 :  15 - 0xf
      13'h1F3: dout <= 8'b00010000; //  499 :  16 - 0x10
      13'h1F4: dout <= 8'b00100000; //  500 :  32 - 0x20
      13'h1F5: dout <= 8'b00100011; //  501 :  35 - 0x23
      13'h1F6: dout <= 8'b00100100; //  502 :  36 - 0x24
      13'h1F7: dout <= 8'b00100100; //  503 :  36 - 0x24
      13'h1F8: dout <= 8'b00000000; //  504 :   0 - 0x0
      13'h1F9: dout <= 8'b00000000; //  505 :   0 - 0x0
      13'h1FA: dout <= 8'b00000000; //  506 :   0 - 0x0
      13'h1FB: dout <= 8'b00000000; //  507 :   0 - 0x0
      13'h1FC: dout <= 8'b00000000; //  508 :   0 - 0x0
      13'h1FD: dout <= 8'b00000000; //  509 :   0 - 0x0
      13'h1FE: dout <= 8'b00000000; //  510 :   0 - 0x0
      13'h1FF: dout <= 8'b00000000; //  511 :   0 - 0x0
      13'h200: dout <= 8'b00000000; //  512 :   0 - 0x0 -- Sprite 0x20
      13'h201: dout <= 8'b00000000; //  513 :   0 - 0x0
      13'h202: dout <= 8'b00000000; //  514 :   0 - 0x0
      13'h203: dout <= 8'b00000000; //  515 :   0 - 0x0
      13'h204: dout <= 8'b00000000; //  516 :   0 - 0x0
      13'h205: dout <= 8'b00000000; //  517 :   0 - 0x0
      13'h206: dout <= 8'b00000000; //  518 :   0 - 0x0
      13'h207: dout <= 8'b00000000; //  519 :   0 - 0x0
      13'h208: dout <= 8'b00000000; //  520 :   0 - 0x0
      13'h209: dout <= 8'b00000000; //  521 :   0 - 0x0
      13'h20A: dout <= 8'b00000000; //  522 :   0 - 0x0
      13'h20B: dout <= 8'b00000000; //  523 :   0 - 0x0
      13'h20C: dout <= 8'b00000000; //  524 :   0 - 0x0
      13'h20D: dout <= 8'b00000000; //  525 :   0 - 0x0
      13'h20E: dout <= 8'b00000000; //  526 :   0 - 0x0
      13'h20F: dout <= 8'b00000000; //  527 :   0 - 0x0
      13'h210: dout <= 8'b00000000; //  528 :   0 - 0x0 -- Sprite 0x21
      13'h211: dout <= 8'b00000000; //  529 :   0 - 0x0
      13'h212: dout <= 8'b11110000; //  530 : 240 - 0xf0
      13'h213: dout <= 8'b00001000; //  531 :   8 - 0x8
      13'h214: dout <= 8'b00001000; //  532 :   8 - 0x8
      13'h215: dout <= 8'b11110000; //  533 : 240 - 0xf0
      13'h216: dout <= 8'b00000000; //  534 :   0 - 0x0
      13'h217: dout <= 8'b00000000; //  535 :   0 - 0x0
      13'h218: dout <= 8'b00001111; //  536 :  15 - 0xf
      13'h219: dout <= 8'b00001111; //  537 :  15 - 0xf
      13'h21A: dout <= 8'b00001111; //  538 :  15 - 0xf
      13'h21B: dout <= 8'b00000111; //  539 :   7 - 0x7
      13'h21C: dout <= 8'b00000111; //  540 :   7 - 0x7
      13'h21D: dout <= 8'b00001111; //  541 :  15 - 0xf
      13'h21E: dout <= 8'b00001111; //  542 :  15 - 0xf
      13'h21F: dout <= 8'b00001111; //  543 :  15 - 0xf
      13'h220: dout <= 8'b00000000; //  544 :   0 - 0x0 -- Sprite 0x22
      13'h221: dout <= 8'b00000000; //  545 :   0 - 0x0
      13'h222: dout <= 8'b00001111; //  546 :  15 - 0xf
      13'h223: dout <= 8'b00010000; //  547 :  16 - 0x10
      13'h224: dout <= 8'b00010000; //  548 :  16 - 0x10
      13'h225: dout <= 8'b00001111; //  549 :  15 - 0xf
      13'h226: dout <= 8'b00000000; //  550 :   0 - 0x0
      13'h227: dout <= 8'b00000000; //  551 :   0 - 0x0
      13'h228: dout <= 8'b11110000; //  552 : 240 - 0xf0
      13'h229: dout <= 8'b11110000; //  553 : 240 - 0xf0
      13'h22A: dout <= 8'b11110000; //  554 : 240 - 0xf0
      13'h22B: dout <= 8'b11100000; //  555 : 224 - 0xe0
      13'h22C: dout <= 8'b11100000; //  556 : 224 - 0xe0
      13'h22D: dout <= 8'b11110000; //  557 : 240 - 0xf0
      13'h22E: dout <= 8'b11110000; //  558 : 240 - 0xf0
      13'h22F: dout <= 8'b11110000; //  559 : 240 - 0xf0
      13'h230: dout <= 8'b11111111; //  560 : 255 - 0xff -- Sprite 0x23
      13'h231: dout <= 8'b11111111; //  561 : 255 - 0xff
      13'h232: dout <= 8'b11100001; //  562 : 225 - 0xe1
      13'h233: dout <= 8'b11100001; //  563 : 225 - 0xe1
      13'h234: dout <= 8'b11100001; //  564 : 225 - 0xe1
      13'h235: dout <= 8'b11100001; //  565 : 225 - 0xe1
      13'h236: dout <= 8'b11100001; //  566 : 225 - 0xe1
      13'h237: dout <= 8'b11100001; //  567 : 225 - 0xe1
      13'h238: dout <= 8'b11111111; //  568 : 255 - 0xff
      13'h239: dout <= 8'b11111111; //  569 : 255 - 0xff
      13'h23A: dout <= 8'b11100001; //  570 : 225 - 0xe1
      13'h23B: dout <= 8'b11100001; //  571 : 225 - 0xe1
      13'h23C: dout <= 8'b11100001; //  572 : 225 - 0xe1
      13'h23D: dout <= 8'b11100001; //  573 : 225 - 0xe1
      13'h23E: dout <= 8'b11100001; //  574 : 225 - 0xe1
      13'h23F: dout <= 8'b11100001; //  575 : 225 - 0xe1
      13'h240: dout <= 8'b10000111; //  576 : 135 - 0x87 -- Sprite 0x24
      13'h241: dout <= 8'b11000111; //  577 : 199 - 0xc7
      13'h242: dout <= 8'b11000000; //  578 : 192 - 0xc0
      13'h243: dout <= 8'b11000111; //  579 : 199 - 0xc7
      13'h244: dout <= 8'b11001111; //  580 : 207 - 0xcf
      13'h245: dout <= 8'b11001110; //  581 : 206 - 0xce
      13'h246: dout <= 8'b11001111; //  582 : 207 - 0xcf
      13'h247: dout <= 8'b11000111; //  583 : 199 - 0xc7
      13'h248: dout <= 8'b10000111; //  584 : 135 - 0x87
      13'h249: dout <= 8'b11000111; //  585 : 199 - 0xc7
      13'h24A: dout <= 8'b11000000; //  586 : 192 - 0xc0
      13'h24B: dout <= 8'b11000111; //  587 : 199 - 0xc7
      13'h24C: dout <= 8'b11001111; //  588 : 207 - 0xcf
      13'h24D: dout <= 8'b11001110; //  589 : 206 - 0xce
      13'h24E: dout <= 8'b11001111; //  590 : 207 - 0xcf
      13'h24F: dout <= 8'b11000111; //  591 : 199 - 0xc7
      13'h250: dout <= 8'b11111000; //  592 : 248 - 0xf8 -- Sprite 0x25
      13'h251: dout <= 8'b11111100; //  593 : 252 - 0xfc
      13'h252: dout <= 8'b00011100; //  594 :  28 - 0x1c
      13'h253: dout <= 8'b11111100; //  595 : 252 - 0xfc
      13'h254: dout <= 8'b11111100; //  596 : 252 - 0xfc
      13'h255: dout <= 8'b00011100; //  597 :  28 - 0x1c
      13'h256: dout <= 8'b11111100; //  598 : 252 - 0xfc
      13'h257: dout <= 8'b11111100; //  599 : 252 - 0xfc
      13'h258: dout <= 8'b11111000; //  600 : 248 - 0xf8
      13'h259: dout <= 8'b11111100; //  601 : 252 - 0xfc
      13'h25A: dout <= 8'b00011100; //  602 :  28 - 0x1c
      13'h25B: dout <= 8'b11111100; //  603 : 252 - 0xfc
      13'h25C: dout <= 8'b11111100; //  604 : 252 - 0xfc
      13'h25D: dout <= 8'b00011100; //  605 :  28 - 0x1c
      13'h25E: dout <= 8'b11111100; //  606 : 252 - 0xfc
      13'h25F: dout <= 8'b11111100; //  607 : 252 - 0xfc
      13'h260: dout <= 8'b11111111; //  608 : 255 - 0xff -- Sprite 0x26
      13'h261: dout <= 8'b11111111; //  609 : 255 - 0xff
      13'h262: dout <= 8'b11100111; //  610 : 231 - 0xe7
      13'h263: dout <= 8'b11100111; //  611 : 231 - 0xe7
      13'h264: dout <= 8'b11100111; //  612 : 231 - 0xe7
      13'h265: dout <= 8'b11100111; //  613 : 231 - 0xe7
      13'h266: dout <= 8'b11100111; //  614 : 231 - 0xe7
      13'h267: dout <= 8'b11100111; //  615 : 231 - 0xe7
      13'h268: dout <= 8'b11111111; //  616 : 255 - 0xff
      13'h269: dout <= 8'b11111111; //  617 : 255 - 0xff
      13'h26A: dout <= 8'b11100111; //  618 : 231 - 0xe7
      13'h26B: dout <= 8'b11100111; //  619 : 231 - 0xe7
      13'h26C: dout <= 8'b11100111; //  620 : 231 - 0xe7
      13'h26D: dout <= 8'b11100111; //  621 : 231 - 0xe7
      13'h26E: dout <= 8'b11100111; //  622 : 231 - 0xe7
      13'h26F: dout <= 8'b11100111; //  623 : 231 - 0xe7
      13'h270: dout <= 8'b11110000; //  624 : 240 - 0xf0 -- Sprite 0x27
      13'h271: dout <= 8'b11111001; //  625 : 249 - 0xf9
      13'h272: dout <= 8'b00111001; //  626 :  57 - 0x39
      13'h273: dout <= 8'b00111001; //  627 :  57 - 0x39
      13'h274: dout <= 8'b00111001; //  628 :  57 - 0x39
      13'h275: dout <= 8'b00111001; //  629 :  57 - 0x39
      13'h276: dout <= 8'b00111001; //  630 :  57 - 0x39
      13'h277: dout <= 8'b00111000; //  631 :  56 - 0x38
      13'h278: dout <= 8'b11110000; //  632 : 240 - 0xf0
      13'h279: dout <= 8'b11111001; //  633 : 249 - 0xf9
      13'h27A: dout <= 8'b00111001; //  634 :  57 - 0x39
      13'h27B: dout <= 8'b00111001; //  635 :  57 - 0x39
      13'h27C: dout <= 8'b00111001; //  636 :  57 - 0x39
      13'h27D: dout <= 8'b00111001; //  637 :  57 - 0x39
      13'h27E: dout <= 8'b00111001; //  638 :  57 - 0x39
      13'h27F: dout <= 8'b00111000; //  639 :  56 - 0x38
      13'h280: dout <= 8'b11111111; //  640 : 255 - 0xff -- Sprite 0x28
      13'h281: dout <= 8'b11111111; //  641 : 255 - 0xff
      13'h282: dout <= 8'b11000000; //  642 : 192 - 0xc0
      13'h283: dout <= 8'b11000000; //  643 : 192 - 0xc0
      13'h284: dout <= 8'b11000000; //  644 : 192 - 0xc0
      13'h285: dout <= 8'b11000000; //  645 : 192 - 0xc0
      13'h286: dout <= 8'b11111111; //  646 : 255 - 0xff
      13'h287: dout <= 8'b11111111; //  647 : 255 - 0xff
      13'h288: dout <= 8'b11111111; //  648 : 255 - 0xff
      13'h289: dout <= 8'b11111111; //  649 : 255 - 0xff
      13'h28A: dout <= 8'b11000000; //  650 : 192 - 0xc0
      13'h28B: dout <= 8'b11000000; //  651 : 192 - 0xc0
      13'h28C: dout <= 8'b11000000; //  652 : 192 - 0xc0
      13'h28D: dout <= 8'b11000000; //  653 : 192 - 0xc0
      13'h28E: dout <= 8'b11111111; //  654 : 255 - 0xff
      13'h28F: dout <= 8'b11111111; //  655 : 255 - 0xff
      13'h290: dout <= 8'b00011111; //  656 :  31 - 0x1f -- Sprite 0x29
      13'h291: dout <= 8'b00111111; //  657 :  63 - 0x3f
      13'h292: dout <= 8'b00110000; //  658 :  48 - 0x30
      13'h293: dout <= 8'b00110000; //  659 :  48 - 0x30
      13'h294: dout <= 8'b00110000; //  660 :  48 - 0x30
      13'h295: dout <= 8'b00110000; //  661 :  48 - 0x30
      13'h296: dout <= 8'b00111111; //  662 :  63 - 0x3f
      13'h297: dout <= 8'b00011111; //  663 :  31 - 0x1f
      13'h298: dout <= 8'b00011111; //  664 :  31 - 0x1f
      13'h299: dout <= 8'b00111111; //  665 :  63 - 0x3f
      13'h29A: dout <= 8'b00110000; //  666 :  48 - 0x30
      13'h29B: dout <= 8'b00110000; //  667 :  48 - 0x30
      13'h29C: dout <= 8'b00110000; //  668 :  48 - 0x30
      13'h29D: dout <= 8'b00110000; //  669 :  48 - 0x30
      13'h29E: dout <= 8'b00111111; //  670 :  63 - 0x3f
      13'h29F: dout <= 8'b00011111; //  671 :  31 - 0x1f
      13'h2A0: dout <= 8'b11100011; //  672 : 227 - 0xe3 -- Sprite 0x2a
      13'h2A1: dout <= 8'b11110011; //  673 : 243 - 0xf3
      13'h2A2: dout <= 8'b01110000; //  674 : 112 - 0x70
      13'h2A3: dout <= 8'b01110000; //  675 : 112 - 0x70
      13'h2A4: dout <= 8'b01110000; //  676 : 112 - 0x70
      13'h2A5: dout <= 8'b01110000; //  677 : 112 - 0x70
      13'h2A6: dout <= 8'b11110000; //  678 : 240 - 0xf0
      13'h2A7: dout <= 8'b11100000; //  679 : 224 - 0xe0
      13'h2A8: dout <= 8'b11100011; //  680 : 227 - 0xe3
      13'h2A9: dout <= 8'b11110011; //  681 : 243 - 0xf3
      13'h2AA: dout <= 8'b01110000; //  682 : 112 - 0x70
      13'h2AB: dout <= 8'b01110000; //  683 : 112 - 0x70
      13'h2AC: dout <= 8'b01110000; //  684 : 112 - 0x70
      13'h2AD: dout <= 8'b01110000; //  685 : 112 - 0x70
      13'h2AE: dout <= 8'b11110000; //  686 : 240 - 0xf0
      13'h2AF: dout <= 8'b11100000; //  687 : 224 - 0xe0
      13'h2B0: dout <= 8'b11111110; //  688 : 254 - 0xfe -- Sprite 0x2b
      13'h2B1: dout <= 8'b11111110; //  689 : 254 - 0xfe
      13'h2B2: dout <= 8'b01110000; //  690 : 112 - 0x70
      13'h2B3: dout <= 8'b01110000; //  691 : 112 - 0x70
      13'h2B4: dout <= 8'b01110000; //  692 : 112 - 0x70
      13'h2B5: dout <= 8'b01110000; //  693 : 112 - 0x70
      13'h2B6: dout <= 8'b01110000; //  694 : 112 - 0x70
      13'h2B7: dout <= 8'b01110000; //  695 : 112 - 0x70
      13'h2B8: dout <= 8'b11111110; //  696 : 254 - 0xfe
      13'h2B9: dout <= 8'b11111110; //  697 : 254 - 0xfe
      13'h2BA: dout <= 8'b01110000; //  698 : 112 - 0x70
      13'h2BB: dout <= 8'b01110000; //  699 : 112 - 0x70
      13'h2BC: dout <= 8'b01110000; //  700 : 112 - 0x70
      13'h2BD: dout <= 8'b01110000; //  701 : 112 - 0x70
      13'h2BE: dout <= 8'b01110000; //  702 : 112 - 0x70
      13'h2BF: dout <= 8'b01110000; //  703 : 112 - 0x70
      13'h2C0: dout <= 8'b00000000; //  704 :   0 - 0x0 -- Sprite 0x2c
      13'h2C1: dout <= 8'b00000000; //  705 :   0 - 0x0
      13'h2C2: dout <= 8'b00000000; //  706 :   0 - 0x0
      13'h2C3: dout <= 8'b00000000; //  707 :   0 - 0x0
      13'h2C4: dout <= 8'b11111111; //  708 : 255 - 0xff
      13'h2C5: dout <= 8'b00000000; //  709 :   0 - 0x0
      13'h2C6: dout <= 8'b00000000; //  710 :   0 - 0x0
      13'h2C7: dout <= 8'b00000000; //  711 :   0 - 0x0
      13'h2C8: dout <= 8'b00000000; //  712 :   0 - 0x0
      13'h2C9: dout <= 8'b00000000; //  713 :   0 - 0x0
      13'h2CA: dout <= 8'b00000000; //  714 :   0 - 0x0
      13'h2CB: dout <= 8'b00000000; //  715 :   0 - 0x0
      13'h2CC: dout <= 8'b00000000; //  716 :   0 - 0x0
      13'h2CD: dout <= 8'b00000000; //  717 :   0 - 0x0
      13'h2CE: dout <= 8'b00000000; //  718 :   0 - 0x0
      13'h2CF: dout <= 8'b00000000; //  719 :   0 - 0x0
      13'h2D0: dout <= 8'b00000000; //  720 :   0 - 0x0 -- Sprite 0x2d
      13'h2D1: dout <= 8'b00000000; //  721 :   0 - 0x0
      13'h2D2: dout <= 8'b00000000; //  722 :   0 - 0x0
      13'h2D3: dout <= 8'b00000000; //  723 :   0 - 0x0
      13'h2D4: dout <= 8'b00000000; //  724 :   0 - 0x0
      13'h2D5: dout <= 8'b00000000; //  725 :   0 - 0x0
      13'h2D6: dout <= 8'b00000000; //  726 :   0 - 0x0
      13'h2D7: dout <= 8'b00000000; //  727 :   0 - 0x0
      13'h2D8: dout <= 8'b11111111; //  728 : 255 - 0xff
      13'h2D9: dout <= 8'b11111111; //  729 : 255 - 0xff
      13'h2DA: dout <= 8'b11111111; //  730 : 255 - 0xff
      13'h2DB: dout <= 8'b11111111; //  731 : 255 - 0xff
      13'h2DC: dout <= 8'b11111111; //  732 : 255 - 0xff
      13'h2DD: dout <= 8'b11111111; //  733 : 255 - 0xff
      13'h2DE: dout <= 8'b11111111; //  734 : 255 - 0xff
      13'h2DF: dout <= 8'b11111111; //  735 : 255 - 0xff
      13'h2E0: dout <= 8'b00000000; //  736 :   0 - 0x0 -- Sprite 0x2e
      13'h2E1: dout <= 8'b00000000; //  737 :   0 - 0x0
      13'h2E2: dout <= 8'b00000000; //  738 :   0 - 0x0
      13'h2E3: dout <= 8'b00011000; //  739 :  24 - 0x18
      13'h2E4: dout <= 8'b00011000; //  740 :  24 - 0x18
      13'h2E5: dout <= 8'b00000000; //  741 :   0 - 0x0
      13'h2E6: dout <= 8'b00000000; //  742 :   0 - 0x0
      13'h2E7: dout <= 8'b00000000; //  743 :   0 - 0x0
      13'h2E8: dout <= 8'b00000000; //  744 :   0 - 0x0
      13'h2E9: dout <= 8'b00000000; //  745 :   0 - 0x0
      13'h2EA: dout <= 8'b00000000; //  746 :   0 - 0x0
      13'h2EB: dout <= 8'b00000000; //  747 :   0 - 0x0
      13'h2EC: dout <= 8'b00000000; //  748 :   0 - 0x0
      13'h2ED: dout <= 8'b00000000; //  749 :   0 - 0x0
      13'h2EE: dout <= 8'b00000000; //  750 :   0 - 0x0
      13'h2EF: dout <= 8'b00000000; //  751 :   0 - 0x0
      13'h2F0: dout <= 8'b00000000; //  752 :   0 - 0x0 -- Sprite 0x2f
      13'h2F1: dout <= 8'b00000000; //  753 :   0 - 0x0
      13'h2F2: dout <= 8'b00000000; //  754 :   0 - 0x0
      13'h2F3: dout <= 8'b00000000; //  755 :   0 - 0x0
      13'h2F4: dout <= 8'b00000000; //  756 :   0 - 0x0
      13'h2F5: dout <= 8'b00000000; //  757 :   0 - 0x0
      13'h2F6: dout <= 8'b00000000; //  758 :   0 - 0x0
      13'h2F7: dout <= 8'b00000000; //  759 :   0 - 0x0
      13'h2F8: dout <= 8'b00000000; //  760 :   0 - 0x0
      13'h2F9: dout <= 8'b00000000; //  761 :   0 - 0x0
      13'h2FA: dout <= 8'b00000000; //  762 :   0 - 0x0
      13'h2FB: dout <= 8'b00011000; //  763 :  24 - 0x18
      13'h2FC: dout <= 8'b00011000; //  764 :  24 - 0x18
      13'h2FD: dout <= 8'b00000000; //  765 :   0 - 0x0
      13'h2FE: dout <= 8'b00000000; //  766 :   0 - 0x0
      13'h2FF: dout <= 8'b00000000; //  767 :   0 - 0x0
      13'h300: dout <= 8'b00011100; //  768 :  28 - 0x1c -- Sprite 0x30
      13'h301: dout <= 8'b00100110; //  769 :  38 - 0x26
      13'h302: dout <= 8'b01100011; //  770 :  99 - 0x63
      13'h303: dout <= 8'b01100011; //  771 :  99 - 0x63
      13'h304: dout <= 8'b01100011; //  772 :  99 - 0x63
      13'h305: dout <= 8'b00110010; //  773 :  50 - 0x32
      13'h306: dout <= 8'b00011100; //  774 :  28 - 0x1c
      13'h307: dout <= 8'b00000000; //  775 :   0 - 0x0
      13'h308: dout <= 8'b00000000; //  776 :   0 - 0x0
      13'h309: dout <= 8'b00000000; //  777 :   0 - 0x0
      13'h30A: dout <= 8'b00000000; //  778 :   0 - 0x0
      13'h30B: dout <= 8'b00000000; //  779 :   0 - 0x0
      13'h30C: dout <= 8'b00000000; //  780 :   0 - 0x0
      13'h30D: dout <= 8'b00000000; //  781 :   0 - 0x0
      13'h30E: dout <= 8'b00000000; //  782 :   0 - 0x0
      13'h30F: dout <= 8'b00000000; //  783 :   0 - 0x0
      13'h310: dout <= 8'b00001100; //  784 :  12 - 0xc -- Sprite 0x31
      13'h311: dout <= 8'b00011100; //  785 :  28 - 0x1c
      13'h312: dout <= 8'b00001100; //  786 :  12 - 0xc
      13'h313: dout <= 8'b00001100; //  787 :  12 - 0xc
      13'h314: dout <= 8'b00001100; //  788 :  12 - 0xc
      13'h315: dout <= 8'b00001100; //  789 :  12 - 0xc
      13'h316: dout <= 8'b00111111; //  790 :  63 - 0x3f
      13'h317: dout <= 8'b00000000; //  791 :   0 - 0x0
      13'h318: dout <= 8'b00000000; //  792 :   0 - 0x0
      13'h319: dout <= 8'b00000000; //  793 :   0 - 0x0
      13'h31A: dout <= 8'b00000000; //  794 :   0 - 0x0
      13'h31B: dout <= 8'b00000000; //  795 :   0 - 0x0
      13'h31C: dout <= 8'b00000000; //  796 :   0 - 0x0
      13'h31D: dout <= 8'b00000000; //  797 :   0 - 0x0
      13'h31E: dout <= 8'b00000000; //  798 :   0 - 0x0
      13'h31F: dout <= 8'b00000000; //  799 :   0 - 0x0
      13'h320: dout <= 8'b00111110; //  800 :  62 - 0x3e -- Sprite 0x32
      13'h321: dout <= 8'b01100011; //  801 :  99 - 0x63
      13'h322: dout <= 8'b00000111; //  802 :   7 - 0x7
      13'h323: dout <= 8'b00011110; //  803 :  30 - 0x1e
      13'h324: dout <= 8'b00111100; //  804 :  60 - 0x3c
      13'h325: dout <= 8'b01110000; //  805 : 112 - 0x70
      13'h326: dout <= 8'b01111111; //  806 : 127 - 0x7f
      13'h327: dout <= 8'b00000000; //  807 :   0 - 0x0
      13'h328: dout <= 8'b00000000; //  808 :   0 - 0x0
      13'h329: dout <= 8'b00000000; //  809 :   0 - 0x0
      13'h32A: dout <= 8'b00000000; //  810 :   0 - 0x0
      13'h32B: dout <= 8'b00000000; //  811 :   0 - 0x0
      13'h32C: dout <= 8'b00000000; //  812 :   0 - 0x0
      13'h32D: dout <= 8'b00000000; //  813 :   0 - 0x0
      13'h32E: dout <= 8'b00000000; //  814 :   0 - 0x0
      13'h32F: dout <= 8'b00000000; //  815 :   0 - 0x0
      13'h330: dout <= 8'b00111111; //  816 :  63 - 0x3f -- Sprite 0x33
      13'h331: dout <= 8'b00000110; //  817 :   6 - 0x6
      13'h332: dout <= 8'b00001100; //  818 :  12 - 0xc
      13'h333: dout <= 8'b00011110; //  819 :  30 - 0x1e
      13'h334: dout <= 8'b00000011; //  820 :   3 - 0x3
      13'h335: dout <= 8'b01100011; //  821 :  99 - 0x63
      13'h336: dout <= 8'b00111110; //  822 :  62 - 0x3e
      13'h337: dout <= 8'b00000000; //  823 :   0 - 0x0
      13'h338: dout <= 8'b00000000; //  824 :   0 - 0x0
      13'h339: dout <= 8'b00000000; //  825 :   0 - 0x0
      13'h33A: dout <= 8'b00000000; //  826 :   0 - 0x0
      13'h33B: dout <= 8'b00000000; //  827 :   0 - 0x0
      13'h33C: dout <= 8'b00000000; //  828 :   0 - 0x0
      13'h33D: dout <= 8'b00000000; //  829 :   0 - 0x0
      13'h33E: dout <= 8'b00000000; //  830 :   0 - 0x0
      13'h33F: dout <= 8'b00000000; //  831 :   0 - 0x0
      13'h340: dout <= 8'b00001110; //  832 :  14 - 0xe -- Sprite 0x34
      13'h341: dout <= 8'b00011110; //  833 :  30 - 0x1e
      13'h342: dout <= 8'b00110110; //  834 :  54 - 0x36
      13'h343: dout <= 8'b01100110; //  835 : 102 - 0x66
      13'h344: dout <= 8'b01111111; //  836 : 127 - 0x7f
      13'h345: dout <= 8'b00000110; //  837 :   6 - 0x6
      13'h346: dout <= 8'b00000110; //  838 :   6 - 0x6
      13'h347: dout <= 8'b00000000; //  839 :   0 - 0x0
      13'h348: dout <= 8'b00000000; //  840 :   0 - 0x0
      13'h349: dout <= 8'b00000000; //  841 :   0 - 0x0
      13'h34A: dout <= 8'b00000000; //  842 :   0 - 0x0
      13'h34B: dout <= 8'b00000000; //  843 :   0 - 0x0
      13'h34C: dout <= 8'b00000000; //  844 :   0 - 0x0
      13'h34D: dout <= 8'b00000000; //  845 :   0 - 0x0
      13'h34E: dout <= 8'b00000000; //  846 :   0 - 0x0
      13'h34F: dout <= 8'b00000000; //  847 :   0 - 0x0
      13'h350: dout <= 8'b01111110; //  848 : 126 - 0x7e -- Sprite 0x35
      13'h351: dout <= 8'b01100000; //  849 :  96 - 0x60
      13'h352: dout <= 8'b01111110; //  850 : 126 - 0x7e
      13'h353: dout <= 8'b00000011; //  851 :   3 - 0x3
      13'h354: dout <= 8'b00000011; //  852 :   3 - 0x3
      13'h355: dout <= 8'b01100011; //  853 :  99 - 0x63
      13'h356: dout <= 8'b00111110; //  854 :  62 - 0x3e
      13'h357: dout <= 8'b00000000; //  855 :   0 - 0x0
      13'h358: dout <= 8'b00000000; //  856 :   0 - 0x0
      13'h359: dout <= 8'b00000000; //  857 :   0 - 0x0
      13'h35A: dout <= 8'b00000000; //  858 :   0 - 0x0
      13'h35B: dout <= 8'b00000000; //  859 :   0 - 0x0
      13'h35C: dout <= 8'b00000000; //  860 :   0 - 0x0
      13'h35D: dout <= 8'b00000000; //  861 :   0 - 0x0
      13'h35E: dout <= 8'b00000000; //  862 :   0 - 0x0
      13'h35F: dout <= 8'b00000000; //  863 :   0 - 0x0
      13'h360: dout <= 8'b00011110; //  864 :  30 - 0x1e -- Sprite 0x36
      13'h361: dout <= 8'b00110000; //  865 :  48 - 0x30
      13'h362: dout <= 8'b01100000; //  866 :  96 - 0x60
      13'h363: dout <= 8'b01111110; //  867 : 126 - 0x7e
      13'h364: dout <= 8'b01100011; //  868 :  99 - 0x63
      13'h365: dout <= 8'b01100011; //  869 :  99 - 0x63
      13'h366: dout <= 8'b00111110; //  870 :  62 - 0x3e
      13'h367: dout <= 8'b00000000; //  871 :   0 - 0x0
      13'h368: dout <= 8'b00000000; //  872 :   0 - 0x0
      13'h369: dout <= 8'b00000000; //  873 :   0 - 0x0
      13'h36A: dout <= 8'b00000000; //  874 :   0 - 0x0
      13'h36B: dout <= 8'b00000000; //  875 :   0 - 0x0
      13'h36C: dout <= 8'b00000000; //  876 :   0 - 0x0
      13'h36D: dout <= 8'b00000000; //  877 :   0 - 0x0
      13'h36E: dout <= 8'b00000000; //  878 :   0 - 0x0
      13'h36F: dout <= 8'b00000000; //  879 :   0 - 0x0
      13'h370: dout <= 8'b01111111; //  880 : 127 - 0x7f -- Sprite 0x37
      13'h371: dout <= 8'b01100011; //  881 :  99 - 0x63
      13'h372: dout <= 8'b00000110; //  882 :   6 - 0x6
      13'h373: dout <= 8'b00001100; //  883 :  12 - 0xc
      13'h374: dout <= 8'b00011000; //  884 :  24 - 0x18
      13'h375: dout <= 8'b00011000; //  885 :  24 - 0x18
      13'h376: dout <= 8'b00011000; //  886 :  24 - 0x18
      13'h377: dout <= 8'b00000000; //  887 :   0 - 0x0
      13'h378: dout <= 8'b00000000; //  888 :   0 - 0x0
      13'h379: dout <= 8'b00000000; //  889 :   0 - 0x0
      13'h37A: dout <= 8'b00000000; //  890 :   0 - 0x0
      13'h37B: dout <= 8'b00000000; //  891 :   0 - 0x0
      13'h37C: dout <= 8'b00000000; //  892 :   0 - 0x0
      13'h37D: dout <= 8'b00000000; //  893 :   0 - 0x0
      13'h37E: dout <= 8'b00000000; //  894 :   0 - 0x0
      13'h37F: dout <= 8'b00000000; //  895 :   0 - 0x0
      13'h380: dout <= 8'b00111100; //  896 :  60 - 0x3c -- Sprite 0x38
      13'h381: dout <= 8'b01100010; //  897 :  98 - 0x62
      13'h382: dout <= 8'b01110010; //  898 : 114 - 0x72
      13'h383: dout <= 8'b00111100; //  899 :  60 - 0x3c
      13'h384: dout <= 8'b01001111; //  900 :  79 - 0x4f
      13'h385: dout <= 8'b01000011; //  901 :  67 - 0x43
      13'h386: dout <= 8'b00111110; //  902 :  62 - 0x3e
      13'h387: dout <= 8'b00000000; //  903 :   0 - 0x0
      13'h388: dout <= 8'b00000000; //  904 :   0 - 0x0
      13'h389: dout <= 8'b00000000; //  905 :   0 - 0x0
      13'h38A: dout <= 8'b00000000; //  906 :   0 - 0x0
      13'h38B: dout <= 8'b00000000; //  907 :   0 - 0x0
      13'h38C: dout <= 8'b00000000; //  908 :   0 - 0x0
      13'h38D: dout <= 8'b00000000; //  909 :   0 - 0x0
      13'h38E: dout <= 8'b00000000; //  910 :   0 - 0x0
      13'h38F: dout <= 8'b00000000; //  911 :   0 - 0x0
      13'h390: dout <= 8'b00111110; //  912 :  62 - 0x3e -- Sprite 0x39
      13'h391: dout <= 8'b01100011; //  913 :  99 - 0x63
      13'h392: dout <= 8'b01100011; //  914 :  99 - 0x63
      13'h393: dout <= 8'b00111111; //  915 :  63 - 0x3f
      13'h394: dout <= 8'b00000011; //  916 :   3 - 0x3
      13'h395: dout <= 8'b00000110; //  917 :   6 - 0x6
      13'h396: dout <= 8'b00111100; //  918 :  60 - 0x3c
      13'h397: dout <= 8'b00000000; //  919 :   0 - 0x0
      13'h398: dout <= 8'b00000000; //  920 :   0 - 0x0
      13'h399: dout <= 8'b00000000; //  921 :   0 - 0x0
      13'h39A: dout <= 8'b00000000; //  922 :   0 - 0x0
      13'h39B: dout <= 8'b00000000; //  923 :   0 - 0x0
      13'h39C: dout <= 8'b00000000; //  924 :   0 - 0x0
      13'h39D: dout <= 8'b00000000; //  925 :   0 - 0x0
      13'h39E: dout <= 8'b00000000; //  926 :   0 - 0x0
      13'h39F: dout <= 8'b00000000; //  927 :   0 - 0x0
      13'h3A0: dout <= 8'b00000000; //  928 :   0 - 0x0 -- Sprite 0x3a
      13'h3A1: dout <= 8'b00000000; //  929 :   0 - 0x0
      13'h3A2: dout <= 8'b00000000; //  930 :   0 - 0x0
      13'h3A3: dout <= 8'b01111110; //  931 : 126 - 0x7e
      13'h3A4: dout <= 8'b00000000; //  932 :   0 - 0x0
      13'h3A5: dout <= 8'b00000000; //  933 :   0 - 0x0
      13'h3A6: dout <= 8'b00000000; //  934 :   0 - 0x0
      13'h3A7: dout <= 8'b00000000; //  935 :   0 - 0x0
      13'h3A8: dout <= 8'b00000000; //  936 :   0 - 0x0
      13'h3A9: dout <= 8'b00000000; //  937 :   0 - 0x0
      13'h3AA: dout <= 8'b00000000; //  938 :   0 - 0x0
      13'h3AB: dout <= 8'b00000000; //  939 :   0 - 0x0
      13'h3AC: dout <= 8'b00000000; //  940 :   0 - 0x0
      13'h3AD: dout <= 8'b00000000; //  941 :   0 - 0x0
      13'h3AE: dout <= 8'b00000000; //  942 :   0 - 0x0
      13'h3AF: dout <= 8'b00000000; //  943 :   0 - 0x0
      13'h3B0: dout <= 8'b00000000; //  944 :   0 - 0x0 -- Sprite 0x3b
      13'h3B1: dout <= 8'b00000010; //  945 :   2 - 0x2
      13'h3B2: dout <= 8'b00000100; //  946 :   4 - 0x4
      13'h3B3: dout <= 8'b00001000; //  947 :   8 - 0x8
      13'h3B4: dout <= 8'b00010000; //  948 :  16 - 0x10
      13'h3B5: dout <= 8'b00100000; //  949 :  32 - 0x20
      13'h3B6: dout <= 8'b00000000; //  950 :   0 - 0x0
      13'h3B7: dout <= 8'b00000000; //  951 :   0 - 0x0
      13'h3B8: dout <= 8'b00000000; //  952 :   0 - 0x0
      13'h3B9: dout <= 8'b00000000; //  953 :   0 - 0x0
      13'h3BA: dout <= 8'b00000000; //  954 :   0 - 0x0
      13'h3BB: dout <= 8'b00000000; //  955 :   0 - 0x0
      13'h3BC: dout <= 8'b00000000; //  956 :   0 - 0x0
      13'h3BD: dout <= 8'b00000000; //  957 :   0 - 0x0
      13'h3BE: dout <= 8'b00000000; //  958 :   0 - 0x0
      13'h3BF: dout <= 8'b00000000; //  959 :   0 - 0x0
      13'h3C0: dout <= 8'b00000000; //  960 :   0 - 0x0 -- Sprite 0x3c
      13'h3C1: dout <= 8'b00000111; //  961 :   7 - 0x7
      13'h3C2: dout <= 8'b00011111; //  962 :  31 - 0x1f
      13'h3C3: dout <= 8'b00111111; //  963 :  63 - 0x3f
      13'h3C4: dout <= 8'b00111111; //  964 :  63 - 0x3f
      13'h3C5: dout <= 8'b00001111; //  965 :  15 - 0xf
      13'h3C6: dout <= 8'b00000011; //  966 :   3 - 0x3
      13'h3C7: dout <= 8'b00000000; //  967 :   0 - 0x0
      13'h3C8: dout <= 8'b00000000; //  968 :   0 - 0x0
      13'h3C9: dout <= 8'b00000111; //  969 :   7 - 0x7
      13'h3CA: dout <= 8'b00011111; //  970 :  31 - 0x1f
      13'h3CB: dout <= 8'b00111111; //  971 :  63 - 0x3f
      13'h3CC: dout <= 8'b00111111; //  972 :  63 - 0x3f
      13'h3CD: dout <= 8'b00001111; //  973 :  15 - 0xf
      13'h3CE: dout <= 8'b00000011; //  974 :   3 - 0x3
      13'h3CF: dout <= 8'b00000000; //  975 :   0 - 0x0
      13'h3D0: dout <= 8'b00000000; //  976 :   0 - 0x0 -- Sprite 0x3d
      13'h3D1: dout <= 8'b11000000; //  977 : 192 - 0xc0
      13'h3D2: dout <= 8'b11110000; //  978 : 240 - 0xf0
      13'h3D3: dout <= 8'b11111000; //  979 : 248 - 0xf8
      13'h3D4: dout <= 8'b11111000; //  980 : 248 - 0xf8
      13'h3D5: dout <= 8'b11111100; //  981 : 252 - 0xfc
      13'h3D6: dout <= 8'b11111100; //  982 : 252 - 0xfc
      13'h3D7: dout <= 8'b11111100; //  983 : 252 - 0xfc
      13'h3D8: dout <= 8'b00000000; //  984 :   0 - 0x0
      13'h3D9: dout <= 8'b11000000; //  985 : 192 - 0xc0
      13'h3DA: dout <= 8'b11110000; //  986 : 240 - 0xf0
      13'h3DB: dout <= 8'b11111000; //  987 : 248 - 0xf8
      13'h3DC: dout <= 8'b11111000; //  988 : 248 - 0xf8
      13'h3DD: dout <= 8'b11111100; //  989 : 252 - 0xfc
      13'h3DE: dout <= 8'b11111100; //  990 : 252 - 0xfc
      13'h3DF: dout <= 8'b11111100; //  991 : 252 - 0xfc
      13'h3E0: dout <= 8'b00000000; //  992 :   0 - 0x0 -- Sprite 0x3e
      13'h3E1: dout <= 8'b00000011; //  993 :   3 - 0x3
      13'h3E2: dout <= 8'b00001111; //  994 :  15 - 0xf
      13'h3E3: dout <= 8'b00111111; //  995 :  63 - 0x3f
      13'h3E4: dout <= 8'b00111111; //  996 :  63 - 0x3f
      13'h3E5: dout <= 8'b00011111; //  997 :  31 - 0x1f
      13'h3E6: dout <= 8'b00000111; //  998 :   7 - 0x7
      13'h3E7: dout <= 8'b00000000; //  999 :   0 - 0x0
      13'h3E8: dout <= 8'b00000000; // 1000 :   0 - 0x0
      13'h3E9: dout <= 8'b00000011; // 1001 :   3 - 0x3
      13'h3EA: dout <= 8'b00001111; // 1002 :  15 - 0xf
      13'h3EB: dout <= 8'b00111111; // 1003 :  63 - 0x3f
      13'h3EC: dout <= 8'b00111111; // 1004 :  63 - 0x3f
      13'h3ED: dout <= 8'b00011111; // 1005 :  31 - 0x1f
      13'h3EE: dout <= 8'b00000111; // 1006 :   7 - 0x7
      13'h3EF: dout <= 8'b00000000; // 1007 :   0 - 0x0
      13'h3F0: dout <= 8'b11111100; // 1008 : 252 - 0xfc -- Sprite 0x3f
      13'h3F1: dout <= 8'b11111100; // 1009 : 252 - 0xfc
      13'h3F2: dout <= 8'b11111100; // 1010 : 252 - 0xfc
      13'h3F3: dout <= 8'b11111000; // 1011 : 248 - 0xf8
      13'h3F4: dout <= 8'b11111000; // 1012 : 248 - 0xf8
      13'h3F5: dout <= 8'b11110000; // 1013 : 240 - 0xf0
      13'h3F6: dout <= 8'b11000000; // 1014 : 192 - 0xc0
      13'h3F7: dout <= 8'b00000000; // 1015 :   0 - 0x0
      13'h3F8: dout <= 8'b11111100; // 1016 : 252 - 0xfc
      13'h3F9: dout <= 8'b11111100; // 1017 : 252 - 0xfc
      13'h3FA: dout <= 8'b11111100; // 1018 : 252 - 0xfc
      13'h3FB: dout <= 8'b11111000; // 1019 : 248 - 0xf8
      13'h3FC: dout <= 8'b11111000; // 1020 : 248 - 0xf8
      13'h3FD: dout <= 8'b11110000; // 1021 : 240 - 0xf0
      13'h3FE: dout <= 8'b11000000; // 1022 : 192 - 0xc0
      13'h3FF: dout <= 8'b00000000; // 1023 :   0 - 0x0
      13'h400: dout <= 8'b00000000; // 1024 :   0 - 0x0 -- Sprite 0x40
      13'h401: dout <= 8'b00000000; // 1025 :   0 - 0x0
      13'h402: dout <= 8'b00000000; // 1026 :   0 - 0x0
      13'h403: dout <= 8'b00000000; // 1027 :   0 - 0x0
      13'h404: dout <= 8'b00000000; // 1028 :   0 - 0x0
      13'h405: dout <= 8'b00000000; // 1029 :   0 - 0x0
      13'h406: dout <= 8'b00000000; // 1030 :   0 - 0x0
      13'h407: dout <= 8'b00000000; // 1031 :   0 - 0x0
      13'h408: dout <= 8'b00000000; // 1032 :   0 - 0x0
      13'h409: dout <= 8'b00000000; // 1033 :   0 - 0x0
      13'h40A: dout <= 8'b00000000; // 1034 :   0 - 0x0
      13'h40B: dout <= 8'b00000000; // 1035 :   0 - 0x0
      13'h40C: dout <= 8'b00000000; // 1036 :   0 - 0x0
      13'h40D: dout <= 8'b00000000; // 1037 :   0 - 0x0
      13'h40E: dout <= 8'b00000000; // 1038 :   0 - 0x0
      13'h40F: dout <= 8'b00000000; // 1039 :   0 - 0x0
      13'h410: dout <= 8'b00011100; // 1040 :  28 - 0x1c -- Sprite 0x41
      13'h411: dout <= 8'b00110110; // 1041 :  54 - 0x36
      13'h412: dout <= 8'b01100011; // 1042 :  99 - 0x63
      13'h413: dout <= 8'b01100011; // 1043 :  99 - 0x63
      13'h414: dout <= 8'b01111111; // 1044 : 127 - 0x7f
      13'h415: dout <= 8'b01100011; // 1045 :  99 - 0x63
      13'h416: dout <= 8'b01100011; // 1046 :  99 - 0x63
      13'h417: dout <= 8'b00000000; // 1047 :   0 - 0x0
      13'h418: dout <= 8'b00000000; // 1048 :   0 - 0x0
      13'h419: dout <= 8'b00000000; // 1049 :   0 - 0x0
      13'h41A: dout <= 8'b00000000; // 1050 :   0 - 0x0
      13'h41B: dout <= 8'b00000000; // 1051 :   0 - 0x0
      13'h41C: dout <= 8'b00000000; // 1052 :   0 - 0x0
      13'h41D: dout <= 8'b00000000; // 1053 :   0 - 0x0
      13'h41E: dout <= 8'b00000000; // 1054 :   0 - 0x0
      13'h41F: dout <= 8'b00000000; // 1055 :   0 - 0x0
      13'h420: dout <= 8'b01111110; // 1056 : 126 - 0x7e -- Sprite 0x42
      13'h421: dout <= 8'b01100011; // 1057 :  99 - 0x63
      13'h422: dout <= 8'b01100011; // 1058 :  99 - 0x63
      13'h423: dout <= 8'b01111110; // 1059 : 126 - 0x7e
      13'h424: dout <= 8'b01100011; // 1060 :  99 - 0x63
      13'h425: dout <= 8'b01100011; // 1061 :  99 - 0x63
      13'h426: dout <= 8'b01111110; // 1062 : 126 - 0x7e
      13'h427: dout <= 8'b00000000; // 1063 :   0 - 0x0
      13'h428: dout <= 8'b00000000; // 1064 :   0 - 0x0
      13'h429: dout <= 8'b00000000; // 1065 :   0 - 0x0
      13'h42A: dout <= 8'b00000000; // 1066 :   0 - 0x0
      13'h42B: dout <= 8'b00000000; // 1067 :   0 - 0x0
      13'h42C: dout <= 8'b00000000; // 1068 :   0 - 0x0
      13'h42D: dout <= 8'b00000000; // 1069 :   0 - 0x0
      13'h42E: dout <= 8'b00000000; // 1070 :   0 - 0x0
      13'h42F: dout <= 8'b00000000; // 1071 :   0 - 0x0
      13'h430: dout <= 8'b00011110; // 1072 :  30 - 0x1e -- Sprite 0x43
      13'h431: dout <= 8'b00110011; // 1073 :  51 - 0x33
      13'h432: dout <= 8'b01100000; // 1074 :  96 - 0x60
      13'h433: dout <= 8'b01100000; // 1075 :  96 - 0x60
      13'h434: dout <= 8'b01100000; // 1076 :  96 - 0x60
      13'h435: dout <= 8'b00110011; // 1077 :  51 - 0x33
      13'h436: dout <= 8'b00011110; // 1078 :  30 - 0x1e
      13'h437: dout <= 8'b00000000; // 1079 :   0 - 0x0
      13'h438: dout <= 8'b00000000; // 1080 :   0 - 0x0
      13'h439: dout <= 8'b00000000; // 1081 :   0 - 0x0
      13'h43A: dout <= 8'b00000000; // 1082 :   0 - 0x0
      13'h43B: dout <= 8'b00000000; // 1083 :   0 - 0x0
      13'h43C: dout <= 8'b00000000; // 1084 :   0 - 0x0
      13'h43D: dout <= 8'b00000000; // 1085 :   0 - 0x0
      13'h43E: dout <= 8'b00000000; // 1086 :   0 - 0x0
      13'h43F: dout <= 8'b00000000; // 1087 :   0 - 0x0
      13'h440: dout <= 8'b01111100; // 1088 : 124 - 0x7c -- Sprite 0x44
      13'h441: dout <= 8'b01100110; // 1089 : 102 - 0x66
      13'h442: dout <= 8'b01100011; // 1090 :  99 - 0x63
      13'h443: dout <= 8'b01100011; // 1091 :  99 - 0x63
      13'h444: dout <= 8'b01100011; // 1092 :  99 - 0x63
      13'h445: dout <= 8'b01100110; // 1093 : 102 - 0x66
      13'h446: dout <= 8'b01111100; // 1094 : 124 - 0x7c
      13'h447: dout <= 8'b00000000; // 1095 :   0 - 0x0
      13'h448: dout <= 8'b00000000; // 1096 :   0 - 0x0
      13'h449: dout <= 8'b00000000; // 1097 :   0 - 0x0
      13'h44A: dout <= 8'b00000000; // 1098 :   0 - 0x0
      13'h44B: dout <= 8'b00000000; // 1099 :   0 - 0x0
      13'h44C: dout <= 8'b00000000; // 1100 :   0 - 0x0
      13'h44D: dout <= 8'b00000000; // 1101 :   0 - 0x0
      13'h44E: dout <= 8'b00000000; // 1102 :   0 - 0x0
      13'h44F: dout <= 8'b00000000; // 1103 :   0 - 0x0
      13'h450: dout <= 8'b01111111; // 1104 : 127 - 0x7f -- Sprite 0x45
      13'h451: dout <= 8'b01100000; // 1105 :  96 - 0x60
      13'h452: dout <= 8'b01100000; // 1106 :  96 - 0x60
      13'h453: dout <= 8'b01111110; // 1107 : 126 - 0x7e
      13'h454: dout <= 8'b01100000; // 1108 :  96 - 0x60
      13'h455: dout <= 8'b01100000; // 1109 :  96 - 0x60
      13'h456: dout <= 8'b01111111; // 1110 : 127 - 0x7f
      13'h457: dout <= 8'b00000000; // 1111 :   0 - 0x0
      13'h458: dout <= 8'b00000000; // 1112 :   0 - 0x0
      13'h459: dout <= 8'b00000000; // 1113 :   0 - 0x0
      13'h45A: dout <= 8'b00000000; // 1114 :   0 - 0x0
      13'h45B: dout <= 8'b00000000; // 1115 :   0 - 0x0
      13'h45C: dout <= 8'b00000000; // 1116 :   0 - 0x0
      13'h45D: dout <= 8'b00000000; // 1117 :   0 - 0x0
      13'h45E: dout <= 8'b00000000; // 1118 :   0 - 0x0
      13'h45F: dout <= 8'b00000000; // 1119 :   0 - 0x0
      13'h460: dout <= 8'b01111111; // 1120 : 127 - 0x7f -- Sprite 0x46
      13'h461: dout <= 8'b01100000; // 1121 :  96 - 0x60
      13'h462: dout <= 8'b01100000; // 1122 :  96 - 0x60
      13'h463: dout <= 8'b01111110; // 1123 : 126 - 0x7e
      13'h464: dout <= 8'b01100000; // 1124 :  96 - 0x60
      13'h465: dout <= 8'b01100000; // 1125 :  96 - 0x60
      13'h466: dout <= 8'b01100000; // 1126 :  96 - 0x60
      13'h467: dout <= 8'b00000000; // 1127 :   0 - 0x0
      13'h468: dout <= 8'b00000000; // 1128 :   0 - 0x0
      13'h469: dout <= 8'b00000000; // 1129 :   0 - 0x0
      13'h46A: dout <= 8'b00000000; // 1130 :   0 - 0x0
      13'h46B: dout <= 8'b00000000; // 1131 :   0 - 0x0
      13'h46C: dout <= 8'b00000000; // 1132 :   0 - 0x0
      13'h46D: dout <= 8'b00000000; // 1133 :   0 - 0x0
      13'h46E: dout <= 8'b00000000; // 1134 :   0 - 0x0
      13'h46F: dout <= 8'b00000000; // 1135 :   0 - 0x0
      13'h470: dout <= 8'b00011111; // 1136 :  31 - 0x1f -- Sprite 0x47
      13'h471: dout <= 8'b00110000; // 1137 :  48 - 0x30
      13'h472: dout <= 8'b01100000; // 1138 :  96 - 0x60
      13'h473: dout <= 8'b01100111; // 1139 : 103 - 0x67
      13'h474: dout <= 8'b01100011; // 1140 :  99 - 0x63
      13'h475: dout <= 8'b00110011; // 1141 :  51 - 0x33
      13'h476: dout <= 8'b00011111; // 1142 :  31 - 0x1f
      13'h477: dout <= 8'b00000000; // 1143 :   0 - 0x0
      13'h478: dout <= 8'b00000000; // 1144 :   0 - 0x0
      13'h479: dout <= 8'b00000000; // 1145 :   0 - 0x0
      13'h47A: dout <= 8'b00000000; // 1146 :   0 - 0x0
      13'h47B: dout <= 8'b00000000; // 1147 :   0 - 0x0
      13'h47C: dout <= 8'b00000000; // 1148 :   0 - 0x0
      13'h47D: dout <= 8'b00000000; // 1149 :   0 - 0x0
      13'h47E: dout <= 8'b00000000; // 1150 :   0 - 0x0
      13'h47F: dout <= 8'b00000000; // 1151 :   0 - 0x0
      13'h480: dout <= 8'b01100011; // 1152 :  99 - 0x63 -- Sprite 0x48
      13'h481: dout <= 8'b01100011; // 1153 :  99 - 0x63
      13'h482: dout <= 8'b01100011; // 1154 :  99 - 0x63
      13'h483: dout <= 8'b01111111; // 1155 : 127 - 0x7f
      13'h484: dout <= 8'b01100011; // 1156 :  99 - 0x63
      13'h485: dout <= 8'b01100011; // 1157 :  99 - 0x63
      13'h486: dout <= 8'b01100011; // 1158 :  99 - 0x63
      13'h487: dout <= 8'b00000000; // 1159 :   0 - 0x0
      13'h488: dout <= 8'b00000000; // 1160 :   0 - 0x0
      13'h489: dout <= 8'b00000000; // 1161 :   0 - 0x0
      13'h48A: dout <= 8'b00000000; // 1162 :   0 - 0x0
      13'h48B: dout <= 8'b00000000; // 1163 :   0 - 0x0
      13'h48C: dout <= 8'b00000000; // 1164 :   0 - 0x0
      13'h48D: dout <= 8'b00000000; // 1165 :   0 - 0x0
      13'h48E: dout <= 8'b00000000; // 1166 :   0 - 0x0
      13'h48F: dout <= 8'b00000000; // 1167 :   0 - 0x0
      13'h490: dout <= 8'b00111111; // 1168 :  63 - 0x3f -- Sprite 0x49
      13'h491: dout <= 8'b00001100; // 1169 :  12 - 0xc
      13'h492: dout <= 8'b00001100; // 1170 :  12 - 0xc
      13'h493: dout <= 8'b00001100; // 1171 :  12 - 0xc
      13'h494: dout <= 8'b00001100; // 1172 :  12 - 0xc
      13'h495: dout <= 8'b00001100; // 1173 :  12 - 0xc
      13'h496: dout <= 8'b00111111; // 1174 :  63 - 0x3f
      13'h497: dout <= 8'b00000000; // 1175 :   0 - 0x0
      13'h498: dout <= 8'b00000000; // 1176 :   0 - 0x0
      13'h499: dout <= 8'b00000000; // 1177 :   0 - 0x0
      13'h49A: dout <= 8'b00000000; // 1178 :   0 - 0x0
      13'h49B: dout <= 8'b00000000; // 1179 :   0 - 0x0
      13'h49C: dout <= 8'b00000000; // 1180 :   0 - 0x0
      13'h49D: dout <= 8'b00000000; // 1181 :   0 - 0x0
      13'h49E: dout <= 8'b00000000; // 1182 :   0 - 0x0
      13'h49F: dout <= 8'b00000000; // 1183 :   0 - 0x0
      13'h4A0: dout <= 8'b00000011; // 1184 :   3 - 0x3 -- Sprite 0x4a
      13'h4A1: dout <= 8'b00000011; // 1185 :   3 - 0x3
      13'h4A2: dout <= 8'b00000011; // 1186 :   3 - 0x3
      13'h4A3: dout <= 8'b00000011; // 1187 :   3 - 0x3
      13'h4A4: dout <= 8'b00000011; // 1188 :   3 - 0x3
      13'h4A5: dout <= 8'b01100011; // 1189 :  99 - 0x63
      13'h4A6: dout <= 8'b00111110; // 1190 :  62 - 0x3e
      13'h4A7: dout <= 8'b00000000; // 1191 :   0 - 0x0
      13'h4A8: dout <= 8'b00000000; // 1192 :   0 - 0x0
      13'h4A9: dout <= 8'b00000000; // 1193 :   0 - 0x0
      13'h4AA: dout <= 8'b00000000; // 1194 :   0 - 0x0
      13'h4AB: dout <= 8'b00000000; // 1195 :   0 - 0x0
      13'h4AC: dout <= 8'b00000000; // 1196 :   0 - 0x0
      13'h4AD: dout <= 8'b00000000; // 1197 :   0 - 0x0
      13'h4AE: dout <= 8'b00000000; // 1198 :   0 - 0x0
      13'h4AF: dout <= 8'b00000000; // 1199 :   0 - 0x0
      13'h4B0: dout <= 8'b01100011; // 1200 :  99 - 0x63 -- Sprite 0x4b
      13'h4B1: dout <= 8'b01100110; // 1201 : 102 - 0x66
      13'h4B2: dout <= 8'b01101100; // 1202 : 108 - 0x6c
      13'h4B3: dout <= 8'b01111000; // 1203 : 120 - 0x78
      13'h4B4: dout <= 8'b01111100; // 1204 : 124 - 0x7c
      13'h4B5: dout <= 8'b01100110; // 1205 : 102 - 0x66
      13'h4B6: dout <= 8'b01100011; // 1206 :  99 - 0x63
      13'h4B7: dout <= 8'b00000000; // 1207 :   0 - 0x0
      13'h4B8: dout <= 8'b00000000; // 1208 :   0 - 0x0
      13'h4B9: dout <= 8'b00000000; // 1209 :   0 - 0x0
      13'h4BA: dout <= 8'b00000000; // 1210 :   0 - 0x0
      13'h4BB: dout <= 8'b00000000; // 1211 :   0 - 0x0
      13'h4BC: dout <= 8'b00000000; // 1212 :   0 - 0x0
      13'h4BD: dout <= 8'b00000000; // 1213 :   0 - 0x0
      13'h4BE: dout <= 8'b00000000; // 1214 :   0 - 0x0
      13'h4BF: dout <= 8'b00000000; // 1215 :   0 - 0x0
      13'h4C0: dout <= 8'b01100000; // 1216 :  96 - 0x60 -- Sprite 0x4c
      13'h4C1: dout <= 8'b01100000; // 1217 :  96 - 0x60
      13'h4C2: dout <= 8'b01100000; // 1218 :  96 - 0x60
      13'h4C3: dout <= 8'b01100000; // 1219 :  96 - 0x60
      13'h4C4: dout <= 8'b01100000; // 1220 :  96 - 0x60
      13'h4C5: dout <= 8'b01100000; // 1221 :  96 - 0x60
      13'h4C6: dout <= 8'b01111111; // 1222 : 127 - 0x7f
      13'h4C7: dout <= 8'b00000000; // 1223 :   0 - 0x0
      13'h4C8: dout <= 8'b00000000; // 1224 :   0 - 0x0
      13'h4C9: dout <= 8'b00000000; // 1225 :   0 - 0x0
      13'h4CA: dout <= 8'b00000000; // 1226 :   0 - 0x0
      13'h4CB: dout <= 8'b00000000; // 1227 :   0 - 0x0
      13'h4CC: dout <= 8'b00000000; // 1228 :   0 - 0x0
      13'h4CD: dout <= 8'b00000000; // 1229 :   0 - 0x0
      13'h4CE: dout <= 8'b00000000; // 1230 :   0 - 0x0
      13'h4CF: dout <= 8'b00000000; // 1231 :   0 - 0x0
      13'h4D0: dout <= 8'b01100011; // 1232 :  99 - 0x63 -- Sprite 0x4d
      13'h4D1: dout <= 8'b01110111; // 1233 : 119 - 0x77
      13'h4D2: dout <= 8'b01111111; // 1234 : 127 - 0x7f
      13'h4D3: dout <= 8'b01111111; // 1235 : 127 - 0x7f
      13'h4D4: dout <= 8'b01101011; // 1236 : 107 - 0x6b
      13'h4D5: dout <= 8'b01100011; // 1237 :  99 - 0x63
      13'h4D6: dout <= 8'b01100011; // 1238 :  99 - 0x63
      13'h4D7: dout <= 8'b00000000; // 1239 :   0 - 0x0
      13'h4D8: dout <= 8'b00000000; // 1240 :   0 - 0x0
      13'h4D9: dout <= 8'b00000000; // 1241 :   0 - 0x0
      13'h4DA: dout <= 8'b00000000; // 1242 :   0 - 0x0
      13'h4DB: dout <= 8'b00000000; // 1243 :   0 - 0x0
      13'h4DC: dout <= 8'b00000000; // 1244 :   0 - 0x0
      13'h4DD: dout <= 8'b00000000; // 1245 :   0 - 0x0
      13'h4DE: dout <= 8'b00000000; // 1246 :   0 - 0x0
      13'h4DF: dout <= 8'b00000000; // 1247 :   0 - 0x0
      13'h4E0: dout <= 8'b01100011; // 1248 :  99 - 0x63 -- Sprite 0x4e
      13'h4E1: dout <= 8'b01110011; // 1249 : 115 - 0x73
      13'h4E2: dout <= 8'b01111011; // 1250 : 123 - 0x7b
      13'h4E3: dout <= 8'b01111111; // 1251 : 127 - 0x7f
      13'h4E4: dout <= 8'b01101111; // 1252 : 111 - 0x6f
      13'h4E5: dout <= 8'b01100111; // 1253 : 103 - 0x67
      13'h4E6: dout <= 8'b01100011; // 1254 :  99 - 0x63
      13'h4E7: dout <= 8'b00000000; // 1255 :   0 - 0x0
      13'h4E8: dout <= 8'b00000000; // 1256 :   0 - 0x0
      13'h4E9: dout <= 8'b00000000; // 1257 :   0 - 0x0
      13'h4EA: dout <= 8'b00000000; // 1258 :   0 - 0x0
      13'h4EB: dout <= 8'b00000000; // 1259 :   0 - 0x0
      13'h4EC: dout <= 8'b00000000; // 1260 :   0 - 0x0
      13'h4ED: dout <= 8'b00000000; // 1261 :   0 - 0x0
      13'h4EE: dout <= 8'b00000000; // 1262 :   0 - 0x0
      13'h4EF: dout <= 8'b00000000; // 1263 :   0 - 0x0
      13'h4F0: dout <= 8'b00111110; // 1264 :  62 - 0x3e -- Sprite 0x4f
      13'h4F1: dout <= 8'b01100011; // 1265 :  99 - 0x63
      13'h4F2: dout <= 8'b01100011; // 1266 :  99 - 0x63
      13'h4F3: dout <= 8'b01100011; // 1267 :  99 - 0x63
      13'h4F4: dout <= 8'b01100011; // 1268 :  99 - 0x63
      13'h4F5: dout <= 8'b01100011; // 1269 :  99 - 0x63
      13'h4F6: dout <= 8'b00111110; // 1270 :  62 - 0x3e
      13'h4F7: dout <= 8'b00000000; // 1271 :   0 - 0x0
      13'h4F8: dout <= 8'b00000000; // 1272 :   0 - 0x0
      13'h4F9: dout <= 8'b00000000; // 1273 :   0 - 0x0
      13'h4FA: dout <= 8'b00000000; // 1274 :   0 - 0x0
      13'h4FB: dout <= 8'b00000000; // 1275 :   0 - 0x0
      13'h4FC: dout <= 8'b00000000; // 1276 :   0 - 0x0
      13'h4FD: dout <= 8'b00000000; // 1277 :   0 - 0x0
      13'h4FE: dout <= 8'b00000000; // 1278 :   0 - 0x0
      13'h4FF: dout <= 8'b00000000; // 1279 :   0 - 0x0
      13'h500: dout <= 8'b01111110; // 1280 : 126 - 0x7e -- Sprite 0x50
      13'h501: dout <= 8'b01100011; // 1281 :  99 - 0x63
      13'h502: dout <= 8'b01100011; // 1282 :  99 - 0x63
      13'h503: dout <= 8'b01100011; // 1283 :  99 - 0x63
      13'h504: dout <= 8'b01111110; // 1284 : 126 - 0x7e
      13'h505: dout <= 8'b01100000; // 1285 :  96 - 0x60
      13'h506: dout <= 8'b01100000; // 1286 :  96 - 0x60
      13'h507: dout <= 8'b00000000; // 1287 :   0 - 0x0
      13'h508: dout <= 8'b00000000; // 1288 :   0 - 0x0
      13'h509: dout <= 8'b00000000; // 1289 :   0 - 0x0
      13'h50A: dout <= 8'b00000000; // 1290 :   0 - 0x0
      13'h50B: dout <= 8'b00000000; // 1291 :   0 - 0x0
      13'h50C: dout <= 8'b00000000; // 1292 :   0 - 0x0
      13'h50D: dout <= 8'b00000000; // 1293 :   0 - 0x0
      13'h50E: dout <= 8'b00000000; // 1294 :   0 - 0x0
      13'h50F: dout <= 8'b00000000; // 1295 :   0 - 0x0
      13'h510: dout <= 8'b00111110; // 1296 :  62 - 0x3e -- Sprite 0x51
      13'h511: dout <= 8'b01100011; // 1297 :  99 - 0x63
      13'h512: dout <= 8'b01100011; // 1298 :  99 - 0x63
      13'h513: dout <= 8'b01100011; // 1299 :  99 - 0x63
      13'h514: dout <= 8'b01101111; // 1300 : 111 - 0x6f
      13'h515: dout <= 8'b01100110; // 1301 : 102 - 0x66
      13'h516: dout <= 8'b00111101; // 1302 :  61 - 0x3d
      13'h517: dout <= 8'b00000000; // 1303 :   0 - 0x0
      13'h518: dout <= 8'b00000000; // 1304 :   0 - 0x0
      13'h519: dout <= 8'b00000000; // 1305 :   0 - 0x0
      13'h51A: dout <= 8'b00000000; // 1306 :   0 - 0x0
      13'h51B: dout <= 8'b00000000; // 1307 :   0 - 0x0
      13'h51C: dout <= 8'b00000000; // 1308 :   0 - 0x0
      13'h51D: dout <= 8'b00000000; // 1309 :   0 - 0x0
      13'h51E: dout <= 8'b00000000; // 1310 :   0 - 0x0
      13'h51F: dout <= 8'b00000000; // 1311 :   0 - 0x0
      13'h520: dout <= 8'b01111110; // 1312 : 126 - 0x7e -- Sprite 0x52
      13'h521: dout <= 8'b01100011; // 1313 :  99 - 0x63
      13'h522: dout <= 8'b01100011; // 1314 :  99 - 0x63
      13'h523: dout <= 8'b01100111; // 1315 : 103 - 0x67
      13'h524: dout <= 8'b01111100; // 1316 : 124 - 0x7c
      13'h525: dout <= 8'b01101110; // 1317 : 110 - 0x6e
      13'h526: dout <= 8'b01100111; // 1318 : 103 - 0x67
      13'h527: dout <= 8'b00000000; // 1319 :   0 - 0x0
      13'h528: dout <= 8'b00000000; // 1320 :   0 - 0x0
      13'h529: dout <= 8'b00000000; // 1321 :   0 - 0x0
      13'h52A: dout <= 8'b00000000; // 1322 :   0 - 0x0
      13'h52B: dout <= 8'b00000000; // 1323 :   0 - 0x0
      13'h52C: dout <= 8'b00000000; // 1324 :   0 - 0x0
      13'h52D: dout <= 8'b00000000; // 1325 :   0 - 0x0
      13'h52E: dout <= 8'b00000000; // 1326 :   0 - 0x0
      13'h52F: dout <= 8'b00000000; // 1327 :   0 - 0x0
      13'h530: dout <= 8'b00111100; // 1328 :  60 - 0x3c -- Sprite 0x53
      13'h531: dout <= 8'b01100110; // 1329 : 102 - 0x66
      13'h532: dout <= 8'b01100000; // 1330 :  96 - 0x60
      13'h533: dout <= 8'b00111110; // 1331 :  62 - 0x3e
      13'h534: dout <= 8'b00000011; // 1332 :   3 - 0x3
      13'h535: dout <= 8'b01100011; // 1333 :  99 - 0x63
      13'h536: dout <= 8'b00111110; // 1334 :  62 - 0x3e
      13'h537: dout <= 8'b00000000; // 1335 :   0 - 0x0
      13'h538: dout <= 8'b00000000; // 1336 :   0 - 0x0
      13'h539: dout <= 8'b00000000; // 1337 :   0 - 0x0
      13'h53A: dout <= 8'b00000000; // 1338 :   0 - 0x0
      13'h53B: dout <= 8'b00000000; // 1339 :   0 - 0x0
      13'h53C: dout <= 8'b00000000; // 1340 :   0 - 0x0
      13'h53D: dout <= 8'b00000000; // 1341 :   0 - 0x0
      13'h53E: dout <= 8'b00000000; // 1342 :   0 - 0x0
      13'h53F: dout <= 8'b00000000; // 1343 :   0 - 0x0
      13'h540: dout <= 8'b00111111; // 1344 :  63 - 0x3f -- Sprite 0x54
      13'h541: dout <= 8'b00001100; // 1345 :  12 - 0xc
      13'h542: dout <= 8'b00001100; // 1346 :  12 - 0xc
      13'h543: dout <= 8'b00001100; // 1347 :  12 - 0xc
      13'h544: dout <= 8'b00001100; // 1348 :  12 - 0xc
      13'h545: dout <= 8'b00001100; // 1349 :  12 - 0xc
      13'h546: dout <= 8'b00001100; // 1350 :  12 - 0xc
      13'h547: dout <= 8'b00000000; // 1351 :   0 - 0x0
      13'h548: dout <= 8'b00000000; // 1352 :   0 - 0x0
      13'h549: dout <= 8'b00000000; // 1353 :   0 - 0x0
      13'h54A: dout <= 8'b00000000; // 1354 :   0 - 0x0
      13'h54B: dout <= 8'b00000000; // 1355 :   0 - 0x0
      13'h54C: dout <= 8'b00000000; // 1356 :   0 - 0x0
      13'h54D: dout <= 8'b00000000; // 1357 :   0 - 0x0
      13'h54E: dout <= 8'b00000000; // 1358 :   0 - 0x0
      13'h54F: dout <= 8'b00000000; // 1359 :   0 - 0x0
      13'h550: dout <= 8'b01100011; // 1360 :  99 - 0x63 -- Sprite 0x55
      13'h551: dout <= 8'b01100011; // 1361 :  99 - 0x63
      13'h552: dout <= 8'b01100011; // 1362 :  99 - 0x63
      13'h553: dout <= 8'b01100011; // 1363 :  99 - 0x63
      13'h554: dout <= 8'b01100011; // 1364 :  99 - 0x63
      13'h555: dout <= 8'b01100011; // 1365 :  99 - 0x63
      13'h556: dout <= 8'b00111110; // 1366 :  62 - 0x3e
      13'h557: dout <= 8'b00000000; // 1367 :   0 - 0x0
      13'h558: dout <= 8'b00000000; // 1368 :   0 - 0x0
      13'h559: dout <= 8'b00000000; // 1369 :   0 - 0x0
      13'h55A: dout <= 8'b00000000; // 1370 :   0 - 0x0
      13'h55B: dout <= 8'b00000000; // 1371 :   0 - 0x0
      13'h55C: dout <= 8'b00000000; // 1372 :   0 - 0x0
      13'h55D: dout <= 8'b00000000; // 1373 :   0 - 0x0
      13'h55E: dout <= 8'b00000000; // 1374 :   0 - 0x0
      13'h55F: dout <= 8'b00000000; // 1375 :   0 - 0x0
      13'h560: dout <= 8'b01100011; // 1376 :  99 - 0x63 -- Sprite 0x56
      13'h561: dout <= 8'b01100011; // 1377 :  99 - 0x63
      13'h562: dout <= 8'b01100011; // 1378 :  99 - 0x63
      13'h563: dout <= 8'b01110111; // 1379 : 119 - 0x77
      13'h564: dout <= 8'b00111110; // 1380 :  62 - 0x3e
      13'h565: dout <= 8'b00011100; // 1381 :  28 - 0x1c
      13'h566: dout <= 8'b00001000; // 1382 :   8 - 0x8
      13'h567: dout <= 8'b00000000; // 1383 :   0 - 0x0
      13'h568: dout <= 8'b00000000; // 1384 :   0 - 0x0
      13'h569: dout <= 8'b00000000; // 1385 :   0 - 0x0
      13'h56A: dout <= 8'b00000000; // 1386 :   0 - 0x0
      13'h56B: dout <= 8'b00000000; // 1387 :   0 - 0x0
      13'h56C: dout <= 8'b00000000; // 1388 :   0 - 0x0
      13'h56D: dout <= 8'b00000000; // 1389 :   0 - 0x0
      13'h56E: dout <= 8'b00000000; // 1390 :   0 - 0x0
      13'h56F: dout <= 8'b00000000; // 1391 :   0 - 0x0
      13'h570: dout <= 8'b01100011; // 1392 :  99 - 0x63 -- Sprite 0x57
      13'h571: dout <= 8'b01100011; // 1393 :  99 - 0x63
      13'h572: dout <= 8'b01101011; // 1394 : 107 - 0x6b
      13'h573: dout <= 8'b01111111; // 1395 : 127 - 0x7f
      13'h574: dout <= 8'b01111111; // 1396 : 127 - 0x7f
      13'h575: dout <= 8'b01110111; // 1397 : 119 - 0x77
      13'h576: dout <= 8'b01100011; // 1398 :  99 - 0x63
      13'h577: dout <= 8'b00000000; // 1399 :   0 - 0x0
      13'h578: dout <= 8'b00000000; // 1400 :   0 - 0x0
      13'h579: dout <= 8'b00000000; // 1401 :   0 - 0x0
      13'h57A: dout <= 8'b00000000; // 1402 :   0 - 0x0
      13'h57B: dout <= 8'b00000000; // 1403 :   0 - 0x0
      13'h57C: dout <= 8'b00000000; // 1404 :   0 - 0x0
      13'h57D: dout <= 8'b00000000; // 1405 :   0 - 0x0
      13'h57E: dout <= 8'b00000000; // 1406 :   0 - 0x0
      13'h57F: dout <= 8'b00000000; // 1407 :   0 - 0x0
      13'h580: dout <= 8'b01100011; // 1408 :  99 - 0x63 -- Sprite 0x58
      13'h581: dout <= 8'b01110111; // 1409 : 119 - 0x77
      13'h582: dout <= 8'b00111110; // 1410 :  62 - 0x3e
      13'h583: dout <= 8'b00011100; // 1411 :  28 - 0x1c
      13'h584: dout <= 8'b00111110; // 1412 :  62 - 0x3e
      13'h585: dout <= 8'b01110111; // 1413 : 119 - 0x77
      13'h586: dout <= 8'b01100011; // 1414 :  99 - 0x63
      13'h587: dout <= 8'b00000000; // 1415 :   0 - 0x0
      13'h588: dout <= 8'b00000000; // 1416 :   0 - 0x0
      13'h589: dout <= 8'b00000000; // 1417 :   0 - 0x0
      13'h58A: dout <= 8'b00000000; // 1418 :   0 - 0x0
      13'h58B: dout <= 8'b00000000; // 1419 :   0 - 0x0
      13'h58C: dout <= 8'b00000000; // 1420 :   0 - 0x0
      13'h58D: dout <= 8'b00000000; // 1421 :   0 - 0x0
      13'h58E: dout <= 8'b00000000; // 1422 :   0 - 0x0
      13'h58F: dout <= 8'b00000000; // 1423 :   0 - 0x0
      13'h590: dout <= 8'b00110011; // 1424 :  51 - 0x33 -- Sprite 0x59
      13'h591: dout <= 8'b00110011; // 1425 :  51 - 0x33
      13'h592: dout <= 8'b00110011; // 1426 :  51 - 0x33
      13'h593: dout <= 8'b00011110; // 1427 :  30 - 0x1e
      13'h594: dout <= 8'b00001100; // 1428 :  12 - 0xc
      13'h595: dout <= 8'b00001100; // 1429 :  12 - 0xc
      13'h596: dout <= 8'b00001100; // 1430 :  12 - 0xc
      13'h597: dout <= 8'b00000000; // 1431 :   0 - 0x0
      13'h598: dout <= 8'b00000000; // 1432 :   0 - 0x0
      13'h599: dout <= 8'b00000000; // 1433 :   0 - 0x0
      13'h59A: dout <= 8'b00000000; // 1434 :   0 - 0x0
      13'h59B: dout <= 8'b00000000; // 1435 :   0 - 0x0
      13'h59C: dout <= 8'b00000000; // 1436 :   0 - 0x0
      13'h59D: dout <= 8'b00000000; // 1437 :   0 - 0x0
      13'h59E: dout <= 8'b00000000; // 1438 :   0 - 0x0
      13'h59F: dout <= 8'b00000000; // 1439 :   0 - 0x0
      13'h5A0: dout <= 8'b01111111; // 1440 : 127 - 0x7f -- Sprite 0x5a
      13'h5A1: dout <= 8'b00000111; // 1441 :   7 - 0x7
      13'h5A2: dout <= 8'b00001110; // 1442 :  14 - 0xe
      13'h5A3: dout <= 8'b00011100; // 1443 :  28 - 0x1c
      13'h5A4: dout <= 8'b00111000; // 1444 :  56 - 0x38
      13'h5A5: dout <= 8'b01110000; // 1445 : 112 - 0x70
      13'h5A6: dout <= 8'b01111111; // 1446 : 127 - 0x7f
      13'h5A7: dout <= 8'b00000000; // 1447 :   0 - 0x0
      13'h5A8: dout <= 8'b00000000; // 1448 :   0 - 0x0
      13'h5A9: dout <= 8'b00000000; // 1449 :   0 - 0x0
      13'h5AA: dout <= 8'b00000000; // 1450 :   0 - 0x0
      13'h5AB: dout <= 8'b00000000; // 1451 :   0 - 0x0
      13'h5AC: dout <= 8'b00000000; // 1452 :   0 - 0x0
      13'h5AD: dout <= 8'b00000000; // 1453 :   0 - 0x0
      13'h5AE: dout <= 8'b00000000; // 1454 :   0 - 0x0
      13'h5AF: dout <= 8'b00000000; // 1455 :   0 - 0x0
      13'h5B0: dout <= 8'b00000000; // 1456 :   0 - 0x0 -- Sprite 0x5b
      13'h5B1: dout <= 8'b00000000; // 1457 :   0 - 0x0
      13'h5B2: dout <= 8'b00000000; // 1458 :   0 - 0x0
      13'h5B3: dout <= 8'b00000000; // 1459 :   0 - 0x0
      13'h5B4: dout <= 8'b00000000; // 1460 :   0 - 0x0
      13'h5B5: dout <= 8'b00110000; // 1461 :  48 - 0x30
      13'h5B6: dout <= 8'b00110000; // 1462 :  48 - 0x30
      13'h5B7: dout <= 8'b00000000; // 1463 :   0 - 0x0
      13'h5B8: dout <= 8'b00000000; // 1464 :   0 - 0x0
      13'h5B9: dout <= 8'b00000000; // 1465 :   0 - 0x0
      13'h5BA: dout <= 8'b00000000; // 1466 :   0 - 0x0
      13'h5BB: dout <= 8'b00000000; // 1467 :   0 - 0x0
      13'h5BC: dout <= 8'b00000000; // 1468 :   0 - 0x0
      13'h5BD: dout <= 8'b00000000; // 1469 :   0 - 0x0
      13'h5BE: dout <= 8'b00000000; // 1470 :   0 - 0x0
      13'h5BF: dout <= 8'b00000000; // 1471 :   0 - 0x0
      13'h5C0: dout <= 8'b11000000; // 1472 : 192 - 0xc0 -- Sprite 0x5c
      13'h5C1: dout <= 8'b11110000; // 1473 : 240 - 0xf0
      13'h5C2: dout <= 8'b11111100; // 1474 : 252 - 0xfc
      13'h5C3: dout <= 8'b11111111; // 1475 : 255 - 0xff
      13'h5C4: dout <= 8'b11111100; // 1476 : 252 - 0xfc
      13'h5C5: dout <= 8'b11110000; // 1477 : 240 - 0xf0
      13'h5C6: dout <= 8'b11000000; // 1478 : 192 - 0xc0
      13'h5C7: dout <= 8'b00000000; // 1479 :   0 - 0x0
      13'h5C8: dout <= 8'b00000000; // 1480 :   0 - 0x0
      13'h5C9: dout <= 8'b00000000; // 1481 :   0 - 0x0
      13'h5CA: dout <= 8'b00000000; // 1482 :   0 - 0x0
      13'h5CB: dout <= 8'b00000000; // 1483 :   0 - 0x0
      13'h5CC: dout <= 8'b00000000; // 1484 :   0 - 0x0
      13'h5CD: dout <= 8'b00000000; // 1485 :   0 - 0x0
      13'h5CE: dout <= 8'b00000000; // 1486 :   0 - 0x0
      13'h5CF: dout <= 8'b00000000; // 1487 :   0 - 0x0
      13'h5D0: dout <= 8'b00111100; // 1488 :  60 - 0x3c -- Sprite 0x5d
      13'h5D1: dout <= 8'b01000010; // 1489 :  66 - 0x42
      13'h5D2: dout <= 8'b10011001; // 1490 : 153 - 0x99
      13'h5D3: dout <= 8'b10100001; // 1491 : 161 - 0xa1
      13'h5D4: dout <= 8'b10100001; // 1492 : 161 - 0xa1
      13'h5D5: dout <= 8'b10011001; // 1493 : 153 - 0x99
      13'h5D6: dout <= 8'b01000010; // 1494 :  66 - 0x42
      13'h5D7: dout <= 8'b00111100; // 1495 :  60 - 0x3c
      13'h5D8: dout <= 8'b00000000; // 1496 :   0 - 0x0
      13'h5D9: dout <= 8'b00000000; // 1497 :   0 - 0x0
      13'h5DA: dout <= 8'b00000000; // 1498 :   0 - 0x0
      13'h5DB: dout <= 8'b00000000; // 1499 :   0 - 0x0
      13'h5DC: dout <= 8'b00000000; // 1500 :   0 - 0x0
      13'h5DD: dout <= 8'b00000000; // 1501 :   0 - 0x0
      13'h5DE: dout <= 8'b00000000; // 1502 :   0 - 0x0
      13'h5DF: dout <= 8'b00000000; // 1503 :   0 - 0x0
      13'h5E0: dout <= 8'b00000000; // 1504 :   0 - 0x0 -- Sprite 0x5e
      13'h5E1: dout <= 8'b00000000; // 1505 :   0 - 0x0
      13'h5E2: dout <= 8'b00010000; // 1506 :  16 - 0x10
      13'h5E3: dout <= 8'b00010000; // 1507 :  16 - 0x10
      13'h5E4: dout <= 8'b00010000; // 1508 :  16 - 0x10
      13'h5E5: dout <= 8'b00010000; // 1509 :  16 - 0x10
      13'h5E6: dout <= 8'b00000000; // 1510 :   0 - 0x0
      13'h5E7: dout <= 8'b00000000; // 1511 :   0 - 0x0
      13'h5E8: dout <= 8'b00000000; // 1512 :   0 - 0x0
      13'h5E9: dout <= 8'b00000000; // 1513 :   0 - 0x0
      13'h5EA: dout <= 8'b00010000; // 1514 :  16 - 0x10
      13'h5EB: dout <= 8'b00010000; // 1515 :  16 - 0x10
      13'h5EC: dout <= 8'b00010000; // 1516 :  16 - 0x10
      13'h5ED: dout <= 8'b00010000; // 1517 :  16 - 0x10
      13'h5EE: dout <= 8'b00000000; // 1518 :   0 - 0x0
      13'h5EF: dout <= 8'b00000000; // 1519 :   0 - 0x0
      13'h5F0: dout <= 8'b00110110; // 1520 :  54 - 0x36 -- Sprite 0x5f
      13'h5F1: dout <= 8'b00110110; // 1521 :  54 - 0x36
      13'h5F2: dout <= 8'b00010010; // 1522 :  18 - 0x12
      13'h5F3: dout <= 8'b00000000; // 1523 :   0 - 0x0
      13'h5F4: dout <= 8'b00000000; // 1524 :   0 - 0x0
      13'h5F5: dout <= 8'b00000000; // 1525 :   0 - 0x0
      13'h5F6: dout <= 8'b00000000; // 1526 :   0 - 0x0
      13'h5F7: dout <= 8'b00000000; // 1527 :   0 - 0x0
      13'h5F8: dout <= 8'b00000000; // 1528 :   0 - 0x0
      13'h5F9: dout <= 8'b00000000; // 1529 :   0 - 0x0
      13'h5FA: dout <= 8'b00000000; // 1530 :   0 - 0x0
      13'h5FB: dout <= 8'b00000000; // 1531 :   0 - 0x0
      13'h5FC: dout <= 8'b00000000; // 1532 :   0 - 0x0
      13'h5FD: dout <= 8'b00000000; // 1533 :   0 - 0x0
      13'h5FE: dout <= 8'b00000000; // 1534 :   0 - 0x0
      13'h5FF: dout <= 8'b00000000; // 1535 :   0 - 0x0
      13'h600: dout <= 8'b00000000; // 1536 :   0 - 0x0 -- Sprite 0x60
      13'h601: dout <= 8'b00000000; // 1537 :   0 - 0x0
      13'h602: dout <= 8'b00000000; // 1538 :   0 - 0x0
      13'h603: dout <= 8'b00000000; // 1539 :   0 - 0x0
      13'h604: dout <= 8'b00000000; // 1540 :   0 - 0x0
      13'h605: dout <= 8'b00000001; // 1541 :   1 - 0x1
      13'h606: dout <= 8'b00011110; // 1542 :  30 - 0x1e
      13'h607: dout <= 8'b00111011; // 1543 :  59 - 0x3b
      13'h608: dout <= 8'b00000000; // 1544 :   0 - 0x0
      13'h609: dout <= 8'b00000000; // 1545 :   0 - 0x0
      13'h60A: dout <= 8'b00000000; // 1546 :   0 - 0x0
      13'h60B: dout <= 8'b00000000; // 1547 :   0 - 0x0
      13'h60C: dout <= 8'b00000000; // 1548 :   0 - 0x0
      13'h60D: dout <= 8'b00000000; // 1549 :   0 - 0x0
      13'h60E: dout <= 8'b00000000; // 1550 :   0 - 0x0
      13'h60F: dout <= 8'b00000000; // 1551 :   0 - 0x0
      13'h610: dout <= 8'b00000000; // 1552 :   0 - 0x0 -- Sprite 0x61
      13'h611: dout <= 8'b00000000; // 1553 :   0 - 0x0
      13'h612: dout <= 8'b00001100; // 1554 :  12 - 0xc
      13'h613: dout <= 8'b00111100; // 1555 :  60 - 0x3c
      13'h614: dout <= 8'b11010000; // 1556 : 208 - 0xd0
      13'h615: dout <= 8'b00010000; // 1557 :  16 - 0x10
      13'h616: dout <= 8'b00100000; // 1558 :  32 - 0x20
      13'h617: dout <= 8'b01000000; // 1559 :  64 - 0x40
      13'h618: dout <= 8'b00000000; // 1560 :   0 - 0x0
      13'h619: dout <= 8'b00000000; // 1561 :   0 - 0x0
      13'h61A: dout <= 8'b00000000; // 1562 :   0 - 0x0
      13'h61B: dout <= 8'b00000000; // 1563 :   0 - 0x0
      13'h61C: dout <= 8'b00000000; // 1564 :   0 - 0x0
      13'h61D: dout <= 8'b00000000; // 1565 :   0 - 0x0
      13'h61E: dout <= 8'b00000000; // 1566 :   0 - 0x0
      13'h61F: dout <= 8'b00000000; // 1567 :   0 - 0x0
      13'h620: dout <= 8'b00111110; // 1568 :  62 - 0x3e -- Sprite 0x62
      13'h621: dout <= 8'b00101101; // 1569 :  45 - 0x2d
      13'h622: dout <= 8'b00110101; // 1570 :  53 - 0x35
      13'h623: dout <= 8'b00011101; // 1571 :  29 - 0x1d
      13'h624: dout <= 8'b00000001; // 1572 :   1 - 0x1
      13'h625: dout <= 8'b00000000; // 1573 :   0 - 0x0
      13'h626: dout <= 8'b00000000; // 1574 :   0 - 0x0
      13'h627: dout <= 8'b00000000; // 1575 :   0 - 0x0
      13'h628: dout <= 8'b00000000; // 1576 :   0 - 0x0
      13'h629: dout <= 8'b00000000; // 1577 :   0 - 0x0
      13'h62A: dout <= 8'b00000000; // 1578 :   0 - 0x0
      13'h62B: dout <= 8'b00000000; // 1579 :   0 - 0x0
      13'h62C: dout <= 8'b00000000; // 1580 :   0 - 0x0
      13'h62D: dout <= 8'b00000000; // 1581 :   0 - 0x0
      13'h62E: dout <= 8'b00000000; // 1582 :   0 - 0x0
      13'h62F: dout <= 8'b00000000; // 1583 :   0 - 0x0
      13'h630: dout <= 8'b10110000; // 1584 : 176 - 0xb0 -- Sprite 0x63
      13'h631: dout <= 8'b10111000; // 1585 : 184 - 0xb8
      13'h632: dout <= 8'b11111000; // 1586 : 248 - 0xf8
      13'h633: dout <= 8'b01111000; // 1587 : 120 - 0x78
      13'h634: dout <= 8'b10011000; // 1588 : 152 - 0x98
      13'h635: dout <= 8'b11110000; // 1589 : 240 - 0xf0
      13'h636: dout <= 8'b00000000; // 1590 :   0 - 0x0
      13'h637: dout <= 8'b00000000; // 1591 :   0 - 0x0
      13'h638: dout <= 8'b00000000; // 1592 :   0 - 0x0
      13'h639: dout <= 8'b00000000; // 1593 :   0 - 0x0
      13'h63A: dout <= 8'b00000000; // 1594 :   0 - 0x0
      13'h63B: dout <= 8'b00000000; // 1595 :   0 - 0x0
      13'h63C: dout <= 8'b00000000; // 1596 :   0 - 0x0
      13'h63D: dout <= 8'b00000000; // 1597 :   0 - 0x0
      13'h63E: dout <= 8'b00000000; // 1598 :   0 - 0x0
      13'h63F: dout <= 8'b00000000; // 1599 :   0 - 0x0
      13'h640: dout <= 8'b00000000; // 1600 :   0 - 0x0 -- Sprite 0x64
      13'h641: dout <= 8'b00000000; // 1601 :   0 - 0x0
      13'h642: dout <= 8'b00000111; // 1602 :   7 - 0x7
      13'h643: dout <= 8'b00000011; // 1603 :   3 - 0x3
      13'h644: dout <= 8'b00001101; // 1604 :  13 - 0xd
      13'h645: dout <= 8'b00011110; // 1605 :  30 - 0x1e
      13'h646: dout <= 8'b00010111; // 1606 :  23 - 0x17
      13'h647: dout <= 8'b00011101; // 1607 :  29 - 0x1d
      13'h648: dout <= 8'b00000000; // 1608 :   0 - 0x0
      13'h649: dout <= 8'b00000000; // 1609 :   0 - 0x0
      13'h64A: dout <= 8'b00000000; // 1610 :   0 - 0x0
      13'h64B: dout <= 8'b00000000; // 1611 :   0 - 0x0
      13'h64C: dout <= 8'b00000000; // 1612 :   0 - 0x0
      13'h64D: dout <= 8'b00000000; // 1613 :   0 - 0x0
      13'h64E: dout <= 8'b00000000; // 1614 :   0 - 0x0
      13'h64F: dout <= 8'b00000000; // 1615 :   0 - 0x0
      13'h650: dout <= 8'b00000000; // 1616 :   0 - 0x0 -- Sprite 0x65
      13'h651: dout <= 8'b10000000; // 1617 : 128 - 0x80
      13'h652: dout <= 8'b01110000; // 1618 : 112 - 0x70
      13'h653: dout <= 8'b11100000; // 1619 : 224 - 0xe0
      13'h654: dout <= 8'b11011000; // 1620 : 216 - 0xd8
      13'h655: dout <= 8'b10111100; // 1621 : 188 - 0xbc
      13'h656: dout <= 8'b01110100; // 1622 : 116 - 0x74
      13'h657: dout <= 8'b11011100; // 1623 : 220 - 0xdc
      13'h658: dout <= 8'b00000000; // 1624 :   0 - 0x0
      13'h659: dout <= 8'b00000000; // 1625 :   0 - 0x0
      13'h65A: dout <= 8'b00000000; // 1626 :   0 - 0x0
      13'h65B: dout <= 8'b00000000; // 1627 :   0 - 0x0
      13'h65C: dout <= 8'b00000000; // 1628 :   0 - 0x0
      13'h65D: dout <= 8'b00000000; // 1629 :   0 - 0x0
      13'h65E: dout <= 8'b00000000; // 1630 :   0 - 0x0
      13'h65F: dout <= 8'b00000000; // 1631 :   0 - 0x0
      13'h660: dout <= 8'b00011111; // 1632 :  31 - 0x1f -- Sprite 0x66
      13'h661: dout <= 8'b00001011; // 1633 :  11 - 0xb
      13'h662: dout <= 8'b00001111; // 1634 :  15 - 0xf
      13'h663: dout <= 8'b00000101; // 1635 :   5 - 0x5
      13'h664: dout <= 8'b00000011; // 1636 :   3 - 0x3
      13'h665: dout <= 8'b00000001; // 1637 :   1 - 0x1
      13'h666: dout <= 8'b00000000; // 1638 :   0 - 0x0
      13'h667: dout <= 8'b00000000; // 1639 :   0 - 0x0
      13'h668: dout <= 8'b00000000; // 1640 :   0 - 0x0
      13'h669: dout <= 8'b00000000; // 1641 :   0 - 0x0
      13'h66A: dout <= 8'b00000000; // 1642 :   0 - 0x0
      13'h66B: dout <= 8'b00000000; // 1643 :   0 - 0x0
      13'h66C: dout <= 8'b00000000; // 1644 :   0 - 0x0
      13'h66D: dout <= 8'b00000000; // 1645 :   0 - 0x0
      13'h66E: dout <= 8'b00000000; // 1646 :   0 - 0x0
      13'h66F: dout <= 8'b00000000; // 1647 :   0 - 0x0
      13'h670: dout <= 8'b11111100; // 1648 : 252 - 0xfc -- Sprite 0x67
      13'h671: dout <= 8'b01101000; // 1649 : 104 - 0x68
      13'h672: dout <= 8'b11111000; // 1650 : 248 - 0xf8
      13'h673: dout <= 8'b10110000; // 1651 : 176 - 0xb0
      13'h674: dout <= 8'b11100000; // 1652 : 224 - 0xe0
      13'h675: dout <= 8'b10000000; // 1653 : 128 - 0x80
      13'h676: dout <= 8'b00000000; // 1654 :   0 - 0x0
      13'h677: dout <= 8'b00000000; // 1655 :   0 - 0x0
      13'h678: dout <= 8'b00000000; // 1656 :   0 - 0x0
      13'h679: dout <= 8'b00000000; // 1657 :   0 - 0x0
      13'h67A: dout <= 8'b00000000; // 1658 :   0 - 0x0
      13'h67B: dout <= 8'b00000000; // 1659 :   0 - 0x0
      13'h67C: dout <= 8'b00000000; // 1660 :   0 - 0x0
      13'h67D: dout <= 8'b00000000; // 1661 :   0 - 0x0
      13'h67E: dout <= 8'b00000000; // 1662 :   0 - 0x0
      13'h67F: dout <= 8'b00000000; // 1663 :   0 - 0x0
      13'h680: dout <= 8'b00000000; // 1664 :   0 - 0x0 -- Sprite 0x68
      13'h681: dout <= 8'b00000000; // 1665 :   0 - 0x0
      13'h682: dout <= 8'b00000000; // 1666 :   0 - 0x0
      13'h683: dout <= 8'b00000000; // 1667 :   0 - 0x0
      13'h684: dout <= 8'b00000000; // 1668 :   0 - 0x0
      13'h685: dout <= 8'b00000000; // 1669 :   0 - 0x0
      13'h686: dout <= 8'b00000000; // 1670 :   0 - 0x0
      13'h687: dout <= 8'b00000000; // 1671 :   0 - 0x0
      13'h688: dout <= 8'b00000000; // 1672 :   0 - 0x0
      13'h689: dout <= 8'b00000000; // 1673 :   0 - 0x0
      13'h68A: dout <= 8'b00000000; // 1674 :   0 - 0x0
      13'h68B: dout <= 8'b00000001; // 1675 :   1 - 0x1
      13'h68C: dout <= 8'b00000001; // 1676 :   1 - 0x1
      13'h68D: dout <= 8'b00001011; // 1677 :  11 - 0xb
      13'h68E: dout <= 8'b00011100; // 1678 :  28 - 0x1c
      13'h68F: dout <= 8'b00111111; // 1679 :  63 - 0x3f
      13'h690: dout <= 8'b00000000; // 1680 :   0 - 0x0 -- Sprite 0x69
      13'h691: dout <= 8'b00000000; // 1681 :   0 - 0x0
      13'h692: dout <= 8'b00000000; // 1682 :   0 - 0x0
      13'h693: dout <= 8'b00000000; // 1683 :   0 - 0x0
      13'h694: dout <= 8'b00000000; // 1684 :   0 - 0x0
      13'h695: dout <= 8'b00000000; // 1685 :   0 - 0x0
      13'h696: dout <= 8'b00000000; // 1686 :   0 - 0x0
      13'h697: dout <= 8'b00000000; // 1687 :   0 - 0x0
      13'h698: dout <= 8'b00000000; // 1688 :   0 - 0x0
      13'h699: dout <= 8'b00000000; // 1689 :   0 - 0x0
      13'h69A: dout <= 8'b00110000; // 1690 :  48 - 0x30
      13'h69B: dout <= 8'b01111000; // 1691 : 120 - 0x78
      13'h69C: dout <= 8'b10000000; // 1692 : 128 - 0x80
      13'h69D: dout <= 8'b11110000; // 1693 : 240 - 0xf0
      13'h69E: dout <= 8'b11111000; // 1694 : 248 - 0xf8
      13'h69F: dout <= 8'b11111100; // 1695 : 252 - 0xfc
      13'h6A0: dout <= 8'b00000000; // 1696 :   0 - 0x0 -- Sprite 0x6a
      13'h6A1: dout <= 8'b00000000; // 1697 :   0 - 0x0
      13'h6A2: dout <= 8'b00000000; // 1698 :   0 - 0x0
      13'h6A3: dout <= 8'b00000000; // 1699 :   0 - 0x0
      13'h6A4: dout <= 8'b00000000; // 1700 :   0 - 0x0
      13'h6A5: dout <= 8'b00000000; // 1701 :   0 - 0x0
      13'h6A6: dout <= 8'b00000000; // 1702 :   0 - 0x0
      13'h6A7: dout <= 8'b00000000; // 1703 :   0 - 0x0
      13'h6A8: dout <= 8'b00111111; // 1704 :  63 - 0x3f
      13'h6A9: dout <= 8'b00111111; // 1705 :  63 - 0x3f
      13'h6AA: dout <= 8'b00111111; // 1706 :  63 - 0x3f
      13'h6AB: dout <= 8'b00011111; // 1707 :  31 - 0x1f
      13'h6AC: dout <= 8'b00011111; // 1708 :  31 - 0x1f
      13'h6AD: dout <= 8'b00000111; // 1709 :   7 - 0x7
      13'h6AE: dout <= 8'b00000000; // 1710 :   0 - 0x0
      13'h6AF: dout <= 8'b00000000; // 1711 :   0 - 0x0
      13'h6B0: dout <= 8'b00000000; // 1712 :   0 - 0x0 -- Sprite 0x6b
      13'h6B1: dout <= 8'b00000000; // 1713 :   0 - 0x0
      13'h6B2: dout <= 8'b00000000; // 1714 :   0 - 0x0
      13'h6B3: dout <= 8'b00000000; // 1715 :   0 - 0x0
      13'h6B4: dout <= 8'b00000000; // 1716 :   0 - 0x0
      13'h6B5: dout <= 8'b00000000; // 1717 :   0 - 0x0
      13'h6B6: dout <= 8'b00000000; // 1718 :   0 - 0x0
      13'h6B7: dout <= 8'b00000000; // 1719 :   0 - 0x0
      13'h6B8: dout <= 8'b11111100; // 1720 : 252 - 0xfc
      13'h6B9: dout <= 8'b11101100; // 1721 : 236 - 0xec
      13'h6BA: dout <= 8'b11101100; // 1722 : 236 - 0xec
      13'h6BB: dout <= 8'b11011000; // 1723 : 216 - 0xd8
      13'h6BC: dout <= 8'b11111000; // 1724 : 248 - 0xf8
      13'h6BD: dout <= 8'b11100000; // 1725 : 224 - 0xe0
      13'h6BE: dout <= 8'b00000000; // 1726 :   0 - 0x0
      13'h6BF: dout <= 8'b00000000; // 1727 :   0 - 0x0
      13'h6C0: dout <= 8'b00000000; // 1728 :   0 - 0x0 -- Sprite 0x6c
      13'h6C1: dout <= 8'b00000000; // 1729 :   0 - 0x0
      13'h6C2: dout <= 8'b00000001; // 1730 :   1 - 0x1
      13'h6C3: dout <= 8'b00011101; // 1731 :  29 - 0x1d
      13'h6C4: dout <= 8'b00111110; // 1732 :  62 - 0x3e
      13'h6C5: dout <= 8'b00111111; // 1733 :  63 - 0x3f
      13'h6C6: dout <= 8'b00111111; // 1734 :  63 - 0x3f
      13'h6C7: dout <= 8'b00111111; // 1735 :  63 - 0x3f
      13'h6C8: dout <= 8'b00000000; // 1736 :   0 - 0x0
      13'h6C9: dout <= 8'b00000000; // 1737 :   0 - 0x0
      13'h6CA: dout <= 8'b00000001; // 1738 :   1 - 0x1
      13'h6CB: dout <= 8'b00011101; // 1739 :  29 - 0x1d
      13'h6CC: dout <= 8'b00111110; // 1740 :  62 - 0x3e
      13'h6CD: dout <= 8'b00111111; // 1741 :  63 - 0x3f
      13'h6CE: dout <= 8'b00111111; // 1742 :  63 - 0x3f
      13'h6CF: dout <= 8'b00111111; // 1743 :  63 - 0x3f
      13'h6D0: dout <= 8'b00000000; // 1744 :   0 - 0x0 -- Sprite 0x6d
      13'h6D1: dout <= 8'b10000000; // 1745 : 128 - 0x80
      13'h6D2: dout <= 8'b00000000; // 1746 :   0 - 0x0
      13'h6D3: dout <= 8'b01110000; // 1747 : 112 - 0x70
      13'h6D4: dout <= 8'b11111000; // 1748 : 248 - 0xf8
      13'h6D5: dout <= 8'b11111100; // 1749 : 252 - 0xfc
      13'h6D6: dout <= 8'b11111100; // 1750 : 252 - 0xfc
      13'h6D7: dout <= 8'b11111100; // 1751 : 252 - 0xfc
      13'h6D8: dout <= 8'b00000000; // 1752 :   0 - 0x0
      13'h6D9: dout <= 8'b10000000; // 1753 : 128 - 0x80
      13'h6DA: dout <= 8'b00000000; // 1754 :   0 - 0x0
      13'h6DB: dout <= 8'b01110000; // 1755 : 112 - 0x70
      13'h6DC: dout <= 8'b11111000; // 1756 : 248 - 0xf8
      13'h6DD: dout <= 8'b11111100; // 1757 : 252 - 0xfc
      13'h6DE: dout <= 8'b11111100; // 1758 : 252 - 0xfc
      13'h6DF: dout <= 8'b11111100; // 1759 : 252 - 0xfc
      13'h6E0: dout <= 8'b00111111; // 1760 :  63 - 0x3f -- Sprite 0x6e
      13'h6E1: dout <= 8'b00111111; // 1761 :  63 - 0x3f
      13'h6E2: dout <= 8'b00011111; // 1762 :  31 - 0x1f
      13'h6E3: dout <= 8'b00011111; // 1763 :  31 - 0x1f
      13'h6E4: dout <= 8'b00001111; // 1764 :  15 - 0xf
      13'h6E5: dout <= 8'b00000110; // 1765 :   6 - 0x6
      13'h6E6: dout <= 8'b00000000; // 1766 :   0 - 0x0
      13'h6E7: dout <= 8'b00000000; // 1767 :   0 - 0x0
      13'h6E8: dout <= 8'b00111111; // 1768 :  63 - 0x3f
      13'h6E9: dout <= 8'b00111111; // 1769 :  63 - 0x3f
      13'h6EA: dout <= 8'b00011111; // 1770 :  31 - 0x1f
      13'h6EB: dout <= 8'b00011111; // 1771 :  31 - 0x1f
      13'h6EC: dout <= 8'b00001111; // 1772 :  15 - 0xf
      13'h6ED: dout <= 8'b00000110; // 1773 :   6 - 0x6
      13'h6EE: dout <= 8'b00000000; // 1774 :   0 - 0x0
      13'h6EF: dout <= 8'b00000000; // 1775 :   0 - 0x0
      13'h6F0: dout <= 8'b11101100; // 1776 : 236 - 0xec -- Sprite 0x6f
      13'h6F1: dout <= 8'b11101100; // 1777 : 236 - 0xec
      13'h6F2: dout <= 8'b11011000; // 1778 : 216 - 0xd8
      13'h6F3: dout <= 8'b11111000; // 1779 : 248 - 0xf8
      13'h6F4: dout <= 8'b11110000; // 1780 : 240 - 0xf0
      13'h6F5: dout <= 8'b11100000; // 1781 : 224 - 0xe0
      13'h6F6: dout <= 8'b00000000; // 1782 :   0 - 0x0
      13'h6F7: dout <= 8'b00000000; // 1783 :   0 - 0x0
      13'h6F8: dout <= 8'b11101100; // 1784 : 236 - 0xec
      13'h6F9: dout <= 8'b11101100; // 1785 : 236 - 0xec
      13'h6FA: dout <= 8'b11011000; // 1786 : 216 - 0xd8
      13'h6FB: dout <= 8'b11111000; // 1787 : 248 - 0xf8
      13'h6FC: dout <= 8'b11110000; // 1788 : 240 - 0xf0
      13'h6FD: dout <= 8'b11100000; // 1789 : 224 - 0xe0
      13'h6FE: dout <= 8'b00000000; // 1790 :   0 - 0x0
      13'h6FF: dout <= 8'b00000000; // 1791 :   0 - 0x0
      13'h700: dout <= 8'b00000000; // 1792 :   0 - 0x0 -- Sprite 0x70
      13'h701: dout <= 8'b00000100; // 1793 :   4 - 0x4
      13'h702: dout <= 8'b00000011; // 1794 :   3 - 0x3
      13'h703: dout <= 8'b00000000; // 1795 :   0 - 0x0
      13'h704: dout <= 8'b00000001; // 1796 :   1 - 0x1
      13'h705: dout <= 8'b00000111; // 1797 :   7 - 0x7
      13'h706: dout <= 8'b00001111; // 1798 :  15 - 0xf
      13'h707: dout <= 8'b00001100; // 1799 :  12 - 0xc
      13'h708: dout <= 8'b00000000; // 1800 :   0 - 0x0
      13'h709: dout <= 8'b00000000; // 1801 :   0 - 0x0
      13'h70A: dout <= 8'b00000000; // 1802 :   0 - 0x0
      13'h70B: dout <= 8'b00000000; // 1803 :   0 - 0x0
      13'h70C: dout <= 8'b00000000; // 1804 :   0 - 0x0
      13'h70D: dout <= 8'b00000000; // 1805 :   0 - 0x0
      13'h70E: dout <= 8'b00000000; // 1806 :   0 - 0x0
      13'h70F: dout <= 8'b00000000; // 1807 :   0 - 0x0
      13'h710: dout <= 8'b00000000; // 1808 :   0 - 0x0 -- Sprite 0x71
      13'h711: dout <= 8'b00000000; // 1809 :   0 - 0x0
      13'h712: dout <= 8'b11100000; // 1810 : 224 - 0xe0
      13'h713: dout <= 8'b10000000; // 1811 : 128 - 0x80
      13'h714: dout <= 8'b01000000; // 1812 :  64 - 0x40
      13'h715: dout <= 8'b11110000; // 1813 : 240 - 0xf0
      13'h716: dout <= 8'b10011000; // 1814 : 152 - 0x98
      13'h717: dout <= 8'b11111000; // 1815 : 248 - 0xf8
      13'h718: dout <= 8'b00000000; // 1816 :   0 - 0x0
      13'h719: dout <= 8'b00000000; // 1817 :   0 - 0x0
      13'h71A: dout <= 8'b00000000; // 1818 :   0 - 0x0
      13'h71B: dout <= 8'b00000000; // 1819 :   0 - 0x0
      13'h71C: dout <= 8'b00000000; // 1820 :   0 - 0x0
      13'h71D: dout <= 8'b00000000; // 1821 :   0 - 0x0
      13'h71E: dout <= 8'b00000000; // 1822 :   0 - 0x0
      13'h71F: dout <= 8'b00000000; // 1823 :   0 - 0x0
      13'h720: dout <= 8'b00011111; // 1824 :  31 - 0x1f -- Sprite 0x72
      13'h721: dout <= 8'b00010011; // 1825 :  19 - 0x13
      13'h722: dout <= 8'b00011111; // 1826 :  31 - 0x1f
      13'h723: dout <= 8'b00001111; // 1827 :  15 - 0xf
      13'h724: dout <= 8'b00001001; // 1828 :   9 - 0x9
      13'h725: dout <= 8'b00000111; // 1829 :   7 - 0x7
      13'h726: dout <= 8'b00000001; // 1830 :   1 - 0x1
      13'h727: dout <= 8'b00000000; // 1831 :   0 - 0x0
      13'h728: dout <= 8'b00000000; // 1832 :   0 - 0x0
      13'h729: dout <= 8'b00000000; // 1833 :   0 - 0x0
      13'h72A: dout <= 8'b00000000; // 1834 :   0 - 0x0
      13'h72B: dout <= 8'b00000000; // 1835 :   0 - 0x0
      13'h72C: dout <= 8'b00000000; // 1836 :   0 - 0x0
      13'h72D: dout <= 8'b00000000; // 1837 :   0 - 0x0
      13'h72E: dout <= 8'b00000000; // 1838 :   0 - 0x0
      13'h72F: dout <= 8'b00000000; // 1839 :   0 - 0x0
      13'h730: dout <= 8'b11100100; // 1840 : 228 - 0xe4 -- Sprite 0x73
      13'h731: dout <= 8'b00111100; // 1841 :  60 - 0x3c
      13'h732: dout <= 8'b11100100; // 1842 : 228 - 0xe4
      13'h733: dout <= 8'b00111000; // 1843 :  56 - 0x38
      13'h734: dout <= 8'b11111000; // 1844 : 248 - 0xf8
      13'h735: dout <= 8'b11110000; // 1845 : 240 - 0xf0
      13'h736: dout <= 8'b11000000; // 1846 : 192 - 0xc0
      13'h737: dout <= 8'b00000000; // 1847 :   0 - 0x0
      13'h738: dout <= 8'b00000000; // 1848 :   0 - 0x0
      13'h739: dout <= 8'b00000000; // 1849 :   0 - 0x0
      13'h73A: dout <= 8'b00000000; // 1850 :   0 - 0x0
      13'h73B: dout <= 8'b00000000; // 1851 :   0 - 0x0
      13'h73C: dout <= 8'b00000000; // 1852 :   0 - 0x0
      13'h73D: dout <= 8'b00000000; // 1853 :   0 - 0x0
      13'h73E: dout <= 8'b00000000; // 1854 :   0 - 0x0
      13'h73F: dout <= 8'b00000000; // 1855 :   0 - 0x0
      13'h740: dout <= 8'b00000000; // 1856 :   0 - 0x0 -- Sprite 0x74
      13'h741: dout <= 8'b00000000; // 1857 :   0 - 0x0
      13'h742: dout <= 8'b00000000; // 1858 :   0 - 0x0
      13'h743: dout <= 8'b00000000; // 1859 :   0 - 0x0
      13'h744: dout <= 8'b00000000; // 1860 :   0 - 0x0
      13'h745: dout <= 8'b00000000; // 1861 :   0 - 0x0
      13'h746: dout <= 8'b00000000; // 1862 :   0 - 0x0
      13'h747: dout <= 8'b00000000; // 1863 :   0 - 0x0
      13'h748: dout <= 8'b00000000; // 1864 :   0 - 0x0
      13'h749: dout <= 8'b00000000; // 1865 :   0 - 0x0
      13'h74A: dout <= 8'b00000000; // 1866 :   0 - 0x0
      13'h74B: dout <= 8'b00000000; // 1867 :   0 - 0x0
      13'h74C: dout <= 8'b00010001; // 1868 :  17 - 0x11
      13'h74D: dout <= 8'b00010011; // 1869 :  19 - 0x13
      13'h74E: dout <= 8'b00011111; // 1870 :  31 - 0x1f
      13'h74F: dout <= 8'b00011111; // 1871 :  31 - 0x1f
      13'h750: dout <= 8'b00000000; // 1872 :   0 - 0x0 -- Sprite 0x75
      13'h751: dout <= 8'b00000000; // 1873 :   0 - 0x0
      13'h752: dout <= 8'b00000000; // 1874 :   0 - 0x0
      13'h753: dout <= 8'b00000000; // 1875 :   0 - 0x0
      13'h754: dout <= 8'b00000000; // 1876 :   0 - 0x0
      13'h755: dout <= 8'b00000000; // 1877 :   0 - 0x0
      13'h756: dout <= 8'b00000000; // 1878 :   0 - 0x0
      13'h757: dout <= 8'b00000000; // 1879 :   0 - 0x0
      13'h758: dout <= 8'b00000000; // 1880 :   0 - 0x0
      13'h759: dout <= 8'b00000000; // 1881 :   0 - 0x0
      13'h75A: dout <= 8'b00000000; // 1882 :   0 - 0x0
      13'h75B: dout <= 8'b10000000; // 1883 : 128 - 0x80
      13'h75C: dout <= 8'b11000100; // 1884 : 196 - 0xc4
      13'h75D: dout <= 8'b11100100; // 1885 : 228 - 0xe4
      13'h75E: dout <= 8'b11111100; // 1886 : 252 - 0xfc
      13'h75F: dout <= 8'b11111100; // 1887 : 252 - 0xfc
      13'h760: dout <= 8'b00000000; // 1888 :   0 - 0x0 -- Sprite 0x76
      13'h761: dout <= 8'b00000000; // 1889 :   0 - 0x0
      13'h762: dout <= 8'b00000000; // 1890 :   0 - 0x0
      13'h763: dout <= 8'b00000000; // 1891 :   0 - 0x0
      13'h764: dout <= 8'b00000000; // 1892 :   0 - 0x0
      13'h765: dout <= 8'b00000000; // 1893 :   0 - 0x0
      13'h766: dout <= 8'b00000000; // 1894 :   0 - 0x0
      13'h767: dout <= 8'b00000000; // 1895 :   0 - 0x0
      13'h768: dout <= 8'b00011111; // 1896 :  31 - 0x1f
      13'h769: dout <= 8'b00001110; // 1897 :  14 - 0xe
      13'h76A: dout <= 8'b00000110; // 1898 :   6 - 0x6
      13'h76B: dout <= 8'b00000010; // 1899 :   2 - 0x2
      13'h76C: dout <= 8'b00000000; // 1900 :   0 - 0x0
      13'h76D: dout <= 8'b00000000; // 1901 :   0 - 0x0
      13'h76E: dout <= 8'b00000000; // 1902 :   0 - 0x0
      13'h76F: dout <= 8'b00000000; // 1903 :   0 - 0x0
      13'h770: dout <= 8'b00000000; // 1904 :   0 - 0x0 -- Sprite 0x77
      13'h771: dout <= 8'b00000000; // 1905 :   0 - 0x0
      13'h772: dout <= 8'b00000000; // 1906 :   0 - 0x0
      13'h773: dout <= 8'b00000000; // 1907 :   0 - 0x0
      13'h774: dout <= 8'b00000000; // 1908 :   0 - 0x0
      13'h775: dout <= 8'b00000000; // 1909 :   0 - 0x0
      13'h776: dout <= 8'b00000000; // 1910 :   0 - 0x0
      13'h777: dout <= 8'b00000000; // 1911 :   0 - 0x0
      13'h778: dout <= 8'b11111100; // 1912 : 252 - 0xfc
      13'h779: dout <= 8'b10111000; // 1913 : 184 - 0xb8
      13'h77A: dout <= 8'b10110000; // 1914 : 176 - 0xb0
      13'h77B: dout <= 8'b10100000; // 1915 : 160 - 0xa0
      13'h77C: dout <= 8'b10000000; // 1916 : 128 - 0x80
      13'h77D: dout <= 8'b00000000; // 1917 :   0 - 0x0
      13'h77E: dout <= 8'b00000000; // 1918 :   0 - 0x0
      13'h77F: dout <= 8'b00000000; // 1919 :   0 - 0x0
      13'h780: dout <= 8'b00000000; // 1920 :   0 - 0x0 -- Sprite 0x78
      13'h781: dout <= 8'b00000000; // 1921 :   0 - 0x0
      13'h782: dout <= 8'b00000000; // 1922 :   0 - 0x0
      13'h783: dout <= 8'b00000000; // 1923 :   0 - 0x0
      13'h784: dout <= 8'b00000000; // 1924 :   0 - 0x0
      13'h785: dout <= 8'b00000000; // 1925 :   0 - 0x0
      13'h786: dout <= 8'b00000000; // 1926 :   0 - 0x0
      13'h787: dout <= 8'b00000000; // 1927 :   0 - 0x0
      13'h788: dout <= 8'b00000000; // 1928 :   0 - 0x0
      13'h789: dout <= 8'b00000000; // 1929 :   0 - 0x0
      13'h78A: dout <= 8'b00000000; // 1930 :   0 - 0x0
      13'h78B: dout <= 8'b00000001; // 1931 :   1 - 0x1
      13'h78C: dout <= 8'b00000011; // 1932 :   3 - 0x3
      13'h78D: dout <= 8'b00000110; // 1933 :   6 - 0x6
      13'h78E: dout <= 8'b00000110; // 1934 :   6 - 0x6
      13'h78F: dout <= 8'b00001111; // 1935 :  15 - 0xf
      13'h790: dout <= 8'b00000000; // 1936 :   0 - 0x0 -- Sprite 0x79
      13'h791: dout <= 8'b00000000; // 1937 :   0 - 0x0
      13'h792: dout <= 8'b00000000; // 1938 :   0 - 0x0
      13'h793: dout <= 8'b00000000; // 1939 :   0 - 0x0
      13'h794: dout <= 8'b00000000; // 1940 :   0 - 0x0
      13'h795: dout <= 8'b00000000; // 1941 :   0 - 0x0
      13'h796: dout <= 8'b00000000; // 1942 :   0 - 0x0
      13'h797: dout <= 8'b00000000; // 1943 :   0 - 0x0
      13'h798: dout <= 8'b00000000; // 1944 :   0 - 0x0
      13'h799: dout <= 8'b00011000; // 1945 :  24 - 0x18
      13'h79A: dout <= 8'b11110100; // 1946 : 244 - 0xf4
      13'h79B: dout <= 8'b11111000; // 1947 : 248 - 0xf8
      13'h79C: dout <= 8'b00111000; // 1948 :  56 - 0x38
      13'h79D: dout <= 8'b01111100; // 1949 : 124 - 0x7c
      13'h79E: dout <= 8'b11111100; // 1950 : 252 - 0xfc
      13'h79F: dout <= 8'b11111100; // 1951 : 252 - 0xfc
      13'h7A0: dout <= 8'b00000000; // 1952 :   0 - 0x0 -- Sprite 0x7a
      13'h7A1: dout <= 8'b00000000; // 1953 :   0 - 0x0
      13'h7A2: dout <= 8'b00000000; // 1954 :   0 - 0x0
      13'h7A3: dout <= 8'b00000000; // 1955 :   0 - 0x0
      13'h7A4: dout <= 8'b00000000; // 1956 :   0 - 0x0
      13'h7A5: dout <= 8'b00000000; // 1957 :   0 - 0x0
      13'h7A6: dout <= 8'b00000000; // 1958 :   0 - 0x0
      13'h7A7: dout <= 8'b00000000; // 1959 :   0 - 0x0
      13'h7A8: dout <= 8'b00001111; // 1960 :  15 - 0xf
      13'h7A9: dout <= 8'b00011111; // 1961 :  31 - 0x1f
      13'h7AA: dout <= 8'b00110000; // 1962 :  48 - 0x30
      13'h7AB: dout <= 8'b00111000; // 1963 :  56 - 0x38
      13'h7AC: dout <= 8'b00011101; // 1964 :  29 - 0x1d
      13'h7AD: dout <= 8'b00000011; // 1965 :   3 - 0x3
      13'h7AE: dout <= 8'b00000011; // 1966 :   3 - 0x3
      13'h7AF: dout <= 8'b00000000; // 1967 :   0 - 0x0
      13'h7B0: dout <= 8'b00000000; // 1968 :   0 - 0x0 -- Sprite 0x7b
      13'h7B1: dout <= 8'b00000000; // 1969 :   0 - 0x0
      13'h7B2: dout <= 8'b00000000; // 1970 :   0 - 0x0
      13'h7B3: dout <= 8'b00000000; // 1971 :   0 - 0x0
      13'h7B4: dout <= 8'b00000000; // 1972 :   0 - 0x0
      13'h7B5: dout <= 8'b00000000; // 1973 :   0 - 0x0
      13'h7B6: dout <= 8'b00000000; // 1974 :   0 - 0x0
      13'h7B7: dout <= 8'b00000000; // 1975 :   0 - 0x0
      13'h7B8: dout <= 8'b11111100; // 1976 : 252 - 0xfc
      13'h7B9: dout <= 8'b11111100; // 1977 : 252 - 0xfc
      13'h7BA: dout <= 8'b01111100; // 1978 : 124 - 0x7c
      13'h7BB: dout <= 8'b10001110; // 1979 : 142 - 0x8e
      13'h7BC: dout <= 8'b10000110; // 1980 : 134 - 0x86
      13'h7BD: dout <= 8'b10011100; // 1981 : 156 - 0x9c
      13'h7BE: dout <= 8'b01111000; // 1982 : 120 - 0x78
      13'h7BF: dout <= 8'b00000000; // 1983 :   0 - 0x0
      13'h7C0: dout <= 8'b00000000; // 1984 :   0 - 0x0 -- Sprite 0x7c
      13'h7C1: dout <= 8'b00000001; // 1985 :   1 - 0x1
      13'h7C2: dout <= 8'b00000110; // 1986 :   6 - 0x6
      13'h7C3: dout <= 8'b00000111; // 1987 :   7 - 0x7
      13'h7C4: dout <= 8'b00000111; // 1988 :   7 - 0x7
      13'h7C5: dout <= 8'b00000111; // 1989 :   7 - 0x7
      13'h7C6: dout <= 8'b00000001; // 1990 :   1 - 0x1
      13'h7C7: dout <= 8'b00000011; // 1991 :   3 - 0x3
      13'h7C8: dout <= 8'b00000000; // 1992 :   0 - 0x0
      13'h7C9: dout <= 8'b00000001; // 1993 :   1 - 0x1
      13'h7CA: dout <= 8'b00000110; // 1994 :   6 - 0x6
      13'h7CB: dout <= 8'b00000111; // 1995 :   7 - 0x7
      13'h7CC: dout <= 8'b00000111; // 1996 :   7 - 0x7
      13'h7CD: dout <= 8'b00000111; // 1997 :   7 - 0x7
      13'h7CE: dout <= 8'b00000001; // 1998 :   1 - 0x1
      13'h7CF: dout <= 8'b00000011; // 1999 :   3 - 0x3
      13'h7D0: dout <= 8'b00000000; // 2000 :   0 - 0x0 -- Sprite 0x7d
      13'h7D1: dout <= 8'b11000000; // 2001 : 192 - 0xc0
      13'h7D2: dout <= 8'b00110000; // 2002 :  48 - 0x30
      13'h7D3: dout <= 8'b11110000; // 2003 : 240 - 0xf0
      13'h7D4: dout <= 8'b11110000; // 2004 : 240 - 0xf0
      13'h7D5: dout <= 8'b11110000; // 2005 : 240 - 0xf0
      13'h7D6: dout <= 8'b01000000; // 2006 :  64 - 0x40
      13'h7D7: dout <= 8'b01000000; // 2007 :  64 - 0x40
      13'h7D8: dout <= 8'b00000000; // 2008 :   0 - 0x0
      13'h7D9: dout <= 8'b11000000; // 2009 : 192 - 0xc0
      13'h7DA: dout <= 8'b00110000; // 2010 :  48 - 0x30
      13'h7DB: dout <= 8'b11110000; // 2011 : 240 - 0xf0
      13'h7DC: dout <= 8'b11110000; // 2012 : 240 - 0xf0
      13'h7DD: dout <= 8'b11110000; // 2013 : 240 - 0xf0
      13'h7DE: dout <= 8'b01000000; // 2014 :  64 - 0x40
      13'h7DF: dout <= 8'b01000000; // 2015 :  64 - 0x40
      13'h7E0: dout <= 8'b00000001; // 2016 :   1 - 0x1 -- Sprite 0x7e
      13'h7E1: dout <= 8'b00000000; // 2017 :   0 - 0x0
      13'h7E2: dout <= 8'b00000001; // 2018 :   1 - 0x1
      13'h7E3: dout <= 8'b00000011; // 2019 :   3 - 0x3
      13'h7E4: dout <= 8'b00000001; // 2020 :   1 - 0x1
      13'h7E5: dout <= 8'b00000000; // 2021 :   0 - 0x0
      13'h7E6: dout <= 8'b00000000; // 2022 :   0 - 0x0
      13'h7E7: dout <= 8'b00000000; // 2023 :   0 - 0x0
      13'h7E8: dout <= 8'b00000001; // 2024 :   1 - 0x1
      13'h7E9: dout <= 8'b00000000; // 2025 :   0 - 0x0
      13'h7EA: dout <= 8'b00000001; // 2026 :   1 - 0x1
      13'h7EB: dout <= 8'b00000011; // 2027 :   3 - 0x3
      13'h7EC: dout <= 8'b00000001; // 2028 :   1 - 0x1
      13'h7ED: dout <= 8'b00000000; // 2029 :   0 - 0x0
      13'h7EE: dout <= 8'b00000000; // 2030 :   0 - 0x0
      13'h7EF: dout <= 8'b00000000; // 2031 :   0 - 0x0
      13'h7F0: dout <= 8'b01000000; // 2032 :  64 - 0x40 -- Sprite 0x7f
      13'h7F1: dout <= 8'b01000000; // 2033 :  64 - 0x40
      13'h7F2: dout <= 8'b01000000; // 2034 :  64 - 0x40
      13'h7F3: dout <= 8'b01000000; // 2035 :  64 - 0x40
      13'h7F4: dout <= 8'b01000000; // 2036 :  64 - 0x40
      13'h7F5: dout <= 8'b10000000; // 2037 : 128 - 0x80
      13'h7F6: dout <= 8'b00000000; // 2038 :   0 - 0x0
      13'h7F7: dout <= 8'b00000000; // 2039 :   0 - 0x0
      13'h7F8: dout <= 8'b01000000; // 2040 :  64 - 0x40
      13'h7F9: dout <= 8'b01000000; // 2041 :  64 - 0x40
      13'h7FA: dout <= 8'b01000000; // 2042 :  64 - 0x40
      13'h7FB: dout <= 8'b01000000; // 2043 :  64 - 0x40
      13'h7FC: dout <= 8'b01000000; // 2044 :  64 - 0x40
      13'h7FD: dout <= 8'b10000000; // 2045 : 128 - 0x80
      13'h7FE: dout <= 8'b00000000; // 2046 :   0 - 0x0
      13'h7FF: dout <= 8'b00000000; // 2047 :   0 - 0x0
      13'h800: dout <= 8'b11111111; // 2048 : 255 - 0xff -- Sprite 0x80
      13'h801: dout <= 8'b11111111; // 2049 : 255 - 0xff
      13'h802: dout <= 8'b11111111; // 2050 : 255 - 0xff
      13'h803: dout <= 8'b11111111; // 2051 : 255 - 0xff
      13'h804: dout <= 8'b11000000; // 2052 : 192 - 0xc0
      13'h805: dout <= 8'b11000000; // 2053 : 192 - 0xc0
      13'h806: dout <= 8'b11000000; // 2054 : 192 - 0xc0
      13'h807: dout <= 8'b11000111; // 2055 : 199 - 0xc7
      13'h808: dout <= 8'b00000000; // 2056 :   0 - 0x0
      13'h809: dout <= 8'b00000000; // 2057 :   0 - 0x0
      13'h80A: dout <= 8'b00000000; // 2058 :   0 - 0x0
      13'h80B: dout <= 8'b00000000; // 2059 :   0 - 0x0
      13'h80C: dout <= 8'b00000000; // 2060 :   0 - 0x0
      13'h80D: dout <= 8'b00011111; // 2061 :  31 - 0x1f
      13'h80E: dout <= 8'b00010000; // 2062 :  16 - 0x10
      13'h80F: dout <= 8'b00010111; // 2063 :  23 - 0x17
      13'h810: dout <= 8'b11111111; // 2064 : 255 - 0xff -- Sprite 0x81
      13'h811: dout <= 8'b11111111; // 2065 : 255 - 0xff
      13'h812: dout <= 8'b11111111; // 2066 : 255 - 0xff
      13'h813: dout <= 8'b11111111; // 2067 : 255 - 0xff
      13'h814: dout <= 8'b00000000; // 2068 :   0 - 0x0
      13'h815: dout <= 8'b00000000; // 2069 :   0 - 0x0
      13'h816: dout <= 8'b00000000; // 2070 :   0 - 0x0
      13'h817: dout <= 8'b11111111; // 2071 : 255 - 0xff
      13'h818: dout <= 8'b00000000; // 2072 :   0 - 0x0
      13'h819: dout <= 8'b00000000; // 2073 :   0 - 0x0
      13'h81A: dout <= 8'b00000000; // 2074 :   0 - 0x0
      13'h81B: dout <= 8'b00000000; // 2075 :   0 - 0x0
      13'h81C: dout <= 8'b00000000; // 2076 :   0 - 0x0
      13'h81D: dout <= 8'b11111111; // 2077 : 255 - 0xff
      13'h81E: dout <= 8'b00000000; // 2078 :   0 - 0x0
      13'h81F: dout <= 8'b11111111; // 2079 : 255 - 0xff
      13'h820: dout <= 8'b11111111; // 2080 : 255 - 0xff -- Sprite 0x82
      13'h821: dout <= 8'b11111111; // 2081 : 255 - 0xff
      13'h822: dout <= 8'b11111111; // 2082 : 255 - 0xff
      13'h823: dout <= 8'b11111111; // 2083 : 255 - 0xff
      13'h824: dout <= 8'b01111111; // 2084 : 127 - 0x7f
      13'h825: dout <= 8'b00111111; // 2085 :  63 - 0x3f
      13'h826: dout <= 8'b00011111; // 2086 :  31 - 0x1f
      13'h827: dout <= 8'b11001111; // 2087 : 207 - 0xcf
      13'h828: dout <= 8'b00000000; // 2088 :   0 - 0x0
      13'h829: dout <= 8'b00000000; // 2089 :   0 - 0x0
      13'h82A: dout <= 8'b00000000; // 2090 :   0 - 0x0
      13'h82B: dout <= 8'b00000000; // 2091 :   0 - 0x0
      13'h82C: dout <= 8'b00000000; // 2092 :   0 - 0x0
      13'h82D: dout <= 8'b10000000; // 2093 : 128 - 0x80
      13'h82E: dout <= 8'b00000000; // 2094 :   0 - 0x0
      13'h82F: dout <= 8'b11000000; // 2095 : 192 - 0xc0
      13'h830: dout <= 8'b11111111; // 2096 : 255 - 0xff -- Sprite 0x83
      13'h831: dout <= 8'b11111111; // 2097 : 255 - 0xff
      13'h832: dout <= 8'b11111111; // 2098 : 255 - 0xff
      13'h833: dout <= 8'b11110111; // 2099 : 247 - 0xf7
      13'h834: dout <= 8'b11110111; // 2100 : 247 - 0xf7
      13'h835: dout <= 8'b11100010; // 2101 : 226 - 0xe2
      13'h836: dout <= 8'b11100000; // 2102 : 224 - 0xe0
      13'h837: dout <= 8'b11000110; // 2103 : 198 - 0xc6
      13'h838: dout <= 8'b00000000; // 2104 :   0 - 0x0
      13'h839: dout <= 8'b00000000; // 2105 :   0 - 0x0
      13'h83A: dout <= 8'b00000000; // 2106 :   0 - 0x0
      13'h83B: dout <= 8'b00000000; // 2107 :   0 - 0x0
      13'h83C: dout <= 8'b00000000; // 2108 :   0 - 0x0
      13'h83D: dout <= 8'b00001000; // 2109 :   8 - 0x8
      13'h83E: dout <= 8'b00001000; // 2110 :   8 - 0x8
      13'h83F: dout <= 8'b00010110; // 2111 :  22 - 0x16
      13'h840: dout <= 8'b11111111; // 2112 : 255 - 0xff -- Sprite 0x84
      13'h841: dout <= 8'b11111111; // 2113 : 255 - 0xff
      13'h842: dout <= 8'b11111111; // 2114 : 255 - 0xff
      13'h843: dout <= 8'b11111111; // 2115 : 255 - 0xff
      13'h844: dout <= 8'b10111111; // 2116 : 191 - 0xbf
      13'h845: dout <= 8'b10111111; // 2117 : 191 - 0xbf
      13'h846: dout <= 8'b00011111; // 2118 :  31 - 0x1f
      13'h847: dout <= 8'b00011111; // 2119 :  31 - 0x1f
      13'h848: dout <= 8'b00000000; // 2120 :   0 - 0x0
      13'h849: dout <= 8'b00000000; // 2121 :   0 - 0x0
      13'h84A: dout <= 8'b00000000; // 2122 :   0 - 0x0
      13'h84B: dout <= 8'b00000000; // 2123 :   0 - 0x0
      13'h84C: dout <= 8'b00000000; // 2124 :   0 - 0x0
      13'h84D: dout <= 8'b00000000; // 2125 :   0 - 0x0
      13'h84E: dout <= 8'b01000000; // 2126 :  64 - 0x40
      13'h84F: dout <= 8'b11000000; // 2127 : 192 - 0xc0
      13'h850: dout <= 8'b11111111; // 2128 : 255 - 0xff -- Sprite 0x85
      13'h851: dout <= 8'b11111111; // 2129 : 255 - 0xff
      13'h852: dout <= 8'b11111111; // 2130 : 255 - 0xff
      13'h853: dout <= 8'b11111111; // 2131 : 255 - 0xff
      13'h854: dout <= 8'b11111110; // 2132 : 254 - 0xfe
      13'h855: dout <= 8'b11111000; // 2133 : 248 - 0xf8
      13'h856: dout <= 8'b11100000; // 2134 : 224 - 0xe0
      13'h857: dout <= 8'b11000000; // 2135 : 192 - 0xc0
      13'h858: dout <= 8'b00000000; // 2136 :   0 - 0x0
      13'h859: dout <= 8'b00000000; // 2137 :   0 - 0x0
      13'h85A: dout <= 8'b00000000; // 2138 :   0 - 0x0
      13'h85B: dout <= 8'b00000000; // 2139 :   0 - 0x0
      13'h85C: dout <= 8'b00000000; // 2140 :   0 - 0x0
      13'h85D: dout <= 8'b00000001; // 2141 :   1 - 0x1
      13'h85E: dout <= 8'b00000111; // 2142 :   7 - 0x7
      13'h85F: dout <= 8'b00001100; // 2143 :  12 - 0xc
      13'h860: dout <= 8'b11111111; // 2144 : 255 - 0xff -- Sprite 0x86
      13'h861: dout <= 8'b11111111; // 2145 : 255 - 0xff
      13'h862: dout <= 8'b11111111; // 2146 : 255 - 0xff
      13'h863: dout <= 8'b11111111; // 2147 : 255 - 0xff
      13'h864: dout <= 8'b00000111; // 2148 :   7 - 0x7
      13'h865: dout <= 8'b00000000; // 2149 :   0 - 0x0
      13'h866: dout <= 8'b00111111; // 2150 :  63 - 0x3f
      13'h867: dout <= 8'b11111111; // 2151 : 255 - 0xff
      13'h868: dout <= 8'b00000000; // 2152 :   0 - 0x0
      13'h869: dout <= 8'b00000000; // 2153 :   0 - 0x0
      13'h86A: dout <= 8'b00000000; // 2154 :   0 - 0x0
      13'h86B: dout <= 8'b00000000; // 2155 :   0 - 0x0
      13'h86C: dout <= 8'b00000000; // 2156 :   0 - 0x0
      13'h86D: dout <= 8'b11000000; // 2157 : 192 - 0xc0
      13'h86E: dout <= 8'b00111111; // 2158 :  63 - 0x3f
      13'h86F: dout <= 8'b11111111; // 2159 : 255 - 0xff
      13'h870: dout <= 8'b11111111; // 2160 : 255 - 0xff -- Sprite 0x87
      13'h871: dout <= 8'b11111111; // 2161 : 255 - 0xff
      13'h872: dout <= 8'b11111111; // 2162 : 255 - 0xff
      13'h873: dout <= 8'b11111111; // 2163 : 255 - 0xff
      13'h874: dout <= 8'b11111111; // 2164 : 255 - 0xff
      13'h875: dout <= 8'b11111111; // 2165 : 255 - 0xff
      13'h876: dout <= 8'b00111111; // 2166 :  63 - 0x3f
      13'h877: dout <= 8'b11001111; // 2167 : 207 - 0xcf
      13'h878: dout <= 8'b00000000; // 2168 :   0 - 0x0
      13'h879: dout <= 8'b00000000; // 2169 :   0 - 0x0
      13'h87A: dout <= 8'b00000000; // 2170 :   0 - 0x0
      13'h87B: dout <= 8'b00000000; // 2171 :   0 - 0x0
      13'h87C: dout <= 8'b00000000; // 2172 :   0 - 0x0
      13'h87D: dout <= 8'b00000000; // 2173 :   0 - 0x0
      13'h87E: dout <= 8'b00000000; // 2174 :   0 - 0x0
      13'h87F: dout <= 8'b11000000; // 2175 : 192 - 0xc0
      13'h880: dout <= 8'b11111111; // 2176 : 255 - 0xff -- Sprite 0x88
      13'h881: dout <= 8'b11111111; // 2177 : 255 - 0xff
      13'h882: dout <= 8'b11111111; // 2178 : 255 - 0xff
      13'h883: dout <= 8'b11111111; // 2179 : 255 - 0xff
      13'h884: dout <= 8'b11111111; // 2180 : 255 - 0xff
      13'h885: dout <= 8'b11111111; // 2181 : 255 - 0xff
      13'h886: dout <= 8'b11111111; // 2182 : 255 - 0xff
      13'h887: dout <= 8'b11111111; // 2183 : 255 - 0xff
      13'h888: dout <= 8'b00000000; // 2184 :   0 - 0x0
      13'h889: dout <= 8'b00000000; // 2185 :   0 - 0x0
      13'h88A: dout <= 8'b00000000; // 2186 :   0 - 0x0
      13'h88B: dout <= 8'b00000000; // 2187 :   0 - 0x0
      13'h88C: dout <= 8'b00000000; // 2188 :   0 - 0x0
      13'h88D: dout <= 8'b00000000; // 2189 :   0 - 0x0
      13'h88E: dout <= 8'b00000000; // 2190 :   0 - 0x0
      13'h88F: dout <= 8'b00000000; // 2191 :   0 - 0x0
      13'h890: dout <= 8'b11111111; // 2192 : 255 - 0xff -- Sprite 0x89
      13'h891: dout <= 8'b11111111; // 2193 : 255 - 0xff
      13'h892: dout <= 8'b11111111; // 2194 : 255 - 0xff
      13'h893: dout <= 8'b01110111; // 2195 : 119 - 0x77
      13'h894: dout <= 8'b00010011; // 2196 :  19 - 0x13
      13'h895: dout <= 8'b00000001; // 2197 :   1 - 0x1
      13'h896: dout <= 8'b00010000; // 2198 :  16 - 0x10
      13'h897: dout <= 8'b00011000; // 2199 :  24 - 0x18
      13'h898: dout <= 8'b00000000; // 2200 :   0 - 0x0
      13'h899: dout <= 8'b00000000; // 2201 :   0 - 0x0
      13'h89A: dout <= 8'b00000000; // 2202 :   0 - 0x0
      13'h89B: dout <= 8'b00000000; // 2203 :   0 - 0x0
      13'h89C: dout <= 8'b00000000; // 2204 :   0 - 0x0
      13'h89D: dout <= 8'b01000100; // 2205 :  68 - 0x44
      13'h89E: dout <= 8'b01010110; // 2206 :  86 - 0x56
      13'h89F: dout <= 8'b01011011; // 2207 :  91 - 0x5b
      13'h8A0: dout <= 8'b11111111; // 2208 : 255 - 0xff -- Sprite 0x8a
      13'h8A1: dout <= 8'b11111111; // 2209 : 255 - 0xff
      13'h8A2: dout <= 8'b11111111; // 2210 : 255 - 0xff
      13'h8A3: dout <= 8'b11111111; // 2211 : 255 - 0xff
      13'h8A4: dout <= 8'b11111111; // 2212 : 255 - 0xff
      13'h8A5: dout <= 8'b11111111; // 2213 : 255 - 0xff
      13'h8A6: dout <= 8'b11111111; // 2214 : 255 - 0xff
      13'h8A7: dout <= 8'b01111111; // 2215 : 127 - 0x7f
      13'h8A8: dout <= 8'b00000000; // 2216 :   0 - 0x0
      13'h8A9: dout <= 8'b00000000; // 2217 :   0 - 0x0
      13'h8AA: dout <= 8'b00000000; // 2218 :   0 - 0x0
      13'h8AB: dout <= 8'b00000000; // 2219 :   0 - 0x0
      13'h8AC: dout <= 8'b00000000; // 2220 :   0 - 0x0
      13'h8AD: dout <= 8'b00000000; // 2221 :   0 - 0x0
      13'h8AE: dout <= 8'b00000000; // 2222 :   0 - 0x0
      13'h8AF: dout <= 8'b00000000; // 2223 :   0 - 0x0
      13'h8B0: dout <= 8'b11111111; // 2224 : 255 - 0xff -- Sprite 0x8b
      13'h8B1: dout <= 8'b11111111; // 2225 : 255 - 0xff
      13'h8B2: dout <= 8'b11111111; // 2226 : 255 - 0xff
      13'h8B3: dout <= 8'b11110111; // 2227 : 247 - 0xf7
      13'h8B4: dout <= 8'b11100101; // 2228 : 229 - 0xe5
      13'h8B5: dout <= 8'b11000001; // 2229 : 193 - 0xc1
      13'h8B6: dout <= 8'b10000100; // 2230 : 132 - 0x84
      13'h8B7: dout <= 8'b00001100; // 2231 :  12 - 0xc
      13'h8B8: dout <= 8'b00000000; // 2232 :   0 - 0x0
      13'h8B9: dout <= 8'b00000000; // 2233 :   0 - 0x0
      13'h8BA: dout <= 8'b00000000; // 2234 :   0 - 0x0
      13'h8BB: dout <= 8'b00000000; // 2235 :   0 - 0x0
      13'h8BC: dout <= 8'b00000000; // 2236 :   0 - 0x0
      13'h8BD: dout <= 8'b00010000; // 2237 :  16 - 0x10
      13'h8BE: dout <= 8'b00110100; // 2238 :  52 - 0x34
      13'h8BF: dout <= 8'b01101101; // 2239 : 109 - 0x6d
      13'h8C0: dout <= 8'b11111111; // 2240 : 255 - 0xff -- Sprite 0x8c
      13'h8C1: dout <= 8'b11111111; // 2241 : 255 - 0xff
      13'h8C2: dout <= 8'b11111111; // 2242 : 255 - 0xff
      13'h8C3: dout <= 8'b11111111; // 2243 : 255 - 0xff
      13'h8C4: dout <= 8'b11111111; // 2244 : 255 - 0xff
      13'h8C5: dout <= 8'b01111111; // 2245 : 127 - 0x7f
      13'h8C6: dout <= 8'b01111110; // 2246 : 126 - 0x7e
      13'h8C7: dout <= 8'b01111110; // 2247 : 126 - 0x7e
      13'h8C8: dout <= 8'b00000000; // 2248 :   0 - 0x0
      13'h8C9: dout <= 8'b00000000; // 2249 :   0 - 0x0
      13'h8CA: dout <= 8'b00000000; // 2250 :   0 - 0x0
      13'h8CB: dout <= 8'b00000000; // 2251 :   0 - 0x0
      13'h8CC: dout <= 8'b00000000; // 2252 :   0 - 0x0
      13'h8CD: dout <= 8'b00000000; // 2253 :   0 - 0x0
      13'h8CE: dout <= 8'b00000000; // 2254 :   0 - 0x0
      13'h8CF: dout <= 8'b00000000; // 2255 :   0 - 0x0
      13'h8D0: dout <= 8'b11111111; // 2256 : 255 - 0xff -- Sprite 0x8d
      13'h8D1: dout <= 8'b11111111; // 2257 : 255 - 0xff
      13'h8D2: dout <= 8'b10111111; // 2258 : 191 - 0xbf
      13'h8D3: dout <= 8'b10110111; // 2259 : 183 - 0xb7
      13'h8D4: dout <= 8'b00010111; // 2260 :  23 - 0x17
      13'h8D5: dout <= 8'b00000011; // 2261 :   3 - 0x3
      13'h8D6: dout <= 8'b00100011; // 2262 :  35 - 0x23
      13'h8D7: dout <= 8'b00100001; // 2263 :  33 - 0x21
      13'h8D8: dout <= 8'b00000000; // 2264 :   0 - 0x0
      13'h8D9: dout <= 8'b00000000; // 2265 :   0 - 0x0
      13'h8DA: dout <= 8'b00000000; // 2266 :   0 - 0x0
      13'h8DB: dout <= 8'b00000000; // 2267 :   0 - 0x0
      13'h8DC: dout <= 8'b01000000; // 2268 :  64 - 0x40
      13'h8DD: dout <= 8'b01001000; // 2269 :  72 - 0x48
      13'h8DE: dout <= 8'b10101000; // 2270 : 168 - 0xa8
      13'h8DF: dout <= 8'b10101100; // 2271 : 172 - 0xac
      13'h8E0: dout <= 8'b11111111; // 2272 : 255 - 0xff -- Sprite 0x8e
      13'h8E1: dout <= 8'b11111111; // 2273 : 255 - 0xff
      13'h8E2: dout <= 8'b11111011; // 2274 : 251 - 0xfb
      13'h8E3: dout <= 8'b11111001; // 2275 : 249 - 0xf9
      13'h8E4: dout <= 8'b11111000; // 2276 : 248 - 0xf8
      13'h8E5: dout <= 8'b11111000; // 2277 : 248 - 0xf8
      13'h8E6: dout <= 8'b11111000; // 2278 : 248 - 0xf8
      13'h8E7: dout <= 8'b11111000; // 2279 : 248 - 0xf8
      13'h8E8: dout <= 8'b00000000; // 2280 :   0 - 0x0
      13'h8E9: dout <= 8'b00000000; // 2281 :   0 - 0x0
      13'h8EA: dout <= 8'b00000000; // 2282 :   0 - 0x0
      13'h8EB: dout <= 8'b00000000; // 2283 :   0 - 0x0
      13'h8EC: dout <= 8'b00000010; // 2284 :   2 - 0x2
      13'h8ED: dout <= 8'b00000010; // 2285 :   2 - 0x2
      13'h8EE: dout <= 8'b00000010; // 2286 :   2 - 0x2
      13'h8EF: dout <= 8'b00000010; // 2287 :   2 - 0x2
      13'h8F0: dout <= 8'b11111111; // 2288 : 255 - 0xff -- Sprite 0x8f
      13'h8F1: dout <= 8'b11111111; // 2289 : 255 - 0xff
      13'h8F2: dout <= 8'b01111000; // 2290 : 120 - 0x78
      13'h8F3: dout <= 8'b00111000; // 2291 :  56 - 0x38
      13'h8F4: dout <= 8'b00011000; // 2292 :  24 - 0x18
      13'h8F5: dout <= 8'b00001000; // 2293 :   8 - 0x8
      13'h8F6: dout <= 8'b10000000; // 2294 : 128 - 0x80
      13'h8F7: dout <= 8'b11000000; // 2295 : 192 - 0xc0
      13'h8F8: dout <= 8'b00000000; // 2296 :   0 - 0x0
      13'h8F9: dout <= 8'b00000000; // 2297 :   0 - 0x0
      13'h8FA: dout <= 8'b00000000; // 2298 :   0 - 0x0
      13'h8FB: dout <= 8'b00000011; // 2299 :   3 - 0x3
      13'h8FC: dout <= 8'b01000011; // 2300 :  67 - 0x43
      13'h8FD: dout <= 8'b01100010; // 2301 :  98 - 0x62
      13'h8FE: dout <= 8'b10110010; // 2302 : 178 - 0xb2
      13'h8FF: dout <= 8'b11011010; // 2303 : 218 - 0xda
      13'h900: dout <= 8'b11111111; // 2304 : 255 - 0xff -- Sprite 0x90
      13'h901: dout <= 8'b11111111; // 2305 : 255 - 0xff
      13'h902: dout <= 8'b00000001; // 2306 :   1 - 0x1
      13'h903: dout <= 8'b00000001; // 2307 :   1 - 0x1
      13'h904: dout <= 8'b00000001; // 2308 :   1 - 0x1
      13'h905: dout <= 8'b00000000; // 2309 :   0 - 0x0
      13'h906: dout <= 8'b11111111; // 2310 : 255 - 0xff
      13'h907: dout <= 8'b11111111; // 2311 : 255 - 0xff
      13'h908: dout <= 8'b00000000; // 2312 :   0 - 0x0
      13'h909: dout <= 8'b00000000; // 2313 :   0 - 0x0
      13'h90A: dout <= 8'b00000000; // 2314 :   0 - 0x0
      13'h90B: dout <= 8'b11111100; // 2315 : 252 - 0xfc
      13'h90C: dout <= 8'b11111100; // 2316 : 252 - 0xfc
      13'h90D: dout <= 8'b00000000; // 2317 :   0 - 0x0
      13'h90E: dout <= 8'b11111111; // 2318 : 255 - 0xff
      13'h90F: dout <= 8'b11111111; // 2319 : 255 - 0xff
      13'h910: dout <= 8'b11111111; // 2320 : 255 - 0xff -- Sprite 0x91
      13'h911: dout <= 8'b11111111; // 2321 : 255 - 0xff
      13'h912: dout <= 8'b11111111; // 2322 : 255 - 0xff
      13'h913: dout <= 8'b11111111; // 2323 : 255 - 0xff
      13'h914: dout <= 8'b11111111; // 2324 : 255 - 0xff
      13'h915: dout <= 8'b11111111; // 2325 : 255 - 0xff
      13'h916: dout <= 8'b01111111; // 2326 : 127 - 0x7f
      13'h917: dout <= 8'b00111111; // 2327 :  63 - 0x3f
      13'h918: dout <= 8'b00000000; // 2328 :   0 - 0x0
      13'h919: dout <= 8'b00000000; // 2329 :   0 - 0x0
      13'h91A: dout <= 8'b00000000; // 2330 :   0 - 0x0
      13'h91B: dout <= 8'b00000000; // 2331 :   0 - 0x0
      13'h91C: dout <= 8'b00000000; // 2332 :   0 - 0x0
      13'h91D: dout <= 8'b00000000; // 2333 :   0 - 0x0
      13'h91E: dout <= 8'b00000000; // 2334 :   0 - 0x0
      13'h91F: dout <= 8'b00000000; // 2335 :   0 - 0x0
      13'h920: dout <= 8'b11000111; // 2336 : 199 - 0xc7 -- Sprite 0x92
      13'h921: dout <= 8'b11000111; // 2337 : 199 - 0xc7
      13'h922: dout <= 8'b11000111; // 2338 : 199 - 0xc7
      13'h923: dout <= 8'b11000111; // 2339 : 199 - 0xc7
      13'h924: dout <= 8'b11000111; // 2340 : 199 - 0xc7
      13'h925: dout <= 8'b11000111; // 2341 : 199 - 0xc7
      13'h926: dout <= 8'b11000111; // 2342 : 199 - 0xc7
      13'h927: dout <= 8'b11000111; // 2343 : 199 - 0xc7
      13'h928: dout <= 8'b00010111; // 2344 :  23 - 0x17
      13'h929: dout <= 8'b00010111; // 2345 :  23 - 0x17
      13'h92A: dout <= 8'b00010111; // 2346 :  23 - 0x17
      13'h92B: dout <= 8'b00010111; // 2347 :  23 - 0x17
      13'h92C: dout <= 8'b00010111; // 2348 :  23 - 0x17
      13'h92D: dout <= 8'b00010111; // 2349 :  23 - 0x17
      13'h92E: dout <= 8'b00010111; // 2350 :  23 - 0x17
      13'h92F: dout <= 8'b00010111; // 2351 :  23 - 0x17
      13'h930: dout <= 8'b11111111; // 2352 : 255 - 0xff -- Sprite 0x93
      13'h931: dout <= 8'b11111111; // 2353 : 255 - 0xff
      13'h932: dout <= 8'b11111111; // 2354 : 255 - 0xff
      13'h933: dout <= 8'b11111111; // 2355 : 255 - 0xff
      13'h934: dout <= 8'b11111001; // 2356 : 249 - 0xf9
      13'h935: dout <= 8'b11111001; // 2357 : 249 - 0xf9
      13'h936: dout <= 8'b11111111; // 2358 : 255 - 0xff
      13'h937: dout <= 8'b11111111; // 2359 : 255 - 0xff
      13'h938: dout <= 8'b11111111; // 2360 : 255 - 0xff
      13'h939: dout <= 8'b11111111; // 2361 : 255 - 0xff
      13'h93A: dout <= 8'b11111111; // 2362 : 255 - 0xff
      13'h93B: dout <= 8'b11111111; // 2363 : 255 - 0xff
      13'h93C: dout <= 8'b11111001; // 2364 : 249 - 0xf9
      13'h93D: dout <= 8'b11111001; // 2365 : 249 - 0xf9
      13'h93E: dout <= 8'b11111111; // 2366 : 255 - 0xff
      13'h93F: dout <= 8'b11111111; // 2367 : 255 - 0xff
      13'h940: dout <= 8'b11110111; // 2368 : 247 - 0xf7 -- Sprite 0x94
      13'h941: dout <= 8'b11111011; // 2369 : 251 - 0xfb
      13'h942: dout <= 8'b11111011; // 2370 : 251 - 0xfb
      13'h943: dout <= 8'b11111101; // 2371 : 253 - 0xfd
      13'h944: dout <= 8'b11111100; // 2372 : 252 - 0xfc
      13'h945: dout <= 8'b11111100; // 2373 : 252 - 0xfc
      13'h946: dout <= 8'b01111100; // 2374 : 124 - 0x7c
      13'h947: dout <= 8'b01111100; // 2375 : 124 - 0x7c
      13'h948: dout <= 8'b11110000; // 2376 : 240 - 0xf0
      13'h949: dout <= 8'b11111000; // 2377 : 248 - 0xf8
      13'h94A: dout <= 8'b11111000; // 2378 : 248 - 0xf8
      13'h94B: dout <= 8'b11111100; // 2379 : 252 - 0xfc
      13'h94C: dout <= 8'b11111100; // 2380 : 252 - 0xfc
      13'h94D: dout <= 8'b11111100; // 2381 : 252 - 0xfc
      13'h94E: dout <= 8'b01111100; // 2382 : 124 - 0x7c
      13'h94F: dout <= 8'b01111100; // 2383 : 124 - 0x7c
      13'h950: dout <= 8'b11000111; // 2384 : 199 - 0xc7 -- Sprite 0x95
      13'h951: dout <= 8'b10001111; // 2385 : 143 - 0x8f
      13'h952: dout <= 8'b10001111; // 2386 : 143 - 0x8f
      13'h953: dout <= 8'b00011111; // 2387 :  31 - 0x1f
      13'h954: dout <= 8'b00011111; // 2388 :  31 - 0x1f
      13'h955: dout <= 8'b00111111; // 2389 :  63 - 0x3f
      13'h956: dout <= 8'b00111111; // 2390 :  63 - 0x3f
      13'h957: dout <= 8'b01111111; // 2391 : 127 - 0x7f
      13'h958: dout <= 8'b00010111; // 2392 :  23 - 0x17
      13'h959: dout <= 8'b00101111; // 2393 :  47 - 0x2f
      13'h95A: dout <= 8'b00101111; // 2394 :  47 - 0x2f
      13'h95B: dout <= 8'b01011111; // 2395 :  95 - 0x5f
      13'h95C: dout <= 8'b01011111; // 2396 :  95 - 0x5f
      13'h95D: dout <= 8'b10111111; // 2397 : 191 - 0xbf
      13'h95E: dout <= 8'b10111111; // 2398 : 191 - 0xbf
      13'h95F: dout <= 8'b01111111; // 2399 : 127 - 0x7f
      13'h960: dout <= 8'b00001111; // 2400 :  15 - 0xf -- Sprite 0x96
      13'h961: dout <= 8'b00001111; // 2401 :  15 - 0xf
      13'h962: dout <= 8'b10000111; // 2402 : 135 - 0x87
      13'h963: dout <= 8'b10000111; // 2403 : 135 - 0x87
      13'h964: dout <= 8'b11000010; // 2404 : 194 - 0xc2
      13'h965: dout <= 8'b11000010; // 2405 : 194 - 0xc2
      13'h966: dout <= 8'b11100000; // 2406 : 224 - 0xe0
      13'h967: dout <= 8'b11100000; // 2407 : 224 - 0xe0
      13'h968: dout <= 8'b01100000; // 2408 :  96 - 0x60
      13'h969: dout <= 8'b01100000; // 2409 :  96 - 0x60
      13'h96A: dout <= 8'b10110000; // 2410 : 176 - 0xb0
      13'h96B: dout <= 8'b10110000; // 2411 : 176 - 0xb0
      13'h96C: dout <= 8'b11011000; // 2412 : 216 - 0xd8
      13'h96D: dout <= 8'b11011000; // 2413 : 216 - 0xd8
      13'h96E: dout <= 8'b11101100; // 2414 : 236 - 0xec
      13'h96F: dout <= 8'b11101100; // 2415 : 236 - 0xec
      13'h970: dout <= 8'b10000011; // 2416 : 131 - 0x83 -- Sprite 0x97
      13'h971: dout <= 8'b10001111; // 2417 : 143 - 0x8f
      13'h972: dout <= 8'b00001111; // 2418 :  15 - 0xf
      13'h973: dout <= 8'b00011111; // 2419 :  31 - 0x1f
      13'h974: dout <= 8'b00011111; // 2420 :  31 - 0x1f
      13'h975: dout <= 8'b00111111; // 2421 :  63 - 0x3f
      13'h976: dout <= 8'b00111111; // 2422 :  63 - 0x3f
      13'h977: dout <= 8'b00111111; // 2423 :  63 - 0x3f
      13'h978: dout <= 8'b00110011; // 2424 :  51 - 0x33
      13'h979: dout <= 8'b00101111; // 2425 :  47 - 0x2f
      13'h97A: dout <= 8'b01101111; // 2426 : 111 - 0x6f
      13'h97B: dout <= 8'b01011111; // 2427 :  95 - 0x5f
      13'h97C: dout <= 8'b11011111; // 2428 : 223 - 0xdf
      13'h97D: dout <= 8'b10111111; // 2429 : 191 - 0xbf
      13'h97E: dout <= 8'b10111111; // 2430 : 191 - 0xbf
      13'h97F: dout <= 8'b10111111; // 2431 : 191 - 0xbf
      13'h980: dout <= 8'b11111111; // 2432 : 255 - 0xff -- Sprite 0x98
      13'h981: dout <= 8'b11111111; // 2433 : 255 - 0xff
      13'h982: dout <= 8'b11111111; // 2434 : 255 - 0xff
      13'h983: dout <= 8'b11111110; // 2435 : 254 - 0xfe
      13'h984: dout <= 8'b11111001; // 2436 : 249 - 0xf9
      13'h985: dout <= 8'b11100111; // 2437 : 231 - 0xe7
      13'h986: dout <= 8'b11111100; // 2438 : 252 - 0xfc
      13'h987: dout <= 8'b11110000; // 2439 : 240 - 0xf0
      13'h988: dout <= 8'b11111111; // 2440 : 255 - 0xff
      13'h989: dout <= 8'b11111111; // 2441 : 255 - 0xff
      13'h98A: dout <= 8'b11111111; // 2442 : 255 - 0xff
      13'h98B: dout <= 8'b11111110; // 2443 : 254 - 0xfe
      13'h98C: dout <= 8'b11111001; // 2444 : 249 - 0xf9
      13'h98D: dout <= 8'b11100111; // 2445 : 231 - 0xe7
      13'h98E: dout <= 8'b11111100; // 2446 : 252 - 0xfc
      13'h98F: dout <= 8'b11110011; // 2447 : 243 - 0xf3
      13'h990: dout <= 8'b11110111; // 2448 : 247 - 0xf7 -- Sprite 0x99
      13'h991: dout <= 8'b11111011; // 2449 : 251 - 0xfb
      13'h992: dout <= 8'b11111011; // 2450 : 251 - 0xfb
      13'h993: dout <= 8'b01110011; // 2451 : 115 - 0x73
      13'h994: dout <= 8'b11000001; // 2452 : 193 - 0xc1
      13'h995: dout <= 8'b00000011; // 2453 :   3 - 0x3
      13'h996: dout <= 8'b00001111; // 2454 :  15 - 0xf
      13'h997: dout <= 8'b00111111; // 2455 :  63 - 0x3f
      13'h998: dout <= 8'b11110000; // 2456 : 240 - 0xf0
      13'h999: dout <= 8'b11111000; // 2457 : 248 - 0xf8
      13'h99A: dout <= 8'b11111000; // 2458 : 248 - 0xf8
      13'h99B: dout <= 8'b01110000; // 2459 : 112 - 0x70
      13'h99C: dout <= 8'b11001100; // 2460 : 204 - 0xcc
      13'h99D: dout <= 8'b00110000; // 2461 :  48 - 0x30
      13'h99E: dout <= 8'b11000000; // 2462 : 192 - 0xc0
      13'h99F: dout <= 8'b00000000; // 2463 :   0 - 0x0
      13'h9A0: dout <= 8'b11111111; // 2464 : 255 - 0xff -- Sprite 0x9a
      13'h9A1: dout <= 8'b11111111; // 2465 : 255 - 0xff
      13'h9A2: dout <= 8'b11111111; // 2466 : 255 - 0xff
      13'h9A3: dout <= 8'b10000000; // 2467 : 128 - 0x80
      13'h9A4: dout <= 8'b10000000; // 2468 : 128 - 0x80
      13'h9A5: dout <= 8'b10000000; // 2469 : 128 - 0x80
      13'h9A6: dout <= 8'b10001111; // 2470 : 143 - 0x8f
      13'h9A7: dout <= 8'b10001111; // 2471 : 143 - 0x8f
      13'h9A8: dout <= 8'b00000000; // 2472 :   0 - 0x0
      13'h9A9: dout <= 8'b00000000; // 2473 :   0 - 0x0
      13'h9AA: dout <= 8'b00000000; // 2474 :   0 - 0x0
      13'h9AB: dout <= 8'b00000000; // 2475 :   0 - 0x0
      13'h9AC: dout <= 8'b00111111; // 2476 :  63 - 0x3f
      13'h9AD: dout <= 8'b00100000; // 2477 :  32 - 0x20
      13'h9AE: dout <= 8'b00101111; // 2478 :  47 - 0x2f
      13'h9AF: dout <= 8'b00101111; // 2479 :  47 - 0x2f
      13'h9B0: dout <= 8'b11111111; // 2480 : 255 - 0xff -- Sprite 0x9b
      13'h9B1: dout <= 8'b11111111; // 2481 : 255 - 0xff
      13'h9B2: dout <= 8'b11111111; // 2482 : 255 - 0xff
      13'h9B3: dout <= 8'b00001111; // 2483 :  15 - 0xf
      13'h9B4: dout <= 8'b00001111; // 2484 :  15 - 0xf
      13'h9B5: dout <= 8'b00000111; // 2485 :   7 - 0x7
      13'h9B6: dout <= 8'b11110111; // 2486 : 247 - 0xf7
      13'h9B7: dout <= 8'b11110001; // 2487 : 241 - 0xf1
      13'h9B8: dout <= 8'b00000000; // 2488 :   0 - 0x0
      13'h9B9: dout <= 8'b00000000; // 2489 :   0 - 0x0
      13'h9BA: dout <= 8'b00000000; // 2490 :   0 - 0x0
      13'h9BB: dout <= 8'b00000000; // 2491 :   0 - 0x0
      13'h9BC: dout <= 8'b11100000; // 2492 : 224 - 0xe0
      13'h9BD: dout <= 8'b00000000; // 2493 :   0 - 0x0
      13'h9BE: dout <= 8'b11110000; // 2494 : 240 - 0xf0
      13'h9BF: dout <= 8'b11110000; // 2495 : 240 - 0xf0
      13'h9C0: dout <= 8'b00011100; // 2496 :  28 - 0x1c -- Sprite 0x9c
      13'h9C1: dout <= 8'b00011110; // 2497 :  30 - 0x1e
      13'h9C2: dout <= 8'b00011111; // 2498 :  31 - 0x1f
      13'h9C3: dout <= 8'b00011111; // 2499 :  31 - 0x1f
      13'h9C4: dout <= 8'b00011111; // 2500 :  31 - 0x1f
      13'h9C5: dout <= 8'b00011111; // 2501 :  31 - 0x1f
      13'h9C6: dout <= 8'b00011111; // 2502 :  31 - 0x1f
      13'h9C7: dout <= 8'b00011111; // 2503 :  31 - 0x1f
      13'h9C8: dout <= 8'b01011101; // 2504 :  93 - 0x5d
      13'h9C9: dout <= 8'b01011110; // 2505 :  94 - 0x5e
      13'h9CA: dout <= 8'b01011111; // 2506 :  95 - 0x5f
      13'h9CB: dout <= 8'b01011111; // 2507 :  95 - 0x5f
      13'h9CC: dout <= 8'b01011111; // 2508 :  95 - 0x5f
      13'h9CD: dout <= 8'b01011111; // 2509 :  95 - 0x5f
      13'h9CE: dout <= 8'b01011111; // 2510 :  95 - 0x5f
      13'h9CF: dout <= 8'b01011111; // 2511 :  95 - 0x5f
      13'h9D0: dout <= 8'b00111110; // 2512 :  62 - 0x3e -- Sprite 0x9d
      13'h9D1: dout <= 8'b00011100; // 2513 :  28 - 0x1c
      13'h9D2: dout <= 8'b00001000; // 2514 :   8 - 0x8
      13'h9D3: dout <= 8'b10000000; // 2515 : 128 - 0x80
      13'h9D4: dout <= 8'b11000001; // 2516 : 193 - 0xc1
      13'h9D5: dout <= 8'b11100011; // 2517 : 227 - 0xe3
      13'h9D6: dout <= 8'b11110111; // 2518 : 247 - 0xf7
      13'h9D7: dout <= 8'b11111111; // 2519 : 255 - 0xff
      13'h9D8: dout <= 8'b10000000; // 2520 : 128 - 0x80
      13'h9D9: dout <= 8'b11000001; // 2521 : 193 - 0xc1
      13'h9DA: dout <= 8'b01100011; // 2522 :  99 - 0x63
      13'h9DB: dout <= 8'b10110110; // 2523 : 182 - 0xb6
      13'h9DC: dout <= 8'b11011001; // 2524 : 217 - 0xd9
      13'h9DD: dout <= 8'b11101011; // 2525 : 235 - 0xeb
      13'h9DE: dout <= 8'b11110111; // 2526 : 247 - 0xf7
      13'h9DF: dout <= 8'b11111111; // 2527 : 255 - 0xff
      13'h9E0: dout <= 8'b00011100; // 2528 :  28 - 0x1c -- Sprite 0x9e
      13'h9E1: dout <= 8'b00111100; // 2529 :  60 - 0x3c
      13'h9E2: dout <= 8'b01111100; // 2530 : 124 - 0x7c
      13'h9E3: dout <= 8'b11111100; // 2531 : 252 - 0xfc
      13'h9E4: dout <= 8'b11111100; // 2532 : 252 - 0xfc
      13'h9E5: dout <= 8'b11111100; // 2533 : 252 - 0xfc
      13'h9E6: dout <= 8'b11111100; // 2534 : 252 - 0xfc
      13'h9E7: dout <= 8'b11111100; // 2535 : 252 - 0xfc
      13'h9E8: dout <= 8'b11011101; // 2536 : 221 - 0xdd
      13'h9E9: dout <= 8'b10111101; // 2537 : 189 - 0xbd
      13'h9EA: dout <= 8'b01111101; // 2538 : 125 - 0x7d
      13'h9EB: dout <= 8'b11111101; // 2539 : 253 - 0xfd
      13'h9EC: dout <= 8'b11111101; // 2540 : 253 - 0xfd
      13'h9ED: dout <= 8'b11111101; // 2541 : 253 - 0xfd
      13'h9EE: dout <= 8'b11111101; // 2542 : 253 - 0xfd
      13'h9EF: dout <= 8'b11111101; // 2543 : 253 - 0xfd
      13'h9F0: dout <= 8'b01111100; // 2544 : 124 - 0x7c -- Sprite 0x9f
      13'h9F1: dout <= 8'b01111100; // 2545 : 124 - 0x7c
      13'h9F2: dout <= 8'b01111000; // 2546 : 120 - 0x78
      13'h9F3: dout <= 8'b01111000; // 2547 : 120 - 0x78
      13'h9F4: dout <= 8'b01110001; // 2548 : 113 - 0x71
      13'h9F5: dout <= 8'b01110001; // 2549 : 113 - 0x71
      13'h9F6: dout <= 8'b01100011; // 2550 :  99 - 0x63
      13'h9F7: dout <= 8'b01100011; // 2551 :  99 - 0x63
      13'h9F8: dout <= 8'b00000001; // 2552 :   1 - 0x1
      13'h9F9: dout <= 8'b00000001; // 2553 :   1 - 0x1
      13'h9FA: dout <= 8'b00000010; // 2554 :   2 - 0x2
      13'h9FB: dout <= 8'b00000010; // 2555 :   2 - 0x2
      13'h9FC: dout <= 8'b00000101; // 2556 :   5 - 0x5
      13'h9FD: dout <= 8'b00000101; // 2557 :   5 - 0x5
      13'h9FE: dout <= 8'b00001011; // 2558 :  11 - 0xb
      13'h9FF: dout <= 8'b00001011; // 2559 :  11 - 0xb
      13'hA00: dout <= 8'b01110001; // 2560 : 113 - 0x71 -- Sprite 0xa0
      13'hA01: dout <= 8'b01110000; // 2561 : 112 - 0x70
      13'hA02: dout <= 8'b11111000; // 2562 : 248 - 0xf8
      13'hA03: dout <= 8'b11111000; // 2563 : 248 - 0xf8
      13'hA04: dout <= 8'b11111100; // 2564 : 252 - 0xfc
      13'hA05: dout <= 8'b11111100; // 2565 : 252 - 0xfc
      13'hA06: dout <= 8'b11111110; // 2566 : 254 - 0xfe
      13'hA07: dout <= 8'b11111110; // 2567 : 254 - 0xfe
      13'hA08: dout <= 8'b01110100; // 2568 : 116 - 0x74
      13'hA09: dout <= 8'b01110110; // 2569 : 118 - 0x76
      13'hA0A: dout <= 8'b11111010; // 2570 : 250 - 0xfa
      13'hA0B: dout <= 8'b11111011; // 2571 : 251 - 0xfb
      13'hA0C: dout <= 8'b11111101; // 2572 : 253 - 0xfd
      13'hA0D: dout <= 8'b11111101; // 2573 : 253 - 0xfd
      13'hA0E: dout <= 8'b11111110; // 2574 : 254 - 0xfe
      13'hA0F: dout <= 8'b11111110; // 2575 : 254 - 0xfe
      13'hA10: dout <= 8'b11111000; // 2576 : 248 - 0xf8 -- Sprite 0xa1
      13'hA11: dout <= 8'b11111000; // 2577 : 248 - 0xf8
      13'hA12: dout <= 8'b11111000; // 2578 : 248 - 0xf8
      13'hA13: dout <= 8'b01111000; // 2579 : 120 - 0x78
      13'hA14: dout <= 8'b01111000; // 2580 : 120 - 0x78
      13'hA15: dout <= 8'b00111000; // 2581 :  56 - 0x38
      13'hA16: dout <= 8'b00111000; // 2582 :  56 - 0x38
      13'hA17: dout <= 8'b00011000; // 2583 :  24 - 0x18
      13'hA18: dout <= 8'b00000010; // 2584 :   2 - 0x2
      13'hA19: dout <= 8'b00000010; // 2585 :   2 - 0x2
      13'hA1A: dout <= 8'b00000010; // 2586 :   2 - 0x2
      13'hA1B: dout <= 8'b00000010; // 2587 :   2 - 0x2
      13'hA1C: dout <= 8'b00000010; // 2588 :   2 - 0x2
      13'hA1D: dout <= 8'b10000010; // 2589 : 130 - 0x82
      13'hA1E: dout <= 8'b10000010; // 2590 : 130 - 0x82
      13'hA1F: dout <= 8'b11000010; // 2591 : 194 - 0xc2
      13'hA20: dout <= 8'b11100000; // 2592 : 224 - 0xe0 -- Sprite 0xa2
      13'hA21: dout <= 8'b11110000; // 2593 : 240 - 0xf0
      13'hA22: dout <= 8'b11111000; // 2594 : 248 - 0xf8
      13'hA23: dout <= 8'b11111000; // 2595 : 248 - 0xf8
      13'hA24: dout <= 8'b11111100; // 2596 : 252 - 0xfc
      13'hA25: dout <= 8'b11111100; // 2597 : 252 - 0xfc
      13'hA26: dout <= 8'b11111110; // 2598 : 254 - 0xfe
      13'hA27: dout <= 8'b11111111; // 2599 : 255 - 0xff
      13'hA28: dout <= 8'b11101010; // 2600 : 234 - 0xea
      13'hA29: dout <= 8'b11110110; // 2601 : 246 - 0xf6
      13'hA2A: dout <= 8'b11111010; // 2602 : 250 - 0xfa
      13'hA2B: dout <= 8'b11111010; // 2603 : 250 - 0xfa
      13'hA2C: dout <= 8'b11111100; // 2604 : 252 - 0xfc
      13'hA2D: dout <= 8'b11111100; // 2605 : 252 - 0xfc
      13'hA2E: dout <= 8'b11111110; // 2606 : 254 - 0xfe
      13'hA2F: dout <= 8'b11111111; // 2607 : 255 - 0xff
      13'hA30: dout <= 8'b11111111; // 2608 : 255 - 0xff -- Sprite 0xa3
      13'hA31: dout <= 8'b11111111; // 2609 : 255 - 0xff
      13'hA32: dout <= 8'b11111111; // 2610 : 255 - 0xff
      13'hA33: dout <= 8'b11111111; // 2611 : 255 - 0xff
      13'hA34: dout <= 8'b11111111; // 2612 : 255 - 0xff
      13'hA35: dout <= 8'b11111111; // 2613 : 255 - 0xff
      13'hA36: dout <= 8'b11111111; // 2614 : 255 - 0xff
      13'hA37: dout <= 8'b11111111; // 2615 : 255 - 0xff
      13'hA38: dout <= 8'b11111111; // 2616 : 255 - 0xff
      13'hA39: dout <= 8'b11111111; // 2617 : 255 - 0xff
      13'hA3A: dout <= 8'b11111111; // 2618 : 255 - 0xff
      13'hA3B: dout <= 8'b11111111; // 2619 : 255 - 0xff
      13'hA3C: dout <= 8'b11111111; // 2620 : 255 - 0xff
      13'hA3D: dout <= 8'b11111111; // 2621 : 255 - 0xff
      13'hA3E: dout <= 8'b11111111; // 2622 : 255 - 0xff
      13'hA3F: dout <= 8'b11111111; // 2623 : 255 - 0xff
      13'hA40: dout <= 8'b00011111; // 2624 :  31 - 0x1f -- Sprite 0xa4
      13'hA41: dout <= 8'b00011111; // 2625 :  31 - 0x1f
      13'hA42: dout <= 8'b00011111; // 2626 :  31 - 0x1f
      13'hA43: dout <= 8'b00011111; // 2627 :  31 - 0x1f
      13'hA44: dout <= 8'b00011111; // 2628 :  31 - 0x1f
      13'hA45: dout <= 8'b00011111; // 2629 :  31 - 0x1f
      13'hA46: dout <= 8'b00011111; // 2630 :  31 - 0x1f
      13'hA47: dout <= 8'b00011111; // 2631 :  31 - 0x1f
      13'hA48: dout <= 8'b01000000; // 2632 :  64 - 0x40
      13'hA49: dout <= 8'b01000000; // 2633 :  64 - 0x40
      13'hA4A: dout <= 8'b01000000; // 2634 :  64 - 0x40
      13'hA4B: dout <= 8'b01000000; // 2635 :  64 - 0x40
      13'hA4C: dout <= 8'b01000000; // 2636 :  64 - 0x40
      13'hA4D: dout <= 8'b01000000; // 2637 :  64 - 0x40
      13'hA4E: dout <= 8'b01000000; // 2638 :  64 - 0x40
      13'hA4F: dout <= 8'b01000000; // 2639 :  64 - 0x40
      13'hA50: dout <= 8'b11111000; // 2640 : 248 - 0xf8 -- Sprite 0xa5
      13'hA51: dout <= 8'b11111111; // 2641 : 255 - 0xff
      13'hA52: dout <= 8'b11111111; // 2642 : 255 - 0xff
      13'hA53: dout <= 8'b11111000; // 2643 : 248 - 0xf8
      13'hA54: dout <= 8'b11111000; // 2644 : 248 - 0xf8
      13'hA55: dout <= 8'b11111000; // 2645 : 248 - 0xf8
      13'hA56: dout <= 8'b11111000; // 2646 : 248 - 0xf8
      13'hA57: dout <= 8'b11111000; // 2647 : 248 - 0xf8
      13'hA58: dout <= 8'b11111000; // 2648 : 248 - 0xf8
      13'hA59: dout <= 8'b11111111; // 2649 : 255 - 0xff
      13'hA5A: dout <= 8'b11111111; // 2650 : 255 - 0xff
      13'hA5B: dout <= 8'b11111000; // 2651 : 248 - 0xf8
      13'hA5C: dout <= 8'b11111011; // 2652 : 251 - 0xfb
      13'hA5D: dout <= 8'b11111010; // 2653 : 250 - 0xfa
      13'hA5E: dout <= 8'b11111010; // 2654 : 250 - 0xfa
      13'hA5F: dout <= 8'b11111010; // 2655 : 250 - 0xfa
      13'hA60: dout <= 8'b11111100; // 2656 : 252 - 0xfc -- Sprite 0xa6
      13'hA61: dout <= 8'b11111000; // 2657 : 248 - 0xf8
      13'hA62: dout <= 8'b11110000; // 2658 : 240 - 0xf0
      13'hA63: dout <= 8'b00000001; // 2659 :   1 - 0x1
      13'hA64: dout <= 8'b00000001; // 2660 :   1 - 0x1
      13'hA65: dout <= 8'b00000011; // 2661 :   3 - 0x3
      13'hA66: dout <= 8'b11000011; // 2662 : 195 - 0xc3
      13'hA67: dout <= 8'b10000111; // 2663 : 135 - 0x87
      13'hA68: dout <= 8'b11111100; // 2664 : 252 - 0xfc
      13'hA69: dout <= 8'b11111010; // 2665 : 250 - 0xfa
      13'hA6A: dout <= 8'b11110110; // 2666 : 246 - 0xf6
      13'hA6B: dout <= 8'b00001101; // 2667 :  13 - 0xd
      13'hA6C: dout <= 8'b11111001; // 2668 : 249 - 0xf9
      13'hA6D: dout <= 8'b00000011; // 2669 :   3 - 0x3
      13'hA6E: dout <= 8'b00010011; // 2670 :  19 - 0x13
      13'hA6F: dout <= 8'b00110111; // 2671 :  55 - 0x37
      13'hA70: dout <= 8'b01111111; // 2672 : 127 - 0x7f -- Sprite 0xa7
      13'hA71: dout <= 8'b11111001; // 2673 : 249 - 0xf9
      13'hA72: dout <= 8'b11111001; // 2674 : 249 - 0xf9
      13'hA73: dout <= 8'b11111111; // 2675 : 255 - 0xff
      13'hA74: dout <= 8'b11111110; // 2676 : 254 - 0xfe
      13'hA75: dout <= 8'b11111100; // 2677 : 252 - 0xfc
      13'hA76: dout <= 8'b11111111; // 2678 : 255 - 0xff
      13'hA77: dout <= 8'b11111111; // 2679 : 255 - 0xff
      13'hA78: dout <= 8'b01111111; // 2680 : 127 - 0x7f
      13'hA79: dout <= 8'b11111001; // 2681 : 249 - 0xf9
      13'hA7A: dout <= 8'b11111001; // 2682 : 249 - 0xf9
      13'hA7B: dout <= 8'b11111111; // 2683 : 255 - 0xff
      13'hA7C: dout <= 8'b11111110; // 2684 : 254 - 0xfe
      13'hA7D: dout <= 8'b11111100; // 2685 : 252 - 0xfc
      13'hA7E: dout <= 8'b11111111; // 2686 : 255 - 0xff
      13'hA7F: dout <= 8'b11111111; // 2687 : 255 - 0xff
      13'hA80: dout <= 8'b11110000; // 2688 : 240 - 0xf0 -- Sprite 0xa8
      13'hA81: dout <= 8'b11110000; // 2689 : 240 - 0xf0
      13'hA82: dout <= 8'b11111000; // 2690 : 248 - 0xf8
      13'hA83: dout <= 8'b01111000; // 2691 : 120 - 0x78
      13'hA84: dout <= 8'b11111100; // 2692 : 252 - 0xfc
      13'hA85: dout <= 8'b11110100; // 2693 : 244 - 0xf4
      13'hA86: dout <= 8'b11110110; // 2694 : 246 - 0xf6
      13'hA87: dout <= 8'b11111010; // 2695 : 250 - 0xfa
      13'hA88: dout <= 8'b11110110; // 2696 : 246 - 0xf6
      13'hA89: dout <= 8'b11110110; // 2697 : 246 - 0xf6
      13'hA8A: dout <= 8'b11111011; // 2698 : 251 - 0xfb
      13'hA8B: dout <= 8'b01111011; // 2699 : 123 - 0x7b
      13'hA8C: dout <= 8'b11111101; // 2700 : 253 - 0xfd
      13'hA8D: dout <= 8'b11110101; // 2701 : 245 - 0xf5
      13'hA8E: dout <= 8'b11110110; // 2702 : 246 - 0xf6
      13'hA8F: dout <= 8'b11111010; // 2703 : 250 - 0xfa
      13'hA90: dout <= 8'b00111111; // 2704 :  63 - 0x3f -- Sprite 0xa9
      13'hA91: dout <= 8'b00111111; // 2705 :  63 - 0x3f
      13'hA92: dout <= 8'b00111111; // 2706 :  63 - 0x3f
      13'hA93: dout <= 8'b00111111; // 2707 :  63 - 0x3f
      13'hA94: dout <= 8'b00111111; // 2708 :  63 - 0x3f
      13'hA95: dout <= 8'b00011111; // 2709 :  31 - 0x1f
      13'hA96: dout <= 8'b00001111; // 2710 :  15 - 0xf
      13'hA97: dout <= 8'b00000111; // 2711 :   7 - 0x7
      13'hA98: dout <= 8'b10111111; // 2712 : 191 - 0xbf
      13'hA99: dout <= 8'b10111111; // 2713 : 191 - 0xbf
      13'hA9A: dout <= 8'b00111111; // 2714 :  63 - 0x3f
      13'hA9B: dout <= 8'b00111111; // 2715 :  63 - 0x3f
      13'hA9C: dout <= 8'b10111111; // 2716 : 191 - 0xbf
      13'hA9D: dout <= 8'b10011111; // 2717 : 159 - 0x9f
      13'hA9E: dout <= 8'b11001111; // 2718 : 207 - 0xcf
      13'hA9F: dout <= 8'b11010111; // 2719 : 215 - 0xd7
      13'hAA0: dout <= 8'b11100000; // 2720 : 224 - 0xe0 -- Sprite 0xaa
      13'hAA1: dout <= 8'b11111000; // 2721 : 248 - 0xf8
      13'hAA2: dout <= 8'b11111111; // 2722 : 255 - 0xff
      13'hAA3: dout <= 8'b11110011; // 2723 : 243 - 0xf3
      13'hAA4: dout <= 8'b11111100; // 2724 : 252 - 0xfc
      13'hAA5: dout <= 8'b11111111; // 2725 : 255 - 0xff
      13'hAA6: dout <= 8'b11111111; // 2726 : 255 - 0xff
      13'hAA7: dout <= 8'b11111111; // 2727 : 255 - 0xff
      13'hAA8: dout <= 8'b11100100; // 2728 : 228 - 0xe4
      13'hAA9: dout <= 8'b11111000; // 2729 : 248 - 0xf8
      13'hAAA: dout <= 8'b11111111; // 2730 : 255 - 0xff
      13'hAAB: dout <= 8'b11110011; // 2731 : 243 - 0xf3
      13'hAAC: dout <= 8'b11111100; // 2732 : 252 - 0xfc
      13'hAAD: dout <= 8'b11111111; // 2733 : 255 - 0xff
      13'hAAE: dout <= 8'b11111111; // 2734 : 255 - 0xff
      13'hAAF: dout <= 8'b11111111; // 2735 : 255 - 0xff
      13'hAB0: dout <= 8'b11111111; // 2736 : 255 - 0xff -- Sprite 0xab
      13'hAB1: dout <= 8'b11111111; // 2737 : 255 - 0xff
      13'hAB2: dout <= 8'b00111111; // 2738 :  63 - 0x3f
      13'hAB3: dout <= 8'b11001111; // 2739 : 207 - 0xcf
      13'hAB4: dout <= 8'b11110011; // 2740 : 243 - 0xf3
      13'hAB5: dout <= 8'b00111101; // 2741 :  61 - 0x3d
      13'hAB6: dout <= 8'b11011000; // 2742 : 216 - 0xd8
      13'hAB7: dout <= 8'b10110000; // 2743 : 176 - 0xb0
      13'hAB8: dout <= 8'b00000000; // 2744 :   0 - 0x0
      13'hAB9: dout <= 8'b00000000; // 2745 :   0 - 0x0
      13'hABA: dout <= 8'b00000000; // 2746 :   0 - 0x0
      13'hABB: dout <= 8'b11000000; // 2747 : 192 - 0xc0
      13'hABC: dout <= 8'b11110000; // 2748 : 240 - 0xf0
      13'hABD: dout <= 8'b00111100; // 2749 :  60 - 0x3c
      13'hABE: dout <= 8'b11011000; // 2750 : 216 - 0xd8
      13'hABF: dout <= 8'b10110110; // 2751 : 182 - 0xb6
      13'hAC0: dout <= 8'b10001111; // 2752 : 143 - 0x8f -- Sprite 0xac
      13'hAC1: dout <= 8'b11101111; // 2753 : 239 - 0xef
      13'hAC2: dout <= 8'b11100000; // 2754 : 224 - 0xe0
      13'hAC3: dout <= 8'b11111000; // 2755 : 248 - 0xf8
      13'hAC4: dout <= 8'b11111000; // 2756 : 248 - 0xf8
      13'hAC5: dout <= 8'b11111111; // 2757 : 255 - 0xff
      13'hAC6: dout <= 8'b11111111; // 2758 : 255 - 0xff
      13'hAC7: dout <= 8'b11111111; // 2759 : 255 - 0xff
      13'hAC8: dout <= 8'b00001111; // 2760 :  15 - 0xf
      13'hAC9: dout <= 8'b00001111; // 2761 :  15 - 0xf
      13'hACA: dout <= 8'b00000000; // 2762 :   0 - 0x0
      13'hACB: dout <= 8'b00000011; // 2763 :   3 - 0x3
      13'hACC: dout <= 8'b00000000; // 2764 :   0 - 0x0
      13'hACD: dout <= 8'b00000000; // 2765 :   0 - 0x0
      13'hACE: dout <= 8'b00000000; // 2766 :   0 - 0x0
      13'hACF: dout <= 8'b00000000; // 2767 :   0 - 0x0
      13'hAD0: dout <= 8'b11110001; // 2768 : 241 - 0xf1 -- Sprite 0xad
      13'hAD1: dout <= 8'b11110001; // 2769 : 241 - 0xf1
      13'hAD2: dout <= 8'b00000001; // 2770 :   1 - 0x1
      13'hAD3: dout <= 8'b00000001; // 2771 :   1 - 0x1
      13'hAD4: dout <= 8'b00000001; // 2772 :   1 - 0x1
      13'hAD5: dout <= 8'b11111111; // 2773 : 255 - 0xff
      13'hAD6: dout <= 8'b11111111; // 2774 : 255 - 0xff
      13'hAD7: dout <= 8'b11111111; // 2775 : 255 - 0xff
      13'hAD8: dout <= 8'b11110100; // 2776 : 244 - 0xf4
      13'hAD9: dout <= 8'b11110100; // 2777 : 244 - 0xf4
      13'hADA: dout <= 8'b00000100; // 2778 :   4 - 0x4
      13'hADB: dout <= 8'b11111100; // 2779 : 252 - 0xfc
      13'hADC: dout <= 8'b00000000; // 2780 :   0 - 0x0
      13'hADD: dout <= 8'b00000000; // 2781 :   0 - 0x0
      13'hADE: dout <= 8'b00000000; // 2782 :   0 - 0x0
      13'hADF: dout <= 8'b00000000; // 2783 :   0 - 0x0
      13'hAE0: dout <= 8'b00011111; // 2784 :  31 - 0x1f -- Sprite 0xae
      13'hAE1: dout <= 8'b00011111; // 2785 :  31 - 0x1f
      13'hAE2: dout <= 8'b00011111; // 2786 :  31 - 0x1f
      13'hAE3: dout <= 8'b00011111; // 2787 :  31 - 0x1f
      13'hAE4: dout <= 8'b00011111; // 2788 :  31 - 0x1f
      13'hAE5: dout <= 8'b00011111; // 2789 :  31 - 0x1f
      13'hAE6: dout <= 8'b00011111; // 2790 :  31 - 0x1f
      13'hAE7: dout <= 8'b00011111; // 2791 :  31 - 0x1f
      13'hAE8: dout <= 8'b01011111; // 2792 :  95 - 0x5f
      13'hAE9: dout <= 8'b01011111; // 2793 :  95 - 0x5f
      13'hAEA: dout <= 8'b01011111; // 2794 :  95 - 0x5f
      13'hAEB: dout <= 8'b01011111; // 2795 :  95 - 0x5f
      13'hAEC: dout <= 8'b01011111; // 2796 :  95 - 0x5f
      13'hAED: dout <= 8'b01011111; // 2797 :  95 - 0x5f
      13'hAEE: dout <= 8'b01011111; // 2798 :  95 - 0x5f
      13'hAEF: dout <= 8'b01011111; // 2799 :  95 - 0x5f
      13'hAF0: dout <= 8'b11111100; // 2800 : 252 - 0xfc -- Sprite 0xaf
      13'hAF1: dout <= 8'b11111100; // 2801 : 252 - 0xfc
      13'hAF2: dout <= 8'b11111100; // 2802 : 252 - 0xfc
      13'hAF3: dout <= 8'b11111100; // 2803 : 252 - 0xfc
      13'hAF4: dout <= 8'b11110100; // 2804 : 244 - 0xf4
      13'hAF5: dout <= 8'b11110100; // 2805 : 244 - 0xf4
      13'hAF6: dout <= 8'b11110100; // 2806 : 244 - 0xf4
      13'hAF7: dout <= 8'b11110100; // 2807 : 244 - 0xf4
      13'hAF8: dout <= 8'b11111101; // 2808 : 253 - 0xfd
      13'hAF9: dout <= 8'b11111101; // 2809 : 253 - 0xfd
      13'hAFA: dout <= 8'b11111101; // 2810 : 253 - 0xfd
      13'hAFB: dout <= 8'b11111101; // 2811 : 253 - 0xfd
      13'hAFC: dout <= 8'b11110101; // 2812 : 245 - 0xf5
      13'hAFD: dout <= 8'b11110101; // 2813 : 245 - 0xf5
      13'hAFE: dout <= 8'b11110101; // 2814 : 245 - 0xf5
      13'hAFF: dout <= 8'b11110101; // 2815 : 245 - 0xf5
      13'hB00: dout <= 8'b00001100; // 2816 :  12 - 0xc -- Sprite 0xb0
      13'hB01: dout <= 8'b00011100; // 2817 :  28 - 0x1c
      13'hB02: dout <= 8'b00001100; // 2818 :  12 - 0xc
      13'hB03: dout <= 8'b00001100; // 2819 :  12 - 0xc
      13'hB04: dout <= 8'b00001100; // 2820 :  12 - 0xc
      13'hB05: dout <= 8'b00001100; // 2821 :  12 - 0xc
      13'hB06: dout <= 8'b00111111; // 2822 :  63 - 0x3f
      13'hB07: dout <= 8'b00000000; // 2823 :   0 - 0x0
      13'hB08: dout <= 8'b00001100; // 2824 :  12 - 0xc
      13'hB09: dout <= 8'b00011100; // 2825 :  28 - 0x1c
      13'hB0A: dout <= 8'b00001100; // 2826 :  12 - 0xc
      13'hB0B: dout <= 8'b00001100; // 2827 :  12 - 0xc
      13'hB0C: dout <= 8'b00001100; // 2828 :  12 - 0xc
      13'hB0D: dout <= 8'b00001100; // 2829 :  12 - 0xc
      13'hB0E: dout <= 8'b00111111; // 2830 :  63 - 0x3f
      13'hB0F: dout <= 8'b00000000; // 2831 :   0 - 0x0
      13'hB10: dout <= 8'b00111110; // 2832 :  62 - 0x3e -- Sprite 0xb1
      13'hB11: dout <= 8'b01100011; // 2833 :  99 - 0x63
      13'hB12: dout <= 8'b00000111; // 2834 :   7 - 0x7
      13'hB13: dout <= 8'b00011110; // 2835 :  30 - 0x1e
      13'hB14: dout <= 8'b00111100; // 2836 :  60 - 0x3c
      13'hB15: dout <= 8'b01110000; // 2837 : 112 - 0x70
      13'hB16: dout <= 8'b01111111; // 2838 : 127 - 0x7f
      13'hB17: dout <= 8'b00000000; // 2839 :   0 - 0x0
      13'hB18: dout <= 8'b00111110; // 2840 :  62 - 0x3e
      13'hB19: dout <= 8'b01100011; // 2841 :  99 - 0x63
      13'hB1A: dout <= 8'b00000111; // 2842 :   7 - 0x7
      13'hB1B: dout <= 8'b00011110; // 2843 :  30 - 0x1e
      13'hB1C: dout <= 8'b00111100; // 2844 :  60 - 0x3c
      13'hB1D: dout <= 8'b01110000; // 2845 : 112 - 0x70
      13'hB1E: dout <= 8'b01111111; // 2846 : 127 - 0x7f
      13'hB1F: dout <= 8'b00000000; // 2847 :   0 - 0x0
      13'hB20: dout <= 8'b01111110; // 2848 : 126 - 0x7e -- Sprite 0xb2
      13'hB21: dout <= 8'b01100011; // 2849 :  99 - 0x63
      13'hB22: dout <= 8'b01100011; // 2850 :  99 - 0x63
      13'hB23: dout <= 8'b01100011; // 2851 :  99 - 0x63
      13'hB24: dout <= 8'b01111110; // 2852 : 126 - 0x7e
      13'hB25: dout <= 8'b01100000; // 2853 :  96 - 0x60
      13'hB26: dout <= 8'b01100000; // 2854 :  96 - 0x60
      13'hB27: dout <= 8'b00000000; // 2855 :   0 - 0x0
      13'hB28: dout <= 8'b01111110; // 2856 : 126 - 0x7e
      13'hB29: dout <= 8'b01100011; // 2857 :  99 - 0x63
      13'hB2A: dout <= 8'b01100011; // 2858 :  99 - 0x63
      13'hB2B: dout <= 8'b01100011; // 2859 :  99 - 0x63
      13'hB2C: dout <= 8'b01111110; // 2860 : 126 - 0x7e
      13'hB2D: dout <= 8'b01100000; // 2861 :  96 - 0x60
      13'hB2E: dout <= 8'b01100000; // 2862 :  96 - 0x60
      13'hB2F: dout <= 8'b00000000; // 2863 :   0 - 0x0
      13'hB30: dout <= 8'b01100011; // 2864 :  99 - 0x63 -- Sprite 0xb3
      13'hB31: dout <= 8'b01100011; // 2865 :  99 - 0x63
      13'hB32: dout <= 8'b01100011; // 2866 :  99 - 0x63
      13'hB33: dout <= 8'b01100011; // 2867 :  99 - 0x63
      13'hB34: dout <= 8'b01100011; // 2868 :  99 - 0x63
      13'hB35: dout <= 8'b01100011; // 2869 :  99 - 0x63
      13'hB36: dout <= 8'b00111110; // 2870 :  62 - 0x3e
      13'hB37: dout <= 8'b00000000; // 2871 :   0 - 0x0
      13'hB38: dout <= 8'b01100011; // 2872 :  99 - 0x63
      13'hB39: dout <= 8'b01100011; // 2873 :  99 - 0x63
      13'hB3A: dout <= 8'b01100011; // 2874 :  99 - 0x63
      13'hB3B: dout <= 8'b01100011; // 2875 :  99 - 0x63
      13'hB3C: dout <= 8'b01100011; // 2876 :  99 - 0x63
      13'hB3D: dout <= 8'b01100011; // 2877 :  99 - 0x63
      13'hB3E: dout <= 8'b00111110; // 2878 :  62 - 0x3e
      13'hB3F: dout <= 8'b00000000; // 2879 :   0 - 0x0
      13'hB40: dout <= 8'b01100011; // 2880 :  99 - 0x63 -- Sprite 0xb4
      13'hB41: dout <= 8'b01100011; // 2881 :  99 - 0x63
      13'hB42: dout <= 8'b01100011; // 2882 :  99 - 0x63
      13'hB43: dout <= 8'b01111111; // 2883 : 127 - 0x7f
      13'hB44: dout <= 8'b01100011; // 2884 :  99 - 0x63
      13'hB45: dout <= 8'b01100011; // 2885 :  99 - 0x63
      13'hB46: dout <= 8'b01100011; // 2886 :  99 - 0x63
      13'hB47: dout <= 8'b00000000; // 2887 :   0 - 0x0
      13'hB48: dout <= 8'b01100011; // 2888 :  99 - 0x63
      13'hB49: dout <= 8'b01100011; // 2889 :  99 - 0x63
      13'hB4A: dout <= 8'b01100011; // 2890 :  99 - 0x63
      13'hB4B: dout <= 8'b01111111; // 2891 : 127 - 0x7f
      13'hB4C: dout <= 8'b01100011; // 2892 :  99 - 0x63
      13'hB4D: dout <= 8'b01100011; // 2893 :  99 - 0x63
      13'hB4E: dout <= 8'b01100011; // 2894 :  99 - 0x63
      13'hB4F: dout <= 8'b00000000; // 2895 :   0 - 0x0
      13'hB50: dout <= 8'b00111111; // 2896 :  63 - 0x3f -- Sprite 0xb5
      13'hB51: dout <= 8'b00001100; // 2897 :  12 - 0xc
      13'hB52: dout <= 8'b00001100; // 2898 :  12 - 0xc
      13'hB53: dout <= 8'b00001100; // 2899 :  12 - 0xc
      13'hB54: dout <= 8'b00001100; // 2900 :  12 - 0xc
      13'hB55: dout <= 8'b00001100; // 2901 :  12 - 0xc
      13'hB56: dout <= 8'b00111111; // 2902 :  63 - 0x3f
      13'hB57: dout <= 8'b00000000; // 2903 :   0 - 0x0
      13'hB58: dout <= 8'b00111111; // 2904 :  63 - 0x3f
      13'hB59: dout <= 8'b00001100; // 2905 :  12 - 0xc
      13'hB5A: dout <= 8'b00001100; // 2906 :  12 - 0xc
      13'hB5B: dout <= 8'b00001100; // 2907 :  12 - 0xc
      13'hB5C: dout <= 8'b00001100; // 2908 :  12 - 0xc
      13'hB5D: dout <= 8'b00001100; // 2909 :  12 - 0xc
      13'hB5E: dout <= 8'b00111111; // 2910 :  63 - 0x3f
      13'hB5F: dout <= 8'b00000000; // 2911 :   0 - 0x0
      13'hB60: dout <= 8'b00000000; // 2912 :   0 - 0x0 -- Sprite 0xb6
      13'hB61: dout <= 8'b00000000; // 2913 :   0 - 0x0
      13'hB62: dout <= 8'b00000000; // 2914 :   0 - 0x0
      13'hB63: dout <= 8'b01111110; // 2915 : 126 - 0x7e
      13'hB64: dout <= 8'b00000000; // 2916 :   0 - 0x0
      13'hB65: dout <= 8'b00000000; // 2917 :   0 - 0x0
      13'hB66: dout <= 8'b00000000; // 2918 :   0 - 0x0
      13'hB67: dout <= 8'b00000000; // 2919 :   0 - 0x0
      13'hB68: dout <= 8'b00000000; // 2920 :   0 - 0x0
      13'hB69: dout <= 8'b00000000; // 2921 :   0 - 0x0
      13'hB6A: dout <= 8'b00000000; // 2922 :   0 - 0x0
      13'hB6B: dout <= 8'b01111110; // 2923 : 126 - 0x7e
      13'hB6C: dout <= 8'b00000000; // 2924 :   0 - 0x0
      13'hB6D: dout <= 8'b00000000; // 2925 :   0 - 0x0
      13'hB6E: dout <= 8'b00000000; // 2926 :   0 - 0x0
      13'hB6F: dout <= 8'b00000000; // 2927 :   0 - 0x0
      13'hB70: dout <= 8'b00111100; // 2928 :  60 - 0x3c -- Sprite 0xb7
      13'hB71: dout <= 8'b01100110; // 2929 : 102 - 0x66
      13'hB72: dout <= 8'b01100000; // 2930 :  96 - 0x60
      13'hB73: dout <= 8'b00111110; // 2931 :  62 - 0x3e
      13'hB74: dout <= 8'b00000011; // 2932 :   3 - 0x3
      13'hB75: dout <= 8'b01100011; // 2933 :  99 - 0x63
      13'hB76: dout <= 8'b00111110; // 2934 :  62 - 0x3e
      13'hB77: dout <= 8'b00000000; // 2935 :   0 - 0x0
      13'hB78: dout <= 8'b00111100; // 2936 :  60 - 0x3c
      13'hB79: dout <= 8'b01100110; // 2937 : 102 - 0x66
      13'hB7A: dout <= 8'b01100000; // 2938 :  96 - 0x60
      13'hB7B: dout <= 8'b00111110; // 2939 :  62 - 0x3e
      13'hB7C: dout <= 8'b00000011; // 2940 :   3 - 0x3
      13'hB7D: dout <= 8'b01100011; // 2941 :  99 - 0x63
      13'hB7E: dout <= 8'b00111110; // 2942 :  62 - 0x3e
      13'hB7F: dout <= 8'b00000000; // 2943 :   0 - 0x0
      13'hB80: dout <= 8'b00011110; // 2944 :  30 - 0x1e -- Sprite 0xb8
      13'hB81: dout <= 8'b00110011; // 2945 :  51 - 0x33
      13'hB82: dout <= 8'b01100000; // 2946 :  96 - 0x60
      13'hB83: dout <= 8'b01100000; // 2947 :  96 - 0x60
      13'hB84: dout <= 8'b01100000; // 2948 :  96 - 0x60
      13'hB85: dout <= 8'b00110011; // 2949 :  51 - 0x33
      13'hB86: dout <= 8'b00011110; // 2950 :  30 - 0x1e
      13'hB87: dout <= 8'b00000000; // 2951 :   0 - 0x0
      13'hB88: dout <= 8'b00011110; // 2952 :  30 - 0x1e
      13'hB89: dout <= 8'b00110011; // 2953 :  51 - 0x33
      13'hB8A: dout <= 8'b01100000; // 2954 :  96 - 0x60
      13'hB8B: dout <= 8'b01100000; // 2955 :  96 - 0x60
      13'hB8C: dout <= 8'b01100000; // 2956 :  96 - 0x60
      13'hB8D: dout <= 8'b00110011; // 2957 :  51 - 0x33
      13'hB8E: dout <= 8'b00011110; // 2958 :  30 - 0x1e
      13'hB8F: dout <= 8'b00000000; // 2959 :   0 - 0x0
      13'hB90: dout <= 8'b00111110; // 2960 :  62 - 0x3e -- Sprite 0xb9
      13'hB91: dout <= 8'b01100011; // 2961 :  99 - 0x63
      13'hB92: dout <= 8'b01100011; // 2962 :  99 - 0x63
      13'hB93: dout <= 8'b01100011; // 2963 :  99 - 0x63
      13'hB94: dout <= 8'b01100011; // 2964 :  99 - 0x63
      13'hB95: dout <= 8'b01100011; // 2965 :  99 - 0x63
      13'hB96: dout <= 8'b00111110; // 2966 :  62 - 0x3e
      13'hB97: dout <= 8'b00000000; // 2967 :   0 - 0x0
      13'hB98: dout <= 8'b00111110; // 2968 :  62 - 0x3e
      13'hB99: dout <= 8'b01100011; // 2969 :  99 - 0x63
      13'hB9A: dout <= 8'b01100011; // 2970 :  99 - 0x63
      13'hB9B: dout <= 8'b01100011; // 2971 :  99 - 0x63
      13'hB9C: dout <= 8'b01100011; // 2972 :  99 - 0x63
      13'hB9D: dout <= 8'b01100011; // 2973 :  99 - 0x63
      13'hB9E: dout <= 8'b00111110; // 2974 :  62 - 0x3e
      13'hB9F: dout <= 8'b00000000; // 2975 :   0 - 0x0
      13'hBA0: dout <= 8'b01111110; // 2976 : 126 - 0x7e -- Sprite 0xba
      13'hBA1: dout <= 8'b01100011; // 2977 :  99 - 0x63
      13'hBA2: dout <= 8'b01100011; // 2978 :  99 - 0x63
      13'hBA3: dout <= 8'b01100111; // 2979 : 103 - 0x67
      13'hBA4: dout <= 8'b01111100; // 2980 : 124 - 0x7c
      13'hBA5: dout <= 8'b01101110; // 2981 : 110 - 0x6e
      13'hBA6: dout <= 8'b01100111; // 2982 : 103 - 0x67
      13'hBA7: dout <= 8'b00000000; // 2983 :   0 - 0x0
      13'hBA8: dout <= 8'b01111110; // 2984 : 126 - 0x7e
      13'hBA9: dout <= 8'b01100011; // 2985 :  99 - 0x63
      13'hBAA: dout <= 8'b01100011; // 2986 :  99 - 0x63
      13'hBAB: dout <= 8'b01100111; // 2987 : 103 - 0x67
      13'hBAC: dout <= 8'b01111100; // 2988 : 124 - 0x7c
      13'hBAD: dout <= 8'b01101110; // 2989 : 110 - 0x6e
      13'hBAE: dout <= 8'b01100111; // 2990 : 103 - 0x67
      13'hBAF: dout <= 8'b00000000; // 2991 :   0 - 0x0
      13'hBB0: dout <= 8'b01111111; // 2992 : 127 - 0x7f -- Sprite 0xbb
      13'hBB1: dout <= 8'b01100000; // 2993 :  96 - 0x60
      13'hBB2: dout <= 8'b01100000; // 2994 :  96 - 0x60
      13'hBB3: dout <= 8'b01111110; // 2995 : 126 - 0x7e
      13'hBB4: dout <= 8'b01100000; // 2996 :  96 - 0x60
      13'hBB5: dout <= 8'b01100000; // 2997 :  96 - 0x60
      13'hBB6: dout <= 8'b01111111; // 2998 : 127 - 0x7f
      13'hBB7: dout <= 8'b00000000; // 2999 :   0 - 0x0
      13'hBB8: dout <= 8'b01111111; // 3000 : 127 - 0x7f
      13'hBB9: dout <= 8'b01100000; // 3001 :  96 - 0x60
      13'hBBA: dout <= 8'b01100000; // 3002 :  96 - 0x60
      13'hBBB: dout <= 8'b01111110; // 3003 : 126 - 0x7e
      13'hBBC: dout <= 8'b01100000; // 3004 :  96 - 0x60
      13'hBBD: dout <= 8'b01100000; // 3005 :  96 - 0x60
      13'hBBE: dout <= 8'b01111111; // 3006 : 127 - 0x7f
      13'hBBF: dout <= 8'b00000000; // 3007 :   0 - 0x0
      13'hBC0: dout <= 8'b00000000; // 3008 :   0 - 0x0 -- Sprite 0xbc
      13'hBC1: dout <= 8'b00100010; // 3009 :  34 - 0x22
      13'hBC2: dout <= 8'b01100101; // 3010 : 101 - 0x65
      13'hBC3: dout <= 8'b00100101; // 3011 :  37 - 0x25
      13'hBC4: dout <= 8'b00100101; // 3012 :  37 - 0x25
      13'hBC5: dout <= 8'b01110010; // 3013 : 114 - 0x72
      13'hBC6: dout <= 8'b00000000; // 3014 :   0 - 0x0
      13'hBC7: dout <= 8'b00000000; // 3015 :   0 - 0x0
      13'hBC8: dout <= 8'b00000000; // 3016 :   0 - 0x0
      13'hBC9: dout <= 8'b00000000; // 3017 :   0 - 0x0
      13'hBCA: dout <= 8'b00000000; // 3018 :   0 - 0x0
      13'hBCB: dout <= 8'b00000000; // 3019 :   0 - 0x0
      13'hBCC: dout <= 8'b00000000; // 3020 :   0 - 0x0
      13'hBCD: dout <= 8'b00000000; // 3021 :   0 - 0x0
      13'hBCE: dout <= 8'b00000000; // 3022 :   0 - 0x0
      13'hBCF: dout <= 8'b00000000; // 3023 :   0 - 0x0
      13'hBD0: dout <= 8'b00000000; // 3024 :   0 - 0x0 -- Sprite 0xbd
      13'hBD1: dout <= 8'b01110010; // 3025 : 114 - 0x72
      13'hBD2: dout <= 8'b01000101; // 3026 :  69 - 0x45
      13'hBD3: dout <= 8'b01100101; // 3027 : 101 - 0x65
      13'hBD4: dout <= 8'b00010101; // 3028 :  21 - 0x15
      13'hBD5: dout <= 8'b01100010; // 3029 :  98 - 0x62
      13'hBD6: dout <= 8'b00000000; // 3030 :   0 - 0x0
      13'hBD7: dout <= 8'b00000000; // 3031 :   0 - 0x0
      13'hBD8: dout <= 8'b00000000; // 3032 :   0 - 0x0
      13'hBD9: dout <= 8'b00000000; // 3033 :   0 - 0x0
      13'hBDA: dout <= 8'b00000000; // 3034 :   0 - 0x0
      13'hBDB: dout <= 8'b00000000; // 3035 :   0 - 0x0
      13'hBDC: dout <= 8'b00000000; // 3036 :   0 - 0x0
      13'hBDD: dout <= 8'b00000000; // 3037 :   0 - 0x0
      13'hBDE: dout <= 8'b00000000; // 3038 :   0 - 0x0
      13'hBDF: dout <= 8'b00000000; // 3039 :   0 - 0x0
      13'hBE0: dout <= 8'b00000000; // 3040 :   0 - 0x0 -- Sprite 0xbe
      13'hBE1: dout <= 8'b01100111; // 3041 : 103 - 0x67
      13'hBE2: dout <= 8'b01010010; // 3042 :  82 - 0x52
      13'hBE3: dout <= 8'b01100010; // 3043 :  98 - 0x62
      13'hBE4: dout <= 8'b01000010; // 3044 :  66 - 0x42
      13'hBE5: dout <= 8'b01000010; // 3045 :  66 - 0x42
      13'hBE6: dout <= 8'b00000000; // 3046 :   0 - 0x0
      13'hBE7: dout <= 8'b00000000; // 3047 :   0 - 0x0
      13'hBE8: dout <= 8'b00000000; // 3048 :   0 - 0x0
      13'hBE9: dout <= 8'b00000000; // 3049 :   0 - 0x0
      13'hBEA: dout <= 8'b00000000; // 3050 :   0 - 0x0
      13'hBEB: dout <= 8'b00000000; // 3051 :   0 - 0x0
      13'hBEC: dout <= 8'b00000000; // 3052 :   0 - 0x0
      13'hBED: dout <= 8'b00000000; // 3053 :   0 - 0x0
      13'hBEE: dout <= 8'b00000000; // 3054 :   0 - 0x0
      13'hBEF: dout <= 8'b00000000; // 3055 :   0 - 0x0
      13'hBF0: dout <= 8'b00000000; // 3056 :   0 - 0x0 -- Sprite 0xbf
      13'hBF1: dout <= 8'b01100000; // 3057 :  96 - 0x60
      13'hBF2: dout <= 8'b10000000; // 3058 : 128 - 0x80
      13'hBF3: dout <= 8'b01000000; // 3059 :  64 - 0x40
      13'hBF4: dout <= 8'b00100000; // 3060 :  32 - 0x20
      13'hBF5: dout <= 8'b11000110; // 3061 : 198 - 0xc6
      13'hBF6: dout <= 8'b00000000; // 3062 :   0 - 0x0
      13'hBF7: dout <= 8'b00000000; // 3063 :   0 - 0x0
      13'hBF8: dout <= 8'b00000000; // 3064 :   0 - 0x0
      13'hBF9: dout <= 8'b00000000; // 3065 :   0 - 0x0
      13'hBFA: dout <= 8'b00000000; // 3066 :   0 - 0x0
      13'hBFB: dout <= 8'b00000000; // 3067 :   0 - 0x0
      13'hBFC: dout <= 8'b00000000; // 3068 :   0 - 0x0
      13'hBFD: dout <= 8'b00000000; // 3069 :   0 - 0x0
      13'hBFE: dout <= 8'b00000000; // 3070 :   0 - 0x0
      13'hBFF: dout <= 8'b00000000; // 3071 :   0 - 0x0
      13'hC00: dout <= 8'b01100011; // 3072 :  99 - 0x63 -- Sprite 0xc0
      13'hC01: dout <= 8'b01100110; // 3073 : 102 - 0x66
      13'hC02: dout <= 8'b01101100; // 3074 : 108 - 0x6c
      13'hC03: dout <= 8'b01111000; // 3075 : 120 - 0x78
      13'hC04: dout <= 8'b01111100; // 3076 : 124 - 0x7c
      13'hC05: dout <= 8'b01100110; // 3077 : 102 - 0x66
      13'hC06: dout <= 8'b01100011; // 3078 :  99 - 0x63
      13'hC07: dout <= 8'b00000000; // 3079 :   0 - 0x0
      13'hC08: dout <= 8'b01100011; // 3080 :  99 - 0x63
      13'hC09: dout <= 8'b01100110; // 3081 : 102 - 0x66
      13'hC0A: dout <= 8'b01101100; // 3082 : 108 - 0x6c
      13'hC0B: dout <= 8'b01111000; // 3083 : 120 - 0x78
      13'hC0C: dout <= 8'b01111100; // 3084 : 124 - 0x7c
      13'hC0D: dout <= 8'b01100110; // 3085 : 102 - 0x66
      13'hC0E: dout <= 8'b01100011; // 3086 :  99 - 0x63
      13'hC0F: dout <= 8'b00000000; // 3087 :   0 - 0x0
      13'hC10: dout <= 8'b00111111; // 3088 :  63 - 0x3f -- Sprite 0xc1
      13'hC11: dout <= 8'b00001100; // 3089 :  12 - 0xc
      13'hC12: dout <= 8'b00001100; // 3090 :  12 - 0xc
      13'hC13: dout <= 8'b00001100; // 3091 :  12 - 0xc
      13'hC14: dout <= 8'b00001100; // 3092 :  12 - 0xc
      13'hC15: dout <= 8'b00001100; // 3093 :  12 - 0xc
      13'hC16: dout <= 8'b00111111; // 3094 :  63 - 0x3f
      13'hC17: dout <= 8'b00000000; // 3095 :   0 - 0x0
      13'hC18: dout <= 8'b00111111; // 3096 :  63 - 0x3f
      13'hC19: dout <= 8'b00001100; // 3097 :  12 - 0xc
      13'hC1A: dout <= 8'b00001100; // 3098 :  12 - 0xc
      13'hC1B: dout <= 8'b00001100; // 3099 :  12 - 0xc
      13'hC1C: dout <= 8'b00001100; // 3100 :  12 - 0xc
      13'hC1D: dout <= 8'b00001100; // 3101 :  12 - 0xc
      13'hC1E: dout <= 8'b00111111; // 3102 :  63 - 0x3f
      13'hC1F: dout <= 8'b00000000; // 3103 :   0 - 0x0
      13'hC20: dout <= 8'b01100011; // 3104 :  99 - 0x63 -- Sprite 0xc2
      13'hC21: dout <= 8'b01110111; // 3105 : 119 - 0x77
      13'hC22: dout <= 8'b01111111; // 3106 : 127 - 0x7f
      13'hC23: dout <= 8'b01111111; // 3107 : 127 - 0x7f
      13'hC24: dout <= 8'b01101011; // 3108 : 107 - 0x6b
      13'hC25: dout <= 8'b01100011; // 3109 :  99 - 0x63
      13'hC26: dout <= 8'b01100011; // 3110 :  99 - 0x63
      13'hC27: dout <= 8'b00000000; // 3111 :   0 - 0x0
      13'hC28: dout <= 8'b01100011; // 3112 :  99 - 0x63
      13'hC29: dout <= 8'b01110111; // 3113 : 119 - 0x77
      13'hC2A: dout <= 8'b01111111; // 3114 : 127 - 0x7f
      13'hC2B: dout <= 8'b01111111; // 3115 : 127 - 0x7f
      13'hC2C: dout <= 8'b01101011; // 3116 : 107 - 0x6b
      13'hC2D: dout <= 8'b01100011; // 3117 :  99 - 0x63
      13'hC2E: dout <= 8'b01100011; // 3118 :  99 - 0x63
      13'hC2F: dout <= 8'b00000000; // 3119 :   0 - 0x0
      13'hC30: dout <= 8'b00011100; // 3120 :  28 - 0x1c -- Sprite 0xc3
      13'hC31: dout <= 8'b00110110; // 3121 :  54 - 0x36
      13'hC32: dout <= 8'b01100011; // 3122 :  99 - 0x63
      13'hC33: dout <= 8'b01100011; // 3123 :  99 - 0x63
      13'hC34: dout <= 8'b01111111; // 3124 : 127 - 0x7f
      13'hC35: dout <= 8'b01100011; // 3125 :  99 - 0x63
      13'hC36: dout <= 8'b01100011; // 3126 :  99 - 0x63
      13'hC37: dout <= 8'b00000000; // 3127 :   0 - 0x0
      13'hC38: dout <= 8'b00011100; // 3128 :  28 - 0x1c
      13'hC39: dout <= 8'b00110110; // 3129 :  54 - 0x36
      13'hC3A: dout <= 8'b01100011; // 3130 :  99 - 0x63
      13'hC3B: dout <= 8'b01100011; // 3131 :  99 - 0x63
      13'hC3C: dout <= 8'b01111111; // 3132 : 127 - 0x7f
      13'hC3D: dout <= 8'b01100011; // 3133 :  99 - 0x63
      13'hC3E: dout <= 8'b01100011; // 3134 :  99 - 0x63
      13'hC3F: dout <= 8'b00000000; // 3135 :   0 - 0x0
      13'hC40: dout <= 8'b00011111; // 3136 :  31 - 0x1f -- Sprite 0xc4
      13'hC41: dout <= 8'b00110000; // 3137 :  48 - 0x30
      13'hC42: dout <= 8'b01100000; // 3138 :  96 - 0x60
      13'hC43: dout <= 8'b01100111; // 3139 : 103 - 0x67
      13'hC44: dout <= 8'b01100011; // 3140 :  99 - 0x63
      13'hC45: dout <= 8'b00110011; // 3141 :  51 - 0x33
      13'hC46: dout <= 8'b00011111; // 3142 :  31 - 0x1f
      13'hC47: dout <= 8'b00000000; // 3143 :   0 - 0x0
      13'hC48: dout <= 8'b00011111; // 3144 :  31 - 0x1f
      13'hC49: dout <= 8'b00110000; // 3145 :  48 - 0x30
      13'hC4A: dout <= 8'b01100000; // 3146 :  96 - 0x60
      13'hC4B: dout <= 8'b01100111; // 3147 : 103 - 0x67
      13'hC4C: dout <= 8'b01100011; // 3148 :  99 - 0x63
      13'hC4D: dout <= 8'b00110011; // 3149 :  51 - 0x33
      13'hC4E: dout <= 8'b00011111; // 3150 :  31 - 0x1f
      13'hC4F: dout <= 8'b00000000; // 3151 :   0 - 0x0
      13'hC50: dout <= 8'b01100011; // 3152 :  99 - 0x63 -- Sprite 0xc5
      13'hC51: dout <= 8'b01100011; // 3153 :  99 - 0x63
      13'hC52: dout <= 8'b01100011; // 3154 :  99 - 0x63
      13'hC53: dout <= 8'b01100011; // 3155 :  99 - 0x63
      13'hC54: dout <= 8'b01100011; // 3156 :  99 - 0x63
      13'hC55: dout <= 8'b01100011; // 3157 :  99 - 0x63
      13'hC56: dout <= 8'b00111110; // 3158 :  62 - 0x3e
      13'hC57: dout <= 8'b00000000; // 3159 :   0 - 0x0
      13'hC58: dout <= 8'b01100011; // 3160 :  99 - 0x63
      13'hC59: dout <= 8'b01100011; // 3161 :  99 - 0x63
      13'hC5A: dout <= 8'b01100011; // 3162 :  99 - 0x63
      13'hC5B: dout <= 8'b01100011; // 3163 :  99 - 0x63
      13'hC5C: dout <= 8'b01100011; // 3164 :  99 - 0x63
      13'hC5D: dout <= 8'b01100011; // 3165 :  99 - 0x63
      13'hC5E: dout <= 8'b00111110; // 3166 :  62 - 0x3e
      13'hC5F: dout <= 8'b00000000; // 3167 :   0 - 0x0
      13'hC60: dout <= 8'b01111110; // 3168 : 126 - 0x7e -- Sprite 0xc6
      13'hC61: dout <= 8'b01100011; // 3169 :  99 - 0x63
      13'hC62: dout <= 8'b01100011; // 3170 :  99 - 0x63
      13'hC63: dout <= 8'b01100111; // 3171 : 103 - 0x67
      13'hC64: dout <= 8'b01111100; // 3172 : 124 - 0x7c
      13'hC65: dout <= 8'b01101110; // 3173 : 110 - 0x6e
      13'hC66: dout <= 8'b01100111; // 3174 : 103 - 0x67
      13'hC67: dout <= 8'b00000000; // 3175 :   0 - 0x0
      13'hC68: dout <= 8'b01111110; // 3176 : 126 - 0x7e
      13'hC69: dout <= 8'b01100011; // 3177 :  99 - 0x63
      13'hC6A: dout <= 8'b01100011; // 3178 :  99 - 0x63
      13'hC6B: dout <= 8'b01100111; // 3179 : 103 - 0x67
      13'hC6C: dout <= 8'b01111100; // 3180 : 124 - 0x7c
      13'hC6D: dout <= 8'b01101110; // 3181 : 110 - 0x6e
      13'hC6E: dout <= 8'b01100111; // 3182 : 103 - 0x67
      13'hC6F: dout <= 8'b00000000; // 3183 :   0 - 0x0
      13'hC70: dout <= 8'b01111111; // 3184 : 127 - 0x7f -- Sprite 0xc7
      13'hC71: dout <= 8'b01100000; // 3185 :  96 - 0x60
      13'hC72: dout <= 8'b01100000; // 3186 :  96 - 0x60
      13'hC73: dout <= 8'b01111110; // 3187 : 126 - 0x7e
      13'hC74: dout <= 8'b01100000; // 3188 :  96 - 0x60
      13'hC75: dout <= 8'b01100000; // 3189 :  96 - 0x60
      13'hC76: dout <= 8'b01111111; // 3190 : 127 - 0x7f
      13'hC77: dout <= 8'b00000000; // 3191 :   0 - 0x0
      13'hC78: dout <= 8'b01111111; // 3192 : 127 - 0x7f
      13'hC79: dout <= 8'b01100000; // 3193 :  96 - 0x60
      13'hC7A: dout <= 8'b01100000; // 3194 :  96 - 0x60
      13'hC7B: dout <= 8'b01111110; // 3195 : 126 - 0x7e
      13'hC7C: dout <= 8'b01100000; // 3196 :  96 - 0x60
      13'hC7D: dout <= 8'b01100000; // 3197 :  96 - 0x60
      13'hC7E: dout <= 8'b01111111; // 3198 : 127 - 0x7f
      13'hC7F: dout <= 8'b00000000; // 3199 :   0 - 0x0
      13'hC80: dout <= 8'b00110110; // 3200 :  54 - 0x36 -- Sprite 0xc8
      13'hC81: dout <= 8'b00110110; // 3201 :  54 - 0x36
      13'hC82: dout <= 8'b00010010; // 3202 :  18 - 0x12
      13'hC83: dout <= 8'b00000000; // 3203 :   0 - 0x0
      13'hC84: dout <= 8'b00000000; // 3204 :   0 - 0x0
      13'hC85: dout <= 8'b00000000; // 3205 :   0 - 0x0
      13'hC86: dout <= 8'b00000000; // 3206 :   0 - 0x0
      13'hC87: dout <= 8'b00000000; // 3207 :   0 - 0x0
      13'hC88: dout <= 8'b00110110; // 3208 :  54 - 0x36
      13'hC89: dout <= 8'b00110110; // 3209 :  54 - 0x36
      13'hC8A: dout <= 8'b00010010; // 3210 :  18 - 0x12
      13'hC8B: dout <= 8'b00000000; // 3211 :   0 - 0x0
      13'hC8C: dout <= 8'b00000000; // 3212 :   0 - 0x0
      13'hC8D: dout <= 8'b00000000; // 3213 :   0 - 0x0
      13'hC8E: dout <= 8'b00000000; // 3214 :   0 - 0x0
      13'hC8F: dout <= 8'b00000000; // 3215 :   0 - 0x0
      13'hC90: dout <= 8'b00111110; // 3216 :  62 - 0x3e -- Sprite 0xc9
      13'hC91: dout <= 8'b01100011; // 3217 :  99 - 0x63
      13'hC92: dout <= 8'b01100011; // 3218 :  99 - 0x63
      13'hC93: dout <= 8'b01100011; // 3219 :  99 - 0x63
      13'hC94: dout <= 8'b01100011; // 3220 :  99 - 0x63
      13'hC95: dout <= 8'b01100011; // 3221 :  99 - 0x63
      13'hC96: dout <= 8'b00111110; // 3222 :  62 - 0x3e
      13'hC97: dout <= 8'b00000000; // 3223 :   0 - 0x0
      13'hC98: dout <= 8'b00111110; // 3224 :  62 - 0x3e
      13'hC99: dout <= 8'b01100011; // 3225 :  99 - 0x63
      13'hC9A: dout <= 8'b01100011; // 3226 :  99 - 0x63
      13'hC9B: dout <= 8'b01100011; // 3227 :  99 - 0x63
      13'hC9C: dout <= 8'b01100011; // 3228 :  99 - 0x63
      13'hC9D: dout <= 8'b01100011; // 3229 :  99 - 0x63
      13'hC9E: dout <= 8'b00111110; // 3230 :  62 - 0x3e
      13'hC9F: dout <= 8'b00000000; // 3231 :   0 - 0x0
      13'hCA0: dout <= 8'b00111100; // 3232 :  60 - 0x3c -- Sprite 0xca
      13'hCA1: dout <= 8'b01100110; // 3233 : 102 - 0x66
      13'hCA2: dout <= 8'b01100000; // 3234 :  96 - 0x60
      13'hCA3: dout <= 8'b00111110; // 3235 :  62 - 0x3e
      13'hCA4: dout <= 8'b00000011; // 3236 :   3 - 0x3
      13'hCA5: dout <= 8'b01100011; // 3237 :  99 - 0x63
      13'hCA6: dout <= 8'b00111110; // 3238 :  62 - 0x3e
      13'hCA7: dout <= 8'b00000000; // 3239 :   0 - 0x0
      13'hCA8: dout <= 8'b00111100; // 3240 :  60 - 0x3c
      13'hCA9: dout <= 8'b01100110; // 3241 : 102 - 0x66
      13'hCAA: dout <= 8'b01100000; // 3242 :  96 - 0x60
      13'hCAB: dout <= 8'b00111110; // 3243 :  62 - 0x3e
      13'hCAC: dout <= 8'b00000011; // 3244 :   3 - 0x3
      13'hCAD: dout <= 8'b01100011; // 3245 :  99 - 0x63
      13'hCAE: dout <= 8'b00111110; // 3246 :  62 - 0x3e
      13'hCAF: dout <= 8'b00000000; // 3247 :   0 - 0x0
      13'hCB0: dout <= 8'b00000000; // 3248 :   0 - 0x0 -- Sprite 0xcb
      13'hCB1: dout <= 8'b00000000; // 3249 :   0 - 0x0
      13'hCB2: dout <= 8'b00000000; // 3250 :   0 - 0x0
      13'hCB3: dout <= 8'b00000000; // 3251 :   0 - 0x0
      13'hCB4: dout <= 8'b00000000; // 3252 :   0 - 0x0
      13'hCB5: dout <= 8'b00000000; // 3253 :   0 - 0x0
      13'hCB6: dout <= 8'b00000000; // 3254 :   0 - 0x0
      13'hCB7: dout <= 8'b00000000; // 3255 :   0 - 0x0
      13'hCB8: dout <= 8'b00000000; // 3256 :   0 - 0x0
      13'hCB9: dout <= 8'b00111000; // 3257 :  56 - 0x38
      13'hCBA: dout <= 8'b01111100; // 3258 : 124 - 0x7c
      13'hCBB: dout <= 8'b11111110; // 3259 : 254 - 0xfe
      13'hCBC: dout <= 8'b11111110; // 3260 : 254 - 0xfe
      13'hCBD: dout <= 8'b11111110; // 3261 : 254 - 0xfe
      13'hCBE: dout <= 8'b01111100; // 3262 : 124 - 0x7c
      13'hCBF: dout <= 8'b00111000; // 3263 :  56 - 0x38
      13'hCC0: dout <= 8'b00000000; // 3264 :   0 - 0x0 -- Sprite 0xcc
      13'hCC1: dout <= 8'b00000000; // 3265 :   0 - 0x0
      13'hCC2: dout <= 8'b00000000; // 3266 :   0 - 0x0
      13'hCC3: dout <= 8'b00000000; // 3267 :   0 - 0x0
      13'hCC4: dout <= 8'b00000000; // 3268 :   0 - 0x0
      13'hCC5: dout <= 8'b00000000; // 3269 :   0 - 0x0
      13'hCC6: dout <= 8'b00000000; // 3270 :   0 - 0x0
      13'hCC7: dout <= 8'b00000000; // 3271 :   0 - 0x0
      13'hCC8: dout <= 8'b00000000; // 3272 :   0 - 0x0
      13'hCC9: dout <= 8'b00000000; // 3273 :   0 - 0x0
      13'hCCA: dout <= 8'b00000000; // 3274 :   0 - 0x0
      13'hCCB: dout <= 8'b00000000; // 3275 :   0 - 0x0
      13'hCCC: dout <= 8'b00000000; // 3276 :   0 - 0x0
      13'hCCD: dout <= 8'b00000000; // 3277 :   0 - 0x0
      13'hCCE: dout <= 8'b00000000; // 3278 :   0 - 0x0
      13'hCCF: dout <= 8'b00000000; // 3279 :   0 - 0x0
      13'hCD0: dout <= 8'b00000000; // 3280 :   0 - 0x0 -- Sprite 0xcd
      13'hCD1: dout <= 8'b00000000; // 3281 :   0 - 0x0
      13'hCD2: dout <= 8'b00000000; // 3282 :   0 - 0x0
      13'hCD3: dout <= 8'b00000000; // 3283 :   0 - 0x0
      13'hCD4: dout <= 8'b00000000; // 3284 :   0 - 0x0
      13'hCD5: dout <= 8'b00000000; // 3285 :   0 - 0x0
      13'hCD6: dout <= 8'b00000000; // 3286 :   0 - 0x0
      13'hCD7: dout <= 8'b00000000; // 3287 :   0 - 0x0
      13'hCD8: dout <= 8'b00000000; // 3288 :   0 - 0x0
      13'hCD9: dout <= 8'b00000000; // 3289 :   0 - 0x0
      13'hCDA: dout <= 8'b00000000; // 3290 :   0 - 0x0
      13'hCDB: dout <= 8'b00000000; // 3291 :   0 - 0x0
      13'hCDC: dout <= 8'b00000000; // 3292 :   0 - 0x0
      13'hCDD: dout <= 8'b00000000; // 3293 :   0 - 0x0
      13'hCDE: dout <= 8'b00000000; // 3294 :   0 - 0x0
      13'hCDF: dout <= 8'b00000000; // 3295 :   0 - 0x0
      13'hCE0: dout <= 8'b00000000; // 3296 :   0 - 0x0 -- Sprite 0xce
      13'hCE1: dout <= 8'b00000000; // 3297 :   0 - 0x0
      13'hCE2: dout <= 8'b00000000; // 3298 :   0 - 0x0
      13'hCE3: dout <= 8'b00000000; // 3299 :   0 - 0x0
      13'hCE4: dout <= 8'b00000000; // 3300 :   0 - 0x0
      13'hCE5: dout <= 8'b00000000; // 3301 :   0 - 0x0
      13'hCE6: dout <= 8'b00000000; // 3302 :   0 - 0x0
      13'hCE7: dout <= 8'b00000000; // 3303 :   0 - 0x0
      13'hCE8: dout <= 8'b00000000; // 3304 :   0 - 0x0
      13'hCE9: dout <= 8'b00000000; // 3305 :   0 - 0x0
      13'hCEA: dout <= 8'b00000000; // 3306 :   0 - 0x0
      13'hCEB: dout <= 8'b00000000; // 3307 :   0 - 0x0
      13'hCEC: dout <= 8'b00000000; // 3308 :   0 - 0x0
      13'hCED: dout <= 8'b00000000; // 3309 :   0 - 0x0
      13'hCEE: dout <= 8'b00000000; // 3310 :   0 - 0x0
      13'hCEF: dout <= 8'b00000000; // 3311 :   0 - 0x0
      13'hCF0: dout <= 8'b00000000; // 3312 :   0 - 0x0 -- Sprite 0xcf
      13'hCF1: dout <= 8'b00000000; // 3313 :   0 - 0x0
      13'hCF2: dout <= 8'b00000000; // 3314 :   0 - 0x0
      13'hCF3: dout <= 8'b00000000; // 3315 :   0 - 0x0
      13'hCF4: dout <= 8'b00000000; // 3316 :   0 - 0x0
      13'hCF5: dout <= 8'b00000000; // 3317 :   0 - 0x0
      13'hCF6: dout <= 8'b00000000; // 3318 :   0 - 0x0
      13'hCF7: dout <= 8'b00000000; // 3319 :   0 - 0x0
      13'hCF8: dout <= 8'b00000000; // 3320 :   0 - 0x0
      13'hCF9: dout <= 8'b00000000; // 3321 :   0 - 0x0
      13'hCFA: dout <= 8'b00000000; // 3322 :   0 - 0x0
      13'hCFB: dout <= 8'b00000000; // 3323 :   0 - 0x0
      13'hCFC: dout <= 8'b00000000; // 3324 :   0 - 0x0
      13'hCFD: dout <= 8'b00000000; // 3325 :   0 - 0x0
      13'hCFE: dout <= 8'b00000000; // 3326 :   0 - 0x0
      13'hCFF: dout <= 8'b00000000; // 3327 :   0 - 0x0
      13'hD00: dout <= 8'b01000111; // 3328 :  71 - 0x47 -- Sprite 0xd0
      13'hD01: dout <= 8'b01000111; // 3329 :  71 - 0x47
      13'hD02: dout <= 8'b00001111; // 3330 :  15 - 0xf
      13'hD03: dout <= 8'b00001111; // 3331 :  15 - 0xf
      13'hD04: dout <= 8'b00011111; // 3332 :  31 - 0x1f
      13'hD05: dout <= 8'b00011111; // 3333 :  31 - 0x1f
      13'hD06: dout <= 8'b00111111; // 3334 :  63 - 0x3f
      13'hD07: dout <= 8'b00111111; // 3335 :  63 - 0x3f
      13'hD08: dout <= 8'b00010111; // 3336 :  23 - 0x17
      13'hD09: dout <= 8'b00010111; // 3337 :  23 - 0x17
      13'hD0A: dout <= 8'b00101111; // 3338 :  47 - 0x2f
      13'hD0B: dout <= 8'b00101111; // 3339 :  47 - 0x2f
      13'hD0C: dout <= 8'b01011111; // 3340 :  95 - 0x5f
      13'hD0D: dout <= 8'b01011111; // 3341 :  95 - 0x5f
      13'hD0E: dout <= 8'b00111111; // 3342 :  63 - 0x3f
      13'hD0F: dout <= 8'b00111111; // 3343 :  63 - 0x3f
      13'hD10: dout <= 8'b11111111; // 3344 : 255 - 0xff -- Sprite 0xd1
      13'hD11: dout <= 8'b11001111; // 3345 : 207 - 0xcf
      13'hD12: dout <= 8'b11001111; // 3346 : 207 - 0xcf
      13'hD13: dout <= 8'b11111011; // 3347 : 251 - 0xfb
      13'hD14: dout <= 8'b11110111; // 3348 : 247 - 0xf7
      13'hD15: dout <= 8'b11100111; // 3349 : 231 - 0xe7
      13'hD16: dout <= 8'b11111111; // 3350 : 255 - 0xff
      13'hD17: dout <= 8'b11111111; // 3351 : 255 - 0xff
      13'hD18: dout <= 8'b11111111; // 3352 : 255 - 0xff
      13'hD19: dout <= 8'b11001111; // 3353 : 207 - 0xcf
      13'hD1A: dout <= 8'b11001111; // 3354 : 207 - 0xcf
      13'hD1B: dout <= 8'b11111011; // 3355 : 251 - 0xfb
      13'hD1C: dout <= 8'b11110111; // 3356 : 247 - 0xf7
      13'hD1D: dout <= 8'b11100111; // 3357 : 231 - 0xe7
      13'hD1E: dout <= 8'b11111111; // 3358 : 255 - 0xff
      13'hD1F: dout <= 8'b11111111; // 3359 : 255 - 0xff
      13'hD20: dout <= 8'b00011000; // 3360 :  24 - 0x18 -- Sprite 0xd2
      13'hD21: dout <= 8'b00001000; // 3361 :   8 - 0x8
      13'hD22: dout <= 8'b10001000; // 3362 : 136 - 0x88
      13'hD23: dout <= 8'b10000000; // 3363 : 128 - 0x80
      13'hD24: dout <= 8'b01000000; // 3364 :  64 - 0x40
      13'hD25: dout <= 8'b01000000; // 3365 :  64 - 0x40
      13'hD26: dout <= 8'b10100000; // 3366 : 160 - 0xa0
      13'hD27: dout <= 8'b10100000; // 3367 : 160 - 0xa0
      13'hD28: dout <= 8'b01000010; // 3368 :  66 - 0x42
      13'hD29: dout <= 8'b01100010; // 3369 :  98 - 0x62
      13'hD2A: dout <= 8'b10100010; // 3370 : 162 - 0xa2
      13'hD2B: dout <= 8'b10110010; // 3371 : 178 - 0xb2
      13'hD2C: dout <= 8'b01010010; // 3372 :  82 - 0x52
      13'hD2D: dout <= 8'b01011010; // 3373 :  90 - 0x5a
      13'hD2E: dout <= 8'b10101010; // 3374 : 170 - 0xaa
      13'hD2F: dout <= 8'b10101100; // 3375 : 172 - 0xac
      13'hD30: dout <= 8'b11111111; // 3376 : 255 - 0xff -- Sprite 0xd3
      13'hD31: dout <= 8'b11111111; // 3377 : 255 - 0xff
      13'hD32: dout <= 8'b11111111; // 3378 : 255 - 0xff
      13'hD33: dout <= 8'b11111111; // 3379 : 255 - 0xff
      13'hD34: dout <= 8'b11111101; // 3380 : 253 - 0xfd
      13'hD35: dout <= 8'b11111101; // 3381 : 253 - 0xfd
      13'hD36: dout <= 8'b11111101; // 3382 : 253 - 0xfd
      13'hD37: dout <= 8'b11111101; // 3383 : 253 - 0xfd
      13'hD38: dout <= 8'b11111111; // 3384 : 255 - 0xff
      13'hD39: dout <= 8'b11111111; // 3385 : 255 - 0xff
      13'hD3A: dout <= 8'b11111111; // 3386 : 255 - 0xff
      13'hD3B: dout <= 8'b11111111; // 3387 : 255 - 0xff
      13'hD3C: dout <= 8'b11111101; // 3388 : 253 - 0xfd
      13'hD3D: dout <= 8'b11111101; // 3389 : 253 - 0xfd
      13'hD3E: dout <= 8'b11111101; // 3390 : 253 - 0xfd
      13'hD3F: dout <= 8'b11111101; // 3391 : 253 - 0xfd
      13'hD40: dout <= 8'b11000111; // 3392 : 199 - 0xc7 -- Sprite 0xd4
      13'hD41: dout <= 8'b11110111; // 3393 : 247 - 0xf7
      13'hD42: dout <= 8'b11110000; // 3394 : 240 - 0xf0
      13'hD43: dout <= 8'b11111000; // 3395 : 248 - 0xf8
      13'hD44: dout <= 8'b11111000; // 3396 : 248 - 0xf8
      13'hD45: dout <= 8'b11111111; // 3397 : 255 - 0xff
      13'hD46: dout <= 8'b11111111; // 3398 : 255 - 0xff
      13'hD47: dout <= 8'b11111111; // 3399 : 255 - 0xff
      13'hD48: dout <= 8'b00000111; // 3400 :   7 - 0x7
      13'hD49: dout <= 8'b00000111; // 3401 :   7 - 0x7
      13'hD4A: dout <= 8'b00000000; // 3402 :   0 - 0x0
      13'hD4B: dout <= 8'b00000011; // 3403 :   3 - 0x3
      13'hD4C: dout <= 8'b00000000; // 3404 :   0 - 0x0
      13'hD4D: dout <= 8'b00000000; // 3405 :   0 - 0x0
      13'hD4E: dout <= 8'b00000000; // 3406 :   0 - 0x0
      13'hD4F: dout <= 8'b00000000; // 3407 :   0 - 0x0
      13'hD50: dout <= 8'b11111000; // 3408 : 248 - 0xf8 -- Sprite 0xd5
      13'hD51: dout <= 8'b11111000; // 3409 : 248 - 0xf8
      13'hD52: dout <= 8'b00000000; // 3410 :   0 - 0x0
      13'hD53: dout <= 8'b00000000; // 3411 :   0 - 0x0
      13'hD54: dout <= 8'b00000000; // 3412 :   0 - 0x0
      13'hD55: dout <= 8'b11111111; // 3413 : 255 - 0xff
      13'hD56: dout <= 8'b11111111; // 3414 : 255 - 0xff
      13'hD57: dout <= 8'b11111111; // 3415 : 255 - 0xff
      13'hD58: dout <= 8'b11111010; // 3416 : 250 - 0xfa
      13'hD59: dout <= 8'b11111010; // 3417 : 250 - 0xfa
      13'hD5A: dout <= 8'b00000010; // 3418 :   2 - 0x2
      13'hD5B: dout <= 8'b11111110; // 3419 : 254 - 0xfe
      13'hD5C: dout <= 8'b00000000; // 3420 :   0 - 0x0
      13'hD5D: dout <= 8'b00000000; // 3421 :   0 - 0x0
      13'hD5E: dout <= 8'b00000000; // 3422 :   0 - 0x0
      13'hD5F: dout <= 8'b00000000; // 3423 :   0 - 0x0
      13'hD60: dout <= 8'b10001111; // 3424 : 143 - 0x8f -- Sprite 0xd6
      13'hD61: dout <= 8'b11101111; // 3425 : 239 - 0xef
      13'hD62: dout <= 8'b11000000; // 3426 : 192 - 0xc0
      13'hD63: dout <= 8'b11110000; // 3427 : 240 - 0xf0
      13'hD64: dout <= 8'b11100000; // 3428 : 224 - 0xe0
      13'hD65: dout <= 8'b11111111; // 3429 : 255 - 0xff
      13'hD66: dout <= 8'b11111111; // 3430 : 255 - 0xff
      13'hD67: dout <= 8'b11111111; // 3431 : 255 - 0xff
      13'hD68: dout <= 8'b00001111; // 3432 :  15 - 0xf
      13'hD69: dout <= 8'b00001111; // 3433 :  15 - 0xf
      13'hD6A: dout <= 8'b00000000; // 3434 :   0 - 0x0
      13'hD6B: dout <= 8'b00000111; // 3435 :   7 - 0x7
      13'hD6C: dout <= 8'b00000000; // 3436 :   0 - 0x0
      13'hD6D: dout <= 8'b00000000; // 3437 :   0 - 0x0
      13'hD6E: dout <= 8'b00000000; // 3438 :   0 - 0x0
      13'hD6F: dout <= 8'b00000000; // 3439 :   0 - 0x0
      13'hD70: dout <= 8'b11111111; // 3440 : 255 - 0xff -- Sprite 0xd7
      13'hD71: dout <= 8'b11111111; // 3441 : 255 - 0xff
      13'hD72: dout <= 8'b00000000; // 3442 :   0 - 0x0
      13'hD73: dout <= 8'b00000000; // 3443 :   0 - 0x0
      13'hD74: dout <= 8'b00000000; // 3444 :   0 - 0x0
      13'hD75: dout <= 8'b11111111; // 3445 : 255 - 0xff
      13'hD76: dout <= 8'b11111111; // 3446 : 255 - 0xff
      13'hD77: dout <= 8'b11111111; // 3447 : 255 - 0xff
      13'hD78: dout <= 8'b11111111; // 3448 : 255 - 0xff
      13'hD79: dout <= 8'b11111111; // 3449 : 255 - 0xff
      13'hD7A: dout <= 8'b00000000; // 3450 :   0 - 0x0
      13'hD7B: dout <= 8'b11111111; // 3451 : 255 - 0xff
      13'hD7C: dout <= 8'b00000000; // 3452 :   0 - 0x0
      13'hD7D: dout <= 8'b00000000; // 3453 :   0 - 0x0
      13'hD7E: dout <= 8'b00000000; // 3454 :   0 - 0x0
      13'hD7F: dout <= 8'b00000000; // 3455 :   0 - 0x0
      13'hD80: dout <= 8'b11000011; // 3456 : 195 - 0xc3 -- Sprite 0xd8
      13'hD81: dout <= 8'b11111111; // 3457 : 255 - 0xff
      13'hD82: dout <= 8'b00000000; // 3458 :   0 - 0x0
      13'hD83: dout <= 8'b00000000; // 3459 :   0 - 0x0
      13'hD84: dout <= 8'b00000000; // 3460 :   0 - 0x0
      13'hD85: dout <= 8'b11111111; // 3461 : 255 - 0xff
      13'hD86: dout <= 8'b11111111; // 3462 : 255 - 0xff
      13'hD87: dout <= 8'b11111111; // 3463 : 255 - 0xff
      13'hD88: dout <= 8'b11000011; // 3464 : 195 - 0xc3
      13'hD89: dout <= 8'b11111111; // 3465 : 255 - 0xff
      13'hD8A: dout <= 8'b00000000; // 3466 :   0 - 0x0
      13'hD8B: dout <= 8'b11111111; // 3467 : 255 - 0xff
      13'hD8C: dout <= 8'b00000000; // 3468 :   0 - 0x0
      13'hD8D: dout <= 8'b00000000; // 3469 :   0 - 0x0
      13'hD8E: dout <= 8'b00000000; // 3470 :   0 - 0x0
      13'hD8F: dout <= 8'b00000000; // 3471 :   0 - 0x0
      13'hD90: dout <= 8'b00000011; // 3472 :   3 - 0x3 -- Sprite 0xd9
      13'hD91: dout <= 8'b10000001; // 3473 : 129 - 0x81
      13'hD92: dout <= 8'b00000000; // 3474 :   0 - 0x0
      13'hD93: dout <= 8'b00000000; // 3475 :   0 - 0x0
      13'hD94: dout <= 8'b00000011; // 3476 :   3 - 0x3
      13'hD95: dout <= 8'b11111111; // 3477 : 255 - 0xff
      13'hD96: dout <= 8'b11111111; // 3478 : 255 - 0xff
      13'hD97: dout <= 8'b11111111; // 3479 : 255 - 0xff
      13'hD98: dout <= 8'b01101011; // 3480 : 107 - 0x6b
      13'hD99: dout <= 8'b10110101; // 3481 : 181 - 0xb5
      13'hD9A: dout <= 8'b00110110; // 3482 :  54 - 0x36
      13'hD9B: dout <= 8'b11111000; // 3483 : 248 - 0xf8
      13'hD9C: dout <= 8'b00000000; // 3484 :   0 - 0x0
      13'hD9D: dout <= 8'b00000000; // 3485 :   0 - 0x0
      13'hD9E: dout <= 8'b00000000; // 3486 :   0 - 0x0
      13'hD9F: dout <= 8'b00000000; // 3487 :   0 - 0x0
      13'hDA0: dout <= 8'b11111111; // 3488 : 255 - 0xff -- Sprite 0xda
      13'hDA1: dout <= 8'b11111111; // 3489 : 255 - 0xff
      13'hDA2: dout <= 8'b01111110; // 3490 : 126 - 0x7e
      13'hDA3: dout <= 8'b00000000; // 3491 :   0 - 0x0
      13'hDA4: dout <= 8'b00000000; // 3492 :   0 - 0x0
      13'hDA5: dout <= 8'b11100000; // 3493 : 224 - 0xe0
      13'hDA6: dout <= 8'b11111111; // 3494 : 255 - 0xff
      13'hDA7: dout <= 8'b11111111; // 3495 : 255 - 0xff
      13'hDA8: dout <= 8'b11111111; // 3496 : 255 - 0xff
      13'hDA9: dout <= 8'b11111111; // 3497 : 255 - 0xff
      13'hDAA: dout <= 8'b01111110; // 3498 : 126 - 0x7e
      13'hDAB: dout <= 8'b10000001; // 3499 : 129 - 0x81
      13'hDAC: dout <= 8'b00011111; // 3500 :  31 - 0x1f
      13'hDAD: dout <= 8'b00000000; // 3501 :   0 - 0x0
      13'hDAE: dout <= 8'b00000000; // 3502 :   0 - 0x0
      13'hDAF: dout <= 8'b00000000; // 3503 :   0 - 0x0
      13'hDB0: dout <= 8'b01100001; // 3504 :  97 - 0x61 -- Sprite 0xdb
      13'hDB1: dout <= 8'b11000011; // 3505 : 195 - 0xc3
      13'hDB2: dout <= 8'b00000111; // 3506 :   7 - 0x7
      13'hDB3: dout <= 8'b00001111; // 3507 :  15 - 0xf
      13'hDB4: dout <= 8'b00011111; // 3508 :  31 - 0x1f
      13'hDB5: dout <= 8'b01111111; // 3509 : 127 - 0x7f
      13'hDB6: dout <= 8'b11111111; // 3510 : 255 - 0xff
      13'hDB7: dout <= 8'b11111111; // 3511 : 255 - 0xff
      13'hDB8: dout <= 8'b01101100; // 3512 : 108 - 0x6c
      13'hDB9: dout <= 8'b11011000; // 3513 : 216 - 0xd8
      13'hDBA: dout <= 8'b00110000; // 3514 :  48 - 0x30
      13'hDBB: dout <= 8'b11100000; // 3515 : 224 - 0xe0
      13'hDBC: dout <= 8'b10000000; // 3516 : 128 - 0x80
      13'hDBD: dout <= 8'b00000000; // 3517 :   0 - 0x0
      13'hDBE: dout <= 8'b00000000; // 3518 :   0 - 0x0
      13'hDBF: dout <= 8'b00000000; // 3519 :   0 - 0x0
      13'hDC0: dout <= 8'b00011111; // 3520 :  31 - 0x1f -- Sprite 0xdc
      13'hDC1: dout <= 8'b11011111; // 3521 : 223 - 0xdf
      13'hDC2: dout <= 8'b11000000; // 3522 : 192 - 0xc0
      13'hDC3: dout <= 8'b11110000; // 3523 : 240 - 0xf0
      13'hDC4: dout <= 8'b11110000; // 3524 : 240 - 0xf0
      13'hDC5: dout <= 8'b11111111; // 3525 : 255 - 0xff
      13'hDC6: dout <= 8'b11111111; // 3526 : 255 - 0xff
      13'hDC7: dout <= 8'b11111111; // 3527 : 255 - 0xff
      13'hDC8: dout <= 8'b00011111; // 3528 :  31 - 0x1f
      13'hDC9: dout <= 8'b00011111; // 3529 :  31 - 0x1f
      13'hDCA: dout <= 8'b00000000; // 3530 :   0 - 0x0
      13'hDCB: dout <= 8'b00000111; // 3531 :   7 - 0x7
      13'hDCC: dout <= 8'b00000000; // 3532 :   0 - 0x0
      13'hDCD: dout <= 8'b00000000; // 3533 :   0 - 0x0
      13'hDCE: dout <= 8'b00000000; // 3534 :   0 - 0x0
      13'hDCF: dout <= 8'b00000000; // 3535 :   0 - 0x0
      13'hDD0: dout <= 8'b10000100; // 3536 : 132 - 0x84 -- Sprite 0xdd
      13'hDD1: dout <= 8'b11111100; // 3537 : 252 - 0xfc
      13'hDD2: dout <= 8'b00000000; // 3538 :   0 - 0x0
      13'hDD3: dout <= 8'b00000000; // 3539 :   0 - 0x0
      13'hDD4: dout <= 8'b00000000; // 3540 :   0 - 0x0
      13'hDD5: dout <= 8'b11111111; // 3541 : 255 - 0xff
      13'hDD6: dout <= 8'b11111111; // 3542 : 255 - 0xff
      13'hDD7: dout <= 8'b11111111; // 3543 : 255 - 0xff
      13'hDD8: dout <= 8'b10000101; // 3544 : 133 - 0x85
      13'hDD9: dout <= 8'b11111101; // 3545 : 253 - 0xfd
      13'hDDA: dout <= 8'b00000001; // 3546 :   1 - 0x1
      13'hDDB: dout <= 8'b11111111; // 3547 : 255 - 0xff
      13'hDDC: dout <= 8'b00000000; // 3548 :   0 - 0x0
      13'hDDD: dout <= 8'b00000000; // 3549 :   0 - 0x0
      13'hDDE: dout <= 8'b00000000; // 3550 :   0 - 0x0
      13'hDDF: dout <= 8'b00000000; // 3551 :   0 - 0x0
      13'hDE0: dout <= 8'b01111111; // 3552 : 127 - 0x7f -- Sprite 0xde
      13'hDE1: dout <= 8'b01111111; // 3553 : 127 - 0x7f
      13'hDE2: dout <= 8'b00000000; // 3554 :   0 - 0x0
      13'hDE3: dout <= 8'b00000000; // 3555 :   0 - 0x0
      13'hDE4: dout <= 8'b00000000; // 3556 :   0 - 0x0
      13'hDE5: dout <= 8'b11111111; // 3557 : 255 - 0xff
      13'hDE6: dout <= 8'b11111111; // 3558 : 255 - 0xff
      13'hDE7: dout <= 8'b11111111; // 3559 : 255 - 0xff
      13'hDE8: dout <= 8'b01111111; // 3560 : 127 - 0x7f
      13'hDE9: dout <= 8'b01111111; // 3561 : 127 - 0x7f
      13'hDEA: dout <= 8'b00000000; // 3562 :   0 - 0x0
      13'hDEB: dout <= 8'b01011111; // 3563 :  95 - 0x5f
      13'hDEC: dout <= 8'b00000000; // 3564 :   0 - 0x0
      13'hDED: dout <= 8'b00000000; // 3565 :   0 - 0x0
      13'hDEE: dout <= 8'b00000000; // 3566 :   0 - 0x0
      13'hDEF: dout <= 8'b00000000; // 3567 :   0 - 0x0
      13'hDF0: dout <= 8'b11111100; // 3568 : 252 - 0xfc -- Sprite 0xdf
      13'hDF1: dout <= 8'b11111111; // 3569 : 255 - 0xff
      13'hDF2: dout <= 8'b00000000; // 3570 :   0 - 0x0
      13'hDF3: dout <= 8'b00000000; // 3571 :   0 - 0x0
      13'hDF4: dout <= 8'b00000000; // 3572 :   0 - 0x0
      13'hDF5: dout <= 8'b11111111; // 3573 : 255 - 0xff
      13'hDF6: dout <= 8'b11111111; // 3574 : 255 - 0xff
      13'hDF7: dout <= 8'b11111111; // 3575 : 255 - 0xff
      13'hDF8: dout <= 8'b11111100; // 3576 : 252 - 0xfc
      13'hDF9: dout <= 8'b11111111; // 3577 : 255 - 0xff
      13'hDFA: dout <= 8'b00000000; // 3578 :   0 - 0x0
      13'hDFB: dout <= 8'b11111111; // 3579 : 255 - 0xff
      13'hDFC: dout <= 8'b00000000; // 3580 :   0 - 0x0
      13'hDFD: dout <= 8'b00000000; // 3581 :   0 - 0x0
      13'hDFE: dout <= 8'b00000000; // 3582 :   0 - 0x0
      13'hDFF: dout <= 8'b00000000; // 3583 :   0 - 0x0
      13'hE00: dout <= 8'b00110000; // 3584 :  48 - 0x30 -- Sprite 0xe0
      13'hE01: dout <= 8'b11110000; // 3585 : 240 - 0xf0
      13'hE02: dout <= 8'b00000000; // 3586 :   0 - 0x0
      13'hE03: dout <= 8'b00000000; // 3587 :   0 - 0x0
      13'hE04: dout <= 8'b00000000; // 3588 :   0 - 0x0
      13'hE05: dout <= 8'b11111111; // 3589 : 255 - 0xff
      13'hE06: dout <= 8'b11111111; // 3590 : 255 - 0xff
      13'hE07: dout <= 8'b11111111; // 3591 : 255 - 0xff
      13'hE08: dout <= 8'b00110100; // 3592 :  52 - 0x34
      13'hE09: dout <= 8'b11110110; // 3593 : 246 - 0xf6
      13'hE0A: dout <= 8'b00000010; // 3594 :   2 - 0x2
      13'hE0B: dout <= 8'b11111111; // 3595 : 255 - 0xff
      13'hE0C: dout <= 8'b00000000; // 3596 :   0 - 0x0
      13'hE0D: dout <= 8'b00000000; // 3597 :   0 - 0x0
      13'hE0E: dout <= 8'b00000000; // 3598 :   0 - 0x0
      13'hE0F: dout <= 8'b00000000; // 3599 :   0 - 0x0
      13'hE10: dout <= 8'b11111111; // 3600 : 255 - 0xff -- Sprite 0xe1
      13'hE11: dout <= 8'b11111111; // 3601 : 255 - 0xff
      13'hE12: dout <= 8'b00000000; // 3602 :   0 - 0x0
      13'hE13: dout <= 8'b00000000; // 3603 :   0 - 0x0
      13'hE14: dout <= 8'b00000000; // 3604 :   0 - 0x0
      13'hE15: dout <= 8'b11111111; // 3605 : 255 - 0xff
      13'hE16: dout <= 8'b11111111; // 3606 : 255 - 0xff
      13'hE17: dout <= 8'b11111111; // 3607 : 255 - 0xff
      13'hE18: dout <= 8'b11111111; // 3608 : 255 - 0xff
      13'hE19: dout <= 8'b11111111; // 3609 : 255 - 0xff
      13'hE1A: dout <= 8'b00000000; // 3610 :   0 - 0x0
      13'hE1B: dout <= 8'b01111111; // 3611 : 127 - 0x7f
      13'hE1C: dout <= 8'b00000000; // 3612 :   0 - 0x0
      13'hE1D: dout <= 8'b00000000; // 3613 :   0 - 0x0
      13'hE1E: dout <= 8'b00000000; // 3614 :   0 - 0x0
      13'hE1F: dout <= 8'b00000000; // 3615 :   0 - 0x0
      13'hE20: dout <= 8'b11100001; // 3616 : 225 - 0xe1 -- Sprite 0xe2
      13'hE21: dout <= 8'b11111111; // 3617 : 255 - 0xff
      13'hE22: dout <= 8'b00000000; // 3618 :   0 - 0x0
      13'hE23: dout <= 8'b00000000; // 3619 :   0 - 0x0
      13'hE24: dout <= 8'b00000000; // 3620 :   0 - 0x0
      13'hE25: dout <= 8'b11111111; // 3621 : 255 - 0xff
      13'hE26: dout <= 8'b11111111; // 3622 : 255 - 0xff
      13'hE27: dout <= 8'b11111111; // 3623 : 255 - 0xff
      13'hE28: dout <= 8'b11100001; // 3624 : 225 - 0xe1
      13'hE29: dout <= 8'b11111111; // 3625 : 255 - 0xff
      13'hE2A: dout <= 8'b00000000; // 3626 :   0 - 0x0
      13'hE2B: dout <= 8'b11111111; // 3627 : 255 - 0xff
      13'hE2C: dout <= 8'b00000000; // 3628 :   0 - 0x0
      13'hE2D: dout <= 8'b00000000; // 3629 :   0 - 0x0
      13'hE2E: dout <= 8'b00000000; // 3630 :   0 - 0x0
      13'hE2F: dout <= 8'b00000000; // 3631 :   0 - 0x0
      13'hE30: dout <= 8'b00011111; // 3632 :  31 - 0x1f -- Sprite 0xe3
      13'hE31: dout <= 8'b00011111; // 3633 :  31 - 0x1f
      13'hE32: dout <= 8'b00011111; // 3634 :  31 - 0x1f
      13'hE33: dout <= 8'b00011111; // 3635 :  31 - 0x1f
      13'hE34: dout <= 8'b00011111; // 3636 :  31 - 0x1f
      13'hE35: dout <= 8'b11111111; // 3637 : 255 - 0xff
      13'hE36: dout <= 8'b11111111; // 3638 : 255 - 0xff
      13'hE37: dout <= 8'b11111111; // 3639 : 255 - 0xff
      13'hE38: dout <= 8'b01000000; // 3640 :  64 - 0x40
      13'hE39: dout <= 8'b01000000; // 3641 :  64 - 0x40
      13'hE3A: dout <= 8'b01000000; // 3642 :  64 - 0x40
      13'hE3B: dout <= 8'b11000000; // 3643 : 192 - 0xc0
      13'hE3C: dout <= 8'b00000000; // 3644 :   0 - 0x0
      13'hE3D: dout <= 8'b00000000; // 3645 :   0 - 0x0
      13'hE3E: dout <= 8'b00000000; // 3646 :   0 - 0x0
      13'hE3F: dout <= 8'b00000000; // 3647 :   0 - 0x0
      13'hE40: dout <= 8'b00000000; // 3648 :   0 - 0x0 -- Sprite 0xe4
      13'hE41: dout <= 8'b00011111; // 3649 :  31 - 0x1f
      13'hE42: dout <= 8'b00111111; // 3650 :  63 - 0x3f
      13'hE43: dout <= 8'b01111000; // 3651 : 120 - 0x78
      13'hE44: dout <= 8'b01110111; // 3652 : 119 - 0x77
      13'hE45: dout <= 8'b01101111; // 3653 : 111 - 0x6f
      13'hE46: dout <= 8'b01101111; // 3654 : 111 - 0x6f
      13'hE47: dout <= 8'b01101111; // 3655 : 111 - 0x6f
      13'hE48: dout <= 8'b00000000; // 3656 :   0 - 0x0
      13'hE49: dout <= 8'b00000000; // 3657 :   0 - 0x0
      13'hE4A: dout <= 8'b00000000; // 3658 :   0 - 0x0
      13'hE4B: dout <= 8'b00000000; // 3659 :   0 - 0x0
      13'hE4C: dout <= 8'b00000111; // 3660 :   7 - 0x7
      13'hE4D: dout <= 8'b00001111; // 3661 :  15 - 0xf
      13'hE4E: dout <= 8'b00001111; // 3662 :  15 - 0xf
      13'hE4F: dout <= 8'b00001111; // 3663 :  15 - 0xf
      13'hE50: dout <= 8'b00000000; // 3664 :   0 - 0x0 -- Sprite 0xe5
      13'hE51: dout <= 8'b11111000; // 3665 : 248 - 0xf8
      13'hE52: dout <= 8'b11111100; // 3666 : 252 - 0xfc
      13'hE53: dout <= 8'b00011110; // 3667 :  30 - 0x1e
      13'hE54: dout <= 8'b11101110; // 3668 : 238 - 0xee
      13'hE55: dout <= 8'b11110110; // 3669 : 246 - 0xf6
      13'hE56: dout <= 8'b11110110; // 3670 : 246 - 0xf6
      13'hE57: dout <= 8'b11110110; // 3671 : 246 - 0xf6
      13'hE58: dout <= 8'b00000000; // 3672 :   0 - 0x0
      13'hE59: dout <= 8'b00000000; // 3673 :   0 - 0x0
      13'hE5A: dout <= 8'b00000000; // 3674 :   0 - 0x0
      13'hE5B: dout <= 8'b00000000; // 3675 :   0 - 0x0
      13'hE5C: dout <= 8'b11100000; // 3676 : 224 - 0xe0
      13'hE5D: dout <= 8'b11110000; // 3677 : 240 - 0xf0
      13'hE5E: dout <= 8'b11110000; // 3678 : 240 - 0xf0
      13'hE5F: dout <= 8'b11110000; // 3679 : 240 - 0xf0
      13'hE60: dout <= 8'b11110110; // 3680 : 246 - 0xf6 -- Sprite 0xe6
      13'hE61: dout <= 8'b11110110; // 3681 : 246 - 0xf6
      13'hE62: dout <= 8'b11110110; // 3682 : 246 - 0xf6
      13'hE63: dout <= 8'b11101110; // 3683 : 238 - 0xee
      13'hE64: dout <= 8'b00011110; // 3684 :  30 - 0x1e
      13'hE65: dout <= 8'b11111100; // 3685 : 252 - 0xfc
      13'hE66: dout <= 8'b11111000; // 3686 : 248 - 0xf8
      13'hE67: dout <= 8'b00000000; // 3687 :   0 - 0x0
      13'hE68: dout <= 8'b11110000; // 3688 : 240 - 0xf0
      13'hE69: dout <= 8'b11110000; // 3689 : 240 - 0xf0
      13'hE6A: dout <= 8'b11110000; // 3690 : 240 - 0xf0
      13'hE6B: dout <= 8'b11100000; // 3691 : 224 - 0xe0
      13'hE6C: dout <= 8'b00000000; // 3692 :   0 - 0x0
      13'hE6D: dout <= 8'b00000000; // 3693 :   0 - 0x0
      13'hE6E: dout <= 8'b00000000; // 3694 :   0 - 0x0
      13'hE6F: dout <= 8'b00000000; // 3695 :   0 - 0x0
      13'hE70: dout <= 8'b01101111; // 3696 : 111 - 0x6f -- Sprite 0xe7
      13'hE71: dout <= 8'b01101111; // 3697 : 111 - 0x6f
      13'hE72: dout <= 8'b01101111; // 3698 : 111 - 0x6f
      13'hE73: dout <= 8'b01110111; // 3699 : 119 - 0x77
      13'hE74: dout <= 8'b01111000; // 3700 : 120 - 0x78
      13'hE75: dout <= 8'b00111111; // 3701 :  63 - 0x3f
      13'hE76: dout <= 8'b00011111; // 3702 :  31 - 0x1f
      13'hE77: dout <= 8'b00000000; // 3703 :   0 - 0x0
      13'hE78: dout <= 8'b00001111; // 3704 :  15 - 0xf
      13'hE79: dout <= 8'b00001111; // 3705 :  15 - 0xf
      13'hE7A: dout <= 8'b00001111; // 3706 :  15 - 0xf
      13'hE7B: dout <= 8'b00000111; // 3707 :   7 - 0x7
      13'hE7C: dout <= 8'b00000000; // 3708 :   0 - 0x0
      13'hE7D: dout <= 8'b00000000; // 3709 :   0 - 0x0
      13'hE7E: dout <= 8'b00000000; // 3710 :   0 - 0x0
      13'hE7F: dout <= 8'b00000000; // 3711 :   0 - 0x0
      13'hE80: dout <= 8'b00000000; // 3712 :   0 - 0x0 -- Sprite 0xe8
      13'hE81: dout <= 8'b11111111; // 3713 : 255 - 0xff
      13'hE82: dout <= 8'b11111111; // 3714 : 255 - 0xff
      13'hE83: dout <= 8'b00000000; // 3715 :   0 - 0x0
      13'hE84: dout <= 8'b11111111; // 3716 : 255 - 0xff
      13'hE85: dout <= 8'b11111111; // 3717 : 255 - 0xff
      13'hE86: dout <= 8'b11111111; // 3718 : 255 - 0xff
      13'hE87: dout <= 8'b11111111; // 3719 : 255 - 0xff
      13'hE88: dout <= 8'b00000000; // 3720 :   0 - 0x0
      13'hE89: dout <= 8'b00000000; // 3721 :   0 - 0x0
      13'hE8A: dout <= 8'b00000000; // 3722 :   0 - 0x0
      13'hE8B: dout <= 8'b00000000; // 3723 :   0 - 0x0
      13'hE8C: dout <= 8'b11111111; // 3724 : 255 - 0xff
      13'hE8D: dout <= 8'b11111111; // 3725 : 255 - 0xff
      13'hE8E: dout <= 8'b11111111; // 3726 : 255 - 0xff
      13'hE8F: dout <= 8'b11111111; // 3727 : 255 - 0xff
      13'hE90: dout <= 8'b11110110; // 3728 : 246 - 0xf6 -- Sprite 0xe9
      13'hE91: dout <= 8'b11110110; // 3729 : 246 - 0xf6
      13'hE92: dout <= 8'b11110110; // 3730 : 246 - 0xf6
      13'hE93: dout <= 8'b11110110; // 3731 : 246 - 0xf6
      13'hE94: dout <= 8'b11110110; // 3732 : 246 - 0xf6
      13'hE95: dout <= 8'b11110110; // 3733 : 246 - 0xf6
      13'hE96: dout <= 8'b11110110; // 3734 : 246 - 0xf6
      13'hE97: dout <= 8'b11110110; // 3735 : 246 - 0xf6
      13'hE98: dout <= 8'b11110000; // 3736 : 240 - 0xf0
      13'hE99: dout <= 8'b11110000; // 3737 : 240 - 0xf0
      13'hE9A: dout <= 8'b11110000; // 3738 : 240 - 0xf0
      13'hE9B: dout <= 8'b11110000; // 3739 : 240 - 0xf0
      13'hE9C: dout <= 8'b11110000; // 3740 : 240 - 0xf0
      13'hE9D: dout <= 8'b11110000; // 3741 : 240 - 0xf0
      13'hE9E: dout <= 8'b11110000; // 3742 : 240 - 0xf0
      13'hE9F: dout <= 8'b11110000; // 3743 : 240 - 0xf0
      13'hEA0: dout <= 8'b11111111; // 3744 : 255 - 0xff -- Sprite 0xea
      13'hEA1: dout <= 8'b11111111; // 3745 : 255 - 0xff
      13'hEA2: dout <= 8'b11111111; // 3746 : 255 - 0xff
      13'hEA3: dout <= 8'b11111111; // 3747 : 255 - 0xff
      13'hEA4: dout <= 8'b00000000; // 3748 :   0 - 0x0
      13'hEA5: dout <= 8'b11111111; // 3749 : 255 - 0xff
      13'hEA6: dout <= 8'b11111111; // 3750 : 255 - 0xff
      13'hEA7: dout <= 8'b00000000; // 3751 :   0 - 0x0
      13'hEA8: dout <= 8'b11111111; // 3752 : 255 - 0xff
      13'hEA9: dout <= 8'b11111111; // 3753 : 255 - 0xff
      13'hEAA: dout <= 8'b11111111; // 3754 : 255 - 0xff
      13'hEAB: dout <= 8'b11111111; // 3755 : 255 - 0xff
      13'hEAC: dout <= 8'b00000000; // 3756 :   0 - 0x0
      13'hEAD: dout <= 8'b00000000; // 3757 :   0 - 0x0
      13'hEAE: dout <= 8'b00000000; // 3758 :   0 - 0x0
      13'hEAF: dout <= 8'b00000000; // 3759 :   0 - 0x0
      13'hEB0: dout <= 8'b01101111; // 3760 : 111 - 0x6f -- Sprite 0xeb
      13'hEB1: dout <= 8'b01101111; // 3761 : 111 - 0x6f
      13'hEB2: dout <= 8'b01101111; // 3762 : 111 - 0x6f
      13'hEB3: dout <= 8'b01101111; // 3763 : 111 - 0x6f
      13'hEB4: dout <= 8'b01101111; // 3764 : 111 - 0x6f
      13'hEB5: dout <= 8'b01101111; // 3765 : 111 - 0x6f
      13'hEB6: dout <= 8'b01101111; // 3766 : 111 - 0x6f
      13'hEB7: dout <= 8'b01101111; // 3767 : 111 - 0x6f
      13'hEB8: dout <= 8'b00001111; // 3768 :  15 - 0xf
      13'hEB9: dout <= 8'b00001111; // 3769 :  15 - 0xf
      13'hEBA: dout <= 8'b00001111; // 3770 :  15 - 0xf
      13'hEBB: dout <= 8'b00001111; // 3771 :  15 - 0xf
      13'hEBC: dout <= 8'b00001111; // 3772 :  15 - 0xf
      13'hEBD: dout <= 8'b00001111; // 3773 :  15 - 0xf
      13'hEBE: dout <= 8'b00001111; // 3774 :  15 - 0xf
      13'hEBF: dout <= 8'b00001111; // 3775 :  15 - 0xf
      13'hEC0: dout <= 8'b00000000; // 3776 :   0 - 0x0 -- Sprite 0xec
      13'hEC1: dout <= 8'b00000000; // 3777 :   0 - 0x0
      13'hEC2: dout <= 8'b00000000; // 3778 :   0 - 0x0
      13'hEC3: dout <= 8'b00000000; // 3779 :   0 - 0x0
      13'hEC4: dout <= 8'b00000000; // 3780 :   0 - 0x0
      13'hEC5: dout <= 8'b00000000; // 3781 :   0 - 0x0
      13'hEC6: dout <= 8'b00000000; // 3782 :   0 - 0x0
      13'hEC7: dout <= 8'b00000000; // 3783 :   0 - 0x0
      13'hEC8: dout <= 8'b00000000; // 3784 :   0 - 0x0
      13'hEC9: dout <= 8'b00000000; // 3785 :   0 - 0x0
      13'hECA: dout <= 8'b00000000; // 3786 :   0 - 0x0
      13'hECB: dout <= 8'b00000000; // 3787 :   0 - 0x0
      13'hECC: dout <= 8'b00000000; // 3788 :   0 - 0x0
      13'hECD: dout <= 8'b00000000; // 3789 :   0 - 0x0
      13'hECE: dout <= 8'b00000000; // 3790 :   0 - 0x0
      13'hECF: dout <= 8'b00000000; // 3791 :   0 - 0x0
      13'hED0: dout <= 8'b00000000; // 3792 :   0 - 0x0 -- Sprite 0xed
      13'hED1: dout <= 8'b00000000; // 3793 :   0 - 0x0
      13'hED2: dout <= 8'b00000000; // 3794 :   0 - 0x0
      13'hED3: dout <= 8'b00000000; // 3795 :   0 - 0x0
      13'hED4: dout <= 8'b00000000; // 3796 :   0 - 0x0
      13'hED5: dout <= 8'b00000000; // 3797 :   0 - 0x0
      13'hED6: dout <= 8'b00000000; // 3798 :   0 - 0x0
      13'hED7: dout <= 8'b00000000; // 3799 :   0 - 0x0
      13'hED8: dout <= 8'b00000000; // 3800 :   0 - 0x0
      13'hED9: dout <= 8'b00000000; // 3801 :   0 - 0x0
      13'hEDA: dout <= 8'b00000000; // 3802 :   0 - 0x0
      13'hEDB: dout <= 8'b00000000; // 3803 :   0 - 0x0
      13'hEDC: dout <= 8'b00000000; // 3804 :   0 - 0x0
      13'hEDD: dout <= 8'b00000000; // 3805 :   0 - 0x0
      13'hEDE: dout <= 8'b00000000; // 3806 :   0 - 0x0
      13'hEDF: dout <= 8'b00000000; // 3807 :   0 - 0x0
      13'hEE0: dout <= 8'b00000000; // 3808 :   0 - 0x0 -- Sprite 0xee
      13'hEE1: dout <= 8'b00000000; // 3809 :   0 - 0x0
      13'hEE2: dout <= 8'b00000000; // 3810 :   0 - 0x0
      13'hEE3: dout <= 8'b00000000; // 3811 :   0 - 0x0
      13'hEE4: dout <= 8'b00000000; // 3812 :   0 - 0x0
      13'hEE5: dout <= 8'b00000000; // 3813 :   0 - 0x0
      13'hEE6: dout <= 8'b00000000; // 3814 :   0 - 0x0
      13'hEE7: dout <= 8'b00000000; // 3815 :   0 - 0x0
      13'hEE8: dout <= 8'b00000000; // 3816 :   0 - 0x0
      13'hEE9: dout <= 8'b00000000; // 3817 :   0 - 0x0
      13'hEEA: dout <= 8'b00000000; // 3818 :   0 - 0x0
      13'hEEB: dout <= 8'b00000000; // 3819 :   0 - 0x0
      13'hEEC: dout <= 8'b00000000; // 3820 :   0 - 0x0
      13'hEED: dout <= 8'b00000000; // 3821 :   0 - 0x0
      13'hEEE: dout <= 8'b00000000; // 3822 :   0 - 0x0
      13'hEEF: dout <= 8'b00000000; // 3823 :   0 - 0x0
      13'hEF0: dout <= 8'b00000000; // 3824 :   0 - 0x0 -- Sprite 0xef
      13'hEF1: dout <= 8'b00000000; // 3825 :   0 - 0x0
      13'hEF2: dout <= 8'b00000000; // 3826 :   0 - 0x0
      13'hEF3: dout <= 8'b00000000; // 3827 :   0 - 0x0
      13'hEF4: dout <= 8'b00000000; // 3828 :   0 - 0x0
      13'hEF5: dout <= 8'b00000000; // 3829 :   0 - 0x0
      13'hEF6: dout <= 8'b00000000; // 3830 :   0 - 0x0
      13'hEF7: dout <= 8'b00000000; // 3831 :   0 - 0x0
      13'hEF8: dout <= 8'b00000000; // 3832 :   0 - 0x0
      13'hEF9: dout <= 8'b00000000; // 3833 :   0 - 0x0
      13'hEFA: dout <= 8'b00000000; // 3834 :   0 - 0x0
      13'hEFB: dout <= 8'b00000000; // 3835 :   0 - 0x0
      13'hEFC: dout <= 8'b00000000; // 3836 :   0 - 0x0
      13'hEFD: dout <= 8'b00000000; // 3837 :   0 - 0x0
      13'hEFE: dout <= 8'b00000000; // 3838 :   0 - 0x0
      13'hEFF: dout <= 8'b00000000; // 3839 :   0 - 0x0
      13'hF00: dout <= 8'b11111111; // 3840 : 255 - 0xff -- Sprite 0xf0
      13'hF01: dout <= 8'b11111111; // 3841 : 255 - 0xff
      13'hF02: dout <= 8'b11111111; // 3842 : 255 - 0xff
      13'hF03: dout <= 8'b11111111; // 3843 : 255 - 0xff
      13'hF04: dout <= 8'b11111111; // 3844 : 255 - 0xff
      13'hF05: dout <= 8'b11111111; // 3845 : 255 - 0xff
      13'hF06: dout <= 8'b11111111; // 3846 : 255 - 0xff
      13'hF07: dout <= 8'b11111111; // 3847 : 255 - 0xff
      13'hF08: dout <= 8'b11111111; // 3848 : 255 - 0xff
      13'hF09: dout <= 8'b11111111; // 3849 : 255 - 0xff
      13'hF0A: dout <= 8'b11111111; // 3850 : 255 - 0xff
      13'hF0B: dout <= 8'b11111111; // 3851 : 255 - 0xff
      13'hF0C: dout <= 8'b11111111; // 3852 : 255 - 0xff
      13'hF0D: dout <= 8'b11111111; // 3853 : 255 - 0xff
      13'hF0E: dout <= 8'b11111111; // 3854 : 255 - 0xff
      13'hF0F: dout <= 8'b11111111; // 3855 : 255 - 0xff
      13'hF10: dout <= 8'b11111111; // 3856 : 255 - 0xff -- Sprite 0xf1
      13'hF11: dout <= 8'b11111111; // 3857 : 255 - 0xff
      13'hF12: dout <= 8'b11111111; // 3858 : 255 - 0xff
      13'hF13: dout <= 8'b11111111; // 3859 : 255 - 0xff
      13'hF14: dout <= 8'b11111111; // 3860 : 255 - 0xff
      13'hF15: dout <= 8'b11111111; // 3861 : 255 - 0xff
      13'hF16: dout <= 8'b11111111; // 3862 : 255 - 0xff
      13'hF17: dout <= 8'b11111111; // 3863 : 255 - 0xff
      13'hF18: dout <= 8'b11111111; // 3864 : 255 - 0xff
      13'hF19: dout <= 8'b11111111; // 3865 : 255 - 0xff
      13'hF1A: dout <= 8'b11111111; // 3866 : 255 - 0xff
      13'hF1B: dout <= 8'b11111111; // 3867 : 255 - 0xff
      13'hF1C: dout <= 8'b11111111; // 3868 : 255 - 0xff
      13'hF1D: dout <= 8'b11111111; // 3869 : 255 - 0xff
      13'hF1E: dout <= 8'b11111111; // 3870 : 255 - 0xff
      13'hF1F: dout <= 8'b11111111; // 3871 : 255 - 0xff
      13'hF20: dout <= 8'b11111111; // 3872 : 255 - 0xff -- Sprite 0xf2
      13'hF21: dout <= 8'b11111111; // 3873 : 255 - 0xff
      13'hF22: dout <= 8'b11111111; // 3874 : 255 - 0xff
      13'hF23: dout <= 8'b11111111; // 3875 : 255 - 0xff
      13'hF24: dout <= 8'b11111111; // 3876 : 255 - 0xff
      13'hF25: dout <= 8'b11111111; // 3877 : 255 - 0xff
      13'hF26: dout <= 8'b11111111; // 3878 : 255 - 0xff
      13'hF27: dout <= 8'b11111111; // 3879 : 255 - 0xff
      13'hF28: dout <= 8'b11111111; // 3880 : 255 - 0xff
      13'hF29: dout <= 8'b11111111; // 3881 : 255 - 0xff
      13'hF2A: dout <= 8'b11111111; // 3882 : 255 - 0xff
      13'hF2B: dout <= 8'b11111111; // 3883 : 255 - 0xff
      13'hF2C: dout <= 8'b11111111; // 3884 : 255 - 0xff
      13'hF2D: dout <= 8'b11111111; // 3885 : 255 - 0xff
      13'hF2E: dout <= 8'b11111111; // 3886 : 255 - 0xff
      13'hF2F: dout <= 8'b11111111; // 3887 : 255 - 0xff
      13'hF30: dout <= 8'b11111111; // 3888 : 255 - 0xff -- Sprite 0xf3
      13'hF31: dout <= 8'b11111111; // 3889 : 255 - 0xff
      13'hF32: dout <= 8'b11111111; // 3890 : 255 - 0xff
      13'hF33: dout <= 8'b11111111; // 3891 : 255 - 0xff
      13'hF34: dout <= 8'b11111111; // 3892 : 255 - 0xff
      13'hF35: dout <= 8'b11111111; // 3893 : 255 - 0xff
      13'hF36: dout <= 8'b11111111; // 3894 : 255 - 0xff
      13'hF37: dout <= 8'b11111111; // 3895 : 255 - 0xff
      13'hF38: dout <= 8'b11111111; // 3896 : 255 - 0xff
      13'hF39: dout <= 8'b11111111; // 3897 : 255 - 0xff
      13'hF3A: dout <= 8'b11111111; // 3898 : 255 - 0xff
      13'hF3B: dout <= 8'b11111111; // 3899 : 255 - 0xff
      13'hF3C: dout <= 8'b11111111; // 3900 : 255 - 0xff
      13'hF3D: dout <= 8'b11111111; // 3901 : 255 - 0xff
      13'hF3E: dout <= 8'b11111111; // 3902 : 255 - 0xff
      13'hF3F: dout <= 8'b11111111; // 3903 : 255 - 0xff
      13'hF40: dout <= 8'b11111111; // 3904 : 255 - 0xff -- Sprite 0xf4
      13'hF41: dout <= 8'b11111111; // 3905 : 255 - 0xff
      13'hF42: dout <= 8'b11111111; // 3906 : 255 - 0xff
      13'hF43: dout <= 8'b11111111; // 3907 : 255 - 0xff
      13'hF44: dout <= 8'b11111111; // 3908 : 255 - 0xff
      13'hF45: dout <= 8'b11111111; // 3909 : 255 - 0xff
      13'hF46: dout <= 8'b11111111; // 3910 : 255 - 0xff
      13'hF47: dout <= 8'b11111111; // 3911 : 255 - 0xff
      13'hF48: dout <= 8'b11111111; // 3912 : 255 - 0xff
      13'hF49: dout <= 8'b11111111; // 3913 : 255 - 0xff
      13'hF4A: dout <= 8'b11111111; // 3914 : 255 - 0xff
      13'hF4B: dout <= 8'b11111111; // 3915 : 255 - 0xff
      13'hF4C: dout <= 8'b11111111; // 3916 : 255 - 0xff
      13'hF4D: dout <= 8'b11111111; // 3917 : 255 - 0xff
      13'hF4E: dout <= 8'b11111111; // 3918 : 255 - 0xff
      13'hF4F: dout <= 8'b11111111; // 3919 : 255 - 0xff
      13'hF50: dout <= 8'b11111111; // 3920 : 255 - 0xff -- Sprite 0xf5
      13'hF51: dout <= 8'b11111111; // 3921 : 255 - 0xff
      13'hF52: dout <= 8'b11111111; // 3922 : 255 - 0xff
      13'hF53: dout <= 8'b11111111; // 3923 : 255 - 0xff
      13'hF54: dout <= 8'b11111111; // 3924 : 255 - 0xff
      13'hF55: dout <= 8'b11111111; // 3925 : 255 - 0xff
      13'hF56: dout <= 8'b11111111; // 3926 : 255 - 0xff
      13'hF57: dout <= 8'b11111111; // 3927 : 255 - 0xff
      13'hF58: dout <= 8'b11111111; // 3928 : 255 - 0xff
      13'hF59: dout <= 8'b11111111; // 3929 : 255 - 0xff
      13'hF5A: dout <= 8'b11111111; // 3930 : 255 - 0xff
      13'hF5B: dout <= 8'b11111111; // 3931 : 255 - 0xff
      13'hF5C: dout <= 8'b11111111; // 3932 : 255 - 0xff
      13'hF5D: dout <= 8'b11111111; // 3933 : 255 - 0xff
      13'hF5E: dout <= 8'b11111111; // 3934 : 255 - 0xff
      13'hF5F: dout <= 8'b11111111; // 3935 : 255 - 0xff
      13'hF60: dout <= 8'b11111111; // 3936 : 255 - 0xff -- Sprite 0xf6
      13'hF61: dout <= 8'b11111111; // 3937 : 255 - 0xff
      13'hF62: dout <= 8'b11111111; // 3938 : 255 - 0xff
      13'hF63: dout <= 8'b11111111; // 3939 : 255 - 0xff
      13'hF64: dout <= 8'b11111111; // 3940 : 255 - 0xff
      13'hF65: dout <= 8'b11111111; // 3941 : 255 - 0xff
      13'hF66: dout <= 8'b11111111; // 3942 : 255 - 0xff
      13'hF67: dout <= 8'b11111111; // 3943 : 255 - 0xff
      13'hF68: dout <= 8'b11111111; // 3944 : 255 - 0xff
      13'hF69: dout <= 8'b11111111; // 3945 : 255 - 0xff
      13'hF6A: dout <= 8'b11111111; // 3946 : 255 - 0xff
      13'hF6B: dout <= 8'b11111111; // 3947 : 255 - 0xff
      13'hF6C: dout <= 8'b11111111; // 3948 : 255 - 0xff
      13'hF6D: dout <= 8'b11111111; // 3949 : 255 - 0xff
      13'hF6E: dout <= 8'b11111111; // 3950 : 255 - 0xff
      13'hF6F: dout <= 8'b11111111; // 3951 : 255 - 0xff
      13'hF70: dout <= 8'b11111111; // 3952 : 255 - 0xff -- Sprite 0xf7
      13'hF71: dout <= 8'b11111111; // 3953 : 255 - 0xff
      13'hF72: dout <= 8'b11111111; // 3954 : 255 - 0xff
      13'hF73: dout <= 8'b11111111; // 3955 : 255 - 0xff
      13'hF74: dout <= 8'b11111111; // 3956 : 255 - 0xff
      13'hF75: dout <= 8'b11111111; // 3957 : 255 - 0xff
      13'hF76: dout <= 8'b11111111; // 3958 : 255 - 0xff
      13'hF77: dout <= 8'b11111111; // 3959 : 255 - 0xff
      13'hF78: dout <= 8'b11111111; // 3960 : 255 - 0xff
      13'hF79: dout <= 8'b11111111; // 3961 : 255 - 0xff
      13'hF7A: dout <= 8'b11111111; // 3962 : 255 - 0xff
      13'hF7B: dout <= 8'b11111111; // 3963 : 255 - 0xff
      13'hF7C: dout <= 8'b11111111; // 3964 : 255 - 0xff
      13'hF7D: dout <= 8'b11111111; // 3965 : 255 - 0xff
      13'hF7E: dout <= 8'b11111111; // 3966 : 255 - 0xff
      13'hF7F: dout <= 8'b11111111; // 3967 : 255 - 0xff
      13'hF80: dout <= 8'b11111111; // 3968 : 255 - 0xff -- Sprite 0xf8
      13'hF81: dout <= 8'b11111111; // 3969 : 255 - 0xff
      13'hF82: dout <= 8'b11111111; // 3970 : 255 - 0xff
      13'hF83: dout <= 8'b11111111; // 3971 : 255 - 0xff
      13'hF84: dout <= 8'b11111111; // 3972 : 255 - 0xff
      13'hF85: dout <= 8'b11111111; // 3973 : 255 - 0xff
      13'hF86: dout <= 8'b11111111; // 3974 : 255 - 0xff
      13'hF87: dout <= 8'b11111111; // 3975 : 255 - 0xff
      13'hF88: dout <= 8'b11111111; // 3976 : 255 - 0xff
      13'hF89: dout <= 8'b11111111; // 3977 : 255 - 0xff
      13'hF8A: dout <= 8'b11111111; // 3978 : 255 - 0xff
      13'hF8B: dout <= 8'b11111111; // 3979 : 255 - 0xff
      13'hF8C: dout <= 8'b11111111; // 3980 : 255 - 0xff
      13'hF8D: dout <= 8'b11111111; // 3981 : 255 - 0xff
      13'hF8E: dout <= 8'b11111111; // 3982 : 255 - 0xff
      13'hF8F: dout <= 8'b11111111; // 3983 : 255 - 0xff
      13'hF90: dout <= 8'b11111111; // 3984 : 255 - 0xff -- Sprite 0xf9
      13'hF91: dout <= 8'b11111111; // 3985 : 255 - 0xff
      13'hF92: dout <= 8'b11111111; // 3986 : 255 - 0xff
      13'hF93: dout <= 8'b11111111; // 3987 : 255 - 0xff
      13'hF94: dout <= 8'b11111111; // 3988 : 255 - 0xff
      13'hF95: dout <= 8'b11111111; // 3989 : 255 - 0xff
      13'hF96: dout <= 8'b11111111; // 3990 : 255 - 0xff
      13'hF97: dout <= 8'b11111111; // 3991 : 255 - 0xff
      13'hF98: dout <= 8'b11111111; // 3992 : 255 - 0xff
      13'hF99: dout <= 8'b11111111; // 3993 : 255 - 0xff
      13'hF9A: dout <= 8'b11111111; // 3994 : 255 - 0xff
      13'hF9B: dout <= 8'b11111111; // 3995 : 255 - 0xff
      13'hF9C: dout <= 8'b11111111; // 3996 : 255 - 0xff
      13'hF9D: dout <= 8'b11111111; // 3997 : 255 - 0xff
      13'hF9E: dout <= 8'b11111111; // 3998 : 255 - 0xff
      13'hF9F: dout <= 8'b11111111; // 3999 : 255 - 0xff
      13'hFA0: dout <= 8'b11111111; // 4000 : 255 - 0xff -- Sprite 0xfa
      13'hFA1: dout <= 8'b11111111; // 4001 : 255 - 0xff
      13'hFA2: dout <= 8'b11111111; // 4002 : 255 - 0xff
      13'hFA3: dout <= 8'b11111111; // 4003 : 255 - 0xff
      13'hFA4: dout <= 8'b11111111; // 4004 : 255 - 0xff
      13'hFA5: dout <= 8'b11111111; // 4005 : 255 - 0xff
      13'hFA6: dout <= 8'b11111111; // 4006 : 255 - 0xff
      13'hFA7: dout <= 8'b11111111; // 4007 : 255 - 0xff
      13'hFA8: dout <= 8'b11111111; // 4008 : 255 - 0xff
      13'hFA9: dout <= 8'b11111111; // 4009 : 255 - 0xff
      13'hFAA: dout <= 8'b11111111; // 4010 : 255 - 0xff
      13'hFAB: dout <= 8'b11111111; // 4011 : 255 - 0xff
      13'hFAC: dout <= 8'b11111111; // 4012 : 255 - 0xff
      13'hFAD: dout <= 8'b11111111; // 4013 : 255 - 0xff
      13'hFAE: dout <= 8'b11111111; // 4014 : 255 - 0xff
      13'hFAF: dout <= 8'b11111111; // 4015 : 255 - 0xff
      13'hFB0: dout <= 8'b11111111; // 4016 : 255 - 0xff -- Sprite 0xfb
      13'hFB1: dout <= 8'b11111111; // 4017 : 255 - 0xff
      13'hFB2: dout <= 8'b11111111; // 4018 : 255 - 0xff
      13'hFB3: dout <= 8'b11111111; // 4019 : 255 - 0xff
      13'hFB4: dout <= 8'b11111111; // 4020 : 255 - 0xff
      13'hFB5: dout <= 8'b11111111; // 4021 : 255 - 0xff
      13'hFB6: dout <= 8'b11111111; // 4022 : 255 - 0xff
      13'hFB7: dout <= 8'b11111111; // 4023 : 255 - 0xff
      13'hFB8: dout <= 8'b11111111; // 4024 : 255 - 0xff
      13'hFB9: dout <= 8'b11111111; // 4025 : 255 - 0xff
      13'hFBA: dout <= 8'b11111111; // 4026 : 255 - 0xff
      13'hFBB: dout <= 8'b11111111; // 4027 : 255 - 0xff
      13'hFBC: dout <= 8'b11111111; // 4028 : 255 - 0xff
      13'hFBD: dout <= 8'b11111111; // 4029 : 255 - 0xff
      13'hFBE: dout <= 8'b11111111; // 4030 : 255 - 0xff
      13'hFBF: dout <= 8'b11111111; // 4031 : 255 - 0xff
      13'hFC0: dout <= 8'b11111111; // 4032 : 255 - 0xff -- Sprite 0xfc
      13'hFC1: dout <= 8'b11111111; // 4033 : 255 - 0xff
      13'hFC2: dout <= 8'b11111111; // 4034 : 255 - 0xff
      13'hFC3: dout <= 8'b11111111; // 4035 : 255 - 0xff
      13'hFC4: dout <= 8'b11111111; // 4036 : 255 - 0xff
      13'hFC5: dout <= 8'b11111111; // 4037 : 255 - 0xff
      13'hFC6: dout <= 8'b11111111; // 4038 : 255 - 0xff
      13'hFC7: dout <= 8'b11111111; // 4039 : 255 - 0xff
      13'hFC8: dout <= 8'b11111111; // 4040 : 255 - 0xff
      13'hFC9: dout <= 8'b11111111; // 4041 : 255 - 0xff
      13'hFCA: dout <= 8'b11111111; // 4042 : 255 - 0xff
      13'hFCB: dout <= 8'b11111111; // 4043 : 255 - 0xff
      13'hFCC: dout <= 8'b11111111; // 4044 : 255 - 0xff
      13'hFCD: dout <= 8'b11111111; // 4045 : 255 - 0xff
      13'hFCE: dout <= 8'b11111111; // 4046 : 255 - 0xff
      13'hFCF: dout <= 8'b11111111; // 4047 : 255 - 0xff
      13'hFD0: dout <= 8'b11111111; // 4048 : 255 - 0xff -- Sprite 0xfd
      13'hFD1: dout <= 8'b11111111; // 4049 : 255 - 0xff
      13'hFD2: dout <= 8'b11111111; // 4050 : 255 - 0xff
      13'hFD3: dout <= 8'b11111111; // 4051 : 255 - 0xff
      13'hFD4: dout <= 8'b11111111; // 4052 : 255 - 0xff
      13'hFD5: dout <= 8'b11111111; // 4053 : 255 - 0xff
      13'hFD6: dout <= 8'b11111111; // 4054 : 255 - 0xff
      13'hFD7: dout <= 8'b11111111; // 4055 : 255 - 0xff
      13'hFD8: dout <= 8'b11111111; // 4056 : 255 - 0xff
      13'hFD9: dout <= 8'b11111111; // 4057 : 255 - 0xff
      13'hFDA: dout <= 8'b11111111; // 4058 : 255 - 0xff
      13'hFDB: dout <= 8'b11111111; // 4059 : 255 - 0xff
      13'hFDC: dout <= 8'b11111111; // 4060 : 255 - 0xff
      13'hFDD: dout <= 8'b11111111; // 4061 : 255 - 0xff
      13'hFDE: dout <= 8'b11111111; // 4062 : 255 - 0xff
      13'hFDF: dout <= 8'b11111111; // 4063 : 255 - 0xff
      13'hFE0: dout <= 8'b11111111; // 4064 : 255 - 0xff -- Sprite 0xfe
      13'hFE1: dout <= 8'b11111111; // 4065 : 255 - 0xff
      13'hFE2: dout <= 8'b11111111; // 4066 : 255 - 0xff
      13'hFE3: dout <= 8'b11111111; // 4067 : 255 - 0xff
      13'hFE4: dout <= 8'b11111111; // 4068 : 255 - 0xff
      13'hFE5: dout <= 8'b11111111; // 4069 : 255 - 0xff
      13'hFE6: dout <= 8'b11111111; // 4070 : 255 - 0xff
      13'hFE7: dout <= 8'b11111111; // 4071 : 255 - 0xff
      13'hFE8: dout <= 8'b11111111; // 4072 : 255 - 0xff
      13'hFE9: dout <= 8'b11111111; // 4073 : 255 - 0xff
      13'hFEA: dout <= 8'b11111111; // 4074 : 255 - 0xff
      13'hFEB: dout <= 8'b11111111; // 4075 : 255 - 0xff
      13'hFEC: dout <= 8'b11111111; // 4076 : 255 - 0xff
      13'hFED: dout <= 8'b11111111; // 4077 : 255 - 0xff
      13'hFEE: dout <= 8'b11111111; // 4078 : 255 - 0xff
      13'hFEF: dout <= 8'b11111111; // 4079 : 255 - 0xff
      13'hFF0: dout <= 8'b11111111; // 4080 : 255 - 0xff -- Sprite 0xff
      13'hFF1: dout <= 8'b11111111; // 4081 : 255 - 0xff
      13'hFF2: dout <= 8'b11111111; // 4082 : 255 - 0xff
      13'hFF3: dout <= 8'b11111111; // 4083 : 255 - 0xff
      13'hFF4: dout <= 8'b11111111; // 4084 : 255 - 0xff
      13'hFF5: dout <= 8'b11111111; // 4085 : 255 - 0xff
      13'hFF6: dout <= 8'b11111111; // 4086 : 255 - 0xff
      13'hFF7: dout <= 8'b11111111; // 4087 : 255 - 0xff
      13'hFF8: dout <= 8'b11111111; // 4088 : 255 - 0xff
      13'hFF9: dout <= 8'b11111111; // 4089 : 255 - 0xff
      13'hFFA: dout <= 8'b11111111; // 4090 : 255 - 0xff
      13'hFFB: dout <= 8'b11111111; // 4091 : 255 - 0xff
      13'hFFC: dout <= 8'b11111111; // 4092 : 255 - 0xff
      13'hFFD: dout <= 8'b11111111; // 4093 : 255 - 0xff
      13'hFFE: dout <= 8'b11111111; // 4094 : 255 - 0xff
      13'hFFF: dout <= 8'b11111111; // 4095 : 255 - 0xff
          // Pattern Table 1---------
      13'h1000: dout <= 8'b00000000; // 4096 :   0 - 0x0 -- Background 0x0
      13'h1001: dout <= 8'b00000011; // 4097 :   3 - 0x3
      13'h1002: dout <= 8'b00001111; // 4098 :  15 - 0xf
      13'h1003: dout <= 8'b00011111; // 4099 :  31 - 0x1f
      13'h1004: dout <= 8'b00111111; // 4100 :  63 - 0x3f
      13'h1005: dout <= 8'b00111111; // 4101 :  63 - 0x3f
      13'h1006: dout <= 8'b01111111; // 4102 : 127 - 0x7f
      13'h1007: dout <= 8'b01111111; // 4103 : 127 - 0x7f
      13'h1008: dout <= 8'b00000000; // 4104 :   0 - 0x0
      13'h1009: dout <= 8'b00000000; // 4105 :   0 - 0x0
      13'h100A: dout <= 8'b00000000; // 4106 :   0 - 0x0
      13'h100B: dout <= 8'b00000000; // 4107 :   0 - 0x0
      13'h100C: dout <= 8'b00000000; // 4108 :   0 - 0x0
      13'h100D: dout <= 8'b00000000; // 4109 :   0 - 0x0
      13'h100E: dout <= 8'b00000000; // 4110 :   0 - 0x0
      13'h100F: dout <= 8'b00000000; // 4111 :   0 - 0x0
      13'h1010: dout <= 8'b00000000; // 4112 :   0 - 0x0 -- Background 0x1
      13'h1011: dout <= 8'b11000000; // 4113 : 192 - 0xc0
      13'h1012: dout <= 8'b11110000; // 4114 : 240 - 0xf0
      13'h1013: dout <= 8'b11111000; // 4115 : 248 - 0xf8
      13'h1014: dout <= 8'b11111000; // 4116 : 248 - 0xf8
      13'h1015: dout <= 8'b11111100; // 4117 : 252 - 0xfc
      13'h1016: dout <= 8'b11111100; // 4118 : 252 - 0xfc
      13'h1017: dout <= 8'b11111100; // 4119 : 252 - 0xfc
      13'h1018: dout <= 8'b00000000; // 4120 :   0 - 0x0
      13'h1019: dout <= 8'b00000000; // 4121 :   0 - 0x0
      13'h101A: dout <= 8'b00000000; // 4122 :   0 - 0x0
      13'h101B: dout <= 8'b00000000; // 4123 :   0 - 0x0
      13'h101C: dout <= 8'b00000000; // 4124 :   0 - 0x0
      13'h101D: dout <= 8'b00000000; // 4125 :   0 - 0x0
      13'h101E: dout <= 8'b00000000; // 4126 :   0 - 0x0
      13'h101F: dout <= 8'b00000000; // 4127 :   0 - 0x0
      13'h1020: dout <= 8'b00000000; // 4128 :   0 - 0x0 -- Background 0x2
      13'h1021: dout <= 8'b00000111; // 4129 :   7 - 0x7
      13'h1022: dout <= 8'b00011111; // 4130 :  31 - 0x1f
      13'h1023: dout <= 8'b00111111; // 4131 :  63 - 0x3f
      13'h1024: dout <= 8'b00111111; // 4132 :  63 - 0x3f
      13'h1025: dout <= 8'b00001111; // 4133 :  15 - 0xf
      13'h1026: dout <= 8'b00000011; // 4134 :   3 - 0x3
      13'h1027: dout <= 8'b00000000; // 4135 :   0 - 0x0
      13'h1028: dout <= 8'b00000000; // 4136 :   0 - 0x0
      13'h1029: dout <= 8'b00000000; // 4137 :   0 - 0x0
      13'h102A: dout <= 8'b00000000; // 4138 :   0 - 0x0
      13'h102B: dout <= 8'b00000000; // 4139 :   0 - 0x0
      13'h102C: dout <= 8'b00000000; // 4140 :   0 - 0x0
      13'h102D: dout <= 8'b00000000; // 4141 :   0 - 0x0
      13'h102E: dout <= 8'b00000000; // 4142 :   0 - 0x0
      13'h102F: dout <= 8'b00000000; // 4143 :   0 - 0x0
      13'h1030: dout <= 8'b00000000; // 4144 :   0 - 0x0 -- Background 0x3
      13'h1031: dout <= 8'b00000000; // 4145 :   0 - 0x0
      13'h1032: dout <= 8'b00000111; // 4146 :   7 - 0x7
      13'h1033: dout <= 8'b00011111; // 4147 :  31 - 0x1f
      13'h1034: dout <= 8'b00111111; // 4148 :  63 - 0x3f
      13'h1035: dout <= 8'b00111111; // 4149 :  63 - 0x3f
      13'h1036: dout <= 8'b01111111; // 4150 : 127 - 0x7f
      13'h1037: dout <= 8'b01111111; // 4151 : 127 - 0x7f
      13'h1038: dout <= 8'b00000000; // 4152 :   0 - 0x0
      13'h1039: dout <= 8'b00000000; // 4153 :   0 - 0x0
      13'h103A: dout <= 8'b00000000; // 4154 :   0 - 0x0
      13'h103B: dout <= 8'b00000000; // 4155 :   0 - 0x0
      13'h103C: dout <= 8'b00000000; // 4156 :   0 - 0x0
      13'h103D: dout <= 8'b00000000; // 4157 :   0 - 0x0
      13'h103E: dout <= 8'b00000000; // 4158 :   0 - 0x0
      13'h103F: dout <= 8'b00000000; // 4159 :   0 - 0x0
      13'h1040: dout <= 8'b01111110; // 4160 : 126 - 0x7e -- Background 0x4
      13'h1041: dout <= 8'b01111110; // 4161 : 126 - 0x7e
      13'h1042: dout <= 8'b01111100; // 4162 : 124 - 0x7c
      13'h1043: dout <= 8'b00111100; // 4163 :  60 - 0x3c
      13'h1044: dout <= 8'b00111000; // 4164 :  56 - 0x38
      13'h1045: dout <= 8'b00011000; // 4165 :  24 - 0x18
      13'h1046: dout <= 8'b00000000; // 4166 :   0 - 0x0
      13'h1047: dout <= 8'b00000000; // 4167 :   0 - 0x0
      13'h1048: dout <= 8'b00000000; // 4168 :   0 - 0x0
      13'h1049: dout <= 8'b00000000; // 4169 :   0 - 0x0
      13'h104A: dout <= 8'b00000000; // 4170 :   0 - 0x0
      13'h104B: dout <= 8'b00000000; // 4171 :   0 - 0x0
      13'h104C: dout <= 8'b00000000; // 4172 :   0 - 0x0
      13'h104D: dout <= 8'b00000000; // 4173 :   0 - 0x0
      13'h104E: dout <= 8'b00000000; // 4174 :   0 - 0x0
      13'h104F: dout <= 8'b00000000; // 4175 :   0 - 0x0
      13'h1050: dout <= 8'b00000000; // 4176 :   0 - 0x0 -- Background 0x5
      13'h1051: dout <= 8'b11000000; // 4177 : 192 - 0xc0
      13'h1052: dout <= 8'b11110000; // 4178 : 240 - 0xf0
      13'h1053: dout <= 8'b11111000; // 4179 : 248 - 0xf8
      13'h1054: dout <= 8'b11111000; // 4180 : 248 - 0xf8
      13'h1055: dout <= 8'b11111100; // 4181 : 252 - 0xfc
      13'h1056: dout <= 8'b01111100; // 4182 : 124 - 0x7c
      13'h1057: dout <= 8'b00111100; // 4183 :  60 - 0x3c
      13'h1058: dout <= 8'b00000000; // 4184 :   0 - 0x0
      13'h1059: dout <= 8'b00000000; // 4185 :   0 - 0x0
      13'h105A: dout <= 8'b00000000; // 4186 :   0 - 0x0
      13'h105B: dout <= 8'b00000000; // 4187 :   0 - 0x0
      13'h105C: dout <= 8'b00000000; // 4188 :   0 - 0x0
      13'h105D: dout <= 8'b00000000; // 4189 :   0 - 0x0
      13'h105E: dout <= 8'b00000000; // 4190 :   0 - 0x0
      13'h105F: dout <= 8'b00000000; // 4191 :   0 - 0x0
      13'h1060: dout <= 8'b00000000; // 4192 :   0 - 0x0 -- Background 0x6
      13'h1061: dout <= 8'b00000111; // 4193 :   7 - 0x7
      13'h1062: dout <= 8'b00000111; // 4194 :   7 - 0x7
      13'h1063: dout <= 8'b00000011; // 4195 :   3 - 0x3
      13'h1064: dout <= 8'b00000001; // 4196 :   1 - 0x1
      13'h1065: dout <= 8'b00000000; // 4197 :   0 - 0x0
      13'h1066: dout <= 8'b00000000; // 4198 :   0 - 0x0
      13'h1067: dout <= 8'b00000000; // 4199 :   0 - 0x0
      13'h1068: dout <= 8'b00000000; // 4200 :   0 - 0x0
      13'h1069: dout <= 8'b00000000; // 4201 :   0 - 0x0
      13'h106A: dout <= 8'b00000000; // 4202 :   0 - 0x0
      13'h106B: dout <= 8'b00000000; // 4203 :   0 - 0x0
      13'h106C: dout <= 8'b00000000; // 4204 :   0 - 0x0
      13'h106D: dout <= 8'b00000000; // 4205 :   0 - 0x0
      13'h106E: dout <= 8'b00000000; // 4206 :   0 - 0x0
      13'h106F: dout <= 8'b00000000; // 4207 :   0 - 0x0
      13'h1070: dout <= 8'b00000000; // 4208 :   0 - 0x0 -- Background 0x7
      13'h1071: dout <= 8'b00000000; // 4209 :   0 - 0x0
      13'h1072: dout <= 8'b00000111; // 4210 :   7 - 0x7
      13'h1073: dout <= 8'b00011111; // 4211 :  31 - 0x1f
      13'h1074: dout <= 8'b00111111; // 4212 :  63 - 0x3f
      13'h1075: dout <= 8'b00111111; // 4213 :  63 - 0x3f
      13'h1076: dout <= 8'b01111110; // 4214 : 126 - 0x7e
      13'h1077: dout <= 8'b01111100; // 4215 : 124 - 0x7c
      13'h1078: dout <= 8'b00000000; // 4216 :   0 - 0x0
      13'h1079: dout <= 8'b00000000; // 4217 :   0 - 0x0
      13'h107A: dout <= 8'b00000000; // 4218 :   0 - 0x0
      13'h107B: dout <= 8'b00000000; // 4219 :   0 - 0x0
      13'h107C: dout <= 8'b00000000; // 4220 :   0 - 0x0
      13'h107D: dout <= 8'b00000000; // 4221 :   0 - 0x0
      13'h107E: dout <= 8'b00000000; // 4222 :   0 - 0x0
      13'h107F: dout <= 8'b00000000; // 4223 :   0 - 0x0
      13'h1080: dout <= 8'b01111000; // 4224 : 120 - 0x78 -- Background 0x8
      13'h1081: dout <= 8'b01110000; // 4225 : 112 - 0x70
      13'h1082: dout <= 8'b01100000; // 4226 :  96 - 0x60
      13'h1083: dout <= 8'b00000000; // 4227 :   0 - 0x0
      13'h1084: dout <= 8'b00000000; // 4228 :   0 - 0x0
      13'h1085: dout <= 8'b00000000; // 4229 :   0 - 0x0
      13'h1086: dout <= 8'b00000000; // 4230 :   0 - 0x0
      13'h1087: dout <= 8'b00000000; // 4231 :   0 - 0x0
      13'h1088: dout <= 8'b00000000; // 4232 :   0 - 0x0
      13'h1089: dout <= 8'b00000000; // 4233 :   0 - 0x0
      13'h108A: dout <= 8'b00000000; // 4234 :   0 - 0x0
      13'h108B: dout <= 8'b00000000; // 4235 :   0 - 0x0
      13'h108C: dout <= 8'b00000000; // 4236 :   0 - 0x0
      13'h108D: dout <= 8'b00000000; // 4237 :   0 - 0x0
      13'h108E: dout <= 8'b00000000; // 4238 :   0 - 0x0
      13'h108F: dout <= 8'b00000000; // 4239 :   0 - 0x0
      13'h1090: dout <= 8'b00000000; // 4240 :   0 - 0x0 -- Background 0x9
      13'h1091: dout <= 8'b00000000; // 4241 :   0 - 0x0
      13'h1092: dout <= 8'b00000000; // 4242 :   0 - 0x0
      13'h1093: dout <= 8'b00000000; // 4243 :   0 - 0x0
      13'h1094: dout <= 8'b00000000; // 4244 :   0 - 0x0
      13'h1095: dout <= 8'b01000000; // 4245 :  64 - 0x40
      13'h1096: dout <= 8'b11110000; // 4246 : 240 - 0xf0
      13'h1097: dout <= 8'b11111000; // 4247 : 248 - 0xf8
      13'h1098: dout <= 8'b00000000; // 4248 :   0 - 0x0
      13'h1099: dout <= 8'b00000000; // 4249 :   0 - 0x0
      13'h109A: dout <= 8'b00000000; // 4250 :   0 - 0x0
      13'h109B: dout <= 8'b00000000; // 4251 :   0 - 0x0
      13'h109C: dout <= 8'b00000000; // 4252 :   0 - 0x0
      13'h109D: dout <= 8'b00000000; // 4253 :   0 - 0x0
      13'h109E: dout <= 8'b00000000; // 4254 :   0 - 0x0
      13'h109F: dout <= 8'b00000000; // 4255 :   0 - 0x0
      13'h10A0: dout <= 8'b11111110; // 4256 : 254 - 0xfe -- Background 0xa
      13'h10A1: dout <= 8'b01111111; // 4257 : 127 - 0x7f
      13'h10A2: dout <= 8'b01111111; // 4258 : 127 - 0x7f
      13'h10A3: dout <= 8'b00111111; // 4259 :  63 - 0x3f
      13'h10A4: dout <= 8'b00001110; // 4260 :  14 - 0xe
      13'h10A5: dout <= 8'b00000000; // 4261 :   0 - 0x0
      13'h10A6: dout <= 8'b00000000; // 4262 :   0 - 0x0
      13'h10A7: dout <= 8'b00000000; // 4263 :   0 - 0x0
      13'h10A8: dout <= 8'b00000000; // 4264 :   0 - 0x0
      13'h10A9: dout <= 8'b00000000; // 4265 :   0 - 0x0
      13'h10AA: dout <= 8'b00000000; // 4266 :   0 - 0x0
      13'h10AB: dout <= 8'b00000000; // 4267 :   0 - 0x0
      13'h10AC: dout <= 8'b00000000; // 4268 :   0 - 0x0
      13'h10AD: dout <= 8'b00000000; // 4269 :   0 - 0x0
      13'h10AE: dout <= 8'b00000000; // 4270 :   0 - 0x0
      13'h10AF: dout <= 8'b00000000; // 4271 :   0 - 0x0
      13'h10B0: dout <= 8'b00000000; // 4272 :   0 - 0x0 -- Background 0xb
      13'h10B1: dout <= 8'b00000000; // 4273 :   0 - 0x0
      13'h10B2: dout <= 8'b00000000; // 4274 :   0 - 0x0
      13'h10B3: dout <= 8'b00000000; // 4275 :   0 - 0x0
      13'h10B4: dout <= 8'b00000000; // 4276 :   0 - 0x0
      13'h10B5: dout <= 8'b00000000; // 4277 :   0 - 0x0
      13'h10B6: dout <= 8'b00000000; // 4278 :   0 - 0x0
      13'h10B7: dout <= 8'b11100000; // 4279 : 224 - 0xe0
      13'h10B8: dout <= 8'b00000000; // 4280 :   0 - 0x0
      13'h10B9: dout <= 8'b00000000; // 4281 :   0 - 0x0
      13'h10BA: dout <= 8'b00000000; // 4282 :   0 - 0x0
      13'h10BB: dout <= 8'b00000000; // 4283 :   0 - 0x0
      13'h10BC: dout <= 8'b00000000; // 4284 :   0 - 0x0
      13'h10BD: dout <= 8'b00000000; // 4285 :   0 - 0x0
      13'h10BE: dout <= 8'b00000000; // 4286 :   0 - 0x0
      13'h10BF: dout <= 8'b00000000; // 4287 :   0 - 0x0
      13'h10C0: dout <= 8'b11111100; // 4288 : 252 - 0xfc -- Background 0xc
      13'h10C1: dout <= 8'b11111111; // 4289 : 255 - 0xff
      13'h10C2: dout <= 8'b01111111; // 4290 : 127 - 0x7f
      13'h10C3: dout <= 8'b00111111; // 4291 :  63 - 0x3f
      13'h10C4: dout <= 8'b00001110; // 4292 :  14 - 0xe
      13'h10C5: dout <= 8'b00000000; // 4293 :   0 - 0x0
      13'h10C6: dout <= 8'b00000000; // 4294 :   0 - 0x0
      13'h10C7: dout <= 8'b00000000; // 4295 :   0 - 0x0
      13'h10C8: dout <= 8'b00000000; // 4296 :   0 - 0x0
      13'h10C9: dout <= 8'b00000000; // 4297 :   0 - 0x0
      13'h10CA: dout <= 8'b00000000; // 4298 :   0 - 0x0
      13'h10CB: dout <= 8'b00000000; // 4299 :   0 - 0x0
      13'h10CC: dout <= 8'b00000000; // 4300 :   0 - 0x0
      13'h10CD: dout <= 8'b00000000; // 4301 :   0 - 0x0
      13'h10CE: dout <= 8'b00000000; // 4302 :   0 - 0x0
      13'h10CF: dout <= 8'b00000000; // 4303 :   0 - 0x0
      13'h10D0: dout <= 8'b11110000; // 4304 : 240 - 0xf0 -- Background 0xd
      13'h10D1: dout <= 8'b11111111; // 4305 : 255 - 0xff
      13'h10D2: dout <= 8'b11111111; // 4306 : 255 - 0xff
      13'h10D3: dout <= 8'b01111111; // 4307 : 127 - 0x7f
      13'h10D4: dout <= 8'b00011110; // 4308 :  30 - 0x1e
      13'h10D5: dout <= 8'b00000000; // 4309 :   0 - 0x0
      13'h10D6: dout <= 8'b00000000; // 4310 :   0 - 0x0
      13'h10D7: dout <= 8'b00000000; // 4311 :   0 - 0x0
      13'h10D8: dout <= 8'b00000000; // 4312 :   0 - 0x0
      13'h10D9: dout <= 8'b00000000; // 4313 :   0 - 0x0
      13'h10DA: dout <= 8'b00000000; // 4314 :   0 - 0x0
      13'h10DB: dout <= 8'b00000000; // 4315 :   0 - 0x0
      13'h10DC: dout <= 8'b00000000; // 4316 :   0 - 0x0
      13'h10DD: dout <= 8'b00000000; // 4317 :   0 - 0x0
      13'h10DE: dout <= 8'b00000000; // 4318 :   0 - 0x0
      13'h10DF: dout <= 8'b00000000; // 4319 :   0 - 0x0
      13'h10E0: dout <= 8'b00000000; // 4320 :   0 - 0x0 -- Background 0xe
      13'h10E1: dout <= 8'b00001111; // 4321 :  15 - 0xf
      13'h10E2: dout <= 8'b11111111; // 4322 : 255 - 0xff
      13'h10E3: dout <= 8'b11111111; // 4323 : 255 - 0xff
      13'h10E4: dout <= 8'b01111111; // 4324 : 127 - 0x7f
      13'h10E5: dout <= 8'b00011110; // 4325 :  30 - 0x1e
      13'h10E6: dout <= 8'b00000000; // 4326 :   0 - 0x0
      13'h10E7: dout <= 8'b00000000; // 4327 :   0 - 0x0
      13'h10E8: dout <= 8'b00000000; // 4328 :   0 - 0x0
      13'h10E9: dout <= 8'b00000000; // 4329 :   0 - 0x0
      13'h10EA: dout <= 8'b00000000; // 4330 :   0 - 0x0
      13'h10EB: dout <= 8'b00000000; // 4331 :   0 - 0x0
      13'h10EC: dout <= 8'b00000000; // 4332 :   0 - 0x0
      13'h10ED: dout <= 8'b00000000; // 4333 :   0 - 0x0
      13'h10EE: dout <= 8'b00000000; // 4334 :   0 - 0x0
      13'h10EF: dout <= 8'b00000000; // 4335 :   0 - 0x0
      13'h10F0: dout <= 8'b00000000; // 4336 :   0 - 0x0 -- Background 0xf
      13'h10F1: dout <= 8'b00000011; // 4337 :   3 - 0x3
      13'h10F2: dout <= 8'b00001111; // 4338 :  15 - 0xf
      13'h10F3: dout <= 8'b01111111; // 4339 : 127 - 0x7f
      13'h10F4: dout <= 8'b11111111; // 4340 : 255 - 0xff
      13'h10F5: dout <= 8'b01111110; // 4341 : 126 - 0x7e
      13'h10F6: dout <= 8'b00011100; // 4342 :  28 - 0x1c
      13'h10F7: dout <= 8'b00000000; // 4343 :   0 - 0x0
      13'h10F8: dout <= 8'b00000000; // 4344 :   0 - 0x0
      13'h10F9: dout <= 8'b00000000; // 4345 :   0 - 0x0
      13'h10FA: dout <= 8'b00000000; // 4346 :   0 - 0x0
      13'h10FB: dout <= 8'b00000000; // 4347 :   0 - 0x0
      13'h10FC: dout <= 8'b00000000; // 4348 :   0 - 0x0
      13'h10FD: dout <= 8'b00000000; // 4349 :   0 - 0x0
      13'h10FE: dout <= 8'b00000000; // 4350 :   0 - 0x0
      13'h10FF: dout <= 8'b00000000; // 4351 :   0 - 0x0
      13'h1100: dout <= 8'b00000000; // 4352 :   0 - 0x0 -- Background 0x10
      13'h1101: dout <= 8'b00000001; // 4353 :   1 - 0x1
      13'h1102: dout <= 8'b00000011; // 4354 :   3 - 0x3
      13'h1103: dout <= 8'b00001111; // 4355 :  15 - 0xf
      13'h1104: dout <= 8'b00011111; // 4356 :  31 - 0x1f
      13'h1105: dout <= 8'b01111111; // 4357 : 127 - 0x7f
      13'h1106: dout <= 8'b01111110; // 4358 : 126 - 0x7e
      13'h1107: dout <= 8'b00111100; // 4359 :  60 - 0x3c
      13'h1108: dout <= 8'b00000000; // 4360 :   0 - 0x0
      13'h1109: dout <= 8'b00000000; // 4361 :   0 - 0x0
      13'h110A: dout <= 8'b00000000; // 4362 :   0 - 0x0
      13'h110B: dout <= 8'b00000000; // 4363 :   0 - 0x0
      13'h110C: dout <= 8'b00000000; // 4364 :   0 - 0x0
      13'h110D: dout <= 8'b00000000; // 4365 :   0 - 0x0
      13'h110E: dout <= 8'b00000000; // 4366 :   0 - 0x0
      13'h110F: dout <= 8'b00000000; // 4367 :   0 - 0x0
      13'h1110: dout <= 8'b00000000; // 4368 :   0 - 0x0 -- Background 0x11
      13'h1111: dout <= 8'b00000001; // 4369 :   1 - 0x1
      13'h1112: dout <= 8'b00000011; // 4370 :   3 - 0x3
      13'h1113: dout <= 8'b00000111; // 4371 :   7 - 0x7
      13'h1114: dout <= 8'b00000111; // 4372 :   7 - 0x7
      13'h1115: dout <= 8'b00001111; // 4373 :  15 - 0xf
      13'h1116: dout <= 8'b00011111; // 4374 :  31 - 0x1f
      13'h1117: dout <= 8'b00001110; // 4375 :  14 - 0xe
      13'h1118: dout <= 8'b00000000; // 4376 :   0 - 0x0
      13'h1119: dout <= 8'b00000000; // 4377 :   0 - 0x0
      13'h111A: dout <= 8'b00000000; // 4378 :   0 - 0x0
      13'h111B: dout <= 8'b00000000; // 4379 :   0 - 0x0
      13'h111C: dout <= 8'b00000000; // 4380 :   0 - 0x0
      13'h111D: dout <= 8'b00000000; // 4381 :   0 - 0x0
      13'h111E: dout <= 8'b00000000; // 4382 :   0 - 0x0
      13'h111F: dout <= 8'b00000000; // 4383 :   0 - 0x0
      13'h1120: dout <= 8'b00000000; // 4384 :   0 - 0x0 -- Background 0x12
      13'h1121: dout <= 8'b00000000; // 4385 :   0 - 0x0
      13'h1122: dout <= 8'b00000001; // 4386 :   1 - 0x1
      13'h1123: dout <= 8'b00000011; // 4387 :   3 - 0x3
      13'h1124: dout <= 8'b00000011; // 4388 :   3 - 0x3
      13'h1125: dout <= 8'b00000011; // 4389 :   3 - 0x3
      13'h1126: dout <= 8'b00000111; // 4390 :   7 - 0x7
      13'h1127: dout <= 8'b00000010; // 4391 :   2 - 0x2
      13'h1128: dout <= 8'b00000000; // 4392 :   0 - 0x0
      13'h1129: dout <= 8'b00000000; // 4393 :   0 - 0x0
      13'h112A: dout <= 8'b00000000; // 4394 :   0 - 0x0
      13'h112B: dout <= 8'b00000000; // 4395 :   0 - 0x0
      13'h112C: dout <= 8'b00000000; // 4396 :   0 - 0x0
      13'h112D: dout <= 8'b00000000; // 4397 :   0 - 0x0
      13'h112E: dout <= 8'b00000000; // 4398 :   0 - 0x0
      13'h112F: dout <= 8'b00000000; // 4399 :   0 - 0x0
      13'h1130: dout <= 8'b00000000; // 4400 :   0 - 0x0 -- Background 0x13
      13'h1131: dout <= 8'b00000000; // 4401 :   0 - 0x0
      13'h1132: dout <= 8'b00000001; // 4402 :   1 - 0x1
      13'h1133: dout <= 8'b00000001; // 4403 :   1 - 0x1
      13'h1134: dout <= 8'b00000001; // 4404 :   1 - 0x1
      13'h1135: dout <= 8'b00000001; // 4405 :   1 - 0x1
      13'h1136: dout <= 8'b00000001; // 4406 :   1 - 0x1
      13'h1137: dout <= 8'b00000001; // 4407 :   1 - 0x1
      13'h1138: dout <= 8'b00000000; // 4408 :   0 - 0x0
      13'h1139: dout <= 8'b00000000; // 4409 :   0 - 0x0
      13'h113A: dout <= 8'b00000000; // 4410 :   0 - 0x0
      13'h113B: dout <= 8'b00000000; // 4411 :   0 - 0x0
      13'h113C: dout <= 8'b00000000; // 4412 :   0 - 0x0
      13'h113D: dout <= 8'b00000000; // 4413 :   0 - 0x0
      13'h113E: dout <= 8'b00000000; // 4414 :   0 - 0x0
      13'h113F: dout <= 8'b00000000; // 4415 :   0 - 0x0
      13'h1140: dout <= 8'b00000000; // 4416 :   0 - 0x0 -- Background 0x14
      13'h1141: dout <= 8'b00000000; // 4417 :   0 - 0x0
      13'h1142: dout <= 8'b00000000; // 4418 :   0 - 0x0
      13'h1143: dout <= 8'b00000000; // 4419 :   0 - 0x0
      13'h1144: dout <= 8'b00000000; // 4420 :   0 - 0x0
      13'h1145: dout <= 8'b00000000; // 4421 :   0 - 0x0
      13'h1146: dout <= 8'b00000100; // 4422 :   4 - 0x4
      13'h1147: dout <= 8'b00000010; // 4423 :   2 - 0x2
      13'h1148: dout <= 8'b00000000; // 4424 :   0 - 0x0
      13'h1149: dout <= 8'b00000000; // 4425 :   0 - 0x0
      13'h114A: dout <= 8'b00000000; // 4426 :   0 - 0x0
      13'h114B: dout <= 8'b00000000; // 4427 :   0 - 0x0
      13'h114C: dout <= 8'b00000000; // 4428 :   0 - 0x0
      13'h114D: dout <= 8'b00000000; // 4429 :   0 - 0x0
      13'h114E: dout <= 8'b00000000; // 4430 :   0 - 0x0
      13'h114F: dout <= 8'b00000000; // 4431 :   0 - 0x0
      13'h1150: dout <= 8'b00000000; // 4432 :   0 - 0x0 -- Background 0x15
      13'h1151: dout <= 8'b00000000; // 4433 :   0 - 0x0
      13'h1152: dout <= 8'b00000000; // 4434 :   0 - 0x0
      13'h1153: dout <= 8'b00000000; // 4435 :   0 - 0x0
      13'h1154: dout <= 8'b00000000; // 4436 :   0 - 0x0
      13'h1155: dout <= 8'b00000000; // 4437 :   0 - 0x0
      13'h1156: dout <= 8'b00100000; // 4438 :  32 - 0x20
      13'h1157: dout <= 8'b01001000; // 4439 :  72 - 0x48
      13'h1158: dout <= 8'b00000000; // 4440 :   0 - 0x0
      13'h1159: dout <= 8'b00000000; // 4441 :   0 - 0x0
      13'h115A: dout <= 8'b00000000; // 4442 :   0 - 0x0
      13'h115B: dout <= 8'b00000000; // 4443 :   0 - 0x0
      13'h115C: dout <= 8'b00000000; // 4444 :   0 - 0x0
      13'h115D: dout <= 8'b00000000; // 4445 :   0 - 0x0
      13'h115E: dout <= 8'b00000000; // 4446 :   0 - 0x0
      13'h115F: dout <= 8'b00000000; // 4447 :   0 - 0x0
      13'h1160: dout <= 8'b00010000; // 4448 :  16 - 0x10 -- Background 0x16
      13'h1161: dout <= 8'b00001000; // 4449 :   8 - 0x8
      13'h1162: dout <= 8'b00000000; // 4450 :   0 - 0x0
      13'h1163: dout <= 8'b00110000; // 4451 :  48 - 0x30
      13'h1164: dout <= 8'b00000000; // 4452 :   0 - 0x0
      13'h1165: dout <= 8'b00001000; // 4453 :   8 - 0x8
      13'h1166: dout <= 8'b00010010; // 4454 :  18 - 0x12
      13'h1167: dout <= 8'b00000100; // 4455 :   4 - 0x4
      13'h1168: dout <= 8'b00000000; // 4456 :   0 - 0x0
      13'h1169: dout <= 8'b00000000; // 4457 :   0 - 0x0
      13'h116A: dout <= 8'b00000000; // 4458 :   0 - 0x0
      13'h116B: dout <= 8'b00000000; // 4459 :   0 - 0x0
      13'h116C: dout <= 8'b00000000; // 4460 :   0 - 0x0
      13'h116D: dout <= 8'b00000000; // 4461 :   0 - 0x0
      13'h116E: dout <= 8'b00000000; // 4462 :   0 - 0x0
      13'h116F: dout <= 8'b00000000; // 4463 :   0 - 0x0
      13'h1170: dout <= 8'b00010000; // 4464 :  16 - 0x10 -- Background 0x17
      13'h1171: dout <= 8'b00000000; // 4465 :   0 - 0x0
      13'h1172: dout <= 8'b00001100; // 4466 :  12 - 0xc
      13'h1173: dout <= 8'b00000000; // 4467 :   0 - 0x0
      13'h1174: dout <= 8'b00010000; // 4468 :  16 - 0x10
      13'h1175: dout <= 8'b00001000; // 4469 :   8 - 0x8
      13'h1176: dout <= 8'b01000000; // 4470 :  64 - 0x40
      13'h1177: dout <= 8'b00100000; // 4471 :  32 - 0x20
      13'h1178: dout <= 8'b00000000; // 4472 :   0 - 0x0
      13'h1179: dout <= 8'b00000000; // 4473 :   0 - 0x0
      13'h117A: dout <= 8'b00000000; // 4474 :   0 - 0x0
      13'h117B: dout <= 8'b00000000; // 4475 :   0 - 0x0
      13'h117C: dout <= 8'b00000000; // 4476 :   0 - 0x0
      13'h117D: dout <= 8'b00000000; // 4477 :   0 - 0x0
      13'h117E: dout <= 8'b00000000; // 4478 :   0 - 0x0
      13'h117F: dout <= 8'b00000000; // 4479 :   0 - 0x0
      13'h1180: dout <= 8'b00000000; // 4480 :   0 - 0x0 -- Background 0x18
      13'h1181: dout <= 8'b00000000; // 4481 :   0 - 0x0
      13'h1182: dout <= 8'b00000011; // 4482 :   3 - 0x3
      13'h1183: dout <= 8'b00000011; // 4483 :   3 - 0x3
      13'h1184: dout <= 8'b00000001; // 4484 :   1 - 0x1
      13'h1185: dout <= 8'b00100001; // 4485 :  33 - 0x21
      13'h1186: dout <= 8'b00100001; // 4486 :  33 - 0x21
      13'h1187: dout <= 8'b01110011; // 4487 : 115 - 0x73
      13'h1188: dout <= 8'b00000000; // 4488 :   0 - 0x0
      13'h1189: dout <= 8'b00000000; // 4489 :   0 - 0x0
      13'h118A: dout <= 8'b00000011; // 4490 :   3 - 0x3
      13'h118B: dout <= 8'b00000011; // 4491 :   3 - 0x3
      13'h118C: dout <= 8'b00010011; // 4492 :  19 - 0x13
      13'h118D: dout <= 8'b00111111; // 4493 :  63 - 0x3f
      13'h118E: dout <= 8'b00111111; // 4494 :  63 - 0x3f
      13'h118F: dout <= 8'b01111111; // 4495 : 127 - 0x7f
      13'h1190: dout <= 8'b01111111; // 4496 : 127 - 0x7f -- Background 0x19
      13'h1191: dout <= 8'b01111111; // 4497 : 127 - 0x7f
      13'h1192: dout <= 8'b01111111; // 4498 : 127 - 0x7f
      13'h1193: dout <= 8'b01111111; // 4499 : 127 - 0x7f
      13'h1194: dout <= 8'b01101110; // 4500 : 110 - 0x6e
      13'h1195: dout <= 8'b01000110; // 4501 :  70 - 0x46
      13'h1196: dout <= 8'b00000000; // 4502 :   0 - 0x0
      13'h1197: dout <= 8'b00000000; // 4503 :   0 - 0x0
      13'h1198: dout <= 8'b01111111; // 4504 : 127 - 0x7f
      13'h1199: dout <= 8'b01111111; // 4505 : 127 - 0x7f
      13'h119A: dout <= 8'b01111111; // 4506 : 127 - 0x7f
      13'h119B: dout <= 8'b01111111; // 4507 : 127 - 0x7f
      13'h119C: dout <= 8'b01101110; // 4508 : 110 - 0x6e
      13'h119D: dout <= 8'b01000110; // 4509 :  70 - 0x46
      13'h119E: dout <= 8'b00000000; // 4510 :   0 - 0x0
      13'h119F: dout <= 8'b00000000; // 4511 :   0 - 0x0
      13'h11A0: dout <= 8'b01111111; // 4512 : 127 - 0x7f -- Background 0x1a
      13'h11A1: dout <= 8'b01111111; // 4513 : 127 - 0x7f
      13'h11A2: dout <= 8'b01111111; // 4514 : 127 - 0x7f
      13'h11A3: dout <= 8'b01111111; // 4515 : 127 - 0x7f
      13'h11A4: dout <= 8'b01111011; // 4516 : 123 - 0x7b
      13'h11A5: dout <= 8'b00110001; // 4517 :  49 - 0x31
      13'h11A6: dout <= 8'b00000000; // 4518 :   0 - 0x0
      13'h11A7: dout <= 8'b00000000; // 4519 :   0 - 0x0
      13'h11A8: dout <= 8'b01111111; // 4520 : 127 - 0x7f
      13'h11A9: dout <= 8'b01111111; // 4521 : 127 - 0x7f
      13'h11AA: dout <= 8'b01111111; // 4522 : 127 - 0x7f
      13'h11AB: dout <= 8'b01111111; // 4523 : 127 - 0x7f
      13'h11AC: dout <= 8'b01111011; // 4524 : 123 - 0x7b
      13'h11AD: dout <= 8'b00110001; // 4525 :  49 - 0x31
      13'h11AE: dout <= 8'b00000000; // 4526 :   0 - 0x0
      13'h11AF: dout <= 8'b00000000; // 4527 :   0 - 0x0
      13'h11B0: dout <= 8'b00000000; // 4528 :   0 - 0x0 -- Background 0x1b
      13'h11B1: dout <= 8'b00000011; // 4529 :   3 - 0x3
      13'h11B2: dout <= 8'b00001111; // 4530 :  15 - 0xf
      13'h11B3: dout <= 8'b00011111; // 4531 :  31 - 0x1f
      13'h11B4: dout <= 8'b00100111; // 4532 :  39 - 0x27
      13'h11B5: dout <= 8'b00000011; // 4533 :   3 - 0x3
      13'h11B6: dout <= 8'b00000011; // 4534 :   3 - 0x3
      13'h11B7: dout <= 8'b01000011; // 4535 :  67 - 0x43
      13'h11B8: dout <= 8'b00000000; // 4536 :   0 - 0x0
      13'h11B9: dout <= 8'b00000011; // 4537 :   3 - 0x3
      13'h11BA: dout <= 8'b00001111; // 4538 :  15 - 0xf
      13'h11BB: dout <= 8'b00011111; // 4539 :  31 - 0x1f
      13'h11BC: dout <= 8'b00111111; // 4540 :  63 - 0x3f
      13'h11BD: dout <= 8'b00111111; // 4541 :  63 - 0x3f
      13'h11BE: dout <= 8'b00001111; // 4542 :  15 - 0xf
      13'h11BF: dout <= 8'b01001111; // 4543 :  79 - 0x4f
      13'h11C0: dout <= 8'b00000000; // 4544 :   0 - 0x0 -- Background 0x1c
      13'h11C1: dout <= 8'b11000000; // 4545 : 192 - 0xc0
      13'h11C2: dout <= 8'b11110000; // 4546 : 240 - 0xf0
      13'h11C3: dout <= 8'b11111000; // 4547 : 248 - 0xf8
      13'h11C4: dout <= 8'b10011100; // 4548 : 156 - 0x9c
      13'h11C5: dout <= 8'b00001100; // 4549 :  12 - 0xc
      13'h11C6: dout <= 8'b00001100; // 4550 :  12 - 0xc
      13'h11C7: dout <= 8'b00001110; // 4551 :  14 - 0xe
      13'h11C8: dout <= 8'b00000000; // 4552 :   0 - 0x0
      13'h11C9: dout <= 8'b11000000; // 4553 : 192 - 0xc0
      13'h11CA: dout <= 8'b11110000; // 4554 : 240 - 0xf0
      13'h11CB: dout <= 8'b11111000; // 4555 : 248 - 0xf8
      13'h11CC: dout <= 8'b11111100; // 4556 : 252 - 0xfc
      13'h11CD: dout <= 8'b11111100; // 4557 : 252 - 0xfc
      13'h11CE: dout <= 8'b00111100; // 4558 :  60 - 0x3c
      13'h11CF: dout <= 8'b00111110; // 4559 :  62 - 0x3e
      13'h11D0: dout <= 8'b01100111; // 4560 : 103 - 0x67 -- Background 0x1d
      13'h11D1: dout <= 8'b01111111; // 4561 : 127 - 0x7f
      13'h11D2: dout <= 8'b01111111; // 4562 : 127 - 0x7f
      13'h11D3: dout <= 8'b01111111; // 4563 : 127 - 0x7f
      13'h11D4: dout <= 8'b01101110; // 4564 : 110 - 0x6e
      13'h11D5: dout <= 8'b01000110; // 4565 :  70 - 0x46
      13'h11D6: dout <= 8'b00000000; // 4566 :   0 - 0x0
      13'h11D7: dout <= 8'b00000000; // 4567 :   0 - 0x0
      13'h11D8: dout <= 8'b01111111; // 4568 : 127 - 0x7f
      13'h11D9: dout <= 8'b01111111; // 4569 : 127 - 0x7f
      13'h11DA: dout <= 8'b01111111; // 4570 : 127 - 0x7f
      13'h11DB: dout <= 8'b01111111; // 4571 : 127 - 0x7f
      13'h11DC: dout <= 8'b01101110; // 4572 : 110 - 0x6e
      13'h11DD: dout <= 8'b01000110; // 4573 :  70 - 0x46
      13'h11DE: dout <= 8'b00000000; // 4574 :   0 - 0x0
      13'h11DF: dout <= 8'b00000000; // 4575 :   0 - 0x0
      13'h11E0: dout <= 8'b01100111; // 4576 : 103 - 0x67 -- Background 0x1e
      13'h11E1: dout <= 8'b01111111; // 4577 : 127 - 0x7f
      13'h11E2: dout <= 8'b01111111; // 4578 : 127 - 0x7f
      13'h11E3: dout <= 8'b01111111; // 4579 : 127 - 0x7f
      13'h11E4: dout <= 8'b01111011; // 4580 : 123 - 0x7b
      13'h11E5: dout <= 8'b00110001; // 4581 :  49 - 0x31
      13'h11E6: dout <= 8'b00000000; // 4582 :   0 - 0x0
      13'h11E7: dout <= 8'b00000000; // 4583 :   0 - 0x0
      13'h11E8: dout <= 8'b01111111; // 4584 : 127 - 0x7f
      13'h11E9: dout <= 8'b01111111; // 4585 : 127 - 0x7f
      13'h11EA: dout <= 8'b01111111; // 4586 : 127 - 0x7f
      13'h11EB: dout <= 8'b01111111; // 4587 : 127 - 0x7f
      13'h11EC: dout <= 8'b01111011; // 4588 : 123 - 0x7b
      13'h11ED: dout <= 8'b00110001; // 4589 :  49 - 0x31
      13'h11EE: dout <= 8'b00000000; // 4590 :   0 - 0x0
      13'h11EF: dout <= 8'b00000000; // 4591 :   0 - 0x0
      13'h11F0: dout <= 8'b10011110; // 4592 : 158 - 0x9e -- Background 0x1f
      13'h11F1: dout <= 8'b11111110; // 4593 : 254 - 0xfe
      13'h11F2: dout <= 8'b11111110; // 4594 : 254 - 0xfe
      13'h11F3: dout <= 8'b11111110; // 4595 : 254 - 0xfe
      13'h11F4: dout <= 8'b01110110; // 4596 : 118 - 0x76
      13'h11F5: dout <= 8'b01100010; // 4597 :  98 - 0x62
      13'h11F6: dout <= 8'b00000000; // 4598 :   0 - 0x0
      13'h11F7: dout <= 8'b00000000; // 4599 :   0 - 0x0
      13'h11F8: dout <= 8'b11111110; // 4600 : 254 - 0xfe
      13'h11F9: dout <= 8'b11111110; // 4601 : 254 - 0xfe
      13'h11FA: dout <= 8'b11111110; // 4602 : 254 - 0xfe
      13'h11FB: dout <= 8'b11111110; // 4603 : 254 - 0xfe
      13'h11FC: dout <= 8'b01110110; // 4604 : 118 - 0x76
      13'h11FD: dout <= 8'b01100010; // 4605 :  98 - 0x62
      13'h11FE: dout <= 8'b00000000; // 4606 :   0 - 0x0
      13'h11FF: dout <= 8'b00000000; // 4607 :   0 - 0x0
      13'h1200: dout <= 8'b10011110; // 4608 : 158 - 0x9e -- Background 0x20
      13'h1201: dout <= 8'b11111110; // 4609 : 254 - 0xfe
      13'h1202: dout <= 8'b11111110; // 4610 : 254 - 0xfe
      13'h1203: dout <= 8'b11111110; // 4611 : 254 - 0xfe
      13'h1204: dout <= 8'b11011110; // 4612 : 222 - 0xde
      13'h1205: dout <= 8'b10001100; // 4613 : 140 - 0x8c
      13'h1206: dout <= 8'b00000000; // 4614 :   0 - 0x0
      13'h1207: dout <= 8'b00000000; // 4615 :   0 - 0x0
      13'h1208: dout <= 8'b11111110; // 4616 : 254 - 0xfe
      13'h1209: dout <= 8'b11111110; // 4617 : 254 - 0xfe
      13'h120A: dout <= 8'b11111110; // 4618 : 254 - 0xfe
      13'h120B: dout <= 8'b11111110; // 4619 : 254 - 0xfe
      13'h120C: dout <= 8'b11011110; // 4620 : 222 - 0xde
      13'h120D: dout <= 8'b10001100; // 4621 : 140 - 0x8c
      13'h120E: dout <= 8'b00000000; // 4622 :   0 - 0x0
      13'h120F: dout <= 8'b00000000; // 4623 :   0 - 0x0
      13'h1210: dout <= 8'b00000000; // 4624 :   0 - 0x0 -- Background 0x21
      13'h1211: dout <= 8'b00000011; // 4625 :   3 - 0x3
      13'h1212: dout <= 8'b00001111; // 4626 :  15 - 0xf
      13'h1213: dout <= 8'b00011111; // 4627 :  31 - 0x1f
      13'h1214: dout <= 8'b00111111; // 4628 :  63 - 0x3f
      13'h1215: dout <= 8'b00110011; // 4629 :  51 - 0x33
      13'h1216: dout <= 8'b00100001; // 4630 :  33 - 0x21
      13'h1217: dout <= 8'b01100001; // 4631 :  97 - 0x61
      13'h1218: dout <= 8'b00000000; // 4632 :   0 - 0x0
      13'h1219: dout <= 8'b00000011; // 4633 :   3 - 0x3
      13'h121A: dout <= 8'b00001111; // 4634 :  15 - 0xf
      13'h121B: dout <= 8'b00011111; // 4635 :  31 - 0x1f
      13'h121C: dout <= 8'b00111111; // 4636 :  63 - 0x3f
      13'h121D: dout <= 8'b00111111; // 4637 :  63 - 0x3f
      13'h121E: dout <= 8'b00111111; // 4638 :  63 - 0x3f
      13'h121F: dout <= 8'b01111111; // 4639 : 127 - 0x7f
      13'h1220: dout <= 8'b01100001; // 4640 :  97 - 0x61 -- Background 0x22
      13'h1221: dout <= 8'b01110011; // 4641 : 115 - 0x73
      13'h1222: dout <= 8'b01111111; // 4642 : 127 - 0x7f
      13'h1223: dout <= 8'b01111111; // 4643 : 127 - 0x7f
      13'h1224: dout <= 8'b01101110; // 4644 : 110 - 0x6e
      13'h1225: dout <= 8'b01000110; // 4645 :  70 - 0x46
      13'h1226: dout <= 8'b00000000; // 4646 :   0 - 0x0
      13'h1227: dout <= 8'b00000000; // 4647 :   0 - 0x0
      13'h1228: dout <= 8'b01110011; // 4648 : 115 - 0x73
      13'h1229: dout <= 8'b01110011; // 4649 : 115 - 0x73
      13'h122A: dout <= 8'b01111111; // 4650 : 127 - 0x7f
      13'h122B: dout <= 8'b01111111; // 4651 : 127 - 0x7f
      13'h122C: dout <= 8'b01101110; // 4652 : 110 - 0x6e
      13'h122D: dout <= 8'b01000110; // 4653 :  70 - 0x46
      13'h122E: dout <= 8'b00000000; // 4654 :   0 - 0x0
      13'h122F: dout <= 8'b00000000; // 4655 :   0 - 0x0
      13'h1230: dout <= 8'b01100001; // 4656 :  97 - 0x61 -- Background 0x23
      13'h1231: dout <= 8'b01110011; // 4657 : 115 - 0x73
      13'h1232: dout <= 8'b01111111; // 4658 : 127 - 0x7f
      13'h1233: dout <= 8'b01111111; // 4659 : 127 - 0x7f
      13'h1234: dout <= 8'b01110111; // 4660 : 119 - 0x77
      13'h1235: dout <= 8'b00100011; // 4661 :  35 - 0x23
      13'h1236: dout <= 8'b00000000; // 4662 :   0 - 0x0
      13'h1237: dout <= 8'b00000000; // 4663 :   0 - 0x0
      13'h1238: dout <= 8'b01110011; // 4664 : 115 - 0x73
      13'h1239: dout <= 8'b01110011; // 4665 : 115 - 0x73
      13'h123A: dout <= 8'b01111111; // 4666 : 127 - 0x7f
      13'h123B: dout <= 8'b01111111; // 4667 : 127 - 0x7f
      13'h123C: dout <= 8'b01110111; // 4668 : 119 - 0x77
      13'h123D: dout <= 8'b00100011; // 4669 :  35 - 0x23
      13'h123E: dout <= 8'b00000000; // 4670 :   0 - 0x0
      13'h123F: dout <= 8'b00000000; // 4671 :   0 - 0x0
      13'h1240: dout <= 8'b00000000; // 4672 :   0 - 0x0 -- Background 0x24
      13'h1241: dout <= 8'b00000011; // 4673 :   3 - 0x3
      13'h1242: dout <= 8'b00001111; // 4674 :  15 - 0xf
      13'h1243: dout <= 8'b00011111; // 4675 :  31 - 0x1f
      13'h1244: dout <= 8'b00111111; // 4676 :  63 - 0x3f
      13'h1245: dout <= 8'b00111111; // 4677 :  63 - 0x3f
      13'h1246: dout <= 8'b00111111; // 4678 :  63 - 0x3f
      13'h1247: dout <= 8'b01111111; // 4679 : 127 - 0x7f
      13'h1248: dout <= 8'b00000000; // 4680 :   0 - 0x0
      13'h1249: dout <= 8'b00000000; // 4681 :   0 - 0x0
      13'h124A: dout <= 8'b00000000; // 4682 :   0 - 0x0
      13'h124B: dout <= 8'b00000000; // 4683 :   0 - 0x0
      13'h124C: dout <= 8'b00000000; // 4684 :   0 - 0x0
      13'h124D: dout <= 8'b00000110; // 4685 :   6 - 0x6
      13'h124E: dout <= 8'b00000110; // 4686 :   6 - 0x6
      13'h124F: dout <= 8'b00000000; // 4687 :   0 - 0x0
      13'h1250: dout <= 8'b01111111; // 4688 : 127 - 0x7f -- Background 0x25
      13'h1251: dout <= 8'b01111111; // 4689 : 127 - 0x7f
      13'h1252: dout <= 8'b01111111; // 4690 : 127 - 0x7f
      13'h1253: dout <= 8'b01111111; // 4691 : 127 - 0x7f
      13'h1254: dout <= 8'b01101110; // 4692 : 110 - 0x6e
      13'h1255: dout <= 8'b01000110; // 4693 :  70 - 0x46
      13'h1256: dout <= 8'b00000000; // 4694 :   0 - 0x0
      13'h1257: dout <= 8'b00000000; // 4695 :   0 - 0x0
      13'h1258: dout <= 8'b00000000; // 4696 :   0 - 0x0
      13'h1259: dout <= 8'b00011001; // 4697 :  25 - 0x19
      13'h125A: dout <= 8'b00100110; // 4698 :  38 - 0x26
      13'h125B: dout <= 8'b00000000; // 4699 :   0 - 0x0
      13'h125C: dout <= 8'b00000000; // 4700 :   0 - 0x0
      13'h125D: dout <= 8'b00000000; // 4701 :   0 - 0x0
      13'h125E: dout <= 8'b00000000; // 4702 :   0 - 0x0
      13'h125F: dout <= 8'b00000000; // 4703 :   0 - 0x0
      13'h1260: dout <= 8'b01111111; // 4704 : 127 - 0x7f -- Background 0x26
      13'h1261: dout <= 8'b01111111; // 4705 : 127 - 0x7f
      13'h1262: dout <= 8'b01111111; // 4706 : 127 - 0x7f
      13'h1263: dout <= 8'b01111111; // 4707 : 127 - 0x7f
      13'h1264: dout <= 8'b01111011; // 4708 : 123 - 0x7b
      13'h1265: dout <= 8'b00110001; // 4709 :  49 - 0x31
      13'h1266: dout <= 8'b00000000; // 4710 :   0 - 0x0
      13'h1267: dout <= 8'b00000000; // 4711 :   0 - 0x0
      13'h1268: dout <= 8'b00000000; // 4712 :   0 - 0x0
      13'h1269: dout <= 8'b00011001; // 4713 :  25 - 0x19
      13'h126A: dout <= 8'b00100110; // 4714 :  38 - 0x26
      13'h126B: dout <= 8'b00000000; // 4715 :   0 - 0x0
      13'h126C: dout <= 8'b00000000; // 4716 :   0 - 0x0
      13'h126D: dout <= 8'b00000000; // 4717 :   0 - 0x0
      13'h126E: dout <= 8'b00000000; // 4718 :   0 - 0x0
      13'h126F: dout <= 8'b00000000; // 4719 :   0 - 0x0
      13'h1270: dout <= 8'b00000000; // 4720 :   0 - 0x0 -- Background 0x27
      13'h1271: dout <= 8'b00000000; // 4721 :   0 - 0x0
      13'h1272: dout <= 8'b00000000; // 4722 :   0 - 0x0
      13'h1273: dout <= 8'b00000000; // 4723 :   0 - 0x0
      13'h1274: dout <= 8'b00000000; // 4724 :   0 - 0x0
      13'h1275: dout <= 8'b00000000; // 4725 :   0 - 0x0
      13'h1276: dout <= 8'b00000000; // 4726 :   0 - 0x0
      13'h1277: dout <= 8'b00000000; // 4727 :   0 - 0x0
      13'h1278: dout <= 8'b00000000; // 4728 :   0 - 0x0
      13'h1279: dout <= 8'b00001100; // 4729 :  12 - 0xc
      13'h127A: dout <= 8'b00010010; // 4730 :  18 - 0x12
      13'h127B: dout <= 8'b00010010; // 4731 :  18 - 0x12
      13'h127C: dout <= 8'b00011110; // 4732 :  30 - 0x1e
      13'h127D: dout <= 8'b00001100; // 4733 :  12 - 0xc
      13'h127E: dout <= 8'b00000000; // 4734 :   0 - 0x0
      13'h127F: dout <= 8'b00000000; // 4735 :   0 - 0x0
      13'h1280: dout <= 8'b00000000; // 4736 :   0 - 0x0 -- Background 0x28
      13'h1281: dout <= 8'b00000000; // 4737 :   0 - 0x0
      13'h1282: dout <= 8'b00000000; // 4738 :   0 - 0x0
      13'h1283: dout <= 8'b00000000; // 4739 :   0 - 0x0
      13'h1284: dout <= 8'b00000000; // 4740 :   0 - 0x0
      13'h1285: dout <= 8'b00000000; // 4741 :   0 - 0x0
      13'h1286: dout <= 8'b00000000; // 4742 :   0 - 0x0
      13'h1287: dout <= 8'b00000000; // 4743 :   0 - 0x0
      13'h1288: dout <= 8'b00000000; // 4744 :   0 - 0x0
      13'h1289: dout <= 8'b00000000; // 4745 :   0 - 0x0
      13'h128A: dout <= 8'b00000000; // 4746 :   0 - 0x0
      13'h128B: dout <= 8'b00000000; // 4747 :   0 - 0x0
      13'h128C: dout <= 8'b00000000; // 4748 :   0 - 0x0
      13'h128D: dout <= 8'b00111000; // 4749 :  56 - 0x38
      13'h128E: dout <= 8'b01001101; // 4750 :  77 - 0x4d
      13'h128F: dout <= 8'b01001101; // 4751 :  77 - 0x4d
      13'h1290: dout <= 8'b00000000; // 4752 :   0 - 0x0 -- Background 0x29
      13'h1291: dout <= 8'b00000000; // 4753 :   0 - 0x0
      13'h1292: dout <= 8'b00000000; // 4754 :   0 - 0x0
      13'h1293: dout <= 8'b00000000; // 4755 :   0 - 0x0
      13'h1294: dout <= 8'b00000000; // 4756 :   0 - 0x0
      13'h1295: dout <= 8'b00000000; // 4757 :   0 - 0x0
      13'h1296: dout <= 8'b00000000; // 4758 :   0 - 0x0
      13'h1297: dout <= 8'b00000000; // 4759 :   0 - 0x0
      13'h1298: dout <= 8'b00000000; // 4760 :   0 - 0x0
      13'h1299: dout <= 8'b00000000; // 4761 :   0 - 0x0
      13'h129A: dout <= 8'b00000000; // 4762 :   0 - 0x0
      13'h129B: dout <= 8'b00000000; // 4763 :   0 - 0x0
      13'h129C: dout <= 8'b00000000; // 4764 :   0 - 0x0
      13'h129D: dout <= 8'b11100000; // 4765 : 224 - 0xe0
      13'h129E: dout <= 8'b00110000; // 4766 :  48 - 0x30
      13'h129F: dout <= 8'b00110000; // 4767 :  48 - 0x30
      13'h12A0: dout <= 8'b00000000; // 4768 :   0 - 0x0 -- Background 0x2a
      13'h12A1: dout <= 8'b00000000; // 4769 :   0 - 0x0
      13'h12A2: dout <= 8'b00000000; // 4770 :   0 - 0x0
      13'h12A3: dout <= 8'b00000000; // 4771 :   0 - 0x0
      13'h12A4: dout <= 8'b00000000; // 4772 :   0 - 0x0
      13'h12A5: dout <= 8'b00000000; // 4773 :   0 - 0x0
      13'h12A6: dout <= 8'b00000000; // 4774 :   0 - 0x0
      13'h12A7: dout <= 8'b00000000; // 4775 :   0 - 0x0
      13'h12A8: dout <= 8'b00111000; // 4776 :  56 - 0x38
      13'h12A9: dout <= 8'b00000000; // 4777 :   0 - 0x0
      13'h12AA: dout <= 8'b00000000; // 4778 :   0 - 0x0
      13'h12AB: dout <= 8'b00000000; // 4779 :   0 - 0x0
      13'h12AC: dout <= 8'b00000000; // 4780 :   0 - 0x0
      13'h12AD: dout <= 8'b00000000; // 4781 :   0 - 0x0
      13'h12AE: dout <= 8'b00000000; // 4782 :   0 - 0x0
      13'h12AF: dout <= 8'b00000000; // 4783 :   0 - 0x0
      13'h12B0: dout <= 8'b00000000; // 4784 :   0 - 0x0 -- Background 0x2b
      13'h12B1: dout <= 8'b00000000; // 4785 :   0 - 0x0
      13'h12B2: dout <= 8'b00000000; // 4786 :   0 - 0x0
      13'h12B3: dout <= 8'b00000000; // 4787 :   0 - 0x0
      13'h12B4: dout <= 8'b00000000; // 4788 :   0 - 0x0
      13'h12B5: dout <= 8'b00000000; // 4789 :   0 - 0x0
      13'h12B6: dout <= 8'b00000000; // 4790 :   0 - 0x0
      13'h12B7: dout <= 8'b00000000; // 4791 :   0 - 0x0
      13'h12B8: dout <= 8'b11100000; // 4792 : 224 - 0xe0
      13'h12B9: dout <= 8'b00000000; // 4793 :   0 - 0x0
      13'h12BA: dout <= 8'b00000000; // 4794 :   0 - 0x0
      13'h12BB: dout <= 8'b00000000; // 4795 :   0 - 0x0
      13'h12BC: dout <= 8'b00000000; // 4796 :   0 - 0x0
      13'h12BD: dout <= 8'b00000000; // 4797 :   0 - 0x0
      13'h12BE: dout <= 8'b00000000; // 4798 :   0 - 0x0
      13'h12BF: dout <= 8'b00000000; // 4799 :   0 - 0x0
      13'h12C0: dout <= 8'b00000000; // 4800 :   0 - 0x0 -- Background 0x2c
      13'h12C1: dout <= 8'b00000000; // 4801 :   0 - 0x0
      13'h12C2: dout <= 8'b00000000; // 4802 :   0 - 0x0
      13'h12C3: dout <= 8'b00000000; // 4803 :   0 - 0x0
      13'h12C4: dout <= 8'b00000000; // 4804 :   0 - 0x0
      13'h12C5: dout <= 8'b00000000; // 4805 :   0 - 0x0
      13'h12C6: dout <= 8'b00000000; // 4806 :   0 - 0x0
      13'h12C7: dout <= 8'b00000000; // 4807 :   0 - 0x0
      13'h12C8: dout <= 8'b00000000; // 4808 :   0 - 0x0
      13'h12C9: dout <= 8'b00000000; // 4809 :   0 - 0x0
      13'h12CA: dout <= 8'b00000000; // 4810 :   0 - 0x0
      13'h12CB: dout <= 8'b00000000; // 4811 :   0 - 0x0
      13'h12CC: dout <= 8'b00000000; // 4812 :   0 - 0x0
      13'h12CD: dout <= 8'b00000000; // 4813 :   0 - 0x0
      13'h12CE: dout <= 8'b00001100; // 4814 :  12 - 0xc
      13'h12CF: dout <= 8'b00011110; // 4815 :  30 - 0x1e
      13'h12D0: dout <= 8'b00000000; // 4816 :   0 - 0x0 -- Background 0x2d
      13'h12D1: dout <= 8'b00000000; // 4817 :   0 - 0x0
      13'h12D2: dout <= 8'b00000000; // 4818 :   0 - 0x0
      13'h12D3: dout <= 8'b00000000; // 4819 :   0 - 0x0
      13'h12D4: dout <= 8'b00000000; // 4820 :   0 - 0x0
      13'h12D5: dout <= 8'b00000000; // 4821 :   0 - 0x0
      13'h12D6: dout <= 8'b00000000; // 4822 :   0 - 0x0
      13'h12D7: dout <= 8'b00000000; // 4823 :   0 - 0x0
      13'h12D8: dout <= 8'b00010010; // 4824 :  18 - 0x12
      13'h12D9: dout <= 8'b00010010; // 4825 :  18 - 0x12
      13'h12DA: dout <= 8'b00001100; // 4826 :  12 - 0xc
      13'h12DB: dout <= 8'b00000000; // 4827 :   0 - 0x0
      13'h12DC: dout <= 8'b00000000; // 4828 :   0 - 0x0
      13'h12DD: dout <= 8'b00000000; // 4829 :   0 - 0x0
      13'h12DE: dout <= 8'b00000000; // 4830 :   0 - 0x0
      13'h12DF: dout <= 8'b00000000; // 4831 :   0 - 0x0
      13'h12E0: dout <= 8'b00000000; // 4832 :   0 - 0x0 -- Background 0x2e
      13'h12E1: dout <= 8'b00000000; // 4833 :   0 - 0x0
      13'h12E2: dout <= 8'b00000000; // 4834 :   0 - 0x0
      13'h12E3: dout <= 8'b00000000; // 4835 :   0 - 0x0
      13'h12E4: dout <= 8'b00000000; // 4836 :   0 - 0x0
      13'h12E5: dout <= 8'b00000000; // 4837 :   0 - 0x0
      13'h12E6: dout <= 8'b00000000; // 4838 :   0 - 0x0
      13'h12E7: dout <= 8'b00000000; // 4839 :   0 - 0x0
      13'h12E8: dout <= 8'b00000000; // 4840 :   0 - 0x0
      13'h12E9: dout <= 8'b00000000; // 4841 :   0 - 0x0
      13'h12EA: dout <= 8'b00000000; // 4842 :   0 - 0x0
      13'h12EB: dout <= 8'b00010001; // 4843 :  17 - 0x11
      13'h12EC: dout <= 8'b00110010; // 4844 :  50 - 0x32
      13'h12ED: dout <= 8'b00010010; // 4845 :  18 - 0x12
      13'h12EE: dout <= 8'b00010010; // 4846 :  18 - 0x12
      13'h12EF: dout <= 8'b00010010; // 4847 :  18 - 0x12
      13'h12F0: dout <= 8'b00000000; // 4848 :   0 - 0x0 -- Background 0x2f
      13'h12F1: dout <= 8'b00000000; // 4849 :   0 - 0x0
      13'h12F2: dout <= 8'b00000000; // 4850 :   0 - 0x0
      13'h12F3: dout <= 8'b00000000; // 4851 :   0 - 0x0
      13'h12F4: dout <= 8'b00000000; // 4852 :   0 - 0x0
      13'h12F5: dout <= 8'b00000000; // 4853 :   0 - 0x0
      13'h12F6: dout <= 8'b00000000; // 4854 :   0 - 0x0
      13'h12F7: dout <= 8'b00000000; // 4855 :   0 - 0x0
      13'h12F8: dout <= 8'b00000000; // 4856 :   0 - 0x0
      13'h12F9: dout <= 8'b00000000; // 4857 :   0 - 0x0
      13'h12FA: dout <= 8'b00000000; // 4858 :   0 - 0x0
      13'h12FB: dout <= 8'b10001100; // 4859 : 140 - 0x8c
      13'h12FC: dout <= 8'b01010010; // 4860 :  82 - 0x52
      13'h12FD: dout <= 8'b01010010; // 4861 :  82 - 0x52
      13'h12FE: dout <= 8'b01010010; // 4862 :  82 - 0x52
      13'h12FF: dout <= 8'b01010010; // 4863 :  82 - 0x52
      13'h1300: dout <= 8'b00000000; // 4864 :   0 - 0x0 -- Background 0x30
      13'h1301: dout <= 8'b00000000; // 4865 :   0 - 0x0
      13'h1302: dout <= 8'b00000000; // 4866 :   0 - 0x0
      13'h1303: dout <= 8'b00000000; // 4867 :   0 - 0x0
      13'h1304: dout <= 8'b00000000; // 4868 :   0 - 0x0
      13'h1305: dout <= 8'b00000000; // 4869 :   0 - 0x0
      13'h1306: dout <= 8'b00000000; // 4870 :   0 - 0x0
      13'h1307: dout <= 8'b00000000; // 4871 :   0 - 0x0
      13'h1308: dout <= 8'b00010010; // 4872 :  18 - 0x12
      13'h1309: dout <= 8'b00111001; // 4873 :  57 - 0x39
      13'h130A: dout <= 8'b00000000; // 4874 :   0 - 0x0
      13'h130B: dout <= 8'b00000000; // 4875 :   0 - 0x0
      13'h130C: dout <= 8'b00000000; // 4876 :   0 - 0x0
      13'h130D: dout <= 8'b00000000; // 4877 :   0 - 0x0
      13'h130E: dout <= 8'b00000000; // 4878 :   0 - 0x0
      13'h130F: dout <= 8'b00000000; // 4879 :   0 - 0x0
      13'h1310: dout <= 8'b00000000; // 4880 :   0 - 0x0 -- Background 0x31
      13'h1311: dout <= 8'b00000000; // 4881 :   0 - 0x0
      13'h1312: dout <= 8'b00000000; // 4882 :   0 - 0x0
      13'h1313: dout <= 8'b00000000; // 4883 :   0 - 0x0
      13'h1314: dout <= 8'b00000000; // 4884 :   0 - 0x0
      13'h1315: dout <= 8'b00000000; // 4885 :   0 - 0x0
      13'h1316: dout <= 8'b00000000; // 4886 :   0 - 0x0
      13'h1317: dout <= 8'b00000000; // 4887 :   0 - 0x0
      13'h1318: dout <= 8'b01010010; // 4888 :  82 - 0x52
      13'h1319: dout <= 8'b10001100; // 4889 : 140 - 0x8c
      13'h131A: dout <= 8'b00000000; // 4890 :   0 - 0x0
      13'h131B: dout <= 8'b00000000; // 4891 :   0 - 0x0
      13'h131C: dout <= 8'b00000000; // 4892 :   0 - 0x0
      13'h131D: dout <= 8'b00000000; // 4893 :   0 - 0x0
      13'h131E: dout <= 8'b00000000; // 4894 :   0 - 0x0
      13'h131F: dout <= 8'b00000000; // 4895 :   0 - 0x0
      13'h1320: dout <= 8'b00000000; // 4896 :   0 - 0x0 -- Background 0x32
      13'h1321: dout <= 8'b00000000; // 4897 :   0 - 0x0
      13'h1322: dout <= 8'b00000000; // 4898 :   0 - 0x0
      13'h1323: dout <= 8'b00000000; // 4899 :   0 - 0x0
      13'h1324: dout <= 8'b00000000; // 4900 :   0 - 0x0
      13'h1325: dout <= 8'b00000000; // 4901 :   0 - 0x0
      13'h1326: dout <= 8'b00000000; // 4902 :   0 - 0x0
      13'h1327: dout <= 8'b00000000; // 4903 :   0 - 0x0
      13'h1328: dout <= 8'b00000000; // 4904 :   0 - 0x0
      13'h1329: dout <= 8'b00000000; // 4905 :   0 - 0x0
      13'h132A: dout <= 8'b00000000; // 4906 :   0 - 0x0
      13'h132B: dout <= 8'b01110001; // 4907 : 113 - 0x71
      13'h132C: dout <= 8'b10001010; // 4908 : 138 - 0x8a
      13'h132D: dout <= 8'b00001010; // 4909 :  10 - 0xa
      13'h132E: dout <= 8'b00010010; // 4910 :  18 - 0x12
      13'h132F: dout <= 8'b00100010; // 4911 :  34 - 0x22
      13'h1330: dout <= 8'b00000000; // 4912 :   0 - 0x0 -- Background 0x33
      13'h1331: dout <= 8'b00000000; // 4913 :   0 - 0x0
      13'h1332: dout <= 8'b00000000; // 4914 :   0 - 0x0
      13'h1333: dout <= 8'b00000000; // 4915 :   0 - 0x0
      13'h1334: dout <= 8'b00000000; // 4916 :   0 - 0x0
      13'h1335: dout <= 8'b00000000; // 4917 :   0 - 0x0
      13'h1336: dout <= 8'b00000000; // 4918 :   0 - 0x0
      13'h1337: dout <= 8'b00000000; // 4919 :   0 - 0x0
      13'h1338: dout <= 8'b01000010; // 4920 :  66 - 0x42
      13'h1339: dout <= 8'b11111001; // 4921 : 249 - 0xf9
      13'h133A: dout <= 8'b00000000; // 4922 :   0 - 0x0
      13'h133B: dout <= 8'b00000000; // 4923 :   0 - 0x0
      13'h133C: dout <= 8'b00000000; // 4924 :   0 - 0x0
      13'h133D: dout <= 8'b00000000; // 4925 :   0 - 0x0
      13'h133E: dout <= 8'b00000000; // 4926 :   0 - 0x0
      13'h133F: dout <= 8'b00000000; // 4927 :   0 - 0x0
      13'h1340: dout <= 8'b00000000; // 4928 :   0 - 0x0 -- Background 0x34
      13'h1341: dout <= 8'b00000000; // 4929 :   0 - 0x0
      13'h1342: dout <= 8'b00000000; // 4930 :   0 - 0x0
      13'h1343: dout <= 8'b00000000; // 4931 :   0 - 0x0
      13'h1344: dout <= 8'b00000000; // 4932 :   0 - 0x0
      13'h1345: dout <= 8'b00000000; // 4933 :   0 - 0x0
      13'h1346: dout <= 8'b00000000; // 4934 :   0 - 0x0
      13'h1347: dout <= 8'b00000000; // 4935 :   0 - 0x0
      13'h1348: dout <= 8'b00000000; // 4936 :   0 - 0x0
      13'h1349: dout <= 8'b00000000; // 4937 :   0 - 0x0
      13'h134A: dout <= 8'b00000000; // 4938 :   0 - 0x0
      13'h134B: dout <= 8'b00110001; // 4939 :  49 - 0x31
      13'h134C: dout <= 8'b01001010; // 4940 :  74 - 0x4a
      13'h134D: dout <= 8'b00001010; // 4941 :  10 - 0xa
      13'h134E: dout <= 8'b00110010; // 4942 :  50 - 0x32
      13'h134F: dout <= 8'b00001010; // 4943 :  10 - 0xa
      13'h1350: dout <= 8'b00000000; // 4944 :   0 - 0x0 -- Background 0x35
      13'h1351: dout <= 8'b00000000; // 4945 :   0 - 0x0
      13'h1352: dout <= 8'b00000000; // 4946 :   0 - 0x0
      13'h1353: dout <= 8'b00000000; // 4947 :   0 - 0x0
      13'h1354: dout <= 8'b00000000; // 4948 :   0 - 0x0
      13'h1355: dout <= 8'b00000000; // 4949 :   0 - 0x0
      13'h1356: dout <= 8'b00000000; // 4950 :   0 - 0x0
      13'h1357: dout <= 8'b00000000; // 4951 :   0 - 0x0
      13'h1358: dout <= 8'b01001010; // 4952 :  74 - 0x4a
      13'h1359: dout <= 8'b00110001; // 4953 :  49 - 0x31
      13'h135A: dout <= 8'b00000000; // 4954 :   0 - 0x0
      13'h135B: dout <= 8'b00000000; // 4955 :   0 - 0x0
      13'h135C: dout <= 8'b00000000; // 4956 :   0 - 0x0
      13'h135D: dout <= 8'b00000000; // 4957 :   0 - 0x0
      13'h135E: dout <= 8'b00000000; // 4958 :   0 - 0x0
      13'h135F: dout <= 8'b00000000; // 4959 :   0 - 0x0
      13'h1360: dout <= 8'b00000000; // 4960 :   0 - 0x0 -- Background 0x36
      13'h1361: dout <= 8'b00000000; // 4961 :   0 - 0x0
      13'h1362: dout <= 8'b00000000; // 4962 :   0 - 0x0
      13'h1363: dout <= 8'b00000000; // 4963 :   0 - 0x0
      13'h1364: dout <= 8'b00000000; // 4964 :   0 - 0x0
      13'h1365: dout <= 8'b00000000; // 4965 :   0 - 0x0
      13'h1366: dout <= 8'b00000000; // 4966 :   0 - 0x0
      13'h1367: dout <= 8'b00000000; // 4967 :   0 - 0x0
      13'h1368: dout <= 8'b00000000; // 4968 :   0 - 0x0
      13'h1369: dout <= 8'b00000000; // 4969 :   0 - 0x0
      13'h136A: dout <= 8'b00000000; // 4970 :   0 - 0x0
      13'h136B: dout <= 8'b00010001; // 4971 :  17 - 0x11
      13'h136C: dout <= 8'b00110010; // 4972 :  50 - 0x32
      13'h136D: dout <= 8'b01010010; // 4973 :  82 - 0x52
      13'h136E: dout <= 8'b10010010; // 4974 : 146 - 0x92
      13'h136F: dout <= 8'b11111010; // 4975 : 250 - 0xfa
      13'h1370: dout <= 8'b00000000; // 4976 :   0 - 0x0 -- Background 0x37
      13'h1371: dout <= 8'b00000000; // 4977 :   0 - 0x0
      13'h1372: dout <= 8'b00000000; // 4978 :   0 - 0x0
      13'h1373: dout <= 8'b00000000; // 4979 :   0 - 0x0
      13'h1374: dout <= 8'b00000000; // 4980 :   0 - 0x0
      13'h1375: dout <= 8'b00000000; // 4981 :   0 - 0x0
      13'h1376: dout <= 8'b00000000; // 4982 :   0 - 0x0
      13'h1377: dout <= 8'b00000000; // 4983 :   0 - 0x0
      13'h1378: dout <= 8'b00010010; // 4984 :  18 - 0x12
      13'h1379: dout <= 8'b00010001; // 4985 :  17 - 0x11
      13'h137A: dout <= 8'b00000000; // 4986 :   0 - 0x0
      13'h137B: dout <= 8'b00000000; // 4987 :   0 - 0x0
      13'h137C: dout <= 8'b00000000; // 4988 :   0 - 0x0
      13'h137D: dout <= 8'b00000000; // 4989 :   0 - 0x0
      13'h137E: dout <= 8'b00000000; // 4990 :   0 - 0x0
      13'h137F: dout <= 8'b00000000; // 4991 :   0 - 0x0
      13'h1380: dout <= 8'b00000000; // 4992 :   0 - 0x0 -- Background 0x38
      13'h1381: dout <= 8'b00000000; // 4993 :   0 - 0x0
      13'h1382: dout <= 8'b00000000; // 4994 :   0 - 0x0
      13'h1383: dout <= 8'b00000000; // 4995 :   0 - 0x0
      13'h1384: dout <= 8'b00000000; // 4996 :   0 - 0x0
      13'h1385: dout <= 8'b00000000; // 4997 :   0 - 0x0
      13'h1386: dout <= 8'b00000000; // 4998 :   0 - 0x0
      13'h1387: dout <= 8'b00000000; // 4999 :   0 - 0x0
      13'h1388: dout <= 8'b00000000; // 5000 :   0 - 0x0
      13'h1389: dout <= 8'b00000000; // 5001 :   0 - 0x0
      13'h138A: dout <= 8'b00000000; // 5002 :   0 - 0x0
      13'h138B: dout <= 8'b01110001; // 5003 : 113 - 0x71
      13'h138C: dout <= 8'b01000010; // 5004 :  66 - 0x42
      13'h138D: dout <= 8'b01000010; // 5005 :  66 - 0x42
      13'h138E: dout <= 8'b01110010; // 5006 : 114 - 0x72
      13'h138F: dout <= 8'b00001010; // 5007 :  10 - 0xa
      13'h1390: dout <= 8'b00000000; // 5008 :   0 - 0x0 -- Background 0x39
      13'h1391: dout <= 8'b00000000; // 5009 :   0 - 0x0
      13'h1392: dout <= 8'b00000000; // 5010 :   0 - 0x0
      13'h1393: dout <= 8'b00000000; // 5011 :   0 - 0x0
      13'h1394: dout <= 8'b00000000; // 5012 :   0 - 0x0
      13'h1395: dout <= 8'b00000000; // 5013 :   0 - 0x0
      13'h1396: dout <= 8'b00000000; // 5014 :   0 - 0x0
      13'h1397: dout <= 8'b00000000; // 5015 :   0 - 0x0
      13'h1398: dout <= 8'b00001010; // 5016 :  10 - 0xa
      13'h1399: dout <= 8'b01110001; // 5017 : 113 - 0x71
      13'h139A: dout <= 8'b00000000; // 5018 :   0 - 0x0
      13'h139B: dout <= 8'b00000000; // 5019 :   0 - 0x0
      13'h139C: dout <= 8'b00000000; // 5020 :   0 - 0x0
      13'h139D: dout <= 8'b00000000; // 5021 :   0 - 0x0
      13'h139E: dout <= 8'b00000000; // 5022 :   0 - 0x0
      13'h139F: dout <= 8'b00000000; // 5023 :   0 - 0x0
      13'h13A0: dout <= 8'b00000000; // 5024 :   0 - 0x0 -- Background 0x3a
      13'h13A1: dout <= 8'b00000000; // 5025 :   0 - 0x0
      13'h13A2: dout <= 8'b00000000; // 5026 :   0 - 0x0
      13'h13A3: dout <= 8'b00000000; // 5027 :   0 - 0x0
      13'h13A4: dout <= 8'b00000000; // 5028 :   0 - 0x0
      13'h13A5: dout <= 8'b00000000; // 5029 :   0 - 0x0
      13'h13A6: dout <= 8'b00000000; // 5030 :   0 - 0x0
      13'h13A7: dout <= 8'b00000000; // 5031 :   0 - 0x0
      13'h13A8: dout <= 8'b00000000; // 5032 :   0 - 0x0
      13'h13A9: dout <= 8'b00000000; // 5033 :   0 - 0x0
      13'h13AA: dout <= 8'b00000000; // 5034 :   0 - 0x0
      13'h13AB: dout <= 8'b01110001; // 5035 : 113 - 0x71
      13'h13AC: dout <= 8'b00001010; // 5036 :  10 - 0xa
      13'h13AD: dout <= 8'b00010010; // 5037 :  18 - 0x12
      13'h13AE: dout <= 8'b00010010; // 5038 :  18 - 0x12
      13'h13AF: dout <= 8'b00100010; // 5039 :  34 - 0x22
      13'h13B0: dout <= 8'b00000000; // 5040 :   0 - 0x0 -- Background 0x3b
      13'h13B1: dout <= 8'b00000000; // 5041 :   0 - 0x0
      13'h13B2: dout <= 8'b00000000; // 5042 :   0 - 0x0
      13'h13B3: dout <= 8'b00000000; // 5043 :   0 - 0x0
      13'h13B4: dout <= 8'b00000000; // 5044 :   0 - 0x0
      13'h13B5: dout <= 8'b00000000; // 5045 :   0 - 0x0
      13'h13B6: dout <= 8'b00000000; // 5046 :   0 - 0x0
      13'h13B7: dout <= 8'b00000000; // 5047 :   0 - 0x0
      13'h13B8: dout <= 8'b00100010; // 5048 :  34 - 0x22
      13'h13B9: dout <= 8'b00100001; // 5049 :  33 - 0x21
      13'h13BA: dout <= 8'b00000000; // 5050 :   0 - 0x0
      13'h13BB: dout <= 8'b00000000; // 5051 :   0 - 0x0
      13'h13BC: dout <= 8'b00000000; // 5052 :   0 - 0x0
      13'h13BD: dout <= 8'b00000000; // 5053 :   0 - 0x0
      13'h13BE: dout <= 8'b00000000; // 5054 :   0 - 0x0
      13'h13BF: dout <= 8'b00000000; // 5055 :   0 - 0x0
      13'h13C0: dout <= 8'b00000000; // 5056 :   0 - 0x0 -- Background 0x3c
      13'h13C1: dout <= 8'b00000000; // 5057 :   0 - 0x0
      13'h13C2: dout <= 8'b00000000; // 5058 :   0 - 0x0
      13'h13C3: dout <= 8'b00000000; // 5059 :   0 - 0x0
      13'h13C4: dout <= 8'b00000000; // 5060 :   0 - 0x0
      13'h13C5: dout <= 8'b00000000; // 5061 :   0 - 0x0
      13'h13C6: dout <= 8'b00000000; // 5062 :   0 - 0x0
      13'h13C7: dout <= 8'b00000000; // 5063 :   0 - 0x0
      13'h13C8: dout <= 8'b00000000; // 5064 :   0 - 0x0
      13'h13C9: dout <= 8'b00000000; // 5065 :   0 - 0x0
      13'h13CA: dout <= 8'b00000000; // 5066 :   0 - 0x0
      13'h13CB: dout <= 8'b01110001; // 5067 : 113 - 0x71
      13'h13CC: dout <= 8'b10001010; // 5068 : 138 - 0x8a
      13'h13CD: dout <= 8'b10001010; // 5069 : 138 - 0x8a
      13'h13CE: dout <= 8'b01110010; // 5070 : 114 - 0x72
      13'h13CF: dout <= 8'b10001010; // 5071 : 138 - 0x8a
      13'h13D0: dout <= 8'b00000000; // 5072 :   0 - 0x0 -- Background 0x3d
      13'h13D1: dout <= 8'b00000000; // 5073 :   0 - 0x0
      13'h13D2: dout <= 8'b00000000; // 5074 :   0 - 0x0
      13'h13D3: dout <= 8'b00000000; // 5075 :   0 - 0x0
      13'h13D4: dout <= 8'b00000000; // 5076 :   0 - 0x0
      13'h13D5: dout <= 8'b00000000; // 5077 :   0 - 0x0
      13'h13D6: dout <= 8'b00000000; // 5078 :   0 - 0x0
      13'h13D7: dout <= 8'b00000000; // 5079 :   0 - 0x0
      13'h13D8: dout <= 8'b10001010; // 5080 : 138 - 0x8a
      13'h13D9: dout <= 8'b01110001; // 5081 : 113 - 0x71
      13'h13DA: dout <= 8'b00000000; // 5082 :   0 - 0x0
      13'h13DB: dout <= 8'b00000000; // 5083 :   0 - 0x0
      13'h13DC: dout <= 8'b00000000; // 5084 :   0 - 0x0
      13'h13DD: dout <= 8'b00000000; // 5085 :   0 - 0x0
      13'h13DE: dout <= 8'b00000000; // 5086 :   0 - 0x0
      13'h13DF: dout <= 8'b00000000; // 5087 :   0 - 0x0
      13'h13E0: dout <= 8'b00000000; // 5088 :   0 - 0x0 -- Background 0x3e
      13'h13E1: dout <= 8'b00000000; // 5089 :   0 - 0x0
      13'h13E2: dout <= 8'b00000000; // 5090 :   0 - 0x0
      13'h13E3: dout <= 8'b00000000; // 5091 :   0 - 0x0
      13'h13E4: dout <= 8'b00000000; // 5092 :   0 - 0x0
      13'h13E5: dout <= 8'b00000000; // 5093 :   0 - 0x0
      13'h13E6: dout <= 8'b00000000; // 5094 :   0 - 0x0
      13'h13E7: dout <= 8'b00000000; // 5095 :   0 - 0x0
      13'h13E8: dout <= 8'b00000000; // 5096 :   0 - 0x0
      13'h13E9: dout <= 8'b00000000; // 5097 :   0 - 0x0
      13'h13EA: dout <= 8'b00000000; // 5098 :   0 - 0x0
      13'h13EB: dout <= 8'b10011000; // 5099 : 152 - 0x98
      13'h13EC: dout <= 8'b10100101; // 5100 : 165 - 0xa5
      13'h13ED: dout <= 8'b10100101; // 5101 : 165 - 0xa5
      13'h13EE: dout <= 8'b10100101; // 5102 : 165 - 0xa5
      13'h13EF: dout <= 8'b10100101; // 5103 : 165 - 0xa5
      13'h13F0: dout <= 8'b00000000; // 5104 :   0 - 0x0 -- Background 0x3f
      13'h13F1: dout <= 8'b00000000; // 5105 :   0 - 0x0
      13'h13F2: dout <= 8'b00000000; // 5106 :   0 - 0x0
      13'h13F3: dout <= 8'b00000000; // 5107 :   0 - 0x0
      13'h13F4: dout <= 8'b00000000; // 5108 :   0 - 0x0
      13'h13F5: dout <= 8'b00000000; // 5109 :   0 - 0x0
      13'h13F6: dout <= 8'b00000000; // 5110 :   0 - 0x0
      13'h13F7: dout <= 8'b00000000; // 5111 :   0 - 0x0
      13'h13F8: dout <= 8'b00000000; // 5112 :   0 - 0x0
      13'h13F9: dout <= 8'b00000000; // 5113 :   0 - 0x0
      13'h13FA: dout <= 8'b00000000; // 5114 :   0 - 0x0
      13'h13FB: dout <= 8'b11000110; // 5115 : 198 - 0xc6
      13'h13FC: dout <= 8'b00101001; // 5116 :  41 - 0x29
      13'h13FD: dout <= 8'b00101001; // 5117 :  41 - 0x29
      13'h13FE: dout <= 8'b00101001; // 5118 :  41 - 0x29
      13'h13FF: dout <= 8'b00101001; // 5119 :  41 - 0x29
      13'h1400: dout <= 8'b00000000; // 5120 :   0 - 0x0 -- Background 0x40
      13'h1401: dout <= 8'b00000000; // 5121 :   0 - 0x0
      13'h1402: dout <= 8'b00000000; // 5122 :   0 - 0x0
      13'h1403: dout <= 8'b00000000; // 5123 :   0 - 0x0
      13'h1404: dout <= 8'b00000000; // 5124 :   0 - 0x0
      13'h1405: dout <= 8'b00000000; // 5125 :   0 - 0x0
      13'h1406: dout <= 8'b00000000; // 5126 :   0 - 0x0
      13'h1407: dout <= 8'b00000000; // 5127 :   0 - 0x0
      13'h1408: dout <= 8'b10100101; // 5128 : 165 - 0xa5
      13'h1409: dout <= 8'b10011000; // 5129 : 152 - 0x98
      13'h140A: dout <= 8'b00000000; // 5130 :   0 - 0x0
      13'h140B: dout <= 8'b00000000; // 5131 :   0 - 0x0
      13'h140C: dout <= 8'b00000000; // 5132 :   0 - 0x0
      13'h140D: dout <= 8'b00000000; // 5133 :   0 - 0x0
      13'h140E: dout <= 8'b00000000; // 5134 :   0 - 0x0
      13'h140F: dout <= 8'b00000000; // 5135 :   0 - 0x0
      13'h1410: dout <= 8'b00000000; // 5136 :   0 - 0x0 -- Background 0x41
      13'h1411: dout <= 8'b00000000; // 5137 :   0 - 0x0
      13'h1412: dout <= 8'b00000000; // 5138 :   0 - 0x0
      13'h1413: dout <= 8'b00000000; // 5139 :   0 - 0x0
      13'h1414: dout <= 8'b00000000; // 5140 :   0 - 0x0
      13'h1415: dout <= 8'b00000000; // 5141 :   0 - 0x0
      13'h1416: dout <= 8'b00000000; // 5142 :   0 - 0x0
      13'h1417: dout <= 8'b00000000; // 5143 :   0 - 0x0
      13'h1418: dout <= 8'b00101001; // 5144 :  41 - 0x29
      13'h1419: dout <= 8'b11000110; // 5145 : 198 - 0xc6
      13'h141A: dout <= 8'b00000000; // 5146 :   0 - 0x0
      13'h141B: dout <= 8'b00000000; // 5147 :   0 - 0x0
      13'h141C: dout <= 8'b00000000; // 5148 :   0 - 0x0
      13'h141D: dout <= 8'b00000000; // 5149 :   0 - 0x0
      13'h141E: dout <= 8'b00000000; // 5150 :   0 - 0x0
      13'h141F: dout <= 8'b00000000; // 5151 :   0 - 0x0
      13'h1420: dout <= 8'b00000000; // 5152 :   0 - 0x0 -- Background 0x42
      13'h1421: dout <= 8'b00000000; // 5153 :   0 - 0x0
      13'h1422: dout <= 8'b00000000; // 5154 :   0 - 0x0
      13'h1423: dout <= 8'b00000000; // 5155 :   0 - 0x0
      13'h1424: dout <= 8'b00000000; // 5156 :   0 - 0x0
      13'h1425: dout <= 8'b00000000; // 5157 :   0 - 0x0
      13'h1426: dout <= 8'b00000000; // 5158 :   0 - 0x0
      13'h1427: dout <= 8'b00000000; // 5159 :   0 - 0x0
      13'h1428: dout <= 8'b00000000; // 5160 :   0 - 0x0
      13'h1429: dout <= 8'b00000000; // 5161 :   0 - 0x0
      13'h142A: dout <= 8'b00000000; // 5162 :   0 - 0x0
      13'h142B: dout <= 8'b10011100; // 5163 : 156 - 0x9c
      13'h142C: dout <= 8'b10100001; // 5164 : 161 - 0xa1
      13'h142D: dout <= 8'b10100001; // 5165 : 161 - 0xa1
      13'h142E: dout <= 8'b10111101; // 5166 : 189 - 0xbd
      13'h142F: dout <= 8'b10100101; // 5167 : 165 - 0xa5
      13'h1430: dout <= 8'b00000000; // 5168 :   0 - 0x0 -- Background 0x43
      13'h1431: dout <= 8'b00000000; // 5169 :   0 - 0x0
      13'h1432: dout <= 8'b00000000; // 5170 :   0 - 0x0
      13'h1433: dout <= 8'b00000000; // 5171 :   0 - 0x0
      13'h1434: dout <= 8'b00000000; // 5172 :   0 - 0x0
      13'h1435: dout <= 8'b00000000; // 5173 :   0 - 0x0
      13'h1436: dout <= 8'b00000000; // 5174 :   0 - 0x0
      13'h1437: dout <= 8'b00000000; // 5175 :   0 - 0x0
      13'h1438: dout <= 8'b10100101; // 5176 : 165 - 0xa5
      13'h1439: dout <= 8'b10011000; // 5177 : 152 - 0x98
      13'h143A: dout <= 8'b00000000; // 5178 :   0 - 0x0
      13'h143B: dout <= 8'b00000000; // 5179 :   0 - 0x0
      13'h143C: dout <= 8'b00000000; // 5180 :   0 - 0x0
      13'h143D: dout <= 8'b00000000; // 5181 :   0 - 0x0
      13'h143E: dout <= 8'b00000000; // 5182 :   0 - 0x0
      13'h143F: dout <= 8'b00000000; // 5183 :   0 - 0x0
      13'h1440: dout <= 8'b00000000; // 5184 :   0 - 0x0 -- Background 0x44
      13'h1441: dout <= 8'b00000000; // 5185 :   0 - 0x0
      13'h1442: dout <= 8'b00000000; // 5186 :   0 - 0x0
      13'h1443: dout <= 8'b00000000; // 5187 :   0 - 0x0
      13'h1444: dout <= 8'b00000000; // 5188 :   0 - 0x0
      13'h1445: dout <= 8'b00000000; // 5189 :   0 - 0x0
      13'h1446: dout <= 8'b00000000; // 5190 :   0 - 0x0
      13'h1447: dout <= 8'b00000000; // 5191 :   0 - 0x0
      13'h1448: dout <= 8'b00000000; // 5192 :   0 - 0x0
      13'h1449: dout <= 8'b00000000; // 5193 :   0 - 0x0
      13'h144A: dout <= 8'b00000000; // 5194 :   0 - 0x0
      13'h144B: dout <= 8'b01100010; // 5195 :  98 - 0x62
      13'h144C: dout <= 8'b10010101; // 5196 : 149 - 0x95
      13'h144D: dout <= 8'b00010101; // 5197 :  21 - 0x15
      13'h144E: dout <= 8'b00100101; // 5198 :  37 - 0x25
      13'h144F: dout <= 8'b01000101; // 5199 :  69 - 0x45
      13'h1450: dout <= 8'b00000000; // 5200 :   0 - 0x0 -- Background 0x45
      13'h1451: dout <= 8'b00000000; // 5201 :   0 - 0x0
      13'h1452: dout <= 8'b00000000; // 5202 :   0 - 0x0
      13'h1453: dout <= 8'b00000000; // 5203 :   0 - 0x0
      13'h1454: dout <= 8'b00000000; // 5204 :   0 - 0x0
      13'h1455: dout <= 8'b00000000; // 5205 :   0 - 0x0
      13'h1456: dout <= 8'b00000000; // 5206 :   0 - 0x0
      13'h1457: dout <= 8'b00000000; // 5207 :   0 - 0x0
      13'h1458: dout <= 8'b00000000; // 5208 :   0 - 0x0
      13'h1459: dout <= 8'b00000000; // 5209 :   0 - 0x0
      13'h145A: dout <= 8'b00000000; // 5210 :   0 - 0x0
      13'h145B: dout <= 8'b00100010; // 5211 :  34 - 0x22
      13'h145C: dout <= 8'b01010101; // 5212 :  85 - 0x55
      13'h145D: dout <= 8'b01010101; // 5213 :  85 - 0x55
      13'h145E: dout <= 8'b01010101; // 5214 :  85 - 0x55
      13'h145F: dout <= 8'b01010101; // 5215 :  85 - 0x55
      13'h1460: dout <= 8'b00000000; // 5216 :   0 - 0x0 -- Background 0x46
      13'h1461: dout <= 8'b00000000; // 5217 :   0 - 0x0
      13'h1462: dout <= 8'b00000000; // 5218 :   0 - 0x0
      13'h1463: dout <= 8'b00000000; // 5219 :   0 - 0x0
      13'h1464: dout <= 8'b00000000; // 5220 :   0 - 0x0
      13'h1465: dout <= 8'b00000000; // 5221 :   0 - 0x0
      13'h1466: dout <= 8'b00000000; // 5222 :   0 - 0x0
      13'h1467: dout <= 8'b00000000; // 5223 :   0 - 0x0
      13'h1468: dout <= 8'b10000101; // 5224 : 133 - 0x85
      13'h1469: dout <= 8'b11110010; // 5225 : 242 - 0xf2
      13'h146A: dout <= 8'b00000000; // 5226 :   0 - 0x0
      13'h146B: dout <= 8'b00000000; // 5227 :   0 - 0x0
      13'h146C: dout <= 8'b00000000; // 5228 :   0 - 0x0
      13'h146D: dout <= 8'b00000000; // 5229 :   0 - 0x0
      13'h146E: dout <= 8'b00000000; // 5230 :   0 - 0x0
      13'h146F: dout <= 8'b00000000; // 5231 :   0 - 0x0
      13'h1470: dout <= 8'b00000000; // 5232 :   0 - 0x0 -- Background 0x47
      13'h1471: dout <= 8'b00000000; // 5233 :   0 - 0x0
      13'h1472: dout <= 8'b00000000; // 5234 :   0 - 0x0
      13'h1473: dout <= 8'b00000000; // 5235 :   0 - 0x0
      13'h1474: dout <= 8'b00000000; // 5236 :   0 - 0x0
      13'h1475: dout <= 8'b00000000; // 5237 :   0 - 0x0
      13'h1476: dout <= 8'b00000000; // 5238 :   0 - 0x0
      13'h1477: dout <= 8'b00000000; // 5239 :   0 - 0x0
      13'h1478: dout <= 8'b01010101; // 5240 :  85 - 0x55
      13'h1479: dout <= 8'b00100010; // 5241 :  34 - 0x22
      13'h147A: dout <= 8'b00000000; // 5242 :   0 - 0x0
      13'h147B: dout <= 8'b00000000; // 5243 :   0 - 0x0
      13'h147C: dout <= 8'b00000000; // 5244 :   0 - 0x0
      13'h147D: dout <= 8'b00000000; // 5245 :   0 - 0x0
      13'h147E: dout <= 8'b00000000; // 5246 :   0 - 0x0
      13'h147F: dout <= 8'b00000000; // 5247 :   0 - 0x0
      13'h1480: dout <= 8'b00000000; // 5248 :   0 - 0x0 -- Background 0x48
      13'h1481: dout <= 8'b00000000; // 5249 :   0 - 0x0
      13'h1482: dout <= 8'b00000000; // 5250 :   0 - 0x0
      13'h1483: dout <= 8'b00000000; // 5251 :   0 - 0x0
      13'h1484: dout <= 8'b00000000; // 5252 :   0 - 0x0
      13'h1485: dout <= 8'b00000000; // 5253 :   0 - 0x0
      13'h1486: dout <= 8'b00000000; // 5254 :   0 - 0x0
      13'h1487: dout <= 8'b00000000; // 5255 :   0 - 0x0
      13'h1488: dout <= 8'b00000000; // 5256 :   0 - 0x0
      13'h1489: dout <= 8'b00000000; // 5257 :   0 - 0x0
      13'h148A: dout <= 8'b00000000; // 5258 :   0 - 0x0
      13'h148B: dout <= 8'b01100010; // 5259 :  98 - 0x62
      13'h148C: dout <= 8'b10010101; // 5260 : 149 - 0x95
      13'h148D: dout <= 8'b00010101; // 5261 :  21 - 0x15
      13'h148E: dout <= 8'b01100101; // 5262 : 101 - 0x65
      13'h148F: dout <= 8'b00010101; // 5263 :  21 - 0x15
      13'h1490: dout <= 8'b00000000; // 5264 :   0 - 0x0 -- Background 0x49
      13'h1491: dout <= 8'b00000000; // 5265 :   0 - 0x0
      13'h1492: dout <= 8'b00000000; // 5266 :   0 - 0x0
      13'h1493: dout <= 8'b00000000; // 5267 :   0 - 0x0
      13'h1494: dout <= 8'b00000000; // 5268 :   0 - 0x0
      13'h1495: dout <= 8'b00000000; // 5269 :   0 - 0x0
      13'h1496: dout <= 8'b00000000; // 5270 :   0 - 0x0
      13'h1497: dout <= 8'b00000000; // 5271 :   0 - 0x0
      13'h1498: dout <= 8'b10010101; // 5272 : 149 - 0x95
      13'h1499: dout <= 8'b01100010; // 5273 :  98 - 0x62
      13'h149A: dout <= 8'b00000000; // 5274 :   0 - 0x0
      13'h149B: dout <= 8'b00000000; // 5275 :   0 - 0x0
      13'h149C: dout <= 8'b00000000; // 5276 :   0 - 0x0
      13'h149D: dout <= 8'b00000000; // 5277 :   0 - 0x0
      13'h149E: dout <= 8'b00000000; // 5278 :   0 - 0x0
      13'h149F: dout <= 8'b00000000; // 5279 :   0 - 0x0
      13'h14A0: dout <= 8'b00000000; // 5280 :   0 - 0x0 -- Background 0x4a
      13'h14A1: dout <= 8'b00000000; // 5281 :   0 - 0x0
      13'h14A2: dout <= 8'b00000000; // 5282 :   0 - 0x0
      13'h14A3: dout <= 8'b00000000; // 5283 :   0 - 0x0
      13'h14A4: dout <= 8'b00000000; // 5284 :   0 - 0x0
      13'h14A5: dout <= 8'b00000000; // 5285 :   0 - 0x0
      13'h14A6: dout <= 8'b00000000; // 5286 :   0 - 0x0
      13'h14A7: dout <= 8'b00000000; // 5287 :   0 - 0x0
      13'h14A8: dout <= 8'b00000000; // 5288 :   0 - 0x0
      13'h14A9: dout <= 8'b00000000; // 5289 :   0 - 0x0
      13'h14AA: dout <= 8'b00000000; // 5290 :   0 - 0x0
      13'h14AB: dout <= 8'b11100010; // 5291 : 226 - 0xe2
      13'h14AC: dout <= 8'b10000101; // 5292 : 133 - 0x85
      13'h14AD: dout <= 8'b10000101; // 5293 : 133 - 0x85
      13'h14AE: dout <= 8'b11100101; // 5294 : 229 - 0xe5
      13'h14AF: dout <= 8'b00010101; // 5295 :  21 - 0x15
      13'h14B0: dout <= 8'b00000000; // 5296 :   0 - 0x0 -- Background 0x4b
      13'h14B1: dout <= 8'b00000000; // 5297 :   0 - 0x0
      13'h14B2: dout <= 8'b00000000; // 5298 :   0 - 0x0
      13'h14B3: dout <= 8'b00000000; // 5299 :   0 - 0x0
      13'h14B4: dout <= 8'b00000000; // 5300 :   0 - 0x0
      13'h14B5: dout <= 8'b00000000; // 5301 :   0 - 0x0
      13'h14B6: dout <= 8'b00000000; // 5302 :   0 - 0x0
      13'h14B7: dout <= 8'b00000000; // 5303 :   0 - 0x0
      13'h14B8: dout <= 8'b00010101; // 5304 :  21 - 0x15
      13'h14B9: dout <= 8'b11100010; // 5305 : 226 - 0xe2
      13'h14BA: dout <= 8'b00000000; // 5306 :   0 - 0x0
      13'h14BB: dout <= 8'b00000000; // 5307 :   0 - 0x0
      13'h14BC: dout <= 8'b00000000; // 5308 :   0 - 0x0
      13'h14BD: dout <= 8'b00000000; // 5309 :   0 - 0x0
      13'h14BE: dout <= 8'b00000000; // 5310 :   0 - 0x0
      13'h14BF: dout <= 8'b00000000; // 5311 :   0 - 0x0
      13'h14C0: dout <= 8'b00000000; // 5312 :   0 - 0x0 -- Background 0x4c
      13'h14C1: dout <= 8'b00000000; // 5313 :   0 - 0x0
      13'h14C2: dout <= 8'b00000000; // 5314 :   0 - 0x0
      13'h14C3: dout <= 8'b00000000; // 5315 :   0 - 0x0
      13'h14C4: dout <= 8'b00000000; // 5316 :   0 - 0x0
      13'h14C5: dout <= 8'b00000000; // 5317 :   0 - 0x0
      13'h14C6: dout <= 8'b00000000; // 5318 :   0 - 0x0
      13'h14C7: dout <= 8'b00000000; // 5319 :   0 - 0x0
      13'h14C8: dout <= 8'b00000000; // 5320 :   0 - 0x0
      13'h14C9: dout <= 8'b00000000; // 5321 :   0 - 0x0
      13'h14CA: dout <= 8'b00000000; // 5322 :   0 - 0x0
      13'h14CB: dout <= 8'b00000000; // 5323 :   0 - 0x0
      13'h14CC: dout <= 8'b00000000; // 5324 :   0 - 0x0
      13'h14CD: dout <= 8'b00000000; // 5325 :   0 - 0x0
      13'h14CE: dout <= 8'b00000000; // 5326 :   0 - 0x0
      13'h14CF: dout <= 8'b00000000; // 5327 :   0 - 0x0
      13'h14D0: dout <= 8'b00000000; // 5328 :   0 - 0x0 -- Background 0x4d
      13'h14D1: dout <= 8'b00000000; // 5329 :   0 - 0x0
      13'h14D2: dout <= 8'b00000000; // 5330 :   0 - 0x0
      13'h14D3: dout <= 8'b00000001; // 5331 :   1 - 0x1
      13'h14D4: dout <= 8'b00000011; // 5332 :   3 - 0x3
      13'h14D5: dout <= 8'b00000111; // 5333 :   7 - 0x7
      13'h14D6: dout <= 8'b00001111; // 5334 :  15 - 0xf
      13'h14D7: dout <= 8'b00011111; // 5335 :  31 - 0x1f
      13'h14D8: dout <= 8'b00000000; // 5336 :   0 - 0x0
      13'h14D9: dout <= 8'b00000000; // 5337 :   0 - 0x0
      13'h14DA: dout <= 8'b00000000; // 5338 :   0 - 0x0
      13'h14DB: dout <= 8'b00000000; // 5339 :   0 - 0x0
      13'h14DC: dout <= 8'b00000000; // 5340 :   0 - 0x0
      13'h14DD: dout <= 8'b00000000; // 5341 :   0 - 0x0
      13'h14DE: dout <= 8'b00000000; // 5342 :   0 - 0x0
      13'h14DF: dout <= 8'b00000000; // 5343 :   0 - 0x0
      13'h14E0: dout <= 8'b00000000; // 5344 :   0 - 0x0 -- Background 0x4e
      13'h14E1: dout <= 8'b00001111; // 5345 :  15 - 0xf
      13'h14E2: dout <= 8'b01111111; // 5346 : 127 - 0x7f
      13'h14E3: dout <= 8'b11111111; // 5347 : 255 - 0xff
      13'h14E4: dout <= 8'b11111111; // 5348 : 255 - 0xff
      13'h14E5: dout <= 8'b11111111; // 5349 : 255 - 0xff
      13'h14E6: dout <= 8'b11111111; // 5350 : 255 - 0xff
      13'h14E7: dout <= 8'b11111111; // 5351 : 255 - 0xff
      13'h14E8: dout <= 8'b00000000; // 5352 :   0 - 0x0
      13'h14E9: dout <= 8'b00000000; // 5353 :   0 - 0x0
      13'h14EA: dout <= 8'b00000000; // 5354 :   0 - 0x0
      13'h14EB: dout <= 8'b00000000; // 5355 :   0 - 0x0
      13'h14EC: dout <= 8'b00000000; // 5356 :   0 - 0x0
      13'h14ED: dout <= 8'b00000000; // 5357 :   0 - 0x0
      13'h14EE: dout <= 8'b00000000; // 5358 :   0 - 0x0
      13'h14EF: dout <= 8'b00000000; // 5359 :   0 - 0x0
      13'h14F0: dout <= 8'b00011111; // 5360 :  31 - 0x1f -- Background 0x4f
      13'h14F1: dout <= 8'b00111111; // 5361 :  63 - 0x3f
      13'h14F2: dout <= 8'b00111111; // 5362 :  63 - 0x3f
      13'h14F3: dout <= 8'b00111111; // 5363 :  63 - 0x3f
      13'h14F4: dout <= 8'b01111111; // 5364 : 127 - 0x7f
      13'h14F5: dout <= 8'b01111111; // 5365 : 127 - 0x7f
      13'h14F6: dout <= 8'b01111111; // 5366 : 127 - 0x7f
      13'h14F7: dout <= 8'b01111111; // 5367 : 127 - 0x7f
      13'h14F8: dout <= 8'b00000000; // 5368 :   0 - 0x0
      13'h14F9: dout <= 8'b00000000; // 5369 :   0 - 0x0
      13'h14FA: dout <= 8'b00000000; // 5370 :   0 - 0x0
      13'h14FB: dout <= 8'b00000000; // 5371 :   0 - 0x0
      13'h14FC: dout <= 8'b00000000; // 5372 :   0 - 0x0
      13'h14FD: dout <= 8'b00000000; // 5373 :   0 - 0x0
      13'h14FE: dout <= 8'b00000000; // 5374 :   0 - 0x0
      13'h14FF: dout <= 8'b00000000; // 5375 :   0 - 0x0
      13'h1500: dout <= 8'b11111111; // 5376 : 255 - 0xff -- Background 0x50
      13'h1501: dout <= 8'b11111111; // 5377 : 255 - 0xff
      13'h1502: dout <= 8'b11111111; // 5378 : 255 - 0xff
      13'h1503: dout <= 8'b11111111; // 5379 : 255 - 0xff
      13'h1504: dout <= 8'b11111111; // 5380 : 255 - 0xff
      13'h1505: dout <= 8'b11111111; // 5381 : 255 - 0xff
      13'h1506: dout <= 8'b11111111; // 5382 : 255 - 0xff
      13'h1507: dout <= 8'b11111111; // 5383 : 255 - 0xff
      13'h1508: dout <= 8'b00000000; // 5384 :   0 - 0x0
      13'h1509: dout <= 8'b00000000; // 5385 :   0 - 0x0
      13'h150A: dout <= 8'b00000000; // 5386 :   0 - 0x0
      13'h150B: dout <= 8'b00000000; // 5387 :   0 - 0x0
      13'h150C: dout <= 8'b00000000; // 5388 :   0 - 0x0
      13'h150D: dout <= 8'b00000000; // 5389 :   0 - 0x0
      13'h150E: dout <= 8'b00000000; // 5390 :   0 - 0x0
      13'h150F: dout <= 8'b00000000; // 5391 :   0 - 0x0
      13'h1510: dout <= 8'b11111111; // 5392 : 255 - 0xff -- Background 0x51
      13'h1511: dout <= 8'b11111111; // 5393 : 255 - 0xff
      13'h1512: dout <= 8'b11111111; // 5394 : 255 - 0xff
      13'h1513: dout <= 8'b11111111; // 5395 : 255 - 0xff
      13'h1514: dout <= 8'b11111111; // 5396 : 255 - 0xff
      13'h1515: dout <= 8'b11111111; // 5397 : 255 - 0xff
      13'h1516: dout <= 8'b11111111; // 5398 : 255 - 0xff
      13'h1517: dout <= 8'b11111110; // 5399 : 254 - 0xfe
      13'h1518: dout <= 8'b00000000; // 5400 :   0 - 0x0
      13'h1519: dout <= 8'b00000000; // 5401 :   0 - 0x0
      13'h151A: dout <= 8'b00000000; // 5402 :   0 - 0x0
      13'h151B: dout <= 8'b00000000; // 5403 :   0 - 0x0
      13'h151C: dout <= 8'b00000000; // 5404 :   0 - 0x0
      13'h151D: dout <= 8'b00000000; // 5405 :   0 - 0x0
      13'h151E: dout <= 8'b00000000; // 5406 :   0 - 0x0
      13'h151F: dout <= 8'b00000000; // 5407 :   0 - 0x0
      13'h1520: dout <= 8'b00000000; // 5408 :   0 - 0x0 -- Background 0x52
      13'h1521: dout <= 8'b00000000; // 5409 :   0 - 0x0
      13'h1522: dout <= 8'b00000000; // 5410 :   0 - 0x0
      13'h1523: dout <= 8'b10000000; // 5411 : 128 - 0x80
      13'h1524: dout <= 8'b11000000; // 5412 : 192 - 0xc0
      13'h1525: dout <= 8'b11100000; // 5413 : 224 - 0xe0
      13'h1526: dout <= 8'b11110000; // 5414 : 240 - 0xf0
      13'h1527: dout <= 8'b11110000; // 5415 : 240 - 0xf0
      13'h1528: dout <= 8'b00000000; // 5416 :   0 - 0x0
      13'h1529: dout <= 8'b00000000; // 5417 :   0 - 0x0
      13'h152A: dout <= 8'b00000000; // 5418 :   0 - 0x0
      13'h152B: dout <= 8'b00000000; // 5419 :   0 - 0x0
      13'h152C: dout <= 8'b00000000; // 5420 :   0 - 0x0
      13'h152D: dout <= 8'b00000000; // 5421 :   0 - 0x0
      13'h152E: dout <= 8'b00000000; // 5422 :   0 - 0x0
      13'h152F: dout <= 8'b00000000; // 5423 :   0 - 0x0
      13'h1530: dout <= 8'b11111111; // 5424 : 255 - 0xff -- Background 0x53
      13'h1531: dout <= 8'b11111111; // 5425 : 255 - 0xff
      13'h1532: dout <= 8'b11111110; // 5426 : 254 - 0xfe
      13'h1533: dout <= 8'b11111100; // 5427 : 252 - 0xfc
      13'h1534: dout <= 8'b11110000; // 5428 : 240 - 0xf0
      13'h1535: dout <= 8'b11100000; // 5429 : 224 - 0xe0
      13'h1536: dout <= 8'b10000000; // 5430 : 128 - 0x80
      13'h1537: dout <= 8'b00000000; // 5431 :   0 - 0x0
      13'h1538: dout <= 8'b00000000; // 5432 :   0 - 0x0
      13'h1539: dout <= 8'b00000000; // 5433 :   0 - 0x0
      13'h153A: dout <= 8'b00000000; // 5434 :   0 - 0x0
      13'h153B: dout <= 8'b00000000; // 5435 :   0 - 0x0
      13'h153C: dout <= 8'b00000000; // 5436 :   0 - 0x0
      13'h153D: dout <= 8'b00000000; // 5437 :   0 - 0x0
      13'h153E: dout <= 8'b00000000; // 5438 :   0 - 0x0
      13'h153F: dout <= 8'b00000000; // 5439 :   0 - 0x0
      13'h1540: dout <= 8'b11000000; // 5440 : 192 - 0xc0 -- Background 0x54
      13'h1541: dout <= 8'b10000000; // 5441 : 128 - 0x80
      13'h1542: dout <= 8'b00000000; // 5442 :   0 - 0x0
      13'h1543: dout <= 8'b00000000; // 5443 :   0 - 0x0
      13'h1544: dout <= 8'b00000000; // 5444 :   0 - 0x0
      13'h1545: dout <= 8'b00000000; // 5445 :   0 - 0x0
      13'h1546: dout <= 8'b00000000; // 5446 :   0 - 0x0
      13'h1547: dout <= 8'b00000000; // 5447 :   0 - 0x0
      13'h1548: dout <= 8'b00000000; // 5448 :   0 - 0x0
      13'h1549: dout <= 8'b00000000; // 5449 :   0 - 0x0
      13'h154A: dout <= 8'b00000000; // 5450 :   0 - 0x0
      13'h154B: dout <= 8'b00000000; // 5451 :   0 - 0x0
      13'h154C: dout <= 8'b00000000; // 5452 :   0 - 0x0
      13'h154D: dout <= 8'b00000000; // 5453 :   0 - 0x0
      13'h154E: dout <= 8'b00000000; // 5454 :   0 - 0x0
      13'h154F: dout <= 8'b00000000; // 5455 :   0 - 0x0
      13'h1550: dout <= 8'b00000000; // 5456 :   0 - 0x0 -- Background 0x55
      13'h1551: dout <= 8'b11110000; // 5457 : 240 - 0xf0
      13'h1552: dout <= 8'b11111110; // 5458 : 254 - 0xfe
      13'h1553: dout <= 8'b11111110; // 5459 : 254 - 0xfe
      13'h1554: dout <= 8'b11111110; // 5460 : 254 - 0xfe
      13'h1555: dout <= 8'b11111100; // 5461 : 252 - 0xfc
      13'h1556: dout <= 8'b11111000; // 5462 : 248 - 0xf8
      13'h1557: dout <= 8'b11111000; // 5463 : 248 - 0xf8
      13'h1558: dout <= 8'b00000000; // 5464 :   0 - 0x0
      13'h1559: dout <= 8'b00000000; // 5465 :   0 - 0x0
      13'h155A: dout <= 8'b00000000; // 5466 :   0 - 0x0
      13'h155B: dout <= 8'b00000000; // 5467 :   0 - 0x0
      13'h155C: dout <= 8'b00000000; // 5468 :   0 - 0x0
      13'h155D: dout <= 8'b00000000; // 5469 :   0 - 0x0
      13'h155E: dout <= 8'b00000000; // 5470 :   0 - 0x0
      13'h155F: dout <= 8'b00000000; // 5471 :   0 - 0x0
      13'h1560: dout <= 8'b11110000; // 5472 : 240 - 0xf0 -- Background 0x56
      13'h1561: dout <= 8'b11100000; // 5473 : 224 - 0xe0
      13'h1562: dout <= 8'b11100000; // 5474 : 224 - 0xe0
      13'h1563: dout <= 8'b11000000; // 5475 : 192 - 0xc0
      13'h1564: dout <= 8'b10000000; // 5476 : 128 - 0x80
      13'h1565: dout <= 8'b10000000; // 5477 : 128 - 0x80
      13'h1566: dout <= 8'b00000000; // 5478 :   0 - 0x0
      13'h1567: dout <= 8'b00000000; // 5479 :   0 - 0x0
      13'h1568: dout <= 8'b00000000; // 5480 :   0 - 0x0
      13'h1569: dout <= 8'b00000000; // 5481 :   0 - 0x0
      13'h156A: dout <= 8'b00000000; // 5482 :   0 - 0x0
      13'h156B: dout <= 8'b00000000; // 5483 :   0 - 0x0
      13'h156C: dout <= 8'b00000000; // 5484 :   0 - 0x0
      13'h156D: dout <= 8'b00000000; // 5485 :   0 - 0x0
      13'h156E: dout <= 8'b00000000; // 5486 :   0 - 0x0
      13'h156F: dout <= 8'b00000000; // 5487 :   0 - 0x0
      13'h1570: dout <= 8'b00000000; // 5488 :   0 - 0x0 -- Background 0x57
      13'h1571: dout <= 8'b00000000; // 5489 :   0 - 0x0
      13'h1572: dout <= 8'b00000000; // 5490 :   0 - 0x0
      13'h1573: dout <= 8'b00000000; // 5491 :   0 - 0x0
      13'h1574: dout <= 8'b00000000; // 5492 :   0 - 0x0
      13'h1575: dout <= 8'b00000000; // 5493 :   0 - 0x0
      13'h1576: dout <= 8'b00000000; // 5494 :   0 - 0x0
      13'h1577: dout <= 8'b00000100; // 5495 :   4 - 0x4
      13'h1578: dout <= 8'b00000000; // 5496 :   0 - 0x0
      13'h1579: dout <= 8'b00000000; // 5497 :   0 - 0x0
      13'h157A: dout <= 8'b00000000; // 5498 :   0 - 0x0
      13'h157B: dout <= 8'b00000000; // 5499 :   0 - 0x0
      13'h157C: dout <= 8'b00000000; // 5500 :   0 - 0x0
      13'h157D: dout <= 8'b00000000; // 5501 :   0 - 0x0
      13'h157E: dout <= 8'b00000000; // 5502 :   0 - 0x0
      13'h157F: dout <= 8'b00000100; // 5503 :   4 - 0x4
      13'h1580: dout <= 8'b00000110; // 5504 :   6 - 0x6 -- Background 0x58
      13'h1581: dout <= 8'b00000110; // 5505 :   6 - 0x6
      13'h1582: dout <= 8'b00000111; // 5506 :   7 - 0x7
      13'h1583: dout <= 8'b00000111; // 5507 :   7 - 0x7
      13'h1584: dout <= 8'b00000111; // 5508 :   7 - 0x7
      13'h1585: dout <= 8'b00000111; // 5509 :   7 - 0x7
      13'h1586: dout <= 8'b00000000; // 5510 :   0 - 0x0
      13'h1587: dout <= 8'b00000000; // 5511 :   0 - 0x0
      13'h1588: dout <= 8'b00000110; // 5512 :   6 - 0x6
      13'h1589: dout <= 8'b00000110; // 5513 :   6 - 0x6
      13'h158A: dout <= 8'b00000111; // 5514 :   7 - 0x7
      13'h158B: dout <= 8'b00000111; // 5515 :   7 - 0x7
      13'h158C: dout <= 8'b00000111; // 5516 :   7 - 0x7
      13'h158D: dout <= 8'b00000111; // 5517 :   7 - 0x7
      13'h158E: dout <= 8'b00000000; // 5518 :   0 - 0x0
      13'h158F: dout <= 8'b00000000; // 5519 :   0 - 0x0
      13'h1590: dout <= 8'b00000000; // 5520 :   0 - 0x0 -- Background 0x59
      13'h1591: dout <= 8'b00000000; // 5521 :   0 - 0x0
      13'h1592: dout <= 8'b00000000; // 5522 :   0 - 0x0
      13'h1593: dout <= 8'b00000000; // 5523 :   0 - 0x0
      13'h1594: dout <= 8'b00000000; // 5524 :   0 - 0x0
      13'h1595: dout <= 8'b00000000; // 5525 :   0 - 0x0
      13'h1596: dout <= 8'b00000000; // 5526 :   0 - 0x0
      13'h1597: dout <= 8'b00010000; // 5527 :  16 - 0x10
      13'h1598: dout <= 8'b00000000; // 5528 :   0 - 0x0
      13'h1599: dout <= 8'b00000000; // 5529 :   0 - 0x0
      13'h159A: dout <= 8'b00000000; // 5530 :   0 - 0x0
      13'h159B: dout <= 8'b00000000; // 5531 :   0 - 0x0
      13'h159C: dout <= 8'b00000000; // 5532 :   0 - 0x0
      13'h159D: dout <= 8'b00000000; // 5533 :   0 - 0x0
      13'h159E: dout <= 8'b00000000; // 5534 :   0 - 0x0
      13'h159F: dout <= 8'b00010000; // 5535 :  16 - 0x10
      13'h15A0: dout <= 8'b00011100; // 5536 :  28 - 0x1c -- Background 0x5a
      13'h15A1: dout <= 8'b00011110; // 5537 :  30 - 0x1e
      13'h15A2: dout <= 8'b00011111; // 5538 :  31 - 0x1f
      13'h15A3: dout <= 8'b00011111; // 5539 :  31 - 0x1f
      13'h15A4: dout <= 8'b00011111; // 5540 :  31 - 0x1f
      13'h15A5: dout <= 8'b00011111; // 5541 :  31 - 0x1f
      13'h15A6: dout <= 8'b00000000; // 5542 :   0 - 0x0
      13'h15A7: dout <= 8'b00000000; // 5543 :   0 - 0x0
      13'h15A8: dout <= 8'b00011100; // 5544 :  28 - 0x1c
      13'h15A9: dout <= 8'b00011110; // 5545 :  30 - 0x1e
      13'h15AA: dout <= 8'b00011111; // 5546 :  31 - 0x1f
      13'h15AB: dout <= 8'b00011111; // 5547 :  31 - 0x1f
      13'h15AC: dout <= 8'b00011111; // 5548 :  31 - 0x1f
      13'h15AD: dout <= 8'b00011111; // 5549 :  31 - 0x1f
      13'h15AE: dout <= 8'b00000000; // 5550 :   0 - 0x0
      13'h15AF: dout <= 8'b00000000; // 5551 :   0 - 0x0
      13'h15B0: dout <= 8'b00000000; // 5552 :   0 - 0x0 -- Background 0x5b
      13'h15B1: dout <= 8'b00000000; // 5553 :   0 - 0x0
      13'h15B2: dout <= 8'b00000000; // 5554 :   0 - 0x0
      13'h15B3: dout <= 8'b00000000; // 5555 :   0 - 0x0
      13'h15B4: dout <= 8'b00000000; // 5556 :   0 - 0x0
      13'h15B5: dout <= 8'b00000000; // 5557 :   0 - 0x0
      13'h15B6: dout <= 8'b00000000; // 5558 :   0 - 0x0
      13'h15B7: dout <= 8'b11000000; // 5559 : 192 - 0xc0
      13'h15B8: dout <= 8'b00000000; // 5560 :   0 - 0x0
      13'h15B9: dout <= 8'b00000000; // 5561 :   0 - 0x0
      13'h15BA: dout <= 8'b00000000; // 5562 :   0 - 0x0
      13'h15BB: dout <= 8'b00000000; // 5563 :   0 - 0x0
      13'h15BC: dout <= 8'b00000000; // 5564 :   0 - 0x0
      13'h15BD: dout <= 8'b00000000; // 5565 :   0 - 0x0
      13'h15BE: dout <= 8'b00000000; // 5566 :   0 - 0x0
      13'h15BF: dout <= 8'b11000000; // 5567 : 192 - 0xc0
      13'h15C0: dout <= 8'b11110000; // 5568 : 240 - 0xf0 -- Background 0x5c
      13'h15C1: dout <= 8'b11111100; // 5569 : 252 - 0xfc
      13'h15C2: dout <= 8'b11111111; // 5570 : 255 - 0xff
      13'h15C3: dout <= 8'b11111111; // 5571 : 255 - 0xff
      13'h15C4: dout <= 8'b11111111; // 5572 : 255 - 0xff
      13'h15C5: dout <= 8'b11111111; // 5573 : 255 - 0xff
      13'h15C6: dout <= 8'b00000000; // 5574 :   0 - 0x0
      13'h15C7: dout <= 8'b00000000; // 5575 :   0 - 0x0
      13'h15C8: dout <= 8'b11110000; // 5576 : 240 - 0xf0
      13'h15C9: dout <= 8'b11111100; // 5577 : 252 - 0xfc
      13'h15CA: dout <= 8'b11111111; // 5578 : 255 - 0xff
      13'h15CB: dout <= 8'b11111111; // 5579 : 255 - 0xff
      13'h15CC: dout <= 8'b11111111; // 5580 : 255 - 0xff
      13'h15CD: dout <= 8'b11111111; // 5581 : 255 - 0xff
      13'h15CE: dout <= 8'b00000000; // 5582 :   0 - 0x0
      13'h15CF: dout <= 8'b00000000; // 5583 :   0 - 0x0
      13'h15D0: dout <= 8'b00000000; // 5584 :   0 - 0x0 -- Background 0x5d
      13'h15D1: dout <= 8'b00000000; // 5585 :   0 - 0x0
      13'h15D2: dout <= 8'b00000001; // 5586 :   1 - 0x1
      13'h15D3: dout <= 8'b00000011; // 5587 :   3 - 0x3
      13'h15D4: dout <= 8'b00001111; // 5588 :  15 - 0xf
      13'h15D5: dout <= 8'b00001111; // 5589 :  15 - 0xf
      13'h15D6: dout <= 8'b00000000; // 5590 :   0 - 0x0
      13'h15D7: dout <= 8'b00000000; // 5591 :   0 - 0x0
      13'h15D8: dout <= 8'b00000000; // 5592 :   0 - 0x0
      13'h15D9: dout <= 8'b00000000; // 5593 :   0 - 0x0
      13'h15DA: dout <= 8'b00000001; // 5594 :   1 - 0x1
      13'h15DB: dout <= 8'b00000011; // 5595 :   3 - 0x3
      13'h15DC: dout <= 8'b00001111; // 5596 :  15 - 0xf
      13'h15DD: dout <= 8'b00001111; // 5597 :  15 - 0xf
      13'h15DE: dout <= 8'b00000000; // 5598 :   0 - 0x0
      13'h15DF: dout <= 8'b00000000; // 5599 :   0 - 0x0
      13'h15E0: dout <= 8'b11111100; // 5600 : 252 - 0xfc -- Background 0x5e
      13'h15E1: dout <= 8'b11111100; // 5601 : 252 - 0xfc
      13'h15E2: dout <= 8'b11111100; // 5602 : 252 - 0xfc
      13'h15E3: dout <= 8'b11111100; // 5603 : 252 - 0xfc
      13'h15E4: dout <= 8'b11111000; // 5604 : 248 - 0xf8
      13'h15E5: dout <= 8'b11111100; // 5605 : 252 - 0xfc
      13'h15E6: dout <= 8'b00111100; // 5606 :  60 - 0x3c
      13'h15E7: dout <= 8'b00000000; // 5607 :   0 - 0x0
      13'h15E8: dout <= 8'b11111000; // 5608 : 248 - 0xf8
      13'h15E9: dout <= 8'b11110000; // 5609 : 240 - 0xf0
      13'h15EA: dout <= 8'b11100000; // 5610 : 224 - 0xe0
      13'h15EB: dout <= 8'b11110000; // 5611 : 240 - 0xf0
      13'h15EC: dout <= 8'b11100000; // 5612 : 224 - 0xe0
      13'h15ED: dout <= 8'b11000000; // 5613 : 192 - 0xc0
      13'h15EE: dout <= 8'b00000000; // 5614 :   0 - 0x0
      13'h15EF: dout <= 8'b00000000; // 5615 :   0 - 0x0
      13'h15F0: dout <= 8'b00000100; // 5616 :   4 - 0x4 -- Background 0x5f
      13'h15F1: dout <= 8'b00001100; // 5617 :  12 - 0xc
      13'h15F2: dout <= 8'b00011100; // 5618 :  28 - 0x1c
      13'h15F3: dout <= 8'b00001100; // 5619 :  12 - 0xc
      13'h15F4: dout <= 8'b00011000; // 5620 :  24 - 0x18
      13'h15F5: dout <= 8'b00111100; // 5621 :  60 - 0x3c
      13'h15F6: dout <= 8'b00111100; // 5622 :  60 - 0x3c
      13'h15F7: dout <= 8'b00000000; // 5623 :   0 - 0x0
      13'h15F8: dout <= 8'b00000000; // 5624 :   0 - 0x0
      13'h15F9: dout <= 8'b00000000; // 5625 :   0 - 0x0
      13'h15FA: dout <= 8'b00000000; // 5626 :   0 - 0x0
      13'h15FB: dout <= 8'b00000000; // 5627 :   0 - 0x0
      13'h15FC: dout <= 8'b00000000; // 5628 :   0 - 0x0
      13'h15FD: dout <= 8'b00000000; // 5629 :   0 - 0x0
      13'h15FE: dout <= 8'b00000000; // 5630 :   0 - 0x0
      13'h15FF: dout <= 8'b00000000; // 5631 :   0 - 0x0
      13'h1600: dout <= 8'b00000000; // 5632 :   0 - 0x0 -- Background 0x60
      13'h1601: dout <= 8'b00000011; // 5633 :   3 - 0x3
      13'h1602: dout <= 8'b00001111; // 5634 :  15 - 0xf
      13'h1603: dout <= 8'b00010011; // 5635 :  19 - 0x13
      13'h1604: dout <= 8'b00100001; // 5636 :  33 - 0x21
      13'h1605: dout <= 8'b00100001; // 5637 :  33 - 0x21
      13'h1606: dout <= 8'b00100001; // 5638 :  33 - 0x21
      13'h1607: dout <= 8'b01110011; // 5639 : 115 - 0x73
      13'h1608: dout <= 8'b00000000; // 5640 :   0 - 0x0
      13'h1609: dout <= 8'b00000011; // 5641 :   3 - 0x3
      13'h160A: dout <= 8'b00001111; // 5642 :  15 - 0xf
      13'h160B: dout <= 8'b00011111; // 5643 :  31 - 0x1f
      13'h160C: dout <= 8'b00111111; // 5644 :  63 - 0x3f
      13'h160D: dout <= 8'b00111111; // 5645 :  63 - 0x3f
      13'h160E: dout <= 8'b00111001; // 5646 :  57 - 0x39
      13'h160F: dout <= 8'b01111011; // 5647 : 123 - 0x7b
      13'h1610: dout <= 8'b00000000; // 5648 :   0 - 0x0 -- Background 0x61
      13'h1611: dout <= 8'b11000000; // 5649 : 192 - 0xc0
      13'h1612: dout <= 8'b11110000; // 5650 : 240 - 0xf0
      13'h1613: dout <= 8'b11001000; // 5651 : 200 - 0xc8
      13'h1614: dout <= 8'b10000100; // 5652 : 132 - 0x84
      13'h1615: dout <= 8'b10000100; // 5653 : 132 - 0x84
      13'h1616: dout <= 8'b10000100; // 5654 : 132 - 0x84
      13'h1617: dout <= 8'b11001110; // 5655 : 206 - 0xce
      13'h1618: dout <= 8'b00000000; // 5656 :   0 - 0x0
      13'h1619: dout <= 8'b11000000; // 5657 : 192 - 0xc0
      13'h161A: dout <= 8'b11110000; // 5658 : 240 - 0xf0
      13'h161B: dout <= 8'b11111000; // 5659 : 248 - 0xf8
      13'h161C: dout <= 8'b11111100; // 5660 : 252 - 0xfc
      13'h161D: dout <= 8'b11111100; // 5661 : 252 - 0xfc
      13'h161E: dout <= 8'b11100100; // 5662 : 228 - 0xe4
      13'h161F: dout <= 8'b11101110; // 5663 : 238 - 0xee
      13'h1620: dout <= 8'b10010100; // 5664 : 148 - 0x94 -- Background 0x62
      13'h1621: dout <= 8'b11101010; // 5665 : 234 - 0xea
      13'h1622: dout <= 8'b11011110; // 5666 : 222 - 0xde
      13'h1623: dout <= 8'b11101110; // 5667 : 238 - 0xee
      13'h1624: dout <= 8'b11011110; // 5668 : 222 - 0xde
      13'h1625: dout <= 8'b01100110; // 5669 : 102 - 0x66
      13'h1626: dout <= 8'b01000010; // 5670 :  66 - 0x42
      13'h1627: dout <= 8'b00000000; // 5671 :   0 - 0x0
      13'h1628: dout <= 8'b11111110; // 5672 : 254 - 0xfe
      13'h1629: dout <= 8'b11111110; // 5673 : 254 - 0xfe
      13'h162A: dout <= 8'b11111110; // 5674 : 254 - 0xfe
      13'h162B: dout <= 8'b11111110; // 5675 : 254 - 0xfe
      13'h162C: dout <= 8'b11111110; // 5676 : 254 - 0xfe
      13'h162D: dout <= 8'b01100110; // 5677 : 102 - 0x66
      13'h162E: dout <= 8'b01000010; // 5678 :  66 - 0x42
      13'h162F: dout <= 8'b00000000; // 5679 :   0 - 0x0
      13'h1630: dout <= 8'b10010100; // 5680 : 148 - 0x94 -- Background 0x63
      13'h1631: dout <= 8'b11101010; // 5681 : 234 - 0xea
      13'h1632: dout <= 8'b11011110; // 5682 : 222 - 0xde
      13'h1633: dout <= 8'b11101110; // 5683 : 238 - 0xee
      13'h1634: dout <= 8'b11011110; // 5684 : 222 - 0xde
      13'h1635: dout <= 8'b11001110; // 5685 : 206 - 0xce
      13'h1636: dout <= 8'b10001100; // 5686 : 140 - 0x8c
      13'h1637: dout <= 8'b00000000; // 5687 :   0 - 0x0
      13'h1638: dout <= 8'b11111110; // 5688 : 254 - 0xfe
      13'h1639: dout <= 8'b11111110; // 5689 : 254 - 0xfe
      13'h163A: dout <= 8'b11111110; // 5690 : 254 - 0xfe
      13'h163B: dout <= 8'b11111110; // 5691 : 254 - 0xfe
      13'h163C: dout <= 8'b11111110; // 5692 : 254 - 0xfe
      13'h163D: dout <= 8'b11011110; // 5693 : 222 - 0xde
      13'h163E: dout <= 8'b10001100; // 5694 : 140 - 0x8c
      13'h163F: dout <= 8'b00000000; // 5695 :   0 - 0x0
      13'h1640: dout <= 8'b00000000; // 5696 :   0 - 0x0 -- Background 0x64
      13'h1641: dout <= 8'b00000000; // 5697 :   0 - 0x0
      13'h1642: dout <= 8'b00000000; // 5698 :   0 - 0x0
      13'h1643: dout <= 8'b00000000; // 5699 :   0 - 0x0
      13'h1644: dout <= 8'b00000000; // 5700 :   0 - 0x0
      13'h1645: dout <= 8'b00000000; // 5701 :   0 - 0x0
      13'h1646: dout <= 8'b00000000; // 5702 :   0 - 0x0
      13'h1647: dout <= 8'b00000001; // 5703 :   1 - 0x1
      13'h1648: dout <= 8'b00000000; // 5704 :   0 - 0x0
      13'h1649: dout <= 8'b00000000; // 5705 :   0 - 0x0
      13'h164A: dout <= 8'b00000000; // 5706 :   0 - 0x0
      13'h164B: dout <= 8'b00000000; // 5707 :   0 - 0x0
      13'h164C: dout <= 8'b00000000; // 5708 :   0 - 0x0
      13'h164D: dout <= 8'b00000000; // 5709 :   0 - 0x0
      13'h164E: dout <= 8'b00000000; // 5710 :   0 - 0x0
      13'h164F: dout <= 8'b00000000; // 5711 :   0 - 0x0
      13'h1650: dout <= 8'b00000000; // 5712 :   0 - 0x0 -- Background 0x65
      13'h1651: dout <= 8'b00000000; // 5713 :   0 - 0x0
      13'h1652: dout <= 8'b00000000; // 5714 :   0 - 0x0
      13'h1653: dout <= 8'b00000000; // 5715 :   0 - 0x0
      13'h1654: dout <= 8'b00000000; // 5716 :   0 - 0x0
      13'h1655: dout <= 8'b00110110; // 5717 :  54 - 0x36
      13'h1656: dout <= 8'b00110110; // 5718 :  54 - 0x36
      13'h1657: dout <= 8'b10010000; // 5719 : 144 - 0x90
      13'h1658: dout <= 8'b00000000; // 5720 :   0 - 0x0
      13'h1659: dout <= 8'b00000000; // 5721 :   0 - 0x0
      13'h165A: dout <= 8'b00000000; // 5722 :   0 - 0x0
      13'h165B: dout <= 8'b00000000; // 5723 :   0 - 0x0
      13'h165C: dout <= 8'b01101100; // 5724 : 108 - 0x6c
      13'h165D: dout <= 8'b11111110; // 5725 : 254 - 0xfe
      13'h165E: dout <= 8'b11111110; // 5726 : 254 - 0xfe
      13'h165F: dout <= 8'b11111100; // 5727 : 252 - 0xfc
      13'h1660: dout <= 8'b00000001; // 5728 :   1 - 0x1 -- Background 0x66
      13'h1661: dout <= 8'b00000011; // 5729 :   3 - 0x3
      13'h1662: dout <= 8'b00000111; // 5730 :   7 - 0x7
      13'h1663: dout <= 8'b00000111; // 5731 :   7 - 0x7
      13'h1664: dout <= 8'b00011111; // 5732 :  31 - 0x1f
      13'h1665: dout <= 8'b00011111; // 5733 :  31 - 0x1f
      13'h1666: dout <= 8'b00011100; // 5734 :  28 - 0x1c
      13'h1667: dout <= 8'b00000000; // 5735 :   0 - 0x0
      13'h1668: dout <= 8'b00000000; // 5736 :   0 - 0x0
      13'h1669: dout <= 8'b00000000; // 5737 :   0 - 0x0
      13'h166A: dout <= 8'b00000000; // 5738 :   0 - 0x0
      13'h166B: dout <= 8'b00000000; // 5739 :   0 - 0x0
      13'h166C: dout <= 8'b00000000; // 5740 :   0 - 0x0
      13'h166D: dout <= 8'b00000000; // 5741 :   0 - 0x0
      13'h166E: dout <= 8'b00000000; // 5742 :   0 - 0x0
      13'h166F: dout <= 8'b00000000; // 5743 :   0 - 0x0
      13'h1670: dout <= 8'b11111000; // 5744 : 248 - 0xf8 -- Background 0x67
      13'h1671: dout <= 8'b11111000; // 5745 : 248 - 0xf8
      13'h1672: dout <= 8'b11111000; // 5746 : 248 - 0xf8
      13'h1673: dout <= 8'b11111000; // 5747 : 248 - 0xf8
      13'h1674: dout <= 8'b11111110; // 5748 : 254 - 0xfe
      13'h1675: dout <= 8'b11111110; // 5749 : 254 - 0xfe
      13'h1676: dout <= 8'b00001110; // 5750 :  14 - 0xe
      13'h1677: dout <= 8'b00000000; // 5751 :   0 - 0x0
      13'h1678: dout <= 8'b00000000; // 5752 :   0 - 0x0
      13'h1679: dout <= 8'b00000000; // 5753 :   0 - 0x0
      13'h167A: dout <= 8'b00000000; // 5754 :   0 - 0x0
      13'h167B: dout <= 8'b00000000; // 5755 :   0 - 0x0
      13'h167C: dout <= 8'b00000000; // 5756 :   0 - 0x0
      13'h167D: dout <= 8'b00000000; // 5757 :   0 - 0x0
      13'h167E: dout <= 8'b00000000; // 5758 :   0 - 0x0
      13'h167F: dout <= 8'b00000000; // 5759 :   0 - 0x0
      13'h1680: dout <= 8'b00000111; // 5760 :   7 - 0x7 -- Background 0x68
      13'h1681: dout <= 8'b00001111; // 5761 :  15 - 0xf
      13'h1682: dout <= 8'b00011111; // 5762 :  31 - 0x1f
      13'h1683: dout <= 8'b00011111; // 5763 :  31 - 0x1f
      13'h1684: dout <= 8'b00111111; // 5764 :  63 - 0x3f
      13'h1685: dout <= 8'b00111111; // 5765 :  63 - 0x3f
      13'h1686: dout <= 8'b00111000; // 5766 :  56 - 0x38
      13'h1687: dout <= 8'b00000000; // 5767 :   0 - 0x0
      13'h1688: dout <= 8'b00000000; // 5768 :   0 - 0x0
      13'h1689: dout <= 8'b00000000; // 5769 :   0 - 0x0
      13'h168A: dout <= 8'b00000000; // 5770 :   0 - 0x0
      13'h168B: dout <= 8'b00000000; // 5771 :   0 - 0x0
      13'h168C: dout <= 8'b00000000; // 5772 :   0 - 0x0
      13'h168D: dout <= 8'b00000000; // 5773 :   0 - 0x0
      13'h168E: dout <= 8'b00000000; // 5774 :   0 - 0x0
      13'h168F: dout <= 8'b00000000; // 5775 :   0 - 0x0
      13'h1690: dout <= 8'b11111000; // 5776 : 248 - 0xf8 -- Background 0x69
      13'h1691: dout <= 8'b11110000; // 5777 : 240 - 0xf0
      13'h1692: dout <= 8'b11110000; // 5778 : 240 - 0xf0
      13'h1693: dout <= 8'b11100000; // 5779 : 224 - 0xe0
      13'h1694: dout <= 8'b11111000; // 5780 : 248 - 0xf8
      13'h1695: dout <= 8'b11111000; // 5781 : 248 - 0xf8
      13'h1696: dout <= 8'b00111000; // 5782 :  56 - 0x38
      13'h1697: dout <= 8'b00000000; // 5783 :   0 - 0x0
      13'h1698: dout <= 8'b00000000; // 5784 :   0 - 0x0
      13'h1699: dout <= 8'b00000000; // 5785 :   0 - 0x0
      13'h169A: dout <= 8'b00000000; // 5786 :   0 - 0x0
      13'h169B: dout <= 8'b00000000; // 5787 :   0 - 0x0
      13'h169C: dout <= 8'b00000000; // 5788 :   0 - 0x0
      13'h169D: dout <= 8'b00000000; // 5789 :   0 - 0x0
      13'h169E: dout <= 8'b00000000; // 5790 :   0 - 0x0
      13'h169F: dout <= 8'b00000000; // 5791 :   0 - 0x0
      13'h16A0: dout <= 8'b00000000; // 5792 :   0 - 0x0 -- Background 0x6a
      13'h16A1: dout <= 8'b00011111; // 5793 :  31 - 0x1f
      13'h16A2: dout <= 8'b01111111; // 5794 : 127 - 0x7f
      13'h16A3: dout <= 8'b00111111; // 5795 :  63 - 0x3f
      13'h16A4: dout <= 8'b00001111; // 5796 :  15 - 0xf
      13'h16A5: dout <= 8'b00000111; // 5797 :   7 - 0x7
      13'h16A6: dout <= 8'b00000000; // 5798 :   0 - 0x0
      13'h16A7: dout <= 8'b00000000; // 5799 :   0 - 0x0
      13'h16A8: dout <= 8'b00000000; // 5800 :   0 - 0x0
      13'h16A9: dout <= 8'b00011111; // 5801 :  31 - 0x1f
      13'h16AA: dout <= 8'b01111111; // 5802 : 127 - 0x7f
      13'h16AB: dout <= 8'b00111111; // 5803 :  63 - 0x3f
      13'h16AC: dout <= 8'b00001111; // 5804 :  15 - 0xf
      13'h16AD: dout <= 8'b00000111; // 5805 :   7 - 0x7
      13'h16AE: dout <= 8'b00000000; // 5806 :   0 - 0x0
      13'h16AF: dout <= 8'b00000000; // 5807 :   0 - 0x0
      13'h16B0: dout <= 8'b00000000; // 5808 :   0 - 0x0 -- Background 0x6b
      13'h16B1: dout <= 8'b00000000; // 5809 :   0 - 0x0
      13'h16B2: dout <= 8'b11000000; // 5810 : 192 - 0xc0
      13'h16B3: dout <= 8'b11110000; // 5811 : 240 - 0xf0
      13'h16B4: dout <= 8'b11111000; // 5812 : 248 - 0xf8
      13'h16B5: dout <= 8'b11111000; // 5813 : 248 - 0xf8
      13'h16B6: dout <= 8'b11100000; // 5814 : 224 - 0xe0
      13'h16B7: dout <= 8'b00000000; // 5815 :   0 - 0x0
      13'h16B8: dout <= 8'b00000000; // 5816 :   0 - 0x0
      13'h16B9: dout <= 8'b00000000; // 5817 :   0 - 0x0
      13'h16BA: dout <= 8'b11000000; // 5818 : 192 - 0xc0
      13'h16BB: dout <= 8'b11110000; // 5819 : 240 - 0xf0
      13'h16BC: dout <= 8'b11111000; // 5820 : 248 - 0xf8
      13'h16BD: dout <= 8'b11111000; // 5821 : 248 - 0xf8
      13'h16BE: dout <= 8'b11100000; // 5822 : 224 - 0xe0
      13'h16BF: dout <= 8'b00000000; // 5823 :   0 - 0x0
      13'h16C0: dout <= 8'b00000000; // 5824 :   0 - 0x0 -- Background 0x6c
      13'h16C1: dout <= 8'b00000000; // 5825 :   0 - 0x0
      13'h16C2: dout <= 8'b00000000; // 5826 :   0 - 0x0
      13'h16C3: dout <= 8'b00000000; // 5827 :   0 - 0x0
      13'h16C4: dout <= 8'b00000000; // 5828 :   0 - 0x0
      13'h16C5: dout <= 8'b00000000; // 5829 :   0 - 0x0
      13'h16C6: dout <= 8'b00000000; // 5830 :   0 - 0x0
      13'h16C7: dout <= 8'b00000000; // 5831 :   0 - 0x0
      13'h16C8: dout <= 8'b00000000; // 5832 :   0 - 0x0
      13'h16C9: dout <= 8'b00000000; // 5833 :   0 - 0x0
      13'h16CA: dout <= 8'b00000000; // 5834 :   0 - 0x0
      13'h16CB: dout <= 8'b00000000; // 5835 :   0 - 0x0
      13'h16CC: dout <= 8'b00000000; // 5836 :   0 - 0x0
      13'h16CD: dout <= 8'b00000000; // 5837 :   0 - 0x0
      13'h16CE: dout <= 8'b00000000; // 5838 :   0 - 0x0
      13'h16CF: dout <= 8'b00000000; // 5839 :   0 - 0x0
      13'h16D0: dout <= 8'b00000000; // 5840 :   0 - 0x0 -- Background 0x6d
      13'h16D1: dout <= 8'b00000000; // 5841 :   0 - 0x0
      13'h16D2: dout <= 8'b00000000; // 5842 :   0 - 0x0
      13'h16D3: dout <= 8'b00000000; // 5843 :   0 - 0x0
      13'h16D4: dout <= 8'b00000000; // 5844 :   0 - 0x0
      13'h16D5: dout <= 8'b00000000; // 5845 :   0 - 0x0
      13'h16D6: dout <= 8'b00000000; // 5846 :   0 - 0x0
      13'h16D7: dout <= 8'b00000000; // 5847 :   0 - 0x0
      13'h16D8: dout <= 8'b00000000; // 5848 :   0 - 0x0
      13'h16D9: dout <= 8'b00000000; // 5849 :   0 - 0x0
      13'h16DA: dout <= 8'b00000000; // 5850 :   0 - 0x0
      13'h16DB: dout <= 8'b00000000; // 5851 :   0 - 0x0
      13'h16DC: dout <= 8'b00000000; // 5852 :   0 - 0x0
      13'h16DD: dout <= 8'b00000000; // 5853 :   0 - 0x0
      13'h16DE: dout <= 8'b00000000; // 5854 :   0 - 0x0
      13'h16DF: dout <= 8'b00000000; // 5855 :   0 - 0x0
      13'h16E0: dout <= 8'b00000000; // 5856 :   0 - 0x0 -- Background 0x6e
      13'h16E1: dout <= 8'b00000000; // 5857 :   0 - 0x0
      13'h16E2: dout <= 8'b00000000; // 5858 :   0 - 0x0
      13'h16E3: dout <= 8'b00000000; // 5859 :   0 - 0x0
      13'h16E4: dout <= 8'b00000000; // 5860 :   0 - 0x0
      13'h16E5: dout <= 8'b00000000; // 5861 :   0 - 0x0
      13'h16E6: dout <= 8'b00000000; // 5862 :   0 - 0x0
      13'h16E7: dout <= 8'b00000000; // 5863 :   0 - 0x0
      13'h16E8: dout <= 8'b00000000; // 5864 :   0 - 0x0
      13'h16E9: dout <= 8'b00000000; // 5865 :   0 - 0x0
      13'h16EA: dout <= 8'b00000000; // 5866 :   0 - 0x0
      13'h16EB: dout <= 8'b00000000; // 5867 :   0 - 0x0
      13'h16EC: dout <= 8'b00000000; // 5868 :   0 - 0x0
      13'h16ED: dout <= 8'b00000000; // 5869 :   0 - 0x0
      13'h16EE: dout <= 8'b00000000; // 5870 :   0 - 0x0
      13'h16EF: dout <= 8'b00000000; // 5871 :   0 - 0x0
      13'h16F0: dout <= 8'b00000000; // 5872 :   0 - 0x0 -- Background 0x6f
      13'h16F1: dout <= 8'b00000000; // 5873 :   0 - 0x0
      13'h16F2: dout <= 8'b00000000; // 5874 :   0 - 0x0
      13'h16F3: dout <= 8'b00000000; // 5875 :   0 - 0x0
      13'h16F4: dout <= 8'b00000000; // 5876 :   0 - 0x0
      13'h16F5: dout <= 8'b00000000; // 5877 :   0 - 0x0
      13'h16F6: dout <= 8'b00000000; // 5878 :   0 - 0x0
      13'h16F7: dout <= 8'b00000000; // 5879 :   0 - 0x0
      13'h16F8: dout <= 8'b00000000; // 5880 :   0 - 0x0
      13'h16F9: dout <= 8'b00000000; // 5881 :   0 - 0x0
      13'h16FA: dout <= 8'b00000000; // 5882 :   0 - 0x0
      13'h16FB: dout <= 8'b00000000; // 5883 :   0 - 0x0
      13'h16FC: dout <= 8'b00000000; // 5884 :   0 - 0x0
      13'h16FD: dout <= 8'b00000000; // 5885 :   0 - 0x0
      13'h16FE: dout <= 8'b00000000; // 5886 :   0 - 0x0
      13'h16FF: dout <= 8'b00000000; // 5887 :   0 - 0x0
      13'h1700: dout <= 8'b11111111; // 5888 : 255 - 0xff -- Background 0x70
      13'h1701: dout <= 8'b11111111; // 5889 : 255 - 0xff
      13'h1702: dout <= 8'b11111111; // 5890 : 255 - 0xff
      13'h1703: dout <= 8'b11111111; // 5891 : 255 - 0xff
      13'h1704: dout <= 8'b11111111; // 5892 : 255 - 0xff
      13'h1705: dout <= 8'b11111111; // 5893 : 255 - 0xff
      13'h1706: dout <= 8'b11111111; // 5894 : 255 - 0xff
      13'h1707: dout <= 8'b11111111; // 5895 : 255 - 0xff
      13'h1708: dout <= 8'b11111111; // 5896 : 255 - 0xff
      13'h1709: dout <= 8'b11111111; // 5897 : 255 - 0xff
      13'h170A: dout <= 8'b11111111; // 5898 : 255 - 0xff
      13'h170B: dout <= 8'b11111111; // 5899 : 255 - 0xff
      13'h170C: dout <= 8'b11111111; // 5900 : 255 - 0xff
      13'h170D: dout <= 8'b11111111; // 5901 : 255 - 0xff
      13'h170E: dout <= 8'b11111111; // 5902 : 255 - 0xff
      13'h170F: dout <= 8'b11111111; // 5903 : 255 - 0xff
      13'h1710: dout <= 8'b11111111; // 5904 : 255 - 0xff -- Background 0x71
      13'h1711: dout <= 8'b11111111; // 5905 : 255 - 0xff
      13'h1712: dout <= 8'b11111111; // 5906 : 255 - 0xff
      13'h1713: dout <= 8'b11111111; // 5907 : 255 - 0xff
      13'h1714: dout <= 8'b11111111; // 5908 : 255 - 0xff
      13'h1715: dout <= 8'b11111111; // 5909 : 255 - 0xff
      13'h1716: dout <= 8'b11111111; // 5910 : 255 - 0xff
      13'h1717: dout <= 8'b11111111; // 5911 : 255 - 0xff
      13'h1718: dout <= 8'b11111111; // 5912 : 255 - 0xff
      13'h1719: dout <= 8'b11111111; // 5913 : 255 - 0xff
      13'h171A: dout <= 8'b11111111; // 5914 : 255 - 0xff
      13'h171B: dout <= 8'b11111111; // 5915 : 255 - 0xff
      13'h171C: dout <= 8'b11111111; // 5916 : 255 - 0xff
      13'h171D: dout <= 8'b11111111; // 5917 : 255 - 0xff
      13'h171E: dout <= 8'b11111111; // 5918 : 255 - 0xff
      13'h171F: dout <= 8'b11111111; // 5919 : 255 - 0xff
      13'h1720: dout <= 8'b11111111; // 5920 : 255 - 0xff -- Background 0x72
      13'h1721: dout <= 8'b11111111; // 5921 : 255 - 0xff
      13'h1722: dout <= 8'b11111111; // 5922 : 255 - 0xff
      13'h1723: dout <= 8'b11111111; // 5923 : 255 - 0xff
      13'h1724: dout <= 8'b11111111; // 5924 : 255 - 0xff
      13'h1725: dout <= 8'b11111111; // 5925 : 255 - 0xff
      13'h1726: dout <= 8'b11111111; // 5926 : 255 - 0xff
      13'h1727: dout <= 8'b11111111; // 5927 : 255 - 0xff
      13'h1728: dout <= 8'b11111111; // 5928 : 255 - 0xff
      13'h1729: dout <= 8'b11111111; // 5929 : 255 - 0xff
      13'h172A: dout <= 8'b11111111; // 5930 : 255 - 0xff
      13'h172B: dout <= 8'b11111111; // 5931 : 255 - 0xff
      13'h172C: dout <= 8'b11111111; // 5932 : 255 - 0xff
      13'h172D: dout <= 8'b11111111; // 5933 : 255 - 0xff
      13'h172E: dout <= 8'b11111111; // 5934 : 255 - 0xff
      13'h172F: dout <= 8'b11111111; // 5935 : 255 - 0xff
      13'h1730: dout <= 8'b11111111; // 5936 : 255 - 0xff -- Background 0x73
      13'h1731: dout <= 8'b11111111; // 5937 : 255 - 0xff
      13'h1732: dout <= 8'b11111111; // 5938 : 255 - 0xff
      13'h1733: dout <= 8'b11111111; // 5939 : 255 - 0xff
      13'h1734: dout <= 8'b11111111; // 5940 : 255 - 0xff
      13'h1735: dout <= 8'b11111111; // 5941 : 255 - 0xff
      13'h1736: dout <= 8'b11111111; // 5942 : 255 - 0xff
      13'h1737: dout <= 8'b11111111; // 5943 : 255 - 0xff
      13'h1738: dout <= 8'b11111111; // 5944 : 255 - 0xff
      13'h1739: dout <= 8'b11111111; // 5945 : 255 - 0xff
      13'h173A: dout <= 8'b11111111; // 5946 : 255 - 0xff
      13'h173B: dout <= 8'b11111111; // 5947 : 255 - 0xff
      13'h173C: dout <= 8'b11111111; // 5948 : 255 - 0xff
      13'h173D: dout <= 8'b11111111; // 5949 : 255 - 0xff
      13'h173E: dout <= 8'b11111111; // 5950 : 255 - 0xff
      13'h173F: dout <= 8'b11111111; // 5951 : 255 - 0xff
      13'h1740: dout <= 8'b11111111; // 5952 : 255 - 0xff -- Background 0x74
      13'h1741: dout <= 8'b11111111; // 5953 : 255 - 0xff
      13'h1742: dout <= 8'b11111111; // 5954 : 255 - 0xff
      13'h1743: dout <= 8'b11111111; // 5955 : 255 - 0xff
      13'h1744: dout <= 8'b11111111; // 5956 : 255 - 0xff
      13'h1745: dout <= 8'b11111111; // 5957 : 255 - 0xff
      13'h1746: dout <= 8'b11111111; // 5958 : 255 - 0xff
      13'h1747: dout <= 8'b11111111; // 5959 : 255 - 0xff
      13'h1748: dout <= 8'b11111111; // 5960 : 255 - 0xff
      13'h1749: dout <= 8'b11111111; // 5961 : 255 - 0xff
      13'h174A: dout <= 8'b11111111; // 5962 : 255 - 0xff
      13'h174B: dout <= 8'b11111111; // 5963 : 255 - 0xff
      13'h174C: dout <= 8'b11111111; // 5964 : 255 - 0xff
      13'h174D: dout <= 8'b11111111; // 5965 : 255 - 0xff
      13'h174E: dout <= 8'b11111111; // 5966 : 255 - 0xff
      13'h174F: dout <= 8'b11111111; // 5967 : 255 - 0xff
      13'h1750: dout <= 8'b11111111; // 5968 : 255 - 0xff -- Background 0x75
      13'h1751: dout <= 8'b11111111; // 5969 : 255 - 0xff
      13'h1752: dout <= 8'b11111111; // 5970 : 255 - 0xff
      13'h1753: dout <= 8'b11111111; // 5971 : 255 - 0xff
      13'h1754: dout <= 8'b11111111; // 5972 : 255 - 0xff
      13'h1755: dout <= 8'b11111111; // 5973 : 255 - 0xff
      13'h1756: dout <= 8'b11111111; // 5974 : 255 - 0xff
      13'h1757: dout <= 8'b11111111; // 5975 : 255 - 0xff
      13'h1758: dout <= 8'b11111111; // 5976 : 255 - 0xff
      13'h1759: dout <= 8'b11111111; // 5977 : 255 - 0xff
      13'h175A: dout <= 8'b11111111; // 5978 : 255 - 0xff
      13'h175B: dout <= 8'b11111111; // 5979 : 255 - 0xff
      13'h175C: dout <= 8'b11111111; // 5980 : 255 - 0xff
      13'h175D: dout <= 8'b11111111; // 5981 : 255 - 0xff
      13'h175E: dout <= 8'b11111111; // 5982 : 255 - 0xff
      13'h175F: dout <= 8'b11111111; // 5983 : 255 - 0xff
      13'h1760: dout <= 8'b11111111; // 5984 : 255 - 0xff -- Background 0x76
      13'h1761: dout <= 8'b11111111; // 5985 : 255 - 0xff
      13'h1762: dout <= 8'b11111111; // 5986 : 255 - 0xff
      13'h1763: dout <= 8'b11111111; // 5987 : 255 - 0xff
      13'h1764: dout <= 8'b11111111; // 5988 : 255 - 0xff
      13'h1765: dout <= 8'b11111111; // 5989 : 255 - 0xff
      13'h1766: dout <= 8'b11111111; // 5990 : 255 - 0xff
      13'h1767: dout <= 8'b11111111; // 5991 : 255 - 0xff
      13'h1768: dout <= 8'b11111111; // 5992 : 255 - 0xff
      13'h1769: dout <= 8'b11111111; // 5993 : 255 - 0xff
      13'h176A: dout <= 8'b11111111; // 5994 : 255 - 0xff
      13'h176B: dout <= 8'b11111111; // 5995 : 255 - 0xff
      13'h176C: dout <= 8'b11111111; // 5996 : 255 - 0xff
      13'h176D: dout <= 8'b11111111; // 5997 : 255 - 0xff
      13'h176E: dout <= 8'b11111111; // 5998 : 255 - 0xff
      13'h176F: dout <= 8'b11111111; // 5999 : 255 - 0xff
      13'h1770: dout <= 8'b11111111; // 6000 : 255 - 0xff -- Background 0x77
      13'h1771: dout <= 8'b11111111; // 6001 : 255 - 0xff
      13'h1772: dout <= 8'b11111111; // 6002 : 255 - 0xff
      13'h1773: dout <= 8'b11111111; // 6003 : 255 - 0xff
      13'h1774: dout <= 8'b11111111; // 6004 : 255 - 0xff
      13'h1775: dout <= 8'b11111111; // 6005 : 255 - 0xff
      13'h1776: dout <= 8'b11111111; // 6006 : 255 - 0xff
      13'h1777: dout <= 8'b11111111; // 6007 : 255 - 0xff
      13'h1778: dout <= 8'b11111111; // 6008 : 255 - 0xff
      13'h1779: dout <= 8'b11111111; // 6009 : 255 - 0xff
      13'h177A: dout <= 8'b11111111; // 6010 : 255 - 0xff
      13'h177B: dout <= 8'b11111111; // 6011 : 255 - 0xff
      13'h177C: dout <= 8'b11111111; // 6012 : 255 - 0xff
      13'h177D: dout <= 8'b11111111; // 6013 : 255 - 0xff
      13'h177E: dout <= 8'b11111111; // 6014 : 255 - 0xff
      13'h177F: dout <= 8'b11111111; // 6015 : 255 - 0xff
      13'h1780: dout <= 8'b11111111; // 6016 : 255 - 0xff -- Background 0x78
      13'h1781: dout <= 8'b11111111; // 6017 : 255 - 0xff
      13'h1782: dout <= 8'b11111111; // 6018 : 255 - 0xff
      13'h1783: dout <= 8'b11111111; // 6019 : 255 - 0xff
      13'h1784: dout <= 8'b11111111; // 6020 : 255 - 0xff
      13'h1785: dout <= 8'b11111111; // 6021 : 255 - 0xff
      13'h1786: dout <= 8'b11111111; // 6022 : 255 - 0xff
      13'h1787: dout <= 8'b11111111; // 6023 : 255 - 0xff
      13'h1788: dout <= 8'b11111111; // 6024 : 255 - 0xff
      13'h1789: dout <= 8'b11111111; // 6025 : 255 - 0xff
      13'h178A: dout <= 8'b11111111; // 6026 : 255 - 0xff
      13'h178B: dout <= 8'b11111111; // 6027 : 255 - 0xff
      13'h178C: dout <= 8'b11111111; // 6028 : 255 - 0xff
      13'h178D: dout <= 8'b11111111; // 6029 : 255 - 0xff
      13'h178E: dout <= 8'b11111111; // 6030 : 255 - 0xff
      13'h178F: dout <= 8'b11111111; // 6031 : 255 - 0xff
      13'h1790: dout <= 8'b11111111; // 6032 : 255 - 0xff -- Background 0x79
      13'h1791: dout <= 8'b11111111; // 6033 : 255 - 0xff
      13'h1792: dout <= 8'b11111111; // 6034 : 255 - 0xff
      13'h1793: dout <= 8'b11111111; // 6035 : 255 - 0xff
      13'h1794: dout <= 8'b11111111; // 6036 : 255 - 0xff
      13'h1795: dout <= 8'b11111111; // 6037 : 255 - 0xff
      13'h1796: dout <= 8'b11111111; // 6038 : 255 - 0xff
      13'h1797: dout <= 8'b11111111; // 6039 : 255 - 0xff
      13'h1798: dout <= 8'b11111111; // 6040 : 255 - 0xff
      13'h1799: dout <= 8'b11111111; // 6041 : 255 - 0xff
      13'h179A: dout <= 8'b11111111; // 6042 : 255 - 0xff
      13'h179B: dout <= 8'b11111111; // 6043 : 255 - 0xff
      13'h179C: dout <= 8'b11111111; // 6044 : 255 - 0xff
      13'h179D: dout <= 8'b11111111; // 6045 : 255 - 0xff
      13'h179E: dout <= 8'b11111111; // 6046 : 255 - 0xff
      13'h179F: dout <= 8'b11111111; // 6047 : 255 - 0xff
      13'h17A0: dout <= 8'b11111111; // 6048 : 255 - 0xff -- Background 0x7a
      13'h17A1: dout <= 8'b11111111; // 6049 : 255 - 0xff
      13'h17A2: dout <= 8'b11111111; // 6050 : 255 - 0xff
      13'h17A3: dout <= 8'b11111111; // 6051 : 255 - 0xff
      13'h17A4: dout <= 8'b11111111; // 6052 : 255 - 0xff
      13'h17A5: dout <= 8'b11111111; // 6053 : 255 - 0xff
      13'h17A6: dout <= 8'b11111111; // 6054 : 255 - 0xff
      13'h17A7: dout <= 8'b11111111; // 6055 : 255 - 0xff
      13'h17A8: dout <= 8'b11111111; // 6056 : 255 - 0xff
      13'h17A9: dout <= 8'b11111111; // 6057 : 255 - 0xff
      13'h17AA: dout <= 8'b11111111; // 6058 : 255 - 0xff
      13'h17AB: dout <= 8'b11111111; // 6059 : 255 - 0xff
      13'h17AC: dout <= 8'b11111111; // 6060 : 255 - 0xff
      13'h17AD: dout <= 8'b11111111; // 6061 : 255 - 0xff
      13'h17AE: dout <= 8'b11111111; // 6062 : 255 - 0xff
      13'h17AF: dout <= 8'b11111111; // 6063 : 255 - 0xff
      13'h17B0: dout <= 8'b11111111; // 6064 : 255 - 0xff -- Background 0x7b
      13'h17B1: dout <= 8'b11111111; // 6065 : 255 - 0xff
      13'h17B2: dout <= 8'b11111111; // 6066 : 255 - 0xff
      13'h17B3: dout <= 8'b11111111; // 6067 : 255 - 0xff
      13'h17B4: dout <= 8'b11111111; // 6068 : 255 - 0xff
      13'h17B5: dout <= 8'b11111111; // 6069 : 255 - 0xff
      13'h17B6: dout <= 8'b11111111; // 6070 : 255 - 0xff
      13'h17B7: dout <= 8'b11111111; // 6071 : 255 - 0xff
      13'h17B8: dout <= 8'b11111111; // 6072 : 255 - 0xff
      13'h17B9: dout <= 8'b11111111; // 6073 : 255 - 0xff
      13'h17BA: dout <= 8'b11111111; // 6074 : 255 - 0xff
      13'h17BB: dout <= 8'b11111111; // 6075 : 255 - 0xff
      13'h17BC: dout <= 8'b11111111; // 6076 : 255 - 0xff
      13'h17BD: dout <= 8'b11111111; // 6077 : 255 - 0xff
      13'h17BE: dout <= 8'b11111111; // 6078 : 255 - 0xff
      13'h17BF: dout <= 8'b11111111; // 6079 : 255 - 0xff
      13'h17C0: dout <= 8'b11111111; // 6080 : 255 - 0xff -- Background 0x7c
      13'h17C1: dout <= 8'b11111111; // 6081 : 255 - 0xff
      13'h17C2: dout <= 8'b11111111; // 6082 : 255 - 0xff
      13'h17C3: dout <= 8'b11111111; // 6083 : 255 - 0xff
      13'h17C4: dout <= 8'b11111111; // 6084 : 255 - 0xff
      13'h17C5: dout <= 8'b11111111; // 6085 : 255 - 0xff
      13'h17C6: dout <= 8'b11111111; // 6086 : 255 - 0xff
      13'h17C7: dout <= 8'b11111111; // 6087 : 255 - 0xff
      13'h17C8: dout <= 8'b11111111; // 6088 : 255 - 0xff
      13'h17C9: dout <= 8'b11111111; // 6089 : 255 - 0xff
      13'h17CA: dout <= 8'b11111111; // 6090 : 255 - 0xff
      13'h17CB: dout <= 8'b11111111; // 6091 : 255 - 0xff
      13'h17CC: dout <= 8'b11111111; // 6092 : 255 - 0xff
      13'h17CD: dout <= 8'b11111111; // 6093 : 255 - 0xff
      13'h17CE: dout <= 8'b11111111; // 6094 : 255 - 0xff
      13'h17CF: dout <= 8'b11111111; // 6095 : 255 - 0xff
      13'h17D0: dout <= 8'b11111111; // 6096 : 255 - 0xff -- Background 0x7d
      13'h17D1: dout <= 8'b11111111; // 6097 : 255 - 0xff
      13'h17D2: dout <= 8'b11111111; // 6098 : 255 - 0xff
      13'h17D3: dout <= 8'b11111111; // 6099 : 255 - 0xff
      13'h17D4: dout <= 8'b11111111; // 6100 : 255 - 0xff
      13'h17D5: dout <= 8'b11111111; // 6101 : 255 - 0xff
      13'h17D6: dout <= 8'b11111111; // 6102 : 255 - 0xff
      13'h17D7: dout <= 8'b11111111; // 6103 : 255 - 0xff
      13'h17D8: dout <= 8'b11111111; // 6104 : 255 - 0xff
      13'h17D9: dout <= 8'b11111111; // 6105 : 255 - 0xff
      13'h17DA: dout <= 8'b11111111; // 6106 : 255 - 0xff
      13'h17DB: dout <= 8'b11111111; // 6107 : 255 - 0xff
      13'h17DC: dout <= 8'b11111111; // 6108 : 255 - 0xff
      13'h17DD: dout <= 8'b11111111; // 6109 : 255 - 0xff
      13'h17DE: dout <= 8'b11111111; // 6110 : 255 - 0xff
      13'h17DF: dout <= 8'b11111111; // 6111 : 255 - 0xff
      13'h17E0: dout <= 8'b11111111; // 6112 : 255 - 0xff -- Background 0x7e
      13'h17E1: dout <= 8'b11111111; // 6113 : 255 - 0xff
      13'h17E2: dout <= 8'b11111111; // 6114 : 255 - 0xff
      13'h17E3: dout <= 8'b11111111; // 6115 : 255 - 0xff
      13'h17E4: dout <= 8'b11111111; // 6116 : 255 - 0xff
      13'h17E5: dout <= 8'b11111111; // 6117 : 255 - 0xff
      13'h17E6: dout <= 8'b11111111; // 6118 : 255 - 0xff
      13'h17E7: dout <= 8'b11111111; // 6119 : 255 - 0xff
      13'h17E8: dout <= 8'b11111111; // 6120 : 255 - 0xff
      13'h17E9: dout <= 8'b11111111; // 6121 : 255 - 0xff
      13'h17EA: dout <= 8'b11111111; // 6122 : 255 - 0xff
      13'h17EB: dout <= 8'b11111111; // 6123 : 255 - 0xff
      13'h17EC: dout <= 8'b11111111; // 6124 : 255 - 0xff
      13'h17ED: dout <= 8'b11111111; // 6125 : 255 - 0xff
      13'h17EE: dout <= 8'b11111111; // 6126 : 255 - 0xff
      13'h17EF: dout <= 8'b11111111; // 6127 : 255 - 0xff
      13'h17F0: dout <= 8'b11111111; // 6128 : 255 - 0xff -- Background 0x7f
      13'h17F1: dout <= 8'b11111111; // 6129 : 255 - 0xff
      13'h17F2: dout <= 8'b11111111; // 6130 : 255 - 0xff
      13'h17F3: dout <= 8'b11111111; // 6131 : 255 - 0xff
      13'h17F4: dout <= 8'b11111111; // 6132 : 255 - 0xff
      13'h17F5: dout <= 8'b11111111; // 6133 : 255 - 0xff
      13'h17F6: dout <= 8'b11111111; // 6134 : 255 - 0xff
      13'h17F7: dout <= 8'b11111111; // 6135 : 255 - 0xff
      13'h17F8: dout <= 8'b11111111; // 6136 : 255 - 0xff
      13'h17F9: dout <= 8'b11111111; // 6137 : 255 - 0xff
      13'h17FA: dout <= 8'b11111111; // 6138 : 255 - 0xff
      13'h17FB: dout <= 8'b11111111; // 6139 : 255 - 0xff
      13'h17FC: dout <= 8'b11111111; // 6140 : 255 - 0xff
      13'h17FD: dout <= 8'b11111111; // 6141 : 255 - 0xff
      13'h17FE: dout <= 8'b11111111; // 6142 : 255 - 0xff
      13'h17FF: dout <= 8'b11111111; // 6143 : 255 - 0xff
      13'h1800: dout <= 8'b11111111; // 6144 : 255 - 0xff -- Background 0x80
      13'h1801: dout <= 8'b11111111; // 6145 : 255 - 0xff
      13'h1802: dout <= 8'b11111111; // 6146 : 255 - 0xff
      13'h1803: dout <= 8'b11111111; // 6147 : 255 - 0xff
      13'h1804: dout <= 8'b11111111; // 6148 : 255 - 0xff
      13'h1805: dout <= 8'b11111111; // 6149 : 255 - 0xff
      13'h1806: dout <= 8'b11111111; // 6150 : 255 - 0xff
      13'h1807: dout <= 8'b11111111; // 6151 : 255 - 0xff
      13'h1808: dout <= 8'b11111111; // 6152 : 255 - 0xff
      13'h1809: dout <= 8'b11111111; // 6153 : 255 - 0xff
      13'h180A: dout <= 8'b11111111; // 6154 : 255 - 0xff
      13'h180B: dout <= 8'b11111111; // 6155 : 255 - 0xff
      13'h180C: dout <= 8'b11111111; // 6156 : 255 - 0xff
      13'h180D: dout <= 8'b11111111; // 6157 : 255 - 0xff
      13'h180E: dout <= 8'b11111111; // 6158 : 255 - 0xff
      13'h180F: dout <= 8'b11111111; // 6159 : 255 - 0xff
      13'h1810: dout <= 8'b11111111; // 6160 : 255 - 0xff -- Background 0x81
      13'h1811: dout <= 8'b11111111; // 6161 : 255 - 0xff
      13'h1812: dout <= 8'b11111111; // 6162 : 255 - 0xff
      13'h1813: dout <= 8'b11111111; // 6163 : 255 - 0xff
      13'h1814: dout <= 8'b11111111; // 6164 : 255 - 0xff
      13'h1815: dout <= 8'b11111111; // 6165 : 255 - 0xff
      13'h1816: dout <= 8'b11111111; // 6166 : 255 - 0xff
      13'h1817: dout <= 8'b11111111; // 6167 : 255 - 0xff
      13'h1818: dout <= 8'b11111111; // 6168 : 255 - 0xff
      13'h1819: dout <= 8'b11111111; // 6169 : 255 - 0xff
      13'h181A: dout <= 8'b11111111; // 6170 : 255 - 0xff
      13'h181B: dout <= 8'b11111111; // 6171 : 255 - 0xff
      13'h181C: dout <= 8'b11111111; // 6172 : 255 - 0xff
      13'h181D: dout <= 8'b11111111; // 6173 : 255 - 0xff
      13'h181E: dout <= 8'b11111111; // 6174 : 255 - 0xff
      13'h181F: dout <= 8'b11111111; // 6175 : 255 - 0xff
      13'h1820: dout <= 8'b11111111; // 6176 : 255 - 0xff -- Background 0x82
      13'h1821: dout <= 8'b11111111; // 6177 : 255 - 0xff
      13'h1822: dout <= 8'b11111111; // 6178 : 255 - 0xff
      13'h1823: dout <= 8'b11111111; // 6179 : 255 - 0xff
      13'h1824: dout <= 8'b11111111; // 6180 : 255 - 0xff
      13'h1825: dout <= 8'b11111111; // 6181 : 255 - 0xff
      13'h1826: dout <= 8'b11111111; // 6182 : 255 - 0xff
      13'h1827: dout <= 8'b11111111; // 6183 : 255 - 0xff
      13'h1828: dout <= 8'b11111111; // 6184 : 255 - 0xff
      13'h1829: dout <= 8'b11111111; // 6185 : 255 - 0xff
      13'h182A: dout <= 8'b11111111; // 6186 : 255 - 0xff
      13'h182B: dout <= 8'b11111111; // 6187 : 255 - 0xff
      13'h182C: dout <= 8'b11111111; // 6188 : 255 - 0xff
      13'h182D: dout <= 8'b11111111; // 6189 : 255 - 0xff
      13'h182E: dout <= 8'b11111111; // 6190 : 255 - 0xff
      13'h182F: dout <= 8'b11111111; // 6191 : 255 - 0xff
      13'h1830: dout <= 8'b11111111; // 6192 : 255 - 0xff -- Background 0x83
      13'h1831: dout <= 8'b11111111; // 6193 : 255 - 0xff
      13'h1832: dout <= 8'b11111111; // 6194 : 255 - 0xff
      13'h1833: dout <= 8'b11111111; // 6195 : 255 - 0xff
      13'h1834: dout <= 8'b11111111; // 6196 : 255 - 0xff
      13'h1835: dout <= 8'b11111111; // 6197 : 255 - 0xff
      13'h1836: dout <= 8'b11111111; // 6198 : 255 - 0xff
      13'h1837: dout <= 8'b11111111; // 6199 : 255 - 0xff
      13'h1838: dout <= 8'b11111111; // 6200 : 255 - 0xff
      13'h1839: dout <= 8'b11111111; // 6201 : 255 - 0xff
      13'h183A: dout <= 8'b11111111; // 6202 : 255 - 0xff
      13'h183B: dout <= 8'b11111111; // 6203 : 255 - 0xff
      13'h183C: dout <= 8'b11111111; // 6204 : 255 - 0xff
      13'h183D: dout <= 8'b11111111; // 6205 : 255 - 0xff
      13'h183E: dout <= 8'b11111111; // 6206 : 255 - 0xff
      13'h183F: dout <= 8'b11111111; // 6207 : 255 - 0xff
      13'h1840: dout <= 8'b11111111; // 6208 : 255 - 0xff -- Background 0x84
      13'h1841: dout <= 8'b11111111; // 6209 : 255 - 0xff
      13'h1842: dout <= 8'b11111111; // 6210 : 255 - 0xff
      13'h1843: dout <= 8'b11111111; // 6211 : 255 - 0xff
      13'h1844: dout <= 8'b11111111; // 6212 : 255 - 0xff
      13'h1845: dout <= 8'b11111111; // 6213 : 255 - 0xff
      13'h1846: dout <= 8'b11111111; // 6214 : 255 - 0xff
      13'h1847: dout <= 8'b11111111; // 6215 : 255 - 0xff
      13'h1848: dout <= 8'b11111111; // 6216 : 255 - 0xff
      13'h1849: dout <= 8'b11111111; // 6217 : 255 - 0xff
      13'h184A: dout <= 8'b11111111; // 6218 : 255 - 0xff
      13'h184B: dout <= 8'b11111111; // 6219 : 255 - 0xff
      13'h184C: dout <= 8'b11111111; // 6220 : 255 - 0xff
      13'h184D: dout <= 8'b11111111; // 6221 : 255 - 0xff
      13'h184E: dout <= 8'b11111111; // 6222 : 255 - 0xff
      13'h184F: dout <= 8'b11111111; // 6223 : 255 - 0xff
      13'h1850: dout <= 8'b11111111; // 6224 : 255 - 0xff -- Background 0x85
      13'h1851: dout <= 8'b11111111; // 6225 : 255 - 0xff
      13'h1852: dout <= 8'b11111111; // 6226 : 255 - 0xff
      13'h1853: dout <= 8'b11111111; // 6227 : 255 - 0xff
      13'h1854: dout <= 8'b11111111; // 6228 : 255 - 0xff
      13'h1855: dout <= 8'b11111111; // 6229 : 255 - 0xff
      13'h1856: dout <= 8'b11111111; // 6230 : 255 - 0xff
      13'h1857: dout <= 8'b11111111; // 6231 : 255 - 0xff
      13'h1858: dout <= 8'b11111111; // 6232 : 255 - 0xff
      13'h1859: dout <= 8'b11111111; // 6233 : 255 - 0xff
      13'h185A: dout <= 8'b11111111; // 6234 : 255 - 0xff
      13'h185B: dout <= 8'b11111111; // 6235 : 255 - 0xff
      13'h185C: dout <= 8'b11111111; // 6236 : 255 - 0xff
      13'h185D: dout <= 8'b11111111; // 6237 : 255 - 0xff
      13'h185E: dout <= 8'b11111111; // 6238 : 255 - 0xff
      13'h185F: dout <= 8'b11111111; // 6239 : 255 - 0xff
      13'h1860: dout <= 8'b11111111; // 6240 : 255 - 0xff -- Background 0x86
      13'h1861: dout <= 8'b11111111; // 6241 : 255 - 0xff
      13'h1862: dout <= 8'b11111111; // 6242 : 255 - 0xff
      13'h1863: dout <= 8'b11111111; // 6243 : 255 - 0xff
      13'h1864: dout <= 8'b11111111; // 6244 : 255 - 0xff
      13'h1865: dout <= 8'b11111111; // 6245 : 255 - 0xff
      13'h1866: dout <= 8'b11111111; // 6246 : 255 - 0xff
      13'h1867: dout <= 8'b11111111; // 6247 : 255 - 0xff
      13'h1868: dout <= 8'b11111111; // 6248 : 255 - 0xff
      13'h1869: dout <= 8'b11111111; // 6249 : 255 - 0xff
      13'h186A: dout <= 8'b11111111; // 6250 : 255 - 0xff
      13'h186B: dout <= 8'b11111111; // 6251 : 255 - 0xff
      13'h186C: dout <= 8'b11111111; // 6252 : 255 - 0xff
      13'h186D: dout <= 8'b11111111; // 6253 : 255 - 0xff
      13'h186E: dout <= 8'b11111111; // 6254 : 255 - 0xff
      13'h186F: dout <= 8'b11111111; // 6255 : 255 - 0xff
      13'h1870: dout <= 8'b11111111; // 6256 : 255 - 0xff -- Background 0x87
      13'h1871: dout <= 8'b11111111; // 6257 : 255 - 0xff
      13'h1872: dout <= 8'b11111111; // 6258 : 255 - 0xff
      13'h1873: dout <= 8'b11111111; // 6259 : 255 - 0xff
      13'h1874: dout <= 8'b11111111; // 6260 : 255 - 0xff
      13'h1875: dout <= 8'b11111111; // 6261 : 255 - 0xff
      13'h1876: dout <= 8'b11111111; // 6262 : 255 - 0xff
      13'h1877: dout <= 8'b11111111; // 6263 : 255 - 0xff
      13'h1878: dout <= 8'b11111111; // 6264 : 255 - 0xff
      13'h1879: dout <= 8'b11111111; // 6265 : 255 - 0xff
      13'h187A: dout <= 8'b11111111; // 6266 : 255 - 0xff
      13'h187B: dout <= 8'b11111111; // 6267 : 255 - 0xff
      13'h187C: dout <= 8'b11111111; // 6268 : 255 - 0xff
      13'h187D: dout <= 8'b11111111; // 6269 : 255 - 0xff
      13'h187E: dout <= 8'b11111111; // 6270 : 255 - 0xff
      13'h187F: dout <= 8'b11111111; // 6271 : 255 - 0xff
      13'h1880: dout <= 8'b11111111; // 6272 : 255 - 0xff -- Background 0x88
      13'h1881: dout <= 8'b11111111; // 6273 : 255 - 0xff
      13'h1882: dout <= 8'b11111111; // 6274 : 255 - 0xff
      13'h1883: dout <= 8'b11111111; // 6275 : 255 - 0xff
      13'h1884: dout <= 8'b11111111; // 6276 : 255 - 0xff
      13'h1885: dout <= 8'b11111111; // 6277 : 255 - 0xff
      13'h1886: dout <= 8'b11111111; // 6278 : 255 - 0xff
      13'h1887: dout <= 8'b11111111; // 6279 : 255 - 0xff
      13'h1888: dout <= 8'b11111111; // 6280 : 255 - 0xff
      13'h1889: dout <= 8'b11111111; // 6281 : 255 - 0xff
      13'h188A: dout <= 8'b11111111; // 6282 : 255 - 0xff
      13'h188B: dout <= 8'b11111111; // 6283 : 255 - 0xff
      13'h188C: dout <= 8'b11111111; // 6284 : 255 - 0xff
      13'h188D: dout <= 8'b11111111; // 6285 : 255 - 0xff
      13'h188E: dout <= 8'b11111111; // 6286 : 255 - 0xff
      13'h188F: dout <= 8'b11111111; // 6287 : 255 - 0xff
      13'h1890: dout <= 8'b11111111; // 6288 : 255 - 0xff -- Background 0x89
      13'h1891: dout <= 8'b11111111; // 6289 : 255 - 0xff
      13'h1892: dout <= 8'b11111111; // 6290 : 255 - 0xff
      13'h1893: dout <= 8'b11111111; // 6291 : 255 - 0xff
      13'h1894: dout <= 8'b11111111; // 6292 : 255 - 0xff
      13'h1895: dout <= 8'b11111111; // 6293 : 255 - 0xff
      13'h1896: dout <= 8'b11111111; // 6294 : 255 - 0xff
      13'h1897: dout <= 8'b11111111; // 6295 : 255 - 0xff
      13'h1898: dout <= 8'b11111111; // 6296 : 255 - 0xff
      13'h1899: dout <= 8'b11111111; // 6297 : 255 - 0xff
      13'h189A: dout <= 8'b11111111; // 6298 : 255 - 0xff
      13'h189B: dout <= 8'b11111111; // 6299 : 255 - 0xff
      13'h189C: dout <= 8'b11111111; // 6300 : 255 - 0xff
      13'h189D: dout <= 8'b11111111; // 6301 : 255 - 0xff
      13'h189E: dout <= 8'b11111111; // 6302 : 255 - 0xff
      13'h189F: dout <= 8'b11111111; // 6303 : 255 - 0xff
      13'h18A0: dout <= 8'b11111111; // 6304 : 255 - 0xff -- Background 0x8a
      13'h18A1: dout <= 8'b11111111; // 6305 : 255 - 0xff
      13'h18A2: dout <= 8'b11111111; // 6306 : 255 - 0xff
      13'h18A3: dout <= 8'b11111111; // 6307 : 255 - 0xff
      13'h18A4: dout <= 8'b11111111; // 6308 : 255 - 0xff
      13'h18A5: dout <= 8'b11111111; // 6309 : 255 - 0xff
      13'h18A6: dout <= 8'b11111111; // 6310 : 255 - 0xff
      13'h18A7: dout <= 8'b11111111; // 6311 : 255 - 0xff
      13'h18A8: dout <= 8'b11111111; // 6312 : 255 - 0xff
      13'h18A9: dout <= 8'b11111111; // 6313 : 255 - 0xff
      13'h18AA: dout <= 8'b11111111; // 6314 : 255 - 0xff
      13'h18AB: dout <= 8'b11111111; // 6315 : 255 - 0xff
      13'h18AC: dout <= 8'b11111111; // 6316 : 255 - 0xff
      13'h18AD: dout <= 8'b11111111; // 6317 : 255 - 0xff
      13'h18AE: dout <= 8'b11111111; // 6318 : 255 - 0xff
      13'h18AF: dout <= 8'b11111111; // 6319 : 255 - 0xff
      13'h18B0: dout <= 8'b11111111; // 6320 : 255 - 0xff -- Background 0x8b
      13'h18B1: dout <= 8'b11111111; // 6321 : 255 - 0xff
      13'h18B2: dout <= 8'b11111111; // 6322 : 255 - 0xff
      13'h18B3: dout <= 8'b11111111; // 6323 : 255 - 0xff
      13'h18B4: dout <= 8'b11111111; // 6324 : 255 - 0xff
      13'h18B5: dout <= 8'b11111111; // 6325 : 255 - 0xff
      13'h18B6: dout <= 8'b11111111; // 6326 : 255 - 0xff
      13'h18B7: dout <= 8'b11111111; // 6327 : 255 - 0xff
      13'h18B8: dout <= 8'b11111111; // 6328 : 255 - 0xff
      13'h18B9: dout <= 8'b11111111; // 6329 : 255 - 0xff
      13'h18BA: dout <= 8'b11111111; // 6330 : 255 - 0xff
      13'h18BB: dout <= 8'b11111111; // 6331 : 255 - 0xff
      13'h18BC: dout <= 8'b11111111; // 6332 : 255 - 0xff
      13'h18BD: dout <= 8'b11111111; // 6333 : 255 - 0xff
      13'h18BE: dout <= 8'b11111111; // 6334 : 255 - 0xff
      13'h18BF: dout <= 8'b11111111; // 6335 : 255 - 0xff
      13'h18C0: dout <= 8'b11111111; // 6336 : 255 - 0xff -- Background 0x8c
      13'h18C1: dout <= 8'b11111111; // 6337 : 255 - 0xff
      13'h18C2: dout <= 8'b11111111; // 6338 : 255 - 0xff
      13'h18C3: dout <= 8'b11111111; // 6339 : 255 - 0xff
      13'h18C4: dout <= 8'b11111111; // 6340 : 255 - 0xff
      13'h18C5: dout <= 8'b11111111; // 6341 : 255 - 0xff
      13'h18C6: dout <= 8'b11111111; // 6342 : 255 - 0xff
      13'h18C7: dout <= 8'b11111111; // 6343 : 255 - 0xff
      13'h18C8: dout <= 8'b11111111; // 6344 : 255 - 0xff
      13'h18C9: dout <= 8'b11111111; // 6345 : 255 - 0xff
      13'h18CA: dout <= 8'b11111111; // 6346 : 255 - 0xff
      13'h18CB: dout <= 8'b11111111; // 6347 : 255 - 0xff
      13'h18CC: dout <= 8'b11111111; // 6348 : 255 - 0xff
      13'h18CD: dout <= 8'b11111111; // 6349 : 255 - 0xff
      13'h18CE: dout <= 8'b11111111; // 6350 : 255 - 0xff
      13'h18CF: dout <= 8'b11111111; // 6351 : 255 - 0xff
      13'h18D0: dout <= 8'b11111111; // 6352 : 255 - 0xff -- Background 0x8d
      13'h18D1: dout <= 8'b11111111; // 6353 : 255 - 0xff
      13'h18D2: dout <= 8'b11111111; // 6354 : 255 - 0xff
      13'h18D3: dout <= 8'b11111111; // 6355 : 255 - 0xff
      13'h18D4: dout <= 8'b11111111; // 6356 : 255 - 0xff
      13'h18D5: dout <= 8'b11111111; // 6357 : 255 - 0xff
      13'h18D6: dout <= 8'b11111111; // 6358 : 255 - 0xff
      13'h18D7: dout <= 8'b11111111; // 6359 : 255 - 0xff
      13'h18D8: dout <= 8'b11111111; // 6360 : 255 - 0xff
      13'h18D9: dout <= 8'b11111111; // 6361 : 255 - 0xff
      13'h18DA: dout <= 8'b11111111; // 6362 : 255 - 0xff
      13'h18DB: dout <= 8'b11111111; // 6363 : 255 - 0xff
      13'h18DC: dout <= 8'b11111111; // 6364 : 255 - 0xff
      13'h18DD: dout <= 8'b11111111; // 6365 : 255 - 0xff
      13'h18DE: dout <= 8'b11111111; // 6366 : 255 - 0xff
      13'h18DF: dout <= 8'b11111111; // 6367 : 255 - 0xff
      13'h18E0: dout <= 8'b11111111; // 6368 : 255 - 0xff -- Background 0x8e
      13'h18E1: dout <= 8'b11111111; // 6369 : 255 - 0xff
      13'h18E2: dout <= 8'b11111111; // 6370 : 255 - 0xff
      13'h18E3: dout <= 8'b11111111; // 6371 : 255 - 0xff
      13'h18E4: dout <= 8'b11111111; // 6372 : 255 - 0xff
      13'h18E5: dout <= 8'b11111111; // 6373 : 255 - 0xff
      13'h18E6: dout <= 8'b11111111; // 6374 : 255 - 0xff
      13'h18E7: dout <= 8'b11111111; // 6375 : 255 - 0xff
      13'h18E8: dout <= 8'b11111111; // 6376 : 255 - 0xff
      13'h18E9: dout <= 8'b11111111; // 6377 : 255 - 0xff
      13'h18EA: dout <= 8'b11111111; // 6378 : 255 - 0xff
      13'h18EB: dout <= 8'b11111111; // 6379 : 255 - 0xff
      13'h18EC: dout <= 8'b11111111; // 6380 : 255 - 0xff
      13'h18ED: dout <= 8'b11111111; // 6381 : 255 - 0xff
      13'h18EE: dout <= 8'b11111111; // 6382 : 255 - 0xff
      13'h18EF: dout <= 8'b11111111; // 6383 : 255 - 0xff
      13'h18F0: dout <= 8'b11111111; // 6384 : 255 - 0xff -- Background 0x8f
      13'h18F1: dout <= 8'b11111111; // 6385 : 255 - 0xff
      13'h18F2: dout <= 8'b11111111; // 6386 : 255 - 0xff
      13'h18F3: dout <= 8'b11111111; // 6387 : 255 - 0xff
      13'h18F4: dout <= 8'b11111111; // 6388 : 255 - 0xff
      13'h18F5: dout <= 8'b11111111; // 6389 : 255 - 0xff
      13'h18F6: dout <= 8'b11111111; // 6390 : 255 - 0xff
      13'h18F7: dout <= 8'b11111111; // 6391 : 255 - 0xff
      13'h18F8: dout <= 8'b11111111; // 6392 : 255 - 0xff
      13'h18F9: dout <= 8'b11111111; // 6393 : 255 - 0xff
      13'h18FA: dout <= 8'b11111111; // 6394 : 255 - 0xff
      13'h18FB: dout <= 8'b11111111; // 6395 : 255 - 0xff
      13'h18FC: dout <= 8'b11111111; // 6396 : 255 - 0xff
      13'h18FD: dout <= 8'b11111111; // 6397 : 255 - 0xff
      13'h18FE: dout <= 8'b11111111; // 6398 : 255 - 0xff
      13'h18FF: dout <= 8'b11111111; // 6399 : 255 - 0xff
      13'h1900: dout <= 8'b00000000; // 6400 :   0 - 0x0 -- Background 0x90
      13'h1901: dout <= 8'b00000000; // 6401 :   0 - 0x0
      13'h1902: dout <= 8'b00000000; // 6402 :   0 - 0x0
      13'h1903: dout <= 8'b00000000; // 6403 :   0 - 0x0
      13'h1904: dout <= 8'b00000000; // 6404 :   0 - 0x0
      13'h1905: dout <= 8'b00000001; // 6405 :   1 - 0x1
      13'h1906: dout <= 8'b00011110; // 6406 :  30 - 0x1e
      13'h1907: dout <= 8'b00111011; // 6407 :  59 - 0x3b
      13'h1908: dout <= 8'b00000000; // 6408 :   0 - 0x0
      13'h1909: dout <= 8'b00000000; // 6409 :   0 - 0x0
      13'h190A: dout <= 8'b00000000; // 6410 :   0 - 0x0
      13'h190B: dout <= 8'b00000000; // 6411 :   0 - 0x0
      13'h190C: dout <= 8'b00000000; // 6412 :   0 - 0x0
      13'h190D: dout <= 8'b00000000; // 6413 :   0 - 0x0
      13'h190E: dout <= 8'b00000000; // 6414 :   0 - 0x0
      13'h190F: dout <= 8'b00000000; // 6415 :   0 - 0x0
      13'h1910: dout <= 8'b00000000; // 6416 :   0 - 0x0 -- Background 0x91
      13'h1911: dout <= 8'b00000000; // 6417 :   0 - 0x0
      13'h1912: dout <= 8'b00001100; // 6418 :  12 - 0xc
      13'h1913: dout <= 8'b00111100; // 6419 :  60 - 0x3c
      13'h1914: dout <= 8'b11010000; // 6420 : 208 - 0xd0
      13'h1915: dout <= 8'b00010000; // 6421 :  16 - 0x10
      13'h1916: dout <= 8'b00100000; // 6422 :  32 - 0x20
      13'h1917: dout <= 8'b01000000; // 6423 :  64 - 0x40
      13'h1918: dout <= 8'b00000000; // 6424 :   0 - 0x0
      13'h1919: dout <= 8'b00000000; // 6425 :   0 - 0x0
      13'h191A: dout <= 8'b00000000; // 6426 :   0 - 0x0
      13'h191B: dout <= 8'b00000000; // 6427 :   0 - 0x0
      13'h191C: dout <= 8'b00000000; // 6428 :   0 - 0x0
      13'h191D: dout <= 8'b00000000; // 6429 :   0 - 0x0
      13'h191E: dout <= 8'b00000000; // 6430 :   0 - 0x0
      13'h191F: dout <= 8'b00000000; // 6431 :   0 - 0x0
      13'h1920: dout <= 8'b00111110; // 6432 :  62 - 0x3e -- Background 0x92
      13'h1921: dout <= 8'b00101101; // 6433 :  45 - 0x2d
      13'h1922: dout <= 8'b00110101; // 6434 :  53 - 0x35
      13'h1923: dout <= 8'b00011101; // 6435 :  29 - 0x1d
      13'h1924: dout <= 8'b00000001; // 6436 :   1 - 0x1
      13'h1925: dout <= 8'b00000000; // 6437 :   0 - 0x0
      13'h1926: dout <= 8'b00000000; // 6438 :   0 - 0x0
      13'h1927: dout <= 8'b00000000; // 6439 :   0 - 0x0
      13'h1928: dout <= 8'b00000000; // 6440 :   0 - 0x0
      13'h1929: dout <= 8'b00000000; // 6441 :   0 - 0x0
      13'h192A: dout <= 8'b00000000; // 6442 :   0 - 0x0
      13'h192B: dout <= 8'b00000000; // 6443 :   0 - 0x0
      13'h192C: dout <= 8'b00000000; // 6444 :   0 - 0x0
      13'h192D: dout <= 8'b00000000; // 6445 :   0 - 0x0
      13'h192E: dout <= 8'b00000000; // 6446 :   0 - 0x0
      13'h192F: dout <= 8'b00000000; // 6447 :   0 - 0x0
      13'h1930: dout <= 8'b10110000; // 6448 : 176 - 0xb0 -- Background 0x93
      13'h1931: dout <= 8'b10111000; // 6449 : 184 - 0xb8
      13'h1932: dout <= 8'b11111000; // 6450 : 248 - 0xf8
      13'h1933: dout <= 8'b01111000; // 6451 : 120 - 0x78
      13'h1934: dout <= 8'b10011000; // 6452 : 152 - 0x98
      13'h1935: dout <= 8'b11110000; // 6453 : 240 - 0xf0
      13'h1936: dout <= 8'b00000000; // 6454 :   0 - 0x0
      13'h1937: dout <= 8'b00000000; // 6455 :   0 - 0x0
      13'h1938: dout <= 8'b00000000; // 6456 :   0 - 0x0
      13'h1939: dout <= 8'b00000000; // 6457 :   0 - 0x0
      13'h193A: dout <= 8'b00000000; // 6458 :   0 - 0x0
      13'h193B: dout <= 8'b00000000; // 6459 :   0 - 0x0
      13'h193C: dout <= 8'b00000000; // 6460 :   0 - 0x0
      13'h193D: dout <= 8'b00000000; // 6461 :   0 - 0x0
      13'h193E: dout <= 8'b00000000; // 6462 :   0 - 0x0
      13'h193F: dout <= 8'b00000000; // 6463 :   0 - 0x0
      13'h1940: dout <= 8'b00000000; // 6464 :   0 - 0x0 -- Background 0x94
      13'h1941: dout <= 8'b00000000; // 6465 :   0 - 0x0
      13'h1942: dout <= 8'b00000111; // 6466 :   7 - 0x7
      13'h1943: dout <= 8'b00000011; // 6467 :   3 - 0x3
      13'h1944: dout <= 8'b00001101; // 6468 :  13 - 0xd
      13'h1945: dout <= 8'b00011110; // 6469 :  30 - 0x1e
      13'h1946: dout <= 8'b00010111; // 6470 :  23 - 0x17
      13'h1947: dout <= 8'b00011101; // 6471 :  29 - 0x1d
      13'h1948: dout <= 8'b00000000; // 6472 :   0 - 0x0
      13'h1949: dout <= 8'b00000000; // 6473 :   0 - 0x0
      13'h194A: dout <= 8'b00000000; // 6474 :   0 - 0x0
      13'h194B: dout <= 8'b00000000; // 6475 :   0 - 0x0
      13'h194C: dout <= 8'b00000000; // 6476 :   0 - 0x0
      13'h194D: dout <= 8'b00000000; // 6477 :   0 - 0x0
      13'h194E: dout <= 8'b00000000; // 6478 :   0 - 0x0
      13'h194F: dout <= 8'b00000000; // 6479 :   0 - 0x0
      13'h1950: dout <= 8'b00000000; // 6480 :   0 - 0x0 -- Background 0x95
      13'h1951: dout <= 8'b10000000; // 6481 : 128 - 0x80
      13'h1952: dout <= 8'b01110000; // 6482 : 112 - 0x70
      13'h1953: dout <= 8'b11100000; // 6483 : 224 - 0xe0
      13'h1954: dout <= 8'b11011000; // 6484 : 216 - 0xd8
      13'h1955: dout <= 8'b10111100; // 6485 : 188 - 0xbc
      13'h1956: dout <= 8'b01110100; // 6486 : 116 - 0x74
      13'h1957: dout <= 8'b11011100; // 6487 : 220 - 0xdc
      13'h1958: dout <= 8'b00000000; // 6488 :   0 - 0x0
      13'h1959: dout <= 8'b00000000; // 6489 :   0 - 0x0
      13'h195A: dout <= 8'b00000000; // 6490 :   0 - 0x0
      13'h195B: dout <= 8'b00000000; // 6491 :   0 - 0x0
      13'h195C: dout <= 8'b00000000; // 6492 :   0 - 0x0
      13'h195D: dout <= 8'b00000000; // 6493 :   0 - 0x0
      13'h195E: dout <= 8'b00000000; // 6494 :   0 - 0x0
      13'h195F: dout <= 8'b00000000; // 6495 :   0 - 0x0
      13'h1960: dout <= 8'b00011111; // 6496 :  31 - 0x1f -- Background 0x96
      13'h1961: dout <= 8'b00001011; // 6497 :  11 - 0xb
      13'h1962: dout <= 8'b00001111; // 6498 :  15 - 0xf
      13'h1963: dout <= 8'b00000101; // 6499 :   5 - 0x5
      13'h1964: dout <= 8'b00000011; // 6500 :   3 - 0x3
      13'h1965: dout <= 8'b00000001; // 6501 :   1 - 0x1
      13'h1966: dout <= 8'b00000000; // 6502 :   0 - 0x0
      13'h1967: dout <= 8'b00000000; // 6503 :   0 - 0x0
      13'h1968: dout <= 8'b00000000; // 6504 :   0 - 0x0
      13'h1969: dout <= 8'b00000000; // 6505 :   0 - 0x0
      13'h196A: dout <= 8'b00000000; // 6506 :   0 - 0x0
      13'h196B: dout <= 8'b00000000; // 6507 :   0 - 0x0
      13'h196C: dout <= 8'b00000000; // 6508 :   0 - 0x0
      13'h196D: dout <= 8'b00000000; // 6509 :   0 - 0x0
      13'h196E: dout <= 8'b00000000; // 6510 :   0 - 0x0
      13'h196F: dout <= 8'b00000000; // 6511 :   0 - 0x0
      13'h1970: dout <= 8'b11111100; // 6512 : 252 - 0xfc -- Background 0x97
      13'h1971: dout <= 8'b01101000; // 6513 : 104 - 0x68
      13'h1972: dout <= 8'b11111000; // 6514 : 248 - 0xf8
      13'h1973: dout <= 8'b10110000; // 6515 : 176 - 0xb0
      13'h1974: dout <= 8'b11100000; // 6516 : 224 - 0xe0
      13'h1975: dout <= 8'b10000000; // 6517 : 128 - 0x80
      13'h1976: dout <= 8'b00000000; // 6518 :   0 - 0x0
      13'h1977: dout <= 8'b00000000; // 6519 :   0 - 0x0
      13'h1978: dout <= 8'b00000000; // 6520 :   0 - 0x0
      13'h1979: dout <= 8'b00000000; // 6521 :   0 - 0x0
      13'h197A: dout <= 8'b00000000; // 6522 :   0 - 0x0
      13'h197B: dout <= 8'b00000000; // 6523 :   0 - 0x0
      13'h197C: dout <= 8'b00000000; // 6524 :   0 - 0x0
      13'h197D: dout <= 8'b00000000; // 6525 :   0 - 0x0
      13'h197E: dout <= 8'b00000000; // 6526 :   0 - 0x0
      13'h197F: dout <= 8'b00000000; // 6527 :   0 - 0x0
      13'h1980: dout <= 8'b00000000; // 6528 :   0 - 0x0 -- Background 0x98
      13'h1981: dout <= 8'b00000000; // 6529 :   0 - 0x0
      13'h1982: dout <= 8'b00000000; // 6530 :   0 - 0x0
      13'h1983: dout <= 8'b00000001; // 6531 :   1 - 0x1
      13'h1984: dout <= 8'b00000001; // 6532 :   1 - 0x1
      13'h1985: dout <= 8'b00001011; // 6533 :  11 - 0xb
      13'h1986: dout <= 8'b00011100; // 6534 :  28 - 0x1c
      13'h1987: dout <= 8'b00111111; // 6535 :  63 - 0x3f
      13'h1988: dout <= 8'b00000000; // 6536 :   0 - 0x0
      13'h1989: dout <= 8'b00000000; // 6537 :   0 - 0x0
      13'h198A: dout <= 8'b00000000; // 6538 :   0 - 0x0
      13'h198B: dout <= 8'b00000000; // 6539 :   0 - 0x0
      13'h198C: dout <= 8'b00000000; // 6540 :   0 - 0x0
      13'h198D: dout <= 8'b00000000; // 6541 :   0 - 0x0
      13'h198E: dout <= 8'b00000000; // 6542 :   0 - 0x0
      13'h198F: dout <= 8'b00000000; // 6543 :   0 - 0x0
      13'h1990: dout <= 8'b00000000; // 6544 :   0 - 0x0 -- Background 0x99
      13'h1991: dout <= 8'b00000000; // 6545 :   0 - 0x0
      13'h1992: dout <= 8'b00110000; // 6546 :  48 - 0x30
      13'h1993: dout <= 8'b01111000; // 6547 : 120 - 0x78
      13'h1994: dout <= 8'b10000000; // 6548 : 128 - 0x80
      13'h1995: dout <= 8'b11110000; // 6549 : 240 - 0xf0
      13'h1996: dout <= 8'b11111000; // 6550 : 248 - 0xf8
      13'h1997: dout <= 8'b11111100; // 6551 : 252 - 0xfc
      13'h1998: dout <= 8'b00000000; // 6552 :   0 - 0x0
      13'h1999: dout <= 8'b00000000; // 6553 :   0 - 0x0
      13'h199A: dout <= 8'b00000000; // 6554 :   0 - 0x0
      13'h199B: dout <= 8'b00000000; // 6555 :   0 - 0x0
      13'h199C: dout <= 8'b00000000; // 6556 :   0 - 0x0
      13'h199D: dout <= 8'b00000000; // 6557 :   0 - 0x0
      13'h199E: dout <= 8'b00000000; // 6558 :   0 - 0x0
      13'h199F: dout <= 8'b00000000; // 6559 :   0 - 0x0
      13'h19A0: dout <= 8'b00111111; // 6560 :  63 - 0x3f -- Background 0x9a
      13'h19A1: dout <= 8'b00111111; // 6561 :  63 - 0x3f
      13'h19A2: dout <= 8'b00111111; // 6562 :  63 - 0x3f
      13'h19A3: dout <= 8'b00011111; // 6563 :  31 - 0x1f
      13'h19A4: dout <= 8'b00011111; // 6564 :  31 - 0x1f
      13'h19A5: dout <= 8'b00000111; // 6565 :   7 - 0x7
      13'h19A6: dout <= 8'b00000000; // 6566 :   0 - 0x0
      13'h19A7: dout <= 8'b00000000; // 6567 :   0 - 0x0
      13'h19A8: dout <= 8'b00000000; // 6568 :   0 - 0x0
      13'h19A9: dout <= 8'b00000000; // 6569 :   0 - 0x0
      13'h19AA: dout <= 8'b00000000; // 6570 :   0 - 0x0
      13'h19AB: dout <= 8'b00000000; // 6571 :   0 - 0x0
      13'h19AC: dout <= 8'b00000000; // 6572 :   0 - 0x0
      13'h19AD: dout <= 8'b00000000; // 6573 :   0 - 0x0
      13'h19AE: dout <= 8'b00000000; // 6574 :   0 - 0x0
      13'h19AF: dout <= 8'b00000000; // 6575 :   0 - 0x0
      13'h19B0: dout <= 8'b11111100; // 6576 : 252 - 0xfc -- Background 0x9b
      13'h19B1: dout <= 8'b11101100; // 6577 : 236 - 0xec
      13'h19B2: dout <= 8'b11101100; // 6578 : 236 - 0xec
      13'h19B3: dout <= 8'b11011000; // 6579 : 216 - 0xd8
      13'h19B4: dout <= 8'b11111000; // 6580 : 248 - 0xf8
      13'h19B5: dout <= 8'b11100000; // 6581 : 224 - 0xe0
      13'h19B6: dout <= 8'b00000000; // 6582 :   0 - 0x0
      13'h19B7: dout <= 8'b00000000; // 6583 :   0 - 0x0
      13'h19B8: dout <= 8'b00000000; // 6584 :   0 - 0x0
      13'h19B9: dout <= 8'b00000000; // 6585 :   0 - 0x0
      13'h19BA: dout <= 8'b00000000; // 6586 :   0 - 0x0
      13'h19BB: dout <= 8'b00000000; // 6587 :   0 - 0x0
      13'h19BC: dout <= 8'b00000000; // 6588 :   0 - 0x0
      13'h19BD: dout <= 8'b00000000; // 6589 :   0 - 0x0
      13'h19BE: dout <= 8'b00000000; // 6590 :   0 - 0x0
      13'h19BF: dout <= 8'b00000000; // 6591 :   0 - 0x0
      13'h19C0: dout <= 8'b00000000; // 6592 :   0 - 0x0 -- Background 0x9c
      13'h19C1: dout <= 8'b00000000; // 6593 :   0 - 0x0
      13'h19C2: dout <= 8'b00000001; // 6594 :   1 - 0x1
      13'h19C3: dout <= 8'b00011101; // 6595 :  29 - 0x1d
      13'h19C4: dout <= 8'b00111110; // 6596 :  62 - 0x3e
      13'h19C5: dout <= 8'b00111111; // 6597 :  63 - 0x3f
      13'h19C6: dout <= 8'b00111111; // 6598 :  63 - 0x3f
      13'h19C7: dout <= 8'b00111111; // 6599 :  63 - 0x3f
      13'h19C8: dout <= 8'b00000000; // 6600 :   0 - 0x0
      13'h19C9: dout <= 8'b00000000; // 6601 :   0 - 0x0
      13'h19CA: dout <= 8'b00000000; // 6602 :   0 - 0x0
      13'h19CB: dout <= 8'b00000000; // 6603 :   0 - 0x0
      13'h19CC: dout <= 8'b00000000; // 6604 :   0 - 0x0
      13'h19CD: dout <= 8'b00000000; // 6605 :   0 - 0x0
      13'h19CE: dout <= 8'b00000000; // 6606 :   0 - 0x0
      13'h19CF: dout <= 8'b00000000; // 6607 :   0 - 0x0
      13'h19D0: dout <= 8'b00000000; // 6608 :   0 - 0x0 -- Background 0x9d
      13'h19D1: dout <= 8'b10000000; // 6609 : 128 - 0x80
      13'h19D2: dout <= 8'b00000000; // 6610 :   0 - 0x0
      13'h19D3: dout <= 8'b01110000; // 6611 : 112 - 0x70
      13'h19D4: dout <= 8'b11111000; // 6612 : 248 - 0xf8
      13'h19D5: dout <= 8'b11111100; // 6613 : 252 - 0xfc
      13'h19D6: dout <= 8'b11111100; // 6614 : 252 - 0xfc
      13'h19D7: dout <= 8'b11111100; // 6615 : 252 - 0xfc
      13'h19D8: dout <= 8'b00000000; // 6616 :   0 - 0x0
      13'h19D9: dout <= 8'b00000000; // 6617 :   0 - 0x0
      13'h19DA: dout <= 8'b00000000; // 6618 :   0 - 0x0
      13'h19DB: dout <= 8'b00000000; // 6619 :   0 - 0x0
      13'h19DC: dout <= 8'b00000000; // 6620 :   0 - 0x0
      13'h19DD: dout <= 8'b00000000; // 6621 :   0 - 0x0
      13'h19DE: dout <= 8'b00000000; // 6622 :   0 - 0x0
      13'h19DF: dout <= 8'b00000000; // 6623 :   0 - 0x0
      13'h19E0: dout <= 8'b00111111; // 6624 :  63 - 0x3f -- Background 0x9e
      13'h19E1: dout <= 8'b00111111; // 6625 :  63 - 0x3f
      13'h19E2: dout <= 8'b00011111; // 6626 :  31 - 0x1f
      13'h19E3: dout <= 8'b00011111; // 6627 :  31 - 0x1f
      13'h19E4: dout <= 8'b00001111; // 6628 :  15 - 0xf
      13'h19E5: dout <= 8'b00000110; // 6629 :   6 - 0x6
      13'h19E6: dout <= 8'b00000000; // 6630 :   0 - 0x0
      13'h19E7: dout <= 8'b00000000; // 6631 :   0 - 0x0
      13'h19E8: dout <= 8'b00000000; // 6632 :   0 - 0x0
      13'h19E9: dout <= 8'b00000000; // 6633 :   0 - 0x0
      13'h19EA: dout <= 8'b00000000; // 6634 :   0 - 0x0
      13'h19EB: dout <= 8'b00000000; // 6635 :   0 - 0x0
      13'h19EC: dout <= 8'b00000000; // 6636 :   0 - 0x0
      13'h19ED: dout <= 8'b00000000; // 6637 :   0 - 0x0
      13'h19EE: dout <= 8'b00000000; // 6638 :   0 - 0x0
      13'h19EF: dout <= 8'b00000000; // 6639 :   0 - 0x0
      13'h19F0: dout <= 8'b11101100; // 6640 : 236 - 0xec -- Background 0x9f
      13'h19F1: dout <= 8'b11101100; // 6641 : 236 - 0xec
      13'h19F2: dout <= 8'b11011000; // 6642 : 216 - 0xd8
      13'h19F3: dout <= 8'b11111000; // 6643 : 248 - 0xf8
      13'h19F4: dout <= 8'b11110000; // 6644 : 240 - 0xf0
      13'h19F5: dout <= 8'b11100000; // 6645 : 224 - 0xe0
      13'h19F6: dout <= 8'b00000000; // 6646 :   0 - 0x0
      13'h19F7: dout <= 8'b00000000; // 6647 :   0 - 0x0
      13'h19F8: dout <= 8'b00000000; // 6648 :   0 - 0x0
      13'h19F9: dout <= 8'b00000000; // 6649 :   0 - 0x0
      13'h19FA: dout <= 8'b00000000; // 6650 :   0 - 0x0
      13'h19FB: dout <= 8'b00000000; // 6651 :   0 - 0x0
      13'h19FC: dout <= 8'b00000000; // 6652 :   0 - 0x0
      13'h19FD: dout <= 8'b00000000; // 6653 :   0 - 0x0
      13'h19FE: dout <= 8'b00000000; // 6654 :   0 - 0x0
      13'h19FF: dout <= 8'b00000000; // 6655 :   0 - 0x0
      13'h1A00: dout <= 8'b00000000; // 6656 :   0 - 0x0 -- Background 0xa0
      13'h1A01: dout <= 8'b00000100; // 6657 :   4 - 0x4
      13'h1A02: dout <= 8'b00000011; // 6658 :   3 - 0x3
      13'h1A03: dout <= 8'b00000000; // 6659 :   0 - 0x0
      13'h1A04: dout <= 8'b00000001; // 6660 :   1 - 0x1
      13'h1A05: dout <= 8'b00000111; // 6661 :   7 - 0x7
      13'h1A06: dout <= 8'b00001111; // 6662 :  15 - 0xf
      13'h1A07: dout <= 8'b00001100; // 6663 :  12 - 0xc
      13'h1A08: dout <= 8'b00000000; // 6664 :   0 - 0x0
      13'h1A09: dout <= 8'b00000000; // 6665 :   0 - 0x0
      13'h1A0A: dout <= 8'b00000000; // 6666 :   0 - 0x0
      13'h1A0B: dout <= 8'b00000000; // 6667 :   0 - 0x0
      13'h1A0C: dout <= 8'b00000000; // 6668 :   0 - 0x0
      13'h1A0D: dout <= 8'b00000000; // 6669 :   0 - 0x0
      13'h1A0E: dout <= 8'b00000000; // 6670 :   0 - 0x0
      13'h1A0F: dout <= 8'b00000000; // 6671 :   0 - 0x0
      13'h1A10: dout <= 8'b00000000; // 6672 :   0 - 0x0 -- Background 0xa1
      13'h1A11: dout <= 8'b00000000; // 6673 :   0 - 0x0
      13'h1A12: dout <= 8'b11100000; // 6674 : 224 - 0xe0
      13'h1A13: dout <= 8'b10000000; // 6675 : 128 - 0x80
      13'h1A14: dout <= 8'b01000000; // 6676 :  64 - 0x40
      13'h1A15: dout <= 8'b11110000; // 6677 : 240 - 0xf0
      13'h1A16: dout <= 8'b10011000; // 6678 : 152 - 0x98
      13'h1A17: dout <= 8'b11111000; // 6679 : 248 - 0xf8
      13'h1A18: dout <= 8'b00000000; // 6680 :   0 - 0x0
      13'h1A19: dout <= 8'b00000000; // 6681 :   0 - 0x0
      13'h1A1A: dout <= 8'b00000000; // 6682 :   0 - 0x0
      13'h1A1B: dout <= 8'b00000000; // 6683 :   0 - 0x0
      13'h1A1C: dout <= 8'b00000000; // 6684 :   0 - 0x0
      13'h1A1D: dout <= 8'b00000000; // 6685 :   0 - 0x0
      13'h1A1E: dout <= 8'b00000000; // 6686 :   0 - 0x0
      13'h1A1F: dout <= 8'b00000000; // 6687 :   0 - 0x0
      13'h1A20: dout <= 8'b00011111; // 6688 :  31 - 0x1f -- Background 0xa2
      13'h1A21: dout <= 8'b00010011; // 6689 :  19 - 0x13
      13'h1A22: dout <= 8'b00011111; // 6690 :  31 - 0x1f
      13'h1A23: dout <= 8'b00001111; // 6691 :  15 - 0xf
      13'h1A24: dout <= 8'b00001001; // 6692 :   9 - 0x9
      13'h1A25: dout <= 8'b00000111; // 6693 :   7 - 0x7
      13'h1A26: dout <= 8'b00000001; // 6694 :   1 - 0x1
      13'h1A27: dout <= 8'b00000000; // 6695 :   0 - 0x0
      13'h1A28: dout <= 8'b00000000; // 6696 :   0 - 0x0
      13'h1A29: dout <= 8'b00000000; // 6697 :   0 - 0x0
      13'h1A2A: dout <= 8'b00000000; // 6698 :   0 - 0x0
      13'h1A2B: dout <= 8'b00000000; // 6699 :   0 - 0x0
      13'h1A2C: dout <= 8'b00000000; // 6700 :   0 - 0x0
      13'h1A2D: dout <= 8'b00000000; // 6701 :   0 - 0x0
      13'h1A2E: dout <= 8'b00000000; // 6702 :   0 - 0x0
      13'h1A2F: dout <= 8'b00000000; // 6703 :   0 - 0x0
      13'h1A30: dout <= 8'b11100100; // 6704 : 228 - 0xe4 -- Background 0xa3
      13'h1A31: dout <= 8'b00111100; // 6705 :  60 - 0x3c
      13'h1A32: dout <= 8'b11100100; // 6706 : 228 - 0xe4
      13'h1A33: dout <= 8'b00111000; // 6707 :  56 - 0x38
      13'h1A34: dout <= 8'b11111000; // 6708 : 248 - 0xf8
      13'h1A35: dout <= 8'b11110000; // 6709 : 240 - 0xf0
      13'h1A36: dout <= 8'b11000000; // 6710 : 192 - 0xc0
      13'h1A37: dout <= 8'b00000000; // 6711 :   0 - 0x0
      13'h1A38: dout <= 8'b00000000; // 6712 :   0 - 0x0
      13'h1A39: dout <= 8'b00000000; // 6713 :   0 - 0x0
      13'h1A3A: dout <= 8'b00000000; // 6714 :   0 - 0x0
      13'h1A3B: dout <= 8'b00000000; // 6715 :   0 - 0x0
      13'h1A3C: dout <= 8'b00000000; // 6716 :   0 - 0x0
      13'h1A3D: dout <= 8'b00000000; // 6717 :   0 - 0x0
      13'h1A3E: dout <= 8'b00000000; // 6718 :   0 - 0x0
      13'h1A3F: dout <= 8'b00000000; // 6719 :   0 - 0x0
      13'h1A40: dout <= 8'b00000000; // 6720 :   0 - 0x0 -- Background 0xa4
      13'h1A41: dout <= 8'b00000000; // 6721 :   0 - 0x0
      13'h1A42: dout <= 8'b00000000; // 6722 :   0 - 0x0
      13'h1A43: dout <= 8'b00000000; // 6723 :   0 - 0x0
      13'h1A44: dout <= 8'b00010001; // 6724 :  17 - 0x11
      13'h1A45: dout <= 8'b00010011; // 6725 :  19 - 0x13
      13'h1A46: dout <= 8'b00011111; // 6726 :  31 - 0x1f
      13'h1A47: dout <= 8'b00011111; // 6727 :  31 - 0x1f
      13'h1A48: dout <= 8'b00000000; // 6728 :   0 - 0x0
      13'h1A49: dout <= 8'b00000000; // 6729 :   0 - 0x0
      13'h1A4A: dout <= 8'b00000000; // 6730 :   0 - 0x0
      13'h1A4B: dout <= 8'b00000000; // 6731 :   0 - 0x0
      13'h1A4C: dout <= 8'b00000000; // 6732 :   0 - 0x0
      13'h1A4D: dout <= 8'b00000000; // 6733 :   0 - 0x0
      13'h1A4E: dout <= 8'b00000000; // 6734 :   0 - 0x0
      13'h1A4F: dout <= 8'b00000000; // 6735 :   0 - 0x0
      13'h1A50: dout <= 8'b00000000; // 6736 :   0 - 0x0 -- Background 0xa5
      13'h1A51: dout <= 8'b00000000; // 6737 :   0 - 0x0
      13'h1A52: dout <= 8'b00000000; // 6738 :   0 - 0x0
      13'h1A53: dout <= 8'b10000000; // 6739 : 128 - 0x80
      13'h1A54: dout <= 8'b11000100; // 6740 : 196 - 0xc4
      13'h1A55: dout <= 8'b11100100; // 6741 : 228 - 0xe4
      13'h1A56: dout <= 8'b11111100; // 6742 : 252 - 0xfc
      13'h1A57: dout <= 8'b11111100; // 6743 : 252 - 0xfc
      13'h1A58: dout <= 8'b00000000; // 6744 :   0 - 0x0
      13'h1A59: dout <= 8'b00000000; // 6745 :   0 - 0x0
      13'h1A5A: dout <= 8'b00000000; // 6746 :   0 - 0x0
      13'h1A5B: dout <= 8'b00000000; // 6747 :   0 - 0x0
      13'h1A5C: dout <= 8'b00000000; // 6748 :   0 - 0x0
      13'h1A5D: dout <= 8'b00000000; // 6749 :   0 - 0x0
      13'h1A5E: dout <= 8'b00000000; // 6750 :   0 - 0x0
      13'h1A5F: dout <= 8'b00000000; // 6751 :   0 - 0x0
      13'h1A60: dout <= 8'b00011111; // 6752 :  31 - 0x1f -- Background 0xa6
      13'h1A61: dout <= 8'b00001110; // 6753 :  14 - 0xe
      13'h1A62: dout <= 8'b00000110; // 6754 :   6 - 0x6
      13'h1A63: dout <= 8'b00000010; // 6755 :   2 - 0x2
      13'h1A64: dout <= 8'b00000000; // 6756 :   0 - 0x0
      13'h1A65: dout <= 8'b00000000; // 6757 :   0 - 0x0
      13'h1A66: dout <= 8'b00000000; // 6758 :   0 - 0x0
      13'h1A67: dout <= 8'b00000000; // 6759 :   0 - 0x0
      13'h1A68: dout <= 8'b00000000; // 6760 :   0 - 0x0
      13'h1A69: dout <= 8'b00000000; // 6761 :   0 - 0x0
      13'h1A6A: dout <= 8'b00000000; // 6762 :   0 - 0x0
      13'h1A6B: dout <= 8'b00000000; // 6763 :   0 - 0x0
      13'h1A6C: dout <= 8'b00000000; // 6764 :   0 - 0x0
      13'h1A6D: dout <= 8'b00000000; // 6765 :   0 - 0x0
      13'h1A6E: dout <= 8'b00000000; // 6766 :   0 - 0x0
      13'h1A6F: dout <= 8'b00000000; // 6767 :   0 - 0x0
      13'h1A70: dout <= 8'b11111100; // 6768 : 252 - 0xfc -- Background 0xa7
      13'h1A71: dout <= 8'b10111000; // 6769 : 184 - 0xb8
      13'h1A72: dout <= 8'b10110000; // 6770 : 176 - 0xb0
      13'h1A73: dout <= 8'b10100000; // 6771 : 160 - 0xa0
      13'h1A74: dout <= 8'b10000000; // 6772 : 128 - 0x80
      13'h1A75: dout <= 8'b00000000; // 6773 :   0 - 0x0
      13'h1A76: dout <= 8'b00000000; // 6774 :   0 - 0x0
      13'h1A77: dout <= 8'b00000000; // 6775 :   0 - 0x0
      13'h1A78: dout <= 8'b00000000; // 6776 :   0 - 0x0
      13'h1A79: dout <= 8'b00000000; // 6777 :   0 - 0x0
      13'h1A7A: dout <= 8'b00000000; // 6778 :   0 - 0x0
      13'h1A7B: dout <= 8'b00000000; // 6779 :   0 - 0x0
      13'h1A7C: dout <= 8'b00000000; // 6780 :   0 - 0x0
      13'h1A7D: dout <= 8'b00000000; // 6781 :   0 - 0x0
      13'h1A7E: dout <= 8'b00000000; // 6782 :   0 - 0x0
      13'h1A7F: dout <= 8'b00000000; // 6783 :   0 - 0x0
      13'h1A80: dout <= 8'b00000000; // 6784 :   0 - 0x0 -- Background 0xa8
      13'h1A81: dout <= 8'b00000000; // 6785 :   0 - 0x0
      13'h1A82: dout <= 8'b00000000; // 6786 :   0 - 0x0
      13'h1A83: dout <= 8'b00000001; // 6787 :   1 - 0x1
      13'h1A84: dout <= 8'b00000011; // 6788 :   3 - 0x3
      13'h1A85: dout <= 8'b00000110; // 6789 :   6 - 0x6
      13'h1A86: dout <= 8'b00000110; // 6790 :   6 - 0x6
      13'h1A87: dout <= 8'b00001111; // 6791 :  15 - 0xf
      13'h1A88: dout <= 8'b00000000; // 6792 :   0 - 0x0
      13'h1A89: dout <= 8'b00000000; // 6793 :   0 - 0x0
      13'h1A8A: dout <= 8'b00000000; // 6794 :   0 - 0x0
      13'h1A8B: dout <= 8'b00000000; // 6795 :   0 - 0x0
      13'h1A8C: dout <= 8'b00000000; // 6796 :   0 - 0x0
      13'h1A8D: dout <= 8'b00000000; // 6797 :   0 - 0x0
      13'h1A8E: dout <= 8'b00000000; // 6798 :   0 - 0x0
      13'h1A8F: dout <= 8'b00000000; // 6799 :   0 - 0x0
      13'h1A90: dout <= 8'b00000000; // 6800 :   0 - 0x0 -- Background 0xa9
      13'h1A91: dout <= 8'b00011000; // 6801 :  24 - 0x18
      13'h1A92: dout <= 8'b11110100; // 6802 : 244 - 0xf4
      13'h1A93: dout <= 8'b11111000; // 6803 : 248 - 0xf8
      13'h1A94: dout <= 8'b00111000; // 6804 :  56 - 0x38
      13'h1A95: dout <= 8'b01111100; // 6805 : 124 - 0x7c
      13'h1A96: dout <= 8'b11111100; // 6806 : 252 - 0xfc
      13'h1A97: dout <= 8'b11111100; // 6807 : 252 - 0xfc
      13'h1A98: dout <= 8'b00000000; // 6808 :   0 - 0x0
      13'h1A99: dout <= 8'b00000000; // 6809 :   0 - 0x0
      13'h1A9A: dout <= 8'b00000000; // 6810 :   0 - 0x0
      13'h1A9B: dout <= 8'b00000000; // 6811 :   0 - 0x0
      13'h1A9C: dout <= 8'b00000000; // 6812 :   0 - 0x0
      13'h1A9D: dout <= 8'b00000000; // 6813 :   0 - 0x0
      13'h1A9E: dout <= 8'b00000000; // 6814 :   0 - 0x0
      13'h1A9F: dout <= 8'b00000000; // 6815 :   0 - 0x0
      13'h1AA0: dout <= 8'b00001111; // 6816 :  15 - 0xf -- Background 0xaa
      13'h1AA1: dout <= 8'b00011111; // 6817 :  31 - 0x1f
      13'h1AA2: dout <= 8'b00110000; // 6818 :  48 - 0x30
      13'h1AA3: dout <= 8'b00111000; // 6819 :  56 - 0x38
      13'h1AA4: dout <= 8'b00011101; // 6820 :  29 - 0x1d
      13'h1AA5: dout <= 8'b00000011; // 6821 :   3 - 0x3
      13'h1AA6: dout <= 8'b00000011; // 6822 :   3 - 0x3
      13'h1AA7: dout <= 8'b00000000; // 6823 :   0 - 0x0
      13'h1AA8: dout <= 8'b00000000; // 6824 :   0 - 0x0
      13'h1AA9: dout <= 8'b00000000; // 6825 :   0 - 0x0
      13'h1AAA: dout <= 8'b00000000; // 6826 :   0 - 0x0
      13'h1AAB: dout <= 8'b00000000; // 6827 :   0 - 0x0
      13'h1AAC: dout <= 8'b00000000; // 6828 :   0 - 0x0
      13'h1AAD: dout <= 8'b00000000; // 6829 :   0 - 0x0
      13'h1AAE: dout <= 8'b00000000; // 6830 :   0 - 0x0
      13'h1AAF: dout <= 8'b00000000; // 6831 :   0 - 0x0
      13'h1AB0: dout <= 8'b11111100; // 6832 : 252 - 0xfc -- Background 0xab
      13'h1AB1: dout <= 8'b11111100; // 6833 : 252 - 0xfc
      13'h1AB2: dout <= 8'b01111100; // 6834 : 124 - 0x7c
      13'h1AB3: dout <= 8'b10001110; // 6835 : 142 - 0x8e
      13'h1AB4: dout <= 8'b10000110; // 6836 : 134 - 0x86
      13'h1AB5: dout <= 8'b10011100; // 6837 : 156 - 0x9c
      13'h1AB6: dout <= 8'b01111000; // 6838 : 120 - 0x78
      13'h1AB7: dout <= 8'b00000000; // 6839 :   0 - 0x0
      13'h1AB8: dout <= 8'b00000000; // 6840 :   0 - 0x0
      13'h1AB9: dout <= 8'b00000000; // 6841 :   0 - 0x0
      13'h1ABA: dout <= 8'b00000000; // 6842 :   0 - 0x0
      13'h1ABB: dout <= 8'b00000000; // 6843 :   0 - 0x0
      13'h1ABC: dout <= 8'b00000000; // 6844 :   0 - 0x0
      13'h1ABD: dout <= 8'b00000000; // 6845 :   0 - 0x0
      13'h1ABE: dout <= 8'b00000000; // 6846 :   0 - 0x0
      13'h1ABF: dout <= 8'b00000000; // 6847 :   0 - 0x0
      13'h1AC0: dout <= 8'b00000000; // 6848 :   0 - 0x0 -- Background 0xac
      13'h1AC1: dout <= 8'b00000001; // 6849 :   1 - 0x1
      13'h1AC2: dout <= 8'b00000110; // 6850 :   6 - 0x6
      13'h1AC3: dout <= 8'b00000111; // 6851 :   7 - 0x7
      13'h1AC4: dout <= 8'b00000111; // 6852 :   7 - 0x7
      13'h1AC5: dout <= 8'b00000111; // 6853 :   7 - 0x7
      13'h1AC6: dout <= 8'b00000001; // 6854 :   1 - 0x1
      13'h1AC7: dout <= 8'b00000011; // 6855 :   3 - 0x3
      13'h1AC8: dout <= 8'b00000000; // 6856 :   0 - 0x0
      13'h1AC9: dout <= 8'b00000000; // 6857 :   0 - 0x0
      13'h1ACA: dout <= 8'b00000000; // 6858 :   0 - 0x0
      13'h1ACB: dout <= 8'b00000000; // 6859 :   0 - 0x0
      13'h1ACC: dout <= 8'b00000000; // 6860 :   0 - 0x0
      13'h1ACD: dout <= 8'b00000000; // 6861 :   0 - 0x0
      13'h1ACE: dout <= 8'b00000000; // 6862 :   0 - 0x0
      13'h1ACF: dout <= 8'b00000000; // 6863 :   0 - 0x0
      13'h1AD0: dout <= 8'b00000000; // 6864 :   0 - 0x0 -- Background 0xad
      13'h1AD1: dout <= 8'b11000000; // 6865 : 192 - 0xc0
      13'h1AD2: dout <= 8'b00110000; // 6866 :  48 - 0x30
      13'h1AD3: dout <= 8'b11110000; // 6867 : 240 - 0xf0
      13'h1AD4: dout <= 8'b11110000; // 6868 : 240 - 0xf0
      13'h1AD5: dout <= 8'b11110000; // 6869 : 240 - 0xf0
      13'h1AD6: dout <= 8'b01000000; // 6870 :  64 - 0x40
      13'h1AD7: dout <= 8'b01000000; // 6871 :  64 - 0x40
      13'h1AD8: dout <= 8'b00000000; // 6872 :   0 - 0x0
      13'h1AD9: dout <= 8'b00000000; // 6873 :   0 - 0x0
      13'h1ADA: dout <= 8'b00000000; // 6874 :   0 - 0x0
      13'h1ADB: dout <= 8'b00000000; // 6875 :   0 - 0x0
      13'h1ADC: dout <= 8'b00000000; // 6876 :   0 - 0x0
      13'h1ADD: dout <= 8'b00000000; // 6877 :   0 - 0x0
      13'h1ADE: dout <= 8'b00000000; // 6878 :   0 - 0x0
      13'h1ADF: dout <= 8'b00000000; // 6879 :   0 - 0x0
      13'h1AE0: dout <= 8'b00000001; // 6880 :   1 - 0x1 -- Background 0xae
      13'h1AE1: dout <= 8'b00000000; // 6881 :   0 - 0x0
      13'h1AE2: dout <= 8'b00000001; // 6882 :   1 - 0x1
      13'h1AE3: dout <= 8'b00000011; // 6883 :   3 - 0x3
      13'h1AE4: dout <= 8'b00000001; // 6884 :   1 - 0x1
      13'h1AE5: dout <= 8'b00000000; // 6885 :   0 - 0x0
      13'h1AE6: dout <= 8'b00000000; // 6886 :   0 - 0x0
      13'h1AE7: dout <= 8'b00000000; // 6887 :   0 - 0x0
      13'h1AE8: dout <= 8'b00000000; // 6888 :   0 - 0x0
      13'h1AE9: dout <= 8'b00000000; // 6889 :   0 - 0x0
      13'h1AEA: dout <= 8'b00000000; // 6890 :   0 - 0x0
      13'h1AEB: dout <= 8'b00000000; // 6891 :   0 - 0x0
      13'h1AEC: dout <= 8'b00000000; // 6892 :   0 - 0x0
      13'h1AED: dout <= 8'b00000000; // 6893 :   0 - 0x0
      13'h1AEE: dout <= 8'b00000000; // 6894 :   0 - 0x0
      13'h1AEF: dout <= 8'b00000000; // 6895 :   0 - 0x0
      13'h1AF0: dout <= 8'b01000000; // 6896 :  64 - 0x40 -- Background 0xaf
      13'h1AF1: dout <= 8'b01000000; // 6897 :  64 - 0x40
      13'h1AF2: dout <= 8'b01000000; // 6898 :  64 - 0x40
      13'h1AF3: dout <= 8'b01000000; // 6899 :  64 - 0x40
      13'h1AF4: dout <= 8'b01000000; // 6900 :  64 - 0x40
      13'h1AF5: dout <= 8'b10000000; // 6901 : 128 - 0x80
      13'h1AF6: dout <= 8'b00000000; // 6902 :   0 - 0x0
      13'h1AF7: dout <= 8'b00000000; // 6903 :   0 - 0x0
      13'h1AF8: dout <= 8'b00000000; // 6904 :   0 - 0x0
      13'h1AF9: dout <= 8'b00000000; // 6905 :   0 - 0x0
      13'h1AFA: dout <= 8'b00000000; // 6906 :   0 - 0x0
      13'h1AFB: dout <= 8'b00000000; // 6907 :   0 - 0x0
      13'h1AFC: dout <= 8'b00000000; // 6908 :   0 - 0x0
      13'h1AFD: dout <= 8'b00000000; // 6909 :   0 - 0x0
      13'h1AFE: dout <= 8'b00000000; // 6910 :   0 - 0x0
      13'h1AFF: dout <= 8'b00000000; // 6911 :   0 - 0x0
      13'h1B00: dout <= 8'b01111110; // 6912 : 126 - 0x7e -- Background 0xb0
      13'h1B01: dout <= 8'b01100011; // 6913 :  99 - 0x63
      13'h1B02: dout <= 8'b01100011; // 6914 :  99 - 0x63
      13'h1B03: dout <= 8'b01100011; // 6915 :  99 - 0x63
      13'h1B04: dout <= 8'b01111110; // 6916 : 126 - 0x7e
      13'h1B05: dout <= 8'b01100000; // 6917 :  96 - 0x60
      13'h1B06: dout <= 8'b01100000; // 6918 :  96 - 0x60
      13'h1B07: dout <= 8'b00000000; // 6919 :   0 - 0x0
      13'h1B08: dout <= 8'b01111110; // 6920 : 126 - 0x7e
      13'h1B09: dout <= 8'b01100011; // 6921 :  99 - 0x63
      13'h1B0A: dout <= 8'b01100011; // 6922 :  99 - 0x63
      13'h1B0B: dout <= 8'b01100011; // 6923 :  99 - 0x63
      13'h1B0C: dout <= 8'b01111110; // 6924 : 126 - 0x7e
      13'h1B0D: dout <= 8'b01100000; // 6925 :  96 - 0x60
      13'h1B0E: dout <= 8'b01100000; // 6926 :  96 - 0x60
      13'h1B0F: dout <= 8'b00000000; // 6927 :   0 - 0x0
      13'h1B10: dout <= 8'b01100000; // 6928 :  96 - 0x60 -- Background 0xb1
      13'h1B11: dout <= 8'b01100000; // 6929 :  96 - 0x60
      13'h1B12: dout <= 8'b01100000; // 6930 :  96 - 0x60
      13'h1B13: dout <= 8'b01100000; // 6931 :  96 - 0x60
      13'h1B14: dout <= 8'b01100000; // 6932 :  96 - 0x60
      13'h1B15: dout <= 8'b01100000; // 6933 :  96 - 0x60
      13'h1B16: dout <= 8'b01111111; // 6934 : 127 - 0x7f
      13'h1B17: dout <= 8'b00000000; // 6935 :   0 - 0x0
      13'h1B18: dout <= 8'b01100000; // 6936 :  96 - 0x60
      13'h1B19: dout <= 8'b01100000; // 6937 :  96 - 0x60
      13'h1B1A: dout <= 8'b01100000; // 6938 :  96 - 0x60
      13'h1B1B: dout <= 8'b01100000; // 6939 :  96 - 0x60
      13'h1B1C: dout <= 8'b01100000; // 6940 :  96 - 0x60
      13'h1B1D: dout <= 8'b01100000; // 6941 :  96 - 0x60
      13'h1B1E: dout <= 8'b01111111; // 6942 : 127 - 0x7f
      13'h1B1F: dout <= 8'b00000000; // 6943 :   0 - 0x0
      13'h1B20: dout <= 8'b00011100; // 6944 :  28 - 0x1c -- Background 0xb2
      13'h1B21: dout <= 8'b00110110; // 6945 :  54 - 0x36
      13'h1B22: dout <= 8'b01100011; // 6946 :  99 - 0x63
      13'h1B23: dout <= 8'b01100011; // 6947 :  99 - 0x63
      13'h1B24: dout <= 8'b01111111; // 6948 : 127 - 0x7f
      13'h1B25: dout <= 8'b01100011; // 6949 :  99 - 0x63
      13'h1B26: dout <= 8'b01100011; // 6950 :  99 - 0x63
      13'h1B27: dout <= 8'b00000000; // 6951 :   0 - 0x0
      13'h1B28: dout <= 8'b00011100; // 6952 :  28 - 0x1c
      13'h1B29: dout <= 8'b00110110; // 6953 :  54 - 0x36
      13'h1B2A: dout <= 8'b01100011; // 6954 :  99 - 0x63
      13'h1B2B: dout <= 8'b01100011; // 6955 :  99 - 0x63
      13'h1B2C: dout <= 8'b01111111; // 6956 : 127 - 0x7f
      13'h1B2D: dout <= 8'b01100011; // 6957 :  99 - 0x63
      13'h1B2E: dout <= 8'b01100011; // 6958 :  99 - 0x63
      13'h1B2F: dout <= 8'b00000000; // 6959 :   0 - 0x0
      13'h1B30: dout <= 8'b00110011; // 6960 :  51 - 0x33 -- Background 0xb3
      13'h1B31: dout <= 8'b00110011; // 6961 :  51 - 0x33
      13'h1B32: dout <= 8'b00110011; // 6962 :  51 - 0x33
      13'h1B33: dout <= 8'b00011110; // 6963 :  30 - 0x1e
      13'h1B34: dout <= 8'b00001100; // 6964 :  12 - 0xc
      13'h1B35: dout <= 8'b00001100; // 6965 :  12 - 0xc
      13'h1B36: dout <= 8'b00001100; // 6966 :  12 - 0xc
      13'h1B37: dout <= 8'b00000000; // 6967 :   0 - 0x0
      13'h1B38: dout <= 8'b00110011; // 6968 :  51 - 0x33
      13'h1B39: dout <= 8'b00110011; // 6969 :  51 - 0x33
      13'h1B3A: dout <= 8'b00110011; // 6970 :  51 - 0x33
      13'h1B3B: dout <= 8'b00011110; // 6971 :  30 - 0x1e
      13'h1B3C: dout <= 8'b00001100; // 6972 :  12 - 0xc
      13'h1B3D: dout <= 8'b00001100; // 6973 :  12 - 0xc
      13'h1B3E: dout <= 8'b00001100; // 6974 :  12 - 0xc
      13'h1B3F: dout <= 8'b00000000; // 6975 :   0 - 0x0
      13'h1B40: dout <= 8'b01111111; // 6976 : 127 - 0x7f -- Background 0xb4
      13'h1B41: dout <= 8'b01100000; // 6977 :  96 - 0x60
      13'h1B42: dout <= 8'b01100000; // 6978 :  96 - 0x60
      13'h1B43: dout <= 8'b01111110; // 6979 : 126 - 0x7e
      13'h1B44: dout <= 8'b01100000; // 6980 :  96 - 0x60
      13'h1B45: dout <= 8'b01100000; // 6981 :  96 - 0x60
      13'h1B46: dout <= 8'b01111111; // 6982 : 127 - 0x7f
      13'h1B47: dout <= 8'b00000000; // 6983 :   0 - 0x0
      13'h1B48: dout <= 8'b01111111; // 6984 : 127 - 0x7f
      13'h1B49: dout <= 8'b01100000; // 6985 :  96 - 0x60
      13'h1B4A: dout <= 8'b01100000; // 6986 :  96 - 0x60
      13'h1B4B: dout <= 8'b01111110; // 6987 : 126 - 0x7e
      13'h1B4C: dout <= 8'b01100000; // 6988 :  96 - 0x60
      13'h1B4D: dout <= 8'b01100000; // 6989 :  96 - 0x60
      13'h1B4E: dout <= 8'b01111111; // 6990 : 127 - 0x7f
      13'h1B4F: dout <= 8'b00000000; // 6991 :   0 - 0x0
      13'h1B50: dout <= 8'b01111110; // 6992 : 126 - 0x7e -- Background 0xb5
      13'h1B51: dout <= 8'b01100011; // 6993 :  99 - 0x63
      13'h1B52: dout <= 8'b01100011; // 6994 :  99 - 0x63
      13'h1B53: dout <= 8'b01100111; // 6995 : 103 - 0x67
      13'h1B54: dout <= 8'b01111100; // 6996 : 124 - 0x7c
      13'h1B55: dout <= 8'b01101110; // 6997 : 110 - 0x6e
      13'h1B56: dout <= 8'b01100111; // 6998 : 103 - 0x67
      13'h1B57: dout <= 8'b00000000; // 6999 :   0 - 0x0
      13'h1B58: dout <= 8'b01111110; // 7000 : 126 - 0x7e
      13'h1B59: dout <= 8'b01100011; // 7001 :  99 - 0x63
      13'h1B5A: dout <= 8'b01100011; // 7002 :  99 - 0x63
      13'h1B5B: dout <= 8'b01100111; // 7003 : 103 - 0x67
      13'h1B5C: dout <= 8'b01111100; // 7004 : 124 - 0x7c
      13'h1B5D: dout <= 8'b01101110; // 7005 : 110 - 0x6e
      13'h1B5E: dout <= 8'b01100111; // 7006 : 103 - 0x67
      13'h1B5F: dout <= 8'b00000000; // 7007 :   0 - 0x0
      13'h1B60: dout <= 8'b00111110; // 7008 :  62 - 0x3e -- Background 0xb6
      13'h1B61: dout <= 8'b01100011; // 7009 :  99 - 0x63
      13'h1B62: dout <= 8'b01100011; // 7010 :  99 - 0x63
      13'h1B63: dout <= 8'b01100011; // 7011 :  99 - 0x63
      13'h1B64: dout <= 8'b01100011; // 7012 :  99 - 0x63
      13'h1B65: dout <= 8'b01100011; // 7013 :  99 - 0x63
      13'h1B66: dout <= 8'b00111110; // 7014 :  62 - 0x3e
      13'h1B67: dout <= 8'b00000000; // 7015 :   0 - 0x0
      13'h1B68: dout <= 8'b00111110; // 7016 :  62 - 0x3e
      13'h1B69: dout <= 8'b01100011; // 7017 :  99 - 0x63
      13'h1B6A: dout <= 8'b01100011; // 7018 :  99 - 0x63
      13'h1B6B: dout <= 8'b01100011; // 7019 :  99 - 0x63
      13'h1B6C: dout <= 8'b01100011; // 7020 :  99 - 0x63
      13'h1B6D: dout <= 8'b01100011; // 7021 :  99 - 0x63
      13'h1B6E: dout <= 8'b00111110; // 7022 :  62 - 0x3e
      13'h1B6F: dout <= 8'b00000000; // 7023 :   0 - 0x0
      13'h1B70: dout <= 8'b01100011; // 7024 :  99 - 0x63 -- Background 0xb7
      13'h1B71: dout <= 8'b01110011; // 7025 : 115 - 0x73
      13'h1B72: dout <= 8'b01111011; // 7026 : 123 - 0x7b
      13'h1B73: dout <= 8'b01111111; // 7027 : 127 - 0x7f
      13'h1B74: dout <= 8'b01101111; // 7028 : 111 - 0x6f
      13'h1B75: dout <= 8'b01100111; // 7029 : 103 - 0x67
      13'h1B76: dout <= 8'b01100011; // 7030 :  99 - 0x63
      13'h1B77: dout <= 8'b00000000; // 7031 :   0 - 0x0
      13'h1B78: dout <= 8'b01100011; // 7032 :  99 - 0x63
      13'h1B79: dout <= 8'b01110011; // 7033 : 115 - 0x73
      13'h1B7A: dout <= 8'b01111011; // 7034 : 123 - 0x7b
      13'h1B7B: dout <= 8'b01111111; // 7035 : 127 - 0x7f
      13'h1B7C: dout <= 8'b01101111; // 7036 : 111 - 0x6f
      13'h1B7D: dout <= 8'b01100111; // 7037 : 103 - 0x67
      13'h1B7E: dout <= 8'b01100011; // 7038 :  99 - 0x63
      13'h1B7F: dout <= 8'b00000000; // 7039 :   0 - 0x0
      13'h1B80: dout <= 8'b00111111; // 7040 :  63 - 0x3f -- Background 0xb8
      13'h1B81: dout <= 8'b00001100; // 7041 :  12 - 0xc
      13'h1B82: dout <= 8'b00001100; // 7042 :  12 - 0xc
      13'h1B83: dout <= 8'b00001100; // 7043 :  12 - 0xc
      13'h1B84: dout <= 8'b00001100; // 7044 :  12 - 0xc
      13'h1B85: dout <= 8'b00001100; // 7045 :  12 - 0xc
      13'h1B86: dout <= 8'b00001100; // 7046 :  12 - 0xc
      13'h1B87: dout <= 8'b00000000; // 7047 :   0 - 0x0
      13'h1B88: dout <= 8'b00111111; // 7048 :  63 - 0x3f
      13'h1B89: dout <= 8'b00001100; // 7049 :  12 - 0xc
      13'h1B8A: dout <= 8'b00001100; // 7050 :  12 - 0xc
      13'h1B8B: dout <= 8'b00001100; // 7051 :  12 - 0xc
      13'h1B8C: dout <= 8'b00001100; // 7052 :  12 - 0xc
      13'h1B8D: dout <= 8'b00001100; // 7053 :  12 - 0xc
      13'h1B8E: dout <= 8'b00001100; // 7054 :  12 - 0xc
      13'h1B8F: dout <= 8'b00000000; // 7055 :   0 - 0x0
      13'h1B90: dout <= 8'b01100011; // 7056 :  99 - 0x63 -- Background 0xb9
      13'h1B91: dout <= 8'b01100011; // 7057 :  99 - 0x63
      13'h1B92: dout <= 8'b01101011; // 7058 : 107 - 0x6b
      13'h1B93: dout <= 8'b01111111; // 7059 : 127 - 0x7f
      13'h1B94: dout <= 8'b01111111; // 7060 : 127 - 0x7f
      13'h1B95: dout <= 8'b01110111; // 7061 : 119 - 0x77
      13'h1B96: dout <= 8'b01100011; // 7062 :  99 - 0x63
      13'h1B97: dout <= 8'b00000000; // 7063 :   0 - 0x0
      13'h1B98: dout <= 8'b01100011; // 7064 :  99 - 0x63
      13'h1B99: dout <= 8'b01100011; // 7065 :  99 - 0x63
      13'h1B9A: dout <= 8'b01101011; // 7066 : 107 - 0x6b
      13'h1B9B: dout <= 8'b01111111; // 7067 : 127 - 0x7f
      13'h1B9C: dout <= 8'b01111111; // 7068 : 127 - 0x7f
      13'h1B9D: dout <= 8'b01110111; // 7069 : 119 - 0x77
      13'h1B9E: dout <= 8'b01100011; // 7070 :  99 - 0x63
      13'h1B9F: dout <= 8'b00000000; // 7071 :   0 - 0x0
      13'h1BA0: dout <= 8'b01111100; // 7072 : 124 - 0x7c -- Background 0xba
      13'h1BA1: dout <= 8'b01100110; // 7073 : 102 - 0x66
      13'h1BA2: dout <= 8'b01100011; // 7074 :  99 - 0x63
      13'h1BA3: dout <= 8'b01100011; // 7075 :  99 - 0x63
      13'h1BA4: dout <= 8'b01100011; // 7076 :  99 - 0x63
      13'h1BA5: dout <= 8'b01100110; // 7077 : 102 - 0x66
      13'h1BA6: dout <= 8'b01111100; // 7078 : 124 - 0x7c
      13'h1BA7: dout <= 8'b00000000; // 7079 :   0 - 0x0
      13'h1BA8: dout <= 8'b00000000; // 7080 :   0 - 0x0
      13'h1BA9: dout <= 8'b00000000; // 7081 :   0 - 0x0
      13'h1BAA: dout <= 8'b00000000; // 7082 :   0 - 0x0
      13'h1BAB: dout <= 8'b00000000; // 7083 :   0 - 0x0
      13'h1BAC: dout <= 8'b00000000; // 7084 :   0 - 0x0
      13'h1BAD: dout <= 8'b00000000; // 7085 :   0 - 0x0
      13'h1BAE: dout <= 8'b00000000; // 7086 :   0 - 0x0
      13'h1BAF: dout <= 8'b00000000; // 7087 :   0 - 0x0
      13'h1BB0: dout <= 8'b00011100; // 7088 :  28 - 0x1c -- Background 0xbb
      13'h1BB1: dout <= 8'b00011100; // 7089 :  28 - 0x1c
      13'h1BB2: dout <= 8'b00011100; // 7090 :  28 - 0x1c
      13'h1BB3: dout <= 8'b00011000; // 7091 :  24 - 0x18
      13'h1BB4: dout <= 8'b00011000; // 7092 :  24 - 0x18
      13'h1BB5: dout <= 8'b00000000; // 7093 :   0 - 0x0
      13'h1BB6: dout <= 8'b00011000; // 7094 :  24 - 0x18
      13'h1BB7: dout <= 8'b00000000; // 7095 :   0 - 0x0
      13'h1BB8: dout <= 8'b00000000; // 7096 :   0 - 0x0
      13'h1BB9: dout <= 8'b00000000; // 7097 :   0 - 0x0
      13'h1BBA: dout <= 8'b00000000; // 7098 :   0 - 0x0
      13'h1BBB: dout <= 8'b00000000; // 7099 :   0 - 0x0
      13'h1BBC: dout <= 8'b00000000; // 7100 :   0 - 0x0
      13'h1BBD: dout <= 8'b00000000; // 7101 :   0 - 0x0
      13'h1BBE: dout <= 8'b00000000; // 7102 :   0 - 0x0
      13'h1BBF: dout <= 8'b00000000; // 7103 :   0 - 0x0
      13'h1BC0: dout <= 8'b00011111; // 7104 :  31 - 0x1f -- Background 0xbc
      13'h1BC1: dout <= 8'b00110000; // 7105 :  48 - 0x30
      13'h1BC2: dout <= 8'b01100000; // 7106 :  96 - 0x60
      13'h1BC3: dout <= 8'b01100111; // 7107 : 103 - 0x67
      13'h1BC4: dout <= 8'b01100011; // 7108 :  99 - 0x63
      13'h1BC5: dout <= 8'b00110011; // 7109 :  51 - 0x33
      13'h1BC6: dout <= 8'b00011111; // 7110 :  31 - 0x1f
      13'h1BC7: dout <= 8'b00000000; // 7111 :   0 - 0x0
      13'h1BC8: dout <= 8'b00011111; // 7112 :  31 - 0x1f
      13'h1BC9: dout <= 8'b00110000; // 7113 :  48 - 0x30
      13'h1BCA: dout <= 8'b01100000; // 7114 :  96 - 0x60
      13'h1BCB: dout <= 8'b01100111; // 7115 : 103 - 0x67
      13'h1BCC: dout <= 8'b01100011; // 7116 :  99 - 0x63
      13'h1BCD: dout <= 8'b00110011; // 7117 :  51 - 0x33
      13'h1BCE: dout <= 8'b00011111; // 7118 :  31 - 0x1f
      13'h1BCF: dout <= 8'b00000000; // 7119 :   0 - 0x0
      13'h1BD0: dout <= 8'b01100011; // 7120 :  99 - 0x63 -- Background 0xbd
      13'h1BD1: dout <= 8'b01110111; // 7121 : 119 - 0x77
      13'h1BD2: dout <= 8'b01111111; // 7122 : 127 - 0x7f
      13'h1BD3: dout <= 8'b01111111; // 7123 : 127 - 0x7f
      13'h1BD4: dout <= 8'b01101011; // 7124 : 107 - 0x6b
      13'h1BD5: dout <= 8'b01100011; // 7125 :  99 - 0x63
      13'h1BD6: dout <= 8'b01100011; // 7126 :  99 - 0x63
      13'h1BD7: dout <= 8'b00000000; // 7127 :   0 - 0x0
      13'h1BD8: dout <= 8'b01100011; // 7128 :  99 - 0x63
      13'h1BD9: dout <= 8'b01110111; // 7129 : 119 - 0x77
      13'h1BDA: dout <= 8'b01111111; // 7130 : 127 - 0x7f
      13'h1BDB: dout <= 8'b01111111; // 7131 : 127 - 0x7f
      13'h1BDC: dout <= 8'b01101011; // 7132 : 107 - 0x6b
      13'h1BDD: dout <= 8'b01100011; // 7133 :  99 - 0x63
      13'h1BDE: dout <= 8'b01100011; // 7134 :  99 - 0x63
      13'h1BDF: dout <= 8'b00000000; // 7135 :   0 - 0x0
      13'h1BE0: dout <= 8'b01100011; // 7136 :  99 - 0x63 -- Background 0xbe
      13'h1BE1: dout <= 8'b01100011; // 7137 :  99 - 0x63
      13'h1BE2: dout <= 8'b01100011; // 7138 :  99 - 0x63
      13'h1BE3: dout <= 8'b01110111; // 7139 : 119 - 0x77
      13'h1BE4: dout <= 8'b00111110; // 7140 :  62 - 0x3e
      13'h1BE5: dout <= 8'b00011100; // 7141 :  28 - 0x1c
      13'h1BE6: dout <= 8'b00001000; // 7142 :   8 - 0x8
      13'h1BE7: dout <= 8'b00000000; // 7143 :   0 - 0x0
      13'h1BE8: dout <= 8'b01100011; // 7144 :  99 - 0x63
      13'h1BE9: dout <= 8'b01100011; // 7145 :  99 - 0x63
      13'h1BEA: dout <= 8'b01100011; // 7146 :  99 - 0x63
      13'h1BEB: dout <= 8'b01110111; // 7147 : 119 - 0x77
      13'h1BEC: dout <= 8'b00111110; // 7148 :  62 - 0x3e
      13'h1BED: dout <= 8'b00011100; // 7149 :  28 - 0x1c
      13'h1BEE: dout <= 8'b00001000; // 7150 :   8 - 0x8
      13'h1BEF: dout <= 8'b00000000; // 7151 :   0 - 0x0
      13'h1BF0: dout <= 8'b00000000; // 7152 :   0 - 0x0 -- Background 0xbf
      13'h1BF1: dout <= 8'b00000000; // 7153 :   0 - 0x0
      13'h1BF2: dout <= 8'b00000000; // 7154 :   0 - 0x0
      13'h1BF3: dout <= 8'b00000000; // 7155 :   0 - 0x0
      13'h1BF4: dout <= 8'b00000000; // 7156 :   0 - 0x0
      13'h1BF5: dout <= 8'b00000000; // 7157 :   0 - 0x0
      13'h1BF6: dout <= 8'b00000000; // 7158 :   0 - 0x0
      13'h1BF7: dout <= 8'b00000000; // 7159 :   0 - 0x0
      13'h1BF8: dout <= 8'b00000000; // 7160 :   0 - 0x0
      13'h1BF9: dout <= 8'b00000000; // 7161 :   0 - 0x0
      13'h1BFA: dout <= 8'b00000000; // 7162 :   0 - 0x0
      13'h1BFB: dout <= 8'b00000000; // 7163 :   0 - 0x0
      13'h1BFC: dout <= 8'b00000000; // 7164 :   0 - 0x0
      13'h1BFD: dout <= 8'b00000000; // 7165 :   0 - 0x0
      13'h1BFE: dout <= 8'b00000000; // 7166 :   0 - 0x0
      13'h1BFF: dout <= 8'b00000000; // 7167 :   0 - 0x0
      13'h1C00: dout <= 8'b00011111; // 7168 :  31 - 0x1f -- Background 0xc0
      13'h1C01: dout <= 8'b00110000; // 7169 :  48 - 0x30
      13'h1C02: dout <= 8'b01100000; // 7170 :  96 - 0x60
      13'h1C03: dout <= 8'b01100111; // 7171 : 103 - 0x67
      13'h1C04: dout <= 8'b01100011; // 7172 :  99 - 0x63
      13'h1C05: dout <= 8'b00110011; // 7173 :  51 - 0x33
      13'h1C06: dout <= 8'b00011111; // 7174 :  31 - 0x1f
      13'h1C07: dout <= 8'b00000000; // 7175 :   0 - 0x0
      13'h1C08: dout <= 8'b00000000; // 7176 :   0 - 0x0
      13'h1C09: dout <= 8'b00000000; // 7177 :   0 - 0x0
      13'h1C0A: dout <= 8'b00000000; // 7178 :   0 - 0x0
      13'h1C0B: dout <= 8'b00000000; // 7179 :   0 - 0x0
      13'h1C0C: dout <= 8'b00000000; // 7180 :   0 - 0x0
      13'h1C0D: dout <= 8'b00000000; // 7181 :   0 - 0x0
      13'h1C0E: dout <= 8'b00000000; // 7182 :   0 - 0x0
      13'h1C0F: dout <= 8'b00000000; // 7183 :   0 - 0x0
      13'h1C10: dout <= 8'b00011100; // 7184 :  28 - 0x1c -- Background 0xc1
      13'h1C11: dout <= 8'b00110110; // 7185 :  54 - 0x36
      13'h1C12: dout <= 8'b01100011; // 7186 :  99 - 0x63
      13'h1C13: dout <= 8'b01100011; // 7187 :  99 - 0x63
      13'h1C14: dout <= 8'b01111111; // 7188 : 127 - 0x7f
      13'h1C15: dout <= 8'b01100011; // 7189 :  99 - 0x63
      13'h1C16: dout <= 8'b01100011; // 7190 :  99 - 0x63
      13'h1C17: dout <= 8'b00000000; // 7191 :   0 - 0x0
      13'h1C18: dout <= 8'b00000000; // 7192 :   0 - 0x0
      13'h1C19: dout <= 8'b00000000; // 7193 :   0 - 0x0
      13'h1C1A: dout <= 8'b00000000; // 7194 :   0 - 0x0
      13'h1C1B: dout <= 8'b00000000; // 7195 :   0 - 0x0
      13'h1C1C: dout <= 8'b00000000; // 7196 :   0 - 0x0
      13'h1C1D: dout <= 8'b00000000; // 7197 :   0 - 0x0
      13'h1C1E: dout <= 8'b00000000; // 7198 :   0 - 0x0
      13'h1C1F: dout <= 8'b00000000; // 7199 :   0 - 0x0
      13'h1C20: dout <= 8'b01100011; // 7200 :  99 - 0x63 -- Background 0xc2
      13'h1C21: dout <= 8'b01110111; // 7201 : 119 - 0x77
      13'h1C22: dout <= 8'b01111111; // 7202 : 127 - 0x7f
      13'h1C23: dout <= 8'b01111111; // 7203 : 127 - 0x7f
      13'h1C24: dout <= 8'b01101011; // 7204 : 107 - 0x6b
      13'h1C25: dout <= 8'b01100011; // 7205 :  99 - 0x63
      13'h1C26: dout <= 8'b01100011; // 7206 :  99 - 0x63
      13'h1C27: dout <= 8'b00000000; // 7207 :   0 - 0x0
      13'h1C28: dout <= 8'b00000000; // 7208 :   0 - 0x0
      13'h1C29: dout <= 8'b00000000; // 7209 :   0 - 0x0
      13'h1C2A: dout <= 8'b00000000; // 7210 :   0 - 0x0
      13'h1C2B: dout <= 8'b00000000; // 7211 :   0 - 0x0
      13'h1C2C: dout <= 8'b00000000; // 7212 :   0 - 0x0
      13'h1C2D: dout <= 8'b00000000; // 7213 :   0 - 0x0
      13'h1C2E: dout <= 8'b00000000; // 7214 :   0 - 0x0
      13'h1C2F: dout <= 8'b00000000; // 7215 :   0 - 0x0
      13'h1C30: dout <= 8'b01111111; // 7216 : 127 - 0x7f -- Background 0xc3
      13'h1C31: dout <= 8'b01100000; // 7217 :  96 - 0x60
      13'h1C32: dout <= 8'b01100000; // 7218 :  96 - 0x60
      13'h1C33: dout <= 8'b01111110; // 7219 : 126 - 0x7e
      13'h1C34: dout <= 8'b01100000; // 7220 :  96 - 0x60
      13'h1C35: dout <= 8'b01100000; // 7221 :  96 - 0x60
      13'h1C36: dout <= 8'b01111111; // 7222 : 127 - 0x7f
      13'h1C37: dout <= 8'b00000000; // 7223 :   0 - 0x0
      13'h1C38: dout <= 8'b00000000; // 7224 :   0 - 0x0
      13'h1C39: dout <= 8'b00000000; // 7225 :   0 - 0x0
      13'h1C3A: dout <= 8'b00000000; // 7226 :   0 - 0x0
      13'h1C3B: dout <= 8'b00000000; // 7227 :   0 - 0x0
      13'h1C3C: dout <= 8'b00000000; // 7228 :   0 - 0x0
      13'h1C3D: dout <= 8'b00000000; // 7229 :   0 - 0x0
      13'h1C3E: dout <= 8'b00000000; // 7230 :   0 - 0x0
      13'h1C3F: dout <= 8'b00000000; // 7231 :   0 - 0x0
      13'h1C40: dout <= 8'b00111110; // 7232 :  62 - 0x3e -- Background 0xc4
      13'h1C41: dout <= 8'b01100011; // 7233 :  99 - 0x63
      13'h1C42: dout <= 8'b01100011; // 7234 :  99 - 0x63
      13'h1C43: dout <= 8'b01100011; // 7235 :  99 - 0x63
      13'h1C44: dout <= 8'b01100011; // 7236 :  99 - 0x63
      13'h1C45: dout <= 8'b01100011; // 7237 :  99 - 0x63
      13'h1C46: dout <= 8'b00111110; // 7238 :  62 - 0x3e
      13'h1C47: dout <= 8'b00000000; // 7239 :   0 - 0x0
      13'h1C48: dout <= 8'b00000000; // 7240 :   0 - 0x0
      13'h1C49: dout <= 8'b00000000; // 7241 :   0 - 0x0
      13'h1C4A: dout <= 8'b00000000; // 7242 :   0 - 0x0
      13'h1C4B: dout <= 8'b00000000; // 7243 :   0 - 0x0
      13'h1C4C: dout <= 8'b00000000; // 7244 :   0 - 0x0
      13'h1C4D: dout <= 8'b00000000; // 7245 :   0 - 0x0
      13'h1C4E: dout <= 8'b00000000; // 7246 :   0 - 0x0
      13'h1C4F: dout <= 8'b00000000; // 7247 :   0 - 0x0
      13'h1C50: dout <= 8'b01100011; // 7248 :  99 - 0x63 -- Background 0xc5
      13'h1C51: dout <= 8'b01100011; // 7249 :  99 - 0x63
      13'h1C52: dout <= 8'b01100011; // 7250 :  99 - 0x63
      13'h1C53: dout <= 8'b01110111; // 7251 : 119 - 0x77
      13'h1C54: dout <= 8'b00111110; // 7252 :  62 - 0x3e
      13'h1C55: dout <= 8'b00011100; // 7253 :  28 - 0x1c
      13'h1C56: dout <= 8'b00001000; // 7254 :   8 - 0x8
      13'h1C57: dout <= 8'b00000000; // 7255 :   0 - 0x0
      13'h1C58: dout <= 8'b00000000; // 7256 :   0 - 0x0
      13'h1C59: dout <= 8'b00000000; // 7257 :   0 - 0x0
      13'h1C5A: dout <= 8'b00000000; // 7258 :   0 - 0x0
      13'h1C5B: dout <= 8'b00000000; // 7259 :   0 - 0x0
      13'h1C5C: dout <= 8'b00000000; // 7260 :   0 - 0x0
      13'h1C5D: dout <= 8'b00000000; // 7261 :   0 - 0x0
      13'h1C5E: dout <= 8'b00000000; // 7262 :   0 - 0x0
      13'h1C5F: dout <= 8'b00000000; // 7263 :   0 - 0x0
      13'h1C60: dout <= 8'b01111110; // 7264 : 126 - 0x7e -- Background 0xc6
      13'h1C61: dout <= 8'b01100011; // 7265 :  99 - 0x63
      13'h1C62: dout <= 8'b01100011; // 7266 :  99 - 0x63
      13'h1C63: dout <= 8'b01100111; // 7267 : 103 - 0x67
      13'h1C64: dout <= 8'b01111100; // 7268 : 124 - 0x7c
      13'h1C65: dout <= 8'b01101110; // 7269 : 110 - 0x6e
      13'h1C66: dout <= 8'b01100111; // 7270 : 103 - 0x67
      13'h1C67: dout <= 8'b00000000; // 7271 :   0 - 0x0
      13'h1C68: dout <= 8'b00000000; // 7272 :   0 - 0x0
      13'h1C69: dout <= 8'b00000000; // 7273 :   0 - 0x0
      13'h1C6A: dout <= 8'b00000000; // 7274 :   0 - 0x0
      13'h1C6B: dout <= 8'b00000000; // 7275 :   0 - 0x0
      13'h1C6C: dout <= 8'b00000000; // 7276 :   0 - 0x0
      13'h1C6D: dout <= 8'b00000000; // 7277 :   0 - 0x0
      13'h1C6E: dout <= 8'b00000000; // 7278 :   0 - 0x0
      13'h1C6F: dout <= 8'b00000000; // 7279 :   0 - 0x0
      13'h1C70: dout <= 8'b00110011; // 7280 :  51 - 0x33 -- Background 0xc7
      13'h1C71: dout <= 8'b00110011; // 7281 :  51 - 0x33
      13'h1C72: dout <= 8'b00110011; // 7282 :  51 - 0x33
      13'h1C73: dout <= 8'b00011110; // 7283 :  30 - 0x1e
      13'h1C74: dout <= 8'b00001100; // 7284 :  12 - 0xc
      13'h1C75: dout <= 8'b00001100; // 7285 :  12 - 0xc
      13'h1C76: dout <= 8'b00001100; // 7286 :  12 - 0xc
      13'h1C77: dout <= 8'b00000000; // 7287 :   0 - 0x0
      13'h1C78: dout <= 8'b00000000; // 7288 :   0 - 0x0
      13'h1C79: dout <= 8'b00000000; // 7289 :   0 - 0x0
      13'h1C7A: dout <= 8'b00000000; // 7290 :   0 - 0x0
      13'h1C7B: dout <= 8'b00000000; // 7291 :   0 - 0x0
      13'h1C7C: dout <= 8'b00000000; // 7292 :   0 - 0x0
      13'h1C7D: dout <= 8'b00000000; // 7293 :   0 - 0x0
      13'h1C7E: dout <= 8'b00000000; // 7294 :   0 - 0x0
      13'h1C7F: dout <= 8'b00000000; // 7295 :   0 - 0x0
      13'h1C80: dout <= 8'b00000000; // 7296 :   0 - 0x0 -- Background 0xc8
      13'h1C81: dout <= 8'b00000000; // 7297 :   0 - 0x0
      13'h1C82: dout <= 8'b00000000; // 7298 :   0 - 0x0
      13'h1C83: dout <= 8'b00000000; // 7299 :   0 - 0x0
      13'h1C84: dout <= 8'b00000000; // 7300 :   0 - 0x0
      13'h1C85: dout <= 8'b00000000; // 7301 :   0 - 0x0
      13'h1C86: dout <= 8'b00000000; // 7302 :   0 - 0x0
      13'h1C87: dout <= 8'b00000000; // 7303 :   0 - 0x0
      13'h1C88: dout <= 8'b00000000; // 7304 :   0 - 0x0
      13'h1C89: dout <= 8'b00000000; // 7305 :   0 - 0x0
      13'h1C8A: dout <= 8'b00000000; // 7306 :   0 - 0x0
      13'h1C8B: dout <= 8'b00000000; // 7307 :   0 - 0x0
      13'h1C8C: dout <= 8'b00000000; // 7308 :   0 - 0x0
      13'h1C8D: dout <= 8'b00000000; // 7309 :   0 - 0x0
      13'h1C8E: dout <= 8'b00000000; // 7310 :   0 - 0x0
      13'h1C8F: dout <= 8'b00000000; // 7311 :   0 - 0x0
      13'h1C90: dout <= 8'b00000000; // 7312 :   0 - 0x0 -- Background 0xc9
      13'h1C91: dout <= 8'b00000000; // 7313 :   0 - 0x0
      13'h1C92: dout <= 8'b00000000; // 7314 :   0 - 0x0
      13'h1C93: dout <= 8'b00000000; // 7315 :   0 - 0x0
      13'h1C94: dout <= 8'b00000000; // 7316 :   0 - 0x0
      13'h1C95: dout <= 8'b00000000; // 7317 :   0 - 0x0
      13'h1C96: dout <= 8'b00000000; // 7318 :   0 - 0x0
      13'h1C97: dout <= 8'b00000000; // 7319 :   0 - 0x0
      13'h1C98: dout <= 8'b00000000; // 7320 :   0 - 0x0
      13'h1C99: dout <= 8'b00000000; // 7321 :   0 - 0x0
      13'h1C9A: dout <= 8'b00000000; // 7322 :   0 - 0x0
      13'h1C9B: dout <= 8'b00000000; // 7323 :   0 - 0x0
      13'h1C9C: dout <= 8'b00000000; // 7324 :   0 - 0x0
      13'h1C9D: dout <= 8'b00000000; // 7325 :   0 - 0x0
      13'h1C9E: dout <= 8'b00000000; // 7326 :   0 - 0x0
      13'h1C9F: dout <= 8'b00000000; // 7327 :   0 - 0x0
      13'h1CA0: dout <= 8'b00000000; // 7328 :   0 - 0x0 -- Background 0xca
      13'h1CA1: dout <= 8'b00000000; // 7329 :   0 - 0x0
      13'h1CA2: dout <= 8'b00000000; // 7330 :   0 - 0x0
      13'h1CA3: dout <= 8'b00000000; // 7331 :   0 - 0x0
      13'h1CA4: dout <= 8'b00000000; // 7332 :   0 - 0x0
      13'h1CA5: dout <= 8'b00000000; // 7333 :   0 - 0x0
      13'h1CA6: dout <= 8'b00000000; // 7334 :   0 - 0x0
      13'h1CA7: dout <= 8'b00000000; // 7335 :   0 - 0x0
      13'h1CA8: dout <= 8'b00000000; // 7336 :   0 - 0x0
      13'h1CA9: dout <= 8'b00000000; // 7337 :   0 - 0x0
      13'h1CAA: dout <= 8'b00000000; // 7338 :   0 - 0x0
      13'h1CAB: dout <= 8'b00000000; // 7339 :   0 - 0x0
      13'h1CAC: dout <= 8'b00000000; // 7340 :   0 - 0x0
      13'h1CAD: dout <= 8'b00000000; // 7341 :   0 - 0x0
      13'h1CAE: dout <= 8'b00000000; // 7342 :   0 - 0x0
      13'h1CAF: dout <= 8'b00000000; // 7343 :   0 - 0x0
      13'h1CB0: dout <= 8'b00000000; // 7344 :   0 - 0x0 -- Background 0xcb
      13'h1CB1: dout <= 8'b00000000; // 7345 :   0 - 0x0
      13'h1CB2: dout <= 8'b00000000; // 7346 :   0 - 0x0
      13'h1CB3: dout <= 8'b00000000; // 7347 :   0 - 0x0
      13'h1CB4: dout <= 8'b00000000; // 7348 :   0 - 0x0
      13'h1CB5: dout <= 8'b00000000; // 7349 :   0 - 0x0
      13'h1CB6: dout <= 8'b00000000; // 7350 :   0 - 0x0
      13'h1CB7: dout <= 8'b00000000; // 7351 :   0 - 0x0
      13'h1CB8: dout <= 8'b00000000; // 7352 :   0 - 0x0
      13'h1CB9: dout <= 8'b00000000; // 7353 :   0 - 0x0
      13'h1CBA: dout <= 8'b00000000; // 7354 :   0 - 0x0
      13'h1CBB: dout <= 8'b00000000; // 7355 :   0 - 0x0
      13'h1CBC: dout <= 8'b00000000; // 7356 :   0 - 0x0
      13'h1CBD: dout <= 8'b00000000; // 7357 :   0 - 0x0
      13'h1CBE: dout <= 8'b00000000; // 7358 :   0 - 0x0
      13'h1CBF: dout <= 8'b00000000; // 7359 :   0 - 0x0
      13'h1CC0: dout <= 8'b00000000; // 7360 :   0 - 0x0 -- Background 0xcc
      13'h1CC1: dout <= 8'b00000000; // 7361 :   0 - 0x0
      13'h1CC2: dout <= 8'b00000000; // 7362 :   0 - 0x0
      13'h1CC3: dout <= 8'b00000000; // 7363 :   0 - 0x0
      13'h1CC4: dout <= 8'b00000000; // 7364 :   0 - 0x0
      13'h1CC5: dout <= 8'b00000000; // 7365 :   0 - 0x0
      13'h1CC6: dout <= 8'b00000000; // 7366 :   0 - 0x0
      13'h1CC7: dout <= 8'b00000000; // 7367 :   0 - 0x0
      13'h1CC8: dout <= 8'b00000000; // 7368 :   0 - 0x0
      13'h1CC9: dout <= 8'b00000000; // 7369 :   0 - 0x0
      13'h1CCA: dout <= 8'b00000000; // 7370 :   0 - 0x0
      13'h1CCB: dout <= 8'b00000000; // 7371 :   0 - 0x0
      13'h1CCC: dout <= 8'b00000000; // 7372 :   0 - 0x0
      13'h1CCD: dout <= 8'b00000000; // 7373 :   0 - 0x0
      13'h1CCE: dout <= 8'b00000000; // 7374 :   0 - 0x0
      13'h1CCF: dout <= 8'b00000000; // 7375 :   0 - 0x0
      13'h1CD0: dout <= 8'b00000000; // 7376 :   0 - 0x0 -- Background 0xcd
      13'h1CD1: dout <= 8'b00000000; // 7377 :   0 - 0x0
      13'h1CD2: dout <= 8'b00000000; // 7378 :   0 - 0x0
      13'h1CD3: dout <= 8'b00000000; // 7379 :   0 - 0x0
      13'h1CD4: dout <= 8'b00000000; // 7380 :   0 - 0x0
      13'h1CD5: dout <= 8'b00000000; // 7381 :   0 - 0x0
      13'h1CD6: dout <= 8'b00000000; // 7382 :   0 - 0x0
      13'h1CD7: dout <= 8'b00000000; // 7383 :   0 - 0x0
      13'h1CD8: dout <= 8'b00000000; // 7384 :   0 - 0x0
      13'h1CD9: dout <= 8'b00000000; // 7385 :   0 - 0x0
      13'h1CDA: dout <= 8'b00000000; // 7386 :   0 - 0x0
      13'h1CDB: dout <= 8'b00000000; // 7387 :   0 - 0x0
      13'h1CDC: dout <= 8'b00000000; // 7388 :   0 - 0x0
      13'h1CDD: dout <= 8'b00000000; // 7389 :   0 - 0x0
      13'h1CDE: dout <= 8'b00000000; // 7390 :   0 - 0x0
      13'h1CDF: dout <= 8'b00000000; // 7391 :   0 - 0x0
      13'h1CE0: dout <= 8'b00000000; // 7392 :   0 - 0x0 -- Background 0xce
      13'h1CE1: dout <= 8'b00000000; // 7393 :   0 - 0x0
      13'h1CE2: dout <= 8'b00000000; // 7394 :   0 - 0x0
      13'h1CE3: dout <= 8'b00000000; // 7395 :   0 - 0x0
      13'h1CE4: dout <= 8'b00000000; // 7396 :   0 - 0x0
      13'h1CE5: dout <= 8'b00000000; // 7397 :   0 - 0x0
      13'h1CE6: dout <= 8'b00000000; // 7398 :   0 - 0x0
      13'h1CE7: dout <= 8'b00000000; // 7399 :   0 - 0x0
      13'h1CE8: dout <= 8'b00000000; // 7400 :   0 - 0x0
      13'h1CE9: dout <= 8'b00000000; // 7401 :   0 - 0x0
      13'h1CEA: dout <= 8'b00000000; // 7402 :   0 - 0x0
      13'h1CEB: dout <= 8'b00000000; // 7403 :   0 - 0x0
      13'h1CEC: dout <= 8'b00000000; // 7404 :   0 - 0x0
      13'h1CED: dout <= 8'b00000000; // 7405 :   0 - 0x0
      13'h1CEE: dout <= 8'b00000000; // 7406 :   0 - 0x0
      13'h1CEF: dout <= 8'b00000000; // 7407 :   0 - 0x0
      13'h1CF0: dout <= 8'b00000000; // 7408 :   0 - 0x0 -- Background 0xcf
      13'h1CF1: dout <= 8'b00000000; // 7409 :   0 - 0x0
      13'h1CF2: dout <= 8'b00000000; // 7410 :   0 - 0x0
      13'h1CF3: dout <= 8'b00000000; // 7411 :   0 - 0x0
      13'h1CF4: dout <= 8'b00000000; // 7412 :   0 - 0x0
      13'h1CF5: dout <= 8'b00000000; // 7413 :   0 - 0x0
      13'h1CF6: dout <= 8'b00000000; // 7414 :   0 - 0x0
      13'h1CF7: dout <= 8'b00000000; // 7415 :   0 - 0x0
      13'h1CF8: dout <= 8'b00000000; // 7416 :   0 - 0x0
      13'h1CF9: dout <= 8'b00000000; // 7417 :   0 - 0x0
      13'h1CFA: dout <= 8'b00000000; // 7418 :   0 - 0x0
      13'h1CFB: dout <= 8'b00000000; // 7419 :   0 - 0x0
      13'h1CFC: dout <= 8'b00000000; // 7420 :   0 - 0x0
      13'h1CFD: dout <= 8'b00000000; // 7421 :   0 - 0x0
      13'h1CFE: dout <= 8'b00000000; // 7422 :   0 - 0x0
      13'h1CFF: dout <= 8'b00000000; // 7423 :   0 - 0x0
      13'h1D00: dout <= 8'b11111111; // 7424 : 255 - 0xff -- Background 0xd0
      13'h1D01: dout <= 8'b11111111; // 7425 : 255 - 0xff
      13'h1D02: dout <= 8'b11111111; // 7426 : 255 - 0xff
      13'h1D03: dout <= 8'b11111111; // 7427 : 255 - 0xff
      13'h1D04: dout <= 8'b11111111; // 7428 : 255 - 0xff
      13'h1D05: dout <= 8'b11111111; // 7429 : 255 - 0xff
      13'h1D06: dout <= 8'b11111111; // 7430 : 255 - 0xff
      13'h1D07: dout <= 8'b11111111; // 7431 : 255 - 0xff
      13'h1D08: dout <= 8'b11111111; // 7432 : 255 - 0xff
      13'h1D09: dout <= 8'b11111111; // 7433 : 255 - 0xff
      13'h1D0A: dout <= 8'b11111111; // 7434 : 255 - 0xff
      13'h1D0B: dout <= 8'b11111111; // 7435 : 255 - 0xff
      13'h1D0C: dout <= 8'b11111111; // 7436 : 255 - 0xff
      13'h1D0D: dout <= 8'b11111111; // 7437 : 255 - 0xff
      13'h1D0E: dout <= 8'b11111111; // 7438 : 255 - 0xff
      13'h1D0F: dout <= 8'b11111111; // 7439 : 255 - 0xff
      13'h1D10: dout <= 8'b11111111; // 7440 : 255 - 0xff -- Background 0xd1
      13'h1D11: dout <= 8'b11111111; // 7441 : 255 - 0xff
      13'h1D12: dout <= 8'b11111111; // 7442 : 255 - 0xff
      13'h1D13: dout <= 8'b11111111; // 7443 : 255 - 0xff
      13'h1D14: dout <= 8'b11111111; // 7444 : 255 - 0xff
      13'h1D15: dout <= 8'b11111111; // 7445 : 255 - 0xff
      13'h1D16: dout <= 8'b11111111; // 7446 : 255 - 0xff
      13'h1D17: dout <= 8'b11111111; // 7447 : 255 - 0xff
      13'h1D18: dout <= 8'b11111111; // 7448 : 255 - 0xff
      13'h1D19: dout <= 8'b11111111; // 7449 : 255 - 0xff
      13'h1D1A: dout <= 8'b11111111; // 7450 : 255 - 0xff
      13'h1D1B: dout <= 8'b11111111; // 7451 : 255 - 0xff
      13'h1D1C: dout <= 8'b11111111; // 7452 : 255 - 0xff
      13'h1D1D: dout <= 8'b11111111; // 7453 : 255 - 0xff
      13'h1D1E: dout <= 8'b11111111; // 7454 : 255 - 0xff
      13'h1D1F: dout <= 8'b11111111; // 7455 : 255 - 0xff
      13'h1D20: dout <= 8'b11111111; // 7456 : 255 - 0xff -- Background 0xd2
      13'h1D21: dout <= 8'b11111111; // 7457 : 255 - 0xff
      13'h1D22: dout <= 8'b11111111; // 7458 : 255 - 0xff
      13'h1D23: dout <= 8'b11111111; // 7459 : 255 - 0xff
      13'h1D24: dout <= 8'b11111111; // 7460 : 255 - 0xff
      13'h1D25: dout <= 8'b11111111; // 7461 : 255 - 0xff
      13'h1D26: dout <= 8'b11111111; // 7462 : 255 - 0xff
      13'h1D27: dout <= 8'b11111111; // 7463 : 255 - 0xff
      13'h1D28: dout <= 8'b11111111; // 7464 : 255 - 0xff
      13'h1D29: dout <= 8'b11111111; // 7465 : 255 - 0xff
      13'h1D2A: dout <= 8'b11111111; // 7466 : 255 - 0xff
      13'h1D2B: dout <= 8'b11111111; // 7467 : 255 - 0xff
      13'h1D2C: dout <= 8'b11111111; // 7468 : 255 - 0xff
      13'h1D2D: dout <= 8'b11111111; // 7469 : 255 - 0xff
      13'h1D2E: dout <= 8'b11111111; // 7470 : 255 - 0xff
      13'h1D2F: dout <= 8'b11111111; // 7471 : 255 - 0xff
      13'h1D30: dout <= 8'b11111111; // 7472 : 255 - 0xff -- Background 0xd3
      13'h1D31: dout <= 8'b11111111; // 7473 : 255 - 0xff
      13'h1D32: dout <= 8'b11111111; // 7474 : 255 - 0xff
      13'h1D33: dout <= 8'b11111111; // 7475 : 255 - 0xff
      13'h1D34: dout <= 8'b11111111; // 7476 : 255 - 0xff
      13'h1D35: dout <= 8'b11111111; // 7477 : 255 - 0xff
      13'h1D36: dout <= 8'b11111111; // 7478 : 255 - 0xff
      13'h1D37: dout <= 8'b11111111; // 7479 : 255 - 0xff
      13'h1D38: dout <= 8'b11111111; // 7480 : 255 - 0xff
      13'h1D39: dout <= 8'b11111111; // 7481 : 255 - 0xff
      13'h1D3A: dout <= 8'b11111111; // 7482 : 255 - 0xff
      13'h1D3B: dout <= 8'b11111111; // 7483 : 255 - 0xff
      13'h1D3C: dout <= 8'b11111111; // 7484 : 255 - 0xff
      13'h1D3D: dout <= 8'b11111111; // 7485 : 255 - 0xff
      13'h1D3E: dout <= 8'b11111111; // 7486 : 255 - 0xff
      13'h1D3F: dout <= 8'b11111111; // 7487 : 255 - 0xff
      13'h1D40: dout <= 8'b11111111; // 7488 : 255 - 0xff -- Background 0xd4
      13'h1D41: dout <= 8'b11111111; // 7489 : 255 - 0xff
      13'h1D42: dout <= 8'b11111111; // 7490 : 255 - 0xff
      13'h1D43: dout <= 8'b11111111; // 7491 : 255 - 0xff
      13'h1D44: dout <= 8'b11111111; // 7492 : 255 - 0xff
      13'h1D45: dout <= 8'b11111111; // 7493 : 255 - 0xff
      13'h1D46: dout <= 8'b11111111; // 7494 : 255 - 0xff
      13'h1D47: dout <= 8'b11111111; // 7495 : 255 - 0xff
      13'h1D48: dout <= 8'b11111111; // 7496 : 255 - 0xff
      13'h1D49: dout <= 8'b11111111; // 7497 : 255 - 0xff
      13'h1D4A: dout <= 8'b11111111; // 7498 : 255 - 0xff
      13'h1D4B: dout <= 8'b11111111; // 7499 : 255 - 0xff
      13'h1D4C: dout <= 8'b11111111; // 7500 : 255 - 0xff
      13'h1D4D: dout <= 8'b11111111; // 7501 : 255 - 0xff
      13'h1D4E: dout <= 8'b11111111; // 7502 : 255 - 0xff
      13'h1D4F: dout <= 8'b11111111; // 7503 : 255 - 0xff
      13'h1D50: dout <= 8'b11111111; // 7504 : 255 - 0xff -- Background 0xd5
      13'h1D51: dout <= 8'b11111111; // 7505 : 255 - 0xff
      13'h1D52: dout <= 8'b11111111; // 7506 : 255 - 0xff
      13'h1D53: dout <= 8'b11111111; // 7507 : 255 - 0xff
      13'h1D54: dout <= 8'b11111111; // 7508 : 255 - 0xff
      13'h1D55: dout <= 8'b11111111; // 7509 : 255 - 0xff
      13'h1D56: dout <= 8'b11111111; // 7510 : 255 - 0xff
      13'h1D57: dout <= 8'b11111111; // 7511 : 255 - 0xff
      13'h1D58: dout <= 8'b11111111; // 7512 : 255 - 0xff
      13'h1D59: dout <= 8'b11111111; // 7513 : 255 - 0xff
      13'h1D5A: dout <= 8'b11111111; // 7514 : 255 - 0xff
      13'h1D5B: dout <= 8'b11111111; // 7515 : 255 - 0xff
      13'h1D5C: dout <= 8'b11111111; // 7516 : 255 - 0xff
      13'h1D5D: dout <= 8'b11111111; // 7517 : 255 - 0xff
      13'h1D5E: dout <= 8'b11111111; // 7518 : 255 - 0xff
      13'h1D5F: dout <= 8'b11111111; // 7519 : 255 - 0xff
      13'h1D60: dout <= 8'b11111111; // 7520 : 255 - 0xff -- Background 0xd6
      13'h1D61: dout <= 8'b11111111; // 7521 : 255 - 0xff
      13'h1D62: dout <= 8'b11111111; // 7522 : 255 - 0xff
      13'h1D63: dout <= 8'b11111111; // 7523 : 255 - 0xff
      13'h1D64: dout <= 8'b11111111; // 7524 : 255 - 0xff
      13'h1D65: dout <= 8'b11111111; // 7525 : 255 - 0xff
      13'h1D66: dout <= 8'b11111111; // 7526 : 255 - 0xff
      13'h1D67: dout <= 8'b11111111; // 7527 : 255 - 0xff
      13'h1D68: dout <= 8'b11111111; // 7528 : 255 - 0xff
      13'h1D69: dout <= 8'b11111111; // 7529 : 255 - 0xff
      13'h1D6A: dout <= 8'b11111111; // 7530 : 255 - 0xff
      13'h1D6B: dout <= 8'b11111111; // 7531 : 255 - 0xff
      13'h1D6C: dout <= 8'b11111111; // 7532 : 255 - 0xff
      13'h1D6D: dout <= 8'b11111111; // 7533 : 255 - 0xff
      13'h1D6E: dout <= 8'b11111111; // 7534 : 255 - 0xff
      13'h1D6F: dout <= 8'b11111111; // 7535 : 255 - 0xff
      13'h1D70: dout <= 8'b11111111; // 7536 : 255 - 0xff -- Background 0xd7
      13'h1D71: dout <= 8'b11111111; // 7537 : 255 - 0xff
      13'h1D72: dout <= 8'b11111111; // 7538 : 255 - 0xff
      13'h1D73: dout <= 8'b11111111; // 7539 : 255 - 0xff
      13'h1D74: dout <= 8'b11111111; // 7540 : 255 - 0xff
      13'h1D75: dout <= 8'b11111111; // 7541 : 255 - 0xff
      13'h1D76: dout <= 8'b11111111; // 7542 : 255 - 0xff
      13'h1D77: dout <= 8'b11111111; // 7543 : 255 - 0xff
      13'h1D78: dout <= 8'b11111111; // 7544 : 255 - 0xff
      13'h1D79: dout <= 8'b11111111; // 7545 : 255 - 0xff
      13'h1D7A: dout <= 8'b11111111; // 7546 : 255 - 0xff
      13'h1D7B: dout <= 8'b11111111; // 7547 : 255 - 0xff
      13'h1D7C: dout <= 8'b11111111; // 7548 : 255 - 0xff
      13'h1D7D: dout <= 8'b11111111; // 7549 : 255 - 0xff
      13'h1D7E: dout <= 8'b11111111; // 7550 : 255 - 0xff
      13'h1D7F: dout <= 8'b11111111; // 7551 : 255 - 0xff
      13'h1D80: dout <= 8'b11111111; // 7552 : 255 - 0xff -- Background 0xd8
      13'h1D81: dout <= 8'b11111111; // 7553 : 255 - 0xff
      13'h1D82: dout <= 8'b11111111; // 7554 : 255 - 0xff
      13'h1D83: dout <= 8'b11111111; // 7555 : 255 - 0xff
      13'h1D84: dout <= 8'b11111111; // 7556 : 255 - 0xff
      13'h1D85: dout <= 8'b11111111; // 7557 : 255 - 0xff
      13'h1D86: dout <= 8'b11111111; // 7558 : 255 - 0xff
      13'h1D87: dout <= 8'b11111111; // 7559 : 255 - 0xff
      13'h1D88: dout <= 8'b11111111; // 7560 : 255 - 0xff
      13'h1D89: dout <= 8'b11111111; // 7561 : 255 - 0xff
      13'h1D8A: dout <= 8'b11111111; // 7562 : 255 - 0xff
      13'h1D8B: dout <= 8'b11111111; // 7563 : 255 - 0xff
      13'h1D8C: dout <= 8'b11111111; // 7564 : 255 - 0xff
      13'h1D8D: dout <= 8'b11111111; // 7565 : 255 - 0xff
      13'h1D8E: dout <= 8'b11111111; // 7566 : 255 - 0xff
      13'h1D8F: dout <= 8'b11111111; // 7567 : 255 - 0xff
      13'h1D90: dout <= 8'b11111111; // 7568 : 255 - 0xff -- Background 0xd9
      13'h1D91: dout <= 8'b11111111; // 7569 : 255 - 0xff
      13'h1D92: dout <= 8'b11111111; // 7570 : 255 - 0xff
      13'h1D93: dout <= 8'b11111111; // 7571 : 255 - 0xff
      13'h1D94: dout <= 8'b11111111; // 7572 : 255 - 0xff
      13'h1D95: dout <= 8'b11111111; // 7573 : 255 - 0xff
      13'h1D96: dout <= 8'b11111111; // 7574 : 255 - 0xff
      13'h1D97: dout <= 8'b11111111; // 7575 : 255 - 0xff
      13'h1D98: dout <= 8'b11111111; // 7576 : 255 - 0xff
      13'h1D99: dout <= 8'b11111111; // 7577 : 255 - 0xff
      13'h1D9A: dout <= 8'b11111111; // 7578 : 255 - 0xff
      13'h1D9B: dout <= 8'b11111111; // 7579 : 255 - 0xff
      13'h1D9C: dout <= 8'b11111111; // 7580 : 255 - 0xff
      13'h1D9D: dout <= 8'b11111111; // 7581 : 255 - 0xff
      13'h1D9E: dout <= 8'b11111111; // 7582 : 255 - 0xff
      13'h1D9F: dout <= 8'b11111111; // 7583 : 255 - 0xff
      13'h1DA0: dout <= 8'b11111111; // 7584 : 255 - 0xff -- Background 0xda
      13'h1DA1: dout <= 8'b11111111; // 7585 : 255 - 0xff
      13'h1DA2: dout <= 8'b11111111; // 7586 : 255 - 0xff
      13'h1DA3: dout <= 8'b11111111; // 7587 : 255 - 0xff
      13'h1DA4: dout <= 8'b11111111; // 7588 : 255 - 0xff
      13'h1DA5: dout <= 8'b11111111; // 7589 : 255 - 0xff
      13'h1DA6: dout <= 8'b11111111; // 7590 : 255 - 0xff
      13'h1DA7: dout <= 8'b11111111; // 7591 : 255 - 0xff
      13'h1DA8: dout <= 8'b11111111; // 7592 : 255 - 0xff
      13'h1DA9: dout <= 8'b11111111; // 7593 : 255 - 0xff
      13'h1DAA: dout <= 8'b11111111; // 7594 : 255 - 0xff
      13'h1DAB: dout <= 8'b11111111; // 7595 : 255 - 0xff
      13'h1DAC: dout <= 8'b11111111; // 7596 : 255 - 0xff
      13'h1DAD: dout <= 8'b11111111; // 7597 : 255 - 0xff
      13'h1DAE: dout <= 8'b11111111; // 7598 : 255 - 0xff
      13'h1DAF: dout <= 8'b11111111; // 7599 : 255 - 0xff
      13'h1DB0: dout <= 8'b11111111; // 7600 : 255 - 0xff -- Background 0xdb
      13'h1DB1: dout <= 8'b11111111; // 7601 : 255 - 0xff
      13'h1DB2: dout <= 8'b11111111; // 7602 : 255 - 0xff
      13'h1DB3: dout <= 8'b11111111; // 7603 : 255 - 0xff
      13'h1DB4: dout <= 8'b11111111; // 7604 : 255 - 0xff
      13'h1DB5: dout <= 8'b11111111; // 7605 : 255 - 0xff
      13'h1DB6: dout <= 8'b11111111; // 7606 : 255 - 0xff
      13'h1DB7: dout <= 8'b11111111; // 7607 : 255 - 0xff
      13'h1DB8: dout <= 8'b11111111; // 7608 : 255 - 0xff
      13'h1DB9: dout <= 8'b11111111; // 7609 : 255 - 0xff
      13'h1DBA: dout <= 8'b11111111; // 7610 : 255 - 0xff
      13'h1DBB: dout <= 8'b11111111; // 7611 : 255 - 0xff
      13'h1DBC: dout <= 8'b11111111; // 7612 : 255 - 0xff
      13'h1DBD: dout <= 8'b11111111; // 7613 : 255 - 0xff
      13'h1DBE: dout <= 8'b11111111; // 7614 : 255 - 0xff
      13'h1DBF: dout <= 8'b11111111; // 7615 : 255 - 0xff
      13'h1DC0: dout <= 8'b11111111; // 7616 : 255 - 0xff -- Background 0xdc
      13'h1DC1: dout <= 8'b11111111; // 7617 : 255 - 0xff
      13'h1DC2: dout <= 8'b11111111; // 7618 : 255 - 0xff
      13'h1DC3: dout <= 8'b11111111; // 7619 : 255 - 0xff
      13'h1DC4: dout <= 8'b11111111; // 7620 : 255 - 0xff
      13'h1DC5: dout <= 8'b11111111; // 7621 : 255 - 0xff
      13'h1DC6: dout <= 8'b11111111; // 7622 : 255 - 0xff
      13'h1DC7: dout <= 8'b11111111; // 7623 : 255 - 0xff
      13'h1DC8: dout <= 8'b11111111; // 7624 : 255 - 0xff
      13'h1DC9: dout <= 8'b11111111; // 7625 : 255 - 0xff
      13'h1DCA: dout <= 8'b11111111; // 7626 : 255 - 0xff
      13'h1DCB: dout <= 8'b11111111; // 7627 : 255 - 0xff
      13'h1DCC: dout <= 8'b11111111; // 7628 : 255 - 0xff
      13'h1DCD: dout <= 8'b11111111; // 7629 : 255 - 0xff
      13'h1DCE: dout <= 8'b11111111; // 7630 : 255 - 0xff
      13'h1DCF: dout <= 8'b11111111; // 7631 : 255 - 0xff
      13'h1DD0: dout <= 8'b11111111; // 7632 : 255 - 0xff -- Background 0xdd
      13'h1DD1: dout <= 8'b11111111; // 7633 : 255 - 0xff
      13'h1DD2: dout <= 8'b11111111; // 7634 : 255 - 0xff
      13'h1DD3: dout <= 8'b11111111; // 7635 : 255 - 0xff
      13'h1DD4: dout <= 8'b11111111; // 7636 : 255 - 0xff
      13'h1DD5: dout <= 8'b11111111; // 7637 : 255 - 0xff
      13'h1DD6: dout <= 8'b11111111; // 7638 : 255 - 0xff
      13'h1DD7: dout <= 8'b11111111; // 7639 : 255 - 0xff
      13'h1DD8: dout <= 8'b11111111; // 7640 : 255 - 0xff
      13'h1DD9: dout <= 8'b11111111; // 7641 : 255 - 0xff
      13'h1DDA: dout <= 8'b11111111; // 7642 : 255 - 0xff
      13'h1DDB: dout <= 8'b11111111; // 7643 : 255 - 0xff
      13'h1DDC: dout <= 8'b11111111; // 7644 : 255 - 0xff
      13'h1DDD: dout <= 8'b11111111; // 7645 : 255 - 0xff
      13'h1DDE: dout <= 8'b11111111; // 7646 : 255 - 0xff
      13'h1DDF: dout <= 8'b11111111; // 7647 : 255 - 0xff
      13'h1DE0: dout <= 8'b11111111; // 7648 : 255 - 0xff -- Background 0xde
      13'h1DE1: dout <= 8'b11111111; // 7649 : 255 - 0xff
      13'h1DE2: dout <= 8'b11111111; // 7650 : 255 - 0xff
      13'h1DE3: dout <= 8'b11111111; // 7651 : 255 - 0xff
      13'h1DE4: dout <= 8'b11111111; // 7652 : 255 - 0xff
      13'h1DE5: dout <= 8'b11111111; // 7653 : 255 - 0xff
      13'h1DE6: dout <= 8'b11111111; // 7654 : 255 - 0xff
      13'h1DE7: dout <= 8'b11111111; // 7655 : 255 - 0xff
      13'h1DE8: dout <= 8'b11111111; // 7656 : 255 - 0xff
      13'h1DE9: dout <= 8'b11111111; // 7657 : 255 - 0xff
      13'h1DEA: dout <= 8'b11111111; // 7658 : 255 - 0xff
      13'h1DEB: dout <= 8'b11111111; // 7659 : 255 - 0xff
      13'h1DEC: dout <= 8'b11111111; // 7660 : 255 - 0xff
      13'h1DED: dout <= 8'b11111111; // 7661 : 255 - 0xff
      13'h1DEE: dout <= 8'b11111111; // 7662 : 255 - 0xff
      13'h1DEF: dout <= 8'b11111111; // 7663 : 255 - 0xff
      13'h1DF0: dout <= 8'b11111111; // 7664 : 255 - 0xff -- Background 0xdf
      13'h1DF1: dout <= 8'b11111111; // 7665 : 255 - 0xff
      13'h1DF2: dout <= 8'b11111111; // 7666 : 255 - 0xff
      13'h1DF3: dout <= 8'b11111111; // 7667 : 255 - 0xff
      13'h1DF4: dout <= 8'b11111111; // 7668 : 255 - 0xff
      13'h1DF5: dout <= 8'b11111111; // 7669 : 255 - 0xff
      13'h1DF6: dout <= 8'b11111111; // 7670 : 255 - 0xff
      13'h1DF7: dout <= 8'b11111111; // 7671 : 255 - 0xff
      13'h1DF8: dout <= 8'b11111111; // 7672 : 255 - 0xff
      13'h1DF9: dout <= 8'b11111111; // 7673 : 255 - 0xff
      13'h1DFA: dout <= 8'b11111111; // 7674 : 255 - 0xff
      13'h1DFB: dout <= 8'b11111111; // 7675 : 255 - 0xff
      13'h1DFC: dout <= 8'b11111111; // 7676 : 255 - 0xff
      13'h1DFD: dout <= 8'b11111111; // 7677 : 255 - 0xff
      13'h1DFE: dout <= 8'b11111111; // 7678 : 255 - 0xff
      13'h1DFF: dout <= 8'b11111111; // 7679 : 255 - 0xff
      13'h1E00: dout <= 8'b11111111; // 7680 : 255 - 0xff -- Background 0xe0
      13'h1E01: dout <= 8'b11111111; // 7681 : 255 - 0xff
      13'h1E02: dout <= 8'b11111111; // 7682 : 255 - 0xff
      13'h1E03: dout <= 8'b11111111; // 7683 : 255 - 0xff
      13'h1E04: dout <= 8'b11111111; // 7684 : 255 - 0xff
      13'h1E05: dout <= 8'b11111111; // 7685 : 255 - 0xff
      13'h1E06: dout <= 8'b11111111; // 7686 : 255 - 0xff
      13'h1E07: dout <= 8'b11111111; // 7687 : 255 - 0xff
      13'h1E08: dout <= 8'b11111111; // 7688 : 255 - 0xff
      13'h1E09: dout <= 8'b11111111; // 7689 : 255 - 0xff
      13'h1E0A: dout <= 8'b11111111; // 7690 : 255 - 0xff
      13'h1E0B: dout <= 8'b11111111; // 7691 : 255 - 0xff
      13'h1E0C: dout <= 8'b11111111; // 7692 : 255 - 0xff
      13'h1E0D: dout <= 8'b11111111; // 7693 : 255 - 0xff
      13'h1E0E: dout <= 8'b11111111; // 7694 : 255 - 0xff
      13'h1E0F: dout <= 8'b11111111; // 7695 : 255 - 0xff
      13'h1E10: dout <= 8'b11111111; // 7696 : 255 - 0xff -- Background 0xe1
      13'h1E11: dout <= 8'b11111111; // 7697 : 255 - 0xff
      13'h1E12: dout <= 8'b11111111; // 7698 : 255 - 0xff
      13'h1E13: dout <= 8'b11111111; // 7699 : 255 - 0xff
      13'h1E14: dout <= 8'b11111111; // 7700 : 255 - 0xff
      13'h1E15: dout <= 8'b11111111; // 7701 : 255 - 0xff
      13'h1E16: dout <= 8'b11111111; // 7702 : 255 - 0xff
      13'h1E17: dout <= 8'b11111111; // 7703 : 255 - 0xff
      13'h1E18: dout <= 8'b11111111; // 7704 : 255 - 0xff
      13'h1E19: dout <= 8'b11111111; // 7705 : 255 - 0xff
      13'h1E1A: dout <= 8'b11111111; // 7706 : 255 - 0xff
      13'h1E1B: dout <= 8'b11111111; // 7707 : 255 - 0xff
      13'h1E1C: dout <= 8'b11111111; // 7708 : 255 - 0xff
      13'h1E1D: dout <= 8'b11111111; // 7709 : 255 - 0xff
      13'h1E1E: dout <= 8'b11111111; // 7710 : 255 - 0xff
      13'h1E1F: dout <= 8'b11111111; // 7711 : 255 - 0xff
      13'h1E20: dout <= 8'b11111111; // 7712 : 255 - 0xff -- Background 0xe2
      13'h1E21: dout <= 8'b11111111; // 7713 : 255 - 0xff
      13'h1E22: dout <= 8'b11111111; // 7714 : 255 - 0xff
      13'h1E23: dout <= 8'b11111111; // 7715 : 255 - 0xff
      13'h1E24: dout <= 8'b11111111; // 7716 : 255 - 0xff
      13'h1E25: dout <= 8'b11111111; // 7717 : 255 - 0xff
      13'h1E26: dout <= 8'b11111111; // 7718 : 255 - 0xff
      13'h1E27: dout <= 8'b11111111; // 7719 : 255 - 0xff
      13'h1E28: dout <= 8'b11111111; // 7720 : 255 - 0xff
      13'h1E29: dout <= 8'b11111111; // 7721 : 255 - 0xff
      13'h1E2A: dout <= 8'b11111111; // 7722 : 255 - 0xff
      13'h1E2B: dout <= 8'b11111111; // 7723 : 255 - 0xff
      13'h1E2C: dout <= 8'b11111111; // 7724 : 255 - 0xff
      13'h1E2D: dout <= 8'b11111111; // 7725 : 255 - 0xff
      13'h1E2E: dout <= 8'b11111111; // 7726 : 255 - 0xff
      13'h1E2F: dout <= 8'b11111111; // 7727 : 255 - 0xff
      13'h1E30: dout <= 8'b11111111; // 7728 : 255 - 0xff -- Background 0xe3
      13'h1E31: dout <= 8'b11111111; // 7729 : 255 - 0xff
      13'h1E32: dout <= 8'b11111111; // 7730 : 255 - 0xff
      13'h1E33: dout <= 8'b11111111; // 7731 : 255 - 0xff
      13'h1E34: dout <= 8'b11111111; // 7732 : 255 - 0xff
      13'h1E35: dout <= 8'b11111111; // 7733 : 255 - 0xff
      13'h1E36: dout <= 8'b11111111; // 7734 : 255 - 0xff
      13'h1E37: dout <= 8'b11111111; // 7735 : 255 - 0xff
      13'h1E38: dout <= 8'b11111111; // 7736 : 255 - 0xff
      13'h1E39: dout <= 8'b11111111; // 7737 : 255 - 0xff
      13'h1E3A: dout <= 8'b11111111; // 7738 : 255 - 0xff
      13'h1E3B: dout <= 8'b11111111; // 7739 : 255 - 0xff
      13'h1E3C: dout <= 8'b11111111; // 7740 : 255 - 0xff
      13'h1E3D: dout <= 8'b11111111; // 7741 : 255 - 0xff
      13'h1E3E: dout <= 8'b11111111; // 7742 : 255 - 0xff
      13'h1E3F: dout <= 8'b11111111; // 7743 : 255 - 0xff
      13'h1E40: dout <= 8'b11111111; // 7744 : 255 - 0xff -- Background 0xe4
      13'h1E41: dout <= 8'b11111111; // 7745 : 255 - 0xff
      13'h1E42: dout <= 8'b11111111; // 7746 : 255 - 0xff
      13'h1E43: dout <= 8'b11111111; // 7747 : 255 - 0xff
      13'h1E44: dout <= 8'b11111111; // 7748 : 255 - 0xff
      13'h1E45: dout <= 8'b11111111; // 7749 : 255 - 0xff
      13'h1E46: dout <= 8'b11111111; // 7750 : 255 - 0xff
      13'h1E47: dout <= 8'b11111111; // 7751 : 255 - 0xff
      13'h1E48: dout <= 8'b11111111; // 7752 : 255 - 0xff
      13'h1E49: dout <= 8'b11111111; // 7753 : 255 - 0xff
      13'h1E4A: dout <= 8'b11111111; // 7754 : 255 - 0xff
      13'h1E4B: dout <= 8'b11111111; // 7755 : 255 - 0xff
      13'h1E4C: dout <= 8'b11111111; // 7756 : 255 - 0xff
      13'h1E4D: dout <= 8'b11111111; // 7757 : 255 - 0xff
      13'h1E4E: dout <= 8'b11111111; // 7758 : 255 - 0xff
      13'h1E4F: dout <= 8'b11111111; // 7759 : 255 - 0xff
      13'h1E50: dout <= 8'b11111111; // 7760 : 255 - 0xff -- Background 0xe5
      13'h1E51: dout <= 8'b11111111; // 7761 : 255 - 0xff
      13'h1E52: dout <= 8'b11111111; // 7762 : 255 - 0xff
      13'h1E53: dout <= 8'b11111111; // 7763 : 255 - 0xff
      13'h1E54: dout <= 8'b11111111; // 7764 : 255 - 0xff
      13'h1E55: dout <= 8'b11111111; // 7765 : 255 - 0xff
      13'h1E56: dout <= 8'b11111111; // 7766 : 255 - 0xff
      13'h1E57: dout <= 8'b11111111; // 7767 : 255 - 0xff
      13'h1E58: dout <= 8'b11111111; // 7768 : 255 - 0xff
      13'h1E59: dout <= 8'b11111111; // 7769 : 255 - 0xff
      13'h1E5A: dout <= 8'b11111111; // 7770 : 255 - 0xff
      13'h1E5B: dout <= 8'b11111111; // 7771 : 255 - 0xff
      13'h1E5C: dout <= 8'b11111111; // 7772 : 255 - 0xff
      13'h1E5D: dout <= 8'b11111111; // 7773 : 255 - 0xff
      13'h1E5E: dout <= 8'b11111111; // 7774 : 255 - 0xff
      13'h1E5F: dout <= 8'b11111111; // 7775 : 255 - 0xff
      13'h1E60: dout <= 8'b11111111; // 7776 : 255 - 0xff -- Background 0xe6
      13'h1E61: dout <= 8'b11111111; // 7777 : 255 - 0xff
      13'h1E62: dout <= 8'b11111111; // 7778 : 255 - 0xff
      13'h1E63: dout <= 8'b11111111; // 7779 : 255 - 0xff
      13'h1E64: dout <= 8'b11111111; // 7780 : 255 - 0xff
      13'h1E65: dout <= 8'b11111111; // 7781 : 255 - 0xff
      13'h1E66: dout <= 8'b11111111; // 7782 : 255 - 0xff
      13'h1E67: dout <= 8'b11111111; // 7783 : 255 - 0xff
      13'h1E68: dout <= 8'b11111111; // 7784 : 255 - 0xff
      13'h1E69: dout <= 8'b11111111; // 7785 : 255 - 0xff
      13'h1E6A: dout <= 8'b11111111; // 7786 : 255 - 0xff
      13'h1E6B: dout <= 8'b11111111; // 7787 : 255 - 0xff
      13'h1E6C: dout <= 8'b11111111; // 7788 : 255 - 0xff
      13'h1E6D: dout <= 8'b11111111; // 7789 : 255 - 0xff
      13'h1E6E: dout <= 8'b11111111; // 7790 : 255 - 0xff
      13'h1E6F: dout <= 8'b11111111; // 7791 : 255 - 0xff
      13'h1E70: dout <= 8'b11111111; // 7792 : 255 - 0xff -- Background 0xe7
      13'h1E71: dout <= 8'b11111111; // 7793 : 255 - 0xff
      13'h1E72: dout <= 8'b11111111; // 7794 : 255 - 0xff
      13'h1E73: dout <= 8'b11111111; // 7795 : 255 - 0xff
      13'h1E74: dout <= 8'b11111111; // 7796 : 255 - 0xff
      13'h1E75: dout <= 8'b11111111; // 7797 : 255 - 0xff
      13'h1E76: dout <= 8'b11111111; // 7798 : 255 - 0xff
      13'h1E77: dout <= 8'b11111111; // 7799 : 255 - 0xff
      13'h1E78: dout <= 8'b11111111; // 7800 : 255 - 0xff
      13'h1E79: dout <= 8'b11111111; // 7801 : 255 - 0xff
      13'h1E7A: dout <= 8'b11111111; // 7802 : 255 - 0xff
      13'h1E7B: dout <= 8'b11111111; // 7803 : 255 - 0xff
      13'h1E7C: dout <= 8'b11111111; // 7804 : 255 - 0xff
      13'h1E7D: dout <= 8'b11111111; // 7805 : 255 - 0xff
      13'h1E7E: dout <= 8'b11111111; // 7806 : 255 - 0xff
      13'h1E7F: dout <= 8'b11111111; // 7807 : 255 - 0xff
      13'h1E80: dout <= 8'b11111111; // 7808 : 255 - 0xff -- Background 0xe8
      13'h1E81: dout <= 8'b11111111; // 7809 : 255 - 0xff
      13'h1E82: dout <= 8'b11111111; // 7810 : 255 - 0xff
      13'h1E83: dout <= 8'b11111111; // 7811 : 255 - 0xff
      13'h1E84: dout <= 8'b11111111; // 7812 : 255 - 0xff
      13'h1E85: dout <= 8'b11111111; // 7813 : 255 - 0xff
      13'h1E86: dout <= 8'b11111111; // 7814 : 255 - 0xff
      13'h1E87: dout <= 8'b11111111; // 7815 : 255 - 0xff
      13'h1E88: dout <= 8'b11111111; // 7816 : 255 - 0xff
      13'h1E89: dout <= 8'b11111111; // 7817 : 255 - 0xff
      13'h1E8A: dout <= 8'b11111111; // 7818 : 255 - 0xff
      13'h1E8B: dout <= 8'b11111111; // 7819 : 255 - 0xff
      13'h1E8C: dout <= 8'b11111111; // 7820 : 255 - 0xff
      13'h1E8D: dout <= 8'b11111111; // 7821 : 255 - 0xff
      13'h1E8E: dout <= 8'b11111111; // 7822 : 255 - 0xff
      13'h1E8F: dout <= 8'b11111111; // 7823 : 255 - 0xff
      13'h1E90: dout <= 8'b11111111; // 7824 : 255 - 0xff -- Background 0xe9
      13'h1E91: dout <= 8'b11111111; // 7825 : 255 - 0xff
      13'h1E92: dout <= 8'b11111111; // 7826 : 255 - 0xff
      13'h1E93: dout <= 8'b11111111; // 7827 : 255 - 0xff
      13'h1E94: dout <= 8'b11111111; // 7828 : 255 - 0xff
      13'h1E95: dout <= 8'b11111111; // 7829 : 255 - 0xff
      13'h1E96: dout <= 8'b11111111; // 7830 : 255 - 0xff
      13'h1E97: dout <= 8'b11111111; // 7831 : 255 - 0xff
      13'h1E98: dout <= 8'b11111111; // 7832 : 255 - 0xff
      13'h1E99: dout <= 8'b11111111; // 7833 : 255 - 0xff
      13'h1E9A: dout <= 8'b11111111; // 7834 : 255 - 0xff
      13'h1E9B: dout <= 8'b11111111; // 7835 : 255 - 0xff
      13'h1E9C: dout <= 8'b11111111; // 7836 : 255 - 0xff
      13'h1E9D: dout <= 8'b11111111; // 7837 : 255 - 0xff
      13'h1E9E: dout <= 8'b11111111; // 7838 : 255 - 0xff
      13'h1E9F: dout <= 8'b11111111; // 7839 : 255 - 0xff
      13'h1EA0: dout <= 8'b11111111; // 7840 : 255 - 0xff -- Background 0xea
      13'h1EA1: dout <= 8'b11111111; // 7841 : 255 - 0xff
      13'h1EA2: dout <= 8'b11111111; // 7842 : 255 - 0xff
      13'h1EA3: dout <= 8'b11111111; // 7843 : 255 - 0xff
      13'h1EA4: dout <= 8'b11111111; // 7844 : 255 - 0xff
      13'h1EA5: dout <= 8'b11111111; // 7845 : 255 - 0xff
      13'h1EA6: dout <= 8'b11111111; // 7846 : 255 - 0xff
      13'h1EA7: dout <= 8'b11111111; // 7847 : 255 - 0xff
      13'h1EA8: dout <= 8'b11111111; // 7848 : 255 - 0xff
      13'h1EA9: dout <= 8'b11111111; // 7849 : 255 - 0xff
      13'h1EAA: dout <= 8'b11111111; // 7850 : 255 - 0xff
      13'h1EAB: dout <= 8'b11111111; // 7851 : 255 - 0xff
      13'h1EAC: dout <= 8'b11111111; // 7852 : 255 - 0xff
      13'h1EAD: dout <= 8'b11111111; // 7853 : 255 - 0xff
      13'h1EAE: dout <= 8'b11111111; // 7854 : 255 - 0xff
      13'h1EAF: dout <= 8'b11111111; // 7855 : 255 - 0xff
      13'h1EB0: dout <= 8'b11111111; // 7856 : 255 - 0xff -- Background 0xeb
      13'h1EB1: dout <= 8'b11111111; // 7857 : 255 - 0xff
      13'h1EB2: dout <= 8'b11111111; // 7858 : 255 - 0xff
      13'h1EB3: dout <= 8'b11111111; // 7859 : 255 - 0xff
      13'h1EB4: dout <= 8'b11111111; // 7860 : 255 - 0xff
      13'h1EB5: dout <= 8'b11111111; // 7861 : 255 - 0xff
      13'h1EB6: dout <= 8'b11111111; // 7862 : 255 - 0xff
      13'h1EB7: dout <= 8'b11111111; // 7863 : 255 - 0xff
      13'h1EB8: dout <= 8'b11111111; // 7864 : 255 - 0xff
      13'h1EB9: dout <= 8'b11111111; // 7865 : 255 - 0xff
      13'h1EBA: dout <= 8'b11111111; // 7866 : 255 - 0xff
      13'h1EBB: dout <= 8'b11111111; // 7867 : 255 - 0xff
      13'h1EBC: dout <= 8'b11111111; // 7868 : 255 - 0xff
      13'h1EBD: dout <= 8'b11111111; // 7869 : 255 - 0xff
      13'h1EBE: dout <= 8'b11111111; // 7870 : 255 - 0xff
      13'h1EBF: dout <= 8'b11111111; // 7871 : 255 - 0xff
      13'h1EC0: dout <= 8'b11111111; // 7872 : 255 - 0xff -- Background 0xec
      13'h1EC1: dout <= 8'b11111111; // 7873 : 255 - 0xff
      13'h1EC2: dout <= 8'b11111111; // 7874 : 255 - 0xff
      13'h1EC3: dout <= 8'b11111111; // 7875 : 255 - 0xff
      13'h1EC4: dout <= 8'b11111111; // 7876 : 255 - 0xff
      13'h1EC5: dout <= 8'b11111111; // 7877 : 255 - 0xff
      13'h1EC6: dout <= 8'b11111111; // 7878 : 255 - 0xff
      13'h1EC7: dout <= 8'b11111111; // 7879 : 255 - 0xff
      13'h1EC8: dout <= 8'b11111111; // 7880 : 255 - 0xff
      13'h1EC9: dout <= 8'b11111111; // 7881 : 255 - 0xff
      13'h1ECA: dout <= 8'b11111111; // 7882 : 255 - 0xff
      13'h1ECB: dout <= 8'b11111111; // 7883 : 255 - 0xff
      13'h1ECC: dout <= 8'b11111111; // 7884 : 255 - 0xff
      13'h1ECD: dout <= 8'b11111111; // 7885 : 255 - 0xff
      13'h1ECE: dout <= 8'b11111111; // 7886 : 255 - 0xff
      13'h1ECF: dout <= 8'b11111111; // 7887 : 255 - 0xff
      13'h1ED0: dout <= 8'b11111111; // 7888 : 255 - 0xff -- Background 0xed
      13'h1ED1: dout <= 8'b11111111; // 7889 : 255 - 0xff
      13'h1ED2: dout <= 8'b11111111; // 7890 : 255 - 0xff
      13'h1ED3: dout <= 8'b11111111; // 7891 : 255 - 0xff
      13'h1ED4: dout <= 8'b11111111; // 7892 : 255 - 0xff
      13'h1ED5: dout <= 8'b11111111; // 7893 : 255 - 0xff
      13'h1ED6: dout <= 8'b11111111; // 7894 : 255 - 0xff
      13'h1ED7: dout <= 8'b11111111; // 7895 : 255 - 0xff
      13'h1ED8: dout <= 8'b11111111; // 7896 : 255 - 0xff
      13'h1ED9: dout <= 8'b11111111; // 7897 : 255 - 0xff
      13'h1EDA: dout <= 8'b11111111; // 7898 : 255 - 0xff
      13'h1EDB: dout <= 8'b11111111; // 7899 : 255 - 0xff
      13'h1EDC: dout <= 8'b11111111; // 7900 : 255 - 0xff
      13'h1EDD: dout <= 8'b11111111; // 7901 : 255 - 0xff
      13'h1EDE: dout <= 8'b11111111; // 7902 : 255 - 0xff
      13'h1EDF: dout <= 8'b11111111; // 7903 : 255 - 0xff
      13'h1EE0: dout <= 8'b11111111; // 7904 : 255 - 0xff -- Background 0xee
      13'h1EE1: dout <= 8'b11111111; // 7905 : 255 - 0xff
      13'h1EE2: dout <= 8'b11111111; // 7906 : 255 - 0xff
      13'h1EE3: dout <= 8'b11111111; // 7907 : 255 - 0xff
      13'h1EE4: dout <= 8'b11111111; // 7908 : 255 - 0xff
      13'h1EE5: dout <= 8'b11111111; // 7909 : 255 - 0xff
      13'h1EE6: dout <= 8'b11111111; // 7910 : 255 - 0xff
      13'h1EE7: dout <= 8'b11111111; // 7911 : 255 - 0xff
      13'h1EE8: dout <= 8'b11111111; // 7912 : 255 - 0xff
      13'h1EE9: dout <= 8'b11111111; // 7913 : 255 - 0xff
      13'h1EEA: dout <= 8'b11111111; // 7914 : 255 - 0xff
      13'h1EEB: dout <= 8'b11111111; // 7915 : 255 - 0xff
      13'h1EEC: dout <= 8'b11111111; // 7916 : 255 - 0xff
      13'h1EED: dout <= 8'b11111111; // 7917 : 255 - 0xff
      13'h1EEE: dout <= 8'b11111111; // 7918 : 255 - 0xff
      13'h1EEF: dout <= 8'b11111111; // 7919 : 255 - 0xff
      13'h1EF0: dout <= 8'b11111111; // 7920 : 255 - 0xff -- Background 0xef
      13'h1EF1: dout <= 8'b11111111; // 7921 : 255 - 0xff
      13'h1EF2: dout <= 8'b11111111; // 7922 : 255 - 0xff
      13'h1EF3: dout <= 8'b11111111; // 7923 : 255 - 0xff
      13'h1EF4: dout <= 8'b11111111; // 7924 : 255 - 0xff
      13'h1EF5: dout <= 8'b11111111; // 7925 : 255 - 0xff
      13'h1EF6: dout <= 8'b11111111; // 7926 : 255 - 0xff
      13'h1EF7: dout <= 8'b11111111; // 7927 : 255 - 0xff
      13'h1EF8: dout <= 8'b11111111; // 7928 : 255 - 0xff
      13'h1EF9: dout <= 8'b11111111; // 7929 : 255 - 0xff
      13'h1EFA: dout <= 8'b11111111; // 7930 : 255 - 0xff
      13'h1EFB: dout <= 8'b11111111; // 7931 : 255 - 0xff
      13'h1EFC: dout <= 8'b11111111; // 7932 : 255 - 0xff
      13'h1EFD: dout <= 8'b11111111; // 7933 : 255 - 0xff
      13'h1EFE: dout <= 8'b11111111; // 7934 : 255 - 0xff
      13'h1EFF: dout <= 8'b11111111; // 7935 : 255 - 0xff
      13'h1F00: dout <= 8'b11111111; // 7936 : 255 - 0xff -- Background 0xf0
      13'h1F01: dout <= 8'b11111111; // 7937 : 255 - 0xff
      13'h1F02: dout <= 8'b11111111; // 7938 : 255 - 0xff
      13'h1F03: dout <= 8'b11111111; // 7939 : 255 - 0xff
      13'h1F04: dout <= 8'b11111111; // 7940 : 255 - 0xff
      13'h1F05: dout <= 8'b11111111; // 7941 : 255 - 0xff
      13'h1F06: dout <= 8'b11111111; // 7942 : 255 - 0xff
      13'h1F07: dout <= 8'b11111111; // 7943 : 255 - 0xff
      13'h1F08: dout <= 8'b11111111; // 7944 : 255 - 0xff
      13'h1F09: dout <= 8'b11111111; // 7945 : 255 - 0xff
      13'h1F0A: dout <= 8'b11111111; // 7946 : 255 - 0xff
      13'h1F0B: dout <= 8'b11111111; // 7947 : 255 - 0xff
      13'h1F0C: dout <= 8'b11111111; // 7948 : 255 - 0xff
      13'h1F0D: dout <= 8'b11111111; // 7949 : 255 - 0xff
      13'h1F0E: dout <= 8'b11111111; // 7950 : 255 - 0xff
      13'h1F0F: dout <= 8'b11111111; // 7951 : 255 - 0xff
      13'h1F10: dout <= 8'b11111111; // 7952 : 255 - 0xff -- Background 0xf1
      13'h1F11: dout <= 8'b11111111; // 7953 : 255 - 0xff
      13'h1F12: dout <= 8'b11111111; // 7954 : 255 - 0xff
      13'h1F13: dout <= 8'b11111111; // 7955 : 255 - 0xff
      13'h1F14: dout <= 8'b11111111; // 7956 : 255 - 0xff
      13'h1F15: dout <= 8'b11111111; // 7957 : 255 - 0xff
      13'h1F16: dout <= 8'b11111111; // 7958 : 255 - 0xff
      13'h1F17: dout <= 8'b11111111; // 7959 : 255 - 0xff
      13'h1F18: dout <= 8'b11111111; // 7960 : 255 - 0xff
      13'h1F19: dout <= 8'b11111111; // 7961 : 255 - 0xff
      13'h1F1A: dout <= 8'b11111111; // 7962 : 255 - 0xff
      13'h1F1B: dout <= 8'b11111111; // 7963 : 255 - 0xff
      13'h1F1C: dout <= 8'b11111111; // 7964 : 255 - 0xff
      13'h1F1D: dout <= 8'b11111111; // 7965 : 255 - 0xff
      13'h1F1E: dout <= 8'b11111111; // 7966 : 255 - 0xff
      13'h1F1F: dout <= 8'b11111111; // 7967 : 255 - 0xff
      13'h1F20: dout <= 8'b11111111; // 7968 : 255 - 0xff -- Background 0xf2
      13'h1F21: dout <= 8'b11111111; // 7969 : 255 - 0xff
      13'h1F22: dout <= 8'b11111111; // 7970 : 255 - 0xff
      13'h1F23: dout <= 8'b11111111; // 7971 : 255 - 0xff
      13'h1F24: dout <= 8'b11111111; // 7972 : 255 - 0xff
      13'h1F25: dout <= 8'b11111111; // 7973 : 255 - 0xff
      13'h1F26: dout <= 8'b11111111; // 7974 : 255 - 0xff
      13'h1F27: dout <= 8'b11111111; // 7975 : 255 - 0xff
      13'h1F28: dout <= 8'b11111111; // 7976 : 255 - 0xff
      13'h1F29: dout <= 8'b11111111; // 7977 : 255 - 0xff
      13'h1F2A: dout <= 8'b11111111; // 7978 : 255 - 0xff
      13'h1F2B: dout <= 8'b11111111; // 7979 : 255 - 0xff
      13'h1F2C: dout <= 8'b11111111; // 7980 : 255 - 0xff
      13'h1F2D: dout <= 8'b11111111; // 7981 : 255 - 0xff
      13'h1F2E: dout <= 8'b11111111; // 7982 : 255 - 0xff
      13'h1F2F: dout <= 8'b11111111; // 7983 : 255 - 0xff
      13'h1F30: dout <= 8'b11111111; // 7984 : 255 - 0xff -- Background 0xf3
      13'h1F31: dout <= 8'b11111111; // 7985 : 255 - 0xff
      13'h1F32: dout <= 8'b11111111; // 7986 : 255 - 0xff
      13'h1F33: dout <= 8'b11111111; // 7987 : 255 - 0xff
      13'h1F34: dout <= 8'b11111111; // 7988 : 255 - 0xff
      13'h1F35: dout <= 8'b11111111; // 7989 : 255 - 0xff
      13'h1F36: dout <= 8'b11111111; // 7990 : 255 - 0xff
      13'h1F37: dout <= 8'b11111111; // 7991 : 255 - 0xff
      13'h1F38: dout <= 8'b11111111; // 7992 : 255 - 0xff
      13'h1F39: dout <= 8'b11111111; // 7993 : 255 - 0xff
      13'h1F3A: dout <= 8'b11111111; // 7994 : 255 - 0xff
      13'h1F3B: dout <= 8'b11111111; // 7995 : 255 - 0xff
      13'h1F3C: dout <= 8'b11111111; // 7996 : 255 - 0xff
      13'h1F3D: dout <= 8'b11111111; // 7997 : 255 - 0xff
      13'h1F3E: dout <= 8'b11111111; // 7998 : 255 - 0xff
      13'h1F3F: dout <= 8'b11111111; // 7999 : 255 - 0xff
      13'h1F40: dout <= 8'b11111111; // 8000 : 255 - 0xff -- Background 0xf4
      13'h1F41: dout <= 8'b11111111; // 8001 : 255 - 0xff
      13'h1F42: dout <= 8'b11111111; // 8002 : 255 - 0xff
      13'h1F43: dout <= 8'b11111111; // 8003 : 255 - 0xff
      13'h1F44: dout <= 8'b11111111; // 8004 : 255 - 0xff
      13'h1F45: dout <= 8'b11111111; // 8005 : 255 - 0xff
      13'h1F46: dout <= 8'b11111111; // 8006 : 255 - 0xff
      13'h1F47: dout <= 8'b11111111; // 8007 : 255 - 0xff
      13'h1F48: dout <= 8'b11111111; // 8008 : 255 - 0xff
      13'h1F49: dout <= 8'b11111111; // 8009 : 255 - 0xff
      13'h1F4A: dout <= 8'b11111111; // 8010 : 255 - 0xff
      13'h1F4B: dout <= 8'b11111111; // 8011 : 255 - 0xff
      13'h1F4C: dout <= 8'b11111111; // 8012 : 255 - 0xff
      13'h1F4D: dout <= 8'b11111111; // 8013 : 255 - 0xff
      13'h1F4E: dout <= 8'b11111111; // 8014 : 255 - 0xff
      13'h1F4F: dout <= 8'b11111111; // 8015 : 255 - 0xff
      13'h1F50: dout <= 8'b11111111; // 8016 : 255 - 0xff -- Background 0xf5
      13'h1F51: dout <= 8'b11111111; // 8017 : 255 - 0xff
      13'h1F52: dout <= 8'b11111111; // 8018 : 255 - 0xff
      13'h1F53: dout <= 8'b11111111; // 8019 : 255 - 0xff
      13'h1F54: dout <= 8'b11111111; // 8020 : 255 - 0xff
      13'h1F55: dout <= 8'b11111111; // 8021 : 255 - 0xff
      13'h1F56: dout <= 8'b11111111; // 8022 : 255 - 0xff
      13'h1F57: dout <= 8'b11111111; // 8023 : 255 - 0xff
      13'h1F58: dout <= 8'b11111111; // 8024 : 255 - 0xff
      13'h1F59: dout <= 8'b11111111; // 8025 : 255 - 0xff
      13'h1F5A: dout <= 8'b11111111; // 8026 : 255 - 0xff
      13'h1F5B: dout <= 8'b11111111; // 8027 : 255 - 0xff
      13'h1F5C: dout <= 8'b11111111; // 8028 : 255 - 0xff
      13'h1F5D: dout <= 8'b11111111; // 8029 : 255 - 0xff
      13'h1F5E: dout <= 8'b11111111; // 8030 : 255 - 0xff
      13'h1F5F: dout <= 8'b11111111; // 8031 : 255 - 0xff
      13'h1F60: dout <= 8'b11111111; // 8032 : 255 - 0xff -- Background 0xf6
      13'h1F61: dout <= 8'b11111111; // 8033 : 255 - 0xff
      13'h1F62: dout <= 8'b11111111; // 8034 : 255 - 0xff
      13'h1F63: dout <= 8'b11111111; // 8035 : 255 - 0xff
      13'h1F64: dout <= 8'b11111111; // 8036 : 255 - 0xff
      13'h1F65: dout <= 8'b11111111; // 8037 : 255 - 0xff
      13'h1F66: dout <= 8'b11111111; // 8038 : 255 - 0xff
      13'h1F67: dout <= 8'b11111111; // 8039 : 255 - 0xff
      13'h1F68: dout <= 8'b11111111; // 8040 : 255 - 0xff
      13'h1F69: dout <= 8'b11111111; // 8041 : 255 - 0xff
      13'h1F6A: dout <= 8'b11111111; // 8042 : 255 - 0xff
      13'h1F6B: dout <= 8'b11111111; // 8043 : 255 - 0xff
      13'h1F6C: dout <= 8'b11111111; // 8044 : 255 - 0xff
      13'h1F6D: dout <= 8'b11111111; // 8045 : 255 - 0xff
      13'h1F6E: dout <= 8'b11111111; // 8046 : 255 - 0xff
      13'h1F6F: dout <= 8'b11111111; // 8047 : 255 - 0xff
      13'h1F70: dout <= 8'b11111111; // 8048 : 255 - 0xff -- Background 0xf7
      13'h1F71: dout <= 8'b11111111; // 8049 : 255 - 0xff
      13'h1F72: dout <= 8'b11111111; // 8050 : 255 - 0xff
      13'h1F73: dout <= 8'b11111111; // 8051 : 255 - 0xff
      13'h1F74: dout <= 8'b11111111; // 8052 : 255 - 0xff
      13'h1F75: dout <= 8'b11111111; // 8053 : 255 - 0xff
      13'h1F76: dout <= 8'b11111111; // 8054 : 255 - 0xff
      13'h1F77: dout <= 8'b11111111; // 8055 : 255 - 0xff
      13'h1F78: dout <= 8'b11111111; // 8056 : 255 - 0xff
      13'h1F79: dout <= 8'b11111111; // 8057 : 255 - 0xff
      13'h1F7A: dout <= 8'b11111111; // 8058 : 255 - 0xff
      13'h1F7B: dout <= 8'b11111111; // 8059 : 255 - 0xff
      13'h1F7C: dout <= 8'b11111111; // 8060 : 255 - 0xff
      13'h1F7D: dout <= 8'b11111111; // 8061 : 255 - 0xff
      13'h1F7E: dout <= 8'b11111111; // 8062 : 255 - 0xff
      13'h1F7F: dout <= 8'b11111111; // 8063 : 255 - 0xff
      13'h1F80: dout <= 8'b11111111; // 8064 : 255 - 0xff -- Background 0xf8
      13'h1F81: dout <= 8'b11111111; // 8065 : 255 - 0xff
      13'h1F82: dout <= 8'b11111111; // 8066 : 255 - 0xff
      13'h1F83: dout <= 8'b11111111; // 8067 : 255 - 0xff
      13'h1F84: dout <= 8'b11111111; // 8068 : 255 - 0xff
      13'h1F85: dout <= 8'b11111111; // 8069 : 255 - 0xff
      13'h1F86: dout <= 8'b11111111; // 8070 : 255 - 0xff
      13'h1F87: dout <= 8'b11111111; // 8071 : 255 - 0xff
      13'h1F88: dout <= 8'b11111111; // 8072 : 255 - 0xff
      13'h1F89: dout <= 8'b11111111; // 8073 : 255 - 0xff
      13'h1F8A: dout <= 8'b11111111; // 8074 : 255 - 0xff
      13'h1F8B: dout <= 8'b11111111; // 8075 : 255 - 0xff
      13'h1F8C: dout <= 8'b11111111; // 8076 : 255 - 0xff
      13'h1F8D: dout <= 8'b11111111; // 8077 : 255 - 0xff
      13'h1F8E: dout <= 8'b11111111; // 8078 : 255 - 0xff
      13'h1F8F: dout <= 8'b11111111; // 8079 : 255 - 0xff
      13'h1F90: dout <= 8'b11111111; // 8080 : 255 - 0xff -- Background 0xf9
      13'h1F91: dout <= 8'b11111111; // 8081 : 255 - 0xff
      13'h1F92: dout <= 8'b11111111; // 8082 : 255 - 0xff
      13'h1F93: dout <= 8'b11111111; // 8083 : 255 - 0xff
      13'h1F94: dout <= 8'b11111111; // 8084 : 255 - 0xff
      13'h1F95: dout <= 8'b11111111; // 8085 : 255 - 0xff
      13'h1F96: dout <= 8'b11111111; // 8086 : 255 - 0xff
      13'h1F97: dout <= 8'b11111111; // 8087 : 255 - 0xff
      13'h1F98: dout <= 8'b11111111; // 8088 : 255 - 0xff
      13'h1F99: dout <= 8'b11111111; // 8089 : 255 - 0xff
      13'h1F9A: dout <= 8'b11111111; // 8090 : 255 - 0xff
      13'h1F9B: dout <= 8'b11111111; // 8091 : 255 - 0xff
      13'h1F9C: dout <= 8'b11111111; // 8092 : 255 - 0xff
      13'h1F9D: dout <= 8'b11111111; // 8093 : 255 - 0xff
      13'h1F9E: dout <= 8'b11111111; // 8094 : 255 - 0xff
      13'h1F9F: dout <= 8'b11111111; // 8095 : 255 - 0xff
      13'h1FA0: dout <= 8'b11111111; // 8096 : 255 - 0xff -- Background 0xfa
      13'h1FA1: dout <= 8'b11111111; // 8097 : 255 - 0xff
      13'h1FA2: dout <= 8'b11111111; // 8098 : 255 - 0xff
      13'h1FA3: dout <= 8'b11111111; // 8099 : 255 - 0xff
      13'h1FA4: dout <= 8'b11111111; // 8100 : 255 - 0xff
      13'h1FA5: dout <= 8'b11111111; // 8101 : 255 - 0xff
      13'h1FA6: dout <= 8'b11111111; // 8102 : 255 - 0xff
      13'h1FA7: dout <= 8'b11111111; // 8103 : 255 - 0xff
      13'h1FA8: dout <= 8'b11111111; // 8104 : 255 - 0xff
      13'h1FA9: dout <= 8'b11111111; // 8105 : 255 - 0xff
      13'h1FAA: dout <= 8'b11111111; // 8106 : 255 - 0xff
      13'h1FAB: dout <= 8'b11111111; // 8107 : 255 - 0xff
      13'h1FAC: dout <= 8'b11111111; // 8108 : 255 - 0xff
      13'h1FAD: dout <= 8'b11111111; // 8109 : 255 - 0xff
      13'h1FAE: dout <= 8'b11111111; // 8110 : 255 - 0xff
      13'h1FAF: dout <= 8'b11111111; // 8111 : 255 - 0xff
      13'h1FB0: dout <= 8'b11111111; // 8112 : 255 - 0xff -- Background 0xfb
      13'h1FB1: dout <= 8'b11111111; // 8113 : 255 - 0xff
      13'h1FB2: dout <= 8'b11111111; // 8114 : 255 - 0xff
      13'h1FB3: dout <= 8'b11111111; // 8115 : 255 - 0xff
      13'h1FB4: dout <= 8'b11111111; // 8116 : 255 - 0xff
      13'h1FB5: dout <= 8'b11111111; // 8117 : 255 - 0xff
      13'h1FB6: dout <= 8'b11111111; // 8118 : 255 - 0xff
      13'h1FB7: dout <= 8'b11111111; // 8119 : 255 - 0xff
      13'h1FB8: dout <= 8'b11111111; // 8120 : 255 - 0xff
      13'h1FB9: dout <= 8'b11111111; // 8121 : 255 - 0xff
      13'h1FBA: dout <= 8'b11111111; // 8122 : 255 - 0xff
      13'h1FBB: dout <= 8'b11111111; // 8123 : 255 - 0xff
      13'h1FBC: dout <= 8'b11111111; // 8124 : 255 - 0xff
      13'h1FBD: dout <= 8'b11111111; // 8125 : 255 - 0xff
      13'h1FBE: dout <= 8'b11111111; // 8126 : 255 - 0xff
      13'h1FBF: dout <= 8'b11111111; // 8127 : 255 - 0xff
      13'h1FC0: dout <= 8'b11111111; // 8128 : 255 - 0xff -- Background 0xfc
      13'h1FC1: dout <= 8'b11111111; // 8129 : 255 - 0xff
      13'h1FC2: dout <= 8'b11111111; // 8130 : 255 - 0xff
      13'h1FC3: dout <= 8'b11111111; // 8131 : 255 - 0xff
      13'h1FC4: dout <= 8'b11111111; // 8132 : 255 - 0xff
      13'h1FC5: dout <= 8'b11111111; // 8133 : 255 - 0xff
      13'h1FC6: dout <= 8'b11111111; // 8134 : 255 - 0xff
      13'h1FC7: dout <= 8'b11111111; // 8135 : 255 - 0xff
      13'h1FC8: dout <= 8'b11111111; // 8136 : 255 - 0xff
      13'h1FC9: dout <= 8'b11111111; // 8137 : 255 - 0xff
      13'h1FCA: dout <= 8'b11111111; // 8138 : 255 - 0xff
      13'h1FCB: dout <= 8'b11111111; // 8139 : 255 - 0xff
      13'h1FCC: dout <= 8'b11111111; // 8140 : 255 - 0xff
      13'h1FCD: dout <= 8'b11111111; // 8141 : 255 - 0xff
      13'h1FCE: dout <= 8'b11111111; // 8142 : 255 - 0xff
      13'h1FCF: dout <= 8'b11111111; // 8143 : 255 - 0xff
      13'h1FD0: dout <= 8'b11111111; // 8144 : 255 - 0xff -- Background 0xfd
      13'h1FD1: dout <= 8'b11111111; // 8145 : 255 - 0xff
      13'h1FD2: dout <= 8'b11111111; // 8146 : 255 - 0xff
      13'h1FD3: dout <= 8'b11111111; // 8147 : 255 - 0xff
      13'h1FD4: dout <= 8'b11111111; // 8148 : 255 - 0xff
      13'h1FD5: dout <= 8'b11111111; // 8149 : 255 - 0xff
      13'h1FD6: dout <= 8'b11111111; // 8150 : 255 - 0xff
      13'h1FD7: dout <= 8'b11111111; // 8151 : 255 - 0xff
      13'h1FD8: dout <= 8'b11111111; // 8152 : 255 - 0xff
      13'h1FD9: dout <= 8'b11111111; // 8153 : 255 - 0xff
      13'h1FDA: dout <= 8'b11111111; // 8154 : 255 - 0xff
      13'h1FDB: dout <= 8'b11111111; // 8155 : 255 - 0xff
      13'h1FDC: dout <= 8'b11111111; // 8156 : 255 - 0xff
      13'h1FDD: dout <= 8'b11111111; // 8157 : 255 - 0xff
      13'h1FDE: dout <= 8'b11111111; // 8158 : 255 - 0xff
      13'h1FDF: dout <= 8'b11111111; // 8159 : 255 - 0xff
      13'h1FE0: dout <= 8'b11111111; // 8160 : 255 - 0xff -- Background 0xfe
      13'h1FE1: dout <= 8'b11111111; // 8161 : 255 - 0xff
      13'h1FE2: dout <= 8'b11111111; // 8162 : 255 - 0xff
      13'h1FE3: dout <= 8'b11111111; // 8163 : 255 - 0xff
      13'h1FE4: dout <= 8'b11111111; // 8164 : 255 - 0xff
      13'h1FE5: dout <= 8'b11111111; // 8165 : 255 - 0xff
      13'h1FE6: dout <= 8'b11111111; // 8166 : 255 - 0xff
      13'h1FE7: dout <= 8'b11111111; // 8167 : 255 - 0xff
      13'h1FE8: dout <= 8'b11111111; // 8168 : 255 - 0xff
      13'h1FE9: dout <= 8'b11111111; // 8169 : 255 - 0xff
      13'h1FEA: dout <= 8'b11111111; // 8170 : 255 - 0xff
      13'h1FEB: dout <= 8'b11111111; // 8171 : 255 - 0xff
      13'h1FEC: dout <= 8'b11111111; // 8172 : 255 - 0xff
      13'h1FED: dout <= 8'b11111111; // 8173 : 255 - 0xff
      13'h1FEE: dout <= 8'b11111111; // 8174 : 255 - 0xff
      13'h1FEF: dout <= 8'b11111111; // 8175 : 255 - 0xff
      13'h1FF0: dout <= 8'b11111111; // 8176 : 255 - 0xff -- Background 0xff
      13'h1FF1: dout <= 8'b11111111; // 8177 : 255 - 0xff
      13'h1FF2: dout <= 8'b11111111; // 8178 : 255 - 0xff
      13'h1FF3: dout <= 8'b11111111; // 8179 : 255 - 0xff
      13'h1FF4: dout <= 8'b11111111; // 8180 : 255 - 0xff
      13'h1FF5: dout <= 8'b11111111; // 8181 : 255 - 0xff
      13'h1FF6: dout <= 8'b11111111; // 8182 : 255 - 0xff
      13'h1FF7: dout <= 8'b11111111; // 8183 : 255 - 0xff
      13'h1FF8: dout <= 8'b11111111; // 8184 : 255 - 0xff
      13'h1FF9: dout <= 8'b11111111; // 8185 : 255 - 0xff
      13'h1FFA: dout <= 8'b11111111; // 8186 : 255 - 0xff
      13'h1FFB: dout <= 8'b11111111; // 8187 : 255 - 0xff
      13'h1FFC: dout <= 8'b11111111; // 8188 : 255 - 0xff
      13'h1FFD: dout <= 8'b11111111; // 8189 : 255 - 0xff
      13'h1FFE: dout <= 8'b11111111; // 8190 : 255 - 0xff
      13'h1FFF: dout <= 8'b11111111; // 8191 : 255 - 0xff
    endcase
  end

endmodule
