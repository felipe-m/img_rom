--- Autcmatically generated VHDL ROM from a NES memory file----
---   SPRITEs MEMORY (OAM)
-- https://wiki.nesdev.com/w/index.php/PPU_OAM


---  Original memory dump file name: smario_traspas_oam.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_OAM_SMARIO_TRASPAS is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(8-1 downto 0);  --256 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_OAM_SMARIO_TRASPAS;

architecture BEHAVIORAL of ROM_OAM_SMARIO_TRASPAS is
  signal addr_int  : natural range 0 to 2**8-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
    "00011000", --    0 -  0x0  :   24 - 0x18 -- Sprite 0x0
    "11111111", --    1 -  0x1  :  255 - 0xff
    "00100011", --    2 -  0x2  :   35 - 0x23
    "01011000", --    3 -  0x3  :   88 - 0x58
    "10110000", --    4 -  0x4  :  176 - 0xb0 -- Sprite 0x1
    "11111100", --    5 -  0x5  :  252 - 0xfc
    "00000000", --    6 -  0x6  :    0 - 0x0
    "01110000", --    7 -  0x7  :  112 - 0x70
    "10110000", --    8 -  0x8  :  176 - 0xb0 -- Sprite 0x2
    "11111100", --    9 -  0x9  :  252 - 0xfc
    "00000000", --   10 -  0xa  :    0 - 0x0
    "01111000", --   11 -  0xb  :  120 - 0x78
    "10111000", --   12 -  0xc  :  184 - 0xb8 -- Sprite 0x3
    "11111100", --   13 -  0xd  :  252 - 0xfc
    "00000000", --   14 -  0xe  :    0 - 0x0
    "01110000", --   15 -  0xf  :  112 - 0x70
    "10111000", --   16 - 0x10  :  184 - 0xb8 -- Sprite 0x4
    "11111100", --   17 - 0x11  :  252 - 0xfc
    "00000000", --   18 - 0x12  :    0 - 0x0
    "01111000", --   19 - 0x13  :  120 - 0x78
    "11000000", --   20 - 0x14  :  192 - 0xc0 -- Sprite 0x5
    "00111010", --   21 - 0x15  :   58 - 0x3a
    "00000000", --   22 - 0x16  :    0 - 0x0
    "01110000", --   23 - 0x17  :  112 - 0x70
    "11000000", --   24 - 0x18  :  192 - 0xc0 -- Sprite 0x6
    "00110111", --   25 - 0x19  :   55 - 0x37
    "00000000", --   26 - 0x1a  :    0 - 0x0
    "01111000", --   27 - 0x1b  :  120 - 0x78
    "11001000", --   28 - 0x1c  :  200 - 0xc8 -- Sprite 0x7
    "01001111", --   29 - 0x1d  :   79 - 0x4f
    "00000000", --   30 - 0x1e  :    0 - 0x0
    "01110000", --   31 - 0x1f  :  112 - 0x70
    "11001000", --   32 - 0x20  :  200 - 0xc8 -- Sprite 0x8
    "01001111", --   33 - 0x21  :   79 - 0x4f
    "01000000", --   34 - 0x22  :   64 - 0x40
    "01111000", --   35 - 0x23  :  120 - 0x78
    "11111000", --   36 - 0x24  :  248 - 0xf8 -- Sprite 0x9
    "00000000", --   37 - 0x25  :    0 - 0x0
    "00000000", --   38 - 0x26  :    0 - 0x0
    "00000000", --   39 - 0x27  :    0 - 0x0
    "11111000", --   40 - 0x28  :  248 - 0xf8 -- Sprite 0xa
    "11111100", --   41 - 0x29  :  252 - 0xfc
    "00000001", --   42 - 0x2a  :    1 - 0x1
    "01000010", --   43 - 0x2b  :   66 - 0x42
    "11111000", --   44 - 0x2c  :  248 - 0xf8 -- Sprite 0xb
    "11111100", --   45 - 0x2d  :  252 - 0xfc
    "01000001", --   46 - 0x2e  :   65 - 0x41
    "01001010", --   47 - 0x2f  :   74 - 0x4a
    "11111000", --   48 - 0x30  :  248 - 0xf8 -- Sprite 0xc
    "01101111", --   49 - 0x31  :  111 - 0x6f
    "10000001", --   50 - 0x32  :  129 - 0x81
    "01000010", --   51 - 0x33  :   66 - 0x42
    "11111000", --   52 - 0x34  :  248 - 0xf8 -- Sprite 0xd
    "01101111", --   53 - 0x35  :  111 - 0x6f
    "11000001", --   54 - 0x36  :  193 - 0xc1
    "01001010", --   55 - 0x37  :   74 - 0x4a
    "11111000", --   56 - 0x38  :  248 - 0xf8 -- Sprite 0xe
    "01101110", --   57 - 0x39  :  110 - 0x6e
    "10000001", --   58 - 0x3a  :  129 - 0x81
    "01000010", --   59 - 0x3b  :   66 - 0x42
    "11111000", --   60 - 0x3c  :  248 - 0xf8 -- Sprite 0xf
    "01101110", --   61 - 0x3d  :  110 - 0x6e
    "11000001", --   62 - 0x3e  :  193 - 0xc1
    "01001010", --   63 - 0x3f  :   74 - 0x4a
    "11111000", --   64 - 0x40  :  248 - 0xf8 -- Sprite 0x10
    "01110011", --   65 - 0x41  :  115 - 0x73
    "01000011", --   66 - 0x42  :   67 - 0x43
    "10111101", --   67 - 0x43  :  189 - 0xbd
    "11111000", --   68 - 0x44  :  248 - 0xf8 -- Sprite 0x11
    "01110010", --   69 - 0x45  :  114 - 0x72
    "01000011", --   70 - 0x46  :   67 - 0x43
    "11000101", --   71 - 0x47  :  197 - 0xc5
    "11111000", --   72 - 0x48  :  248 - 0xf8 -- Sprite 0x12
    "11110110", --   73 - 0x49  :  246 - 0xf6
    "00000010", --   74 - 0x4a  :    2 - 0x2
    "01011000", --   75 - 0x4b  :   88 - 0x58
    "11111000", --   76 - 0x4c  :  248 - 0xf8 -- Sprite 0x13
    "11111011", --   77 - 0x4d  :  251 - 0xfb
    "00000010", --   78 - 0x4e  :    2 - 0x2
    "01100000", --   79 - 0x4f  :   96 - 0x60
    "11111000", --   80 - 0x50  :  248 - 0xf8 -- Sprite 0x14
    "11111100", --   81 - 0x51  :  252 - 0xfc
    "10000011", --   82 - 0x52  :  131 - 0x83
    "00101111", --   83 - 0x53  :   47 - 0x2f
    "11111000", --   84 - 0x54  :  248 - 0xf8 -- Sprite 0x15
    "11111100", --   85 - 0x55  :  252 - 0xfc
    "11000011", --   86 - 0x56  :  195 - 0xc3
    "00110111", --   87 - 0x57  :   55 - 0x37
    "11111000", --   88 - 0x58  :  248 - 0xf8 -- Sprite 0x16
    "11101111", --   89 - 0x59  :  239 - 0xef
    "10000011", --   90 - 0x5a  :  131 - 0x83
    "00101111", --   91 - 0x5b  :   47 - 0x2f
    "11111000", --   92 - 0x5c  :  248 - 0xf8 -- Sprite 0x17
    "11101111", --   93 - 0x5d  :  239 - 0xef
    "11000011", --   94 - 0x5e  :  195 - 0xc3
    "00110111", --   95 - 0x5f  :   55 - 0x37
    "11111000", --   96 - 0x60  :  248 - 0xf8 -- Sprite 0x18
    "11111100", --   97 - 0x61  :  252 - 0xfc
    "00000001", --   98 - 0x62  :    1 - 0x1
    "01000100", --   99 - 0x63  :   68 - 0x44
    "11111000", --  100 - 0x64  :  248 - 0xf8 -- Sprite 0x19
    "11111100", --  101 - 0x65  :  252 - 0xfc
    "01000001", --  102 - 0x66  :   65 - 0x41
    "01001100", --  103 - 0x67  :   76 - 0x4c
    "11111000", --  104 - 0x68  :  248 - 0xf8 -- Sprite 0x1a
    "01101111", --  105 - 0x69  :  111 - 0x6f
    "10000001", --  106 - 0x6a  :  129 - 0x81
    "01000100", --  107 - 0x6b  :   68 - 0x44
    "11111000", --  108 - 0x6c  :  248 - 0xf8 -- Sprite 0x1b
    "01101111", --  109 - 0x6d  :  111 - 0x6f
    "11000001", --  110 - 0x6e  :  193 - 0xc1
    "01001100", --  111 - 0x6f  :   76 - 0x4c
    "11111000", --  112 - 0x70  :  248 - 0xf8 -- Sprite 0x1c
    "01101110", --  113 - 0x71  :  110 - 0x6e
    "10000001", --  114 - 0x72  :  129 - 0x81
    "01000100", --  115 - 0x73  :   68 - 0x44
    "11111000", --  116 - 0x74  :  248 - 0xf8 -- Sprite 0x1d
    "01101110", --  117 - 0x75  :  110 - 0x6e
    "11000001", --  118 - 0x76  :  193 - 0xc1
    "01001100", --  119 - 0x77  :   76 - 0x4c
    "11111000", --  120 - 0x78  :  248 - 0xf8 -- Sprite 0x1e
    "00000000", --  121 - 0x79  :    0 - 0x0
    "00000000", --  122 - 0x7a  :    0 - 0x0
    "00000000", --  123 - 0x7b  :    0 - 0x0
    "11111000", --  124 - 0x7c  :  248 - 0xf8 -- Sprite 0x1f
    "00000000", --  125 - 0x7d  :    0 - 0x0
    "00000000", --  126 - 0x7e  :    0 - 0x0
    "00000000", --  127 - 0x7f  :    0 - 0x0
    "11111000", --  128 - 0x80  :  248 - 0xf8 -- Sprite 0x20
    "00000000", --  129 - 0x81  :    0 - 0x0
    "00000000", --  130 - 0x82  :    0 - 0x0
    "00000000", --  131 - 0x83  :    0 - 0x0
    "11111000", --  132 - 0x84  :  248 - 0xf8 -- Sprite 0x21
    "00000000", --  133 - 0x85  :    0 - 0x0
    "00000000", --  134 - 0x86  :    0 - 0x0
    "00000000", --  135 - 0x87  :    0 - 0x0
    "11111000", --  136 - 0x88  :  248 - 0xf8 -- Sprite 0x22
    "11111100", --  137 - 0x89  :  252 - 0xfc
    "01000011", --  138 - 0x8a  :   67 - 0x43
    "10111110", --  139 - 0x8b  :  190 - 0xbe
    "11111000", --  140 - 0x8c  :  248 - 0xf8 -- Sprite 0x23
    "11111100", --  141 - 0x8d  :  252 - 0xfc
    "01000011", --  142 - 0x8e  :   67 - 0x43
    "11000110", --  143 - 0x8f  :  198 - 0xc6
    "11111000", --  144 - 0x90  :  248 - 0xf8 -- Sprite 0x24
    "01110001", --  145 - 0x91  :  113 - 0x71
    "01000011", --  146 - 0x92  :   67 - 0x43
    "10111110", --  147 - 0x93  :  190 - 0xbe
    "11111000", --  148 - 0x94  :  248 - 0xf8 -- Sprite 0x25
    "01110000", --  149 - 0x95  :  112 - 0x70
    "01000011", --  150 - 0x96  :   67 - 0x43
    "11000110", --  151 - 0x97  :  198 - 0xc6
    "11111000", --  152 - 0x98  :  248 - 0xf8 -- Sprite 0x26
    "01110011", --  153 - 0x99  :  115 - 0x73
    "01000011", --  154 - 0x9a  :   67 - 0x43
    "10111110", --  155 - 0x9b  :  190 - 0xbe
    "11111000", --  156 - 0x9c  :  248 - 0xf8 -- Sprite 0x27
    "01110010", --  157 - 0x9d  :  114 - 0x72
    "01000011", --  158 - 0x9e  :   67 - 0x43
    "11000110", --  159 - 0x9f  :  198 - 0xc6
    "11111000", --  160 - 0xa0  :  248 - 0xf8 -- Sprite 0x28
    "11111100", --  161 - 0xa1  :  252 - 0xfc
    "00000011", --  162 - 0xa2  :    3 - 0x3
    "00101110", --  163 - 0xa3  :   46 - 0x2e
    "11111000", --  164 - 0xa4  :  248 - 0xf8 -- Sprite 0x29
    "11111100", --  165 - 0xa5  :  252 - 0xfc
    "01000011", --  166 - 0xa6  :   67 - 0x43
    "00110110", --  167 - 0xa7  :   54 - 0x36
    "11111000", --  168 - 0xa8  :  248 - 0xf8 -- Sprite 0x2a
    "11111100", --  169 - 0xa9  :  252 - 0xfc
    "10000011", --  170 - 0xaa  :  131 - 0x83
    "00101110", --  171 - 0xab  :   46 - 0x2e
    "11111000", --  172 - 0xac  :  248 - 0xf8 -- Sprite 0x2b
    "11111100", --  173 - 0xad  :  252 - 0xfc
    "11000011", --  174 - 0xae  :  195 - 0xc3
    "00110110", --  175 - 0xaf  :   54 - 0x36
    "11111000", --  176 - 0xb0  :  248 - 0xf8 -- Sprite 0x2c
    "11101111", --  177 - 0xb1  :  239 - 0xef
    "10000011", --  178 - 0xb2  :  131 - 0x83
    "00101110", --  179 - 0xb3  :   46 - 0x2e
    "11111000", --  180 - 0xb4  :  248 - 0xf8 -- Sprite 0x2d
    "11101111", --  181 - 0xb5  :  239 - 0xef
    "11000011", --  182 - 0xb6  :  195 - 0xc3
    "00110110", --  183 - 0xb7  :   54 - 0x36
    "11111000", --  184 - 0xb8  :  248 - 0xf8 -- Sprite 0x2e
    "11111100", --  185 - 0xb9  :  252 - 0xfc
    "00000001", --  186 - 0xba  :    1 - 0x1
    "01000111", --  187 - 0xbb  :   71 - 0x47
    "11111000", --  188 - 0xbc  :  248 - 0xf8 -- Sprite 0x2f
    "11111100", --  189 - 0xbd  :  252 - 0xfc
    "01000001", --  190 - 0xbe  :   65 - 0x41
    "01001111", --  191 - 0xbf  :   79 - 0x4f
    "11111000", --  192 - 0xc0  :  248 - 0xf8 -- Sprite 0x30
    "01101111", --  193 - 0xc1  :  111 - 0x6f
    "10000001", --  194 - 0xc2  :  129 - 0x81
    "01000111", --  195 - 0xc3  :   71 - 0x47
    "11111000", --  196 - 0xc4  :  248 - 0xf8 -- Sprite 0x31
    "01101111", --  197 - 0xc5  :  111 - 0x6f
    "11000001", --  198 - 0xc6  :  193 - 0xc1
    "01001111", --  199 - 0xc7  :   79 - 0x4f
    "11111000", --  200 - 0xc8  :  248 - 0xf8 -- Sprite 0x32
    "01101110", --  201 - 0xc9  :  110 - 0x6e
    "10000001", --  202 - 0xca  :  129 - 0x81
    "01000111", --  203 - 0xcb  :   71 - 0x47
    "11111000", --  204 - 0xcc  :  248 - 0xf8 -- Sprite 0x33
    "01101110", --  205 - 0xcd  :  110 - 0x6e
    "11000001", --  206 - 0xce  :  193 - 0xc1
    "01001111", --  207 - 0xcf  :   79 - 0x4f
    "11111000", --  208 - 0xd0  :  248 - 0xf8 -- Sprite 0x34
    "11111100", --  209 - 0xd1  :  252 - 0xfc
    "01000011", --  210 - 0xd2  :   67 - 0x43
    "10111110", --  211 - 0xd3  :  190 - 0xbe
    "11111000", --  212 - 0xd4  :  248 - 0xf8 -- Sprite 0x35
    "11111100", --  213 - 0xd5  :  252 - 0xfc
    "01000011", --  214 - 0xd6  :   67 - 0x43
    "11000110", --  215 - 0xd7  :  198 - 0xc6
    "11111000", --  216 - 0xd8  :  248 - 0xf8 -- Sprite 0x36
    "01110001", --  217 - 0xd9  :  113 - 0x71
    "01000011", --  218 - 0xda  :   67 - 0x43
    "10111110", --  219 - 0xdb  :  190 - 0xbe
    "11111000", --  220 - 0xdc  :  248 - 0xf8 -- Sprite 0x37
    "01110000", --  221 - 0xdd  :  112 - 0x70
    "01000011", --  222 - 0xde  :   67 - 0x43
    "11000110", --  223 - 0xdf  :  198 - 0xc6
    "11111000", --  224 - 0xe0  :  248 - 0xf8 -- Sprite 0x38
    "01110011", --  225 - 0xe1  :  115 - 0x73
    "01000011", --  226 - 0xe2  :   67 - 0x43
    "10111110", --  227 - 0xe3  :  190 - 0xbe
    "11111000", --  228 - 0xe4  :  248 - 0xf8 -- Sprite 0x39
    "01110010", --  229 - 0xe5  :  114 - 0x72
    "01000011", --  230 - 0xe6  :   67 - 0x43
    "11000110", --  231 - 0xe7  :  198 - 0xc6
    "11111000", --  232 - 0xe8  :  248 - 0xf8 -- Sprite 0x3a
    "11110110", --  233 - 0xe9  :  246 - 0xf6
    "00000010", --  234 - 0xea  :    2 - 0x2
    "01011000", --  235 - 0xeb  :   88 - 0x58
    "11111000", --  236 - 0xec  :  248 - 0xf8 -- Sprite 0x3b
    "11111011", --  237 - 0xed  :  251 - 0xfb
    "00000010", --  238 - 0xee  :    2 - 0x2
    "01100000", --  239 - 0xef  :   96 - 0x60
    "11111000", --  240 - 0xf0  :  248 - 0xf8 -- Sprite 0x3c
    "11111100", --  241 - 0xf1  :  252 - 0xfc
    "10000011", --  242 - 0xf2  :  131 - 0x83
    "00110000", --  243 - 0xf3  :   48 - 0x30
    "11111000", --  244 - 0xf4  :  248 - 0xf8 -- Sprite 0x3d
    "11111100", --  245 - 0xf5  :  252 - 0xfc
    "11000011", --  246 - 0xf6  :  195 - 0xc3
    "00111000", --  247 - 0xf7  :   56 - 0x38
    "11111000", --  248 - 0xf8  :  248 - 0xf8 -- Sprite 0x3e
    "11101111", --  249 - 0xf9  :  239 - 0xef
    "10000011", --  250 - 0xfa  :  131 - 0x83
    "00110000", --  251 - 0xfb  :   48 - 0x30
    "11111000", --  252 - 0xfc  :  248 - 0xf8 -- Sprite 0x3f
    "11101111", --  253 - 0xfd  :  239 - 0xef
    "11000011", --  254 - 0xfe  :  195 - 0xc3
    "00111000"  --  255 - 0xff  :   56 - 0x38
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
