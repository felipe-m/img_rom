//- Autcmatically generated verilog ROM from a NES memory file----


//-  Original memory dump file name: nespalette.pal --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_COLORS
  (
     //input     clk,   // clock
     input      [6-1:0] addr,  //64 memory positions
     output reg  [12-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                                     //  address:   value 
                                     //    dec  : dec - hex(RGB)
      8'h0: dout  = 12'b010001000100; //    0 : 1092 - 0x444
      8'h1: dout  = 12'b000000000101; //    1 :    5 - 0x005
      8'h2: dout  = 12'b000000000111; //    2 :    7 - 0x007
      8'h3: dout  = 12'b000000000111; //    3 :    7 - 0x007
      8'h4: dout  = 12'b001100000100; //    4 :  772 - 0x304
      8'h5: dout  = 12'b010100000000; //    5 : 1280 - 0x500
      8'h6: dout  = 12'b010100000000; //    6 : 1280 - 0x500
      8'h7: dout  = 12'b010000000000; //    7 : 1024 - 0x400
      8'h8: dout  = 12'b000100000000; //    8 :  256 - 0x100
      8'h9: dout  = 12'b000000010000; //    9 :   16 - 0x010
      8'hA: dout  = 12'b000000010000; //   10 :   16 - 0x010
      8'hB: dout  = 12'b000000010000; //   11 :   16 - 0x010
      8'hC: dout  = 12'b000000010010; //   12 :   18 - 0x012
      8'hD: dout  = 12'b000000000000; //   13 :    0 - 0x000
      8'hE: dout  = 12'b000000000000; //   14 :    0 - 0x000
      8'hF: dout  = 12'b000000000000; //   15 :    0 - 0x000
      8'h10: dout  = 12'b100110011001; //   16 : 2457 - 0x999
      8'h11: dout  = 12'b000001001011; //   17 :   75 - 0x04B
      8'h12: dout  = 12'b000000111110; //   18 :   62 - 0x03E
      8'h13: dout  = 12'b010100011101; //   19 : 1309 - 0x51D
      8'h14: dout  = 12'b100100001010; //   20 : 2314 - 0x90A
      8'h15: dout  = 12'b110000000101; //   21 : 3077 - 0xC05
      8'h16: dout  = 12'b110000000000; //   22 : 3072 - 0xC00
      8'h17: dout  = 12'b101000100000; //   23 : 2592 - 0xA20
      8'h18: dout  = 12'b010100110000; //   24 : 1328 - 0x530
      8'h19: dout  = 12'b000001010000; //   25 :   80 - 0x050
      8'h1A: dout  = 12'b000001100000; //   26 :   96 - 0x060
      8'h1B: dout  = 12'b000001100001; //   27 :   97 - 0x061
      8'h1C: dout  = 12'b000001010110; //   28 :   86 - 0x056
      8'h1D: dout  = 12'b000000000000; //   29 :    0 - 0x000
      8'h1E: dout  = 12'b000000000000; //   30 :    0 - 0x000
      8'h1F: dout  = 12'b000000000000; //   31 :    0 - 0x000
      8'h20: dout  = 12'b111111111111; //   32 : 4095 - 0xFFF
      8'h21: dout  = 12'b000110011111; //   33 :  415 - 0x19F
      8'h22: dout  = 12'b010101111111; //   34 : 1407 - 0x57F
      8'h23: dout  = 12'b100101101111; //   35 : 2415 - 0x96F
      8'h24: dout  = 12'b111101101111; //   36 : 3951 - 0xF6F
      8'h25: dout  = 12'b111101101011; //   37 : 3947 - 0xF6B
      8'h26: dout  = 12'b111101110110; //   38 : 3958 - 0xF76
      8'h27: dout  = 12'b111110000001; //   39 : 3969 - 0xF81
      8'h28: dout  = 12'b110010010000; //   40 : 3216 - 0xC90
      8'h29: dout  = 12'b011110110000; //   41 : 1968 - 0x7B0
      8'h2A: dout  = 12'b001011000010; //   42 :  706 - 0x2C2
      8'h2B: dout  = 12'b000011000111; //   43 :  199 - 0x0C7
      8'h2C: dout  = 12'b000010111101; //   44 :  189 - 0x0BD
      8'h2D: dout  = 12'b001000100010; //   45 :  546 - 0x222
      8'h2E: dout  = 12'b000000000000; //   46 :    0 - 0x000
      8'h2F: dout  = 12'b000000000000; //   47 :    0 - 0x000
      8'h30: dout  = 12'b111111111111; //   48 : 4095 - 0xFFF
      8'h31: dout  = 12'b100111011111; //   49 : 2527 - 0x9DF
      8'h32: dout  = 12'b101011001111; //   50 : 2767 - 0xACF
      8'h33: dout  = 12'b110110111111; //   51 : 3519 - 0xDBF
      8'h34: dout  = 12'b111110111111; //   52 : 4031 - 0xFBF
      8'h35: dout  = 12'b111111001110; //   53 : 4046 - 0xFCE
      8'h36: dout  = 12'b111111001011; //   54 : 4043 - 0xFCB
      8'h37: dout  = 12'b111111001001; //   55 : 4041 - 0xFC9
      8'h38: dout  = 12'b111011011000; //   56 : 3800 - 0xED8
      8'h39: dout  = 12'b110011011000; //   57 : 3288 - 0xCD8
      8'h3A: dout  = 12'b101011101010; //   58 : 2794 - 0xAEA
      8'h3B: dout  = 12'b100111101100; //   59 : 2540 - 0x9EC
      8'h3C: dout  = 12'b100111101110; //   60 : 2542 - 0x9EE
      8'h3D: dout  = 12'b101010101010; //   61 : 2730 - 0xAAA
      8'h3E: dout  = 12'b000000000000; //   62 :    0 - 0x000
      8'h3F: dout  = 12'b000000000000; //   63 :    0 - 0x000
    endcase
  end

endmodule
