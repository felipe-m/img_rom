--- Autcmatically generated VHDL ROM from a NES memory file----
---   NAME TABLE
-- https://wiki.nesdev.com/w/index.php/PPU_nametables
--- Only the first Name Table: 1KiB


---  Original memory dump file name: sprilo_introscr.bin --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_NTABLE_SPRILO_INTROSCREEN is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(10-1 downto 0);  --1024 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_NTABLE_SPRILO_INTROSCREEN;

architecture BEHAVIORAL of ROM_NTABLE_SPRILO_INTROSCREEN is
  signal addr_int  : natural range 0 to 2**10-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
     ------- Name Table 0---------
    "11111010", --    0 -  0x0  :  250 - 0xfa -- line 0x0
    "11111010", --    1 -  0x1  :  250 - 0xfa
    "11111010", --    2 -  0x2  :  250 - 0xfa
    "11101010", --    3 -  0x3  :  234 - 0xea
    "11111010", --    4 -  0x4  :  250 - 0xfa
    "11111010", --    5 -  0x5  :  250 - 0xfa
    "11111010", --    6 -  0x6  :  250 - 0xfa
    "11111010", --    7 -  0x7  :  250 - 0xfa
    "11111010", --    8 -  0x8  :  250 - 0xfa
    "11111010", --    9 -  0x9  :  250 - 0xfa
    "11111010", --   10 -  0xa  :  250 - 0xfa
    "11111010", --   11 -  0xb  :  250 - 0xfa
    "11111010", --   12 -  0xc  :  250 - 0xfa
    "11111010", --   13 -  0xd  :  250 - 0xfa
    "11101010", --   14 -  0xe  :  234 - 0xea
    "11111010", --   15 -  0xf  :  250 - 0xfa
    "11111010", --   16 - 0x10  :  250 - 0xfa
    "11111010", --   17 - 0x11  :  250 - 0xfa
    "11111010", --   18 - 0x12  :  250 - 0xfa
    "11111010", --   19 - 0x13  :  250 - 0xfa
    "11111010", --   20 - 0x14  :  250 - 0xfa
    "11111010", --   21 - 0x15  :  250 - 0xfa
    "11111010", --   22 - 0x16  :  250 - 0xfa
    "11111010", --   23 - 0x17  :  250 - 0xfa
    "11111010", --   24 - 0x18  :  250 - 0xfa
    "11111010", --   25 - 0x19  :  250 - 0xfa
    "11111010", --   26 - 0x1a  :  250 - 0xfa
    "11111010", --   27 - 0x1b  :  250 - 0xfa
    "11111010", --   28 - 0x1c  :  250 - 0xfa
    "11111010", --   29 - 0x1d  :  250 - 0xfa
    "11111010", --   30 - 0x1e  :  250 - 0xfa
    "11111010", --   31 - 0x1f  :  250 - 0xfa
    "11111010", --   32 - 0x20  :  250 - 0xfa -- line 0x1
    "11111010", --   33 - 0x21  :  250 - 0xfa
    "11111010", --   34 - 0x22  :  250 - 0xfa
    "11111010", --   35 - 0x23  :  250 - 0xfa
    "11111010", --   36 - 0x24  :  250 - 0xfa
    "11111010", --   37 - 0x25  :  250 - 0xfa
    "11111010", --   38 - 0x26  :  250 - 0xfa
    "11111001", --   39 - 0x27  :  249 - 0xf9
    "11111001", --   40 - 0x28  :  249 - 0xf9
    "11111010", --   41 - 0x29  :  250 - 0xfa
    "11111010", --   42 - 0x2a  :  250 - 0xfa
    "11111010", --   43 - 0x2b  :  250 - 0xfa
    "11111010", --   44 - 0x2c  :  250 - 0xfa
    "11111010", --   45 - 0x2d  :  250 - 0xfa
    "11111010", --   46 - 0x2e  :  250 - 0xfa
    "11111010", --   47 - 0x2f  :  250 - 0xfa
    "11111010", --   48 - 0x30  :  250 - 0xfa
    "11111010", --   49 - 0x31  :  250 - 0xfa
    "11101001", --   50 - 0x32  :  233 - 0xe9
    "11111010", --   51 - 0x33  :  250 - 0xfa
    "11111010", --   52 - 0x34  :  250 - 0xfa
    "11111010", --   53 - 0x35  :  250 - 0xfa
    "11111010", --   54 - 0x36  :  250 - 0xfa
    "11111010", --   55 - 0x37  :  250 - 0xfa
    "11111010", --   56 - 0x38  :  250 - 0xfa
    "11111010", --   57 - 0x39  :  250 - 0xfa
    "11111001", --   58 - 0x3a  :  249 - 0xf9
    "11111010", --   59 - 0x3b  :  250 - 0xfa
    "11111010", --   60 - 0x3c  :  250 - 0xfa
    "11111010", --   61 - 0x3d  :  250 - 0xfa
    "11111010", --   62 - 0x3e  :  250 - 0xfa
    "11111010", --   63 - 0x3f  :  250 - 0xfa
    "11111010", --   64 - 0x40  :  250 - 0xfa -- line 0x2
    "11111010", --   65 - 0x41  :  250 - 0xfa
    "11111010", --   66 - 0x42  :  250 - 0xfa
    "11111010", --   67 - 0x43  :  250 - 0xfa
    "11111010", --   68 - 0x44  :  250 - 0xfa
    "11111010", --   69 - 0x45  :  250 - 0xfa
    "11111010", --   70 - 0x46  :  250 - 0xfa
    "11111010", --   71 - 0x47  :  250 - 0xfa
    "11111010", --   72 - 0x48  :  250 - 0xfa
    "11111010", --   73 - 0x49  :  250 - 0xfa
    "11111010", --   74 - 0x4a  :  250 - 0xfa
    "11111010", --   75 - 0x4b  :  250 - 0xfa
    "11111010", --   76 - 0x4c  :  250 - 0xfa
    "11111010", --   77 - 0x4d  :  250 - 0xfa
    "11111010", --   78 - 0x4e  :  250 - 0xfa
    "11101001", --   79 - 0x4f  :  233 - 0xe9
    "11111010", --   80 - 0x50  :  250 - 0xfa
    "11111010", --   81 - 0x51  :  250 - 0xfa
    "11111010", --   82 - 0x52  :  250 - 0xfa
    "11111010", --   83 - 0x53  :  250 - 0xfa
    "11111010", --   84 - 0x54  :  250 - 0xfa
    "11111010", --   85 - 0x55  :  250 - 0xfa
    "11111010", --   86 - 0x56  :  250 - 0xfa
    "11111010", --   87 - 0x57  :  250 - 0xfa
    "11111010", --   88 - 0x58  :  250 - 0xfa
    "11111010", --   89 - 0x59  :  250 - 0xfa
    "11111010", --   90 - 0x5a  :  250 - 0xfa
    "11111010", --   91 - 0x5b  :  250 - 0xfa
    "11111010", --   92 - 0x5c  :  250 - 0xfa
    "11111010", --   93 - 0x5d  :  250 - 0xfa
    "11111010", --   94 - 0x5e  :  250 - 0xfa
    "11111010", --   95 - 0x5f  :  250 - 0xfa
    "11111011", --   96 - 0x60  :  251 - 0xfb -- line 0x3
    "11111011", --   97 - 0x61  :  251 - 0xfb
    "11111011", --   98 - 0x62  :  251 - 0xfb
    "11111011", --   99 - 0x63  :  251 - 0xfb
    "11111011", --  100 - 0x64  :  251 - 0xfb
    "11111011", --  101 - 0x65  :  251 - 0xfb
    "11111011", --  102 - 0x66  :  251 - 0xfb
    "11111011", --  103 - 0x67  :  251 - 0xfb
    "11111011", --  104 - 0x68  :  251 - 0xfb
    "11111011", --  105 - 0x69  :  251 - 0xfb
    "11111011", --  106 - 0x6a  :  251 - 0xfb
    "11111011", --  107 - 0x6b  :  251 - 0xfb
    "11111011", --  108 - 0x6c  :  251 - 0xfb
    "11111011", --  109 - 0x6d  :  251 - 0xfb
    "11111011", --  110 - 0x6e  :  251 - 0xfb
    "11111011", --  111 - 0x6f  :  251 - 0xfb
    "11111011", --  112 - 0x70  :  251 - 0xfb
    "11111011", --  113 - 0x71  :  251 - 0xfb
    "11111011", --  114 - 0x72  :  251 - 0xfb
    "11111011", --  115 - 0x73  :  251 - 0xfb
    "11111011", --  116 - 0x74  :  251 - 0xfb
    "11111011", --  117 - 0x75  :  251 - 0xfb
    "11111011", --  118 - 0x76  :  251 - 0xfb
    "11111011", --  119 - 0x77  :  251 - 0xfb
    "11111011", --  120 - 0x78  :  251 - 0xfb
    "11111011", --  121 - 0x79  :  251 - 0xfb
    "11111011", --  122 - 0x7a  :  251 - 0xfb
    "11111011", --  123 - 0x7b  :  251 - 0xfb
    "11111011", --  124 - 0x7c  :  251 - 0xfb
    "11111011", --  125 - 0x7d  :  251 - 0xfb
    "11111011", --  126 - 0x7e  :  251 - 0xfb
    "11111011", --  127 - 0x7f  :  251 - 0xfb
    "11111111", --  128 - 0x80  :  255 - 0xff -- line 0x4
    "11111111", --  129 - 0x81  :  255 - 0xff
    "11111111", --  130 - 0x82  :  255 - 0xff
    "11111111", --  131 - 0x83  :  255 - 0xff
    "11111111", --  132 - 0x84  :  255 - 0xff
    "11111111", --  133 - 0x85  :  255 - 0xff
    "11111111", --  134 - 0x86  :  255 - 0xff
    "11111111", --  135 - 0x87  :  255 - 0xff
    "11111111", --  136 - 0x88  :  255 - 0xff
    "11111111", --  137 - 0x89  :  255 - 0xff
    "11111111", --  138 - 0x8a  :  255 - 0xff
    "11111111", --  139 - 0x8b  :  255 - 0xff
    "11111111", --  140 - 0x8c  :  255 - 0xff
    "11111111", --  141 - 0x8d  :  255 - 0xff
    "11111111", --  142 - 0x8e  :  255 - 0xff
    "11111111", --  143 - 0x8f  :  255 - 0xff
    "11111111", --  144 - 0x90  :  255 - 0xff
    "11111111", --  145 - 0x91  :  255 - 0xff
    "11111111", --  146 - 0x92  :  255 - 0xff
    "11111111", --  147 - 0x93  :  255 - 0xff
    "11111111", --  148 - 0x94  :  255 - 0xff
    "11111111", --  149 - 0x95  :  255 - 0xff
    "11111111", --  150 - 0x96  :  255 - 0xff
    "11111111", --  151 - 0x97  :  255 - 0xff
    "11111111", --  152 - 0x98  :  255 - 0xff
    "11111111", --  153 - 0x99  :  255 - 0xff
    "11111111", --  154 - 0x9a  :  255 - 0xff
    "11111111", --  155 - 0x9b  :  255 - 0xff
    "11111111", --  156 - 0x9c  :  255 - 0xff
    "11111111", --  157 - 0x9d  :  255 - 0xff
    "11111111", --  158 - 0x9e  :  255 - 0xff
    "11111111", --  159 - 0x9f  :  255 - 0xff
    "11111111", --  160 - 0xa0  :  255 - 0xff -- line 0x5
    "11111101", --  161 - 0xa1  :  253 - 0xfd
    "11111111", --  162 - 0xa2  :  255 - 0xff
    "11111101", --  163 - 0xa3  :  253 - 0xfd
    "11111111", --  164 - 0xa4  :  255 - 0xff
    "11111101", --  165 - 0xa5  :  253 - 0xfd
    "11111111", --  166 - 0xa6  :  255 - 0xff
    "11111101", --  167 - 0xa7  :  253 - 0xfd
    "11111111", --  168 - 0xa8  :  255 - 0xff
    "11111101", --  169 - 0xa9  :  253 - 0xfd
    "11111111", --  170 - 0xaa  :  255 - 0xff
    "11111101", --  171 - 0xab  :  253 - 0xfd
    "11111111", --  172 - 0xac  :  255 - 0xff
    "11111101", --  173 - 0xad  :  253 - 0xfd
    "11111111", --  174 - 0xae  :  255 - 0xff
    "11111101", --  175 - 0xaf  :  253 - 0xfd
    "11111111", --  176 - 0xb0  :  255 - 0xff
    "11111101", --  177 - 0xb1  :  253 - 0xfd
    "11111111", --  178 - 0xb2  :  255 - 0xff
    "11111101", --  179 - 0xb3  :  253 - 0xfd
    "11111111", --  180 - 0xb4  :  255 - 0xff
    "11111101", --  181 - 0xb5  :  253 - 0xfd
    "11111111", --  182 - 0xb6  :  255 - 0xff
    "11111101", --  183 - 0xb7  :  253 - 0xfd
    "11111111", --  184 - 0xb8  :  255 - 0xff
    "11111101", --  185 - 0xb9  :  253 - 0xfd
    "11111111", --  186 - 0xba  :  255 - 0xff
    "11111101", --  187 - 0xbb  :  253 - 0xfd
    "11111111", --  188 - 0xbc  :  255 - 0xff
    "11111101", --  189 - 0xbd  :  253 - 0xfd
    "11111111", --  190 - 0xbe  :  255 - 0xff
    "11111101", --  191 - 0xbf  :  253 - 0xfd
    "11111111", --  192 - 0xc0  :  255 - 0xff -- line 0x6
    "11111101", --  193 - 0xc1  :  253 - 0xfd
    "11111111", --  194 - 0xc2  :  255 - 0xff
    "11111101", --  195 - 0xc3  :  253 - 0xfd
    "11111111", --  196 - 0xc4  :  255 - 0xff
    "11111101", --  197 - 0xc5  :  253 - 0xfd
    "11111111", --  198 - 0xc6  :  255 - 0xff
    "11111101", --  199 - 0xc7  :  253 - 0xfd
    "11111111", --  200 - 0xc8  :  255 - 0xff
    "11111101", --  201 - 0xc9  :  253 - 0xfd
    "11111111", --  202 - 0xca  :  255 - 0xff
    "11111101", --  203 - 0xcb  :  253 - 0xfd
    "11111111", --  204 - 0xcc  :  255 - 0xff
    "11111101", --  205 - 0xcd  :  253 - 0xfd
    "11111111", --  206 - 0xce  :  255 - 0xff
    "11111101", --  207 - 0xcf  :  253 - 0xfd
    "11111111", --  208 - 0xd0  :  255 - 0xff
    "11111101", --  209 - 0xd1  :  253 - 0xfd
    "11111111", --  210 - 0xd2  :  255 - 0xff
    "11111101", --  211 - 0xd3  :  253 - 0xfd
    "11111111", --  212 - 0xd4  :  255 - 0xff
    "11111101", --  213 - 0xd5  :  253 - 0xfd
    "11111111", --  214 - 0xd6  :  255 - 0xff
    "11111101", --  215 - 0xd7  :  253 - 0xfd
    "11111111", --  216 - 0xd8  :  255 - 0xff
    "11111101", --  217 - 0xd9  :  253 - 0xfd
    "11111111", --  218 - 0xda  :  255 - 0xff
    "11111101", --  219 - 0xdb  :  253 - 0xfd
    "11111111", --  220 - 0xdc  :  255 - 0xff
    "11111101", --  221 - 0xdd  :  253 - 0xfd
    "11111111", --  222 - 0xde  :  255 - 0xff
    "11111101", --  223 - 0xdf  :  253 - 0xfd
    "11111111", --  224 - 0xe0  :  255 - 0xff -- line 0x7
    "11111111", --  225 - 0xe1  :  255 - 0xff
    "11111111", --  226 - 0xe2  :  255 - 0xff
    "11111111", --  227 - 0xe3  :  255 - 0xff
    "11111111", --  228 - 0xe4  :  255 - 0xff
    "11111111", --  229 - 0xe5  :  255 - 0xff
    "11111111", --  230 - 0xe6  :  255 - 0xff
    "11111111", --  231 - 0xe7  :  255 - 0xff
    "11111111", --  232 - 0xe8  :  255 - 0xff
    "11111111", --  233 - 0xe9  :  255 - 0xff
    "11111111", --  234 - 0xea  :  255 - 0xff
    "11111111", --  235 - 0xeb  :  255 - 0xff
    "11111111", --  236 - 0xec  :  255 - 0xff
    "11111111", --  237 - 0xed  :  255 - 0xff
    "11111111", --  238 - 0xee  :  255 - 0xff
    "11111111", --  239 - 0xef  :  255 - 0xff
    "11111111", --  240 - 0xf0  :  255 - 0xff
    "11111111", --  241 - 0xf1  :  255 - 0xff
    "11111111", --  242 - 0xf2  :  255 - 0xff
    "11111111", --  243 - 0xf3  :  255 - 0xff
    "11111111", --  244 - 0xf4  :  255 - 0xff
    "11111111", --  245 - 0xf5  :  255 - 0xff
    "11111111", --  246 - 0xf6  :  255 - 0xff
    "11111111", --  247 - 0xf7  :  255 - 0xff
    "11111111", --  248 - 0xf8  :  255 - 0xff
    "11111111", --  249 - 0xf9  :  255 - 0xff
    "11111111", --  250 - 0xfa  :  255 - 0xff
    "11111111", --  251 - 0xfb  :  255 - 0xff
    "11111111", --  252 - 0xfc  :  255 - 0xff
    "11111111", --  253 - 0xfd  :  255 - 0xff
    "11111111", --  254 - 0xfe  :  255 - 0xff
    "11111111", --  255 - 0xff  :  255 - 0xff
    "11101011", --  256 - 0x100  :  235 - 0xeb -- line 0x8
    "11101011", --  257 - 0x101  :  235 - 0xeb
    "11101011", --  258 - 0x102  :  235 - 0xeb
    "11101011", --  259 - 0x103  :  235 - 0xeb
    "11101011", --  260 - 0x104  :  235 - 0xeb
    "11101011", --  261 - 0x105  :  235 - 0xeb
    "11101011", --  262 - 0x106  :  235 - 0xeb
    "11101011", --  263 - 0x107  :  235 - 0xeb
    "11101011", --  264 - 0x108  :  235 - 0xeb
    "11101011", --  265 - 0x109  :  235 - 0xeb
    "11101011", --  266 - 0x10a  :  235 - 0xeb
    "11101011", --  267 - 0x10b  :  235 - 0xeb
    "11101011", --  268 - 0x10c  :  235 - 0xeb
    "11101011", --  269 - 0x10d  :  235 - 0xeb
    "11101011", --  270 - 0x10e  :  235 - 0xeb
    "11101011", --  271 - 0x10f  :  235 - 0xeb
    "11101011", --  272 - 0x110  :  235 - 0xeb
    "11101011", --  273 - 0x111  :  235 - 0xeb
    "11101011", --  274 - 0x112  :  235 - 0xeb
    "11101011", --  275 - 0x113  :  235 - 0xeb
    "11101011", --  276 - 0x114  :  235 - 0xeb
    "11101011", --  277 - 0x115  :  235 - 0xeb
    "11101011", --  278 - 0x116  :  235 - 0xeb
    "11101011", --  279 - 0x117  :  235 - 0xeb
    "11101011", --  280 - 0x118  :  235 - 0xeb
    "11101011", --  281 - 0x119  :  235 - 0xeb
    "11101011", --  282 - 0x11a  :  235 - 0xeb
    "11101011", --  283 - 0x11b  :  235 - 0xeb
    "11101011", --  284 - 0x11c  :  235 - 0xeb
    "11101011", --  285 - 0x11d  :  235 - 0xeb
    "11101011", --  286 - 0x11e  :  235 - 0xeb
    "11101011", --  287 - 0x11f  :  235 - 0xeb
    "11111010", --  288 - 0x120  :  250 - 0xfa -- line 0x9
    "11111010", --  289 - 0x121  :  250 - 0xfa
    "11101001", --  290 - 0x122  :  233 - 0xe9
    "11111010", --  291 - 0x123  :  250 - 0xfa
    "11111010", --  292 - 0x124  :  250 - 0xfa
    "11111010", --  293 - 0x125  :  250 - 0xfa
    "11111010", --  294 - 0x126  :  250 - 0xfa
    "11111010", --  295 - 0x127  :  250 - 0xfa
    "11111010", --  296 - 0x128  :  250 - 0xfa
    "11111010", --  297 - 0x129  :  250 - 0xfa
    "11111010", --  298 - 0x12a  :  250 - 0xfa
    "11111010", --  299 - 0x12b  :  250 - 0xfa
    "11111010", --  300 - 0x12c  :  250 - 0xfa
    "11111010", --  301 - 0x12d  :  250 - 0xfa
    "11111010", --  302 - 0x12e  :  250 - 0xfa
    "11111010", --  303 - 0x12f  :  250 - 0xfa
    "11111010", --  304 - 0x130  :  250 - 0xfa
    "11111010", --  305 - 0x131  :  250 - 0xfa
    "11111010", --  306 - 0x132  :  250 - 0xfa
    "11111010", --  307 - 0x133  :  250 - 0xfa
    "11111010", --  308 - 0x134  :  250 - 0xfa
    "11111010", --  309 - 0x135  :  250 - 0xfa
    "11111010", --  310 - 0x136  :  250 - 0xfa
    "11101010", --  311 - 0x137  :  234 - 0xea
    "11111010", --  312 - 0x138  :  250 - 0xfa
    "11111010", --  313 - 0x139  :  250 - 0xfa
    "11111010", --  314 - 0x13a  :  250 - 0xfa
    "11111010", --  315 - 0x13b  :  250 - 0xfa
    "11111010", --  316 - 0x13c  :  250 - 0xfa
    "11111010", --  317 - 0x13d  :  250 - 0xfa
    "11111010", --  318 - 0x13e  :  250 - 0xfa
    "11111010", --  319 - 0x13f  :  250 - 0xfa
    "11111010", --  320 - 0x140  :  250 - 0xfa -- line 0xa
    "11111010", --  321 - 0x141  :  250 - 0xfa
    "11111010", --  322 - 0x142  :  250 - 0xfa
    "11111010", --  323 - 0x143  :  250 - 0xfa
    "11111010", --  324 - 0x144  :  250 - 0xfa
    "11111010", --  325 - 0x145  :  250 - 0xfa
    "11111010", --  326 - 0x146  :  250 - 0xfa
    "11111010", --  327 - 0x147  :  250 - 0xfa
    "11111010", --  328 - 0x148  :  250 - 0xfa
    "11111010", --  329 - 0x149  :  250 - 0xfa
    "11111010", --  330 - 0x14a  :  250 - 0xfa
    "11111010", --  331 - 0x14b  :  250 - 0xfa
    "11111010", --  332 - 0x14c  :  250 - 0xfa
    "11111010", --  333 - 0x14d  :  250 - 0xfa
    "11111010", --  334 - 0x14e  :  250 - 0xfa
    "11111010", --  335 - 0x14f  :  250 - 0xfa
    "11111010", --  336 - 0x150  :  250 - 0xfa
    "11111010", --  337 - 0x151  :  250 - 0xfa
    "11111010", --  338 - 0x152  :  250 - 0xfa
    "11111010", --  339 - 0x153  :  250 - 0xfa
    "11111010", --  340 - 0x154  :  250 - 0xfa
    "11111010", --  341 - 0x155  :  250 - 0xfa
    "11111010", --  342 - 0x156  :  250 - 0xfa
    "11111010", --  343 - 0x157  :  250 - 0xfa
    "11111010", --  344 - 0x158  :  250 - 0xfa
    "11111010", --  345 - 0x159  :  250 - 0xfa
    "11111010", --  346 - 0x15a  :  250 - 0xfa
    "11111010", --  347 - 0x15b  :  250 - 0xfa
    "11111010", --  348 - 0x15c  :  250 - 0xfa
    "11101010", --  349 - 0x15d  :  234 - 0xea
    "11111010", --  350 - 0x15e  :  250 - 0xfa
    "11111010", --  351 - 0x15f  :  250 - 0xfa
    "11111010", --  352 - 0x160  :  250 - 0xfa -- line 0xb
    "11111010", --  353 - 0x161  :  250 - 0xfa
    "11111010", --  354 - 0x162  :  250 - 0xfa
    "11111010", --  355 - 0x163  :  250 - 0xfa
    "11111010", --  356 - 0x164  :  250 - 0xfa
    "11111010", --  357 - 0x165  :  250 - 0xfa
    "11111010", --  358 - 0x166  :  250 - 0xfa
    "11111010", --  359 - 0x167  :  250 - 0xfa
    "11111010", --  360 - 0x168  :  250 - 0xfa
    "11111010", --  361 - 0x169  :  250 - 0xfa
    "11111010", --  362 - 0x16a  :  250 - 0xfa
    "11111010", --  363 - 0x16b  :  250 - 0xfa
    "11111010", --  364 - 0x16c  :  250 - 0xfa
    "11111010", --  365 - 0x16d  :  250 - 0xfa
    "11111010", --  366 - 0x16e  :  250 - 0xfa
    "11111010", --  367 - 0x16f  :  250 - 0xfa
    "11111010", --  368 - 0x170  :  250 - 0xfa
    "11111010", --  369 - 0x171  :  250 - 0xfa
    "11111010", --  370 - 0x172  :  250 - 0xfa
    "11111010", --  371 - 0x173  :  250 - 0xfa
    "11111010", --  372 - 0x174  :  250 - 0xfa
    "11111010", --  373 - 0x175  :  250 - 0xfa
    "11111010", --  374 - 0x176  :  250 - 0xfa
    "11111010", --  375 - 0x177  :  250 - 0xfa
    "11111010", --  376 - 0x178  :  250 - 0xfa
    "11111010", --  377 - 0x179  :  250 - 0xfa
    "11111010", --  378 - 0x17a  :  250 - 0xfa
    "11111010", --  379 - 0x17b  :  250 - 0xfa
    "11111010", --  380 - 0x17c  :  250 - 0xfa
    "11111010", --  381 - 0x17d  :  250 - 0xfa
    "11111010", --  382 - 0x17e  :  250 - 0xfa
    "11111010", --  383 - 0x17f  :  250 - 0xfa
    "11111010", --  384 - 0x180  :  250 - 0xfa -- line 0xc
    "11111010", --  385 - 0x181  :  250 - 0xfa
    "11111010", --  386 - 0x182  :  250 - 0xfa
    "11111010", --  387 - 0x183  :  250 - 0xfa
    "11111010", --  388 - 0x184  :  250 - 0xfa
    "11111010", --  389 - 0x185  :  250 - 0xfa
    "11111010", --  390 - 0x186  :  250 - 0xfa
    "11111010", --  391 - 0x187  :  250 - 0xfa
    "11111010", --  392 - 0x188  :  250 - 0xfa
    "11111010", --  393 - 0x189  :  250 - 0xfa
    "11111010", --  394 - 0x18a  :  250 - 0xfa
    "11111010", --  395 - 0x18b  :  250 - 0xfa
    "11111010", --  396 - 0x18c  :  250 - 0xfa
    "11111010", --  397 - 0x18d  :  250 - 0xfa
    "11111010", --  398 - 0x18e  :  250 - 0xfa
    "11111010", --  399 - 0x18f  :  250 - 0xfa
    "11111010", --  400 - 0x190  :  250 - 0xfa
    "11101001", --  401 - 0x191  :  233 - 0xe9
    "11111001", --  402 - 0x192  :  249 - 0xf9
    "11111010", --  403 - 0x193  :  250 - 0xfa
    "11111010", --  404 - 0x194  :  250 - 0xfa
    "11111010", --  405 - 0x195  :  250 - 0xfa
    "11111010", --  406 - 0x196  :  250 - 0xfa
    "11111010", --  407 - 0x197  :  250 - 0xfa
    "11111010", --  408 - 0x198  :  250 - 0xfa
    "11111010", --  409 - 0x199  :  250 - 0xfa
    "11111010", --  410 - 0x19a  :  250 - 0xfa
    "11111010", --  411 - 0x19b  :  250 - 0xfa
    "11111010", --  412 - 0x19c  :  250 - 0xfa
    "11111010", --  413 - 0x19d  :  250 - 0xfa
    "11111010", --  414 - 0x19e  :  250 - 0xfa
    "11111010", --  415 - 0x19f  :  250 - 0xfa
    "11111010", --  416 - 0x1a0  :  250 - 0xfa -- line 0xd
    "11111010", --  417 - 0x1a1  :  250 - 0xfa
    "11111010", --  418 - 0x1a2  :  250 - 0xfa
    "11111010", --  419 - 0x1a3  :  250 - 0xfa
    "11101010", --  420 - 0x1a4  :  234 - 0xea
    "11111010", --  421 - 0x1a5  :  250 - 0xfa
    "11111010", --  422 - 0x1a6  :  250 - 0xfa
    "11111010", --  423 - 0x1a7  :  250 - 0xfa
    "11111001", --  424 - 0x1a8  :  249 - 0xf9
    "11111010", --  425 - 0x1a9  :  250 - 0xfa
    "11111010", --  426 - 0x1aa  :  250 - 0xfa
    "11111010", --  427 - 0x1ab  :  250 - 0xfa
    "11111010", --  428 - 0x1ac  :  250 - 0xfa
    "11111010", --  429 - 0x1ad  :  250 - 0xfa
    "00011101", --  430 - 0x1ae  :   29 - 0x1d
    "00010001", --  431 - 0x1af  :   17 - 0x11
    "00010100", --  432 - 0x1b0  :   20 - 0x14
    "00010101", --  433 - 0x1b1  :   21 - 0x15
    "11111010", --  434 - 0x1b2  :  250 - 0xfa
    "11111010", --  435 - 0x1b3  :  250 - 0xfa
    "11111010", --  436 - 0x1b4  :  250 - 0xfa
    "11111010", --  437 - 0x1b5  :  250 - 0xfa
    "11111010", --  438 - 0x1b6  :  250 - 0xfa
    "11111010", --  439 - 0x1b7  :  250 - 0xfa
    "11111010", --  440 - 0x1b8  :  250 - 0xfa
    "11111010", --  441 - 0x1b9  :  250 - 0xfa
    "11111010", --  442 - 0x1ba  :  250 - 0xfa
    "11111010", --  443 - 0x1bb  :  250 - 0xfa
    "11111010", --  444 - 0x1bc  :  250 - 0xfa
    "11111010", --  445 - 0x1bd  :  250 - 0xfa
    "11111010", --  446 - 0x1be  :  250 - 0xfa
    "11111010", --  447 - 0x1bf  :  250 - 0xfa
    "11111010", --  448 - 0x1c0  :  250 - 0xfa -- line 0xe
    "11111010", --  449 - 0x1c1  :  250 - 0xfa
    "11111010", --  450 - 0x1c2  :  250 - 0xfa
    "11111010", --  451 - 0x1c3  :  250 - 0xfa
    "11111010", --  452 - 0x1c4  :  250 - 0xfa
    "11111010", --  453 - 0x1c5  :  250 - 0xfa
    "11111010", --  454 - 0x1c6  :  250 - 0xfa
    "11111010", --  455 - 0x1c7  :  250 - 0xfa
    "11111010", --  456 - 0x1c8  :  250 - 0xfa
    "11111010", --  457 - 0x1c9  :  250 - 0xfa
    "11111010", --  458 - 0x1ca  :  250 - 0xfa
    "11111010", --  459 - 0x1cb  :  250 - 0xfa
    "11111010", --  460 - 0x1cc  :  250 - 0xfa
    "11111010", --  461 - 0x1cd  :  250 - 0xfa
    "11111010", --  462 - 0x1ce  :  250 - 0xfa
    "11111010", --  463 - 0x1cf  :  250 - 0xfa
    "11111010", --  464 - 0x1d0  :  250 - 0xfa
    "11111010", --  465 - 0x1d1  :  250 - 0xfa
    "11111010", --  466 - 0x1d2  :  250 - 0xfa
    "11111010", --  467 - 0x1d3  :  250 - 0xfa
    "11111010", --  468 - 0x1d4  :  250 - 0xfa
    "11111010", --  469 - 0x1d5  :  250 - 0xfa
    "11111010", --  470 - 0x1d6  :  250 - 0xfa
    "11111010", --  471 - 0x1d7  :  250 - 0xfa
    "11111010", --  472 - 0x1d8  :  250 - 0xfa
    "11111010", --  473 - 0x1d9  :  250 - 0xfa
    "11111010", --  474 - 0x1da  :  250 - 0xfa
    "11111010", --  475 - 0x1db  :  250 - 0xfa
    "11111010", --  476 - 0x1dc  :  250 - 0xfa
    "11111010", --  477 - 0x1dd  :  250 - 0xfa
    "11111010", --  478 - 0x1de  :  250 - 0xfa
    "11111010", --  479 - 0x1df  :  250 - 0xfa
    "11111010", --  480 - 0x1e0  :  250 - 0xfa -- line 0xf
    "11111001", --  481 - 0x1e1  :  249 - 0xf9
    "11111010", --  482 - 0x1e2  :  250 - 0xfa
    "11111010", --  483 - 0x1e3  :  250 - 0xfa
    "11111010", --  484 - 0x1e4  :  250 - 0xfa
    "11111010", --  485 - 0x1e5  :  250 - 0xfa
    "11111010", --  486 - 0x1e6  :  250 - 0xfa
    "11111010", --  487 - 0x1e7  :  250 - 0xfa
    "11111010", --  488 - 0x1e8  :  250 - 0xfa
    "11111010", --  489 - 0x1e9  :  250 - 0xfa
    "11111010", --  490 - 0x1ea  :  250 - 0xfa
    "11111010", --  491 - 0x1eb  :  250 - 0xfa
    "00010110", --  492 - 0x1ec  :   22 - 0x16
    "00011111", --  493 - 0x1ed  :   31 - 0x1f
    "00100010", --  494 - 0x1ee  :   34 - 0x22
    "11111010", --  495 - 0x1ef  :  250 - 0xfa
    "11111010", --  496 - 0x1f0  :  250 - 0xfa
    "00100100", --  497 - 0x1f1  :   36 - 0x24
    "00011000", --  498 - 0x1f2  :   24 - 0x18
    "00010101", --  499 - 0x1f3  :   21 - 0x15
    "11111010", --  500 - 0x1f4  :  250 - 0xfa
    "11111010", --  501 - 0x1f5  :  250 - 0xfa
    "11111010", --  502 - 0x1f6  :  250 - 0xfa
    "11101001", --  503 - 0x1f7  :  233 - 0xe9
    "11111010", --  504 - 0x1f8  :  250 - 0xfa
    "11111010", --  505 - 0x1f9  :  250 - 0xfa
    "11111010", --  506 - 0x1fa  :  250 - 0xfa
    "11111010", --  507 - 0x1fb  :  250 - 0xfa
    "11111010", --  508 - 0x1fc  :  250 - 0xfa
    "11111010", --  509 - 0x1fd  :  250 - 0xfa
    "11111010", --  510 - 0x1fe  :  250 - 0xfa
    "11111010", --  511 - 0x1ff  :  250 - 0xfa
    "11111010", --  512 - 0x200  :  250 - 0xfa -- line 0x10
    "11111010", --  513 - 0x201  :  250 - 0xfa
    "11111010", --  514 - 0x202  :  250 - 0xfa
    "11111010", --  515 - 0x203  :  250 - 0xfa
    "11111010", --  516 - 0x204  :  250 - 0xfa
    "11111010", --  517 - 0x205  :  250 - 0xfa
    "11111010", --  518 - 0x206  :  250 - 0xfa
    "11111010", --  519 - 0x207  :  250 - 0xfa
    "11111010", --  520 - 0x208  :  250 - 0xfa
    "11101010", --  521 - 0x209  :  234 - 0xea
    "11111010", --  522 - 0x20a  :  250 - 0xfa
    "11111010", --  523 - 0x20b  :  250 - 0xfa
    "11111010", --  524 - 0x20c  :  250 - 0xfa
    "11111010", --  525 - 0x20d  :  250 - 0xfa
    "11111010", --  526 - 0x20e  :  250 - 0xfa
    "11111010", --  527 - 0x20f  :  250 - 0xfa
    "11111010", --  528 - 0x210  :  250 - 0xfa
    "11111010", --  529 - 0x211  :  250 - 0xfa
    "11111010", --  530 - 0x212  :  250 - 0xfa
    "11111010", --  531 - 0x213  :  250 - 0xfa
    "11111010", --  532 - 0x214  :  250 - 0xfa
    "11111010", --  533 - 0x215  :  250 - 0xfa
    "11111010", --  534 - 0x216  :  250 - 0xfa
    "11111010", --  535 - 0x217  :  250 - 0xfa
    "11111010", --  536 - 0x218  :  250 - 0xfa
    "11111010", --  537 - 0x219  :  250 - 0xfa
    "11111010", --  538 - 0x21a  :  250 - 0xfa
    "11111010", --  539 - 0x21b  :  250 - 0xfa
    "11111010", --  540 - 0x21c  :  250 - 0xfa
    "11101010", --  541 - 0x21d  :  234 - 0xea
    "11111010", --  542 - 0x21e  :  250 - 0xfa
    "11111010", --  543 - 0x21f  :  250 - 0xfa
    "11111010", --  544 - 0x220  :  250 - 0xfa -- line 0x11
    "11111010", --  545 - 0x221  :  250 - 0xfa
    "11111010", --  546 - 0x222  :  250 - 0xfa
    "11111010", --  547 - 0x223  :  250 - 0xfa
    "11111010", --  548 - 0x224  :  250 - 0xfa
    "11111010", --  549 - 0x225  :  250 - 0xfa
    "11111010", --  550 - 0x226  :  250 - 0xfa
    "11111010", --  551 - 0x227  :  250 - 0xfa
    "11111010", --  552 - 0x228  :  250 - 0xfa
    "11111010", --  553 - 0x229  :  250 - 0xfa
    "11111010", --  554 - 0x22a  :  250 - 0xfa
    "11111010", --  555 - 0x22b  :  250 - 0xfa
    "11111010", --  556 - 0x22c  :  250 - 0xfa
    "11111010", --  557 - 0x22d  :  250 - 0xfa
    "00000010", --  558 - 0x22e  :    2 - 0x2
    "00000000", --  559 - 0x22f  :    0 - 0x0
    "00000001", --  560 - 0x230  :    1 - 0x1
    "00000111", --  561 - 0x231  :    7 - 0x7
    "11111010", --  562 - 0x232  :  250 - 0xfa
    "11111010", --  563 - 0x233  :  250 - 0xfa
    "11111010", --  564 - 0x234  :  250 - 0xfa
    "11111010", --  565 - 0x235  :  250 - 0xfa
    "11111010", --  566 - 0x236  :  250 - 0xfa
    "11111010", --  567 - 0x237  :  250 - 0xfa
    "11111010", --  568 - 0x238  :  250 - 0xfa
    "11111010", --  569 - 0x239  :  250 - 0xfa
    "11111010", --  570 - 0x23a  :  250 - 0xfa
    "11111010", --  571 - 0x23b  :  250 - 0xfa
    "11111010", --  572 - 0x23c  :  250 - 0xfa
    "11111010", --  573 - 0x23d  :  250 - 0xfa
    "11111010", --  574 - 0x23e  :  250 - 0xfa
    "11111010", --  575 - 0x23f  :  250 - 0xfa
    "11111010", --  576 - 0x240  :  250 - 0xfa -- line 0x12
    "11111010", --  577 - 0x241  :  250 - 0xfa
    "11111010", --  578 - 0x242  :  250 - 0xfa
    "11111010", --  579 - 0x243  :  250 - 0xfa
    "11111001", --  580 - 0x244  :  249 - 0xf9
    "11111010", --  581 - 0x245  :  250 - 0xfa
    "11111010", --  582 - 0x246  :  250 - 0xfa
    "11111010", --  583 - 0x247  :  250 - 0xfa
    "11111010", --  584 - 0x248  :  250 - 0xfa
    "11111010", --  585 - 0x249  :  250 - 0xfa
    "11111010", --  586 - 0x24a  :  250 - 0xfa
    "11111010", --  587 - 0x24b  :  250 - 0xfa
    "11111010", --  588 - 0x24c  :  250 - 0xfa
    "11111010", --  589 - 0x24d  :  250 - 0xfa
    "11111010", --  590 - 0x24e  :  250 - 0xfa
    "11111010", --  591 - 0x24f  :  250 - 0xfa
    "11111010", --  592 - 0x250  :  250 - 0xfa
    "11111010", --  593 - 0x251  :  250 - 0xfa
    "11111010", --  594 - 0x252  :  250 - 0xfa
    "11111010", --  595 - 0x253  :  250 - 0xfa
    "11111010", --  596 - 0x254  :  250 - 0xfa
    "11111010", --  597 - 0x255  :  250 - 0xfa
    "11111010", --  598 - 0x256  :  250 - 0xfa
    "11111010", --  599 - 0x257  :  250 - 0xfa
    "11111010", --  600 - 0x258  :  250 - 0xfa
    "11111010", --  601 - 0x259  :  250 - 0xfa
    "11111010", --  602 - 0x25a  :  250 - 0xfa
    "11111010", --  603 - 0x25b  :  250 - 0xfa
    "11111010", --  604 - 0x25c  :  250 - 0xfa
    "11111010", --  605 - 0x25d  :  250 - 0xfa
    "11111010", --  606 - 0x25e  :  250 - 0xfa
    "11111010", --  607 - 0x25f  :  250 - 0xfa
    "11111010", --  608 - 0x260  :  250 - 0xfa -- line 0x13
    "11111010", --  609 - 0x261  :  250 - 0xfa
    "11111010", --  610 - 0x262  :  250 - 0xfa
    "11111010", --  611 - 0x263  :  250 - 0xfa
    "11111010", --  612 - 0x264  :  250 - 0xfa
    "11111010", --  613 - 0x265  :  250 - 0xfa
    "11111010", --  614 - 0x266  :  250 - 0xfa
    "11111010", --  615 - 0x267  :  250 - 0xfa
    "11111010", --  616 - 0x268  :  250 - 0xfa
    "11111010", --  617 - 0x269  :  250 - 0xfa
    "11111010", --  618 - 0x26a  :  250 - 0xfa
    "11111010", --  619 - 0x26b  :  250 - 0xfa
    "11111010", --  620 - 0x26c  :  250 - 0xfa
    "00010111", --  621 - 0x26d  :   23 - 0x17
    "00011001", --  622 - 0x26e  :   25 - 0x19
    "00100100", --  623 - 0x26f  :   36 - 0x24
    "00011000", --  624 - 0x270  :   24 - 0x18
    "00100101", --  625 - 0x271  :   37 - 0x25
    "00010010", --  626 - 0x272  :   18 - 0x12
    "11111010", --  627 - 0x273  :  250 - 0xfa
    "11111010", --  628 - 0x274  :  250 - 0xfa
    "11111010", --  629 - 0x275  :  250 - 0xfa
    "11111010", --  630 - 0x276  :  250 - 0xfa
    "11101010", --  631 - 0x277  :  234 - 0xea
    "11101001", --  632 - 0x278  :  233 - 0xe9
    "11111010", --  633 - 0x279  :  250 - 0xfa
    "11111010", --  634 - 0x27a  :  250 - 0xfa
    "11111010", --  635 - 0x27b  :  250 - 0xfa
    "11111001", --  636 - 0x27c  :  249 - 0xf9
    "11111010", --  637 - 0x27d  :  250 - 0xfa
    "11111010", --  638 - 0x27e  :  250 - 0xfa
    "11111010", --  639 - 0x27f  :  250 - 0xfa
    "11111010", --  640 - 0x280  :  250 - 0xfa -- line 0x14
    "11111010", --  641 - 0x281  :  250 - 0xfa
    "11111010", --  642 - 0x282  :  250 - 0xfa
    "11111010", --  643 - 0x283  :  250 - 0xfa
    "11111010", --  644 - 0x284  :  250 - 0xfa
    "11111010", --  645 - 0x285  :  250 - 0xfa
    "11111010", --  646 - 0x286  :  250 - 0xfa
    "11111010", --  647 - 0x287  :  250 - 0xfa
    "11111010", --  648 - 0x288  :  250 - 0xfa
    "11111010", --  649 - 0x289  :  250 - 0xfa
    "11111010", --  650 - 0x28a  :  250 - 0xfa
    "11111010", --  651 - 0x28b  :  250 - 0xfa
    "11111010", --  652 - 0x28c  :  250 - 0xfa
    "11111010", --  653 - 0x28d  :  250 - 0xfa
    "11111010", --  654 - 0x28e  :  250 - 0xfa
    "11111010", --  655 - 0x28f  :  250 - 0xfa
    "11111010", --  656 - 0x290  :  250 - 0xfa
    "11111010", --  657 - 0x291  :  250 - 0xfa
    "11111010", --  658 - 0x292  :  250 - 0xfa
    "11111010", --  659 - 0x293  :  250 - 0xfa
    "11111010", --  660 - 0x294  :  250 - 0xfa
    "11111010", --  661 - 0x295  :  250 - 0xfa
    "11111010", --  662 - 0x296  :  250 - 0xfa
    "11111010", --  663 - 0x297  :  250 - 0xfa
    "11111010", --  664 - 0x298  :  250 - 0xfa
    "11111010", --  665 - 0x299  :  250 - 0xfa
    "11111010", --  666 - 0x29a  :  250 - 0xfa
    "11111010", --  667 - 0x29b  :  250 - 0xfa
    "11111010", --  668 - 0x29c  :  250 - 0xfa
    "11111010", --  669 - 0x29d  :  250 - 0xfa
    "11111010", --  670 - 0x29e  :  250 - 0xfa
    "11111010", --  671 - 0x29f  :  250 - 0xfa
    "11111010", --  672 - 0x2a0  :  250 - 0xfa -- line 0x15
    "11111010", --  673 - 0x2a1  :  250 - 0xfa
    "11101010", --  674 - 0x2a2  :  234 - 0xea
    "11111010", --  675 - 0x2a3  :  250 - 0xfa
    "11111010", --  676 - 0x2a4  :  250 - 0xfa
    "11111010", --  677 - 0x2a5  :  250 - 0xfa
    "11111010", --  678 - 0x2a6  :  250 - 0xfa
    "11111010", --  679 - 0x2a7  :  250 - 0xfa
    "11111010", --  680 - 0x2a8  :  250 - 0xfa
    "11111010", --  681 - 0x2a9  :  250 - 0xfa
    "11111010", --  682 - 0x2aa  :  250 - 0xfa
    "11111010", --  683 - 0x2ab  :  250 - 0xfa
    "00010111", --  684 - 0x2ac  :   23 - 0x17
    "00010001", --  685 - 0x2ad  :   17 - 0x11
    "00011101", --  686 - 0x2ae  :   29 - 0x1d
    "00010101", --  687 - 0x2af  :   21 - 0x15
    "11101010", --  688 - 0x2b0  :  234 - 0xea
    "00011111", --  689 - 0x2b1  :   31 - 0x1f
    "00010110", --  690 - 0x2b2  :   22 - 0x16
    "00010110", --  691 - 0x2b3  :   22 - 0x16
    "11111010", --  692 - 0x2b4  :  250 - 0xfa
    "11111010", --  693 - 0x2b5  :  250 - 0xfa
    "11111010", --  694 - 0x2b6  :  250 - 0xfa
    "11111010", --  695 - 0x2b7  :  250 - 0xfa
    "11111010", --  696 - 0x2b8  :  250 - 0xfa
    "11111010", --  697 - 0x2b9  :  250 - 0xfa
    "11111010", --  698 - 0x2ba  :  250 - 0xfa
    "11111010", --  699 - 0x2bb  :  250 - 0xfa
    "11111010", --  700 - 0x2bc  :  250 - 0xfa
    "11111010", --  701 - 0x2bd  :  250 - 0xfa
    "11111010", --  702 - 0x2be  :  250 - 0xfa
    "11111010", --  703 - 0x2bf  :  250 - 0xfa
    "11111010", --  704 - 0x2c0  :  250 - 0xfa -- line 0x16
    "11111010", --  705 - 0x2c1  :  250 - 0xfa
    "11111010", --  706 - 0x2c2  :  250 - 0xfa
    "11111010", --  707 - 0x2c3  :  250 - 0xfa
    "11111010", --  708 - 0x2c4  :  250 - 0xfa
    "11111010", --  709 - 0x2c5  :  250 - 0xfa
    "11111010", --  710 - 0x2c6  :  250 - 0xfa
    "11111010", --  711 - 0x2c7  :  250 - 0xfa
    "11111010", --  712 - 0x2c8  :  250 - 0xfa
    "11111010", --  713 - 0x2c9  :  250 - 0xfa
    "11111010", --  714 - 0x2ca  :  250 - 0xfa
    "11111010", --  715 - 0x2cb  :  250 - 0xfa
    "11111010", --  716 - 0x2cc  :  250 - 0xfa
    "11111010", --  717 - 0x2cd  :  250 - 0xfa
    "11111010", --  718 - 0x2ce  :  250 - 0xfa
    "11111010", --  719 - 0x2cf  :  250 - 0xfa
    "11111010", --  720 - 0x2d0  :  250 - 0xfa
    "11111010", --  721 - 0x2d1  :  250 - 0xfa
    "11111010", --  722 - 0x2d2  :  250 - 0xfa
    "11111010", --  723 - 0x2d3  :  250 - 0xfa
    "11111010", --  724 - 0x2d4  :  250 - 0xfa
    "11111010", --  725 - 0x2d5  :  250 - 0xfa
    "11111010", --  726 - 0x2d6  :  250 - 0xfa
    "11111010", --  727 - 0x2d7  :  250 - 0xfa
    "11111010", --  728 - 0x2d8  :  250 - 0xfa
    "11111010", --  729 - 0x2d9  :  250 - 0xfa
    "11111010", --  730 - 0x2da  :  250 - 0xfa
    "11111010", --  731 - 0x2db  :  250 - 0xfa
    "11111010", --  732 - 0x2dc  :  250 - 0xfa
    "11111010", --  733 - 0x2dd  :  250 - 0xfa
    "11111010", --  734 - 0x2de  :  250 - 0xfa
    "11111010", --  735 - 0x2df  :  250 - 0xfa
    "11111010", --  736 - 0x2e0  :  250 - 0xfa -- line 0x17
    "11111010", --  737 - 0x2e1  :  250 - 0xfa
    "11111010", --  738 - 0x2e2  :  250 - 0xfa
    "11111010", --  739 - 0x2e3  :  250 - 0xfa
    "11111010", --  740 - 0x2e4  :  250 - 0xfa
    "11111010", --  741 - 0x2e5  :  250 - 0xfa
    "11111010", --  742 - 0x2e6  :  250 - 0xfa
    "11111001", --  743 - 0x2e7  :  249 - 0xf9
    "11111010", --  744 - 0x2e8  :  250 - 0xfa
    "11111010", --  745 - 0x2e9  :  250 - 0xfa
    "11111010", --  746 - 0x2ea  :  250 - 0xfa
    "11111010", --  747 - 0x2eb  :  250 - 0xfa
    "11111010", --  748 - 0x2ec  :  250 - 0xfa
    "11111010", --  749 - 0x2ed  :  250 - 0xfa
    "11111010", --  750 - 0x2ee  :  250 - 0xfa
    "00010010", --  751 - 0x2ef  :   18 - 0x12
    "00101001", --  752 - 0x2f0  :   41 - 0x29
    "11111010", --  753 - 0x2f1  :  250 - 0xfa
    "11111010", --  754 - 0x2f2  :  250 - 0xfa
    "11111010", --  755 - 0x2f3  :  250 - 0xfa
    "11111010", --  756 - 0x2f4  :  250 - 0xfa
    "11111010", --  757 - 0x2f5  :  250 - 0xfa
    "11111010", --  758 - 0x2f6  :  250 - 0xfa
    "11111010", --  759 - 0x2f7  :  250 - 0xfa
    "11111010", --  760 - 0x2f8  :  250 - 0xfa
    "11111010", --  761 - 0x2f9  :  250 - 0xfa
    "11111010", --  762 - 0x2fa  :  250 - 0xfa
    "11111010", --  763 - 0x2fb  :  250 - 0xfa
    "11111010", --  764 - 0x2fc  :  250 - 0xfa
    "11111010", --  765 - 0x2fd  :  250 - 0xfa
    "11101010", --  766 - 0x2fe  :  234 - 0xea
    "11111010", --  767 - 0x2ff  :  250 - 0xfa
    "11111010", --  768 - 0x300  :  250 - 0xfa -- line 0x18
    "11111010", --  769 - 0x301  :  250 - 0xfa
    "11111010", --  770 - 0x302  :  250 - 0xfa
    "11111010", --  771 - 0x303  :  250 - 0xfa
    "11111010", --  772 - 0x304  :  250 - 0xfa
    "11111010", --  773 - 0x305  :  250 - 0xfa
    "11111010", --  774 - 0x306  :  250 - 0xfa
    "11111010", --  775 - 0x307  :  250 - 0xfa
    "11111010", --  776 - 0x308  :  250 - 0xfa
    "11111010", --  777 - 0x309  :  250 - 0xfa
    "11111010", --  778 - 0x30a  :  250 - 0xfa
    "11111010", --  779 - 0x30b  :  250 - 0xfa
    "11111010", --  780 - 0x30c  :  250 - 0xfa
    "11111010", --  781 - 0x30d  :  250 - 0xfa
    "11111010", --  782 - 0x30e  :  250 - 0xfa
    "11111010", --  783 - 0x30f  :  250 - 0xfa
    "11111010", --  784 - 0x310  :  250 - 0xfa
    "11111010", --  785 - 0x311  :  250 - 0xfa
    "11111010", --  786 - 0x312  :  250 - 0xfa
    "11111010", --  787 - 0x313  :  250 - 0xfa
    "11111010", --  788 - 0x314  :  250 - 0xfa
    "11111010", --  789 - 0x315  :  250 - 0xfa
    "11111010", --  790 - 0x316  :  250 - 0xfa
    "11111010", --  791 - 0x317  :  250 - 0xfa
    "11111010", --  792 - 0x318  :  250 - 0xfa
    "11111010", --  793 - 0x319  :  250 - 0xfa
    "11111001", --  794 - 0x31a  :  249 - 0xf9
    "11111010", --  795 - 0x31b  :  250 - 0xfa
    "11111010", --  796 - 0x31c  :  250 - 0xfa
    "11111010", --  797 - 0x31d  :  250 - 0xfa
    "11111010", --  798 - 0x31e  :  250 - 0xfa
    "11111010", --  799 - 0x31f  :  250 - 0xfa
    "11111010", --  800 - 0x320  :  250 - 0xfa -- line 0x19
    "11111010", --  801 - 0x321  :  250 - 0xfa
    "11111010", --  802 - 0x322  :  250 - 0xfa
    "11111010", --  803 - 0x323  :  250 - 0xfa
    "11111010", --  804 - 0x324  :  250 - 0xfa
    "11111010", --  805 - 0x325  :  250 - 0xfa
    "11111010", --  806 - 0x326  :  250 - 0xfa
    "11111010", --  807 - 0x327  :  250 - 0xfa
    "11111010", --  808 - 0x328  :  250 - 0xfa
    "00010011", --  809 - 0x329  :   19 - 0x13
    "00010001", --  810 - 0x32a  :   17 - 0x11
    "00011101", --  811 - 0x32b  :   29 - 0x1d
    "00010101", --  812 - 0x32c  :   21 - 0x15
    "00100010", --  813 - 0x32d  :   34 - 0x22
    "00011111", --  814 - 0x32e  :   31 - 0x1f
    "00011110", --  815 - 0x32f  :   30 - 0x1e
    "11111010", --  816 - 0x330  :  250 - 0xfa
    "11111010", --  817 - 0x331  :  250 - 0xfa
    "00010010", --  818 - 0x332  :   18 - 0x12
    "00100010", --  819 - 0x333  :   34 - 0x22
    "00011111", --  820 - 0x334  :   31 - 0x1f
    "00100111", --  821 - 0x335  :   39 - 0x27
    "00011110", --  822 - 0x336  :   30 - 0x1e
    "11111010", --  823 - 0x337  :  250 - 0xfa
    "11111010", --  824 - 0x338  :  250 - 0xfa
    "11111010", --  825 - 0x339  :  250 - 0xfa
    "11111010", --  826 - 0x33a  :  250 - 0xfa
    "11111010", --  827 - 0x33b  :  250 - 0xfa
    "11111010", --  828 - 0x33c  :  250 - 0xfa
    "11111010", --  829 - 0x33d  :  250 - 0xfa
    "11111010", --  830 - 0x33e  :  250 - 0xfa
    "11111010", --  831 - 0x33f  :  250 - 0xfa
    "11111010", --  832 - 0x340  :  250 - 0xfa -- line 0x1a
    "11111010", --  833 - 0x341  :  250 - 0xfa
    "11111010", --  834 - 0x342  :  250 - 0xfa
    "11111010", --  835 - 0x343  :  250 - 0xfa
    "11111010", --  836 - 0x344  :  250 - 0xfa
    "11111010", --  837 - 0x345  :  250 - 0xfa
    "11111010", --  838 - 0x346  :  250 - 0xfa
    "11111010", --  839 - 0x347  :  250 - 0xfa
    "11111010", --  840 - 0x348  :  250 - 0xfa
    "11111010", --  841 - 0x349  :  250 - 0xfa
    "11111010", --  842 - 0x34a  :  250 - 0xfa
    "11111010", --  843 - 0x34b  :  250 - 0xfa
    "11111010", --  844 - 0x34c  :  250 - 0xfa
    "11111010", --  845 - 0x34d  :  250 - 0xfa
    "11111010", --  846 - 0x34e  :  250 - 0xfa
    "11111010", --  847 - 0x34f  :  250 - 0xfa
    "11111010", --  848 - 0x350  :  250 - 0xfa
    "11111010", --  849 - 0x351  :  250 - 0xfa
    "11111010", --  850 - 0x352  :  250 - 0xfa
    "11111010", --  851 - 0x353  :  250 - 0xfa
    "11111010", --  852 - 0x354  :  250 - 0xfa
    "11111010", --  853 - 0x355  :  250 - 0xfa
    "11111010", --  854 - 0x356  :  250 - 0xfa
    "11111010", --  855 - 0x357  :  250 - 0xfa
    "11111010", --  856 - 0x358  :  250 - 0xfa
    "11111010", --  857 - 0x359  :  250 - 0xfa
    "11111010", --  858 - 0x35a  :  250 - 0xfa
    "11111010", --  859 - 0x35b  :  250 - 0xfa
    "11111010", --  860 - 0x35c  :  250 - 0xfa
    "11111010", --  861 - 0x35d  :  250 - 0xfa
    "11111010", --  862 - 0x35e  :  250 - 0xfa
    "11111010", --  863 - 0x35f  :  250 - 0xfa
    "11111010", --  864 - 0x360  :  250 - 0xfa -- line 0x1b
    "11111010", --  865 - 0x361  :  250 - 0xfa
    "11111010", --  866 - 0x362  :  250 - 0xfa
    "11111010", --  867 - 0x363  :  250 - 0xfa
    "11111010", --  868 - 0x364  :  250 - 0xfa
    "11111010", --  869 - 0x365  :  250 - 0xfa
    "11111010", --  870 - 0x366  :  250 - 0xfa
    "11111010", --  871 - 0x367  :  250 - 0xfa
    "11111010", --  872 - 0x368  :  250 - 0xfa
    "00101011", --  873 - 0x369  :   43 - 0x2b
    "00101010", --  874 - 0x36a  :   42 - 0x2a
    "00000110", --  875 - 0x36b  :    6 - 0x6
    "00100110", --  876 - 0x36c  :   38 - 0x26
    "11111010", --  877 - 0x36d  :  250 - 0xfa
    "00010000", --  878 - 0x36e  :   16 - 0x10
    "11111010", --  879 - 0x36f  :  250 - 0xfa
    "00010011", --  880 - 0x370  :   19 - 0x13
    "00011101", --  881 - 0x371  :   29 - 0x1d
    "00100010", --  882 - 0x372  :   34 - 0x22
    "00011110", --  883 - 0x373  :   30 - 0x1e
    "00001010", --  884 - 0x374  :   10 - 0xa
    "00011001", --  885 - 0x375  :   25 - 0x19
    "00011111", --  886 - 0x376  :   31 - 0x1f
    "11111010", --  887 - 0x377  :  250 - 0xfa
    "11111010", --  888 - 0x378  :  250 - 0xfa
    "11111010", --  889 - 0x379  :  250 - 0xfa
    "11101010", --  890 - 0x37a  :  234 - 0xea
    "11111010", --  891 - 0x37b  :  250 - 0xfa
    "11111010", --  892 - 0x37c  :  250 - 0xfa
    "11111010", --  893 - 0x37d  :  250 - 0xfa
    "11111010", --  894 - 0x37e  :  250 - 0xfa
    "11111010", --  895 - 0x37f  :  250 - 0xfa
    "11111010", --  896 - 0x380  :  250 - 0xfa -- line 0x1c
    "11111010", --  897 - 0x381  :  250 - 0xfa
    "11111010", --  898 - 0x382  :  250 - 0xfa
    "11111010", --  899 - 0x383  :  250 - 0xfa
    "11111010", --  900 - 0x384  :  250 - 0xfa
    "11101010", --  901 - 0x385  :  234 - 0xea
    "11111010", --  902 - 0x386  :  250 - 0xfa
    "11111010", --  903 - 0x387  :  250 - 0xfa
    "11111010", --  904 - 0x388  :  250 - 0xfa
    "11101001", --  905 - 0x389  :  233 - 0xe9
    "11111010", --  906 - 0x38a  :  250 - 0xfa
    "11111010", --  907 - 0x38b  :  250 - 0xfa
    "11111010", --  908 - 0x38c  :  250 - 0xfa
    "11111010", --  909 - 0x38d  :  250 - 0xfa
    "11111010", --  910 - 0x38e  :  250 - 0xfa
    "11111010", --  911 - 0x38f  :  250 - 0xfa
    "11111010", --  912 - 0x390  :  250 - 0xfa
    "11111010", --  913 - 0x391  :  250 - 0xfa
    "11111010", --  914 - 0x392  :  250 - 0xfa
    "11111010", --  915 - 0x393  :  250 - 0xfa
    "11111010", --  916 - 0x394  :  250 - 0xfa
    "11111010", --  917 - 0x395  :  250 - 0xfa
    "11111010", --  918 - 0x396  :  250 - 0xfa
    "11111010", --  919 - 0x397  :  250 - 0xfa
    "11111010", --  920 - 0x398  :  250 - 0xfa
    "11111010", --  921 - 0x399  :  250 - 0xfa
    "11111010", --  922 - 0x39a  :  250 - 0xfa
    "11111010", --  923 - 0x39b  :  250 - 0xfa
    "11111010", --  924 - 0x39c  :  250 - 0xfa
    "11111010", --  925 - 0x39d  :  250 - 0xfa
    "11111001", --  926 - 0x39e  :  249 - 0xf9
    "11111010", --  927 - 0x39f  :  250 - 0xfa
    "11111010", --  928 - 0x3a0  :  250 - 0xfa -- line 0x1d
    "11111001", --  929 - 0x3a1  :  249 - 0xf9
    "11111010", --  930 - 0x3a2  :  250 - 0xfa
    "11111010", --  931 - 0x3a3  :  250 - 0xfa
    "11111010", --  932 - 0x3a4  :  250 - 0xfa
    "11111010", --  933 - 0x3a5  :  250 - 0xfa
    "11111010", --  934 - 0x3a6  :  250 - 0xfa
    "11111010", --  935 - 0x3a7  :  250 - 0xfa
    "11111010", --  936 - 0x3a8  :  250 - 0xfa
    "11111010", --  937 - 0x3a9  :  250 - 0xfa
    "11111010", --  938 - 0x3aa  :  250 - 0xfa
    "11111010", --  939 - 0x3ab  :  250 - 0xfa
    "11111010", --  940 - 0x3ac  :  250 - 0xfa
    "11111010", --  941 - 0x3ad  :  250 - 0xfa
    "11111010", --  942 - 0x3ae  :  250 - 0xfa
    "11111010", --  943 - 0x3af  :  250 - 0xfa
    "11111010", --  944 - 0x3b0  :  250 - 0xfa
    "11111010", --  945 - 0x3b1  :  250 - 0xfa
    "11111010", --  946 - 0x3b2  :  250 - 0xfa
    "11111010", --  947 - 0x3b3  :  250 - 0xfa
    "11111010", --  948 - 0x3b4  :  250 - 0xfa
    "11111010", --  949 - 0x3b5  :  250 - 0xfa
    "11111010", --  950 - 0x3b6  :  250 - 0xfa
    "11111010", --  951 - 0x3b7  :  250 - 0xfa
    "11111010", --  952 - 0x3b8  :  250 - 0xfa
    "11111010", --  953 - 0x3b9  :  250 - 0xfa
    "11111010", --  954 - 0x3ba  :  250 - 0xfa
    "11111010", --  955 - 0x3bb  :  250 - 0xfa
    "11111010", --  956 - 0x3bc  :  250 - 0xfa
    "11111010", --  957 - 0x3bd  :  250 - 0xfa
    "11111010", --  958 - 0x3be  :  250 - 0xfa
    "11111010", --  959 - 0x3bf  :  250 - 0xfa
        ---- Attribute Table 0----
    "01010101", --  960 - 0x3c0  :   85 - 0x55
    "01010101", --  961 - 0x3c1  :   85 - 0x55
    "01010101", --  962 - 0x3c2  :   85 - 0x55
    "01010101", --  963 - 0x3c3  :   85 - 0x55
    "01010101", --  964 - 0x3c4  :   85 - 0x55
    "01010101", --  965 - 0x3c5  :   85 - 0x55
    "01010101", --  966 - 0x3c6  :   85 - 0x55
    "01010101", --  967 - 0x3c7  :   85 - 0x55
    "00000000", --  968 - 0x3c8  :    0 - 0x0
    "00000000", --  969 - 0x3c9  :    0 - 0x0
    "00000000", --  970 - 0x3ca  :    0 - 0x0
    "00000000", --  971 - 0x3cb  :    0 - 0x0
    "00000000", --  972 - 0x3cc  :    0 - 0x0
    "00000000", --  973 - 0x3cd  :    0 - 0x0
    "00000000", --  974 - 0x3ce  :    0 - 0x0
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "01010101", --  976 - 0x3d0  :   85 - 0x55
    "01010101", --  977 - 0x3d1  :   85 - 0x55
    "01010101", --  978 - 0x3d2  :   85 - 0x55
    "01010101", --  979 - 0x3d3  :   85 - 0x55
    "01010101", --  980 - 0x3d4  :   85 - 0x55
    "01010101", --  981 - 0x3d5  :   85 - 0x55
    "01010101", --  982 - 0x3d6  :   85 - 0x55
    "01010101", --  983 - 0x3d7  :   85 - 0x55
    "01010101", --  984 - 0x3d8  :   85 - 0x55
    "01010101", --  985 - 0x3d9  :   85 - 0x55
    "01010101", --  986 - 0x3da  :   85 - 0x55
    "01010101", --  987 - 0x3db  :   85 - 0x55
    "01010101", --  988 - 0x3dc  :   85 - 0x55
    "01010101", --  989 - 0x3dd  :   85 - 0x55
    "01010101", --  990 - 0x3de  :   85 - 0x55
    "01010101", --  991 - 0x3df  :   85 - 0x55
    "01010101", --  992 - 0x3e0  :   85 - 0x55
    "01010101", --  993 - 0x3e1  :   85 - 0x55
    "01010101", --  994 - 0x3e2  :   85 - 0x55
    "01010101", --  995 - 0x3e3  :   85 - 0x55
    "01010101", --  996 - 0x3e4  :   85 - 0x55
    "01010101", --  997 - 0x3e5  :   85 - 0x55
    "01010101", --  998 - 0x3e6  :   85 - 0x55
    "01010101", --  999 - 0x3e7  :   85 - 0x55
    "01010101", -- 1000 - 0x3e8  :   85 - 0x55
    "01010101", -- 1001 - 0x3e9  :   85 - 0x55
    "01010101", -- 1002 - 0x3ea  :   85 - 0x55
    "01010101", -- 1003 - 0x3eb  :   85 - 0x55
    "01010101", -- 1004 - 0x3ec  :   85 - 0x55
    "01010101", -- 1005 - 0x3ed  :   85 - 0x55
    "01010101", -- 1006 - 0x3ee  :   85 - 0x55
    "01010101", -- 1007 - 0x3ef  :   85 - 0x55
    "01010101", -- 1008 - 0x3f0  :   85 - 0x55
    "01010101", -- 1009 - 0x3f1  :   85 - 0x55
    "01010101", -- 1010 - 0x3f2  :   85 - 0x55
    "01010101", -- 1011 - 0x3f3  :   85 - 0x55
    "01010101", -- 1012 - 0x3f4  :   85 - 0x55
    "01010101", -- 1013 - 0x3f5  :   85 - 0x55
    "01010101", -- 1014 - 0x3f6  :   85 - 0x55
    "01010101", -- 1015 - 0x3f7  :   85 - 0x55
    "00000101", -- 1016 - 0x3f8  :    5 - 0x5
    "00000101", -- 1017 - 0x3f9  :    5 - 0x5
    "00000101", -- 1018 - 0x3fa  :    5 - 0x5
    "00000101", -- 1019 - 0x3fb  :    5 - 0x5
    "00000101", -- 1020 - 0x3fc  :    5 - 0x5
    "00000101", -- 1021 - 0x3fd  :    5 - 0x5
    "00000101", -- 1022 - 0x3fe  :    5 - 0x5
    "00000101"  -- 1023 - 0x3ff  :    5 - 0x5
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
