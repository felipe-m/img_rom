--- Autcmatically generated VHDL ROM from a NES memory file----
---   SPRITEs MEMORY (OAM)
-- https://wiki.nesdev.com/w/index.php/PPU_OAM


---  Original memory dump file name: donkeykong_oam.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory with clock ------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_OAM_DONKEYKONG is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(8-1 downto 0);  --256 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_OAM_DONKEYKONG;

architecture BEHAVIORAL of ROM_OAM_DONKEYKONG is
  signal addr_int  : natural range 0 to 2**8-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
    "01101011", --    0 -  0x0  :  107 - 0x6b -- Sprite 0x0
    "00000110", --    1 -  0x1  :    6 - 0x6
    "01000000", --    2 -  0x2  :   64 - 0x40
    "01110011", --    3 -  0x3  :  115 - 0x73
    "01110011", --    4 -  0x4  :  115 - 0x73 -- Sprite 0x1
    "00000111", --    5 -  0x5  :    7 - 0x7
    "01000000", --    6 -  0x6  :   64 - 0x40
    "01110011", --    7 -  0x7  :  115 - 0x73
    "01101011", --    8 -  0x8  :  107 - 0x6b -- Sprite 0x2
    "00000100", --    9 -  0x9  :    4 - 0x4
    "01000000", --   10 -  0xa  :   64 - 0x40
    "01111011", --   11 -  0xb  :  123 - 0x7b
    "01110011", --   12 -  0xc  :  115 - 0x73 -- Sprite 0x3
    "00000101", --   13 -  0xd  :    5 - 0x5
    "01000000", --   14 -  0xe  :   64 - 0x40
    "01111011", --   15 -  0xf  :  123 - 0x7b
    "10100101", --   16 - 0x10  :  165 - 0xa5 -- Sprite 0x4
    "10011010", --   17 - 0x11  :  154 - 0x9a
    "01000010", --   18 - 0x12  :   66 - 0x42
    "01001011", --   19 - 0x13  :   75 - 0x4b
    "10101101", --   20 - 0x14  :  173 - 0xad -- Sprite 0x5
    "10011011", --   21 - 0x15  :  155 - 0x9b
    "01000010", --   22 - 0x16  :   66 - 0x42
    "01001011", --   23 - 0x17  :   75 - 0x4b
    "10100101", --   24 - 0x18  :  165 - 0xa5 -- Sprite 0x6
    "10011000", --   25 - 0x19  :  152 - 0x98
    "01000010", --   26 - 0x1a  :   66 - 0x42
    "01010011", --   27 - 0x1b  :   83 - 0x53
    "10101101", --   28 - 0x1c  :  173 - 0xad -- Sprite 0x7
    "10011001", --   29 - 0x1d  :  153 - 0x99
    "01000010", --   30 - 0x1e  :   66 - 0x42
    "01010011", --   31 - 0x1f  :   83 - 0x53
    "11000111", --   32 - 0x20  :  199 - 0xc7 -- Sprite 0x8
    "10011110", --   33 - 0x21  :  158 - 0x9e
    "01000010", --   34 - 0x22  :   66 - 0x42
    "01001100", --   35 - 0x23  :   76 - 0x4c
    "11001111", --   36 - 0x24  :  207 - 0xcf -- Sprite 0x9
    "10011111", --   37 - 0x25  :  159 - 0x9f
    "01000010", --   38 - 0x26  :   66 - 0x42
    "01001100", --   39 - 0x27  :   76 - 0x4c
    "11000111", --   40 - 0x28  :  199 - 0xc7 -- Sprite 0xa
    "10011100", --   41 - 0x29  :  156 - 0x9c
    "01000010", --   42 - 0x2a  :   66 - 0x42
    "01010100", --   43 - 0x2b  :   84 - 0x54
    "11001111", --   44 - 0x2c  :  207 - 0xcf -- Sprite 0xb
    "10011101", --   45 - 0x2d  :  157 - 0x9d
    "01000010", --   46 - 0x2e  :   66 - 0x42
    "01010100", --   47 - 0x2f  :   84 - 0x54
    "10001010", --   48 - 0x30  :  138 - 0x8a -- Sprite 0xc
    "10001000", --   49 - 0x31  :  136 - 0x88
    "00000011", --   50 - 0x32  :    3 - 0x3
    "10111010", --   51 - 0x33  :  186 - 0xba
    "10010010", --   52 - 0x34  :  146 - 0x92 -- Sprite 0xd
    "10001001", --   53 - 0x35  :  137 - 0x89
    "00000011", --   54 - 0x36  :    3 - 0x3
    "10111010", --   55 - 0x37  :  186 - 0xba
    "10001010", --   56 - 0x38  :  138 - 0x8a -- Sprite 0xe
    "10001010", --   57 - 0x39  :  138 - 0x8a
    "00000011", --   58 - 0x3a  :    3 - 0x3
    "11000010", --   59 - 0x3b  :  194 - 0xc2
    "10010010", --   60 - 0x3c  :  146 - 0x92 -- Sprite 0xf
    "10001011", --   61 - 0x3d  :  139 - 0x8b
    "00000011", --   62 - 0x3e  :    3 - 0x3
    "11000010", --   63 - 0x3f  :  194 - 0xc2
    "10000111", --   64 - 0x40  :  135 - 0x87 -- Sprite 0x10
    "10001000", --   65 - 0x41  :  136 - 0x88
    "00000011", --   66 - 0x42  :    3 - 0x3
    "11100110", --   67 - 0x43  :  230 - 0xe6
    "10001111", --   68 - 0x44  :  143 - 0x8f -- Sprite 0x11
    "10001001", --   69 - 0x45  :  137 - 0x89
    "00000011", --   70 - 0x46  :    3 - 0x3
    "11100110", --   71 - 0x47  :  230 - 0xe6
    "10000111", --   72 - 0x48  :  135 - 0x87 -- Sprite 0x12
    "10001010", --   73 - 0x49  :  138 - 0x8a
    "00000011", --   74 - 0x4a  :    3 - 0x3
    "11101110", --   75 - 0x4b  :  238 - 0xee
    "10001111", --   76 - 0x4c  :  143 - 0x8f -- Sprite 0x13
    "10001011", --   77 - 0x4d  :  139 - 0x8b
    "00000011", --   78 - 0x4e  :    3 - 0x3
    "11101110", --   79 - 0x4f  :  238 - 0xee
    "01010011", --   80 - 0x50  :   83 - 0x53 -- Sprite 0x14
    "10000000", --   81 - 0x51  :  128 - 0x80
    "00000011", --   82 - 0x52  :    3 - 0x3
    "00110010", --   83 - 0x53  :   50 - 0x32
    "01011011", --   84 - 0x54  :   91 - 0x5b -- Sprite 0x15
    "10000001", --   85 - 0x55  :  129 - 0x81
    "00000011", --   86 - 0x56  :    3 - 0x3
    "00110010", --   87 - 0x57  :   50 - 0x32
    "01010011", --   88 - 0x58  :   83 - 0x53 -- Sprite 0x16
    "10000010", --   89 - 0x59  :  130 - 0x82
    "00000011", --   90 - 0x5a  :    3 - 0x3
    "00111010", --   91 - 0x5b  :   58 - 0x3a
    "01011011", --   92 - 0x5c  :   91 - 0x5b -- Sprite 0x17
    "10000011", --   93 - 0x5d  :  131 - 0x83
    "00000011", --   94 - 0x5e  :    3 - 0x3
    "00111010", --   95 - 0x5f  :   58 - 0x3a
    "01001001", --   96 - 0x60  :   73 - 0x49 -- Sprite 0x18
    "10001000", --   97 - 0x61  :  136 - 0x88
    "00000011", --   98 - 0x62  :    3 - 0x3
    "11011101", --   99 - 0x63  :  221 - 0xdd
    "01010001", --  100 - 0x64  :   81 - 0x51 -- Sprite 0x19
    "10001001", --  101 - 0x65  :  137 - 0x89
    "00000011", --  102 - 0x66  :    3 - 0x3
    "11011101", --  103 - 0x67  :  221 - 0xdd
    "01001001", --  104 - 0x68  :   73 - 0x49 -- Sprite 0x1a
    "10001010", --  105 - 0x69  :  138 - 0x8a
    "00000011", --  106 - 0x6a  :    3 - 0x3
    "11100101", --  107 - 0x6b  :  229 - 0xe5
    "01010001", --  108 - 0x6c  :   81 - 0x51 -- Sprite 0x1b
    "10001011", --  109 - 0x6d  :  139 - 0x8b
    "00000011", --  110 - 0x6e  :    3 - 0x3
    "11100101", --  111 - 0x6f  :  229 - 0xe5
    "00110010", --  112 - 0x70  :   50 - 0x32 -- Sprite 0x1c
    "10000100", --  113 - 0x71  :  132 - 0x84
    "00000011", --  114 - 0x72  :    3 - 0x3
    "01001101", --  115 - 0x73  :   77 - 0x4d
    "00111010", --  116 - 0x74  :   58 - 0x3a -- Sprite 0x1d
    "10000101", --  117 - 0x75  :  133 - 0x85
    "00000011", --  118 - 0x76  :    3 - 0x3
    "01001101", --  119 - 0x77  :   77 - 0x4d
    "00110010", --  120 - 0x78  :   50 - 0x32 -- Sprite 0x1e
    "10000110", --  121 - 0x79  :  134 - 0x86
    "00000011", --  122 - 0x7a  :    3 - 0x3
    "01010101", --  123 - 0x7b  :   85 - 0x55
    "00111010", --  124 - 0x7c  :   58 - 0x3a -- Sprite 0x1f
    "10000111", --  125 - 0x7d  :  135 - 0x87
    "00000011", --  126 - 0x7e  :    3 - 0x3
    "01010101", --  127 - 0x7f  :   85 - 0x55
    "11111111", --  128 - 0x80  :  255 - 0xff -- Sprite 0x20
    "00000000", --  129 - 0x81  :    0 - 0x0
    "00000011", --  130 - 0x82  :    3 - 0x3
    "00000000", --  131 - 0x83  :    0 - 0x0
    "11111111", --  132 - 0x84  :  255 - 0xff -- Sprite 0x21
    "00000000", --  133 - 0x85  :    0 - 0x0
    "00000011", --  134 - 0x86  :    3 - 0x3
    "00000000", --  135 - 0x87  :    0 - 0x0
    "11111111", --  136 - 0x88  :  255 - 0xff -- Sprite 0x22
    "00000000", --  137 - 0x89  :    0 - 0x0
    "00000011", --  138 - 0x8a  :    3 - 0x3
    "00000000", --  139 - 0x8b  :    0 - 0x0
    "11111111", --  140 - 0x8c  :  255 - 0xff -- Sprite 0x23
    "00000000", --  141 - 0x8d  :    0 - 0x0
    "00000011", --  142 - 0x8e  :    3 - 0x3
    "00000000", --  143 - 0x8f  :    0 - 0x0
    "11111111", --  144 - 0x90  :  255 - 0xff -- Sprite 0x24
    "00000000", --  145 - 0x91  :    0 - 0x0
    "00000011", --  146 - 0x92  :    3 - 0x3
    "00000000", --  147 - 0x93  :    0 - 0x0
    "11111111", --  148 - 0x94  :  255 - 0xff -- Sprite 0x25
    "00000000", --  149 - 0x95  :    0 - 0x0
    "00000011", --  150 - 0x96  :    3 - 0x3
    "00000000", --  151 - 0x97  :    0 - 0x0
    "11111111", --  152 - 0x98  :  255 - 0xff -- Sprite 0x26
    "00000000", --  153 - 0x99  :    0 - 0x0
    "00000011", --  154 - 0x9a  :    3 - 0x3
    "00000000", --  155 - 0x9b  :    0 - 0x0
    "11111111", --  156 - 0x9c  :  255 - 0xff -- Sprite 0x27
    "00000000", --  157 - 0x9d  :    0 - 0x0
    "00000011", --  158 - 0x9e  :    3 - 0x3
    "00000000", --  159 - 0x9f  :    0 - 0x0
    "11111111", --  160 - 0xa0  :  255 - 0xff -- Sprite 0x28
    "00000000", --  161 - 0xa1  :    0 - 0x0
    "00000011", --  162 - 0xa2  :    3 - 0x3
    "00000000", --  163 - 0xa3  :    0 - 0x0
    "11111111", --  164 - 0xa4  :  255 - 0xff -- Sprite 0x29
    "00000000", --  165 - 0xa5  :    0 - 0x0
    "00000011", --  166 - 0xa6  :    3 - 0x3
    "00000000", --  167 - 0xa7  :    0 - 0x0
    "11111111", --  168 - 0xa8  :  255 - 0xff -- Sprite 0x2a
    "00000000", --  169 - 0xa9  :    0 - 0x0
    "00000011", --  170 - 0xaa  :    3 - 0x3
    "00000000", --  171 - 0xab  :    0 - 0x0
    "11111111", --  172 - 0xac  :  255 - 0xff -- Sprite 0x2b
    "00000000", --  173 - 0xad  :    0 - 0x0
    "00000011", --  174 - 0xae  :    3 - 0x3
    "00000000", --  175 - 0xaf  :    0 - 0x0
    "11111111", --  176 - 0xb0  :  255 - 0xff -- Sprite 0x2c
    "00000000", --  177 - 0xb1  :    0 - 0x0
    "00000011", --  178 - 0xb2  :    3 - 0x3
    "00000000", --  179 - 0xb3  :    0 - 0x0
    "11111111", --  180 - 0xb4  :  255 - 0xff -- Sprite 0x2d
    "00000000", --  181 - 0xb5  :    0 - 0x0
    "00000011", --  182 - 0xb6  :    3 - 0x3
    "00000000", --  183 - 0xb7  :    0 - 0x0
    "11111111", --  184 - 0xb8  :  255 - 0xff -- Sprite 0x2e
    "00000000", --  185 - 0xb9  :    0 - 0x0
    "00000011", --  186 - 0xba  :    3 - 0x3
    "00000000", --  187 - 0xbb  :    0 - 0x0
    "11111111", --  188 - 0xbc  :  255 - 0xff -- Sprite 0x2f
    "00000000", --  189 - 0xbd  :    0 - 0x0
    "00000011", --  190 - 0xbe  :    3 - 0x3
    "00000000", --  191 - 0xbf  :    0 - 0x0
    "11111111", --  192 - 0xc0  :  255 - 0xff -- Sprite 0x30
    "11010000", --  193 - 0xc1  :  208 - 0xd0
    "00000001", --  194 - 0xc2  :    1 - 0x1
    "01110100", --  195 - 0xc3  :  116 - 0x74
    "11111111", --  196 - 0xc4  :  255 - 0xff -- Sprite 0x31
    "11010100", --  197 - 0xc5  :  212 - 0xd4
    "00000001", --  198 - 0xc6  :    1 - 0x1
    "01111100", --  199 - 0xc7  :  124 - 0x7c
    "11111111", --  200 - 0xc8  :  255 - 0xff -- Sprite 0x32
    "00000000", --  201 - 0xc9  :    0 - 0x0
    "00000001", --  202 - 0xca  :    1 - 0x1
    "00000000", --  203 - 0xcb  :    0 - 0x0
    "11111111", --  204 - 0xcc  :  255 - 0xff -- Sprite 0x33
    "00000000", --  205 - 0xcd  :    0 - 0x0
    "00000001", --  206 - 0xce  :    1 - 0x1
    "00000000", --  207 - 0xcf  :    0 - 0x0
    "11111111", --  208 - 0xd0  :  255 - 0xff -- Sprite 0x34
    "11110110", --  209 - 0xd1  :  246 - 0xf6
    "00000011", --  210 - 0xd2  :    3 - 0x3
    "10100110", --  211 - 0xd3  :  166 - 0xa6
    "11111111", --  212 - 0xd4  :  255 - 0xff -- Sprite 0x35
    "11110111", --  213 - 0xd5  :  247 - 0xf7
    "00000011", --  214 - 0xd6  :    3 - 0x3
    "10100110", --  215 - 0xd7  :  166 - 0xa6
    "01000110", --  216 - 0xd8  :   70 - 0x46 -- Sprite 0x36
    "11110110", --  217 - 0xd9  :  246 - 0xf6
    "00000011", --  218 - 0xda  :    3 - 0x3
    "00100000", --  219 - 0xdb  :   32 - 0x20
    "01001110", --  220 - 0xdc  :   78 - 0x4e -- Sprite 0x37
    "11110111", --  221 - 0xdd  :  247 - 0xf7
    "00000011", --  222 - 0xde  :    3 - 0x3
    "00100000", --  223 - 0xdf  :   32 - 0x20
    "11000000", --  224 - 0xe0  :  192 - 0xc0 -- Sprite 0x38
    "11111110", --  225 - 0xe1  :  254 - 0xfe
    "00000010", --  226 - 0xe2  :    2 - 0x2
    "00100000", --  227 - 0xe3  :   32 - 0x20
    "11000000", --  228 - 0xe4  :  192 - 0xc0 -- Sprite 0x39
    "11111111", --  229 - 0xe5  :  255 - 0xff
    "00000010", --  230 - 0xe6  :    2 - 0x2
    "00101000", --  231 - 0xe7  :   40 - 0x28
    "00011000", --  232 - 0xe8  :   24 - 0x18 -- Sprite 0x3a
    "11010101", --  233 - 0xe9  :  213 - 0xd5
    "00000001", --  234 - 0xea  :    1 - 0x1
    "01010000", --  235 - 0xeb  :   80 - 0x50
    "00011000", --  236 - 0xec  :   24 - 0x18 -- Sprite 0x3b
    "11010110", --  237 - 0xed  :  214 - 0xd6
    "00000001", --  238 - 0xee  :    1 - 0x1
    "01011000", --  239 - 0xef  :   88 - 0x58
    "00100000", --  240 - 0xf0  :   32 - 0x20 -- Sprite 0x3c
    "11011011", --  241 - 0xf1  :  219 - 0xdb
    "00000001", --  242 - 0xf2  :    1 - 0x1
    "01010000", --  243 - 0xf3  :   80 - 0x50
    "00101000", --  244 - 0xf4  :   40 - 0x28 -- Sprite 0x3d
    "11011100", --  245 - 0xf5  :  220 - 0xdc
    "00000001", --  246 - 0xf6  :    1 - 0x1
    "01010000", --  247 - 0xf7  :   80 - 0x50
    "00100000", --  248 - 0xf8  :   32 - 0x20 -- Sprite 0x3e
    "11011101", --  249 - 0xf9  :  221 - 0xdd
    "00000001", --  250 - 0xfa  :    1 - 0x1
    "01011000", --  251 - 0xfb  :   88 - 0x58
    "00101000", --  252 - 0xfc  :   40 - 0x28 -- Sprite 0x3f
    "11011110", --  253 - 0xfd  :  222 - 0xde
    "00000001", --  254 - 0xfe  :    1 - 0x1
    "01011000"  --  255 - 0xff  :   88 - 0x58
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
