---   Background Pattern table COLOR PLANE 1
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
--- Autcmatically generated VHDL ROM from a NES memory file----


---  Original memory dump file name: donkeykong_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory with clock ------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_DONKEYKONG_BG_PLN1 is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(11-1 downto 0);  --2048 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_DONKEYKONG_BG_PLN1;

architecture BEHAVIORAL of ROM_PTABLE_DONKEYKONG_BG_PLN1 is
  signal addr_int  : natural range 0 to 2**11-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Background pattern Table COLOR PLANE 1
    "00000000", --    0 -  0x0  :    0 - 0x0 -- Background 0x0
    "00000000", --    1 -  0x1  :    0 - 0x0
    "00000000", --    2 -  0x2  :    0 - 0x0
    "00000000", --    3 -  0x3  :    0 - 0x0
    "00000000", --    4 -  0x4  :    0 - 0x0
    "00000000", --    5 -  0x5  :    0 - 0x0
    "00000000", --    6 -  0x6  :    0 - 0x0
    "00000000", --    7 -  0x7  :    0 - 0x0
    "00000000", --    8 -  0x8  :    0 - 0x0 -- Background 0x1
    "00000000", --    9 -  0x9  :    0 - 0x0
    "00000000", --   10 -  0xa  :    0 - 0x0
    "00000000", --   11 -  0xb  :    0 - 0x0
    "00000000", --   12 -  0xc  :    0 - 0x0
    "00000000", --   13 -  0xd  :    0 - 0x0
    "00000000", --   14 -  0xe  :    0 - 0x0
    "00000000", --   15 -  0xf  :    0 - 0x0
    "00000000", --   16 - 0x10  :    0 - 0x0 -- Background 0x2
    "00000000", --   17 - 0x11  :    0 - 0x0
    "00000000", --   18 - 0x12  :    0 - 0x0
    "00000000", --   19 - 0x13  :    0 - 0x0
    "00000000", --   20 - 0x14  :    0 - 0x0
    "00000000", --   21 - 0x15  :    0 - 0x0
    "00000000", --   22 - 0x16  :    0 - 0x0
    "00000000", --   23 - 0x17  :    0 - 0x0
    "00000000", --   24 - 0x18  :    0 - 0x0 -- Background 0x3
    "00000000", --   25 - 0x19  :    0 - 0x0
    "00000000", --   26 - 0x1a  :    0 - 0x0
    "00000000", --   27 - 0x1b  :    0 - 0x0
    "00000000", --   28 - 0x1c  :    0 - 0x0
    "00000000", --   29 - 0x1d  :    0 - 0x0
    "00000000", --   30 - 0x1e  :    0 - 0x0
    "00000000", --   31 - 0x1f  :    0 - 0x0
    "00000000", --   32 - 0x20  :    0 - 0x0 -- Background 0x4
    "00000000", --   33 - 0x21  :    0 - 0x0
    "00000000", --   34 - 0x22  :    0 - 0x0
    "00000000", --   35 - 0x23  :    0 - 0x0
    "00000000", --   36 - 0x24  :    0 - 0x0
    "00000000", --   37 - 0x25  :    0 - 0x0
    "00000000", --   38 - 0x26  :    0 - 0x0
    "00000000", --   39 - 0x27  :    0 - 0x0
    "00000000", --   40 - 0x28  :    0 - 0x0 -- Background 0x5
    "00000000", --   41 - 0x29  :    0 - 0x0
    "00000000", --   42 - 0x2a  :    0 - 0x0
    "00000000", --   43 - 0x2b  :    0 - 0x0
    "00000000", --   44 - 0x2c  :    0 - 0x0
    "00000000", --   45 - 0x2d  :    0 - 0x0
    "00000000", --   46 - 0x2e  :    0 - 0x0
    "00000000", --   47 - 0x2f  :    0 - 0x0
    "00000000", --   48 - 0x30  :    0 - 0x0 -- Background 0x6
    "00000000", --   49 - 0x31  :    0 - 0x0
    "00000000", --   50 - 0x32  :    0 - 0x0
    "00000000", --   51 - 0x33  :    0 - 0x0
    "00000000", --   52 - 0x34  :    0 - 0x0
    "00000000", --   53 - 0x35  :    0 - 0x0
    "00000000", --   54 - 0x36  :    0 - 0x0
    "00000000", --   55 - 0x37  :    0 - 0x0
    "00000000", --   56 - 0x38  :    0 - 0x0 -- Background 0x7
    "00000000", --   57 - 0x39  :    0 - 0x0
    "00000000", --   58 - 0x3a  :    0 - 0x0
    "00000000", --   59 - 0x3b  :    0 - 0x0
    "00000000", --   60 - 0x3c  :    0 - 0x0
    "00000000", --   61 - 0x3d  :    0 - 0x0
    "00000000", --   62 - 0x3e  :    0 - 0x0
    "00000000", --   63 - 0x3f  :    0 - 0x0
    "00000000", --   64 - 0x40  :    0 - 0x0 -- Background 0x8
    "00000000", --   65 - 0x41  :    0 - 0x0
    "00000000", --   66 - 0x42  :    0 - 0x0
    "00000000", --   67 - 0x43  :    0 - 0x0
    "00000000", --   68 - 0x44  :    0 - 0x0
    "00000000", --   69 - 0x45  :    0 - 0x0
    "00000000", --   70 - 0x46  :    0 - 0x0
    "00000000", --   71 - 0x47  :    0 - 0x0
    "00000000", --   72 - 0x48  :    0 - 0x0 -- Background 0x9
    "00000000", --   73 - 0x49  :    0 - 0x0
    "00000000", --   74 - 0x4a  :    0 - 0x0
    "00000000", --   75 - 0x4b  :    0 - 0x0
    "00000000", --   76 - 0x4c  :    0 - 0x0
    "00000000", --   77 - 0x4d  :    0 - 0x0
    "00000000", --   78 - 0x4e  :    0 - 0x0
    "00000000", --   79 - 0x4f  :    0 - 0x0
    "00000000", --   80 - 0x50  :    0 - 0x0 -- Background 0xa
    "00000000", --   81 - 0x51  :    0 - 0x0
    "00000000", --   82 - 0x52  :    0 - 0x0
    "00000000", --   83 - 0x53  :    0 - 0x0
    "00000000", --   84 - 0x54  :    0 - 0x0
    "00000000", --   85 - 0x55  :    0 - 0x0
    "00000000", --   86 - 0x56  :    0 - 0x0
    "00000000", --   87 - 0x57  :    0 - 0x0
    "00000000", --   88 - 0x58  :    0 - 0x0 -- Background 0xb
    "00000000", --   89 - 0x59  :    0 - 0x0
    "00000000", --   90 - 0x5a  :    0 - 0x0
    "00000000", --   91 - 0x5b  :    0 - 0x0
    "00000000", --   92 - 0x5c  :    0 - 0x0
    "00000000", --   93 - 0x5d  :    0 - 0x0
    "00000000", --   94 - 0x5e  :    0 - 0x0
    "00000000", --   95 - 0x5f  :    0 - 0x0
    "00000000", --   96 - 0x60  :    0 - 0x0 -- Background 0xc
    "00000000", --   97 - 0x61  :    0 - 0x0
    "00000000", --   98 - 0x62  :    0 - 0x0
    "00000000", --   99 - 0x63  :    0 - 0x0
    "00000000", --  100 - 0x64  :    0 - 0x0
    "00000000", --  101 - 0x65  :    0 - 0x0
    "00000000", --  102 - 0x66  :    0 - 0x0
    "00000000", --  103 - 0x67  :    0 - 0x0
    "00000000", --  104 - 0x68  :    0 - 0x0 -- Background 0xd
    "00000000", --  105 - 0x69  :    0 - 0x0
    "00000000", --  106 - 0x6a  :    0 - 0x0
    "00000000", --  107 - 0x6b  :    0 - 0x0
    "00000000", --  108 - 0x6c  :    0 - 0x0
    "00000000", --  109 - 0x6d  :    0 - 0x0
    "00000000", --  110 - 0x6e  :    0 - 0x0
    "00000000", --  111 - 0x6f  :    0 - 0x0
    "00000000", --  112 - 0x70  :    0 - 0x0 -- Background 0xe
    "00000000", --  113 - 0x71  :    0 - 0x0
    "00000000", --  114 - 0x72  :    0 - 0x0
    "00000000", --  115 - 0x73  :    0 - 0x0
    "00000000", --  116 - 0x74  :    0 - 0x0
    "00000000", --  117 - 0x75  :    0 - 0x0
    "00000000", --  118 - 0x76  :    0 - 0x0
    "00000000", --  119 - 0x77  :    0 - 0x0
    "00000000", --  120 - 0x78  :    0 - 0x0 -- Background 0xf
    "00000000", --  121 - 0x79  :    0 - 0x0
    "00000000", --  122 - 0x7a  :    0 - 0x0
    "00000000", --  123 - 0x7b  :    0 - 0x0
    "00000000", --  124 - 0x7c  :    0 - 0x0
    "00000000", --  125 - 0x7d  :    0 - 0x0
    "00000000", --  126 - 0x7e  :    0 - 0x0
    "00000000", --  127 - 0x7f  :    0 - 0x0
    "00000000", --  128 - 0x80  :    0 - 0x0 -- Background 0x10
    "00000000", --  129 - 0x81  :    0 - 0x0
    "00000000", --  130 - 0x82  :    0 - 0x0
    "00000000", --  131 - 0x83  :    0 - 0x0
    "00000000", --  132 - 0x84  :    0 - 0x0
    "00000000", --  133 - 0x85  :    0 - 0x0
    "00000000", --  134 - 0x86  :    0 - 0x0
    "00000000", --  135 - 0x87  :    0 - 0x0
    "00000000", --  136 - 0x88  :    0 - 0x0 -- Background 0x11
    "00000000", --  137 - 0x89  :    0 - 0x0
    "00000000", --  138 - 0x8a  :    0 - 0x0
    "00000000", --  139 - 0x8b  :    0 - 0x0
    "00000000", --  140 - 0x8c  :    0 - 0x0
    "00000000", --  141 - 0x8d  :    0 - 0x0
    "00000000", --  142 - 0x8e  :    0 - 0x0
    "00000000", --  143 - 0x8f  :    0 - 0x0
    "00000000", --  144 - 0x90  :    0 - 0x0 -- Background 0x12
    "00000000", --  145 - 0x91  :    0 - 0x0
    "00000000", --  146 - 0x92  :    0 - 0x0
    "00000000", --  147 - 0x93  :    0 - 0x0
    "00000000", --  148 - 0x94  :    0 - 0x0
    "00000000", --  149 - 0x95  :    0 - 0x0
    "00000000", --  150 - 0x96  :    0 - 0x0
    "00000000", --  151 - 0x97  :    0 - 0x0
    "00000000", --  152 - 0x98  :    0 - 0x0 -- Background 0x13
    "00000000", --  153 - 0x99  :    0 - 0x0
    "00000000", --  154 - 0x9a  :    0 - 0x0
    "00000000", --  155 - 0x9b  :    0 - 0x0
    "00000000", --  156 - 0x9c  :    0 - 0x0
    "00000000", --  157 - 0x9d  :    0 - 0x0
    "00000000", --  158 - 0x9e  :    0 - 0x0
    "00000000", --  159 - 0x9f  :    0 - 0x0
    "00000000", --  160 - 0xa0  :    0 - 0x0 -- Background 0x14
    "00000000", --  161 - 0xa1  :    0 - 0x0
    "00000000", --  162 - 0xa2  :    0 - 0x0
    "00000000", --  163 - 0xa3  :    0 - 0x0
    "00000000", --  164 - 0xa4  :    0 - 0x0
    "00000000", --  165 - 0xa5  :    0 - 0x0
    "00000000", --  166 - 0xa6  :    0 - 0x0
    "00000000", --  167 - 0xa7  :    0 - 0x0
    "00000000", --  168 - 0xa8  :    0 - 0x0 -- Background 0x15
    "00000000", --  169 - 0xa9  :    0 - 0x0
    "00000000", --  170 - 0xaa  :    0 - 0x0
    "00000000", --  171 - 0xab  :    0 - 0x0
    "00000000", --  172 - 0xac  :    0 - 0x0
    "00000000", --  173 - 0xad  :    0 - 0x0
    "00000000", --  174 - 0xae  :    0 - 0x0
    "00000000", --  175 - 0xaf  :    0 - 0x0
    "00000000", --  176 - 0xb0  :    0 - 0x0 -- Background 0x16
    "00000000", --  177 - 0xb1  :    0 - 0x0
    "00000000", --  178 - 0xb2  :    0 - 0x0
    "00000000", --  179 - 0xb3  :    0 - 0x0
    "00000000", --  180 - 0xb4  :    0 - 0x0
    "00000000", --  181 - 0xb5  :    0 - 0x0
    "00000000", --  182 - 0xb6  :    0 - 0x0
    "00000000", --  183 - 0xb7  :    0 - 0x0
    "00000000", --  184 - 0xb8  :    0 - 0x0 -- Background 0x17
    "00000000", --  185 - 0xb9  :    0 - 0x0
    "00000000", --  186 - 0xba  :    0 - 0x0
    "00000000", --  187 - 0xbb  :    0 - 0x0
    "00000000", --  188 - 0xbc  :    0 - 0x0
    "00000000", --  189 - 0xbd  :    0 - 0x0
    "00000000", --  190 - 0xbe  :    0 - 0x0
    "00000000", --  191 - 0xbf  :    0 - 0x0
    "00000000", --  192 - 0xc0  :    0 - 0x0 -- Background 0x18
    "00000000", --  193 - 0xc1  :    0 - 0x0
    "00000000", --  194 - 0xc2  :    0 - 0x0
    "00000000", --  195 - 0xc3  :    0 - 0x0
    "00000000", --  196 - 0xc4  :    0 - 0x0
    "00000000", --  197 - 0xc5  :    0 - 0x0
    "00000000", --  198 - 0xc6  :    0 - 0x0
    "00000000", --  199 - 0xc7  :    0 - 0x0
    "00000000", --  200 - 0xc8  :    0 - 0x0 -- Background 0x19
    "00000000", --  201 - 0xc9  :    0 - 0x0
    "00000000", --  202 - 0xca  :    0 - 0x0
    "00000000", --  203 - 0xcb  :    0 - 0x0
    "00000000", --  204 - 0xcc  :    0 - 0x0
    "00000000", --  205 - 0xcd  :    0 - 0x0
    "00000000", --  206 - 0xce  :    0 - 0x0
    "00000000", --  207 - 0xcf  :    0 - 0x0
    "00000000", --  208 - 0xd0  :    0 - 0x0 -- Background 0x1a
    "00000000", --  209 - 0xd1  :    0 - 0x0
    "00000000", --  210 - 0xd2  :    0 - 0x0
    "00000000", --  211 - 0xd3  :    0 - 0x0
    "00000000", --  212 - 0xd4  :    0 - 0x0
    "00000000", --  213 - 0xd5  :    0 - 0x0
    "00000000", --  214 - 0xd6  :    0 - 0x0
    "00000000", --  215 - 0xd7  :    0 - 0x0
    "00000000", --  216 - 0xd8  :    0 - 0x0 -- Background 0x1b
    "00000000", --  217 - 0xd9  :    0 - 0x0
    "00000000", --  218 - 0xda  :    0 - 0x0
    "00000000", --  219 - 0xdb  :    0 - 0x0
    "00000000", --  220 - 0xdc  :    0 - 0x0
    "00000000", --  221 - 0xdd  :    0 - 0x0
    "00000000", --  222 - 0xde  :    0 - 0x0
    "00000000", --  223 - 0xdf  :    0 - 0x0
    "00000000", --  224 - 0xe0  :    0 - 0x0 -- Background 0x1c
    "00000000", --  225 - 0xe1  :    0 - 0x0
    "00000000", --  226 - 0xe2  :    0 - 0x0
    "00000000", --  227 - 0xe3  :    0 - 0x0
    "00000000", --  228 - 0xe4  :    0 - 0x0
    "00000000", --  229 - 0xe5  :    0 - 0x0
    "00000000", --  230 - 0xe6  :    0 - 0x0
    "00000000", --  231 - 0xe7  :    0 - 0x0
    "00000000", --  232 - 0xe8  :    0 - 0x0 -- Background 0x1d
    "00000000", --  233 - 0xe9  :    0 - 0x0
    "00000000", --  234 - 0xea  :    0 - 0x0
    "00000000", --  235 - 0xeb  :    0 - 0x0
    "00000000", --  236 - 0xec  :    0 - 0x0
    "00000000", --  237 - 0xed  :    0 - 0x0
    "00000000", --  238 - 0xee  :    0 - 0x0
    "00000000", --  239 - 0xef  :    0 - 0x0
    "00000000", --  240 - 0xf0  :    0 - 0x0 -- Background 0x1e
    "00000000", --  241 - 0xf1  :    0 - 0x0
    "00000000", --  242 - 0xf2  :    0 - 0x0
    "00000000", --  243 - 0xf3  :    0 - 0x0
    "00000000", --  244 - 0xf4  :    0 - 0x0
    "00000000", --  245 - 0xf5  :    0 - 0x0
    "00000000", --  246 - 0xf6  :    0 - 0x0
    "00000000", --  247 - 0xf7  :    0 - 0x0
    "00000000", --  248 - 0xf8  :    0 - 0x0 -- Background 0x1f
    "00000000", --  249 - 0xf9  :    0 - 0x0
    "00000000", --  250 - 0xfa  :    0 - 0x0
    "00000000", --  251 - 0xfb  :    0 - 0x0
    "00000000", --  252 - 0xfc  :    0 - 0x0
    "00000000", --  253 - 0xfd  :    0 - 0x0
    "00000000", --  254 - 0xfe  :    0 - 0x0
    "00000000", --  255 - 0xff  :    0 - 0x0
    "00000000", --  256 - 0x100  :    0 - 0x0 -- Background 0x20
    "00000000", --  257 - 0x101  :    0 - 0x0
    "00000000", --  258 - 0x102  :    0 - 0x0
    "00000000", --  259 - 0x103  :    0 - 0x0
    "00000000", --  260 - 0x104  :    0 - 0x0
    "00000000", --  261 - 0x105  :    0 - 0x0
    "00000000", --  262 - 0x106  :    0 - 0x0
    "00000000", --  263 - 0x107  :    0 - 0x0
    "00000000", --  264 - 0x108  :    0 - 0x0 -- Background 0x21
    "00000000", --  265 - 0x109  :    0 - 0x0
    "00000000", --  266 - 0x10a  :    0 - 0x0
    "00000000", --  267 - 0x10b  :    0 - 0x0
    "00000000", --  268 - 0x10c  :    0 - 0x0
    "00000000", --  269 - 0x10d  :    0 - 0x0
    "00000000", --  270 - 0x10e  :    0 - 0x0
    "00000000", --  271 - 0x10f  :    0 - 0x0
    "00000000", --  272 - 0x110  :    0 - 0x0 -- Background 0x22
    "00000000", --  273 - 0x111  :    0 - 0x0
    "00000000", --  274 - 0x112  :    0 - 0x0
    "00000000", --  275 - 0x113  :    0 - 0x0
    "00000000", --  276 - 0x114  :    0 - 0x0
    "00000000", --  277 - 0x115  :    0 - 0x0
    "00000000", --  278 - 0x116  :    0 - 0x0
    "00000000", --  279 - 0x117  :    0 - 0x0
    "00000000", --  280 - 0x118  :    0 - 0x0 -- Background 0x23
    "00000000", --  281 - 0x119  :    0 - 0x0
    "00000000", --  282 - 0x11a  :    0 - 0x0
    "00000000", --  283 - 0x11b  :    0 - 0x0
    "00000000", --  284 - 0x11c  :    0 - 0x0
    "00000000", --  285 - 0x11d  :    0 - 0x0
    "00000000", --  286 - 0x11e  :    0 - 0x0
    "00000000", --  287 - 0x11f  :    0 - 0x0
    "00000000", --  288 - 0x120  :    0 - 0x0 -- Background 0x24
    "00000000", --  289 - 0x121  :    0 - 0x0
    "00000000", --  290 - 0x122  :    0 - 0x0
    "00000000", --  291 - 0x123  :    0 - 0x0
    "00000000", --  292 - 0x124  :    0 - 0x0
    "00000000", --  293 - 0x125  :    0 - 0x0
    "00000000", --  294 - 0x126  :    0 - 0x0
    "00000000", --  295 - 0x127  :    0 - 0x0
    "00000000", --  296 - 0x128  :    0 - 0x0 -- Background 0x25
    "00000000", --  297 - 0x129  :    0 - 0x0
    "00000000", --  298 - 0x12a  :    0 - 0x0
    "00000000", --  299 - 0x12b  :    0 - 0x0
    "00000000", --  300 - 0x12c  :    0 - 0x0
    "00000000", --  301 - 0x12d  :    0 - 0x0
    "00000000", --  302 - 0x12e  :    0 - 0x0
    "00000000", --  303 - 0x12f  :    0 - 0x0
    "00000000", --  304 - 0x130  :    0 - 0x0 -- Background 0x26
    "00000000", --  305 - 0x131  :    0 - 0x0
    "00000000", --  306 - 0x132  :    0 - 0x0
    "00000000", --  307 - 0x133  :    0 - 0x0
    "00000000", --  308 - 0x134  :    0 - 0x0
    "00000000", --  309 - 0x135  :    0 - 0x0
    "00000000", --  310 - 0x136  :    0 - 0x0
    "00000000", --  311 - 0x137  :    0 - 0x0
    "00000000", --  312 - 0x138  :    0 - 0x0 -- Background 0x27
    "00000000", --  313 - 0x139  :    0 - 0x0
    "00000000", --  314 - 0x13a  :    0 - 0x0
    "00000000", --  315 - 0x13b  :    0 - 0x0
    "00000000", --  316 - 0x13c  :    0 - 0x0
    "00000000", --  317 - 0x13d  :    0 - 0x0
    "00000000", --  318 - 0x13e  :    0 - 0x0
    "00000000", --  319 - 0x13f  :    0 - 0x0
    "00000000", --  320 - 0x140  :    0 - 0x0 -- Background 0x28
    "00000000", --  321 - 0x141  :    0 - 0x0
    "00000000", --  322 - 0x142  :    0 - 0x0
    "00000000", --  323 - 0x143  :    0 - 0x0
    "00000000", --  324 - 0x144  :    0 - 0x0
    "00000000", --  325 - 0x145  :    0 - 0x0
    "00000000", --  326 - 0x146  :    0 - 0x0
    "00000000", --  327 - 0x147  :    0 - 0x0
    "00000000", --  328 - 0x148  :    0 - 0x0 -- Background 0x29
    "00000000", --  329 - 0x149  :    0 - 0x0
    "00000000", --  330 - 0x14a  :    0 - 0x0
    "00000000", --  331 - 0x14b  :    0 - 0x0
    "00000000", --  332 - 0x14c  :    0 - 0x0
    "00000000", --  333 - 0x14d  :    0 - 0x0
    "00000000", --  334 - 0x14e  :    0 - 0x0
    "00000000", --  335 - 0x14f  :    0 - 0x0
    "00000000", --  336 - 0x150  :    0 - 0x0 -- Background 0x2a
    "00000000", --  337 - 0x151  :    0 - 0x0
    "00000000", --  338 - 0x152  :    0 - 0x0
    "00000000", --  339 - 0x153  :    0 - 0x0
    "00000000", --  340 - 0x154  :    0 - 0x0
    "00000000", --  341 - 0x155  :    0 - 0x0
    "00000000", --  342 - 0x156  :    0 - 0x0
    "00000000", --  343 - 0x157  :    0 - 0x0
    "00000000", --  344 - 0x158  :    0 - 0x0 -- Background 0x2b
    "00000000", --  345 - 0x159  :    0 - 0x0
    "00000000", --  346 - 0x15a  :    0 - 0x0
    "00000000", --  347 - 0x15b  :    0 - 0x0
    "00000000", --  348 - 0x15c  :    0 - 0x0
    "00000000", --  349 - 0x15d  :    0 - 0x0
    "00000000", --  350 - 0x15e  :    0 - 0x0
    "00000000", --  351 - 0x15f  :    0 - 0x0
    "00000000", --  352 - 0x160  :    0 - 0x0 -- Background 0x2c
    "00000000", --  353 - 0x161  :    0 - 0x0
    "00000000", --  354 - 0x162  :    0 - 0x0
    "00000000", --  355 - 0x163  :    0 - 0x0
    "00000000", --  356 - 0x164  :    0 - 0x0
    "00000000", --  357 - 0x165  :    0 - 0x0
    "00000000", --  358 - 0x166  :    0 - 0x0
    "00000000", --  359 - 0x167  :    0 - 0x0
    "00000000", --  360 - 0x168  :    0 - 0x0 -- Background 0x2d
    "00000000", --  361 - 0x169  :    0 - 0x0
    "00000000", --  362 - 0x16a  :    0 - 0x0
    "00000000", --  363 - 0x16b  :    0 - 0x0
    "00000000", --  364 - 0x16c  :    0 - 0x0
    "00000000", --  365 - 0x16d  :    0 - 0x0
    "00000000", --  366 - 0x16e  :    0 - 0x0
    "00000000", --  367 - 0x16f  :    0 - 0x0
    "00000000", --  368 - 0x170  :    0 - 0x0 -- Background 0x2e
    "00000000", --  369 - 0x171  :    0 - 0x0
    "00000000", --  370 - 0x172  :    0 - 0x0
    "00000000", --  371 - 0x173  :    0 - 0x0
    "00000000", --  372 - 0x174  :    0 - 0x0
    "00000000", --  373 - 0x175  :    0 - 0x0
    "00000000", --  374 - 0x176  :    0 - 0x0
    "00000000", --  375 - 0x177  :    0 - 0x0
    "00000000", --  376 - 0x178  :    0 - 0x0 -- Background 0x2f
    "00000000", --  377 - 0x179  :    0 - 0x0
    "00000000", --  378 - 0x17a  :    0 - 0x0
    "00000000", --  379 - 0x17b  :    0 - 0x0
    "00000000", --  380 - 0x17c  :    0 - 0x0
    "00000000", --  381 - 0x17d  :    0 - 0x0
    "00000000", --  382 - 0x17e  :    0 - 0x0
    "00000000", --  383 - 0x17f  :    0 - 0x0
    "00000000", --  384 - 0x180  :    0 - 0x0 -- Background 0x30
    "00000000", --  385 - 0x181  :    0 - 0x0
    "00000000", --  386 - 0x182  :    0 - 0x0
    "00000000", --  387 - 0x183  :    0 - 0x0
    "00000000", --  388 - 0x184  :    0 - 0x0
    "00000000", --  389 - 0x185  :    0 - 0x0
    "00000000", --  390 - 0x186  :    0 - 0x0
    "00000000", --  391 - 0x187  :    0 - 0x0
    "00000000", --  392 - 0x188  :    0 - 0x0 -- Background 0x31
    "00000000", --  393 - 0x189  :    0 - 0x0
    "00000000", --  394 - 0x18a  :    0 - 0x0
    "00000000", --  395 - 0x18b  :    0 - 0x0
    "00000000", --  396 - 0x18c  :    0 - 0x0
    "00000000", --  397 - 0x18d  :    0 - 0x0
    "00000000", --  398 - 0x18e  :    0 - 0x0
    "00000000", --  399 - 0x18f  :    0 - 0x0
    "00000000", --  400 - 0x190  :    0 - 0x0 -- Background 0x32
    "00000000", --  401 - 0x191  :    0 - 0x0
    "00000000", --  402 - 0x192  :    0 - 0x0
    "00000000", --  403 - 0x193  :    0 - 0x0
    "00000000", --  404 - 0x194  :    0 - 0x0
    "00000000", --  405 - 0x195  :    0 - 0x0
    "00000000", --  406 - 0x196  :    0 - 0x0
    "00000000", --  407 - 0x197  :    0 - 0x0
    "00000000", --  408 - 0x198  :    0 - 0x0 -- Background 0x33
    "00000000", --  409 - 0x199  :    0 - 0x0
    "00000000", --  410 - 0x19a  :    0 - 0x0
    "00000000", --  411 - 0x19b  :    0 - 0x0
    "00000000", --  412 - 0x19c  :    0 - 0x0
    "00000000", --  413 - 0x19d  :    0 - 0x0
    "00000000", --  414 - 0x19e  :    0 - 0x0
    "00000000", --  415 - 0x19f  :    0 - 0x0
    "00000000", --  416 - 0x1a0  :    0 - 0x0 -- Background 0x34
    "00000000", --  417 - 0x1a1  :    0 - 0x0
    "00000000", --  418 - 0x1a2  :    0 - 0x0
    "00000000", --  419 - 0x1a3  :    0 - 0x0
    "00000000", --  420 - 0x1a4  :    0 - 0x0
    "00000000", --  421 - 0x1a5  :    0 - 0x0
    "00000000", --  422 - 0x1a6  :    0 - 0x0
    "00000000", --  423 - 0x1a7  :    0 - 0x0
    "00000000", --  424 - 0x1a8  :    0 - 0x0 -- Background 0x35
    "00000000", --  425 - 0x1a9  :    0 - 0x0
    "00000000", --  426 - 0x1aa  :    0 - 0x0
    "00000000", --  427 - 0x1ab  :    0 - 0x0
    "00000000", --  428 - 0x1ac  :    0 - 0x0
    "00000000", --  429 - 0x1ad  :    0 - 0x0
    "00000000", --  430 - 0x1ae  :    0 - 0x0
    "00000000", --  431 - 0x1af  :    0 - 0x0
    "00000000", --  432 - 0x1b0  :    0 - 0x0 -- Background 0x36
    "00000000", --  433 - 0x1b1  :    0 - 0x0
    "00000000", --  434 - 0x1b2  :    0 - 0x0
    "00000000", --  435 - 0x1b3  :    0 - 0x0
    "00000000", --  436 - 0x1b4  :    0 - 0x0
    "00000000", --  437 - 0x1b5  :    0 - 0x0
    "00000000", --  438 - 0x1b6  :    0 - 0x0
    "00000000", --  439 - 0x1b7  :    0 - 0x0
    "00000000", --  440 - 0x1b8  :    0 - 0x0 -- Background 0x37
    "00000000", --  441 - 0x1b9  :    0 - 0x0
    "00000000", --  442 - 0x1ba  :    0 - 0x0
    "00000000", --  443 - 0x1bb  :    0 - 0x0
    "00000000", --  444 - 0x1bc  :    0 - 0x0
    "00000000", --  445 - 0x1bd  :    0 - 0x0
    "00000000", --  446 - 0x1be  :    0 - 0x0
    "00000000", --  447 - 0x1bf  :    0 - 0x0
    "00000000", --  448 - 0x1c0  :    0 - 0x0 -- Background 0x38
    "00000000", --  449 - 0x1c1  :    0 - 0x0
    "00000000", --  450 - 0x1c2  :    0 - 0x0
    "00000000", --  451 - 0x1c3  :    0 - 0x0
    "00000000", --  452 - 0x1c4  :    0 - 0x0
    "00000000", --  453 - 0x1c5  :    0 - 0x0
    "00000000", --  454 - 0x1c6  :    0 - 0x0
    "00000000", --  455 - 0x1c7  :    0 - 0x0
    "00000000", --  456 - 0x1c8  :    0 - 0x0 -- Background 0x39
    "00000000", --  457 - 0x1c9  :    0 - 0x0
    "00000000", --  458 - 0x1ca  :    0 - 0x0
    "00000000", --  459 - 0x1cb  :    0 - 0x0
    "00000000", --  460 - 0x1cc  :    0 - 0x0
    "00000000", --  461 - 0x1cd  :    0 - 0x0
    "00000000", --  462 - 0x1ce  :    0 - 0x0
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "00000000", --  464 - 0x1d0  :    0 - 0x0 -- Background 0x3a
    "00000000", --  465 - 0x1d1  :    0 - 0x0
    "00000000", --  466 - 0x1d2  :    0 - 0x0
    "00000000", --  467 - 0x1d3  :    0 - 0x0
    "00000000", --  468 - 0x1d4  :    0 - 0x0
    "00000000", --  469 - 0x1d5  :    0 - 0x0
    "00000000", --  470 - 0x1d6  :    0 - 0x0
    "00000000", --  471 - 0x1d7  :    0 - 0x0
    "00000000", --  472 - 0x1d8  :    0 - 0x0 -- Background 0x3b
    "00000000", --  473 - 0x1d9  :    0 - 0x0
    "00000000", --  474 - 0x1da  :    0 - 0x0
    "00000000", --  475 - 0x1db  :    0 - 0x0
    "00000000", --  476 - 0x1dc  :    0 - 0x0
    "00000000", --  477 - 0x1dd  :    0 - 0x0
    "00000000", --  478 - 0x1de  :    0 - 0x0
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "00000000", --  480 - 0x1e0  :    0 - 0x0 -- Background 0x3c
    "00000000", --  481 - 0x1e1  :    0 - 0x0
    "00000000", --  482 - 0x1e2  :    0 - 0x0
    "00000000", --  483 - 0x1e3  :    0 - 0x0
    "00000000", --  484 - 0x1e4  :    0 - 0x0
    "00000000", --  485 - 0x1e5  :    0 - 0x0
    "00000000", --  486 - 0x1e6  :    0 - 0x0
    "00000000", --  487 - 0x1e7  :    0 - 0x0
    "00000000", --  488 - 0x1e8  :    0 - 0x0 -- Background 0x3d
    "00000000", --  489 - 0x1e9  :    0 - 0x0
    "00000000", --  490 - 0x1ea  :    0 - 0x0
    "00000000", --  491 - 0x1eb  :    0 - 0x0
    "00000000", --  492 - 0x1ec  :    0 - 0x0
    "00000000", --  493 - 0x1ed  :    0 - 0x0
    "00000000", --  494 - 0x1ee  :    0 - 0x0
    "00000000", --  495 - 0x1ef  :    0 - 0x0
    "00000000", --  496 - 0x1f0  :    0 - 0x0 -- Background 0x3e
    "00000000", --  497 - 0x1f1  :    0 - 0x0
    "00000000", --  498 - 0x1f2  :    0 - 0x0
    "00000000", --  499 - 0x1f3  :    0 - 0x0
    "00000000", --  500 - 0x1f4  :    0 - 0x0
    "00000000", --  501 - 0x1f5  :    0 - 0x0
    "00000000", --  502 - 0x1f6  :    0 - 0x0
    "00000000", --  503 - 0x1f7  :    0 - 0x0
    "10000001", --  504 - 0x1f8  :  129 - 0x81 -- Background 0x3f
    "11111111", --  505 - 0x1f9  :  255 - 0xff
    "10000001", --  506 - 0x1fa  :  129 - 0x81
    "10000001", --  507 - 0x1fb  :  129 - 0x81
    "10000001", --  508 - 0x1fc  :  129 - 0x81
    "11111111", --  509 - 0x1fd  :  255 - 0xff
    "10000001", --  510 - 0x1fe  :  129 - 0x81
    "10000001", --  511 - 0x1ff  :  129 - 0x81
    "10000001", --  512 - 0x200  :  129 - 0x81 -- Background 0x40
    "11111111", --  513 - 0x201  :  255 - 0xff
    "10000001", --  514 - 0x202  :  129 - 0x81
    "10000001", --  515 - 0x203  :  129 - 0x81
    "10000001", --  516 - 0x204  :  129 - 0x81
    "11111111", --  517 - 0x205  :  255 - 0xff
    "10000001", --  518 - 0x206  :  129 - 0x81
    "00000000", --  519 - 0x207  :    0 - 0x0
    "10000001", --  520 - 0x208  :  129 - 0x81 -- Background 0x41
    "11111111", --  521 - 0x209  :  255 - 0xff
    "10000001", --  522 - 0x20a  :  129 - 0x81
    "10000001", --  523 - 0x20b  :  129 - 0x81
    "10000001", --  524 - 0x20c  :  129 - 0x81
    "00000000", --  525 - 0x20d  :    0 - 0x0
    "00000000", --  526 - 0x20e  :    0 - 0x0
    "00000000", --  527 - 0x20f  :    0 - 0x0
    "10000001", --  528 - 0x210  :  129 - 0x81 -- Background 0x42
    "11111111", --  529 - 0x211  :  255 - 0xff
    "10000001", --  530 - 0x212  :  129 - 0x81
    "10000001", --  531 - 0x213  :  129 - 0x81
    "00000000", --  532 - 0x214  :    0 - 0x0
    "00000000", --  533 - 0x215  :    0 - 0x0
    "00000000", --  534 - 0x216  :    0 - 0x0
    "00000000", --  535 - 0x217  :    0 - 0x0
    "10000001", --  536 - 0x218  :  129 - 0x81 -- Background 0x43
    "11111111", --  537 - 0x219  :  255 - 0xff
    "10000001", --  538 - 0x21a  :  129 - 0x81
    "00000000", --  539 - 0x21b  :    0 - 0x0
    "00000000", --  540 - 0x21c  :    0 - 0x0
    "00000000", --  541 - 0x21d  :    0 - 0x0
    "00000000", --  542 - 0x21e  :    0 - 0x0
    "00000000", --  543 - 0x21f  :    0 - 0x0
    "10000001", --  544 - 0x220  :  129 - 0x81 -- Background 0x44
    "11111111", --  545 - 0x221  :  255 - 0xff
    "00000000", --  546 - 0x222  :    0 - 0x0
    "00000000", --  547 - 0x223  :    0 - 0x0
    "00000000", --  548 - 0x224  :    0 - 0x0
    "00000000", --  549 - 0x225  :    0 - 0x0
    "00000000", --  550 - 0x226  :    0 - 0x0
    "00000000", --  551 - 0x227  :    0 - 0x0
    "10000001", --  552 - 0x228  :  129 - 0x81 -- Background 0x45
    "00000000", --  553 - 0x229  :    0 - 0x0
    "00000000", --  554 - 0x22a  :    0 - 0x0
    "00000000", --  555 - 0x22b  :    0 - 0x0
    "00000000", --  556 - 0x22c  :    0 - 0x0
    "00000000", --  557 - 0x22d  :    0 - 0x0
    "00000000", --  558 - 0x22e  :    0 - 0x0
    "00000000", --  559 - 0x22f  :    0 - 0x0
    "00000000", --  560 - 0x230  :    0 - 0x0 -- Background 0x46
    "00000000", --  561 - 0x231  :    0 - 0x0
    "00000000", --  562 - 0x232  :    0 - 0x0
    "00000000", --  563 - 0x233  :    0 - 0x0
    "00000000", --  564 - 0x234  :    0 - 0x0
    "00000000", --  565 - 0x235  :    0 - 0x0
    "00000000", --  566 - 0x236  :    0 - 0x0
    "10000001", --  567 - 0x237  :  129 - 0x81
    "00000000", --  568 - 0x238  :    0 - 0x0 -- Background 0x47
    "00000000", --  569 - 0x239  :    0 - 0x0
    "00000000", --  570 - 0x23a  :    0 - 0x0
    "00000000", --  571 - 0x23b  :    0 - 0x0
    "00000000", --  572 - 0x23c  :    0 - 0x0
    "00000000", --  573 - 0x23d  :    0 - 0x0
    "10000001", --  574 - 0x23e  :  129 - 0x81
    "10000001", --  575 - 0x23f  :  129 - 0x81
    "00000000", --  576 - 0x240  :    0 - 0x0 -- Background 0x48
    "00000000", --  577 - 0x241  :    0 - 0x0
    "00000000", --  578 - 0x242  :    0 - 0x0
    "00000000", --  579 - 0x243  :    0 - 0x0
    "00000000", --  580 - 0x244  :    0 - 0x0
    "11111111", --  581 - 0x245  :  255 - 0xff
    "10000001", --  582 - 0x246  :  129 - 0x81
    "10000001", --  583 - 0x247  :  129 - 0x81
    "00000000", --  584 - 0x248  :    0 - 0x0 -- Background 0x49
    "00000000", --  585 - 0x249  :    0 - 0x0
    "00000000", --  586 - 0x24a  :    0 - 0x0
    "00000000", --  587 - 0x24b  :    0 - 0x0
    "10000001", --  588 - 0x24c  :  129 - 0x81
    "11111111", --  589 - 0x24d  :  255 - 0xff
    "10000001", --  590 - 0x24e  :  129 - 0x81
    "10000001", --  591 - 0x24f  :  129 - 0x81
    "00000000", --  592 - 0x250  :    0 - 0x0 -- Background 0x4a
    "00000000", --  593 - 0x251  :    0 - 0x0
    "00000000", --  594 - 0x252  :    0 - 0x0
    "10000001", --  595 - 0x253  :  129 - 0x81
    "10000001", --  596 - 0x254  :  129 - 0x81
    "11111111", --  597 - 0x255  :  255 - 0xff
    "10000001", --  598 - 0x256  :  129 - 0x81
    "10000001", --  599 - 0x257  :  129 - 0x81
    "00000000", --  600 - 0x258  :    0 - 0x0 -- Background 0x4b
    "00000000", --  601 - 0x259  :    0 - 0x0
    "10000001", --  602 - 0x25a  :  129 - 0x81
    "10000001", --  603 - 0x25b  :  129 - 0x81
    "10000001", --  604 - 0x25c  :  129 - 0x81
    "11111111", --  605 - 0x25d  :  255 - 0xff
    "10000001", --  606 - 0x25e  :  129 - 0x81
    "10000001", --  607 - 0x25f  :  129 - 0x81
    "11111111", --  608 - 0x260  :  255 - 0xff -- Background 0x4c
    "01111111", --  609 - 0x261  :  127 - 0x7f
    "01111111", --  610 - 0x262  :  127 - 0x7f
    "01111111", --  611 - 0x263  :  127 - 0x7f
    "01111111", --  612 - 0x264  :  127 - 0x7f
    "01111111", --  613 - 0x265  :  127 - 0x7f
    "01111111", --  614 - 0x266  :  127 - 0x7f
    "01111111", --  615 - 0x267  :  127 - 0x7f
    "01111111", --  616 - 0x268  :  127 - 0x7f -- Background 0x4d
    "01111111", --  617 - 0x269  :  127 - 0x7f
    "01111111", --  618 - 0x26a  :  127 - 0x7f
    "01111111", --  619 - 0x26b  :  127 - 0x7f
    "01110010", --  620 - 0x26c  :  114 - 0x72
    "01111111", --  621 - 0x26d  :  127 - 0x7f
    "01111111", --  622 - 0x26e  :  127 - 0x7f
    "11111111", --  623 - 0x26f  :  255 - 0xff
    "11111111", --  624 - 0x270  :  255 - 0xff -- Background 0x4e
    "11111110", --  625 - 0x271  :  254 - 0xfe
    "11111110", --  626 - 0x272  :  254 - 0xfe
    "11111110", --  627 - 0x273  :  254 - 0xfe
    "11111110", --  628 - 0x274  :  254 - 0xfe
    "11111110", --  629 - 0x275  :  254 - 0xfe
    "11111110", --  630 - 0x276  :  254 - 0xfe
    "11111110", --  631 - 0x277  :  254 - 0xfe
    "11111110", --  632 - 0x278  :  254 - 0xfe -- Background 0x4f
    "11111110", --  633 - 0x279  :  254 - 0xfe
    "11111110", --  634 - 0x27a  :  254 - 0xfe
    "11111110", --  635 - 0x27b  :  254 - 0xfe
    "01001010", --  636 - 0x27c  :   74 - 0x4a
    "11111110", --  637 - 0x27d  :  254 - 0xfe
    "11111110", --  638 - 0x27e  :  254 - 0xfe
    "11111111", --  639 - 0x27f  :  255 - 0xff
    "00000101", --  640 - 0x280  :    5 - 0x5 -- Background 0x50
    "00001111", --  641 - 0x281  :   15 - 0xf
    "00001011", --  642 - 0x282  :   11 - 0xb
    "00011011", --  643 - 0x283  :   27 - 0x1b
    "00010011", --  644 - 0x284  :   19 - 0x13
    "00010011", --  645 - 0x285  :   19 - 0x13
    "00010011", --  646 - 0x286  :   19 - 0x13
    "00010011", --  647 - 0x287  :   19 - 0x13
    "00010011", --  648 - 0x288  :   19 - 0x13 -- Background 0x51
    "00010011", --  649 - 0x289  :   19 - 0x13
    "00010011", --  650 - 0x28a  :   19 - 0x13
    "00010011", --  651 - 0x28b  :   19 - 0x13
    "00011011", --  652 - 0x28c  :   27 - 0x1b
    "00001011", --  653 - 0x28d  :   11 - 0xb
    "00001111", --  654 - 0x28e  :   15 - 0xf
    "00000101", --  655 - 0x28f  :    5 - 0x5
    "00000101", --  656 - 0x290  :    5 - 0x5 -- Background 0x52
    "00001111", --  657 - 0x291  :   15 - 0xf
    "00001011", --  658 - 0x292  :   11 - 0xb
    "00011011", --  659 - 0x293  :   27 - 0x1b
    "00010011", --  660 - 0x294  :   19 - 0x13
    "00010011", --  661 - 0x295  :   19 - 0x13
    "00010011", --  662 - 0x296  :   19 - 0x13
    "00010011", --  663 - 0x297  :   19 - 0x13
    "00010011", --  664 - 0x298  :   19 - 0x13 -- Background 0x53
    "00010011", --  665 - 0x299  :   19 - 0x13
    "00010011", --  666 - 0x29a  :   19 - 0x13
    "00010011", --  667 - 0x29b  :   19 - 0x13
    "00011011", --  668 - 0x29c  :   27 - 0x1b
    "00001011", --  669 - 0x29d  :   11 - 0xb
    "00001111", --  670 - 0x29e  :   15 - 0xf
    "00000101", --  671 - 0x29f  :    5 - 0x5
    "10100000", --  672 - 0x2a0  :  160 - 0xa0 -- Background 0x54
    "11110001", --  673 - 0x2a1  :  241 - 0xf1
    "11010001", --  674 - 0x2a2  :  209 - 0xd1
    "11011011", --  675 - 0x2a3  :  219 - 0xdb
    "11001010", --  676 - 0x2a4  :  202 - 0xca
    "11001010", --  677 - 0x2a5  :  202 - 0xca
    "11001010", --  678 - 0x2a6  :  202 - 0xca
    "11001010", --  679 - 0x2a7  :  202 - 0xca
    "11001010", --  680 - 0x2a8  :  202 - 0xca -- Background 0x55
    "11001010", --  681 - 0x2a9  :  202 - 0xca
    "11001010", --  682 - 0x2aa  :  202 - 0xca
    "11001010", --  683 - 0x2ab  :  202 - 0xca
    "11011011", --  684 - 0x2ac  :  219 - 0xdb
    "11010001", --  685 - 0x2ad  :  209 - 0xd1
    "11110001", --  686 - 0x2ae  :  241 - 0xf1
    "10100000", --  687 - 0x2af  :  160 - 0xa0
    "10100000", --  688 - 0x2b0  :  160 - 0xa0 -- Background 0x56
    "11110001", --  689 - 0x2b1  :  241 - 0xf1
    "11010001", --  690 - 0x2b2  :  209 - 0xd1
    "11011011", --  691 - 0x2b3  :  219 - 0xdb
    "11001010", --  692 - 0x2b4  :  202 - 0xca
    "11001010", --  693 - 0x2b5  :  202 - 0xca
    "11001010", --  694 - 0x2b6  :  202 - 0xca
    "11001010", --  695 - 0x2b7  :  202 - 0xca
    "11001010", --  696 - 0x2b8  :  202 - 0xca -- Background 0x57
    "11001010", --  697 - 0x2b9  :  202 - 0xca
    "11001010", --  698 - 0x2ba  :  202 - 0xca
    "11001010", --  699 - 0x2bb  :  202 - 0xca
    "11011011", --  700 - 0x2bc  :  219 - 0xdb
    "11010001", --  701 - 0x2bd  :  209 - 0xd1
    "11110000", --  702 - 0x2be  :  240 - 0xf0
    "10100000", --  703 - 0x2bf  :  160 - 0xa0
    "10110100", --  704 - 0x2c0  :  180 - 0xb4 -- Background 0x58
    "11111110", --  705 - 0x2c1  :  254 - 0xfe
    "01111010", --  706 - 0x2c2  :  122 - 0x7a
    "01111011", --  707 - 0x2c3  :  123 - 0x7b
    "01111001", --  708 - 0x2c4  :  121 - 0x79
    "01111001", --  709 - 0x2c5  :  121 - 0x79
    "01111001", --  710 - 0x2c6  :  121 - 0x79
    "01111001", --  711 - 0x2c7  :  121 - 0x79
    "01111001", --  712 - 0x2c8  :  121 - 0x79 -- Background 0x59
    "01111001", --  713 - 0x2c9  :  121 - 0x79
    "01111001", --  714 - 0x2ca  :  121 - 0x79
    "01111001", --  715 - 0x2cb  :  121 - 0x79
    "01111011", --  716 - 0x2cc  :  123 - 0x7b
    "01111010", --  717 - 0x2cd  :  122 - 0x7a
    "11111110", --  718 - 0x2ce  :  254 - 0xfe
    "10110100", --  719 - 0x2cf  :  180 - 0xb4
    "10110100", --  720 - 0x2d0  :  180 - 0xb4 -- Background 0x5a
    "11111110", --  721 - 0x2d1  :  254 - 0xfe
    "01111010", --  722 - 0x2d2  :  122 - 0x7a
    "01111011", --  723 - 0x2d3  :  123 - 0x7b
    "01111001", --  724 - 0x2d4  :  121 - 0x79
    "01111001", --  725 - 0x2d5  :  121 - 0x79
    "01111001", --  726 - 0x2d6  :  121 - 0x79
    "01111001", --  727 - 0x2d7  :  121 - 0x79
    "01111001", --  728 - 0x2d8  :  121 - 0x79 -- Background 0x5b
    "01111001", --  729 - 0x2d9  :  121 - 0x79
    "01111001", --  730 - 0x2da  :  121 - 0x79
    "01111001", --  731 - 0x2db  :  121 - 0x79
    "01111011", --  732 - 0x2dc  :  123 - 0x7b
    "01111010", --  733 - 0x2dd  :  122 - 0x7a
    "11111110", --  734 - 0x2de  :  254 - 0xfe
    "10110100", --  735 - 0x2df  :  180 - 0xb4
    "01111111", --  736 - 0x2e0  :  127 - 0x7f -- Background 0x5c
    "10111111", --  737 - 0x2e1  :  191 - 0xbf
    "11111111", --  738 - 0x2e2  :  255 - 0xff
    "10110010", --  739 - 0x2e3  :  178 - 0xb2
    "10110001", --  740 - 0x2e4  :  177 - 0xb1
    "11111111", --  741 - 0x2e5  :  255 - 0xff
    "10111111", --  742 - 0x2e6  :  191 - 0xbf
    "01111111", --  743 - 0x2e7  :  127 - 0x7f
    "11111110", --  744 - 0x2e8  :  254 - 0xfe -- Background 0x5d
    "11111101", --  745 - 0x2e9  :  253 - 0xfd
    "11111111", --  746 - 0x2ea  :  255 - 0xff
    "11001101", --  747 - 0x2eb  :  205 - 0xcd
    "01101101", --  748 - 0x2ec  :  109 - 0x6d
    "11111111", --  749 - 0x2ed  :  255 - 0xff
    "11111101", --  750 - 0x2ee  :  253 - 0xfd
    "11111110", --  751 - 0x2ef  :  254 - 0xfe
    "11111111", --  752 - 0x2f0  :  255 - 0xff -- Background 0x5e
    "11111111", --  753 - 0x2f1  :  255 - 0xff
    "10101110", --  754 - 0x2f2  :  174 - 0xae
    "11111110", --  755 - 0x2f3  :  254 - 0xfe
    "11111111", --  756 - 0x2f4  :  255 - 0xff
    "00001111", --  757 - 0x2f5  :   15 - 0xf
    "00000111", --  758 - 0x2f6  :    7 - 0x7
    "00000011", --  759 - 0x2f7  :    3 - 0x3
    "11111111", --  760 - 0x2f8  :  255 - 0xff -- Background 0x5f
    "11111111", --  761 - 0x2f9  :  255 - 0xff
    "01110101", --  762 - 0x2fa  :  117 - 0x75
    "01111111", --  763 - 0x2fb  :  127 - 0x7f
    "11111111", --  764 - 0x2fc  :  255 - 0xff
    "11110000", --  765 - 0x2fd  :  240 - 0xf0
    "11100000", --  766 - 0x2fe  :  224 - 0xe0
    "11000000", --  767 - 0x2ff  :  192 - 0xc0
    "00000011", --  768 - 0x300  :    3 - 0x3 -- Background 0x60
    "00000111", --  769 - 0x301  :    7 - 0x7
    "00001111", --  770 - 0x302  :   15 - 0xf
    "11111111", --  771 - 0x303  :  255 - 0xff
    "11111110", --  772 - 0x304  :  254 - 0xfe
    "10101110", --  773 - 0x305  :  174 - 0xae
    "11111111", --  774 - 0x306  :  255 - 0xff
    "11111111", --  775 - 0x307  :  255 - 0xff
    "11000000", --  776 - 0x308  :  192 - 0xc0 -- Background 0x61
    "11100000", --  777 - 0x309  :  224 - 0xe0
    "11110000", --  778 - 0x30a  :  240 - 0xf0
    "11111111", --  779 - 0x30b  :  255 - 0xff
    "01111111", --  780 - 0x30c  :  127 - 0x7f
    "01110101", --  781 - 0x30d  :  117 - 0x75
    "11111111", --  782 - 0x30e  :  255 - 0xff
    "11111111", --  783 - 0x30f  :  255 - 0xff
    "11111111", --  784 - 0x310  :  255 - 0xff -- Background 0x62
    "00000000", --  785 - 0x311  :    0 - 0x0
    "11000011", --  786 - 0x312  :  195 - 0xc3
    "10000001", --  787 - 0x313  :  129 - 0x81
    "10000001", --  788 - 0x314  :  129 - 0x81
    "11000011", --  789 - 0x315  :  195 - 0xc3
    "11111111", --  790 - 0x316  :  255 - 0xff
    "00000000", --  791 - 0x317  :    0 - 0x0
    "10000001", --  792 - 0x318  :  129 - 0x81 -- Background 0x63
    "01100110", --  793 - 0x319  :  102 - 0x66
    "01111110", --  794 - 0x31a  :  126 - 0x7e
    "01111110", --  795 - 0x31b  :  126 - 0x7e
    "01111110", --  796 - 0x31c  :  126 - 0x7e
    "11111111", --  797 - 0x31d  :  255 - 0xff
    "11111111", --  798 - 0x31e  :  255 - 0xff
    "01111110", --  799 - 0x31f  :  126 - 0x7e
    "00000000", --  800 - 0x320  :    0 - 0x0 -- Background 0x64
    "00000000", --  801 - 0x321  :    0 - 0x0
    "00000000", --  802 - 0x322  :    0 - 0x0
    "00000000", --  803 - 0x323  :    0 - 0x0
    "00000000", --  804 - 0x324  :    0 - 0x0
    "00000000", --  805 - 0x325  :    0 - 0x0
    "00000000", --  806 - 0x326  :    0 - 0x0
    "00000000", --  807 - 0x327  :    0 - 0x0
    "00000000", --  808 - 0x328  :    0 - 0x0 -- Background 0x65
    "00000000", --  809 - 0x329  :    0 - 0x0
    "00000000", --  810 - 0x32a  :    0 - 0x0
    "00000000", --  811 - 0x32b  :    0 - 0x0
    "00000000", --  812 - 0x32c  :    0 - 0x0
    "00000000", --  813 - 0x32d  :    0 - 0x0
    "00000000", --  814 - 0x32e  :    0 - 0x0
    "00000000", --  815 - 0x32f  :    0 - 0x0
    "00000000", --  816 - 0x330  :    0 - 0x0 -- Background 0x66
    "00000000", --  817 - 0x331  :    0 - 0x0
    "00000000", --  818 - 0x332  :    0 - 0x0
    "00000000", --  819 - 0x333  :    0 - 0x0
    "00000000", --  820 - 0x334  :    0 - 0x0
    "00000000", --  821 - 0x335  :    0 - 0x0
    "00000000", --  822 - 0x336  :    0 - 0x0
    "00000000", --  823 - 0x337  :    0 - 0x0
    "00000000", --  824 - 0x338  :    0 - 0x0 -- Background 0x67
    "00000000", --  825 - 0x339  :    0 - 0x0
    "00000000", --  826 - 0x33a  :    0 - 0x0
    "00000000", --  827 - 0x33b  :    0 - 0x0
    "00000000", --  828 - 0x33c  :    0 - 0x0
    "00000000", --  829 - 0x33d  :    0 - 0x0
    "00000000", --  830 - 0x33e  :    0 - 0x0
    "00000000", --  831 - 0x33f  :    0 - 0x0
    "00000011", --  832 - 0x340  :    3 - 0x3 -- Background 0x68
    "00000001", --  833 - 0x341  :    1 - 0x1
    "00000000", --  834 - 0x342  :    0 - 0x0
    "00000000", --  835 - 0x343  :    0 - 0x0
    "00000000", --  836 - 0x344  :    0 - 0x0
    "00000000", --  837 - 0x345  :    0 - 0x0
    "00000000", --  838 - 0x346  :    0 - 0x0
    "00000000", --  839 - 0x347  :    0 - 0x0
    "11111111", --  840 - 0x348  :  255 - 0xff -- Background 0x69
    "11111111", --  841 - 0x349  :  255 - 0xff
    "11111111", --  842 - 0x34a  :  255 - 0xff
    "11111111", --  843 - 0x34b  :  255 - 0xff
    "11111111", --  844 - 0x34c  :  255 - 0xff
    "11111111", --  845 - 0x34d  :  255 - 0xff
    "11111111", --  846 - 0x34e  :  255 - 0xff
    "11111111", --  847 - 0x34f  :  255 - 0xff
    "11000000", --  848 - 0x350  :  192 - 0xc0 -- Background 0x6a
    "10000000", --  849 - 0x351  :  128 - 0x80
    "00000000", --  850 - 0x352  :    0 - 0x0
    "00000000", --  851 - 0x353  :    0 - 0x0
    "00000000", --  852 - 0x354  :    0 - 0x0
    "00000000", --  853 - 0x355  :    0 - 0x0
    "00000000", --  854 - 0x356  :    0 - 0x0
    "00000000", --  855 - 0x357  :    0 - 0x0
    "11111111", --  856 - 0x358  :  255 - 0xff -- Background 0x6b
    "11111111", --  857 - 0x359  :  255 - 0xff
    "11111111", --  858 - 0x35a  :  255 - 0xff
    "11111111", --  859 - 0x35b  :  255 - 0xff
    "11111111", --  860 - 0x35c  :  255 - 0xff
    "11111111", --  861 - 0x35d  :  255 - 0xff
    "11111111", --  862 - 0x35e  :  255 - 0xff
    "11111111", --  863 - 0x35f  :  255 - 0xff
    "11111111", --  864 - 0x360  :  255 - 0xff -- Background 0x6c
    "11111111", --  865 - 0x361  :  255 - 0xff
    "11111111", --  866 - 0x362  :  255 - 0xff
    "00011111", --  867 - 0x363  :   31 - 0x1f
    "00011111", --  868 - 0x364  :   31 - 0x1f
    "00111111", --  869 - 0x365  :   63 - 0x3f
    "01111111", --  870 - 0x366  :  127 - 0x7f
    "11111111", --  871 - 0x367  :  255 - 0xff
    "11111111", --  872 - 0x368  :  255 - 0xff -- Background 0x6d
    "11111111", --  873 - 0x369  :  255 - 0xff
    "11111111", --  874 - 0x36a  :  255 - 0xff
    "11111000", --  875 - 0x36b  :  248 - 0xf8
    "11111000", --  876 - 0x36c  :  248 - 0xf8
    "11111100", --  877 - 0x36d  :  252 - 0xfc
    "11111110", --  878 - 0x36e  :  254 - 0xfe
    "11111111", --  879 - 0x36f  :  255 - 0xff
    "00000000", --  880 - 0x370  :    0 - 0x0 -- Background 0x6e
    "00000000", --  881 - 0x371  :    0 - 0x0
    "00000000", --  882 - 0x372  :    0 - 0x0
    "00000000", --  883 - 0x373  :    0 - 0x0
    "00000000", --  884 - 0x374  :    0 - 0x0
    "00111100", --  885 - 0x375  :   60 - 0x3c
    "01000010", --  886 - 0x376  :   66 - 0x42
    "10000001", --  887 - 0x377  :  129 - 0x81
    "10000001", --  888 - 0x378  :  129 - 0x81 -- Background 0x6f
    "10111101", --  889 - 0x379  :  189 - 0xbd
    "01111110", --  890 - 0x37a  :  126 - 0x7e
    "10100101", --  891 - 0x37b  :  165 - 0xa5
    "11011011", --  892 - 0x37c  :  219 - 0xdb
    "11100111", --  893 - 0x37d  :  231 - 0xe7
    "11111111", --  894 - 0x37e  :  255 - 0xff
    "11111111", --  895 - 0x37f  :  255 - 0xff
    "00000000", --  896 - 0x380  :    0 - 0x0 -- Background 0x70
    "00000101", --  897 - 0x381  :    5 - 0x5
    "00011001", --  898 - 0x382  :   25 - 0x19
    "00110011", --  899 - 0x383  :   51 - 0x33
    "01100011", --  900 - 0x384  :   99 - 0x63
    "11000111", --  901 - 0x385  :  199 - 0xc7
    "11000111", --  902 - 0x386  :  199 - 0xc7
    "11000100", --  903 - 0x387  :  196 - 0xc4
    "10000000", --  904 - 0x388  :  128 - 0x80 -- Background 0x71
    "00000000", --  905 - 0x389  :    0 - 0x0
    "00000000", --  906 - 0x38a  :    0 - 0x0
    "00000001", --  907 - 0x38b  :    1 - 0x1
    "00000001", --  908 - 0x38c  :    1 - 0x1
    "00000001", --  909 - 0x38d  :    1 - 0x1
    "00000000", --  910 - 0x38e  :    0 - 0x0
    "00000000", --  911 - 0x38f  :    0 - 0x0
    "00000000", --  912 - 0x390  :    0 - 0x0 -- Background 0x72
    "10100000", --  913 - 0x391  :  160 - 0xa0
    "10011000", --  914 - 0x392  :  152 - 0x98
    "11001100", --  915 - 0x393  :  204 - 0xcc
    "11000110", --  916 - 0x394  :  198 - 0xc6
    "11100011", --  917 - 0x395  :  227 - 0xe3
    "11100011", --  918 - 0x396  :  227 - 0xe3
    "00100011", --  919 - 0x397  :   35 - 0x23
    "00000001", --  920 - 0x398  :    1 - 0x1 -- Background 0x73
    "00000000", --  921 - 0x399  :    0 - 0x0
    "00000000", --  922 - 0x39a  :    0 - 0x0
    "00000000", --  923 - 0x39b  :    0 - 0x0
    "00000000", --  924 - 0x39c  :    0 - 0x0
    "01000000", --  925 - 0x39d  :   64 - 0x40
    "10000000", --  926 - 0x39e  :  128 - 0x80
    "00000000", --  927 - 0x39f  :    0 - 0x0
    "00000001", --  928 - 0x3a0  :    1 - 0x1 -- Background 0x74
    "00000001", --  929 - 0x3a1  :    1 - 0x1
    "00000001", --  930 - 0x3a2  :    1 - 0x1
    "00000001", --  931 - 0x3a3  :    1 - 0x1
    "00000001", --  932 - 0x3a4  :    1 - 0x1
    "00000001", --  933 - 0x3a5  :    1 - 0x1
    "00000001", --  934 - 0x3a6  :    1 - 0x1
    "00000001", --  935 - 0x3a7  :    1 - 0x1
    "10000000", --  936 - 0x3a8  :  128 - 0x80 -- Background 0x75
    "10000000", --  937 - 0x3a9  :  128 - 0x80
    "10000000", --  938 - 0x3aa  :  128 - 0x80
    "10000000", --  939 - 0x3ab  :  128 - 0x80
    "10000000", --  940 - 0x3ac  :  128 - 0x80
    "10000000", --  941 - 0x3ad  :  128 - 0x80
    "10000000", --  942 - 0x3ae  :  128 - 0x80
    "10000000", --  943 - 0x3af  :  128 - 0x80
    "00000001", --  944 - 0x3b0  :    1 - 0x1 -- Background 0x76
    "00000011", --  945 - 0x3b1  :    3 - 0x3
    "00000011", --  946 - 0x3b2  :    3 - 0x3
    "00000111", --  947 - 0x3b3  :    7 - 0x7
    "00000100", --  948 - 0x3b4  :    4 - 0x4
    "00011100", --  949 - 0x3b5  :   28 - 0x1c
    "00111111", --  950 - 0x3b6  :   63 - 0x3f
    "01111111", --  951 - 0x3b7  :  127 - 0x7f
    "01111111", --  952 - 0x3b8  :  127 - 0x7f -- Background 0x77
    "11111111", --  953 - 0x3b9  :  255 - 0xff
    "11111111", --  954 - 0x3ba  :  255 - 0xff
    "01111111", --  955 - 0x3bb  :  127 - 0x7f
    "01111111", --  956 - 0x3bc  :  127 - 0x7f
    "00011111", --  957 - 0x3bd  :   31 - 0x1f
    "00000011", --  958 - 0x3be  :    3 - 0x3
    "00000000", --  959 - 0x3bf  :    0 - 0x0
    "00000000", --  960 - 0x3c0  :    0 - 0x0 -- Background 0x78
    "00000000", --  961 - 0x3c1  :    0 - 0x0
    "00000001", --  962 - 0x3c2  :    1 - 0x1
    "00000001", --  963 - 0x3c3  :    1 - 0x1
    "00000011", --  964 - 0x3c4  :    3 - 0x3
    "00000111", --  965 - 0x3c5  :    7 - 0x7
    "00000111", --  966 - 0x3c6  :    7 - 0x7
    "00001111", --  967 - 0x3c7  :   15 - 0xf
    "11111111", --  968 - 0x3c8  :  255 - 0xff -- Background 0x79
    "11111111", --  969 - 0x3c9  :  255 - 0xff
    "00111111", --  970 - 0x3ca  :   63 - 0x3f
    "00111111", --  971 - 0x3cb  :   63 - 0x3f
    "01111111", --  972 - 0x3cc  :  127 - 0x7f
    "11111110", --  973 - 0x3cd  :  254 - 0xfe
    "11111100", --  974 - 0x3ce  :  252 - 0xfc
    "00110000", --  975 - 0x3cf  :   48 - 0x30
    "11111000", --  976 - 0x3d0  :  248 - 0xf8 -- Background 0x7a
    "11111110", --  977 - 0x3d1  :  254 - 0xfe
    "11111111", --  978 - 0x3d2  :  255 - 0xff
    "11111111", --  979 - 0x3d3  :  255 - 0xff
    "11111111", --  980 - 0x3d4  :  255 - 0xff
    "11111111", --  981 - 0x3d5  :  255 - 0xff
    "11111111", --  982 - 0x3d6  :  255 - 0xff
    "11111111", --  983 - 0x3d7  :  255 - 0xff
    "11111111", --  984 - 0x3d8  :  255 - 0xff -- Background 0x7b
    "11111111", --  985 - 0x3d9  :  255 - 0xff
    "11111111", --  986 - 0x3da  :  255 - 0xff
    "11111111", --  987 - 0x3db  :  255 - 0xff
    "11111111", --  988 - 0x3dc  :  255 - 0xff
    "11111111", --  989 - 0x3dd  :  255 - 0xff
    "11111111", --  990 - 0x3de  :  255 - 0xff
    "01111111", --  991 - 0x3df  :  127 - 0x7f
    "11111111", --  992 - 0x3e0  :  255 - 0xff -- Background 0x7c
    "11111111", --  993 - 0x3e1  :  255 - 0xff
    "11111111", --  994 - 0x3e2  :  255 - 0xff
    "11111111", --  995 - 0x3e3  :  255 - 0xff
    "11111111", --  996 - 0x3e4  :  255 - 0xff
    "11111111", --  997 - 0x3e5  :  255 - 0xff
    "11111111", --  998 - 0x3e6  :  255 - 0xff
    "11111111", --  999 - 0x3e7  :  255 - 0xff
    "11101111", -- 1000 - 0x3e8  :  239 - 0xef -- Background 0x7d
    "11001111", -- 1001 - 0x3e9  :  207 - 0xcf
    "10011111", -- 1002 - 0x3ea  :  159 - 0x9f
    "00011111", -- 1003 - 0x3eb  :   31 - 0x1f
    "00001111", -- 1004 - 0x3ec  :   15 - 0xf
    "01111111", -- 1005 - 0x3ed  :  127 - 0x7f
    "11111111", -- 1006 - 0x3ee  :  255 - 0xff
    "11111111", -- 1007 - 0x3ef  :  255 - 0xff
    "00000000", -- 1008 - 0x3f0  :    0 - 0x0 -- Background 0x7e
    "00000000", -- 1009 - 0x3f1  :    0 - 0x0
    "00000000", -- 1010 - 0x3f2  :    0 - 0x0
    "11110000", -- 1011 - 0x3f3  :  240 - 0xf0
    "11111110", -- 1012 - 0x3f4  :  254 - 0xfe
    "11111111", -- 1013 - 0x3f5  :  255 - 0xff
    "11111111", -- 1014 - 0x3f6  :  255 - 0xff
    "11111111", -- 1015 - 0x3f7  :  255 - 0xff
    "11111111", -- 1016 - 0x3f8  :  255 - 0xff -- Background 0x7f
    "11111111", -- 1017 - 0x3f9  :  255 - 0xff
    "11111111", -- 1018 - 0x3fa  :  255 - 0xff
    "11111111", -- 1019 - 0x3fb  :  255 - 0xff
    "11111111", -- 1020 - 0x3fc  :  255 - 0xff
    "11111111", -- 1021 - 0x3fd  :  255 - 0xff
    "11111111", -- 1022 - 0x3fe  :  255 - 0xff
    "11111111", -- 1023 - 0x3ff  :  255 - 0xff
    "11111111", -- 1024 - 0x400  :  255 - 0xff -- Background 0x80
    "11111111", -- 1025 - 0x401  :  255 - 0xff
    "11111111", -- 1026 - 0x402  :  255 - 0xff
    "11111111", -- 1027 - 0x403  :  255 - 0xff
    "11111111", -- 1028 - 0x404  :  255 - 0xff
    "11111111", -- 1029 - 0x405  :  255 - 0xff
    "11111111", -- 1030 - 0x406  :  255 - 0xff
    "11111111", -- 1031 - 0x407  :  255 - 0xff
    "11111111", -- 1032 - 0x408  :  255 - 0xff -- Background 0x81
    "11111111", -- 1033 - 0x409  :  255 - 0xff
    "11111111", -- 1034 - 0x40a  :  255 - 0xff
    "11110000", -- 1035 - 0x40b  :  240 - 0xf0
    "11110000", -- 1036 - 0x40c  :  240 - 0xf0
    "11111000", -- 1037 - 0x40d  :  248 - 0xf8
    "11111000", -- 1038 - 0x40e  :  248 - 0xf8
    "11111000", -- 1039 - 0x40f  :  248 - 0xf8
    "00000000", -- 1040 - 0x410  :    0 - 0x0 -- Background 0x82
    "00000000", -- 1041 - 0x411  :    0 - 0x0
    "00000000", -- 1042 - 0x412  :    0 - 0x0
    "00000000", -- 1043 - 0x413  :    0 - 0x0
    "00000000", -- 1044 - 0x414  :    0 - 0x0
    "10000000", -- 1045 - 0x415  :  128 - 0x80
    "11000000", -- 1046 - 0x416  :  192 - 0xc0
    "11100000", -- 1047 - 0x417  :  224 - 0xe0
    "11110000", -- 1048 - 0x418  :  240 - 0xf0 -- Background 0x83
    "11110000", -- 1049 - 0x419  :  240 - 0xf0
    "11111000", -- 1050 - 0x41a  :  248 - 0xf8
    "11111000", -- 1051 - 0x41b  :  248 - 0xf8
    "11111000", -- 1052 - 0x41c  :  248 - 0xf8
    "11111100", -- 1053 - 0x41d  :  252 - 0xfc
    "11111100", -- 1054 - 0x41e  :  252 - 0xfc
    "11111110", -- 1055 - 0x41f  :  254 - 0xfe
    "11111111", -- 1056 - 0x420  :  255 - 0xff -- Background 0x84
    "11111111", -- 1057 - 0x421  :  255 - 0xff
    "11111111", -- 1058 - 0x422  :  255 - 0xff
    "11111111", -- 1059 - 0x423  :  255 - 0xff
    "11111111", -- 1060 - 0x424  :  255 - 0xff
    "11111111", -- 1061 - 0x425  :  255 - 0xff
    "11111111", -- 1062 - 0x426  :  255 - 0xff
    "11111111", -- 1063 - 0x427  :  255 - 0xff
    "11111111", -- 1064 - 0x428  :  255 - 0xff -- Background 0x85
    "11111111", -- 1065 - 0x429  :  255 - 0xff
    "11111111", -- 1066 - 0x42a  :  255 - 0xff
    "00001111", -- 1067 - 0x42b  :   15 - 0xf
    "00000111", -- 1068 - 0x42c  :    7 - 0x7
    "00000000", -- 1069 - 0x42d  :    0 - 0x0
    "00000000", -- 1070 - 0x42e  :    0 - 0x0
    "00000000", -- 1071 - 0x42f  :    0 - 0x0
    "00000000", -- 1072 - 0x430  :    0 - 0x0 -- Background 0x86
    "10000000", -- 1073 - 0x431  :  128 - 0x80
    "11000000", -- 1074 - 0x432  :  192 - 0xc0
    "11100000", -- 1075 - 0x433  :  224 - 0xe0
    "11110000", -- 1076 - 0x434  :  240 - 0xf0
    "11110000", -- 1077 - 0x435  :  240 - 0xf0
    "11110000", -- 1078 - 0x436  :  240 - 0xf0
    "11111100", -- 1079 - 0x437  :  252 - 0xfc
    "11111111", -- 1080 - 0x438  :  255 - 0xff -- Background 0x87
    "11111111", -- 1081 - 0x439  :  255 - 0xff
    "11111111", -- 1082 - 0x43a  :  255 - 0xff
    "11111111", -- 1083 - 0x43b  :  255 - 0xff
    "11111111", -- 1084 - 0x43c  :  255 - 0xff
    "00001111", -- 1085 - 0x43d  :   15 - 0xf
    "00011111", -- 1086 - 0x43e  :   31 - 0x1f
    "00111111", -- 1087 - 0x43f  :   63 - 0x3f
    "11000000", -- 1088 - 0x440  :  192 - 0xc0 -- Background 0x88
    "11100000", -- 1089 - 0x441  :  224 - 0xe0
    "11100000", -- 1090 - 0x442  :  224 - 0xe0
    "11100000", -- 1091 - 0x443  :  224 - 0xe0
    "11100000", -- 1092 - 0x444  :  224 - 0xe0
    "11000000", -- 1093 - 0x445  :  192 - 0xc0
    "11000000", -- 1094 - 0x446  :  192 - 0xc0
    "10000000", -- 1095 - 0x447  :  128 - 0x80
    "00000011", -- 1096 - 0x448  :    3 - 0x3 -- Background 0x89
    "00000111", -- 1097 - 0x449  :    7 - 0x7
    "00000111", -- 1098 - 0x44a  :    7 - 0x7
    "00000111", -- 1099 - 0x44b  :    7 - 0x7
    "00000111", -- 1100 - 0x44c  :    7 - 0x7
    "00000011", -- 1101 - 0x44d  :    3 - 0x3
    "00000011", -- 1102 - 0x44e  :    3 - 0x3
    "00000001", -- 1103 - 0x44f  :    1 - 0x1
    "00000000", -- 1104 - 0x450  :    0 - 0x0 -- Background 0x8a
    "00000001", -- 1105 - 0x451  :    1 - 0x1
    "00000011", -- 1106 - 0x452  :    3 - 0x3
    "00000111", -- 1107 - 0x453  :    7 - 0x7
    "00001111", -- 1108 - 0x454  :   15 - 0xf
    "00001111", -- 1109 - 0x455  :   15 - 0xf
    "00001111", -- 1110 - 0x456  :   15 - 0xf
    "00111111", -- 1111 - 0x457  :   63 - 0x3f
    "11111111", -- 1112 - 0x458  :  255 - 0xff -- Background 0x8b
    "11111111", -- 1113 - 0x459  :  255 - 0xff
    "11111111", -- 1114 - 0x45a  :  255 - 0xff
    "11111111", -- 1115 - 0x45b  :  255 - 0xff
    "11111111", -- 1116 - 0x45c  :  255 - 0xff
    "11110000", -- 1117 - 0x45d  :  240 - 0xf0
    "11111000", -- 1118 - 0x45e  :  248 - 0xf8
    "11111100", -- 1119 - 0x45f  :  252 - 0xfc
    "00000000", -- 1120 - 0x460  :    0 - 0x0 -- Background 0x8c
    "00000000", -- 1121 - 0x461  :    0 - 0x0
    "00000000", -- 1122 - 0x462  :    0 - 0x0
    "00000000", -- 1123 - 0x463  :    0 - 0x0
    "00000000", -- 1124 - 0x464  :    0 - 0x0
    "00000001", -- 1125 - 0x465  :    1 - 0x1
    "00000011", -- 1126 - 0x466  :    3 - 0x3
    "00000111", -- 1127 - 0x467  :    7 - 0x7
    "00001111", -- 1128 - 0x468  :   15 - 0xf -- Background 0x8d
    "00001111", -- 1129 - 0x469  :   15 - 0xf
    "00011111", -- 1130 - 0x46a  :   31 - 0x1f
    "00011111", -- 1131 - 0x46b  :   31 - 0x1f
    "00011111", -- 1132 - 0x46c  :   31 - 0x1f
    "00111111", -- 1133 - 0x46d  :   63 - 0x3f
    "00111111", -- 1134 - 0x46e  :   63 - 0x3f
    "01111111", -- 1135 - 0x46f  :  127 - 0x7f
    "11111111", -- 1136 - 0x470  :  255 - 0xff -- Background 0x8e
    "11111111", -- 1137 - 0x471  :  255 - 0xff
    "11111111", -- 1138 - 0x472  :  255 - 0xff
    "11111111", -- 1139 - 0x473  :  255 - 0xff
    "11111111", -- 1140 - 0x474  :  255 - 0xff
    "11111111", -- 1141 - 0x475  :  255 - 0xff
    "11111111", -- 1142 - 0x476  :  255 - 0xff
    "11111111", -- 1143 - 0x477  :  255 - 0xff
    "11111111", -- 1144 - 0x478  :  255 - 0xff -- Background 0x8f
    "11111111", -- 1145 - 0x479  :  255 - 0xff
    "11111111", -- 1146 - 0x47a  :  255 - 0xff
    "11110000", -- 1147 - 0x47b  :  240 - 0xf0
    "11100000", -- 1148 - 0x47c  :  224 - 0xe0
    "00000000", -- 1149 - 0x47d  :    0 - 0x0
    "00000000", -- 1150 - 0x47e  :    0 - 0x0
    "00000000", -- 1151 - 0x47f  :    0 - 0x0
    "00000000", -- 1152 - 0x480  :    0 - 0x0 -- Background 0x90
    "00000000", -- 1153 - 0x481  :    0 - 0x0
    "00000000", -- 1154 - 0x482  :    0 - 0x0
    "00001111", -- 1155 - 0x483  :   15 - 0xf
    "01111111", -- 1156 - 0x484  :  127 - 0x7f
    "11111111", -- 1157 - 0x485  :  255 - 0xff
    "11111111", -- 1158 - 0x486  :  255 - 0xff
    "11111111", -- 1159 - 0x487  :  255 - 0xff
    "11111111", -- 1160 - 0x488  :  255 - 0xff -- Background 0x91
    "11111111", -- 1161 - 0x489  :  255 - 0xff
    "11111111", -- 1162 - 0x48a  :  255 - 0xff
    "11111111", -- 1163 - 0x48b  :  255 - 0xff
    "11111111", -- 1164 - 0x48c  :  255 - 0xff
    "11111111", -- 1165 - 0x48d  :  255 - 0xff
    "11111111", -- 1166 - 0x48e  :  255 - 0xff
    "11111111", -- 1167 - 0x48f  :  255 - 0xff
    "11111111", -- 1168 - 0x490  :  255 - 0xff -- Background 0x92
    "11111111", -- 1169 - 0x491  :  255 - 0xff
    "11111111", -- 1170 - 0x492  :  255 - 0xff
    "11111111", -- 1171 - 0x493  :  255 - 0xff
    "11111111", -- 1172 - 0x494  :  255 - 0xff
    "11111111", -- 1173 - 0x495  :  255 - 0xff
    "11111111", -- 1174 - 0x496  :  255 - 0xff
    "11111111", -- 1175 - 0x497  :  255 - 0xff
    "11111111", -- 1176 - 0x498  :  255 - 0xff -- Background 0x93
    "11111111", -- 1177 - 0x499  :  255 - 0xff
    "11111111", -- 1178 - 0x49a  :  255 - 0xff
    "00001111", -- 1179 - 0x49b  :   15 - 0xf
    "00001111", -- 1180 - 0x49c  :   15 - 0xf
    "00011111", -- 1181 - 0x49d  :   31 - 0x1f
    "00011111", -- 1182 - 0x49e  :   31 - 0x1f
    "00011111", -- 1183 - 0x49f  :   31 - 0x1f
    "00011111", -- 1184 - 0x4a0  :   31 - 0x1f -- Background 0x94
    "01111111", -- 1185 - 0x4a1  :  127 - 0x7f
    "11111111", -- 1186 - 0x4a2  :  255 - 0xff
    "11111111", -- 1187 - 0x4a3  :  255 - 0xff
    "11111111", -- 1188 - 0x4a4  :  255 - 0xff
    "11111111", -- 1189 - 0x4a5  :  255 - 0xff
    "11111111", -- 1190 - 0x4a6  :  255 - 0xff
    "11111111", -- 1191 - 0x4a7  :  255 - 0xff
    "11111111", -- 1192 - 0x4a8  :  255 - 0xff -- Background 0x95
    "11111111", -- 1193 - 0x4a9  :  255 - 0xff
    "11111111", -- 1194 - 0x4aa  :  255 - 0xff
    "11111111", -- 1195 - 0x4ab  :  255 - 0xff
    "11111111", -- 1196 - 0x4ac  :  255 - 0xff
    "11111111", -- 1197 - 0x4ad  :  255 - 0xff
    "11111111", -- 1198 - 0x4ae  :  255 - 0xff
    "11111110", -- 1199 - 0x4af  :  254 - 0xfe
    "11111111", -- 1200 - 0x4b0  :  255 - 0xff -- Background 0x96
    "11111111", -- 1201 - 0x4b1  :  255 - 0xff
    "11111111", -- 1202 - 0x4b2  :  255 - 0xff
    "11111111", -- 1203 - 0x4b3  :  255 - 0xff
    "11111111", -- 1204 - 0x4b4  :  255 - 0xff
    "11111111", -- 1205 - 0x4b5  :  255 - 0xff
    "11111111", -- 1206 - 0x4b6  :  255 - 0xff
    "11111111", -- 1207 - 0x4b7  :  255 - 0xff
    "11110111", -- 1208 - 0x4b8  :  247 - 0xf7 -- Background 0x97
    "11110011", -- 1209 - 0x4b9  :  243 - 0xf3
    "11111001", -- 1210 - 0x4ba  :  249 - 0xf9
    "11111000", -- 1211 - 0x4bb  :  248 - 0xf8
    "11110000", -- 1212 - 0x4bc  :  240 - 0xf0
    "11111110", -- 1213 - 0x4bd  :  254 - 0xfe
    "11111111", -- 1214 - 0x4be  :  255 - 0xff
    "11111111", -- 1215 - 0x4bf  :  255 - 0xff
    "10000000", -- 1216 - 0x4c0  :  128 - 0x80 -- Background 0x98
    "11000000", -- 1217 - 0x4c1  :  192 - 0xc0
    "11000000", -- 1218 - 0x4c2  :  192 - 0xc0
    "11100000", -- 1219 - 0x4c3  :  224 - 0xe0
    "00100000", -- 1220 - 0x4c4  :   32 - 0x20
    "00111000", -- 1221 - 0x4c5  :   56 - 0x38
    "11111100", -- 1222 - 0x4c6  :  252 - 0xfc
    "11111110", -- 1223 - 0x4c7  :  254 - 0xfe
    "11111110", -- 1224 - 0x4c8  :  254 - 0xfe -- Background 0x99
    "11111111", -- 1225 - 0x4c9  :  255 - 0xff
    "11111111", -- 1226 - 0x4ca  :  255 - 0xff
    "11111110", -- 1227 - 0x4cb  :  254 - 0xfe
    "11111100", -- 1228 - 0x4cc  :  252 - 0xfc
    "11111000", -- 1229 - 0x4cd  :  248 - 0xf8
    "11000000", -- 1230 - 0x4ce  :  192 - 0xc0
    "00000000", -- 1231 - 0x4cf  :    0 - 0x0
    "00000000", -- 1232 - 0x4d0  :    0 - 0x0 -- Background 0x9a
    "00000000", -- 1233 - 0x4d1  :    0 - 0x0
    "10000000", -- 1234 - 0x4d2  :  128 - 0x80
    "10000000", -- 1235 - 0x4d3  :  128 - 0x80
    "11000000", -- 1236 - 0x4d4  :  192 - 0xc0
    "11100000", -- 1237 - 0x4d5  :  224 - 0xe0
    "11100000", -- 1238 - 0x4d6  :  224 - 0xe0
    "11110000", -- 1239 - 0x4d7  :  240 - 0xf0
    "11111111", -- 1240 - 0x4d8  :  255 - 0xff -- Background 0x9b
    "11111111", -- 1241 - 0x4d9  :  255 - 0xff
    "11111100", -- 1242 - 0x4da  :  252 - 0xfc
    "11111100", -- 1243 - 0x4db  :  252 - 0xfc
    "11111110", -- 1244 - 0x4dc  :  254 - 0xfe
    "01111110", -- 1245 - 0x4dd  :  126 - 0x7e
    "00111111", -- 1246 - 0x4de  :   63 - 0x3f
    "00001100", -- 1247 - 0x4df  :   12 - 0xc
    "00000000", -- 1248 - 0x4e0  :    0 - 0x0 -- Background 0x9c
    "00000001", -- 1249 - 0x4e1  :    1 - 0x1
    "00000011", -- 1250 - 0x4e2  :    3 - 0x3
    "00000111", -- 1251 - 0x4e3  :    7 - 0x7
    "00000111", -- 1252 - 0x4e4  :    7 - 0x7
    "00000111", -- 1253 - 0x4e5  :    7 - 0x7
    "00001111", -- 1254 - 0x4e6  :   15 - 0xf
    "00001111", -- 1255 - 0x4e7  :   15 - 0xf
    "00001111", -- 1256 - 0x4e8  :   15 - 0xf -- Background 0x9d
    "00001111", -- 1257 - 0x4e9  :   15 - 0xf
    "00000111", -- 1258 - 0x4ea  :    7 - 0x7
    "00000111", -- 1259 - 0x4eb  :    7 - 0x7
    "00000111", -- 1260 - 0x4ec  :    7 - 0x7
    "00000011", -- 1261 - 0x4ed  :    3 - 0x3
    "00000011", -- 1262 - 0x4ee  :    3 - 0x3
    "00000001", -- 1263 - 0x4ef  :    1 - 0x1
    "00000001", -- 1264 - 0x4f0  :    1 - 0x1 -- Background 0x9e
    "00000001", -- 1265 - 0x4f1  :    1 - 0x1
    "00000001", -- 1266 - 0x4f2  :    1 - 0x1
    "00000000", -- 1267 - 0x4f3  :    0 - 0x0
    "00000000", -- 1268 - 0x4f4  :    0 - 0x0
    "00000011", -- 1269 - 0x4f5  :    3 - 0x3
    "00000111", -- 1270 - 0x4f6  :    7 - 0x7
    "00001111", -- 1271 - 0x4f7  :   15 - 0xf
    "00000000", -- 1272 - 0x4f8  :    0 - 0x0 -- Background 0x9f
    "00000000", -- 1273 - 0x4f9  :    0 - 0x0
    "00000000", -- 1274 - 0x4fa  :    0 - 0x0
    "00000000", -- 1275 - 0x4fb  :    0 - 0x0
    "00000001", -- 1276 - 0x4fc  :    1 - 0x1
    "00000011", -- 1277 - 0x4fd  :    3 - 0x3
    "00111111", -- 1278 - 0x4fe  :   63 - 0x3f
    "01111111", -- 1279 - 0x4ff  :  127 - 0x7f
    "11111111", -- 1280 - 0x500  :  255 - 0xff -- Background 0xa0
    "11111111", -- 1281 - 0x501  :  255 - 0xff
    "11111111", -- 1282 - 0x502  :  255 - 0xff
    "11111111", -- 1283 - 0x503  :  255 - 0xff
    "11111111", -- 1284 - 0x504  :  255 - 0xff
    "11111111", -- 1285 - 0x505  :  255 - 0xff
    "11111101", -- 1286 - 0x506  :  253 - 0xfd
    "11111001", -- 1287 - 0x507  :  249 - 0xf9
    "11110011", -- 1288 - 0x508  :  243 - 0xf3 -- Background 0xa1
    "11111111", -- 1289 - 0x509  :  255 - 0xff
    "11111111", -- 1290 - 0x50a  :  255 - 0xff
    "11111111", -- 1291 - 0x50b  :  255 - 0xff
    "11111111", -- 1292 - 0x50c  :  255 - 0xff
    "11111111", -- 1293 - 0x50d  :  255 - 0xff
    "11111111", -- 1294 - 0x50e  :  255 - 0xff
    "11111111", -- 1295 - 0x50f  :  255 - 0xff
    "11111111", -- 1296 - 0x510  :  255 - 0xff -- Background 0xa2
    "11111111", -- 1297 - 0x511  :  255 - 0xff
    "11111111", -- 1298 - 0x512  :  255 - 0xff
    "11111111", -- 1299 - 0x513  :  255 - 0xff
    "11111111", -- 1300 - 0x514  :  255 - 0xff
    "11111111", -- 1301 - 0x515  :  255 - 0xff
    "11111111", -- 1302 - 0x516  :  255 - 0xff
    "11111111", -- 1303 - 0x517  :  255 - 0xff
    "00000111", -- 1304 - 0x518  :    7 - 0x7 -- Background 0xa3
    "00001111", -- 1305 - 0x519  :   15 - 0xf
    "00011111", -- 1306 - 0x51a  :   31 - 0x1f
    "00111111", -- 1307 - 0x51b  :   63 - 0x3f
    "11111100", -- 1308 - 0x51c  :  252 - 0xfc
    "11111100", -- 1309 - 0x51d  :  252 - 0xfc
    "11111111", -- 1310 - 0x51e  :  255 - 0xff
    "11111111", -- 1311 - 0x51f  :  255 - 0xff
    "11111111", -- 1312 - 0x520  :  255 - 0xff -- Background 0xa4
    "11111111", -- 1313 - 0x521  :  255 - 0xff
    "11111111", -- 1314 - 0x522  :  255 - 0xff
    "11111111", -- 1315 - 0x523  :  255 - 0xff
    "11111111", -- 1316 - 0x524  :  255 - 0xff
    "11111111", -- 1317 - 0x525  :  255 - 0xff
    "11111111", -- 1318 - 0x526  :  255 - 0xff
    "11111111", -- 1319 - 0x527  :  255 - 0xff
    "11111111", -- 1320 - 0x528  :  255 - 0xff -- Background 0xa5
    "11111111", -- 1321 - 0x529  :  255 - 0xff
    "11111111", -- 1322 - 0x52a  :  255 - 0xff
    "11111111", -- 1323 - 0x52b  :  255 - 0xff
    "11111111", -- 1324 - 0x52c  :  255 - 0xff
    "11111111", -- 1325 - 0x52d  :  255 - 0xff
    "11111111", -- 1326 - 0x52e  :  255 - 0xff
    "11111111", -- 1327 - 0x52f  :  255 - 0xff
    "11111111", -- 1328 - 0x530  :  255 - 0xff -- Background 0xa6
    "11111111", -- 1329 - 0x531  :  255 - 0xff
    "11110000", -- 1330 - 0x532  :  240 - 0xf0
    "11100000", -- 1331 - 0x533  :  224 - 0xe0
    "11000000", -- 1332 - 0x534  :  192 - 0xc0
    "10000000", -- 1333 - 0x535  :  128 - 0x80
    "10000000", -- 1334 - 0x536  :  128 - 0x80
    "00000000", -- 1335 - 0x537  :    0 - 0x0
    "11110000", -- 1336 - 0x538  :  240 - 0xf0 -- Background 0xa7
    "11111000", -- 1337 - 0x539  :  248 - 0xf8
    "11111100", -- 1338 - 0x53a  :  252 - 0xfc
    "11111110", -- 1339 - 0x53b  :  254 - 0xfe
    "10011111", -- 1340 - 0x53c  :  159 - 0x9f
    "10011111", -- 1341 - 0x53d  :  159 - 0x9f
    "11111111", -- 1342 - 0x53e  :  255 - 0xff
    "11111111", -- 1343 - 0x53f  :  255 - 0xff
    "11111111", -- 1344 - 0x540  :  255 - 0xff -- Background 0xa8
    "11111111", -- 1345 - 0x541  :  255 - 0xff
    "11111111", -- 1346 - 0x542  :  255 - 0xff
    "11111111", -- 1347 - 0x543  :  255 - 0xff
    "11111111", -- 1348 - 0x544  :  255 - 0xff
    "11111111", -- 1349 - 0x545  :  255 - 0xff
    "11111111", -- 1350 - 0x546  :  255 - 0xff
    "11111111", -- 1351 - 0x547  :  255 - 0xff
    "11111111", -- 1352 - 0x548  :  255 - 0xff -- Background 0xa9
    "11111111", -- 1353 - 0x549  :  255 - 0xff
    "11111111", -- 1354 - 0x54a  :  255 - 0xff
    "11111111", -- 1355 - 0x54b  :  255 - 0xff
    "11111111", -- 1356 - 0x54c  :  255 - 0xff
    "11111111", -- 1357 - 0x54d  :  255 - 0xff
    "11111111", -- 1358 - 0x54e  :  255 - 0xff
    "11111111", -- 1359 - 0x54f  :  255 - 0xff
    "11111111", -- 1360 - 0x550  :  255 - 0xff -- Background 0xaa
    "11111111", -- 1361 - 0x551  :  255 - 0xff
    "00001111", -- 1362 - 0x552  :   15 - 0xf
    "00000111", -- 1363 - 0x553  :    7 - 0x7
    "00000011", -- 1364 - 0x554  :    3 - 0x3
    "00000001", -- 1365 - 0x555  :    1 - 0x1
    "00000001", -- 1366 - 0x556  :    1 - 0x1
    "00000000", -- 1367 - 0x557  :    0 - 0x0
    "00000000", -- 1368 - 0x558  :    0 - 0x0 -- Background 0xab
    "00000000", -- 1369 - 0x559  :    0 - 0x0
    "00000000", -- 1370 - 0x55a  :    0 - 0x0
    "00000000", -- 1371 - 0x55b  :    0 - 0x0
    "10000000", -- 1372 - 0x55c  :  128 - 0x80
    "11000000", -- 1373 - 0x55d  :  192 - 0xc0
    "11111100", -- 1374 - 0x55e  :  252 - 0xfc
    "11111110", -- 1375 - 0x55f  :  254 - 0xfe
    "11111111", -- 1376 - 0x560  :  255 - 0xff -- Background 0xac
    "11111111", -- 1377 - 0x561  :  255 - 0xff
    "11111111", -- 1378 - 0x562  :  255 - 0xff
    "11111111", -- 1379 - 0x563  :  255 - 0xff
    "11111111", -- 1380 - 0x564  :  255 - 0xff
    "11111111", -- 1381 - 0x565  :  255 - 0xff
    "10111111", -- 1382 - 0x566  :  191 - 0xbf
    "10011111", -- 1383 - 0x567  :  159 - 0x9f
    "11001111", -- 1384 - 0x568  :  207 - 0xcf -- Background 0xad
    "11111111", -- 1385 - 0x569  :  255 - 0xff
    "11111111", -- 1386 - 0x56a  :  255 - 0xff
    "11111111", -- 1387 - 0x56b  :  255 - 0xff
    "11111111", -- 1388 - 0x56c  :  255 - 0xff
    "11111111", -- 1389 - 0x56d  :  255 - 0xff
    "11111111", -- 1390 - 0x56e  :  255 - 0xff
    "11111111", -- 1391 - 0x56f  :  255 - 0xff
    "11111111", -- 1392 - 0x570  :  255 - 0xff -- Background 0xae
    "11111111", -- 1393 - 0x571  :  255 - 0xff
    "11111111", -- 1394 - 0x572  :  255 - 0xff
    "11111111", -- 1395 - 0x573  :  255 - 0xff
    "11111111", -- 1396 - 0x574  :  255 - 0xff
    "11111111", -- 1397 - 0x575  :  255 - 0xff
    "11111111", -- 1398 - 0x576  :  255 - 0xff
    "11111111", -- 1399 - 0x577  :  255 - 0xff
    "00000000", -- 1400 - 0x578  :    0 - 0x0 -- Background 0xaf
    "10000000", -- 1401 - 0x579  :  128 - 0x80
    "11000000", -- 1402 - 0x57a  :  192 - 0xc0
    "11100000", -- 1403 - 0x57b  :  224 - 0xe0
    "11100000", -- 1404 - 0x57c  :  224 - 0xe0
    "11100000", -- 1405 - 0x57d  :  224 - 0xe0
    "11110000", -- 1406 - 0x57e  :  240 - 0xf0
    "11110000", -- 1407 - 0x57f  :  240 - 0xf0
    "11110000", -- 1408 - 0x580  :  240 - 0xf0 -- Background 0xb0
    "11110000", -- 1409 - 0x581  :  240 - 0xf0
    "11100000", -- 1410 - 0x582  :  224 - 0xe0
    "11100000", -- 1411 - 0x583  :  224 - 0xe0
    "11100000", -- 1412 - 0x584  :  224 - 0xe0
    "11000000", -- 1413 - 0x585  :  192 - 0xc0
    "11000000", -- 1414 - 0x586  :  192 - 0xc0
    "10000000", -- 1415 - 0x587  :  128 - 0x80
    "10000000", -- 1416 - 0x588  :  128 - 0x80 -- Background 0xb1
    "10000000", -- 1417 - 0x589  :  128 - 0x80
    "10000000", -- 1418 - 0x58a  :  128 - 0x80
    "00000000", -- 1419 - 0x58b  :    0 - 0x0
    "00000000", -- 1420 - 0x58c  :    0 - 0x0
    "11000000", -- 1421 - 0x58d  :  192 - 0xc0
    "11100000", -- 1422 - 0x58e  :  224 - 0xe0
    "11110000", -- 1423 - 0x58f  :  240 - 0xf0
    "00000000", -- 1424 - 0x590  :    0 - 0x0 -- Background 0xb2
    "00000000", -- 1425 - 0x591  :    0 - 0x0
    "00000001", -- 1426 - 0x592  :    1 - 0x1
    "00000011", -- 1427 - 0x593  :    3 - 0x3
    "00000111", -- 1428 - 0x594  :    7 - 0x7
    "00000111", -- 1429 - 0x595  :    7 - 0x7
    "00000111", -- 1430 - 0x596  :    7 - 0x7
    "00000111", -- 1431 - 0x597  :    7 - 0x7
    "00000011", -- 1432 - 0x598  :    3 - 0x3 -- Background 0xb3
    "00000001", -- 1433 - 0x599  :    1 - 0x1
    "00000000", -- 1434 - 0x59a  :    0 - 0x0
    "00000000", -- 1435 - 0x59b  :    0 - 0x0
    "00000000", -- 1436 - 0x59c  :    0 - 0x0
    "00000001", -- 1437 - 0x59d  :    1 - 0x1
    "00000011", -- 1438 - 0x59e  :    3 - 0x3
    "00000011", -- 1439 - 0x59f  :    3 - 0x3
    "00000011", -- 1440 - 0x5a0  :    3 - 0x3 -- Background 0xb4
    "00000011", -- 1441 - 0x5a1  :    3 - 0x3
    "00000111", -- 1442 - 0x5a2  :    7 - 0x7
    "00011111", -- 1443 - 0x5a3  :   31 - 0x1f
    "00111111", -- 1444 - 0x5a4  :   63 - 0x3f
    "00111111", -- 1445 - 0x5a5  :   63 - 0x3f
    "00000000", -- 1446 - 0x5a6  :    0 - 0x0
    "00000000", -- 1447 - 0x5a7  :    0 - 0x0
    "00000000", -- 1448 - 0x5a8  :    0 - 0x0 -- Background 0xb5
    "00000000", -- 1449 - 0x5a9  :    0 - 0x0
    "00000000", -- 1450 - 0x5aa  :    0 - 0x0
    "00000000", -- 1451 - 0x5ab  :    0 - 0x0
    "00000001", -- 1452 - 0x5ac  :    1 - 0x1
    "00000011", -- 1453 - 0x5ad  :    3 - 0x3
    "00000011", -- 1454 - 0x5ae  :    3 - 0x3
    "00001111", -- 1455 - 0x5af  :   15 - 0xf
    "00111111", -- 1456 - 0x5b0  :   63 - 0x3f -- Background 0xb6
    "01111111", -- 1457 - 0x5b1  :  127 - 0x7f
    "11111111", -- 1458 - 0x5b2  :  255 - 0xff
    "11111111", -- 1459 - 0x5b3  :  255 - 0xff
    "11111111", -- 1460 - 0x5b4  :  255 - 0xff
    "11111111", -- 1461 - 0x5b5  :  255 - 0xff
    "11111111", -- 1462 - 0x5b6  :  255 - 0xff
    "11111111", -- 1463 - 0x5b7  :  255 - 0xff
    "11111111", -- 1464 - 0x5b8  :  255 - 0xff -- Background 0xb7
    "11111111", -- 1465 - 0x5b9  :  255 - 0xff
    "11111111", -- 1466 - 0x5ba  :  255 - 0xff
    "00011111", -- 1467 - 0x5bb  :   31 - 0x1f
    "01111111", -- 1468 - 0x5bc  :  127 - 0x7f
    "11111111", -- 1469 - 0x5bd  :  255 - 0xff
    "11111111", -- 1470 - 0x5be  :  255 - 0xff
    "11111111", -- 1471 - 0x5bf  :  255 - 0xff
    "11111111", -- 1472 - 0x5c0  :  255 - 0xff -- Background 0xb8
    "11111111", -- 1473 - 0x5c1  :  255 - 0xff
    "11111111", -- 1474 - 0x5c2  :  255 - 0xff
    "11111100", -- 1475 - 0x5c3  :  252 - 0xfc
    "11111000", -- 1476 - 0x5c4  :  248 - 0xf8
    "11111000", -- 1477 - 0x5c5  :  248 - 0xf8
    "00000000", -- 1478 - 0x5c6  :    0 - 0x0
    "00000000", -- 1479 - 0x5c7  :    0 - 0x0
    "11001111", -- 1480 - 0x5c8  :  207 - 0xcf -- Background 0xb9
    "10001000", -- 1481 - 0x5c9  :  136 - 0x88
    "11011101", -- 1482 - 0x5ca  :  221 - 0xdd
    "11001000", -- 1483 - 0x5cb  :  200 - 0xc8
    "11111000", -- 1484 - 0x5cc  :  248 - 0xf8
    "11111111", -- 1485 - 0x5cd  :  255 - 0xff
    "11111111", -- 1486 - 0x5ce  :  255 - 0xff
    "11111111", -- 1487 - 0x5cf  :  255 - 0xff
    "11111111", -- 1488 - 0x5d0  :  255 - 0xff -- Background 0xba
    "11111111", -- 1489 - 0x5d1  :  255 - 0xff
    "11000000", -- 1490 - 0x5d2  :  192 - 0xc0
    "00000000", -- 1491 - 0x5d3  :    0 - 0x0
    "00000000", -- 1492 - 0x5d4  :    0 - 0x0
    "00000000", -- 1493 - 0x5d5  :    0 - 0x0
    "00000000", -- 1494 - 0x5d6  :    0 - 0x0
    "00000000", -- 1495 - 0x5d7  :    0 - 0x0
    "11111001", -- 1496 - 0x5d8  :  249 - 0xf9 -- Background 0xbb
    "10001000", -- 1497 - 0x5d9  :  136 - 0x88
    "11011101", -- 1498 - 0x5da  :  221 - 0xdd
    "10001001", -- 1499 - 0x5db  :  137 - 0x89
    "00001111", -- 1500 - 0x5dc  :   15 - 0xf
    "11111111", -- 1501 - 0x5dd  :  255 - 0xff
    "11111111", -- 1502 - 0x5de  :  255 - 0xff
    "11111111", -- 1503 - 0x5df  :  255 - 0xff
    "00000011", -- 1504 - 0x5e0  :    3 - 0x3 -- Background 0xbc
    "00000111", -- 1505 - 0x5e1  :    7 - 0x7
    "00001111", -- 1506 - 0x5e2  :   15 - 0xf
    "00000111", -- 1507 - 0x5e3  :    7 - 0x7
    "10000111", -- 1508 - 0x5e4  :  135 - 0x87
    "11000011", -- 1509 - 0x5e5  :  195 - 0xc3
    "11100000", -- 1510 - 0x5e6  :  224 - 0xe0
    "11111111", -- 1511 - 0x5e7  :  255 - 0xff
    "11111111", -- 1512 - 0x5e8  :  255 - 0xff -- Background 0xbd
    "11111111", -- 1513 - 0x5e9  :  255 - 0xff
    "11111111", -- 1514 - 0x5ea  :  255 - 0xff
    "11111111", -- 1515 - 0x5eb  :  255 - 0xff
    "11111111", -- 1516 - 0x5ec  :  255 - 0xff
    "11111111", -- 1517 - 0x5ed  :  255 - 0xff
    "11111111", -- 1518 - 0x5ee  :  255 - 0xff
    "11111110", -- 1519 - 0x5ef  :  254 - 0xfe
    "11111100", -- 1520 - 0x5f0  :  252 - 0xfc -- Background 0xbe
    "11111000", -- 1521 - 0x5f1  :  248 - 0xf8
    "11111000", -- 1522 - 0x5f2  :  248 - 0xf8
    "11111000", -- 1523 - 0x5f3  :  248 - 0xf8
    "11111000", -- 1524 - 0x5f4  :  248 - 0xf8
    "11111100", -- 1525 - 0x5f5  :  252 - 0xfc
    "11111110", -- 1526 - 0x5f6  :  254 - 0xfe
    "11111111", -- 1527 - 0x5f7  :  255 - 0xff
    "11111111", -- 1528 - 0x5f8  :  255 - 0xff -- Background 0xbf
    "11111111", -- 1529 - 0x5f9  :  255 - 0xff
    "11111111", -- 1530 - 0x5fa  :  255 - 0xff
    "11111111", -- 1531 - 0x5fb  :  255 - 0xff
    "11111111", -- 1532 - 0x5fc  :  255 - 0xff
    "11111111", -- 1533 - 0x5fd  :  255 - 0xff
    "11111111", -- 1534 - 0x5fe  :  255 - 0xff
    "11111111", -- 1535 - 0x5ff  :  255 - 0xff
    "11000000", -- 1536 - 0x600  :  192 - 0xc0 -- Background 0xc0
    "11110000", -- 1537 - 0x601  :  240 - 0xf0
    "11111100", -- 1538 - 0x602  :  252 - 0xfc
    "11111100", -- 1539 - 0x603  :  252 - 0xfc
    "11111110", -- 1540 - 0x604  :  254 - 0xfe
    "11111110", -- 1541 - 0x605  :  254 - 0xfe
    "11111110", -- 1542 - 0x606  :  254 - 0xfe
    "11111110", -- 1543 - 0x607  :  254 - 0xfe
    "11111111", -- 1544 - 0x608  :  255 - 0xff -- Background 0xc1
    "11111111", -- 1545 - 0x609  :  255 - 0xff
    "11111110", -- 1546 - 0x60a  :  254 - 0xfe
    "11111100", -- 1547 - 0x60b  :  252 - 0xfc
    "11110000", -- 1548 - 0x60c  :  240 - 0xf0
    "11100000", -- 1549 - 0x60d  :  224 - 0xe0
    "10000000", -- 1550 - 0x60e  :  128 - 0x80
    "00000000", -- 1551 - 0x60f  :    0 - 0x0
    "00000011", -- 1552 - 0x610  :    3 - 0x3 -- Background 0xc2
    "00001111", -- 1553 - 0x611  :   15 - 0xf
    "00111111", -- 1554 - 0x612  :   63 - 0x3f
    "00111111", -- 1555 - 0x613  :   63 - 0x3f
    "01111111", -- 1556 - 0x614  :  127 - 0x7f
    "01111111", -- 1557 - 0x615  :  127 - 0x7f
    "01111110", -- 1558 - 0x616  :  126 - 0x7e
    "11111111", -- 1559 - 0x617  :  255 - 0xff
    "11111111", -- 1560 - 0x618  :  255 - 0xff -- Background 0xc3
    "11111111", -- 1561 - 0x619  :  255 - 0xff
    "01111111", -- 1562 - 0x61a  :  127 - 0x7f
    "00111111", -- 1563 - 0x61b  :   63 - 0x3f
    "00001111", -- 1564 - 0x61c  :   15 - 0xf
    "00000111", -- 1565 - 0x61d  :    7 - 0x7
    "00000001", -- 1566 - 0x61e  :    1 - 0x1
    "00000000", -- 1567 - 0x61f  :    0 - 0x0
    "11000000", -- 1568 - 0x620  :  192 - 0xc0 -- Background 0xc4
    "11100000", -- 1569 - 0x621  :  224 - 0xe0
    "11110000", -- 1570 - 0x622  :  240 - 0xf0
    "11100000", -- 1571 - 0x623  :  224 - 0xe0
    "11100001", -- 1572 - 0x624  :  225 - 0xe1
    "11000011", -- 1573 - 0x625  :  195 - 0xc3
    "00000111", -- 1574 - 0x626  :    7 - 0x7
    "11111111", -- 1575 - 0x627  :  255 - 0xff
    "11111111", -- 1576 - 0x628  :  255 - 0xff -- Background 0xc5
    "11111111", -- 1577 - 0x629  :  255 - 0xff
    "11111111", -- 1578 - 0x62a  :  255 - 0xff
    "11111111", -- 1579 - 0x62b  :  255 - 0xff
    "11111111", -- 1580 - 0x62c  :  255 - 0xff
    "11111111", -- 1581 - 0x62d  :  255 - 0xff
    "11111111", -- 1582 - 0x62e  :  255 - 0xff
    "01111111", -- 1583 - 0x62f  :  127 - 0x7f
    "00111111", -- 1584 - 0x630  :   63 - 0x3f -- Background 0xc6
    "00011111", -- 1585 - 0x631  :   31 - 0x1f
    "00011111", -- 1586 - 0x632  :   31 - 0x1f
    "00011111", -- 1587 - 0x633  :   31 - 0x1f
    "00011111", -- 1588 - 0x634  :   31 - 0x1f
    "00111111", -- 1589 - 0x635  :   63 - 0x3f
    "01111111", -- 1590 - 0x636  :  127 - 0x7f
    "11111111", -- 1591 - 0x637  :  255 - 0xff
    "11111111", -- 1592 - 0x638  :  255 - 0xff -- Background 0xc7
    "11111111", -- 1593 - 0x639  :  255 - 0xff
    "11111111", -- 1594 - 0x63a  :  255 - 0xff
    "11111111", -- 1595 - 0x63b  :  255 - 0xff
    "11111111", -- 1596 - 0x63c  :  255 - 0xff
    "11111111", -- 1597 - 0x63d  :  255 - 0xff
    "11111111", -- 1598 - 0x63e  :  255 - 0xff
    "11111111", -- 1599 - 0x63f  :  255 - 0xff
    "11111111", -- 1600 - 0x640  :  255 - 0xff -- Background 0xc8
    "11111111", -- 1601 - 0x641  :  255 - 0xff
    "00000011", -- 1602 - 0x642  :    3 - 0x3
    "00000000", -- 1603 - 0x643  :    0 - 0x0
    "00000000", -- 1604 - 0x644  :    0 - 0x0
    "00000000", -- 1605 - 0x645  :    0 - 0x0
    "00000000", -- 1606 - 0x646  :    0 - 0x0
    "00000000", -- 1607 - 0x647  :    0 - 0x0
    "00000000", -- 1608 - 0x648  :    0 - 0x0 -- Background 0xc9
    "00000000", -- 1609 - 0x649  :    0 - 0x0
    "00000000", -- 1610 - 0x64a  :    0 - 0x0
    "00000000", -- 1611 - 0x64b  :    0 - 0x0
    "10000000", -- 1612 - 0x64c  :  128 - 0x80
    "11000000", -- 1613 - 0x64d  :  192 - 0xc0
    "11000000", -- 1614 - 0x64e  :  192 - 0xc0
    "11110000", -- 1615 - 0x64f  :  240 - 0xf0
    "11111100", -- 1616 - 0x650  :  252 - 0xfc -- Background 0xca
    "11111110", -- 1617 - 0x651  :  254 - 0xfe
    "11111111", -- 1618 - 0x652  :  255 - 0xff
    "11111111", -- 1619 - 0x653  :  255 - 0xff
    "11111111", -- 1620 - 0x654  :  255 - 0xff
    "11111111", -- 1621 - 0x655  :  255 - 0xff
    "11111111", -- 1622 - 0x656  :  255 - 0xff
    "11111111", -- 1623 - 0x657  :  255 - 0xff
    "11111111", -- 1624 - 0x658  :  255 - 0xff -- Background 0xcb
    "11111111", -- 1625 - 0x659  :  255 - 0xff
    "11111111", -- 1626 - 0x65a  :  255 - 0xff
    "11111000", -- 1627 - 0x65b  :  248 - 0xf8
    "11111110", -- 1628 - 0x65c  :  254 - 0xfe
    "11111111", -- 1629 - 0x65d  :  255 - 0xff
    "11111111", -- 1630 - 0x65e  :  255 - 0xff
    "11111111", -- 1631 - 0x65f  :  255 - 0xff
    "11111111", -- 1632 - 0x660  :  255 - 0xff -- Background 0xcc
    "11111111", -- 1633 - 0x661  :  255 - 0xff
    "11111111", -- 1634 - 0x662  :  255 - 0xff
    "00111111", -- 1635 - 0x663  :   63 - 0x3f
    "00011111", -- 1636 - 0x664  :   31 - 0x1f
    "00011111", -- 1637 - 0x665  :   31 - 0x1f
    "00000000", -- 1638 - 0x666  :    0 - 0x0
    "00000000", -- 1639 - 0x667  :    0 - 0x0
    "00000000", -- 1640 - 0x668  :    0 - 0x0 -- Background 0xcd
    "00000000", -- 1641 - 0x669  :    0 - 0x0
    "10000000", -- 1642 - 0x66a  :  128 - 0x80
    "11000000", -- 1643 - 0x66b  :  192 - 0xc0
    "11100000", -- 1644 - 0x66c  :  224 - 0xe0
    "11100000", -- 1645 - 0x66d  :  224 - 0xe0
    "11100000", -- 1646 - 0x66e  :  224 - 0xe0
    "11100000", -- 1647 - 0x66f  :  224 - 0xe0
    "11000000", -- 1648 - 0x670  :  192 - 0xc0 -- Background 0xce
    "10000000", -- 1649 - 0x671  :  128 - 0x80
    "00000000", -- 1650 - 0x672  :    0 - 0x0
    "00000000", -- 1651 - 0x673  :    0 - 0x0
    "00000000", -- 1652 - 0x674  :    0 - 0x0
    "10000000", -- 1653 - 0x675  :  128 - 0x80
    "11000000", -- 1654 - 0x676  :  192 - 0xc0
    "11000000", -- 1655 - 0x677  :  192 - 0xc0
    "11000000", -- 1656 - 0x678  :  192 - 0xc0 -- Background 0xcf
    "11000000", -- 1657 - 0x679  :  192 - 0xc0
    "11100000", -- 1658 - 0x67a  :  224 - 0xe0
    "11111000", -- 1659 - 0x67b  :  248 - 0xf8
    "11111100", -- 1660 - 0x67c  :  252 - 0xfc
    "11111100", -- 1661 - 0x67d  :  252 - 0xfc
    "00000000", -- 1662 - 0x67e  :    0 - 0x0
    "00000000", -- 1663 - 0x67f  :    0 - 0x0
    "00000000", -- 1664 - 0x680  :    0 - 0x0 -- Background 0xd0
    "00000000", -- 1665 - 0x681  :    0 - 0x0
    "00000000", -- 1666 - 0x682  :    0 - 0x0
    "00000000", -- 1667 - 0x683  :    0 - 0x0
    "00000000", -- 1668 - 0x684  :    0 - 0x0
    "00000000", -- 1669 - 0x685  :    0 - 0x0
    "00000000", -- 1670 - 0x686  :    0 - 0x0
    "00000000", -- 1671 - 0x687  :    0 - 0x0
    "00000000", -- 1672 - 0x688  :    0 - 0x0 -- Background 0xd1
    "00000000", -- 1673 - 0x689  :    0 - 0x0
    "00000000", -- 1674 - 0x68a  :    0 - 0x0
    "00000000", -- 1675 - 0x68b  :    0 - 0x0
    "00000000", -- 1676 - 0x68c  :    0 - 0x0
    "00000000", -- 1677 - 0x68d  :    0 - 0x0
    "00000000", -- 1678 - 0x68e  :    0 - 0x0
    "00000000", -- 1679 - 0x68f  :    0 - 0x0
    "00000000", -- 1680 - 0x690  :    0 - 0x0 -- Background 0xd2
    "00000000", -- 1681 - 0x691  :    0 - 0x0
    "00000000", -- 1682 - 0x692  :    0 - 0x0
    "00000000", -- 1683 - 0x693  :    0 - 0x0
    "00000000", -- 1684 - 0x694  :    0 - 0x0
    "00000000", -- 1685 - 0x695  :    0 - 0x0
    "00000000", -- 1686 - 0x696  :    0 - 0x0
    "00000000", -- 1687 - 0x697  :    0 - 0x0
    "00000000", -- 1688 - 0x698  :    0 - 0x0 -- Background 0xd3
    "00000000", -- 1689 - 0x699  :    0 - 0x0
    "00000000", -- 1690 - 0x69a  :    0 - 0x0
    "00000000", -- 1691 - 0x69b  :    0 - 0x0
    "00000000", -- 1692 - 0x69c  :    0 - 0x0
    "00000000", -- 1693 - 0x69d  :    0 - 0x0
    "00000000", -- 1694 - 0x69e  :    0 - 0x0
    "00000000", -- 1695 - 0x69f  :    0 - 0x0
    "00000000", -- 1696 - 0x6a0  :    0 - 0x0 -- Background 0xd4
    "00000000", -- 1697 - 0x6a1  :    0 - 0x0
    "00000000", -- 1698 - 0x6a2  :    0 - 0x0
    "00000000", -- 1699 - 0x6a3  :    0 - 0x0
    "00000011", -- 1700 - 0x6a4  :    3 - 0x3
    "00000111", -- 1701 - 0x6a5  :    7 - 0x7
    "00000011", -- 1702 - 0x6a6  :    3 - 0x3
    "00000111", -- 1703 - 0x6a7  :    7 - 0x7
    "00011111", -- 1704 - 0x6a8  :   31 - 0x1f -- Background 0xd5
    "00111111", -- 1705 - 0x6a9  :   63 - 0x3f
    "01111111", -- 1706 - 0x6aa  :  127 - 0x7f
    "11111111", -- 1707 - 0x6ab  :  255 - 0xff
    "11111111", -- 1708 - 0x6ac  :  255 - 0xff
    "11111111", -- 1709 - 0x6ad  :  255 - 0xff
    "11111111", -- 1710 - 0x6ae  :  255 - 0xff
    "01111111", -- 1711 - 0x6af  :  127 - 0x7f
    "00000000", -- 1712 - 0x6b0  :    0 - 0x0 -- Background 0xd6
    "00000000", -- 1713 - 0x6b1  :    0 - 0x0
    "00000000", -- 1714 - 0x6b2  :    0 - 0x0
    "11000000", -- 1715 - 0x6b3  :  192 - 0xc0
    "11100000", -- 1716 - 0x6b4  :  224 - 0xe0
    "11110000", -- 1717 - 0x6b5  :  240 - 0xf0
    "11110000", -- 1718 - 0x6b6  :  240 - 0xf0
    "11111000", -- 1719 - 0x6b7  :  248 - 0xf8
    "11111100", -- 1720 - 0x6b8  :  252 - 0xfc -- Background 0xd7
    "11111000", -- 1721 - 0x6b9  :  248 - 0xf8
    "11110000", -- 1722 - 0x6ba  :  240 - 0xf0
    "11111111", -- 1723 - 0x6bb  :  255 - 0xff
    "11111111", -- 1724 - 0x6bc  :  255 - 0xff
    "11111111", -- 1725 - 0x6bd  :  255 - 0xff
    "11111111", -- 1726 - 0x6be  :  255 - 0xff
    "11111111", -- 1727 - 0x6bf  :  255 - 0xff
    "00000000", -- 1728 - 0x6c0  :    0 - 0x0 -- Background 0xd8
    "00000000", -- 1729 - 0x6c1  :    0 - 0x0
    "00000000", -- 1730 - 0x6c2  :    0 - 0x0
    "00000000", -- 1731 - 0x6c3  :    0 - 0x0
    "00000011", -- 1732 - 0x6c4  :    3 - 0x3
    "00000111", -- 1733 - 0x6c5  :    7 - 0x7
    "00001111", -- 1734 - 0x6c6  :   15 - 0xf
    "00011111", -- 1735 - 0x6c7  :   31 - 0x1f
    "00111111", -- 1736 - 0x6c8  :   63 - 0x3f -- Background 0xd9
    "00011111", -- 1737 - 0x6c9  :   31 - 0x1f
    "00000111", -- 1738 - 0x6ca  :    7 - 0x7
    "11111111", -- 1739 - 0x6cb  :  255 - 0xff
    "11111111", -- 1740 - 0x6cc  :  255 - 0xff
    "11111111", -- 1741 - 0x6cd  :  255 - 0xff
    "11111111", -- 1742 - 0x6ce  :  255 - 0xff
    "11111111", -- 1743 - 0x6cf  :  255 - 0xff
    "00000000", -- 1744 - 0x6d0  :    0 - 0x0 -- Background 0xda
    "00000000", -- 1745 - 0x6d1  :    0 - 0x0
    "00000000", -- 1746 - 0x6d2  :    0 - 0x0
    "11000000", -- 1747 - 0x6d3  :  192 - 0xc0
    "11000000", -- 1748 - 0x6d4  :  192 - 0xc0
    "11000000", -- 1749 - 0x6d5  :  192 - 0xc0
    "11100000", -- 1750 - 0x6d6  :  224 - 0xe0
    "11111000", -- 1751 - 0x6d7  :  248 - 0xf8
    "11111100", -- 1752 - 0x6d8  :  252 - 0xfc -- Background 0xdb
    "11111110", -- 1753 - 0x6d9  :  254 - 0xfe
    "11111110", -- 1754 - 0x6da  :  254 - 0xfe
    "11111111", -- 1755 - 0x6db  :  255 - 0xff
    "11111111", -- 1756 - 0x6dc  :  255 - 0xff
    "11111111", -- 1757 - 0x6dd  :  255 - 0xff
    "11111111", -- 1758 - 0x6de  :  255 - 0xff
    "11111110", -- 1759 - 0x6df  :  254 - 0xfe
    "00110110", -- 1760 - 0x6e0  :   54 - 0x36 -- Background 0xdc
    "00110110", -- 1761 - 0x6e1  :   54 - 0x36
    "01111110", -- 1762 - 0x6e2  :  126 - 0x7e
    "01111111", -- 1763 - 0x6e3  :  127 - 0x7f
    "01111111", -- 1764 - 0x6e4  :  127 - 0x7f
    "01111111", -- 1765 - 0x6e5  :  127 - 0x7f
    "00111111", -- 1766 - 0x6e6  :   63 - 0x3f
    "00111111", -- 1767 - 0x6e7  :   63 - 0x3f
    "00111111", -- 1768 - 0x6e8  :   63 - 0x3f -- Background 0xdd
    "00011111", -- 1769 - 0x6e9  :   31 - 0x1f
    "00011111", -- 1770 - 0x6ea  :   31 - 0x1f
    "00001111", -- 1771 - 0x6eb  :   15 - 0xf
    "00000111", -- 1772 - 0x6ec  :    7 - 0x7
    "00000011", -- 1773 - 0x6ed  :    3 - 0x3
    "00000000", -- 1774 - 0x6ee  :    0 - 0x0
    "00000000", -- 1775 - 0x6ef  :    0 - 0x0
    "00111111", -- 1776 - 0x6f0  :   63 - 0x3f -- Background 0xde
    "00011111", -- 1777 - 0x6f1  :   31 - 0x1f
    "11011111", -- 1778 - 0x6f2  :  223 - 0xdf
    "11001111", -- 1779 - 0x6f3  :  207 - 0xcf
    "11001111", -- 1780 - 0x6f4  :  207 - 0xcf
    "10011111", -- 1781 - 0x6f5  :  159 - 0x9f
    "11011111", -- 1782 - 0x6f6  :  223 - 0xdf
    "11111111", -- 1783 - 0x6f7  :  255 - 0xff
    "11111111", -- 1784 - 0x6f8  :  255 - 0xff -- Background 0xdf
    "11111111", -- 1785 - 0x6f9  :  255 - 0xff
    "11111111", -- 1786 - 0x6fa  :  255 - 0xff
    "11111111", -- 1787 - 0x6fb  :  255 - 0xff
    "11111111", -- 1788 - 0x6fc  :  255 - 0xff
    "11111111", -- 1789 - 0x6fd  :  255 - 0xff
    "11111111", -- 1790 - 0x6fe  :  255 - 0xff
    "00001111", -- 1791 - 0x6ff  :   15 - 0xf
    "11111111", -- 1792 - 0x700  :  255 - 0xff -- Background 0xe0
    "11111111", -- 1793 - 0x701  :  255 - 0xff
    "11111111", -- 1794 - 0x702  :  255 - 0xff
    "11111111", -- 1795 - 0x703  :  255 - 0xff
    "11111111", -- 1796 - 0x704  :  255 - 0xff
    "11111111", -- 1797 - 0x705  :  255 - 0xff
    "11111111", -- 1798 - 0x706  :  255 - 0xff
    "11111111", -- 1799 - 0x707  :  255 - 0xff
    "11111111", -- 1800 - 0x708  :  255 - 0xff -- Background 0xe1
    "11111001", -- 1801 - 0x709  :  249 - 0xf9
    "11110000", -- 1802 - 0x70a  :  240 - 0xf0
    "11110000", -- 1803 - 0x70b  :  240 - 0xf0
    "10110001", -- 1804 - 0x70c  :  177 - 0xb1
    "11011111", -- 1805 - 0x70d  :  223 - 0xdf
    "11101111", -- 1806 - 0x70e  :  239 - 0xef
    "10000111", -- 1807 - 0x70f  :  135 - 0x87
    "11111111", -- 1808 - 0x710  :  255 - 0xff -- Background 0xe2
    "11111111", -- 1809 - 0x711  :  255 - 0xff
    "11111111", -- 1810 - 0x712  :  255 - 0xff
    "11111111", -- 1811 - 0x713  :  255 - 0xff
    "11111111", -- 1812 - 0x714  :  255 - 0xff
    "11111111", -- 1813 - 0x715  :  255 - 0xff
    "11111111", -- 1814 - 0x716  :  255 - 0xff
    "11111111", -- 1815 - 0x717  :  255 - 0xff
    "11111111", -- 1816 - 0x718  :  255 - 0xff -- Background 0xe3
    "11001111", -- 1817 - 0x719  :  207 - 0xcf
    "10000111", -- 1818 - 0x71a  :  135 - 0x87
    "10000111", -- 1819 - 0x71b  :  135 - 0x87
    "11001110", -- 1820 - 0x71c  :  206 - 0xce
    "11111101", -- 1821 - 0x71d  :  253 - 0xfd
    "11111011", -- 1822 - 0x71e  :  251 - 0xfb
    "11110000", -- 1823 - 0x71f  :  240 - 0xf0
    "11111110", -- 1824 - 0x720  :  254 - 0xfe -- Background 0xe4
    "11111100", -- 1825 - 0x721  :  252 - 0xfc
    "11111100", -- 1826 - 0x722  :  252 - 0xfc
    "11111000", -- 1827 - 0x723  :  248 - 0xf8
    "11111011", -- 1828 - 0x724  :  251 - 0xfb
    "11111101", -- 1829 - 0x725  :  253 - 0xfd
    "11111110", -- 1830 - 0x726  :  254 - 0xfe
    "11111111", -- 1831 - 0x727  :  255 - 0xff
    "11111111", -- 1832 - 0x728  :  255 - 0xff -- Background 0xe5
    "11111111", -- 1833 - 0x729  :  255 - 0xff
    "11111111", -- 1834 - 0x72a  :  255 - 0xff
    "11111111", -- 1835 - 0x72b  :  255 - 0xff
    "11111111", -- 1836 - 0x72c  :  255 - 0xff
    "11111111", -- 1837 - 0x72d  :  255 - 0xff
    "11111111", -- 1838 - 0x72e  :  255 - 0xff
    "11111001", -- 1839 - 0x72f  :  249 - 0xf9
    "00000000", -- 1840 - 0x730  :    0 - 0x0 -- Background 0xe6
    "00000000", -- 1841 - 0x731  :    0 - 0x0
    "00000000", -- 1842 - 0x732  :    0 - 0x0
    "01111000", -- 1843 - 0x733  :  120 - 0x78
    "11111100", -- 1844 - 0x734  :  252 - 0xfc
    "11111100", -- 1845 - 0x735  :  252 - 0xfc
    "11111100", -- 1846 - 0x736  :  252 - 0xfc
    "11111100", -- 1847 - 0x737  :  252 - 0xfc
    "11111110", -- 1848 - 0x738  :  254 - 0xfe -- Background 0xe7
    "11111110", -- 1849 - 0x739  :  254 - 0xfe
    "11111110", -- 1850 - 0x73a  :  254 - 0xfe
    "11111110", -- 1851 - 0x73b  :  254 - 0xfe
    "11111110", -- 1852 - 0x73c  :  254 - 0xfe
    "11111100", -- 1853 - 0x73d  :  252 - 0xfc
    "11111000", -- 1854 - 0x73e  :  248 - 0xf8
    "11110000", -- 1855 - 0x73f  :  240 - 0xf0
    "00000000", -- 1856 - 0x740  :    0 - 0x0 -- Background 0xe8
    "00000000", -- 1857 - 0x741  :    0 - 0x0
    "00000000", -- 1858 - 0x742  :    0 - 0x0
    "00000000", -- 1859 - 0x743  :    0 - 0x0
    "00000000", -- 1860 - 0x744  :    0 - 0x0
    "00000000", -- 1861 - 0x745  :    0 - 0x0
    "00000000", -- 1862 - 0x746  :    0 - 0x0
    "00000000", -- 1863 - 0x747  :    0 - 0x0
    "00000001", -- 1864 - 0x748  :    1 - 0x1 -- Background 0xe9
    "00001111", -- 1865 - 0x749  :   15 - 0xf
    "00011111", -- 1866 - 0x74a  :   31 - 0x1f
    "00011111", -- 1867 - 0x74b  :   31 - 0x1f
    "00111011", -- 1868 - 0x74c  :   59 - 0x3b
    "00110011", -- 1869 - 0x74d  :   51 - 0x33
    "00000001", -- 1870 - 0x74e  :    1 - 0x1
    "00000001", -- 1871 - 0x74f  :    1 - 0x1
    "00000000", -- 1872 - 0x750  :    0 - 0x0 -- Background 0xea
    "00000000", -- 1873 - 0x751  :    0 - 0x0
    "00000000", -- 1874 - 0x752  :    0 - 0x0
    "00110110", -- 1875 - 0x753  :   54 - 0x36
    "01101100", -- 1876 - 0x754  :  108 - 0x6c
    "11111101", -- 1877 - 0x755  :  253 - 0xfd
    "11111111", -- 1878 - 0x756  :  255 - 0xff
    "11111111", -- 1879 - 0x757  :  255 - 0xff
    "11111111", -- 1880 - 0x758  :  255 - 0xff -- Background 0xeb
    "01111111", -- 1881 - 0x759  :  127 - 0x7f
    "01111111", -- 1882 - 0x75a  :  127 - 0x7f
    "01111111", -- 1883 - 0x75b  :  127 - 0x7f
    "01111111", -- 1884 - 0x75c  :  127 - 0x7f
    "00111111", -- 1885 - 0x75d  :   63 - 0x3f
    "00011111", -- 1886 - 0x75e  :   31 - 0x1f
    "00000111", -- 1887 - 0x75f  :    7 - 0x7
    "00000000", -- 1888 - 0x760  :    0 - 0x0 -- Background 0xec
    "00000000", -- 1889 - 0x761  :    0 - 0x0
    "00000000", -- 1890 - 0x762  :    0 - 0x0
    "00000000", -- 1891 - 0x763  :    0 - 0x0
    "00000000", -- 1892 - 0x764  :    0 - 0x0
    "00000000", -- 1893 - 0x765  :    0 - 0x0
    "00000000", -- 1894 - 0x766  :    0 - 0x0
    "11100000", -- 1895 - 0x767  :  224 - 0xe0
    "11111000", -- 1896 - 0x768  :  248 - 0xf8 -- Background 0xed
    "11111111", -- 1897 - 0x769  :  255 - 0xff
    "11111111", -- 1898 - 0x76a  :  255 - 0xff
    "11111111", -- 1899 - 0x76b  :  255 - 0xff
    "11111111", -- 1900 - 0x76c  :  255 - 0xff
    "11111111", -- 1901 - 0x76d  :  255 - 0xff
    "11111111", -- 1902 - 0x76e  :  255 - 0xff
    "11111111", -- 1903 - 0x76f  :  255 - 0xff
    "11111111", -- 1904 - 0x770  :  255 - 0xff -- Background 0xee
    "01111111", -- 1905 - 0x771  :  127 - 0x7f
    "00011111", -- 1906 - 0x772  :   31 - 0x1f
    "00001111", -- 1907 - 0x773  :   15 - 0xf
    "00001111", -- 1908 - 0x774  :   15 - 0xf
    "10011111", -- 1909 - 0x775  :  159 - 0x9f
    "10011111", -- 1910 - 0x776  :  159 - 0x9f
    "10111111", -- 1911 - 0x777  :  191 - 0xbf
    "01111111", -- 1912 - 0x778  :  127 - 0x7f -- Background 0xef
    "11111111", -- 1913 - 0x779  :  255 - 0xff
    "11111111", -- 1914 - 0x77a  :  255 - 0xff
    "11111111", -- 1915 - 0x77b  :  255 - 0xff
    "11111111", -- 1916 - 0x77c  :  255 - 0xff
    "11111111", -- 1917 - 0x77d  :  255 - 0xff
    "11111111", -- 1918 - 0x77e  :  255 - 0xff
    "11001111", -- 1919 - 0x77f  :  207 - 0xcf
    "00000000", -- 1920 - 0x780  :    0 - 0x0 -- Background 0xf0
    "00000000", -- 1921 - 0x781  :    0 - 0x0
    "11110000", -- 1922 - 0x782  :  240 - 0xf0
    "11111111", -- 1923 - 0x783  :  255 - 0xff
    "11111111", -- 1924 - 0x784  :  255 - 0xff
    "11111111", -- 1925 - 0x785  :  255 - 0xff
    "11111111", -- 1926 - 0x786  :  255 - 0xff
    "11111111", -- 1927 - 0x787  :  255 - 0xff
    "11111111", -- 1928 - 0x788  :  255 - 0xff -- Background 0xf1
    "11111111", -- 1929 - 0x789  :  255 - 0xff
    "11111111", -- 1930 - 0x78a  :  255 - 0xff
    "11110001", -- 1931 - 0x78b  :  241 - 0xf1
    "11000100", -- 1932 - 0x78c  :  196 - 0xc4
    "11101110", -- 1933 - 0x78d  :  238 - 0xee
    "11000100", -- 1934 - 0x78e  :  196 - 0xc4
    "10000011", -- 1935 - 0x78f  :  131 - 0x83
    "11000111", -- 1936 - 0x790  :  199 - 0xc7 -- Background 0xf2
    "11111001", -- 1937 - 0x791  :  249 - 0xf9
    "11110000", -- 1938 - 0x792  :  240 - 0xf0
    "11110000", -- 1939 - 0x793  :  240 - 0xf0
    "10110001", -- 1940 - 0x794  :  177 - 0xb1
    "11011111", -- 1941 - 0x795  :  223 - 0xdf
    "11101111", -- 1942 - 0x796  :  239 - 0xef
    "10000111", -- 1943 - 0x797  :  135 - 0x87
    "00000000", -- 1944 - 0x798  :    0 - 0x0 -- Background 0xf3
    "00000000", -- 1945 - 0x799  :    0 - 0x0
    "00000111", -- 1946 - 0x79a  :    7 - 0x7
    "11111111", -- 1947 - 0x79b  :  255 - 0xff
    "11111111", -- 1948 - 0x79c  :  255 - 0xff
    "11111111", -- 1949 - 0x79d  :  255 - 0xff
    "11111111", -- 1950 - 0x79e  :  255 - 0xff
    "11111111", -- 1951 - 0x79f  :  255 - 0xff
    "11111111", -- 1952 - 0x7a0  :  255 - 0xff -- Background 0xf4
    "11111111", -- 1953 - 0x7a1  :  255 - 0xff
    "11111111", -- 1954 - 0x7a2  :  255 - 0xff
    "11000111", -- 1955 - 0x7a3  :  199 - 0xc7
    "01000101", -- 1956 - 0x7a4  :   69 - 0x45
    "11101110", -- 1957 - 0x7a5  :  238 - 0xee
    "01000100", -- 1958 - 0x7a6  :   68 - 0x44
    "11100001", -- 1959 - 0x7a7  :  225 - 0xe1
    "11111111", -- 1960 - 0x7a8  :  255 - 0xff -- Background 0xf5
    "11001111", -- 1961 - 0x7a9  :  207 - 0xcf
    "10000111", -- 1962 - 0x7aa  :  135 - 0x87
    "10000111", -- 1963 - 0x7ab  :  135 - 0x87
    "11001110", -- 1964 - 0x7ac  :  206 - 0xce
    "11111101", -- 1965 - 0x7ad  :  253 - 0xfd
    "11111011", -- 1966 - 0x7ae  :  251 - 0xfb
    "11110000", -- 1967 - 0x7af  :  240 - 0xf0
    "00000000", -- 1968 - 0x7b0  :    0 - 0x0 -- Background 0xf6
    "00000000", -- 1969 - 0x7b1  :    0 - 0x0
    "00000000", -- 1970 - 0x7b2  :    0 - 0x0
    "00000000", -- 1971 - 0x7b3  :    0 - 0x0
    "00000000", -- 1972 - 0x7b4  :    0 - 0x0
    "00000001", -- 1973 - 0x7b5  :    1 - 0x1
    "00000111", -- 1974 - 0x7b6  :    7 - 0x7
    "00001111", -- 1975 - 0x7b7  :   15 - 0xf
    "00111111", -- 1976 - 0x7b8  :   63 - 0x3f -- Background 0xf7
    "11111111", -- 1977 - 0x7b9  :  255 - 0xff
    "11111111", -- 1978 - 0x7ba  :  255 - 0xff
    "11111111", -- 1979 - 0x7bb  :  255 - 0xff
    "11111111", -- 1980 - 0x7bc  :  255 - 0xff
    "11111111", -- 1981 - 0x7bd  :  255 - 0xff
    "11111111", -- 1982 - 0x7be  :  255 - 0xff
    "11111111", -- 1983 - 0x7bf  :  255 - 0xff
    "11111111", -- 1984 - 0x7c0  :  255 - 0xff -- Background 0xf8
    "11111111", -- 1985 - 0x7c1  :  255 - 0xff
    "11111101", -- 1986 - 0x7c2  :  253 - 0xfd
    "11111000", -- 1987 - 0x7c3  :  248 - 0xf8
    "11111111", -- 1988 - 0x7c4  :  255 - 0xff
    "11111111", -- 1989 - 0x7c5  :  255 - 0xff
    "11111110", -- 1990 - 0x7c6  :  254 - 0xfe
    "11111111", -- 1991 - 0x7c7  :  255 - 0xff
    "11111111", -- 1992 - 0x7c8  :  255 - 0xff -- Background 0xf9
    "11111111", -- 1993 - 0x7c9  :  255 - 0xff
    "11111111", -- 1994 - 0x7ca  :  255 - 0xff
    "11111111", -- 1995 - 0x7cb  :  255 - 0xff
    "11111111", -- 1996 - 0x7cc  :  255 - 0xff
    "11111111", -- 1997 - 0x7cd  :  255 - 0xff
    "11111111", -- 1998 - 0x7ce  :  255 - 0xff
    "11111000", -- 1999 - 0x7cf  :  248 - 0xf8
    "00000000", -- 2000 - 0x7d0  :    0 - 0x0 -- Background 0xfa
    "00000000", -- 2001 - 0x7d1  :    0 - 0x0
    "00000000", -- 2002 - 0x7d2  :    0 - 0x0
    "00000000", -- 2003 - 0x7d3  :    0 - 0x0
    "00000000", -- 2004 - 0x7d4  :    0 - 0x0
    "00000000", -- 2005 - 0x7d5  :    0 - 0x0
    "11000000", -- 2006 - 0x7d6  :  192 - 0xc0
    "11110000", -- 2007 - 0x7d7  :  240 - 0xf0
    "11111100", -- 2008 - 0x7d8  :  252 - 0xfc -- Background 0xfb
    "11111110", -- 2009 - 0x7d9  :  254 - 0xfe
    "11101100", -- 2010 - 0x7da  :  236 - 0xec
    "11100000", -- 2011 - 0x7db  :  224 - 0xe0
    "11000000", -- 2012 - 0x7dc  :  192 - 0xc0
    "11000000", -- 2013 - 0x7dd  :  192 - 0xc0
    "10000000", -- 2014 - 0x7de  :  128 - 0x80
    "10000000", -- 2015 - 0x7df  :  128 - 0x80
    "01110000", -- 2016 - 0x7e0  :  112 - 0x70 -- Background 0xfc
    "11111100", -- 2017 - 0x7e1  :  252 - 0xfc
    "11111100", -- 2018 - 0x7e2  :  252 - 0xfc
    "11111100", -- 2019 - 0x7e3  :  252 - 0xfc
    "11111100", -- 2020 - 0x7e4  :  252 - 0xfc
    "11111100", -- 2021 - 0x7e5  :  252 - 0xfc
    "11111110", -- 2022 - 0x7e6  :  254 - 0xfe
    "11111110", -- 2023 - 0x7e7  :  254 - 0xfe
    "11111110", -- 2024 - 0x7e8  :  254 - 0xfe -- Background 0xfd
    "11111100", -- 2025 - 0x7e9  :  252 - 0xfc
    "11111100", -- 2026 - 0x7ea  :  252 - 0xfc
    "11111000", -- 2027 - 0x7eb  :  248 - 0xf8
    "11110000", -- 2028 - 0x7ec  :  240 - 0xf0
    "11100000", -- 2029 - 0x7ed  :  224 - 0xe0
    "10000000", -- 2030 - 0x7ee  :  128 - 0x80
    "00000000", -- 2031 - 0x7ef  :    0 - 0x0
    "00000000", -- 2032 - 0x7f0  :    0 - 0x0 -- Background 0xfe
    "00000000", -- 2033 - 0x7f1  :    0 - 0x0
    "00000000", -- 2034 - 0x7f2  :    0 - 0x0
    "00000000", -- 2035 - 0x7f3  :    0 - 0x0
    "00000000", -- 2036 - 0x7f4  :    0 - 0x0
    "00000000", -- 2037 - 0x7f5  :    0 - 0x0
    "00000000", -- 2038 - 0x7f6  :    0 - 0x0
    "00000000", -- 2039 - 0x7f7  :    0 - 0x0
    "00000000", -- 2040 - 0x7f8  :    0 - 0x0 -- Background 0xff
    "00000000", -- 2041 - 0x7f9  :    0 - 0x0
    "00000000", -- 2042 - 0x7fa  :    0 - 0x0
    "00000000", -- 2043 - 0x7fb  :    0 - 0x0
    "00000000", -- 2044 - 0x7fc  :    0 - 0x0
    "00000000", -- 2045 - 0x7fd  :    0 - 0x0
    "00000000", -- 2046 - 0x7fe  :    0 - 0x0
    "00000000"  -- 2047 - 0x7ff  :    0 - 0x0
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
