//-   Background Pattern table COLOR PLANE 1
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
//- Autcmatically generated verilog ROM from a NES memory file----


//-  Original memory dump file name: donkeykong_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_PTABLE_DONKEYKONG_BG_PLN1
  (
     input     clk,   // clock
     input      [11-1:0] addr,  //2048 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Background pattern Table COLOR PLANE 1
      11'h0: dout <= 8'b00000000; //    0 :   0 - 0x0 -- Background 0x0
      11'h1: dout <= 8'b00000000; //    1 :   0 - 0x0
      11'h2: dout <= 8'b00000000; //    2 :   0 - 0x0
      11'h3: dout <= 8'b00000000; //    3 :   0 - 0x0
      11'h4: dout <= 8'b00000000; //    4 :   0 - 0x0
      11'h5: dout <= 8'b00000000; //    5 :   0 - 0x0
      11'h6: dout <= 8'b00000000; //    6 :   0 - 0x0
      11'h7: dout <= 8'b00000000; //    7 :   0 - 0x0
      11'h8: dout <= 8'b00000000; //    8 :   0 - 0x0 -- Background 0x1
      11'h9: dout <= 8'b00000000; //    9 :   0 - 0x0
      11'hA: dout <= 8'b00000000; //   10 :   0 - 0x0
      11'hB: dout <= 8'b00000000; //   11 :   0 - 0x0
      11'hC: dout <= 8'b00000000; //   12 :   0 - 0x0
      11'hD: dout <= 8'b00000000; //   13 :   0 - 0x0
      11'hE: dout <= 8'b00000000; //   14 :   0 - 0x0
      11'hF: dout <= 8'b00000000; //   15 :   0 - 0x0
      11'h10: dout <= 8'b00000000; //   16 :   0 - 0x0 -- Background 0x2
      11'h11: dout <= 8'b00000000; //   17 :   0 - 0x0
      11'h12: dout <= 8'b00000000; //   18 :   0 - 0x0
      11'h13: dout <= 8'b00000000; //   19 :   0 - 0x0
      11'h14: dout <= 8'b00000000; //   20 :   0 - 0x0
      11'h15: dout <= 8'b00000000; //   21 :   0 - 0x0
      11'h16: dout <= 8'b00000000; //   22 :   0 - 0x0
      11'h17: dout <= 8'b00000000; //   23 :   0 - 0x0
      11'h18: dout <= 8'b00000000; //   24 :   0 - 0x0 -- Background 0x3
      11'h19: dout <= 8'b00000000; //   25 :   0 - 0x0
      11'h1A: dout <= 8'b00000000; //   26 :   0 - 0x0
      11'h1B: dout <= 8'b00000000; //   27 :   0 - 0x0
      11'h1C: dout <= 8'b00000000; //   28 :   0 - 0x0
      11'h1D: dout <= 8'b00000000; //   29 :   0 - 0x0
      11'h1E: dout <= 8'b00000000; //   30 :   0 - 0x0
      11'h1F: dout <= 8'b00000000; //   31 :   0 - 0x0
      11'h20: dout <= 8'b00000000; //   32 :   0 - 0x0 -- Background 0x4
      11'h21: dout <= 8'b00000000; //   33 :   0 - 0x0
      11'h22: dout <= 8'b00000000; //   34 :   0 - 0x0
      11'h23: dout <= 8'b00000000; //   35 :   0 - 0x0
      11'h24: dout <= 8'b00000000; //   36 :   0 - 0x0
      11'h25: dout <= 8'b00000000; //   37 :   0 - 0x0
      11'h26: dout <= 8'b00000000; //   38 :   0 - 0x0
      11'h27: dout <= 8'b00000000; //   39 :   0 - 0x0
      11'h28: dout <= 8'b00000000; //   40 :   0 - 0x0 -- Background 0x5
      11'h29: dout <= 8'b00000000; //   41 :   0 - 0x0
      11'h2A: dout <= 8'b00000000; //   42 :   0 - 0x0
      11'h2B: dout <= 8'b00000000; //   43 :   0 - 0x0
      11'h2C: dout <= 8'b00000000; //   44 :   0 - 0x0
      11'h2D: dout <= 8'b00000000; //   45 :   0 - 0x0
      11'h2E: dout <= 8'b00000000; //   46 :   0 - 0x0
      11'h2F: dout <= 8'b00000000; //   47 :   0 - 0x0
      11'h30: dout <= 8'b00000000; //   48 :   0 - 0x0 -- Background 0x6
      11'h31: dout <= 8'b00000000; //   49 :   0 - 0x0
      11'h32: dout <= 8'b00000000; //   50 :   0 - 0x0
      11'h33: dout <= 8'b00000000; //   51 :   0 - 0x0
      11'h34: dout <= 8'b00000000; //   52 :   0 - 0x0
      11'h35: dout <= 8'b00000000; //   53 :   0 - 0x0
      11'h36: dout <= 8'b00000000; //   54 :   0 - 0x0
      11'h37: dout <= 8'b00000000; //   55 :   0 - 0x0
      11'h38: dout <= 8'b00000000; //   56 :   0 - 0x0 -- Background 0x7
      11'h39: dout <= 8'b00000000; //   57 :   0 - 0x0
      11'h3A: dout <= 8'b00000000; //   58 :   0 - 0x0
      11'h3B: dout <= 8'b00000000; //   59 :   0 - 0x0
      11'h3C: dout <= 8'b00000000; //   60 :   0 - 0x0
      11'h3D: dout <= 8'b00000000; //   61 :   0 - 0x0
      11'h3E: dout <= 8'b00000000; //   62 :   0 - 0x0
      11'h3F: dout <= 8'b00000000; //   63 :   0 - 0x0
      11'h40: dout <= 8'b00000000; //   64 :   0 - 0x0 -- Background 0x8
      11'h41: dout <= 8'b00000000; //   65 :   0 - 0x0
      11'h42: dout <= 8'b00000000; //   66 :   0 - 0x0
      11'h43: dout <= 8'b00000000; //   67 :   0 - 0x0
      11'h44: dout <= 8'b00000000; //   68 :   0 - 0x0
      11'h45: dout <= 8'b00000000; //   69 :   0 - 0x0
      11'h46: dout <= 8'b00000000; //   70 :   0 - 0x0
      11'h47: dout <= 8'b00000000; //   71 :   0 - 0x0
      11'h48: dout <= 8'b00000000; //   72 :   0 - 0x0 -- Background 0x9
      11'h49: dout <= 8'b00000000; //   73 :   0 - 0x0
      11'h4A: dout <= 8'b00000000; //   74 :   0 - 0x0
      11'h4B: dout <= 8'b00000000; //   75 :   0 - 0x0
      11'h4C: dout <= 8'b00000000; //   76 :   0 - 0x0
      11'h4D: dout <= 8'b00000000; //   77 :   0 - 0x0
      11'h4E: dout <= 8'b00000000; //   78 :   0 - 0x0
      11'h4F: dout <= 8'b00000000; //   79 :   0 - 0x0
      11'h50: dout <= 8'b00000000; //   80 :   0 - 0x0 -- Background 0xa
      11'h51: dout <= 8'b00000000; //   81 :   0 - 0x0
      11'h52: dout <= 8'b00000000; //   82 :   0 - 0x0
      11'h53: dout <= 8'b00000000; //   83 :   0 - 0x0
      11'h54: dout <= 8'b00000000; //   84 :   0 - 0x0
      11'h55: dout <= 8'b00000000; //   85 :   0 - 0x0
      11'h56: dout <= 8'b00000000; //   86 :   0 - 0x0
      11'h57: dout <= 8'b00000000; //   87 :   0 - 0x0
      11'h58: dout <= 8'b00000000; //   88 :   0 - 0x0 -- Background 0xb
      11'h59: dout <= 8'b00000000; //   89 :   0 - 0x0
      11'h5A: dout <= 8'b00000000; //   90 :   0 - 0x0
      11'h5B: dout <= 8'b00000000; //   91 :   0 - 0x0
      11'h5C: dout <= 8'b00000000; //   92 :   0 - 0x0
      11'h5D: dout <= 8'b00000000; //   93 :   0 - 0x0
      11'h5E: dout <= 8'b00000000; //   94 :   0 - 0x0
      11'h5F: dout <= 8'b00000000; //   95 :   0 - 0x0
      11'h60: dout <= 8'b00000000; //   96 :   0 - 0x0 -- Background 0xc
      11'h61: dout <= 8'b00000000; //   97 :   0 - 0x0
      11'h62: dout <= 8'b00000000; //   98 :   0 - 0x0
      11'h63: dout <= 8'b00000000; //   99 :   0 - 0x0
      11'h64: dout <= 8'b00000000; //  100 :   0 - 0x0
      11'h65: dout <= 8'b00000000; //  101 :   0 - 0x0
      11'h66: dout <= 8'b00000000; //  102 :   0 - 0x0
      11'h67: dout <= 8'b00000000; //  103 :   0 - 0x0
      11'h68: dout <= 8'b00000000; //  104 :   0 - 0x0 -- Background 0xd
      11'h69: dout <= 8'b00000000; //  105 :   0 - 0x0
      11'h6A: dout <= 8'b00000000; //  106 :   0 - 0x0
      11'h6B: dout <= 8'b00000000; //  107 :   0 - 0x0
      11'h6C: dout <= 8'b00000000; //  108 :   0 - 0x0
      11'h6D: dout <= 8'b00000000; //  109 :   0 - 0x0
      11'h6E: dout <= 8'b00000000; //  110 :   0 - 0x0
      11'h6F: dout <= 8'b00000000; //  111 :   0 - 0x0
      11'h70: dout <= 8'b00000000; //  112 :   0 - 0x0 -- Background 0xe
      11'h71: dout <= 8'b00000000; //  113 :   0 - 0x0
      11'h72: dout <= 8'b00000000; //  114 :   0 - 0x0
      11'h73: dout <= 8'b00000000; //  115 :   0 - 0x0
      11'h74: dout <= 8'b00000000; //  116 :   0 - 0x0
      11'h75: dout <= 8'b00000000; //  117 :   0 - 0x0
      11'h76: dout <= 8'b00000000; //  118 :   0 - 0x0
      11'h77: dout <= 8'b00000000; //  119 :   0 - 0x0
      11'h78: dout <= 8'b00000000; //  120 :   0 - 0x0 -- Background 0xf
      11'h79: dout <= 8'b00000000; //  121 :   0 - 0x0
      11'h7A: dout <= 8'b00000000; //  122 :   0 - 0x0
      11'h7B: dout <= 8'b00000000; //  123 :   0 - 0x0
      11'h7C: dout <= 8'b00000000; //  124 :   0 - 0x0
      11'h7D: dout <= 8'b00000000; //  125 :   0 - 0x0
      11'h7E: dout <= 8'b00000000; //  126 :   0 - 0x0
      11'h7F: dout <= 8'b00000000; //  127 :   0 - 0x0
      11'h80: dout <= 8'b00000000; //  128 :   0 - 0x0 -- Background 0x10
      11'h81: dout <= 8'b00000000; //  129 :   0 - 0x0
      11'h82: dout <= 8'b00000000; //  130 :   0 - 0x0
      11'h83: dout <= 8'b00000000; //  131 :   0 - 0x0
      11'h84: dout <= 8'b00000000; //  132 :   0 - 0x0
      11'h85: dout <= 8'b00000000; //  133 :   0 - 0x0
      11'h86: dout <= 8'b00000000; //  134 :   0 - 0x0
      11'h87: dout <= 8'b00000000; //  135 :   0 - 0x0
      11'h88: dout <= 8'b00000000; //  136 :   0 - 0x0 -- Background 0x11
      11'h89: dout <= 8'b00000000; //  137 :   0 - 0x0
      11'h8A: dout <= 8'b00000000; //  138 :   0 - 0x0
      11'h8B: dout <= 8'b00000000; //  139 :   0 - 0x0
      11'h8C: dout <= 8'b00000000; //  140 :   0 - 0x0
      11'h8D: dout <= 8'b00000000; //  141 :   0 - 0x0
      11'h8E: dout <= 8'b00000000; //  142 :   0 - 0x0
      11'h8F: dout <= 8'b00000000; //  143 :   0 - 0x0
      11'h90: dout <= 8'b00000000; //  144 :   0 - 0x0 -- Background 0x12
      11'h91: dout <= 8'b00000000; //  145 :   0 - 0x0
      11'h92: dout <= 8'b00000000; //  146 :   0 - 0x0
      11'h93: dout <= 8'b00000000; //  147 :   0 - 0x0
      11'h94: dout <= 8'b00000000; //  148 :   0 - 0x0
      11'h95: dout <= 8'b00000000; //  149 :   0 - 0x0
      11'h96: dout <= 8'b00000000; //  150 :   0 - 0x0
      11'h97: dout <= 8'b00000000; //  151 :   0 - 0x0
      11'h98: dout <= 8'b00000000; //  152 :   0 - 0x0 -- Background 0x13
      11'h99: dout <= 8'b00000000; //  153 :   0 - 0x0
      11'h9A: dout <= 8'b00000000; //  154 :   0 - 0x0
      11'h9B: dout <= 8'b00000000; //  155 :   0 - 0x0
      11'h9C: dout <= 8'b00000000; //  156 :   0 - 0x0
      11'h9D: dout <= 8'b00000000; //  157 :   0 - 0x0
      11'h9E: dout <= 8'b00000000; //  158 :   0 - 0x0
      11'h9F: dout <= 8'b00000000; //  159 :   0 - 0x0
      11'hA0: dout <= 8'b00000000; //  160 :   0 - 0x0 -- Background 0x14
      11'hA1: dout <= 8'b00000000; //  161 :   0 - 0x0
      11'hA2: dout <= 8'b00000000; //  162 :   0 - 0x0
      11'hA3: dout <= 8'b00000000; //  163 :   0 - 0x0
      11'hA4: dout <= 8'b00000000; //  164 :   0 - 0x0
      11'hA5: dout <= 8'b00000000; //  165 :   0 - 0x0
      11'hA6: dout <= 8'b00000000; //  166 :   0 - 0x0
      11'hA7: dout <= 8'b00000000; //  167 :   0 - 0x0
      11'hA8: dout <= 8'b00000000; //  168 :   0 - 0x0 -- Background 0x15
      11'hA9: dout <= 8'b00000000; //  169 :   0 - 0x0
      11'hAA: dout <= 8'b00000000; //  170 :   0 - 0x0
      11'hAB: dout <= 8'b00000000; //  171 :   0 - 0x0
      11'hAC: dout <= 8'b00000000; //  172 :   0 - 0x0
      11'hAD: dout <= 8'b00000000; //  173 :   0 - 0x0
      11'hAE: dout <= 8'b00000000; //  174 :   0 - 0x0
      11'hAF: dout <= 8'b00000000; //  175 :   0 - 0x0
      11'hB0: dout <= 8'b00000000; //  176 :   0 - 0x0 -- Background 0x16
      11'hB1: dout <= 8'b00000000; //  177 :   0 - 0x0
      11'hB2: dout <= 8'b00000000; //  178 :   0 - 0x0
      11'hB3: dout <= 8'b00000000; //  179 :   0 - 0x0
      11'hB4: dout <= 8'b00000000; //  180 :   0 - 0x0
      11'hB5: dout <= 8'b00000000; //  181 :   0 - 0x0
      11'hB6: dout <= 8'b00000000; //  182 :   0 - 0x0
      11'hB7: dout <= 8'b00000000; //  183 :   0 - 0x0
      11'hB8: dout <= 8'b00000000; //  184 :   0 - 0x0 -- Background 0x17
      11'hB9: dout <= 8'b00000000; //  185 :   0 - 0x0
      11'hBA: dout <= 8'b00000000; //  186 :   0 - 0x0
      11'hBB: dout <= 8'b00000000; //  187 :   0 - 0x0
      11'hBC: dout <= 8'b00000000; //  188 :   0 - 0x0
      11'hBD: dout <= 8'b00000000; //  189 :   0 - 0x0
      11'hBE: dout <= 8'b00000000; //  190 :   0 - 0x0
      11'hBF: dout <= 8'b00000000; //  191 :   0 - 0x0
      11'hC0: dout <= 8'b00000000; //  192 :   0 - 0x0 -- Background 0x18
      11'hC1: dout <= 8'b00000000; //  193 :   0 - 0x0
      11'hC2: dout <= 8'b00000000; //  194 :   0 - 0x0
      11'hC3: dout <= 8'b00000000; //  195 :   0 - 0x0
      11'hC4: dout <= 8'b00000000; //  196 :   0 - 0x0
      11'hC5: dout <= 8'b00000000; //  197 :   0 - 0x0
      11'hC6: dout <= 8'b00000000; //  198 :   0 - 0x0
      11'hC7: dout <= 8'b00000000; //  199 :   0 - 0x0
      11'hC8: dout <= 8'b00000000; //  200 :   0 - 0x0 -- Background 0x19
      11'hC9: dout <= 8'b00000000; //  201 :   0 - 0x0
      11'hCA: dout <= 8'b00000000; //  202 :   0 - 0x0
      11'hCB: dout <= 8'b00000000; //  203 :   0 - 0x0
      11'hCC: dout <= 8'b00000000; //  204 :   0 - 0x0
      11'hCD: dout <= 8'b00000000; //  205 :   0 - 0x0
      11'hCE: dout <= 8'b00000000; //  206 :   0 - 0x0
      11'hCF: dout <= 8'b00000000; //  207 :   0 - 0x0
      11'hD0: dout <= 8'b00000000; //  208 :   0 - 0x0 -- Background 0x1a
      11'hD1: dout <= 8'b00000000; //  209 :   0 - 0x0
      11'hD2: dout <= 8'b00000000; //  210 :   0 - 0x0
      11'hD3: dout <= 8'b00000000; //  211 :   0 - 0x0
      11'hD4: dout <= 8'b00000000; //  212 :   0 - 0x0
      11'hD5: dout <= 8'b00000000; //  213 :   0 - 0x0
      11'hD6: dout <= 8'b00000000; //  214 :   0 - 0x0
      11'hD7: dout <= 8'b00000000; //  215 :   0 - 0x0
      11'hD8: dout <= 8'b00000000; //  216 :   0 - 0x0 -- Background 0x1b
      11'hD9: dout <= 8'b00000000; //  217 :   0 - 0x0
      11'hDA: dout <= 8'b00000000; //  218 :   0 - 0x0
      11'hDB: dout <= 8'b00000000; //  219 :   0 - 0x0
      11'hDC: dout <= 8'b00000000; //  220 :   0 - 0x0
      11'hDD: dout <= 8'b00000000; //  221 :   0 - 0x0
      11'hDE: dout <= 8'b00000000; //  222 :   0 - 0x0
      11'hDF: dout <= 8'b00000000; //  223 :   0 - 0x0
      11'hE0: dout <= 8'b00000000; //  224 :   0 - 0x0 -- Background 0x1c
      11'hE1: dout <= 8'b00000000; //  225 :   0 - 0x0
      11'hE2: dout <= 8'b00000000; //  226 :   0 - 0x0
      11'hE3: dout <= 8'b00000000; //  227 :   0 - 0x0
      11'hE4: dout <= 8'b00000000; //  228 :   0 - 0x0
      11'hE5: dout <= 8'b00000000; //  229 :   0 - 0x0
      11'hE6: dout <= 8'b00000000; //  230 :   0 - 0x0
      11'hE7: dout <= 8'b00000000; //  231 :   0 - 0x0
      11'hE8: dout <= 8'b00000000; //  232 :   0 - 0x0 -- Background 0x1d
      11'hE9: dout <= 8'b00000000; //  233 :   0 - 0x0
      11'hEA: dout <= 8'b00000000; //  234 :   0 - 0x0
      11'hEB: dout <= 8'b00000000; //  235 :   0 - 0x0
      11'hEC: dout <= 8'b00000000; //  236 :   0 - 0x0
      11'hED: dout <= 8'b00000000; //  237 :   0 - 0x0
      11'hEE: dout <= 8'b00000000; //  238 :   0 - 0x0
      11'hEF: dout <= 8'b00000000; //  239 :   0 - 0x0
      11'hF0: dout <= 8'b00000000; //  240 :   0 - 0x0 -- Background 0x1e
      11'hF1: dout <= 8'b00000000; //  241 :   0 - 0x0
      11'hF2: dout <= 8'b00000000; //  242 :   0 - 0x0
      11'hF3: dout <= 8'b00000000; //  243 :   0 - 0x0
      11'hF4: dout <= 8'b00000000; //  244 :   0 - 0x0
      11'hF5: dout <= 8'b00000000; //  245 :   0 - 0x0
      11'hF6: dout <= 8'b00000000; //  246 :   0 - 0x0
      11'hF7: dout <= 8'b00000000; //  247 :   0 - 0x0
      11'hF8: dout <= 8'b00000000; //  248 :   0 - 0x0 -- Background 0x1f
      11'hF9: dout <= 8'b00000000; //  249 :   0 - 0x0
      11'hFA: dout <= 8'b00000000; //  250 :   0 - 0x0
      11'hFB: dout <= 8'b00000000; //  251 :   0 - 0x0
      11'hFC: dout <= 8'b00000000; //  252 :   0 - 0x0
      11'hFD: dout <= 8'b00000000; //  253 :   0 - 0x0
      11'hFE: dout <= 8'b00000000; //  254 :   0 - 0x0
      11'hFF: dout <= 8'b00000000; //  255 :   0 - 0x0
      11'h100: dout <= 8'b00000000; //  256 :   0 - 0x0 -- Background 0x20
      11'h101: dout <= 8'b00000000; //  257 :   0 - 0x0
      11'h102: dout <= 8'b00000000; //  258 :   0 - 0x0
      11'h103: dout <= 8'b00000000; //  259 :   0 - 0x0
      11'h104: dout <= 8'b00000000; //  260 :   0 - 0x0
      11'h105: dout <= 8'b00000000; //  261 :   0 - 0x0
      11'h106: dout <= 8'b00000000; //  262 :   0 - 0x0
      11'h107: dout <= 8'b00000000; //  263 :   0 - 0x0
      11'h108: dout <= 8'b00000000; //  264 :   0 - 0x0 -- Background 0x21
      11'h109: dout <= 8'b00000000; //  265 :   0 - 0x0
      11'h10A: dout <= 8'b00000000; //  266 :   0 - 0x0
      11'h10B: dout <= 8'b00000000; //  267 :   0 - 0x0
      11'h10C: dout <= 8'b00000000; //  268 :   0 - 0x0
      11'h10D: dout <= 8'b00000000; //  269 :   0 - 0x0
      11'h10E: dout <= 8'b00000000; //  270 :   0 - 0x0
      11'h10F: dout <= 8'b00000000; //  271 :   0 - 0x0
      11'h110: dout <= 8'b00000000; //  272 :   0 - 0x0 -- Background 0x22
      11'h111: dout <= 8'b00000000; //  273 :   0 - 0x0
      11'h112: dout <= 8'b00000000; //  274 :   0 - 0x0
      11'h113: dout <= 8'b00000000; //  275 :   0 - 0x0
      11'h114: dout <= 8'b00000000; //  276 :   0 - 0x0
      11'h115: dout <= 8'b00000000; //  277 :   0 - 0x0
      11'h116: dout <= 8'b00000000; //  278 :   0 - 0x0
      11'h117: dout <= 8'b00000000; //  279 :   0 - 0x0
      11'h118: dout <= 8'b00000000; //  280 :   0 - 0x0 -- Background 0x23
      11'h119: dout <= 8'b00000000; //  281 :   0 - 0x0
      11'h11A: dout <= 8'b00000000; //  282 :   0 - 0x0
      11'h11B: dout <= 8'b00000000; //  283 :   0 - 0x0
      11'h11C: dout <= 8'b00000000; //  284 :   0 - 0x0
      11'h11D: dout <= 8'b00000000; //  285 :   0 - 0x0
      11'h11E: dout <= 8'b00000000; //  286 :   0 - 0x0
      11'h11F: dout <= 8'b00000000; //  287 :   0 - 0x0
      11'h120: dout <= 8'b00000000; //  288 :   0 - 0x0 -- Background 0x24
      11'h121: dout <= 8'b00000000; //  289 :   0 - 0x0
      11'h122: dout <= 8'b00000000; //  290 :   0 - 0x0
      11'h123: dout <= 8'b00000000; //  291 :   0 - 0x0
      11'h124: dout <= 8'b00000000; //  292 :   0 - 0x0
      11'h125: dout <= 8'b00000000; //  293 :   0 - 0x0
      11'h126: dout <= 8'b00000000; //  294 :   0 - 0x0
      11'h127: dout <= 8'b00000000; //  295 :   0 - 0x0
      11'h128: dout <= 8'b00000000; //  296 :   0 - 0x0 -- Background 0x25
      11'h129: dout <= 8'b00000000; //  297 :   0 - 0x0
      11'h12A: dout <= 8'b00000000; //  298 :   0 - 0x0
      11'h12B: dout <= 8'b00000000; //  299 :   0 - 0x0
      11'h12C: dout <= 8'b00000000; //  300 :   0 - 0x0
      11'h12D: dout <= 8'b00000000; //  301 :   0 - 0x0
      11'h12E: dout <= 8'b00000000; //  302 :   0 - 0x0
      11'h12F: dout <= 8'b00000000; //  303 :   0 - 0x0
      11'h130: dout <= 8'b00000000; //  304 :   0 - 0x0 -- Background 0x26
      11'h131: dout <= 8'b00000000; //  305 :   0 - 0x0
      11'h132: dout <= 8'b00000000; //  306 :   0 - 0x0
      11'h133: dout <= 8'b00000000; //  307 :   0 - 0x0
      11'h134: dout <= 8'b00000000; //  308 :   0 - 0x0
      11'h135: dout <= 8'b00000000; //  309 :   0 - 0x0
      11'h136: dout <= 8'b00000000; //  310 :   0 - 0x0
      11'h137: dout <= 8'b00000000; //  311 :   0 - 0x0
      11'h138: dout <= 8'b00000000; //  312 :   0 - 0x0 -- Background 0x27
      11'h139: dout <= 8'b00000000; //  313 :   0 - 0x0
      11'h13A: dout <= 8'b00000000; //  314 :   0 - 0x0
      11'h13B: dout <= 8'b00000000; //  315 :   0 - 0x0
      11'h13C: dout <= 8'b00000000; //  316 :   0 - 0x0
      11'h13D: dout <= 8'b00000000; //  317 :   0 - 0x0
      11'h13E: dout <= 8'b00000000; //  318 :   0 - 0x0
      11'h13F: dout <= 8'b00000000; //  319 :   0 - 0x0
      11'h140: dout <= 8'b00000000; //  320 :   0 - 0x0 -- Background 0x28
      11'h141: dout <= 8'b00000000; //  321 :   0 - 0x0
      11'h142: dout <= 8'b00000000; //  322 :   0 - 0x0
      11'h143: dout <= 8'b00000000; //  323 :   0 - 0x0
      11'h144: dout <= 8'b00000000; //  324 :   0 - 0x0
      11'h145: dout <= 8'b00000000; //  325 :   0 - 0x0
      11'h146: dout <= 8'b00000000; //  326 :   0 - 0x0
      11'h147: dout <= 8'b00000000; //  327 :   0 - 0x0
      11'h148: dout <= 8'b00000000; //  328 :   0 - 0x0 -- Background 0x29
      11'h149: dout <= 8'b00000000; //  329 :   0 - 0x0
      11'h14A: dout <= 8'b00000000; //  330 :   0 - 0x0
      11'h14B: dout <= 8'b00000000; //  331 :   0 - 0x0
      11'h14C: dout <= 8'b00000000; //  332 :   0 - 0x0
      11'h14D: dout <= 8'b00000000; //  333 :   0 - 0x0
      11'h14E: dout <= 8'b00000000; //  334 :   0 - 0x0
      11'h14F: dout <= 8'b00000000; //  335 :   0 - 0x0
      11'h150: dout <= 8'b00000000; //  336 :   0 - 0x0 -- Background 0x2a
      11'h151: dout <= 8'b00000000; //  337 :   0 - 0x0
      11'h152: dout <= 8'b00000000; //  338 :   0 - 0x0
      11'h153: dout <= 8'b00000000; //  339 :   0 - 0x0
      11'h154: dout <= 8'b00000000; //  340 :   0 - 0x0
      11'h155: dout <= 8'b00000000; //  341 :   0 - 0x0
      11'h156: dout <= 8'b00000000; //  342 :   0 - 0x0
      11'h157: dout <= 8'b00000000; //  343 :   0 - 0x0
      11'h158: dout <= 8'b00000000; //  344 :   0 - 0x0 -- Background 0x2b
      11'h159: dout <= 8'b00000000; //  345 :   0 - 0x0
      11'h15A: dout <= 8'b00000000; //  346 :   0 - 0x0
      11'h15B: dout <= 8'b00000000; //  347 :   0 - 0x0
      11'h15C: dout <= 8'b00000000; //  348 :   0 - 0x0
      11'h15D: dout <= 8'b00000000; //  349 :   0 - 0x0
      11'h15E: dout <= 8'b00000000; //  350 :   0 - 0x0
      11'h15F: dout <= 8'b00000000; //  351 :   0 - 0x0
      11'h160: dout <= 8'b00000000; //  352 :   0 - 0x0 -- Background 0x2c
      11'h161: dout <= 8'b00000000; //  353 :   0 - 0x0
      11'h162: dout <= 8'b00000000; //  354 :   0 - 0x0
      11'h163: dout <= 8'b00000000; //  355 :   0 - 0x0
      11'h164: dout <= 8'b00000000; //  356 :   0 - 0x0
      11'h165: dout <= 8'b00000000; //  357 :   0 - 0x0
      11'h166: dout <= 8'b00000000; //  358 :   0 - 0x0
      11'h167: dout <= 8'b00000000; //  359 :   0 - 0x0
      11'h168: dout <= 8'b00000000; //  360 :   0 - 0x0 -- Background 0x2d
      11'h169: dout <= 8'b00000000; //  361 :   0 - 0x0
      11'h16A: dout <= 8'b00000000; //  362 :   0 - 0x0
      11'h16B: dout <= 8'b00000000; //  363 :   0 - 0x0
      11'h16C: dout <= 8'b00000000; //  364 :   0 - 0x0
      11'h16D: dout <= 8'b00000000; //  365 :   0 - 0x0
      11'h16E: dout <= 8'b00000000; //  366 :   0 - 0x0
      11'h16F: dout <= 8'b00000000; //  367 :   0 - 0x0
      11'h170: dout <= 8'b00000000; //  368 :   0 - 0x0 -- Background 0x2e
      11'h171: dout <= 8'b00000000; //  369 :   0 - 0x0
      11'h172: dout <= 8'b00000000; //  370 :   0 - 0x0
      11'h173: dout <= 8'b00000000; //  371 :   0 - 0x0
      11'h174: dout <= 8'b00000000; //  372 :   0 - 0x0
      11'h175: dout <= 8'b00000000; //  373 :   0 - 0x0
      11'h176: dout <= 8'b00000000; //  374 :   0 - 0x0
      11'h177: dout <= 8'b00000000; //  375 :   0 - 0x0
      11'h178: dout <= 8'b00000000; //  376 :   0 - 0x0 -- Background 0x2f
      11'h179: dout <= 8'b00000000; //  377 :   0 - 0x0
      11'h17A: dout <= 8'b00000000; //  378 :   0 - 0x0
      11'h17B: dout <= 8'b00000000; //  379 :   0 - 0x0
      11'h17C: dout <= 8'b00000000; //  380 :   0 - 0x0
      11'h17D: dout <= 8'b00000000; //  381 :   0 - 0x0
      11'h17E: dout <= 8'b00000000; //  382 :   0 - 0x0
      11'h17F: dout <= 8'b00000000; //  383 :   0 - 0x0
      11'h180: dout <= 8'b00000000; //  384 :   0 - 0x0 -- Background 0x30
      11'h181: dout <= 8'b00000000; //  385 :   0 - 0x0
      11'h182: dout <= 8'b00000000; //  386 :   0 - 0x0
      11'h183: dout <= 8'b00000000; //  387 :   0 - 0x0
      11'h184: dout <= 8'b00000000; //  388 :   0 - 0x0
      11'h185: dout <= 8'b00000000; //  389 :   0 - 0x0
      11'h186: dout <= 8'b00000000; //  390 :   0 - 0x0
      11'h187: dout <= 8'b00000000; //  391 :   0 - 0x0
      11'h188: dout <= 8'b00000000; //  392 :   0 - 0x0 -- Background 0x31
      11'h189: dout <= 8'b00000000; //  393 :   0 - 0x0
      11'h18A: dout <= 8'b00000000; //  394 :   0 - 0x0
      11'h18B: dout <= 8'b00000000; //  395 :   0 - 0x0
      11'h18C: dout <= 8'b00000000; //  396 :   0 - 0x0
      11'h18D: dout <= 8'b00000000; //  397 :   0 - 0x0
      11'h18E: dout <= 8'b00000000; //  398 :   0 - 0x0
      11'h18F: dout <= 8'b00000000; //  399 :   0 - 0x0
      11'h190: dout <= 8'b00000000; //  400 :   0 - 0x0 -- Background 0x32
      11'h191: dout <= 8'b00000000; //  401 :   0 - 0x0
      11'h192: dout <= 8'b00000000; //  402 :   0 - 0x0
      11'h193: dout <= 8'b00000000; //  403 :   0 - 0x0
      11'h194: dout <= 8'b00000000; //  404 :   0 - 0x0
      11'h195: dout <= 8'b00000000; //  405 :   0 - 0x0
      11'h196: dout <= 8'b00000000; //  406 :   0 - 0x0
      11'h197: dout <= 8'b00000000; //  407 :   0 - 0x0
      11'h198: dout <= 8'b00000000; //  408 :   0 - 0x0 -- Background 0x33
      11'h199: dout <= 8'b00000000; //  409 :   0 - 0x0
      11'h19A: dout <= 8'b00000000; //  410 :   0 - 0x0
      11'h19B: dout <= 8'b00000000; //  411 :   0 - 0x0
      11'h19C: dout <= 8'b00000000; //  412 :   0 - 0x0
      11'h19D: dout <= 8'b00000000; //  413 :   0 - 0x0
      11'h19E: dout <= 8'b00000000; //  414 :   0 - 0x0
      11'h19F: dout <= 8'b00000000; //  415 :   0 - 0x0
      11'h1A0: dout <= 8'b00000000; //  416 :   0 - 0x0 -- Background 0x34
      11'h1A1: dout <= 8'b00000000; //  417 :   0 - 0x0
      11'h1A2: dout <= 8'b00000000; //  418 :   0 - 0x0
      11'h1A3: dout <= 8'b00000000; //  419 :   0 - 0x0
      11'h1A4: dout <= 8'b00000000; //  420 :   0 - 0x0
      11'h1A5: dout <= 8'b00000000; //  421 :   0 - 0x0
      11'h1A6: dout <= 8'b00000000; //  422 :   0 - 0x0
      11'h1A7: dout <= 8'b00000000; //  423 :   0 - 0x0
      11'h1A8: dout <= 8'b00000000; //  424 :   0 - 0x0 -- Background 0x35
      11'h1A9: dout <= 8'b00000000; //  425 :   0 - 0x0
      11'h1AA: dout <= 8'b00000000; //  426 :   0 - 0x0
      11'h1AB: dout <= 8'b00000000; //  427 :   0 - 0x0
      11'h1AC: dout <= 8'b00000000; //  428 :   0 - 0x0
      11'h1AD: dout <= 8'b00000000; //  429 :   0 - 0x0
      11'h1AE: dout <= 8'b00000000; //  430 :   0 - 0x0
      11'h1AF: dout <= 8'b00000000; //  431 :   0 - 0x0
      11'h1B0: dout <= 8'b00000000; //  432 :   0 - 0x0 -- Background 0x36
      11'h1B1: dout <= 8'b00000000; //  433 :   0 - 0x0
      11'h1B2: dout <= 8'b00000000; //  434 :   0 - 0x0
      11'h1B3: dout <= 8'b00000000; //  435 :   0 - 0x0
      11'h1B4: dout <= 8'b00000000; //  436 :   0 - 0x0
      11'h1B5: dout <= 8'b00000000; //  437 :   0 - 0x0
      11'h1B6: dout <= 8'b00000000; //  438 :   0 - 0x0
      11'h1B7: dout <= 8'b00000000; //  439 :   0 - 0x0
      11'h1B8: dout <= 8'b00000000; //  440 :   0 - 0x0 -- Background 0x37
      11'h1B9: dout <= 8'b00000000; //  441 :   0 - 0x0
      11'h1BA: dout <= 8'b00000000; //  442 :   0 - 0x0
      11'h1BB: dout <= 8'b00000000; //  443 :   0 - 0x0
      11'h1BC: dout <= 8'b00000000; //  444 :   0 - 0x0
      11'h1BD: dout <= 8'b00000000; //  445 :   0 - 0x0
      11'h1BE: dout <= 8'b00000000; //  446 :   0 - 0x0
      11'h1BF: dout <= 8'b00000000; //  447 :   0 - 0x0
      11'h1C0: dout <= 8'b00000000; //  448 :   0 - 0x0 -- Background 0x38
      11'h1C1: dout <= 8'b00000000; //  449 :   0 - 0x0
      11'h1C2: dout <= 8'b00000000; //  450 :   0 - 0x0
      11'h1C3: dout <= 8'b00000000; //  451 :   0 - 0x0
      11'h1C4: dout <= 8'b00000000; //  452 :   0 - 0x0
      11'h1C5: dout <= 8'b00000000; //  453 :   0 - 0x0
      11'h1C6: dout <= 8'b00000000; //  454 :   0 - 0x0
      11'h1C7: dout <= 8'b00000000; //  455 :   0 - 0x0
      11'h1C8: dout <= 8'b00000000; //  456 :   0 - 0x0 -- Background 0x39
      11'h1C9: dout <= 8'b00000000; //  457 :   0 - 0x0
      11'h1CA: dout <= 8'b00000000; //  458 :   0 - 0x0
      11'h1CB: dout <= 8'b00000000; //  459 :   0 - 0x0
      11'h1CC: dout <= 8'b00000000; //  460 :   0 - 0x0
      11'h1CD: dout <= 8'b00000000; //  461 :   0 - 0x0
      11'h1CE: dout <= 8'b00000000; //  462 :   0 - 0x0
      11'h1CF: dout <= 8'b00000000; //  463 :   0 - 0x0
      11'h1D0: dout <= 8'b00000000; //  464 :   0 - 0x0 -- Background 0x3a
      11'h1D1: dout <= 8'b00000000; //  465 :   0 - 0x0
      11'h1D2: dout <= 8'b00000000; //  466 :   0 - 0x0
      11'h1D3: dout <= 8'b00000000; //  467 :   0 - 0x0
      11'h1D4: dout <= 8'b00000000; //  468 :   0 - 0x0
      11'h1D5: dout <= 8'b00000000; //  469 :   0 - 0x0
      11'h1D6: dout <= 8'b00000000; //  470 :   0 - 0x0
      11'h1D7: dout <= 8'b00000000; //  471 :   0 - 0x0
      11'h1D8: dout <= 8'b00000000; //  472 :   0 - 0x0 -- Background 0x3b
      11'h1D9: dout <= 8'b00000000; //  473 :   0 - 0x0
      11'h1DA: dout <= 8'b00000000; //  474 :   0 - 0x0
      11'h1DB: dout <= 8'b00000000; //  475 :   0 - 0x0
      11'h1DC: dout <= 8'b00000000; //  476 :   0 - 0x0
      11'h1DD: dout <= 8'b00000000; //  477 :   0 - 0x0
      11'h1DE: dout <= 8'b00000000; //  478 :   0 - 0x0
      11'h1DF: dout <= 8'b00000000; //  479 :   0 - 0x0
      11'h1E0: dout <= 8'b00000000; //  480 :   0 - 0x0 -- Background 0x3c
      11'h1E1: dout <= 8'b00000000; //  481 :   0 - 0x0
      11'h1E2: dout <= 8'b00000000; //  482 :   0 - 0x0
      11'h1E3: dout <= 8'b00000000; //  483 :   0 - 0x0
      11'h1E4: dout <= 8'b00000000; //  484 :   0 - 0x0
      11'h1E5: dout <= 8'b00000000; //  485 :   0 - 0x0
      11'h1E6: dout <= 8'b00000000; //  486 :   0 - 0x0
      11'h1E7: dout <= 8'b00000000; //  487 :   0 - 0x0
      11'h1E8: dout <= 8'b00000000; //  488 :   0 - 0x0 -- Background 0x3d
      11'h1E9: dout <= 8'b00000000; //  489 :   0 - 0x0
      11'h1EA: dout <= 8'b00000000; //  490 :   0 - 0x0
      11'h1EB: dout <= 8'b00000000; //  491 :   0 - 0x0
      11'h1EC: dout <= 8'b00000000; //  492 :   0 - 0x0
      11'h1ED: dout <= 8'b00000000; //  493 :   0 - 0x0
      11'h1EE: dout <= 8'b00000000; //  494 :   0 - 0x0
      11'h1EF: dout <= 8'b00000000; //  495 :   0 - 0x0
      11'h1F0: dout <= 8'b00000000; //  496 :   0 - 0x0 -- Background 0x3e
      11'h1F1: dout <= 8'b00000000; //  497 :   0 - 0x0
      11'h1F2: dout <= 8'b00000000; //  498 :   0 - 0x0
      11'h1F3: dout <= 8'b00000000; //  499 :   0 - 0x0
      11'h1F4: dout <= 8'b00000000; //  500 :   0 - 0x0
      11'h1F5: dout <= 8'b00000000; //  501 :   0 - 0x0
      11'h1F6: dout <= 8'b00000000; //  502 :   0 - 0x0
      11'h1F7: dout <= 8'b00000000; //  503 :   0 - 0x0
      11'h1F8: dout <= 8'b10000001; //  504 : 129 - 0x81 -- Background 0x3f
      11'h1F9: dout <= 8'b11111111; //  505 : 255 - 0xff
      11'h1FA: dout <= 8'b10000001; //  506 : 129 - 0x81
      11'h1FB: dout <= 8'b10000001; //  507 : 129 - 0x81
      11'h1FC: dout <= 8'b10000001; //  508 : 129 - 0x81
      11'h1FD: dout <= 8'b11111111; //  509 : 255 - 0xff
      11'h1FE: dout <= 8'b10000001; //  510 : 129 - 0x81
      11'h1FF: dout <= 8'b10000001; //  511 : 129 - 0x81
      11'h200: dout <= 8'b10000001; //  512 : 129 - 0x81 -- Background 0x40
      11'h201: dout <= 8'b11111111; //  513 : 255 - 0xff
      11'h202: dout <= 8'b10000001; //  514 : 129 - 0x81
      11'h203: dout <= 8'b10000001; //  515 : 129 - 0x81
      11'h204: dout <= 8'b10000001; //  516 : 129 - 0x81
      11'h205: dout <= 8'b11111111; //  517 : 255 - 0xff
      11'h206: dout <= 8'b10000001; //  518 : 129 - 0x81
      11'h207: dout <= 8'b00000000; //  519 :   0 - 0x0
      11'h208: dout <= 8'b10000001; //  520 : 129 - 0x81 -- Background 0x41
      11'h209: dout <= 8'b11111111; //  521 : 255 - 0xff
      11'h20A: dout <= 8'b10000001; //  522 : 129 - 0x81
      11'h20B: dout <= 8'b10000001; //  523 : 129 - 0x81
      11'h20C: dout <= 8'b10000001; //  524 : 129 - 0x81
      11'h20D: dout <= 8'b00000000; //  525 :   0 - 0x0
      11'h20E: dout <= 8'b00000000; //  526 :   0 - 0x0
      11'h20F: dout <= 8'b00000000; //  527 :   0 - 0x0
      11'h210: dout <= 8'b10000001; //  528 : 129 - 0x81 -- Background 0x42
      11'h211: dout <= 8'b11111111; //  529 : 255 - 0xff
      11'h212: dout <= 8'b10000001; //  530 : 129 - 0x81
      11'h213: dout <= 8'b10000001; //  531 : 129 - 0x81
      11'h214: dout <= 8'b00000000; //  532 :   0 - 0x0
      11'h215: dout <= 8'b00000000; //  533 :   0 - 0x0
      11'h216: dout <= 8'b00000000; //  534 :   0 - 0x0
      11'h217: dout <= 8'b00000000; //  535 :   0 - 0x0
      11'h218: dout <= 8'b10000001; //  536 : 129 - 0x81 -- Background 0x43
      11'h219: dout <= 8'b11111111; //  537 : 255 - 0xff
      11'h21A: dout <= 8'b10000001; //  538 : 129 - 0x81
      11'h21B: dout <= 8'b00000000; //  539 :   0 - 0x0
      11'h21C: dout <= 8'b00000000; //  540 :   0 - 0x0
      11'h21D: dout <= 8'b00000000; //  541 :   0 - 0x0
      11'h21E: dout <= 8'b00000000; //  542 :   0 - 0x0
      11'h21F: dout <= 8'b00000000; //  543 :   0 - 0x0
      11'h220: dout <= 8'b10000001; //  544 : 129 - 0x81 -- Background 0x44
      11'h221: dout <= 8'b11111111; //  545 : 255 - 0xff
      11'h222: dout <= 8'b00000000; //  546 :   0 - 0x0
      11'h223: dout <= 8'b00000000; //  547 :   0 - 0x0
      11'h224: dout <= 8'b00000000; //  548 :   0 - 0x0
      11'h225: dout <= 8'b00000000; //  549 :   0 - 0x0
      11'h226: dout <= 8'b00000000; //  550 :   0 - 0x0
      11'h227: dout <= 8'b00000000; //  551 :   0 - 0x0
      11'h228: dout <= 8'b10000001; //  552 : 129 - 0x81 -- Background 0x45
      11'h229: dout <= 8'b00000000; //  553 :   0 - 0x0
      11'h22A: dout <= 8'b00000000; //  554 :   0 - 0x0
      11'h22B: dout <= 8'b00000000; //  555 :   0 - 0x0
      11'h22C: dout <= 8'b00000000; //  556 :   0 - 0x0
      11'h22D: dout <= 8'b00000000; //  557 :   0 - 0x0
      11'h22E: dout <= 8'b00000000; //  558 :   0 - 0x0
      11'h22F: dout <= 8'b00000000; //  559 :   0 - 0x0
      11'h230: dout <= 8'b00000000; //  560 :   0 - 0x0 -- Background 0x46
      11'h231: dout <= 8'b00000000; //  561 :   0 - 0x0
      11'h232: dout <= 8'b00000000; //  562 :   0 - 0x0
      11'h233: dout <= 8'b00000000; //  563 :   0 - 0x0
      11'h234: dout <= 8'b00000000; //  564 :   0 - 0x0
      11'h235: dout <= 8'b00000000; //  565 :   0 - 0x0
      11'h236: dout <= 8'b00000000; //  566 :   0 - 0x0
      11'h237: dout <= 8'b10000001; //  567 : 129 - 0x81
      11'h238: dout <= 8'b00000000; //  568 :   0 - 0x0 -- Background 0x47
      11'h239: dout <= 8'b00000000; //  569 :   0 - 0x0
      11'h23A: dout <= 8'b00000000; //  570 :   0 - 0x0
      11'h23B: dout <= 8'b00000000; //  571 :   0 - 0x0
      11'h23C: dout <= 8'b00000000; //  572 :   0 - 0x0
      11'h23D: dout <= 8'b00000000; //  573 :   0 - 0x0
      11'h23E: dout <= 8'b10000001; //  574 : 129 - 0x81
      11'h23F: dout <= 8'b10000001; //  575 : 129 - 0x81
      11'h240: dout <= 8'b00000000; //  576 :   0 - 0x0 -- Background 0x48
      11'h241: dout <= 8'b00000000; //  577 :   0 - 0x0
      11'h242: dout <= 8'b00000000; //  578 :   0 - 0x0
      11'h243: dout <= 8'b00000000; //  579 :   0 - 0x0
      11'h244: dout <= 8'b00000000; //  580 :   0 - 0x0
      11'h245: dout <= 8'b11111111; //  581 : 255 - 0xff
      11'h246: dout <= 8'b10000001; //  582 : 129 - 0x81
      11'h247: dout <= 8'b10000001; //  583 : 129 - 0x81
      11'h248: dout <= 8'b00000000; //  584 :   0 - 0x0 -- Background 0x49
      11'h249: dout <= 8'b00000000; //  585 :   0 - 0x0
      11'h24A: dout <= 8'b00000000; //  586 :   0 - 0x0
      11'h24B: dout <= 8'b00000000; //  587 :   0 - 0x0
      11'h24C: dout <= 8'b10000001; //  588 : 129 - 0x81
      11'h24D: dout <= 8'b11111111; //  589 : 255 - 0xff
      11'h24E: dout <= 8'b10000001; //  590 : 129 - 0x81
      11'h24F: dout <= 8'b10000001; //  591 : 129 - 0x81
      11'h250: dout <= 8'b00000000; //  592 :   0 - 0x0 -- Background 0x4a
      11'h251: dout <= 8'b00000000; //  593 :   0 - 0x0
      11'h252: dout <= 8'b00000000; //  594 :   0 - 0x0
      11'h253: dout <= 8'b10000001; //  595 : 129 - 0x81
      11'h254: dout <= 8'b10000001; //  596 : 129 - 0x81
      11'h255: dout <= 8'b11111111; //  597 : 255 - 0xff
      11'h256: dout <= 8'b10000001; //  598 : 129 - 0x81
      11'h257: dout <= 8'b10000001; //  599 : 129 - 0x81
      11'h258: dout <= 8'b00000000; //  600 :   0 - 0x0 -- Background 0x4b
      11'h259: dout <= 8'b00000000; //  601 :   0 - 0x0
      11'h25A: dout <= 8'b10000001; //  602 : 129 - 0x81
      11'h25B: dout <= 8'b10000001; //  603 : 129 - 0x81
      11'h25C: dout <= 8'b10000001; //  604 : 129 - 0x81
      11'h25D: dout <= 8'b11111111; //  605 : 255 - 0xff
      11'h25E: dout <= 8'b10000001; //  606 : 129 - 0x81
      11'h25F: dout <= 8'b10000001; //  607 : 129 - 0x81
      11'h260: dout <= 8'b11111111; //  608 : 255 - 0xff -- Background 0x4c
      11'h261: dout <= 8'b01111111; //  609 : 127 - 0x7f
      11'h262: dout <= 8'b01111111; //  610 : 127 - 0x7f
      11'h263: dout <= 8'b01111111; //  611 : 127 - 0x7f
      11'h264: dout <= 8'b01111111; //  612 : 127 - 0x7f
      11'h265: dout <= 8'b01111111; //  613 : 127 - 0x7f
      11'h266: dout <= 8'b01111111; //  614 : 127 - 0x7f
      11'h267: dout <= 8'b01111111; //  615 : 127 - 0x7f
      11'h268: dout <= 8'b01111111; //  616 : 127 - 0x7f -- Background 0x4d
      11'h269: dout <= 8'b01111111; //  617 : 127 - 0x7f
      11'h26A: dout <= 8'b01111111; //  618 : 127 - 0x7f
      11'h26B: dout <= 8'b01111111; //  619 : 127 - 0x7f
      11'h26C: dout <= 8'b01110010; //  620 : 114 - 0x72
      11'h26D: dout <= 8'b01111111; //  621 : 127 - 0x7f
      11'h26E: dout <= 8'b01111111; //  622 : 127 - 0x7f
      11'h26F: dout <= 8'b11111111; //  623 : 255 - 0xff
      11'h270: dout <= 8'b11111111; //  624 : 255 - 0xff -- Background 0x4e
      11'h271: dout <= 8'b11111110; //  625 : 254 - 0xfe
      11'h272: dout <= 8'b11111110; //  626 : 254 - 0xfe
      11'h273: dout <= 8'b11111110; //  627 : 254 - 0xfe
      11'h274: dout <= 8'b11111110; //  628 : 254 - 0xfe
      11'h275: dout <= 8'b11111110; //  629 : 254 - 0xfe
      11'h276: dout <= 8'b11111110; //  630 : 254 - 0xfe
      11'h277: dout <= 8'b11111110; //  631 : 254 - 0xfe
      11'h278: dout <= 8'b11111110; //  632 : 254 - 0xfe -- Background 0x4f
      11'h279: dout <= 8'b11111110; //  633 : 254 - 0xfe
      11'h27A: dout <= 8'b11111110; //  634 : 254 - 0xfe
      11'h27B: dout <= 8'b11111110; //  635 : 254 - 0xfe
      11'h27C: dout <= 8'b01001010; //  636 :  74 - 0x4a
      11'h27D: dout <= 8'b11111110; //  637 : 254 - 0xfe
      11'h27E: dout <= 8'b11111110; //  638 : 254 - 0xfe
      11'h27F: dout <= 8'b11111111; //  639 : 255 - 0xff
      11'h280: dout <= 8'b00000101; //  640 :   5 - 0x5 -- Background 0x50
      11'h281: dout <= 8'b00001111; //  641 :  15 - 0xf
      11'h282: dout <= 8'b00001011; //  642 :  11 - 0xb
      11'h283: dout <= 8'b00011011; //  643 :  27 - 0x1b
      11'h284: dout <= 8'b00010011; //  644 :  19 - 0x13
      11'h285: dout <= 8'b00010011; //  645 :  19 - 0x13
      11'h286: dout <= 8'b00010011; //  646 :  19 - 0x13
      11'h287: dout <= 8'b00010011; //  647 :  19 - 0x13
      11'h288: dout <= 8'b00010011; //  648 :  19 - 0x13 -- Background 0x51
      11'h289: dout <= 8'b00010011; //  649 :  19 - 0x13
      11'h28A: dout <= 8'b00010011; //  650 :  19 - 0x13
      11'h28B: dout <= 8'b00010011; //  651 :  19 - 0x13
      11'h28C: dout <= 8'b00011011; //  652 :  27 - 0x1b
      11'h28D: dout <= 8'b00001011; //  653 :  11 - 0xb
      11'h28E: dout <= 8'b00001111; //  654 :  15 - 0xf
      11'h28F: dout <= 8'b00000101; //  655 :   5 - 0x5
      11'h290: dout <= 8'b00000101; //  656 :   5 - 0x5 -- Background 0x52
      11'h291: dout <= 8'b00001111; //  657 :  15 - 0xf
      11'h292: dout <= 8'b00001011; //  658 :  11 - 0xb
      11'h293: dout <= 8'b00011011; //  659 :  27 - 0x1b
      11'h294: dout <= 8'b00010011; //  660 :  19 - 0x13
      11'h295: dout <= 8'b00010011; //  661 :  19 - 0x13
      11'h296: dout <= 8'b00010011; //  662 :  19 - 0x13
      11'h297: dout <= 8'b00010011; //  663 :  19 - 0x13
      11'h298: dout <= 8'b00010011; //  664 :  19 - 0x13 -- Background 0x53
      11'h299: dout <= 8'b00010011; //  665 :  19 - 0x13
      11'h29A: dout <= 8'b00010011; //  666 :  19 - 0x13
      11'h29B: dout <= 8'b00010011; //  667 :  19 - 0x13
      11'h29C: dout <= 8'b00011011; //  668 :  27 - 0x1b
      11'h29D: dout <= 8'b00001011; //  669 :  11 - 0xb
      11'h29E: dout <= 8'b00001111; //  670 :  15 - 0xf
      11'h29F: dout <= 8'b00000101; //  671 :   5 - 0x5
      11'h2A0: dout <= 8'b10100000; //  672 : 160 - 0xa0 -- Background 0x54
      11'h2A1: dout <= 8'b11110001; //  673 : 241 - 0xf1
      11'h2A2: dout <= 8'b11010001; //  674 : 209 - 0xd1
      11'h2A3: dout <= 8'b11011011; //  675 : 219 - 0xdb
      11'h2A4: dout <= 8'b11001010; //  676 : 202 - 0xca
      11'h2A5: dout <= 8'b11001010; //  677 : 202 - 0xca
      11'h2A6: dout <= 8'b11001010; //  678 : 202 - 0xca
      11'h2A7: dout <= 8'b11001010; //  679 : 202 - 0xca
      11'h2A8: dout <= 8'b11001010; //  680 : 202 - 0xca -- Background 0x55
      11'h2A9: dout <= 8'b11001010; //  681 : 202 - 0xca
      11'h2AA: dout <= 8'b11001010; //  682 : 202 - 0xca
      11'h2AB: dout <= 8'b11001010; //  683 : 202 - 0xca
      11'h2AC: dout <= 8'b11011011; //  684 : 219 - 0xdb
      11'h2AD: dout <= 8'b11010001; //  685 : 209 - 0xd1
      11'h2AE: dout <= 8'b11110001; //  686 : 241 - 0xf1
      11'h2AF: dout <= 8'b10100000; //  687 : 160 - 0xa0
      11'h2B0: dout <= 8'b10100000; //  688 : 160 - 0xa0 -- Background 0x56
      11'h2B1: dout <= 8'b11110001; //  689 : 241 - 0xf1
      11'h2B2: dout <= 8'b11010001; //  690 : 209 - 0xd1
      11'h2B3: dout <= 8'b11011011; //  691 : 219 - 0xdb
      11'h2B4: dout <= 8'b11001010; //  692 : 202 - 0xca
      11'h2B5: dout <= 8'b11001010; //  693 : 202 - 0xca
      11'h2B6: dout <= 8'b11001010; //  694 : 202 - 0xca
      11'h2B7: dout <= 8'b11001010; //  695 : 202 - 0xca
      11'h2B8: dout <= 8'b11001010; //  696 : 202 - 0xca -- Background 0x57
      11'h2B9: dout <= 8'b11001010; //  697 : 202 - 0xca
      11'h2BA: dout <= 8'b11001010; //  698 : 202 - 0xca
      11'h2BB: dout <= 8'b11001010; //  699 : 202 - 0xca
      11'h2BC: dout <= 8'b11011011; //  700 : 219 - 0xdb
      11'h2BD: dout <= 8'b11010001; //  701 : 209 - 0xd1
      11'h2BE: dout <= 8'b11110000; //  702 : 240 - 0xf0
      11'h2BF: dout <= 8'b10100000; //  703 : 160 - 0xa0
      11'h2C0: dout <= 8'b10110100; //  704 : 180 - 0xb4 -- Background 0x58
      11'h2C1: dout <= 8'b11111110; //  705 : 254 - 0xfe
      11'h2C2: dout <= 8'b01111010; //  706 : 122 - 0x7a
      11'h2C3: dout <= 8'b01111011; //  707 : 123 - 0x7b
      11'h2C4: dout <= 8'b01111001; //  708 : 121 - 0x79
      11'h2C5: dout <= 8'b01111001; //  709 : 121 - 0x79
      11'h2C6: dout <= 8'b01111001; //  710 : 121 - 0x79
      11'h2C7: dout <= 8'b01111001; //  711 : 121 - 0x79
      11'h2C8: dout <= 8'b01111001; //  712 : 121 - 0x79 -- Background 0x59
      11'h2C9: dout <= 8'b01111001; //  713 : 121 - 0x79
      11'h2CA: dout <= 8'b01111001; //  714 : 121 - 0x79
      11'h2CB: dout <= 8'b01111001; //  715 : 121 - 0x79
      11'h2CC: dout <= 8'b01111011; //  716 : 123 - 0x7b
      11'h2CD: dout <= 8'b01111010; //  717 : 122 - 0x7a
      11'h2CE: dout <= 8'b11111110; //  718 : 254 - 0xfe
      11'h2CF: dout <= 8'b10110100; //  719 : 180 - 0xb4
      11'h2D0: dout <= 8'b10110100; //  720 : 180 - 0xb4 -- Background 0x5a
      11'h2D1: dout <= 8'b11111110; //  721 : 254 - 0xfe
      11'h2D2: dout <= 8'b01111010; //  722 : 122 - 0x7a
      11'h2D3: dout <= 8'b01111011; //  723 : 123 - 0x7b
      11'h2D4: dout <= 8'b01111001; //  724 : 121 - 0x79
      11'h2D5: dout <= 8'b01111001; //  725 : 121 - 0x79
      11'h2D6: dout <= 8'b01111001; //  726 : 121 - 0x79
      11'h2D7: dout <= 8'b01111001; //  727 : 121 - 0x79
      11'h2D8: dout <= 8'b01111001; //  728 : 121 - 0x79 -- Background 0x5b
      11'h2D9: dout <= 8'b01111001; //  729 : 121 - 0x79
      11'h2DA: dout <= 8'b01111001; //  730 : 121 - 0x79
      11'h2DB: dout <= 8'b01111001; //  731 : 121 - 0x79
      11'h2DC: dout <= 8'b01111011; //  732 : 123 - 0x7b
      11'h2DD: dout <= 8'b01111010; //  733 : 122 - 0x7a
      11'h2DE: dout <= 8'b11111110; //  734 : 254 - 0xfe
      11'h2DF: dout <= 8'b10110100; //  735 : 180 - 0xb4
      11'h2E0: dout <= 8'b01111111; //  736 : 127 - 0x7f -- Background 0x5c
      11'h2E1: dout <= 8'b10111111; //  737 : 191 - 0xbf
      11'h2E2: dout <= 8'b11111111; //  738 : 255 - 0xff
      11'h2E3: dout <= 8'b10110010; //  739 : 178 - 0xb2
      11'h2E4: dout <= 8'b10110001; //  740 : 177 - 0xb1
      11'h2E5: dout <= 8'b11111111; //  741 : 255 - 0xff
      11'h2E6: dout <= 8'b10111111; //  742 : 191 - 0xbf
      11'h2E7: dout <= 8'b01111111; //  743 : 127 - 0x7f
      11'h2E8: dout <= 8'b11111110; //  744 : 254 - 0xfe -- Background 0x5d
      11'h2E9: dout <= 8'b11111101; //  745 : 253 - 0xfd
      11'h2EA: dout <= 8'b11111111; //  746 : 255 - 0xff
      11'h2EB: dout <= 8'b11001101; //  747 : 205 - 0xcd
      11'h2EC: dout <= 8'b01101101; //  748 : 109 - 0x6d
      11'h2ED: dout <= 8'b11111111; //  749 : 255 - 0xff
      11'h2EE: dout <= 8'b11111101; //  750 : 253 - 0xfd
      11'h2EF: dout <= 8'b11111110; //  751 : 254 - 0xfe
      11'h2F0: dout <= 8'b11111111; //  752 : 255 - 0xff -- Background 0x5e
      11'h2F1: dout <= 8'b11111111; //  753 : 255 - 0xff
      11'h2F2: dout <= 8'b10101110; //  754 : 174 - 0xae
      11'h2F3: dout <= 8'b11111110; //  755 : 254 - 0xfe
      11'h2F4: dout <= 8'b11111111; //  756 : 255 - 0xff
      11'h2F5: dout <= 8'b00001111; //  757 :  15 - 0xf
      11'h2F6: dout <= 8'b00000111; //  758 :   7 - 0x7
      11'h2F7: dout <= 8'b00000011; //  759 :   3 - 0x3
      11'h2F8: dout <= 8'b11111111; //  760 : 255 - 0xff -- Background 0x5f
      11'h2F9: dout <= 8'b11111111; //  761 : 255 - 0xff
      11'h2FA: dout <= 8'b01110101; //  762 : 117 - 0x75
      11'h2FB: dout <= 8'b01111111; //  763 : 127 - 0x7f
      11'h2FC: dout <= 8'b11111111; //  764 : 255 - 0xff
      11'h2FD: dout <= 8'b11110000; //  765 : 240 - 0xf0
      11'h2FE: dout <= 8'b11100000; //  766 : 224 - 0xe0
      11'h2FF: dout <= 8'b11000000; //  767 : 192 - 0xc0
      11'h300: dout <= 8'b00000011; //  768 :   3 - 0x3 -- Background 0x60
      11'h301: dout <= 8'b00000111; //  769 :   7 - 0x7
      11'h302: dout <= 8'b00001111; //  770 :  15 - 0xf
      11'h303: dout <= 8'b11111111; //  771 : 255 - 0xff
      11'h304: dout <= 8'b11111110; //  772 : 254 - 0xfe
      11'h305: dout <= 8'b10101110; //  773 : 174 - 0xae
      11'h306: dout <= 8'b11111111; //  774 : 255 - 0xff
      11'h307: dout <= 8'b11111111; //  775 : 255 - 0xff
      11'h308: dout <= 8'b11000000; //  776 : 192 - 0xc0 -- Background 0x61
      11'h309: dout <= 8'b11100000; //  777 : 224 - 0xe0
      11'h30A: dout <= 8'b11110000; //  778 : 240 - 0xf0
      11'h30B: dout <= 8'b11111111; //  779 : 255 - 0xff
      11'h30C: dout <= 8'b01111111; //  780 : 127 - 0x7f
      11'h30D: dout <= 8'b01110101; //  781 : 117 - 0x75
      11'h30E: dout <= 8'b11111111; //  782 : 255 - 0xff
      11'h30F: dout <= 8'b11111111; //  783 : 255 - 0xff
      11'h310: dout <= 8'b11111111; //  784 : 255 - 0xff -- Background 0x62
      11'h311: dout <= 8'b00000000; //  785 :   0 - 0x0
      11'h312: dout <= 8'b11000011; //  786 : 195 - 0xc3
      11'h313: dout <= 8'b10000001; //  787 : 129 - 0x81
      11'h314: dout <= 8'b10000001; //  788 : 129 - 0x81
      11'h315: dout <= 8'b11000011; //  789 : 195 - 0xc3
      11'h316: dout <= 8'b11111111; //  790 : 255 - 0xff
      11'h317: dout <= 8'b00000000; //  791 :   0 - 0x0
      11'h318: dout <= 8'b10000001; //  792 : 129 - 0x81 -- Background 0x63
      11'h319: dout <= 8'b01100110; //  793 : 102 - 0x66
      11'h31A: dout <= 8'b01111110; //  794 : 126 - 0x7e
      11'h31B: dout <= 8'b01111110; //  795 : 126 - 0x7e
      11'h31C: dout <= 8'b01111110; //  796 : 126 - 0x7e
      11'h31D: dout <= 8'b11111111; //  797 : 255 - 0xff
      11'h31E: dout <= 8'b11111111; //  798 : 255 - 0xff
      11'h31F: dout <= 8'b01111110; //  799 : 126 - 0x7e
      11'h320: dout <= 8'b00000000; //  800 :   0 - 0x0 -- Background 0x64
      11'h321: dout <= 8'b00000000; //  801 :   0 - 0x0
      11'h322: dout <= 8'b00000000; //  802 :   0 - 0x0
      11'h323: dout <= 8'b00000000; //  803 :   0 - 0x0
      11'h324: dout <= 8'b00000000; //  804 :   0 - 0x0
      11'h325: dout <= 8'b00000000; //  805 :   0 - 0x0
      11'h326: dout <= 8'b00000000; //  806 :   0 - 0x0
      11'h327: dout <= 8'b00000000; //  807 :   0 - 0x0
      11'h328: dout <= 8'b00000000; //  808 :   0 - 0x0 -- Background 0x65
      11'h329: dout <= 8'b00000000; //  809 :   0 - 0x0
      11'h32A: dout <= 8'b00000000; //  810 :   0 - 0x0
      11'h32B: dout <= 8'b00000000; //  811 :   0 - 0x0
      11'h32C: dout <= 8'b00000000; //  812 :   0 - 0x0
      11'h32D: dout <= 8'b00000000; //  813 :   0 - 0x0
      11'h32E: dout <= 8'b00000000; //  814 :   0 - 0x0
      11'h32F: dout <= 8'b00000000; //  815 :   0 - 0x0
      11'h330: dout <= 8'b00000000; //  816 :   0 - 0x0 -- Background 0x66
      11'h331: dout <= 8'b00000000; //  817 :   0 - 0x0
      11'h332: dout <= 8'b00000000; //  818 :   0 - 0x0
      11'h333: dout <= 8'b00000000; //  819 :   0 - 0x0
      11'h334: dout <= 8'b00000000; //  820 :   0 - 0x0
      11'h335: dout <= 8'b00000000; //  821 :   0 - 0x0
      11'h336: dout <= 8'b00000000; //  822 :   0 - 0x0
      11'h337: dout <= 8'b00000000; //  823 :   0 - 0x0
      11'h338: dout <= 8'b00000000; //  824 :   0 - 0x0 -- Background 0x67
      11'h339: dout <= 8'b00000000; //  825 :   0 - 0x0
      11'h33A: dout <= 8'b00000000; //  826 :   0 - 0x0
      11'h33B: dout <= 8'b00000000; //  827 :   0 - 0x0
      11'h33C: dout <= 8'b00000000; //  828 :   0 - 0x0
      11'h33D: dout <= 8'b00000000; //  829 :   0 - 0x0
      11'h33E: dout <= 8'b00000000; //  830 :   0 - 0x0
      11'h33F: dout <= 8'b00000000; //  831 :   0 - 0x0
      11'h340: dout <= 8'b00000011; //  832 :   3 - 0x3 -- Background 0x68
      11'h341: dout <= 8'b00000001; //  833 :   1 - 0x1
      11'h342: dout <= 8'b00000000; //  834 :   0 - 0x0
      11'h343: dout <= 8'b00000000; //  835 :   0 - 0x0
      11'h344: dout <= 8'b00000000; //  836 :   0 - 0x0
      11'h345: dout <= 8'b00000000; //  837 :   0 - 0x0
      11'h346: dout <= 8'b00000000; //  838 :   0 - 0x0
      11'h347: dout <= 8'b00000000; //  839 :   0 - 0x0
      11'h348: dout <= 8'b11111111; //  840 : 255 - 0xff -- Background 0x69
      11'h349: dout <= 8'b11111111; //  841 : 255 - 0xff
      11'h34A: dout <= 8'b11111111; //  842 : 255 - 0xff
      11'h34B: dout <= 8'b11111111; //  843 : 255 - 0xff
      11'h34C: dout <= 8'b11111111; //  844 : 255 - 0xff
      11'h34D: dout <= 8'b11111111; //  845 : 255 - 0xff
      11'h34E: dout <= 8'b11111111; //  846 : 255 - 0xff
      11'h34F: dout <= 8'b11111111; //  847 : 255 - 0xff
      11'h350: dout <= 8'b11000000; //  848 : 192 - 0xc0 -- Background 0x6a
      11'h351: dout <= 8'b10000000; //  849 : 128 - 0x80
      11'h352: dout <= 8'b00000000; //  850 :   0 - 0x0
      11'h353: dout <= 8'b00000000; //  851 :   0 - 0x0
      11'h354: dout <= 8'b00000000; //  852 :   0 - 0x0
      11'h355: dout <= 8'b00000000; //  853 :   0 - 0x0
      11'h356: dout <= 8'b00000000; //  854 :   0 - 0x0
      11'h357: dout <= 8'b00000000; //  855 :   0 - 0x0
      11'h358: dout <= 8'b11111111; //  856 : 255 - 0xff -- Background 0x6b
      11'h359: dout <= 8'b11111111; //  857 : 255 - 0xff
      11'h35A: dout <= 8'b11111111; //  858 : 255 - 0xff
      11'h35B: dout <= 8'b11111111; //  859 : 255 - 0xff
      11'h35C: dout <= 8'b11111111; //  860 : 255 - 0xff
      11'h35D: dout <= 8'b11111111; //  861 : 255 - 0xff
      11'h35E: dout <= 8'b11111111; //  862 : 255 - 0xff
      11'h35F: dout <= 8'b11111111; //  863 : 255 - 0xff
      11'h360: dout <= 8'b11111111; //  864 : 255 - 0xff -- Background 0x6c
      11'h361: dout <= 8'b11111111; //  865 : 255 - 0xff
      11'h362: dout <= 8'b11111111; //  866 : 255 - 0xff
      11'h363: dout <= 8'b00011111; //  867 :  31 - 0x1f
      11'h364: dout <= 8'b00011111; //  868 :  31 - 0x1f
      11'h365: dout <= 8'b00111111; //  869 :  63 - 0x3f
      11'h366: dout <= 8'b01111111; //  870 : 127 - 0x7f
      11'h367: dout <= 8'b11111111; //  871 : 255 - 0xff
      11'h368: dout <= 8'b11111111; //  872 : 255 - 0xff -- Background 0x6d
      11'h369: dout <= 8'b11111111; //  873 : 255 - 0xff
      11'h36A: dout <= 8'b11111111; //  874 : 255 - 0xff
      11'h36B: dout <= 8'b11111000; //  875 : 248 - 0xf8
      11'h36C: dout <= 8'b11111000; //  876 : 248 - 0xf8
      11'h36D: dout <= 8'b11111100; //  877 : 252 - 0xfc
      11'h36E: dout <= 8'b11111110; //  878 : 254 - 0xfe
      11'h36F: dout <= 8'b11111111; //  879 : 255 - 0xff
      11'h370: dout <= 8'b00000000; //  880 :   0 - 0x0 -- Background 0x6e
      11'h371: dout <= 8'b00000000; //  881 :   0 - 0x0
      11'h372: dout <= 8'b00000000; //  882 :   0 - 0x0
      11'h373: dout <= 8'b00000000; //  883 :   0 - 0x0
      11'h374: dout <= 8'b00000000; //  884 :   0 - 0x0
      11'h375: dout <= 8'b00111100; //  885 :  60 - 0x3c
      11'h376: dout <= 8'b01000010; //  886 :  66 - 0x42
      11'h377: dout <= 8'b10000001; //  887 : 129 - 0x81
      11'h378: dout <= 8'b10000001; //  888 : 129 - 0x81 -- Background 0x6f
      11'h379: dout <= 8'b10111101; //  889 : 189 - 0xbd
      11'h37A: dout <= 8'b01111110; //  890 : 126 - 0x7e
      11'h37B: dout <= 8'b10100101; //  891 : 165 - 0xa5
      11'h37C: dout <= 8'b11011011; //  892 : 219 - 0xdb
      11'h37D: dout <= 8'b11100111; //  893 : 231 - 0xe7
      11'h37E: dout <= 8'b11111111; //  894 : 255 - 0xff
      11'h37F: dout <= 8'b11111111; //  895 : 255 - 0xff
      11'h380: dout <= 8'b00000000; //  896 :   0 - 0x0 -- Background 0x70
      11'h381: dout <= 8'b00000101; //  897 :   5 - 0x5
      11'h382: dout <= 8'b00011001; //  898 :  25 - 0x19
      11'h383: dout <= 8'b00110011; //  899 :  51 - 0x33
      11'h384: dout <= 8'b01100011; //  900 :  99 - 0x63
      11'h385: dout <= 8'b11000111; //  901 : 199 - 0xc7
      11'h386: dout <= 8'b11000111; //  902 : 199 - 0xc7
      11'h387: dout <= 8'b11000100; //  903 : 196 - 0xc4
      11'h388: dout <= 8'b10000000; //  904 : 128 - 0x80 -- Background 0x71
      11'h389: dout <= 8'b00000000; //  905 :   0 - 0x0
      11'h38A: dout <= 8'b00000000; //  906 :   0 - 0x0
      11'h38B: dout <= 8'b00000001; //  907 :   1 - 0x1
      11'h38C: dout <= 8'b00000001; //  908 :   1 - 0x1
      11'h38D: dout <= 8'b00000001; //  909 :   1 - 0x1
      11'h38E: dout <= 8'b00000000; //  910 :   0 - 0x0
      11'h38F: dout <= 8'b00000000; //  911 :   0 - 0x0
      11'h390: dout <= 8'b00000000; //  912 :   0 - 0x0 -- Background 0x72
      11'h391: dout <= 8'b10100000; //  913 : 160 - 0xa0
      11'h392: dout <= 8'b10011000; //  914 : 152 - 0x98
      11'h393: dout <= 8'b11001100; //  915 : 204 - 0xcc
      11'h394: dout <= 8'b11000110; //  916 : 198 - 0xc6
      11'h395: dout <= 8'b11100011; //  917 : 227 - 0xe3
      11'h396: dout <= 8'b11100011; //  918 : 227 - 0xe3
      11'h397: dout <= 8'b00100011; //  919 :  35 - 0x23
      11'h398: dout <= 8'b00000001; //  920 :   1 - 0x1 -- Background 0x73
      11'h399: dout <= 8'b00000000; //  921 :   0 - 0x0
      11'h39A: dout <= 8'b00000000; //  922 :   0 - 0x0
      11'h39B: dout <= 8'b00000000; //  923 :   0 - 0x0
      11'h39C: dout <= 8'b00000000; //  924 :   0 - 0x0
      11'h39D: dout <= 8'b01000000; //  925 :  64 - 0x40
      11'h39E: dout <= 8'b10000000; //  926 : 128 - 0x80
      11'h39F: dout <= 8'b00000000; //  927 :   0 - 0x0
      11'h3A0: dout <= 8'b00000001; //  928 :   1 - 0x1 -- Background 0x74
      11'h3A1: dout <= 8'b00000001; //  929 :   1 - 0x1
      11'h3A2: dout <= 8'b00000001; //  930 :   1 - 0x1
      11'h3A3: dout <= 8'b00000001; //  931 :   1 - 0x1
      11'h3A4: dout <= 8'b00000001; //  932 :   1 - 0x1
      11'h3A5: dout <= 8'b00000001; //  933 :   1 - 0x1
      11'h3A6: dout <= 8'b00000001; //  934 :   1 - 0x1
      11'h3A7: dout <= 8'b00000001; //  935 :   1 - 0x1
      11'h3A8: dout <= 8'b10000000; //  936 : 128 - 0x80 -- Background 0x75
      11'h3A9: dout <= 8'b10000000; //  937 : 128 - 0x80
      11'h3AA: dout <= 8'b10000000; //  938 : 128 - 0x80
      11'h3AB: dout <= 8'b10000000; //  939 : 128 - 0x80
      11'h3AC: dout <= 8'b10000000; //  940 : 128 - 0x80
      11'h3AD: dout <= 8'b10000000; //  941 : 128 - 0x80
      11'h3AE: dout <= 8'b10000000; //  942 : 128 - 0x80
      11'h3AF: dout <= 8'b10000000; //  943 : 128 - 0x80
      11'h3B0: dout <= 8'b00000001; //  944 :   1 - 0x1 -- Background 0x76
      11'h3B1: dout <= 8'b00000011; //  945 :   3 - 0x3
      11'h3B2: dout <= 8'b00000011; //  946 :   3 - 0x3
      11'h3B3: dout <= 8'b00000111; //  947 :   7 - 0x7
      11'h3B4: dout <= 8'b00000100; //  948 :   4 - 0x4
      11'h3B5: dout <= 8'b00011100; //  949 :  28 - 0x1c
      11'h3B6: dout <= 8'b00111111; //  950 :  63 - 0x3f
      11'h3B7: dout <= 8'b01111111; //  951 : 127 - 0x7f
      11'h3B8: dout <= 8'b01111111; //  952 : 127 - 0x7f -- Background 0x77
      11'h3B9: dout <= 8'b11111111; //  953 : 255 - 0xff
      11'h3BA: dout <= 8'b11111111; //  954 : 255 - 0xff
      11'h3BB: dout <= 8'b01111111; //  955 : 127 - 0x7f
      11'h3BC: dout <= 8'b01111111; //  956 : 127 - 0x7f
      11'h3BD: dout <= 8'b00011111; //  957 :  31 - 0x1f
      11'h3BE: dout <= 8'b00000011; //  958 :   3 - 0x3
      11'h3BF: dout <= 8'b00000000; //  959 :   0 - 0x0
      11'h3C0: dout <= 8'b00000000; //  960 :   0 - 0x0 -- Background 0x78
      11'h3C1: dout <= 8'b00000000; //  961 :   0 - 0x0
      11'h3C2: dout <= 8'b00000001; //  962 :   1 - 0x1
      11'h3C3: dout <= 8'b00000001; //  963 :   1 - 0x1
      11'h3C4: dout <= 8'b00000011; //  964 :   3 - 0x3
      11'h3C5: dout <= 8'b00000111; //  965 :   7 - 0x7
      11'h3C6: dout <= 8'b00000111; //  966 :   7 - 0x7
      11'h3C7: dout <= 8'b00001111; //  967 :  15 - 0xf
      11'h3C8: dout <= 8'b11111111; //  968 : 255 - 0xff -- Background 0x79
      11'h3C9: dout <= 8'b11111111; //  969 : 255 - 0xff
      11'h3CA: dout <= 8'b00111111; //  970 :  63 - 0x3f
      11'h3CB: dout <= 8'b00111111; //  971 :  63 - 0x3f
      11'h3CC: dout <= 8'b01111111; //  972 : 127 - 0x7f
      11'h3CD: dout <= 8'b11111110; //  973 : 254 - 0xfe
      11'h3CE: dout <= 8'b11111100; //  974 : 252 - 0xfc
      11'h3CF: dout <= 8'b00110000; //  975 :  48 - 0x30
      11'h3D0: dout <= 8'b11111000; //  976 : 248 - 0xf8 -- Background 0x7a
      11'h3D1: dout <= 8'b11111110; //  977 : 254 - 0xfe
      11'h3D2: dout <= 8'b11111111; //  978 : 255 - 0xff
      11'h3D3: dout <= 8'b11111111; //  979 : 255 - 0xff
      11'h3D4: dout <= 8'b11111111; //  980 : 255 - 0xff
      11'h3D5: dout <= 8'b11111111; //  981 : 255 - 0xff
      11'h3D6: dout <= 8'b11111111; //  982 : 255 - 0xff
      11'h3D7: dout <= 8'b11111111; //  983 : 255 - 0xff
      11'h3D8: dout <= 8'b11111111; //  984 : 255 - 0xff -- Background 0x7b
      11'h3D9: dout <= 8'b11111111; //  985 : 255 - 0xff
      11'h3DA: dout <= 8'b11111111; //  986 : 255 - 0xff
      11'h3DB: dout <= 8'b11111111; //  987 : 255 - 0xff
      11'h3DC: dout <= 8'b11111111; //  988 : 255 - 0xff
      11'h3DD: dout <= 8'b11111111; //  989 : 255 - 0xff
      11'h3DE: dout <= 8'b11111111; //  990 : 255 - 0xff
      11'h3DF: dout <= 8'b01111111; //  991 : 127 - 0x7f
      11'h3E0: dout <= 8'b11111111; //  992 : 255 - 0xff -- Background 0x7c
      11'h3E1: dout <= 8'b11111111; //  993 : 255 - 0xff
      11'h3E2: dout <= 8'b11111111; //  994 : 255 - 0xff
      11'h3E3: dout <= 8'b11111111; //  995 : 255 - 0xff
      11'h3E4: dout <= 8'b11111111; //  996 : 255 - 0xff
      11'h3E5: dout <= 8'b11111111; //  997 : 255 - 0xff
      11'h3E6: dout <= 8'b11111111; //  998 : 255 - 0xff
      11'h3E7: dout <= 8'b11111111; //  999 : 255 - 0xff
      11'h3E8: dout <= 8'b11101111; // 1000 : 239 - 0xef -- Background 0x7d
      11'h3E9: dout <= 8'b11001111; // 1001 : 207 - 0xcf
      11'h3EA: dout <= 8'b10011111; // 1002 : 159 - 0x9f
      11'h3EB: dout <= 8'b00011111; // 1003 :  31 - 0x1f
      11'h3EC: dout <= 8'b00001111; // 1004 :  15 - 0xf
      11'h3ED: dout <= 8'b01111111; // 1005 : 127 - 0x7f
      11'h3EE: dout <= 8'b11111111; // 1006 : 255 - 0xff
      11'h3EF: dout <= 8'b11111111; // 1007 : 255 - 0xff
      11'h3F0: dout <= 8'b00000000; // 1008 :   0 - 0x0 -- Background 0x7e
      11'h3F1: dout <= 8'b00000000; // 1009 :   0 - 0x0
      11'h3F2: dout <= 8'b00000000; // 1010 :   0 - 0x0
      11'h3F3: dout <= 8'b11110000; // 1011 : 240 - 0xf0
      11'h3F4: dout <= 8'b11111110; // 1012 : 254 - 0xfe
      11'h3F5: dout <= 8'b11111111; // 1013 : 255 - 0xff
      11'h3F6: dout <= 8'b11111111; // 1014 : 255 - 0xff
      11'h3F7: dout <= 8'b11111111; // 1015 : 255 - 0xff
      11'h3F8: dout <= 8'b11111111; // 1016 : 255 - 0xff -- Background 0x7f
      11'h3F9: dout <= 8'b11111111; // 1017 : 255 - 0xff
      11'h3FA: dout <= 8'b11111111; // 1018 : 255 - 0xff
      11'h3FB: dout <= 8'b11111111; // 1019 : 255 - 0xff
      11'h3FC: dout <= 8'b11111111; // 1020 : 255 - 0xff
      11'h3FD: dout <= 8'b11111111; // 1021 : 255 - 0xff
      11'h3FE: dout <= 8'b11111111; // 1022 : 255 - 0xff
      11'h3FF: dout <= 8'b11111111; // 1023 : 255 - 0xff
      11'h400: dout <= 8'b11111111; // 1024 : 255 - 0xff -- Background 0x80
      11'h401: dout <= 8'b11111111; // 1025 : 255 - 0xff
      11'h402: dout <= 8'b11111111; // 1026 : 255 - 0xff
      11'h403: dout <= 8'b11111111; // 1027 : 255 - 0xff
      11'h404: dout <= 8'b11111111; // 1028 : 255 - 0xff
      11'h405: dout <= 8'b11111111; // 1029 : 255 - 0xff
      11'h406: dout <= 8'b11111111; // 1030 : 255 - 0xff
      11'h407: dout <= 8'b11111111; // 1031 : 255 - 0xff
      11'h408: dout <= 8'b11111111; // 1032 : 255 - 0xff -- Background 0x81
      11'h409: dout <= 8'b11111111; // 1033 : 255 - 0xff
      11'h40A: dout <= 8'b11111111; // 1034 : 255 - 0xff
      11'h40B: dout <= 8'b11110000; // 1035 : 240 - 0xf0
      11'h40C: dout <= 8'b11110000; // 1036 : 240 - 0xf0
      11'h40D: dout <= 8'b11111000; // 1037 : 248 - 0xf8
      11'h40E: dout <= 8'b11111000; // 1038 : 248 - 0xf8
      11'h40F: dout <= 8'b11111000; // 1039 : 248 - 0xf8
      11'h410: dout <= 8'b00000000; // 1040 :   0 - 0x0 -- Background 0x82
      11'h411: dout <= 8'b00000000; // 1041 :   0 - 0x0
      11'h412: dout <= 8'b00000000; // 1042 :   0 - 0x0
      11'h413: dout <= 8'b00000000; // 1043 :   0 - 0x0
      11'h414: dout <= 8'b00000000; // 1044 :   0 - 0x0
      11'h415: dout <= 8'b10000000; // 1045 : 128 - 0x80
      11'h416: dout <= 8'b11000000; // 1046 : 192 - 0xc0
      11'h417: dout <= 8'b11100000; // 1047 : 224 - 0xe0
      11'h418: dout <= 8'b11110000; // 1048 : 240 - 0xf0 -- Background 0x83
      11'h419: dout <= 8'b11110000; // 1049 : 240 - 0xf0
      11'h41A: dout <= 8'b11111000; // 1050 : 248 - 0xf8
      11'h41B: dout <= 8'b11111000; // 1051 : 248 - 0xf8
      11'h41C: dout <= 8'b11111000; // 1052 : 248 - 0xf8
      11'h41D: dout <= 8'b11111100; // 1053 : 252 - 0xfc
      11'h41E: dout <= 8'b11111100; // 1054 : 252 - 0xfc
      11'h41F: dout <= 8'b11111110; // 1055 : 254 - 0xfe
      11'h420: dout <= 8'b11111111; // 1056 : 255 - 0xff -- Background 0x84
      11'h421: dout <= 8'b11111111; // 1057 : 255 - 0xff
      11'h422: dout <= 8'b11111111; // 1058 : 255 - 0xff
      11'h423: dout <= 8'b11111111; // 1059 : 255 - 0xff
      11'h424: dout <= 8'b11111111; // 1060 : 255 - 0xff
      11'h425: dout <= 8'b11111111; // 1061 : 255 - 0xff
      11'h426: dout <= 8'b11111111; // 1062 : 255 - 0xff
      11'h427: dout <= 8'b11111111; // 1063 : 255 - 0xff
      11'h428: dout <= 8'b11111111; // 1064 : 255 - 0xff -- Background 0x85
      11'h429: dout <= 8'b11111111; // 1065 : 255 - 0xff
      11'h42A: dout <= 8'b11111111; // 1066 : 255 - 0xff
      11'h42B: dout <= 8'b00001111; // 1067 :  15 - 0xf
      11'h42C: dout <= 8'b00000111; // 1068 :   7 - 0x7
      11'h42D: dout <= 8'b00000000; // 1069 :   0 - 0x0
      11'h42E: dout <= 8'b00000000; // 1070 :   0 - 0x0
      11'h42F: dout <= 8'b00000000; // 1071 :   0 - 0x0
      11'h430: dout <= 8'b00000000; // 1072 :   0 - 0x0 -- Background 0x86
      11'h431: dout <= 8'b10000000; // 1073 : 128 - 0x80
      11'h432: dout <= 8'b11000000; // 1074 : 192 - 0xc0
      11'h433: dout <= 8'b11100000; // 1075 : 224 - 0xe0
      11'h434: dout <= 8'b11110000; // 1076 : 240 - 0xf0
      11'h435: dout <= 8'b11110000; // 1077 : 240 - 0xf0
      11'h436: dout <= 8'b11110000; // 1078 : 240 - 0xf0
      11'h437: dout <= 8'b11111100; // 1079 : 252 - 0xfc
      11'h438: dout <= 8'b11111111; // 1080 : 255 - 0xff -- Background 0x87
      11'h439: dout <= 8'b11111111; // 1081 : 255 - 0xff
      11'h43A: dout <= 8'b11111111; // 1082 : 255 - 0xff
      11'h43B: dout <= 8'b11111111; // 1083 : 255 - 0xff
      11'h43C: dout <= 8'b11111111; // 1084 : 255 - 0xff
      11'h43D: dout <= 8'b00001111; // 1085 :  15 - 0xf
      11'h43E: dout <= 8'b00011111; // 1086 :  31 - 0x1f
      11'h43F: dout <= 8'b00111111; // 1087 :  63 - 0x3f
      11'h440: dout <= 8'b11000000; // 1088 : 192 - 0xc0 -- Background 0x88
      11'h441: dout <= 8'b11100000; // 1089 : 224 - 0xe0
      11'h442: dout <= 8'b11100000; // 1090 : 224 - 0xe0
      11'h443: dout <= 8'b11100000; // 1091 : 224 - 0xe0
      11'h444: dout <= 8'b11100000; // 1092 : 224 - 0xe0
      11'h445: dout <= 8'b11000000; // 1093 : 192 - 0xc0
      11'h446: dout <= 8'b11000000; // 1094 : 192 - 0xc0
      11'h447: dout <= 8'b10000000; // 1095 : 128 - 0x80
      11'h448: dout <= 8'b00000011; // 1096 :   3 - 0x3 -- Background 0x89
      11'h449: dout <= 8'b00000111; // 1097 :   7 - 0x7
      11'h44A: dout <= 8'b00000111; // 1098 :   7 - 0x7
      11'h44B: dout <= 8'b00000111; // 1099 :   7 - 0x7
      11'h44C: dout <= 8'b00000111; // 1100 :   7 - 0x7
      11'h44D: dout <= 8'b00000011; // 1101 :   3 - 0x3
      11'h44E: dout <= 8'b00000011; // 1102 :   3 - 0x3
      11'h44F: dout <= 8'b00000001; // 1103 :   1 - 0x1
      11'h450: dout <= 8'b00000000; // 1104 :   0 - 0x0 -- Background 0x8a
      11'h451: dout <= 8'b00000001; // 1105 :   1 - 0x1
      11'h452: dout <= 8'b00000011; // 1106 :   3 - 0x3
      11'h453: dout <= 8'b00000111; // 1107 :   7 - 0x7
      11'h454: dout <= 8'b00001111; // 1108 :  15 - 0xf
      11'h455: dout <= 8'b00001111; // 1109 :  15 - 0xf
      11'h456: dout <= 8'b00001111; // 1110 :  15 - 0xf
      11'h457: dout <= 8'b00111111; // 1111 :  63 - 0x3f
      11'h458: dout <= 8'b11111111; // 1112 : 255 - 0xff -- Background 0x8b
      11'h459: dout <= 8'b11111111; // 1113 : 255 - 0xff
      11'h45A: dout <= 8'b11111111; // 1114 : 255 - 0xff
      11'h45B: dout <= 8'b11111111; // 1115 : 255 - 0xff
      11'h45C: dout <= 8'b11111111; // 1116 : 255 - 0xff
      11'h45D: dout <= 8'b11110000; // 1117 : 240 - 0xf0
      11'h45E: dout <= 8'b11111000; // 1118 : 248 - 0xf8
      11'h45F: dout <= 8'b11111100; // 1119 : 252 - 0xfc
      11'h460: dout <= 8'b00000000; // 1120 :   0 - 0x0 -- Background 0x8c
      11'h461: dout <= 8'b00000000; // 1121 :   0 - 0x0
      11'h462: dout <= 8'b00000000; // 1122 :   0 - 0x0
      11'h463: dout <= 8'b00000000; // 1123 :   0 - 0x0
      11'h464: dout <= 8'b00000000; // 1124 :   0 - 0x0
      11'h465: dout <= 8'b00000001; // 1125 :   1 - 0x1
      11'h466: dout <= 8'b00000011; // 1126 :   3 - 0x3
      11'h467: dout <= 8'b00000111; // 1127 :   7 - 0x7
      11'h468: dout <= 8'b00001111; // 1128 :  15 - 0xf -- Background 0x8d
      11'h469: dout <= 8'b00001111; // 1129 :  15 - 0xf
      11'h46A: dout <= 8'b00011111; // 1130 :  31 - 0x1f
      11'h46B: dout <= 8'b00011111; // 1131 :  31 - 0x1f
      11'h46C: dout <= 8'b00011111; // 1132 :  31 - 0x1f
      11'h46D: dout <= 8'b00111111; // 1133 :  63 - 0x3f
      11'h46E: dout <= 8'b00111111; // 1134 :  63 - 0x3f
      11'h46F: dout <= 8'b01111111; // 1135 : 127 - 0x7f
      11'h470: dout <= 8'b11111111; // 1136 : 255 - 0xff -- Background 0x8e
      11'h471: dout <= 8'b11111111; // 1137 : 255 - 0xff
      11'h472: dout <= 8'b11111111; // 1138 : 255 - 0xff
      11'h473: dout <= 8'b11111111; // 1139 : 255 - 0xff
      11'h474: dout <= 8'b11111111; // 1140 : 255 - 0xff
      11'h475: dout <= 8'b11111111; // 1141 : 255 - 0xff
      11'h476: dout <= 8'b11111111; // 1142 : 255 - 0xff
      11'h477: dout <= 8'b11111111; // 1143 : 255 - 0xff
      11'h478: dout <= 8'b11111111; // 1144 : 255 - 0xff -- Background 0x8f
      11'h479: dout <= 8'b11111111; // 1145 : 255 - 0xff
      11'h47A: dout <= 8'b11111111; // 1146 : 255 - 0xff
      11'h47B: dout <= 8'b11110000; // 1147 : 240 - 0xf0
      11'h47C: dout <= 8'b11100000; // 1148 : 224 - 0xe0
      11'h47D: dout <= 8'b00000000; // 1149 :   0 - 0x0
      11'h47E: dout <= 8'b00000000; // 1150 :   0 - 0x0
      11'h47F: dout <= 8'b00000000; // 1151 :   0 - 0x0
      11'h480: dout <= 8'b00000000; // 1152 :   0 - 0x0 -- Background 0x90
      11'h481: dout <= 8'b00000000; // 1153 :   0 - 0x0
      11'h482: dout <= 8'b00000000; // 1154 :   0 - 0x0
      11'h483: dout <= 8'b00001111; // 1155 :  15 - 0xf
      11'h484: dout <= 8'b01111111; // 1156 : 127 - 0x7f
      11'h485: dout <= 8'b11111111; // 1157 : 255 - 0xff
      11'h486: dout <= 8'b11111111; // 1158 : 255 - 0xff
      11'h487: dout <= 8'b11111111; // 1159 : 255 - 0xff
      11'h488: dout <= 8'b11111111; // 1160 : 255 - 0xff -- Background 0x91
      11'h489: dout <= 8'b11111111; // 1161 : 255 - 0xff
      11'h48A: dout <= 8'b11111111; // 1162 : 255 - 0xff
      11'h48B: dout <= 8'b11111111; // 1163 : 255 - 0xff
      11'h48C: dout <= 8'b11111111; // 1164 : 255 - 0xff
      11'h48D: dout <= 8'b11111111; // 1165 : 255 - 0xff
      11'h48E: dout <= 8'b11111111; // 1166 : 255 - 0xff
      11'h48F: dout <= 8'b11111111; // 1167 : 255 - 0xff
      11'h490: dout <= 8'b11111111; // 1168 : 255 - 0xff -- Background 0x92
      11'h491: dout <= 8'b11111111; // 1169 : 255 - 0xff
      11'h492: dout <= 8'b11111111; // 1170 : 255 - 0xff
      11'h493: dout <= 8'b11111111; // 1171 : 255 - 0xff
      11'h494: dout <= 8'b11111111; // 1172 : 255 - 0xff
      11'h495: dout <= 8'b11111111; // 1173 : 255 - 0xff
      11'h496: dout <= 8'b11111111; // 1174 : 255 - 0xff
      11'h497: dout <= 8'b11111111; // 1175 : 255 - 0xff
      11'h498: dout <= 8'b11111111; // 1176 : 255 - 0xff -- Background 0x93
      11'h499: dout <= 8'b11111111; // 1177 : 255 - 0xff
      11'h49A: dout <= 8'b11111111; // 1178 : 255 - 0xff
      11'h49B: dout <= 8'b00001111; // 1179 :  15 - 0xf
      11'h49C: dout <= 8'b00001111; // 1180 :  15 - 0xf
      11'h49D: dout <= 8'b00011111; // 1181 :  31 - 0x1f
      11'h49E: dout <= 8'b00011111; // 1182 :  31 - 0x1f
      11'h49F: dout <= 8'b00011111; // 1183 :  31 - 0x1f
      11'h4A0: dout <= 8'b00011111; // 1184 :  31 - 0x1f -- Background 0x94
      11'h4A1: dout <= 8'b01111111; // 1185 : 127 - 0x7f
      11'h4A2: dout <= 8'b11111111; // 1186 : 255 - 0xff
      11'h4A3: dout <= 8'b11111111; // 1187 : 255 - 0xff
      11'h4A4: dout <= 8'b11111111; // 1188 : 255 - 0xff
      11'h4A5: dout <= 8'b11111111; // 1189 : 255 - 0xff
      11'h4A6: dout <= 8'b11111111; // 1190 : 255 - 0xff
      11'h4A7: dout <= 8'b11111111; // 1191 : 255 - 0xff
      11'h4A8: dout <= 8'b11111111; // 1192 : 255 - 0xff -- Background 0x95
      11'h4A9: dout <= 8'b11111111; // 1193 : 255 - 0xff
      11'h4AA: dout <= 8'b11111111; // 1194 : 255 - 0xff
      11'h4AB: dout <= 8'b11111111; // 1195 : 255 - 0xff
      11'h4AC: dout <= 8'b11111111; // 1196 : 255 - 0xff
      11'h4AD: dout <= 8'b11111111; // 1197 : 255 - 0xff
      11'h4AE: dout <= 8'b11111111; // 1198 : 255 - 0xff
      11'h4AF: dout <= 8'b11111110; // 1199 : 254 - 0xfe
      11'h4B0: dout <= 8'b11111111; // 1200 : 255 - 0xff -- Background 0x96
      11'h4B1: dout <= 8'b11111111; // 1201 : 255 - 0xff
      11'h4B2: dout <= 8'b11111111; // 1202 : 255 - 0xff
      11'h4B3: dout <= 8'b11111111; // 1203 : 255 - 0xff
      11'h4B4: dout <= 8'b11111111; // 1204 : 255 - 0xff
      11'h4B5: dout <= 8'b11111111; // 1205 : 255 - 0xff
      11'h4B6: dout <= 8'b11111111; // 1206 : 255 - 0xff
      11'h4B7: dout <= 8'b11111111; // 1207 : 255 - 0xff
      11'h4B8: dout <= 8'b11110111; // 1208 : 247 - 0xf7 -- Background 0x97
      11'h4B9: dout <= 8'b11110011; // 1209 : 243 - 0xf3
      11'h4BA: dout <= 8'b11111001; // 1210 : 249 - 0xf9
      11'h4BB: dout <= 8'b11111000; // 1211 : 248 - 0xf8
      11'h4BC: dout <= 8'b11110000; // 1212 : 240 - 0xf0
      11'h4BD: dout <= 8'b11111110; // 1213 : 254 - 0xfe
      11'h4BE: dout <= 8'b11111111; // 1214 : 255 - 0xff
      11'h4BF: dout <= 8'b11111111; // 1215 : 255 - 0xff
      11'h4C0: dout <= 8'b10000000; // 1216 : 128 - 0x80 -- Background 0x98
      11'h4C1: dout <= 8'b11000000; // 1217 : 192 - 0xc0
      11'h4C2: dout <= 8'b11000000; // 1218 : 192 - 0xc0
      11'h4C3: dout <= 8'b11100000; // 1219 : 224 - 0xe0
      11'h4C4: dout <= 8'b00100000; // 1220 :  32 - 0x20
      11'h4C5: dout <= 8'b00111000; // 1221 :  56 - 0x38
      11'h4C6: dout <= 8'b11111100; // 1222 : 252 - 0xfc
      11'h4C7: dout <= 8'b11111110; // 1223 : 254 - 0xfe
      11'h4C8: dout <= 8'b11111110; // 1224 : 254 - 0xfe -- Background 0x99
      11'h4C9: dout <= 8'b11111111; // 1225 : 255 - 0xff
      11'h4CA: dout <= 8'b11111111; // 1226 : 255 - 0xff
      11'h4CB: dout <= 8'b11111110; // 1227 : 254 - 0xfe
      11'h4CC: dout <= 8'b11111100; // 1228 : 252 - 0xfc
      11'h4CD: dout <= 8'b11111000; // 1229 : 248 - 0xf8
      11'h4CE: dout <= 8'b11000000; // 1230 : 192 - 0xc0
      11'h4CF: dout <= 8'b00000000; // 1231 :   0 - 0x0
      11'h4D0: dout <= 8'b00000000; // 1232 :   0 - 0x0 -- Background 0x9a
      11'h4D1: dout <= 8'b00000000; // 1233 :   0 - 0x0
      11'h4D2: dout <= 8'b10000000; // 1234 : 128 - 0x80
      11'h4D3: dout <= 8'b10000000; // 1235 : 128 - 0x80
      11'h4D4: dout <= 8'b11000000; // 1236 : 192 - 0xc0
      11'h4D5: dout <= 8'b11100000; // 1237 : 224 - 0xe0
      11'h4D6: dout <= 8'b11100000; // 1238 : 224 - 0xe0
      11'h4D7: dout <= 8'b11110000; // 1239 : 240 - 0xf0
      11'h4D8: dout <= 8'b11111111; // 1240 : 255 - 0xff -- Background 0x9b
      11'h4D9: dout <= 8'b11111111; // 1241 : 255 - 0xff
      11'h4DA: dout <= 8'b11111100; // 1242 : 252 - 0xfc
      11'h4DB: dout <= 8'b11111100; // 1243 : 252 - 0xfc
      11'h4DC: dout <= 8'b11111110; // 1244 : 254 - 0xfe
      11'h4DD: dout <= 8'b01111110; // 1245 : 126 - 0x7e
      11'h4DE: dout <= 8'b00111111; // 1246 :  63 - 0x3f
      11'h4DF: dout <= 8'b00001100; // 1247 :  12 - 0xc
      11'h4E0: dout <= 8'b00000000; // 1248 :   0 - 0x0 -- Background 0x9c
      11'h4E1: dout <= 8'b00000001; // 1249 :   1 - 0x1
      11'h4E2: dout <= 8'b00000011; // 1250 :   3 - 0x3
      11'h4E3: dout <= 8'b00000111; // 1251 :   7 - 0x7
      11'h4E4: dout <= 8'b00000111; // 1252 :   7 - 0x7
      11'h4E5: dout <= 8'b00000111; // 1253 :   7 - 0x7
      11'h4E6: dout <= 8'b00001111; // 1254 :  15 - 0xf
      11'h4E7: dout <= 8'b00001111; // 1255 :  15 - 0xf
      11'h4E8: dout <= 8'b00001111; // 1256 :  15 - 0xf -- Background 0x9d
      11'h4E9: dout <= 8'b00001111; // 1257 :  15 - 0xf
      11'h4EA: dout <= 8'b00000111; // 1258 :   7 - 0x7
      11'h4EB: dout <= 8'b00000111; // 1259 :   7 - 0x7
      11'h4EC: dout <= 8'b00000111; // 1260 :   7 - 0x7
      11'h4ED: dout <= 8'b00000011; // 1261 :   3 - 0x3
      11'h4EE: dout <= 8'b00000011; // 1262 :   3 - 0x3
      11'h4EF: dout <= 8'b00000001; // 1263 :   1 - 0x1
      11'h4F0: dout <= 8'b00000001; // 1264 :   1 - 0x1 -- Background 0x9e
      11'h4F1: dout <= 8'b00000001; // 1265 :   1 - 0x1
      11'h4F2: dout <= 8'b00000001; // 1266 :   1 - 0x1
      11'h4F3: dout <= 8'b00000000; // 1267 :   0 - 0x0
      11'h4F4: dout <= 8'b00000000; // 1268 :   0 - 0x0
      11'h4F5: dout <= 8'b00000011; // 1269 :   3 - 0x3
      11'h4F6: dout <= 8'b00000111; // 1270 :   7 - 0x7
      11'h4F7: dout <= 8'b00001111; // 1271 :  15 - 0xf
      11'h4F8: dout <= 8'b00000000; // 1272 :   0 - 0x0 -- Background 0x9f
      11'h4F9: dout <= 8'b00000000; // 1273 :   0 - 0x0
      11'h4FA: dout <= 8'b00000000; // 1274 :   0 - 0x0
      11'h4FB: dout <= 8'b00000000; // 1275 :   0 - 0x0
      11'h4FC: dout <= 8'b00000001; // 1276 :   1 - 0x1
      11'h4FD: dout <= 8'b00000011; // 1277 :   3 - 0x3
      11'h4FE: dout <= 8'b00111111; // 1278 :  63 - 0x3f
      11'h4FF: dout <= 8'b01111111; // 1279 : 127 - 0x7f
      11'h500: dout <= 8'b11111111; // 1280 : 255 - 0xff -- Background 0xa0
      11'h501: dout <= 8'b11111111; // 1281 : 255 - 0xff
      11'h502: dout <= 8'b11111111; // 1282 : 255 - 0xff
      11'h503: dout <= 8'b11111111; // 1283 : 255 - 0xff
      11'h504: dout <= 8'b11111111; // 1284 : 255 - 0xff
      11'h505: dout <= 8'b11111111; // 1285 : 255 - 0xff
      11'h506: dout <= 8'b11111101; // 1286 : 253 - 0xfd
      11'h507: dout <= 8'b11111001; // 1287 : 249 - 0xf9
      11'h508: dout <= 8'b11110011; // 1288 : 243 - 0xf3 -- Background 0xa1
      11'h509: dout <= 8'b11111111; // 1289 : 255 - 0xff
      11'h50A: dout <= 8'b11111111; // 1290 : 255 - 0xff
      11'h50B: dout <= 8'b11111111; // 1291 : 255 - 0xff
      11'h50C: dout <= 8'b11111111; // 1292 : 255 - 0xff
      11'h50D: dout <= 8'b11111111; // 1293 : 255 - 0xff
      11'h50E: dout <= 8'b11111111; // 1294 : 255 - 0xff
      11'h50F: dout <= 8'b11111111; // 1295 : 255 - 0xff
      11'h510: dout <= 8'b11111111; // 1296 : 255 - 0xff -- Background 0xa2
      11'h511: dout <= 8'b11111111; // 1297 : 255 - 0xff
      11'h512: dout <= 8'b11111111; // 1298 : 255 - 0xff
      11'h513: dout <= 8'b11111111; // 1299 : 255 - 0xff
      11'h514: dout <= 8'b11111111; // 1300 : 255 - 0xff
      11'h515: dout <= 8'b11111111; // 1301 : 255 - 0xff
      11'h516: dout <= 8'b11111111; // 1302 : 255 - 0xff
      11'h517: dout <= 8'b11111111; // 1303 : 255 - 0xff
      11'h518: dout <= 8'b00000111; // 1304 :   7 - 0x7 -- Background 0xa3
      11'h519: dout <= 8'b00001111; // 1305 :  15 - 0xf
      11'h51A: dout <= 8'b00011111; // 1306 :  31 - 0x1f
      11'h51B: dout <= 8'b00111111; // 1307 :  63 - 0x3f
      11'h51C: dout <= 8'b11111100; // 1308 : 252 - 0xfc
      11'h51D: dout <= 8'b11111100; // 1309 : 252 - 0xfc
      11'h51E: dout <= 8'b11111111; // 1310 : 255 - 0xff
      11'h51F: dout <= 8'b11111111; // 1311 : 255 - 0xff
      11'h520: dout <= 8'b11111111; // 1312 : 255 - 0xff -- Background 0xa4
      11'h521: dout <= 8'b11111111; // 1313 : 255 - 0xff
      11'h522: dout <= 8'b11111111; // 1314 : 255 - 0xff
      11'h523: dout <= 8'b11111111; // 1315 : 255 - 0xff
      11'h524: dout <= 8'b11111111; // 1316 : 255 - 0xff
      11'h525: dout <= 8'b11111111; // 1317 : 255 - 0xff
      11'h526: dout <= 8'b11111111; // 1318 : 255 - 0xff
      11'h527: dout <= 8'b11111111; // 1319 : 255 - 0xff
      11'h528: dout <= 8'b11111111; // 1320 : 255 - 0xff -- Background 0xa5
      11'h529: dout <= 8'b11111111; // 1321 : 255 - 0xff
      11'h52A: dout <= 8'b11111111; // 1322 : 255 - 0xff
      11'h52B: dout <= 8'b11111111; // 1323 : 255 - 0xff
      11'h52C: dout <= 8'b11111111; // 1324 : 255 - 0xff
      11'h52D: dout <= 8'b11111111; // 1325 : 255 - 0xff
      11'h52E: dout <= 8'b11111111; // 1326 : 255 - 0xff
      11'h52F: dout <= 8'b11111111; // 1327 : 255 - 0xff
      11'h530: dout <= 8'b11111111; // 1328 : 255 - 0xff -- Background 0xa6
      11'h531: dout <= 8'b11111111; // 1329 : 255 - 0xff
      11'h532: dout <= 8'b11110000; // 1330 : 240 - 0xf0
      11'h533: dout <= 8'b11100000; // 1331 : 224 - 0xe0
      11'h534: dout <= 8'b11000000; // 1332 : 192 - 0xc0
      11'h535: dout <= 8'b10000000; // 1333 : 128 - 0x80
      11'h536: dout <= 8'b10000000; // 1334 : 128 - 0x80
      11'h537: dout <= 8'b00000000; // 1335 :   0 - 0x0
      11'h538: dout <= 8'b11110000; // 1336 : 240 - 0xf0 -- Background 0xa7
      11'h539: dout <= 8'b11111000; // 1337 : 248 - 0xf8
      11'h53A: dout <= 8'b11111100; // 1338 : 252 - 0xfc
      11'h53B: dout <= 8'b11111110; // 1339 : 254 - 0xfe
      11'h53C: dout <= 8'b10011111; // 1340 : 159 - 0x9f
      11'h53D: dout <= 8'b10011111; // 1341 : 159 - 0x9f
      11'h53E: dout <= 8'b11111111; // 1342 : 255 - 0xff
      11'h53F: dout <= 8'b11111111; // 1343 : 255 - 0xff
      11'h540: dout <= 8'b11111111; // 1344 : 255 - 0xff -- Background 0xa8
      11'h541: dout <= 8'b11111111; // 1345 : 255 - 0xff
      11'h542: dout <= 8'b11111111; // 1346 : 255 - 0xff
      11'h543: dout <= 8'b11111111; // 1347 : 255 - 0xff
      11'h544: dout <= 8'b11111111; // 1348 : 255 - 0xff
      11'h545: dout <= 8'b11111111; // 1349 : 255 - 0xff
      11'h546: dout <= 8'b11111111; // 1350 : 255 - 0xff
      11'h547: dout <= 8'b11111111; // 1351 : 255 - 0xff
      11'h548: dout <= 8'b11111111; // 1352 : 255 - 0xff -- Background 0xa9
      11'h549: dout <= 8'b11111111; // 1353 : 255 - 0xff
      11'h54A: dout <= 8'b11111111; // 1354 : 255 - 0xff
      11'h54B: dout <= 8'b11111111; // 1355 : 255 - 0xff
      11'h54C: dout <= 8'b11111111; // 1356 : 255 - 0xff
      11'h54D: dout <= 8'b11111111; // 1357 : 255 - 0xff
      11'h54E: dout <= 8'b11111111; // 1358 : 255 - 0xff
      11'h54F: dout <= 8'b11111111; // 1359 : 255 - 0xff
      11'h550: dout <= 8'b11111111; // 1360 : 255 - 0xff -- Background 0xaa
      11'h551: dout <= 8'b11111111; // 1361 : 255 - 0xff
      11'h552: dout <= 8'b00001111; // 1362 :  15 - 0xf
      11'h553: dout <= 8'b00000111; // 1363 :   7 - 0x7
      11'h554: dout <= 8'b00000011; // 1364 :   3 - 0x3
      11'h555: dout <= 8'b00000001; // 1365 :   1 - 0x1
      11'h556: dout <= 8'b00000001; // 1366 :   1 - 0x1
      11'h557: dout <= 8'b00000000; // 1367 :   0 - 0x0
      11'h558: dout <= 8'b00000000; // 1368 :   0 - 0x0 -- Background 0xab
      11'h559: dout <= 8'b00000000; // 1369 :   0 - 0x0
      11'h55A: dout <= 8'b00000000; // 1370 :   0 - 0x0
      11'h55B: dout <= 8'b00000000; // 1371 :   0 - 0x0
      11'h55C: dout <= 8'b10000000; // 1372 : 128 - 0x80
      11'h55D: dout <= 8'b11000000; // 1373 : 192 - 0xc0
      11'h55E: dout <= 8'b11111100; // 1374 : 252 - 0xfc
      11'h55F: dout <= 8'b11111110; // 1375 : 254 - 0xfe
      11'h560: dout <= 8'b11111111; // 1376 : 255 - 0xff -- Background 0xac
      11'h561: dout <= 8'b11111111; // 1377 : 255 - 0xff
      11'h562: dout <= 8'b11111111; // 1378 : 255 - 0xff
      11'h563: dout <= 8'b11111111; // 1379 : 255 - 0xff
      11'h564: dout <= 8'b11111111; // 1380 : 255 - 0xff
      11'h565: dout <= 8'b11111111; // 1381 : 255 - 0xff
      11'h566: dout <= 8'b10111111; // 1382 : 191 - 0xbf
      11'h567: dout <= 8'b10011111; // 1383 : 159 - 0x9f
      11'h568: dout <= 8'b11001111; // 1384 : 207 - 0xcf -- Background 0xad
      11'h569: dout <= 8'b11111111; // 1385 : 255 - 0xff
      11'h56A: dout <= 8'b11111111; // 1386 : 255 - 0xff
      11'h56B: dout <= 8'b11111111; // 1387 : 255 - 0xff
      11'h56C: dout <= 8'b11111111; // 1388 : 255 - 0xff
      11'h56D: dout <= 8'b11111111; // 1389 : 255 - 0xff
      11'h56E: dout <= 8'b11111111; // 1390 : 255 - 0xff
      11'h56F: dout <= 8'b11111111; // 1391 : 255 - 0xff
      11'h570: dout <= 8'b11111111; // 1392 : 255 - 0xff -- Background 0xae
      11'h571: dout <= 8'b11111111; // 1393 : 255 - 0xff
      11'h572: dout <= 8'b11111111; // 1394 : 255 - 0xff
      11'h573: dout <= 8'b11111111; // 1395 : 255 - 0xff
      11'h574: dout <= 8'b11111111; // 1396 : 255 - 0xff
      11'h575: dout <= 8'b11111111; // 1397 : 255 - 0xff
      11'h576: dout <= 8'b11111111; // 1398 : 255 - 0xff
      11'h577: dout <= 8'b11111111; // 1399 : 255 - 0xff
      11'h578: dout <= 8'b00000000; // 1400 :   0 - 0x0 -- Background 0xaf
      11'h579: dout <= 8'b10000000; // 1401 : 128 - 0x80
      11'h57A: dout <= 8'b11000000; // 1402 : 192 - 0xc0
      11'h57B: dout <= 8'b11100000; // 1403 : 224 - 0xe0
      11'h57C: dout <= 8'b11100000; // 1404 : 224 - 0xe0
      11'h57D: dout <= 8'b11100000; // 1405 : 224 - 0xe0
      11'h57E: dout <= 8'b11110000; // 1406 : 240 - 0xf0
      11'h57F: dout <= 8'b11110000; // 1407 : 240 - 0xf0
      11'h580: dout <= 8'b11110000; // 1408 : 240 - 0xf0 -- Background 0xb0
      11'h581: dout <= 8'b11110000; // 1409 : 240 - 0xf0
      11'h582: dout <= 8'b11100000; // 1410 : 224 - 0xe0
      11'h583: dout <= 8'b11100000; // 1411 : 224 - 0xe0
      11'h584: dout <= 8'b11100000; // 1412 : 224 - 0xe0
      11'h585: dout <= 8'b11000000; // 1413 : 192 - 0xc0
      11'h586: dout <= 8'b11000000; // 1414 : 192 - 0xc0
      11'h587: dout <= 8'b10000000; // 1415 : 128 - 0x80
      11'h588: dout <= 8'b10000000; // 1416 : 128 - 0x80 -- Background 0xb1
      11'h589: dout <= 8'b10000000; // 1417 : 128 - 0x80
      11'h58A: dout <= 8'b10000000; // 1418 : 128 - 0x80
      11'h58B: dout <= 8'b00000000; // 1419 :   0 - 0x0
      11'h58C: dout <= 8'b00000000; // 1420 :   0 - 0x0
      11'h58D: dout <= 8'b11000000; // 1421 : 192 - 0xc0
      11'h58E: dout <= 8'b11100000; // 1422 : 224 - 0xe0
      11'h58F: dout <= 8'b11110000; // 1423 : 240 - 0xf0
      11'h590: dout <= 8'b00000000; // 1424 :   0 - 0x0 -- Background 0xb2
      11'h591: dout <= 8'b00000000; // 1425 :   0 - 0x0
      11'h592: dout <= 8'b00000001; // 1426 :   1 - 0x1
      11'h593: dout <= 8'b00000011; // 1427 :   3 - 0x3
      11'h594: dout <= 8'b00000111; // 1428 :   7 - 0x7
      11'h595: dout <= 8'b00000111; // 1429 :   7 - 0x7
      11'h596: dout <= 8'b00000111; // 1430 :   7 - 0x7
      11'h597: dout <= 8'b00000111; // 1431 :   7 - 0x7
      11'h598: dout <= 8'b00000011; // 1432 :   3 - 0x3 -- Background 0xb3
      11'h599: dout <= 8'b00000001; // 1433 :   1 - 0x1
      11'h59A: dout <= 8'b00000000; // 1434 :   0 - 0x0
      11'h59B: dout <= 8'b00000000; // 1435 :   0 - 0x0
      11'h59C: dout <= 8'b00000000; // 1436 :   0 - 0x0
      11'h59D: dout <= 8'b00000001; // 1437 :   1 - 0x1
      11'h59E: dout <= 8'b00000011; // 1438 :   3 - 0x3
      11'h59F: dout <= 8'b00000011; // 1439 :   3 - 0x3
      11'h5A0: dout <= 8'b00000011; // 1440 :   3 - 0x3 -- Background 0xb4
      11'h5A1: dout <= 8'b00000011; // 1441 :   3 - 0x3
      11'h5A2: dout <= 8'b00000111; // 1442 :   7 - 0x7
      11'h5A3: dout <= 8'b00011111; // 1443 :  31 - 0x1f
      11'h5A4: dout <= 8'b00111111; // 1444 :  63 - 0x3f
      11'h5A5: dout <= 8'b00111111; // 1445 :  63 - 0x3f
      11'h5A6: dout <= 8'b00000000; // 1446 :   0 - 0x0
      11'h5A7: dout <= 8'b00000000; // 1447 :   0 - 0x0
      11'h5A8: dout <= 8'b00000000; // 1448 :   0 - 0x0 -- Background 0xb5
      11'h5A9: dout <= 8'b00000000; // 1449 :   0 - 0x0
      11'h5AA: dout <= 8'b00000000; // 1450 :   0 - 0x0
      11'h5AB: dout <= 8'b00000000; // 1451 :   0 - 0x0
      11'h5AC: dout <= 8'b00000001; // 1452 :   1 - 0x1
      11'h5AD: dout <= 8'b00000011; // 1453 :   3 - 0x3
      11'h5AE: dout <= 8'b00000011; // 1454 :   3 - 0x3
      11'h5AF: dout <= 8'b00001111; // 1455 :  15 - 0xf
      11'h5B0: dout <= 8'b00111111; // 1456 :  63 - 0x3f -- Background 0xb6
      11'h5B1: dout <= 8'b01111111; // 1457 : 127 - 0x7f
      11'h5B2: dout <= 8'b11111111; // 1458 : 255 - 0xff
      11'h5B3: dout <= 8'b11111111; // 1459 : 255 - 0xff
      11'h5B4: dout <= 8'b11111111; // 1460 : 255 - 0xff
      11'h5B5: dout <= 8'b11111111; // 1461 : 255 - 0xff
      11'h5B6: dout <= 8'b11111111; // 1462 : 255 - 0xff
      11'h5B7: dout <= 8'b11111111; // 1463 : 255 - 0xff
      11'h5B8: dout <= 8'b11111111; // 1464 : 255 - 0xff -- Background 0xb7
      11'h5B9: dout <= 8'b11111111; // 1465 : 255 - 0xff
      11'h5BA: dout <= 8'b11111111; // 1466 : 255 - 0xff
      11'h5BB: dout <= 8'b00011111; // 1467 :  31 - 0x1f
      11'h5BC: dout <= 8'b01111111; // 1468 : 127 - 0x7f
      11'h5BD: dout <= 8'b11111111; // 1469 : 255 - 0xff
      11'h5BE: dout <= 8'b11111111; // 1470 : 255 - 0xff
      11'h5BF: dout <= 8'b11111111; // 1471 : 255 - 0xff
      11'h5C0: dout <= 8'b11111111; // 1472 : 255 - 0xff -- Background 0xb8
      11'h5C1: dout <= 8'b11111111; // 1473 : 255 - 0xff
      11'h5C2: dout <= 8'b11111111; // 1474 : 255 - 0xff
      11'h5C3: dout <= 8'b11111100; // 1475 : 252 - 0xfc
      11'h5C4: dout <= 8'b11111000; // 1476 : 248 - 0xf8
      11'h5C5: dout <= 8'b11111000; // 1477 : 248 - 0xf8
      11'h5C6: dout <= 8'b00000000; // 1478 :   0 - 0x0
      11'h5C7: dout <= 8'b00000000; // 1479 :   0 - 0x0
      11'h5C8: dout <= 8'b11001111; // 1480 : 207 - 0xcf -- Background 0xb9
      11'h5C9: dout <= 8'b10001000; // 1481 : 136 - 0x88
      11'h5CA: dout <= 8'b11011101; // 1482 : 221 - 0xdd
      11'h5CB: dout <= 8'b11001000; // 1483 : 200 - 0xc8
      11'h5CC: dout <= 8'b11111000; // 1484 : 248 - 0xf8
      11'h5CD: dout <= 8'b11111111; // 1485 : 255 - 0xff
      11'h5CE: dout <= 8'b11111111; // 1486 : 255 - 0xff
      11'h5CF: dout <= 8'b11111111; // 1487 : 255 - 0xff
      11'h5D0: dout <= 8'b11111111; // 1488 : 255 - 0xff -- Background 0xba
      11'h5D1: dout <= 8'b11111111; // 1489 : 255 - 0xff
      11'h5D2: dout <= 8'b11000000; // 1490 : 192 - 0xc0
      11'h5D3: dout <= 8'b00000000; // 1491 :   0 - 0x0
      11'h5D4: dout <= 8'b00000000; // 1492 :   0 - 0x0
      11'h5D5: dout <= 8'b00000000; // 1493 :   0 - 0x0
      11'h5D6: dout <= 8'b00000000; // 1494 :   0 - 0x0
      11'h5D7: dout <= 8'b00000000; // 1495 :   0 - 0x0
      11'h5D8: dout <= 8'b11111001; // 1496 : 249 - 0xf9 -- Background 0xbb
      11'h5D9: dout <= 8'b10001000; // 1497 : 136 - 0x88
      11'h5DA: dout <= 8'b11011101; // 1498 : 221 - 0xdd
      11'h5DB: dout <= 8'b10001001; // 1499 : 137 - 0x89
      11'h5DC: dout <= 8'b00001111; // 1500 :  15 - 0xf
      11'h5DD: dout <= 8'b11111111; // 1501 : 255 - 0xff
      11'h5DE: dout <= 8'b11111111; // 1502 : 255 - 0xff
      11'h5DF: dout <= 8'b11111111; // 1503 : 255 - 0xff
      11'h5E0: dout <= 8'b00000011; // 1504 :   3 - 0x3 -- Background 0xbc
      11'h5E1: dout <= 8'b00000111; // 1505 :   7 - 0x7
      11'h5E2: dout <= 8'b00001111; // 1506 :  15 - 0xf
      11'h5E3: dout <= 8'b00000111; // 1507 :   7 - 0x7
      11'h5E4: dout <= 8'b10000111; // 1508 : 135 - 0x87
      11'h5E5: dout <= 8'b11000011; // 1509 : 195 - 0xc3
      11'h5E6: dout <= 8'b11100000; // 1510 : 224 - 0xe0
      11'h5E7: dout <= 8'b11111111; // 1511 : 255 - 0xff
      11'h5E8: dout <= 8'b11111111; // 1512 : 255 - 0xff -- Background 0xbd
      11'h5E9: dout <= 8'b11111111; // 1513 : 255 - 0xff
      11'h5EA: dout <= 8'b11111111; // 1514 : 255 - 0xff
      11'h5EB: dout <= 8'b11111111; // 1515 : 255 - 0xff
      11'h5EC: dout <= 8'b11111111; // 1516 : 255 - 0xff
      11'h5ED: dout <= 8'b11111111; // 1517 : 255 - 0xff
      11'h5EE: dout <= 8'b11111111; // 1518 : 255 - 0xff
      11'h5EF: dout <= 8'b11111110; // 1519 : 254 - 0xfe
      11'h5F0: dout <= 8'b11111100; // 1520 : 252 - 0xfc -- Background 0xbe
      11'h5F1: dout <= 8'b11111000; // 1521 : 248 - 0xf8
      11'h5F2: dout <= 8'b11111000; // 1522 : 248 - 0xf8
      11'h5F3: dout <= 8'b11111000; // 1523 : 248 - 0xf8
      11'h5F4: dout <= 8'b11111000; // 1524 : 248 - 0xf8
      11'h5F5: dout <= 8'b11111100; // 1525 : 252 - 0xfc
      11'h5F6: dout <= 8'b11111110; // 1526 : 254 - 0xfe
      11'h5F7: dout <= 8'b11111111; // 1527 : 255 - 0xff
      11'h5F8: dout <= 8'b11111111; // 1528 : 255 - 0xff -- Background 0xbf
      11'h5F9: dout <= 8'b11111111; // 1529 : 255 - 0xff
      11'h5FA: dout <= 8'b11111111; // 1530 : 255 - 0xff
      11'h5FB: dout <= 8'b11111111; // 1531 : 255 - 0xff
      11'h5FC: dout <= 8'b11111111; // 1532 : 255 - 0xff
      11'h5FD: dout <= 8'b11111111; // 1533 : 255 - 0xff
      11'h5FE: dout <= 8'b11111111; // 1534 : 255 - 0xff
      11'h5FF: dout <= 8'b11111111; // 1535 : 255 - 0xff
      11'h600: dout <= 8'b11000000; // 1536 : 192 - 0xc0 -- Background 0xc0
      11'h601: dout <= 8'b11110000; // 1537 : 240 - 0xf0
      11'h602: dout <= 8'b11111100; // 1538 : 252 - 0xfc
      11'h603: dout <= 8'b11111100; // 1539 : 252 - 0xfc
      11'h604: dout <= 8'b11111110; // 1540 : 254 - 0xfe
      11'h605: dout <= 8'b11111110; // 1541 : 254 - 0xfe
      11'h606: dout <= 8'b11111110; // 1542 : 254 - 0xfe
      11'h607: dout <= 8'b11111110; // 1543 : 254 - 0xfe
      11'h608: dout <= 8'b11111111; // 1544 : 255 - 0xff -- Background 0xc1
      11'h609: dout <= 8'b11111111; // 1545 : 255 - 0xff
      11'h60A: dout <= 8'b11111110; // 1546 : 254 - 0xfe
      11'h60B: dout <= 8'b11111100; // 1547 : 252 - 0xfc
      11'h60C: dout <= 8'b11110000; // 1548 : 240 - 0xf0
      11'h60D: dout <= 8'b11100000; // 1549 : 224 - 0xe0
      11'h60E: dout <= 8'b10000000; // 1550 : 128 - 0x80
      11'h60F: dout <= 8'b00000000; // 1551 :   0 - 0x0
      11'h610: dout <= 8'b00000011; // 1552 :   3 - 0x3 -- Background 0xc2
      11'h611: dout <= 8'b00001111; // 1553 :  15 - 0xf
      11'h612: dout <= 8'b00111111; // 1554 :  63 - 0x3f
      11'h613: dout <= 8'b00111111; // 1555 :  63 - 0x3f
      11'h614: dout <= 8'b01111111; // 1556 : 127 - 0x7f
      11'h615: dout <= 8'b01111111; // 1557 : 127 - 0x7f
      11'h616: dout <= 8'b01111110; // 1558 : 126 - 0x7e
      11'h617: dout <= 8'b11111111; // 1559 : 255 - 0xff
      11'h618: dout <= 8'b11111111; // 1560 : 255 - 0xff -- Background 0xc3
      11'h619: dout <= 8'b11111111; // 1561 : 255 - 0xff
      11'h61A: dout <= 8'b01111111; // 1562 : 127 - 0x7f
      11'h61B: dout <= 8'b00111111; // 1563 :  63 - 0x3f
      11'h61C: dout <= 8'b00001111; // 1564 :  15 - 0xf
      11'h61D: dout <= 8'b00000111; // 1565 :   7 - 0x7
      11'h61E: dout <= 8'b00000001; // 1566 :   1 - 0x1
      11'h61F: dout <= 8'b00000000; // 1567 :   0 - 0x0
      11'h620: dout <= 8'b11000000; // 1568 : 192 - 0xc0 -- Background 0xc4
      11'h621: dout <= 8'b11100000; // 1569 : 224 - 0xe0
      11'h622: dout <= 8'b11110000; // 1570 : 240 - 0xf0
      11'h623: dout <= 8'b11100000; // 1571 : 224 - 0xe0
      11'h624: dout <= 8'b11100001; // 1572 : 225 - 0xe1
      11'h625: dout <= 8'b11000011; // 1573 : 195 - 0xc3
      11'h626: dout <= 8'b00000111; // 1574 :   7 - 0x7
      11'h627: dout <= 8'b11111111; // 1575 : 255 - 0xff
      11'h628: dout <= 8'b11111111; // 1576 : 255 - 0xff -- Background 0xc5
      11'h629: dout <= 8'b11111111; // 1577 : 255 - 0xff
      11'h62A: dout <= 8'b11111111; // 1578 : 255 - 0xff
      11'h62B: dout <= 8'b11111111; // 1579 : 255 - 0xff
      11'h62C: dout <= 8'b11111111; // 1580 : 255 - 0xff
      11'h62D: dout <= 8'b11111111; // 1581 : 255 - 0xff
      11'h62E: dout <= 8'b11111111; // 1582 : 255 - 0xff
      11'h62F: dout <= 8'b01111111; // 1583 : 127 - 0x7f
      11'h630: dout <= 8'b00111111; // 1584 :  63 - 0x3f -- Background 0xc6
      11'h631: dout <= 8'b00011111; // 1585 :  31 - 0x1f
      11'h632: dout <= 8'b00011111; // 1586 :  31 - 0x1f
      11'h633: dout <= 8'b00011111; // 1587 :  31 - 0x1f
      11'h634: dout <= 8'b00011111; // 1588 :  31 - 0x1f
      11'h635: dout <= 8'b00111111; // 1589 :  63 - 0x3f
      11'h636: dout <= 8'b01111111; // 1590 : 127 - 0x7f
      11'h637: dout <= 8'b11111111; // 1591 : 255 - 0xff
      11'h638: dout <= 8'b11111111; // 1592 : 255 - 0xff -- Background 0xc7
      11'h639: dout <= 8'b11111111; // 1593 : 255 - 0xff
      11'h63A: dout <= 8'b11111111; // 1594 : 255 - 0xff
      11'h63B: dout <= 8'b11111111; // 1595 : 255 - 0xff
      11'h63C: dout <= 8'b11111111; // 1596 : 255 - 0xff
      11'h63D: dout <= 8'b11111111; // 1597 : 255 - 0xff
      11'h63E: dout <= 8'b11111111; // 1598 : 255 - 0xff
      11'h63F: dout <= 8'b11111111; // 1599 : 255 - 0xff
      11'h640: dout <= 8'b11111111; // 1600 : 255 - 0xff -- Background 0xc8
      11'h641: dout <= 8'b11111111; // 1601 : 255 - 0xff
      11'h642: dout <= 8'b00000011; // 1602 :   3 - 0x3
      11'h643: dout <= 8'b00000000; // 1603 :   0 - 0x0
      11'h644: dout <= 8'b00000000; // 1604 :   0 - 0x0
      11'h645: dout <= 8'b00000000; // 1605 :   0 - 0x0
      11'h646: dout <= 8'b00000000; // 1606 :   0 - 0x0
      11'h647: dout <= 8'b00000000; // 1607 :   0 - 0x0
      11'h648: dout <= 8'b00000000; // 1608 :   0 - 0x0 -- Background 0xc9
      11'h649: dout <= 8'b00000000; // 1609 :   0 - 0x0
      11'h64A: dout <= 8'b00000000; // 1610 :   0 - 0x0
      11'h64B: dout <= 8'b00000000; // 1611 :   0 - 0x0
      11'h64C: dout <= 8'b10000000; // 1612 : 128 - 0x80
      11'h64D: dout <= 8'b11000000; // 1613 : 192 - 0xc0
      11'h64E: dout <= 8'b11000000; // 1614 : 192 - 0xc0
      11'h64F: dout <= 8'b11110000; // 1615 : 240 - 0xf0
      11'h650: dout <= 8'b11111100; // 1616 : 252 - 0xfc -- Background 0xca
      11'h651: dout <= 8'b11111110; // 1617 : 254 - 0xfe
      11'h652: dout <= 8'b11111111; // 1618 : 255 - 0xff
      11'h653: dout <= 8'b11111111; // 1619 : 255 - 0xff
      11'h654: dout <= 8'b11111111; // 1620 : 255 - 0xff
      11'h655: dout <= 8'b11111111; // 1621 : 255 - 0xff
      11'h656: dout <= 8'b11111111; // 1622 : 255 - 0xff
      11'h657: dout <= 8'b11111111; // 1623 : 255 - 0xff
      11'h658: dout <= 8'b11111111; // 1624 : 255 - 0xff -- Background 0xcb
      11'h659: dout <= 8'b11111111; // 1625 : 255 - 0xff
      11'h65A: dout <= 8'b11111111; // 1626 : 255 - 0xff
      11'h65B: dout <= 8'b11111000; // 1627 : 248 - 0xf8
      11'h65C: dout <= 8'b11111110; // 1628 : 254 - 0xfe
      11'h65D: dout <= 8'b11111111; // 1629 : 255 - 0xff
      11'h65E: dout <= 8'b11111111; // 1630 : 255 - 0xff
      11'h65F: dout <= 8'b11111111; // 1631 : 255 - 0xff
      11'h660: dout <= 8'b11111111; // 1632 : 255 - 0xff -- Background 0xcc
      11'h661: dout <= 8'b11111111; // 1633 : 255 - 0xff
      11'h662: dout <= 8'b11111111; // 1634 : 255 - 0xff
      11'h663: dout <= 8'b00111111; // 1635 :  63 - 0x3f
      11'h664: dout <= 8'b00011111; // 1636 :  31 - 0x1f
      11'h665: dout <= 8'b00011111; // 1637 :  31 - 0x1f
      11'h666: dout <= 8'b00000000; // 1638 :   0 - 0x0
      11'h667: dout <= 8'b00000000; // 1639 :   0 - 0x0
      11'h668: dout <= 8'b00000000; // 1640 :   0 - 0x0 -- Background 0xcd
      11'h669: dout <= 8'b00000000; // 1641 :   0 - 0x0
      11'h66A: dout <= 8'b10000000; // 1642 : 128 - 0x80
      11'h66B: dout <= 8'b11000000; // 1643 : 192 - 0xc0
      11'h66C: dout <= 8'b11100000; // 1644 : 224 - 0xe0
      11'h66D: dout <= 8'b11100000; // 1645 : 224 - 0xe0
      11'h66E: dout <= 8'b11100000; // 1646 : 224 - 0xe0
      11'h66F: dout <= 8'b11100000; // 1647 : 224 - 0xe0
      11'h670: dout <= 8'b11000000; // 1648 : 192 - 0xc0 -- Background 0xce
      11'h671: dout <= 8'b10000000; // 1649 : 128 - 0x80
      11'h672: dout <= 8'b00000000; // 1650 :   0 - 0x0
      11'h673: dout <= 8'b00000000; // 1651 :   0 - 0x0
      11'h674: dout <= 8'b00000000; // 1652 :   0 - 0x0
      11'h675: dout <= 8'b10000000; // 1653 : 128 - 0x80
      11'h676: dout <= 8'b11000000; // 1654 : 192 - 0xc0
      11'h677: dout <= 8'b11000000; // 1655 : 192 - 0xc0
      11'h678: dout <= 8'b11000000; // 1656 : 192 - 0xc0 -- Background 0xcf
      11'h679: dout <= 8'b11000000; // 1657 : 192 - 0xc0
      11'h67A: dout <= 8'b11100000; // 1658 : 224 - 0xe0
      11'h67B: dout <= 8'b11111000; // 1659 : 248 - 0xf8
      11'h67C: dout <= 8'b11111100; // 1660 : 252 - 0xfc
      11'h67D: dout <= 8'b11111100; // 1661 : 252 - 0xfc
      11'h67E: dout <= 8'b00000000; // 1662 :   0 - 0x0
      11'h67F: dout <= 8'b00000000; // 1663 :   0 - 0x0
      11'h680: dout <= 8'b00000000; // 1664 :   0 - 0x0 -- Background 0xd0
      11'h681: dout <= 8'b00000000; // 1665 :   0 - 0x0
      11'h682: dout <= 8'b00000000; // 1666 :   0 - 0x0
      11'h683: dout <= 8'b00000000; // 1667 :   0 - 0x0
      11'h684: dout <= 8'b00000000; // 1668 :   0 - 0x0
      11'h685: dout <= 8'b00000000; // 1669 :   0 - 0x0
      11'h686: dout <= 8'b00000000; // 1670 :   0 - 0x0
      11'h687: dout <= 8'b00000000; // 1671 :   0 - 0x0
      11'h688: dout <= 8'b00000000; // 1672 :   0 - 0x0 -- Background 0xd1
      11'h689: dout <= 8'b00000000; // 1673 :   0 - 0x0
      11'h68A: dout <= 8'b00000000; // 1674 :   0 - 0x0
      11'h68B: dout <= 8'b00000000; // 1675 :   0 - 0x0
      11'h68C: dout <= 8'b00000000; // 1676 :   0 - 0x0
      11'h68D: dout <= 8'b00000000; // 1677 :   0 - 0x0
      11'h68E: dout <= 8'b00000000; // 1678 :   0 - 0x0
      11'h68F: dout <= 8'b00000000; // 1679 :   0 - 0x0
      11'h690: dout <= 8'b00000000; // 1680 :   0 - 0x0 -- Background 0xd2
      11'h691: dout <= 8'b00000000; // 1681 :   0 - 0x0
      11'h692: dout <= 8'b00000000; // 1682 :   0 - 0x0
      11'h693: dout <= 8'b00000000; // 1683 :   0 - 0x0
      11'h694: dout <= 8'b00000000; // 1684 :   0 - 0x0
      11'h695: dout <= 8'b00000000; // 1685 :   0 - 0x0
      11'h696: dout <= 8'b00000000; // 1686 :   0 - 0x0
      11'h697: dout <= 8'b00000000; // 1687 :   0 - 0x0
      11'h698: dout <= 8'b00000000; // 1688 :   0 - 0x0 -- Background 0xd3
      11'h699: dout <= 8'b00000000; // 1689 :   0 - 0x0
      11'h69A: dout <= 8'b00000000; // 1690 :   0 - 0x0
      11'h69B: dout <= 8'b00000000; // 1691 :   0 - 0x0
      11'h69C: dout <= 8'b00000000; // 1692 :   0 - 0x0
      11'h69D: dout <= 8'b00000000; // 1693 :   0 - 0x0
      11'h69E: dout <= 8'b00000000; // 1694 :   0 - 0x0
      11'h69F: dout <= 8'b00000000; // 1695 :   0 - 0x0
      11'h6A0: dout <= 8'b00000000; // 1696 :   0 - 0x0 -- Background 0xd4
      11'h6A1: dout <= 8'b00000000; // 1697 :   0 - 0x0
      11'h6A2: dout <= 8'b00000000; // 1698 :   0 - 0x0
      11'h6A3: dout <= 8'b00000000; // 1699 :   0 - 0x0
      11'h6A4: dout <= 8'b00000011; // 1700 :   3 - 0x3
      11'h6A5: dout <= 8'b00000111; // 1701 :   7 - 0x7
      11'h6A6: dout <= 8'b00000011; // 1702 :   3 - 0x3
      11'h6A7: dout <= 8'b00000111; // 1703 :   7 - 0x7
      11'h6A8: dout <= 8'b00011111; // 1704 :  31 - 0x1f -- Background 0xd5
      11'h6A9: dout <= 8'b00111111; // 1705 :  63 - 0x3f
      11'h6AA: dout <= 8'b01111111; // 1706 : 127 - 0x7f
      11'h6AB: dout <= 8'b11111111; // 1707 : 255 - 0xff
      11'h6AC: dout <= 8'b11111111; // 1708 : 255 - 0xff
      11'h6AD: dout <= 8'b11111111; // 1709 : 255 - 0xff
      11'h6AE: dout <= 8'b11111111; // 1710 : 255 - 0xff
      11'h6AF: dout <= 8'b01111111; // 1711 : 127 - 0x7f
      11'h6B0: dout <= 8'b00000000; // 1712 :   0 - 0x0 -- Background 0xd6
      11'h6B1: dout <= 8'b00000000; // 1713 :   0 - 0x0
      11'h6B2: dout <= 8'b00000000; // 1714 :   0 - 0x0
      11'h6B3: dout <= 8'b11000000; // 1715 : 192 - 0xc0
      11'h6B4: dout <= 8'b11100000; // 1716 : 224 - 0xe0
      11'h6B5: dout <= 8'b11110000; // 1717 : 240 - 0xf0
      11'h6B6: dout <= 8'b11110000; // 1718 : 240 - 0xf0
      11'h6B7: dout <= 8'b11111000; // 1719 : 248 - 0xf8
      11'h6B8: dout <= 8'b11111100; // 1720 : 252 - 0xfc -- Background 0xd7
      11'h6B9: dout <= 8'b11111000; // 1721 : 248 - 0xf8
      11'h6BA: dout <= 8'b11110000; // 1722 : 240 - 0xf0
      11'h6BB: dout <= 8'b11111111; // 1723 : 255 - 0xff
      11'h6BC: dout <= 8'b11111111; // 1724 : 255 - 0xff
      11'h6BD: dout <= 8'b11111111; // 1725 : 255 - 0xff
      11'h6BE: dout <= 8'b11111111; // 1726 : 255 - 0xff
      11'h6BF: dout <= 8'b11111111; // 1727 : 255 - 0xff
      11'h6C0: dout <= 8'b00000000; // 1728 :   0 - 0x0 -- Background 0xd8
      11'h6C1: dout <= 8'b00000000; // 1729 :   0 - 0x0
      11'h6C2: dout <= 8'b00000000; // 1730 :   0 - 0x0
      11'h6C3: dout <= 8'b00000000; // 1731 :   0 - 0x0
      11'h6C4: dout <= 8'b00000011; // 1732 :   3 - 0x3
      11'h6C5: dout <= 8'b00000111; // 1733 :   7 - 0x7
      11'h6C6: dout <= 8'b00001111; // 1734 :  15 - 0xf
      11'h6C7: dout <= 8'b00011111; // 1735 :  31 - 0x1f
      11'h6C8: dout <= 8'b00111111; // 1736 :  63 - 0x3f -- Background 0xd9
      11'h6C9: dout <= 8'b00011111; // 1737 :  31 - 0x1f
      11'h6CA: dout <= 8'b00000111; // 1738 :   7 - 0x7
      11'h6CB: dout <= 8'b11111111; // 1739 : 255 - 0xff
      11'h6CC: dout <= 8'b11111111; // 1740 : 255 - 0xff
      11'h6CD: dout <= 8'b11111111; // 1741 : 255 - 0xff
      11'h6CE: dout <= 8'b11111111; // 1742 : 255 - 0xff
      11'h6CF: dout <= 8'b11111111; // 1743 : 255 - 0xff
      11'h6D0: dout <= 8'b00000000; // 1744 :   0 - 0x0 -- Background 0xda
      11'h6D1: dout <= 8'b00000000; // 1745 :   0 - 0x0
      11'h6D2: dout <= 8'b00000000; // 1746 :   0 - 0x0
      11'h6D3: dout <= 8'b11000000; // 1747 : 192 - 0xc0
      11'h6D4: dout <= 8'b11000000; // 1748 : 192 - 0xc0
      11'h6D5: dout <= 8'b11000000; // 1749 : 192 - 0xc0
      11'h6D6: dout <= 8'b11100000; // 1750 : 224 - 0xe0
      11'h6D7: dout <= 8'b11111000; // 1751 : 248 - 0xf8
      11'h6D8: dout <= 8'b11111100; // 1752 : 252 - 0xfc -- Background 0xdb
      11'h6D9: dout <= 8'b11111110; // 1753 : 254 - 0xfe
      11'h6DA: dout <= 8'b11111110; // 1754 : 254 - 0xfe
      11'h6DB: dout <= 8'b11111111; // 1755 : 255 - 0xff
      11'h6DC: dout <= 8'b11111111; // 1756 : 255 - 0xff
      11'h6DD: dout <= 8'b11111111; // 1757 : 255 - 0xff
      11'h6DE: dout <= 8'b11111111; // 1758 : 255 - 0xff
      11'h6DF: dout <= 8'b11111110; // 1759 : 254 - 0xfe
      11'h6E0: dout <= 8'b00110110; // 1760 :  54 - 0x36 -- Background 0xdc
      11'h6E1: dout <= 8'b00110110; // 1761 :  54 - 0x36
      11'h6E2: dout <= 8'b01111110; // 1762 : 126 - 0x7e
      11'h6E3: dout <= 8'b01111111; // 1763 : 127 - 0x7f
      11'h6E4: dout <= 8'b01111111; // 1764 : 127 - 0x7f
      11'h6E5: dout <= 8'b01111111; // 1765 : 127 - 0x7f
      11'h6E6: dout <= 8'b00111111; // 1766 :  63 - 0x3f
      11'h6E7: dout <= 8'b00111111; // 1767 :  63 - 0x3f
      11'h6E8: dout <= 8'b00111111; // 1768 :  63 - 0x3f -- Background 0xdd
      11'h6E9: dout <= 8'b00011111; // 1769 :  31 - 0x1f
      11'h6EA: dout <= 8'b00011111; // 1770 :  31 - 0x1f
      11'h6EB: dout <= 8'b00001111; // 1771 :  15 - 0xf
      11'h6EC: dout <= 8'b00000111; // 1772 :   7 - 0x7
      11'h6ED: dout <= 8'b00000011; // 1773 :   3 - 0x3
      11'h6EE: dout <= 8'b00000000; // 1774 :   0 - 0x0
      11'h6EF: dout <= 8'b00000000; // 1775 :   0 - 0x0
      11'h6F0: dout <= 8'b00111111; // 1776 :  63 - 0x3f -- Background 0xde
      11'h6F1: dout <= 8'b00011111; // 1777 :  31 - 0x1f
      11'h6F2: dout <= 8'b11011111; // 1778 : 223 - 0xdf
      11'h6F3: dout <= 8'b11001111; // 1779 : 207 - 0xcf
      11'h6F4: dout <= 8'b11001111; // 1780 : 207 - 0xcf
      11'h6F5: dout <= 8'b10011111; // 1781 : 159 - 0x9f
      11'h6F6: dout <= 8'b11011111; // 1782 : 223 - 0xdf
      11'h6F7: dout <= 8'b11111111; // 1783 : 255 - 0xff
      11'h6F8: dout <= 8'b11111111; // 1784 : 255 - 0xff -- Background 0xdf
      11'h6F9: dout <= 8'b11111111; // 1785 : 255 - 0xff
      11'h6FA: dout <= 8'b11111111; // 1786 : 255 - 0xff
      11'h6FB: dout <= 8'b11111111; // 1787 : 255 - 0xff
      11'h6FC: dout <= 8'b11111111; // 1788 : 255 - 0xff
      11'h6FD: dout <= 8'b11111111; // 1789 : 255 - 0xff
      11'h6FE: dout <= 8'b11111111; // 1790 : 255 - 0xff
      11'h6FF: dout <= 8'b00001111; // 1791 :  15 - 0xf
      11'h700: dout <= 8'b11111111; // 1792 : 255 - 0xff -- Background 0xe0
      11'h701: dout <= 8'b11111111; // 1793 : 255 - 0xff
      11'h702: dout <= 8'b11111111; // 1794 : 255 - 0xff
      11'h703: dout <= 8'b11111111; // 1795 : 255 - 0xff
      11'h704: dout <= 8'b11111111; // 1796 : 255 - 0xff
      11'h705: dout <= 8'b11111111; // 1797 : 255 - 0xff
      11'h706: dout <= 8'b11111111; // 1798 : 255 - 0xff
      11'h707: dout <= 8'b11111111; // 1799 : 255 - 0xff
      11'h708: dout <= 8'b11111111; // 1800 : 255 - 0xff -- Background 0xe1
      11'h709: dout <= 8'b11111001; // 1801 : 249 - 0xf9
      11'h70A: dout <= 8'b11110000; // 1802 : 240 - 0xf0
      11'h70B: dout <= 8'b11110000; // 1803 : 240 - 0xf0
      11'h70C: dout <= 8'b10110001; // 1804 : 177 - 0xb1
      11'h70D: dout <= 8'b11011111; // 1805 : 223 - 0xdf
      11'h70E: dout <= 8'b11101111; // 1806 : 239 - 0xef
      11'h70F: dout <= 8'b10000111; // 1807 : 135 - 0x87
      11'h710: dout <= 8'b11111111; // 1808 : 255 - 0xff -- Background 0xe2
      11'h711: dout <= 8'b11111111; // 1809 : 255 - 0xff
      11'h712: dout <= 8'b11111111; // 1810 : 255 - 0xff
      11'h713: dout <= 8'b11111111; // 1811 : 255 - 0xff
      11'h714: dout <= 8'b11111111; // 1812 : 255 - 0xff
      11'h715: dout <= 8'b11111111; // 1813 : 255 - 0xff
      11'h716: dout <= 8'b11111111; // 1814 : 255 - 0xff
      11'h717: dout <= 8'b11111111; // 1815 : 255 - 0xff
      11'h718: dout <= 8'b11111111; // 1816 : 255 - 0xff -- Background 0xe3
      11'h719: dout <= 8'b11001111; // 1817 : 207 - 0xcf
      11'h71A: dout <= 8'b10000111; // 1818 : 135 - 0x87
      11'h71B: dout <= 8'b10000111; // 1819 : 135 - 0x87
      11'h71C: dout <= 8'b11001110; // 1820 : 206 - 0xce
      11'h71D: dout <= 8'b11111101; // 1821 : 253 - 0xfd
      11'h71E: dout <= 8'b11111011; // 1822 : 251 - 0xfb
      11'h71F: dout <= 8'b11110000; // 1823 : 240 - 0xf0
      11'h720: dout <= 8'b11111110; // 1824 : 254 - 0xfe -- Background 0xe4
      11'h721: dout <= 8'b11111100; // 1825 : 252 - 0xfc
      11'h722: dout <= 8'b11111100; // 1826 : 252 - 0xfc
      11'h723: dout <= 8'b11111000; // 1827 : 248 - 0xf8
      11'h724: dout <= 8'b11111011; // 1828 : 251 - 0xfb
      11'h725: dout <= 8'b11111101; // 1829 : 253 - 0xfd
      11'h726: dout <= 8'b11111110; // 1830 : 254 - 0xfe
      11'h727: dout <= 8'b11111111; // 1831 : 255 - 0xff
      11'h728: dout <= 8'b11111111; // 1832 : 255 - 0xff -- Background 0xe5
      11'h729: dout <= 8'b11111111; // 1833 : 255 - 0xff
      11'h72A: dout <= 8'b11111111; // 1834 : 255 - 0xff
      11'h72B: dout <= 8'b11111111; // 1835 : 255 - 0xff
      11'h72C: dout <= 8'b11111111; // 1836 : 255 - 0xff
      11'h72D: dout <= 8'b11111111; // 1837 : 255 - 0xff
      11'h72E: dout <= 8'b11111111; // 1838 : 255 - 0xff
      11'h72F: dout <= 8'b11111001; // 1839 : 249 - 0xf9
      11'h730: dout <= 8'b00000000; // 1840 :   0 - 0x0 -- Background 0xe6
      11'h731: dout <= 8'b00000000; // 1841 :   0 - 0x0
      11'h732: dout <= 8'b00000000; // 1842 :   0 - 0x0
      11'h733: dout <= 8'b01111000; // 1843 : 120 - 0x78
      11'h734: dout <= 8'b11111100; // 1844 : 252 - 0xfc
      11'h735: dout <= 8'b11111100; // 1845 : 252 - 0xfc
      11'h736: dout <= 8'b11111100; // 1846 : 252 - 0xfc
      11'h737: dout <= 8'b11111100; // 1847 : 252 - 0xfc
      11'h738: dout <= 8'b11111110; // 1848 : 254 - 0xfe -- Background 0xe7
      11'h739: dout <= 8'b11111110; // 1849 : 254 - 0xfe
      11'h73A: dout <= 8'b11111110; // 1850 : 254 - 0xfe
      11'h73B: dout <= 8'b11111110; // 1851 : 254 - 0xfe
      11'h73C: dout <= 8'b11111110; // 1852 : 254 - 0xfe
      11'h73D: dout <= 8'b11111100; // 1853 : 252 - 0xfc
      11'h73E: dout <= 8'b11111000; // 1854 : 248 - 0xf8
      11'h73F: dout <= 8'b11110000; // 1855 : 240 - 0xf0
      11'h740: dout <= 8'b00000000; // 1856 :   0 - 0x0 -- Background 0xe8
      11'h741: dout <= 8'b00000000; // 1857 :   0 - 0x0
      11'h742: dout <= 8'b00000000; // 1858 :   0 - 0x0
      11'h743: dout <= 8'b00000000; // 1859 :   0 - 0x0
      11'h744: dout <= 8'b00000000; // 1860 :   0 - 0x0
      11'h745: dout <= 8'b00000000; // 1861 :   0 - 0x0
      11'h746: dout <= 8'b00000000; // 1862 :   0 - 0x0
      11'h747: dout <= 8'b00000000; // 1863 :   0 - 0x0
      11'h748: dout <= 8'b00000001; // 1864 :   1 - 0x1 -- Background 0xe9
      11'h749: dout <= 8'b00001111; // 1865 :  15 - 0xf
      11'h74A: dout <= 8'b00011111; // 1866 :  31 - 0x1f
      11'h74B: dout <= 8'b00011111; // 1867 :  31 - 0x1f
      11'h74C: dout <= 8'b00111011; // 1868 :  59 - 0x3b
      11'h74D: dout <= 8'b00110011; // 1869 :  51 - 0x33
      11'h74E: dout <= 8'b00000001; // 1870 :   1 - 0x1
      11'h74F: dout <= 8'b00000001; // 1871 :   1 - 0x1
      11'h750: dout <= 8'b00000000; // 1872 :   0 - 0x0 -- Background 0xea
      11'h751: dout <= 8'b00000000; // 1873 :   0 - 0x0
      11'h752: dout <= 8'b00000000; // 1874 :   0 - 0x0
      11'h753: dout <= 8'b00110110; // 1875 :  54 - 0x36
      11'h754: dout <= 8'b01101100; // 1876 : 108 - 0x6c
      11'h755: dout <= 8'b11111101; // 1877 : 253 - 0xfd
      11'h756: dout <= 8'b11111111; // 1878 : 255 - 0xff
      11'h757: dout <= 8'b11111111; // 1879 : 255 - 0xff
      11'h758: dout <= 8'b11111111; // 1880 : 255 - 0xff -- Background 0xeb
      11'h759: dout <= 8'b01111111; // 1881 : 127 - 0x7f
      11'h75A: dout <= 8'b01111111; // 1882 : 127 - 0x7f
      11'h75B: dout <= 8'b01111111; // 1883 : 127 - 0x7f
      11'h75C: dout <= 8'b01111111; // 1884 : 127 - 0x7f
      11'h75D: dout <= 8'b00111111; // 1885 :  63 - 0x3f
      11'h75E: dout <= 8'b00011111; // 1886 :  31 - 0x1f
      11'h75F: dout <= 8'b00000111; // 1887 :   7 - 0x7
      11'h760: dout <= 8'b00000000; // 1888 :   0 - 0x0 -- Background 0xec
      11'h761: dout <= 8'b00000000; // 1889 :   0 - 0x0
      11'h762: dout <= 8'b00000000; // 1890 :   0 - 0x0
      11'h763: dout <= 8'b00000000; // 1891 :   0 - 0x0
      11'h764: dout <= 8'b00000000; // 1892 :   0 - 0x0
      11'h765: dout <= 8'b00000000; // 1893 :   0 - 0x0
      11'h766: dout <= 8'b00000000; // 1894 :   0 - 0x0
      11'h767: dout <= 8'b11100000; // 1895 : 224 - 0xe0
      11'h768: dout <= 8'b11111000; // 1896 : 248 - 0xf8 -- Background 0xed
      11'h769: dout <= 8'b11111111; // 1897 : 255 - 0xff
      11'h76A: dout <= 8'b11111111; // 1898 : 255 - 0xff
      11'h76B: dout <= 8'b11111111; // 1899 : 255 - 0xff
      11'h76C: dout <= 8'b11111111; // 1900 : 255 - 0xff
      11'h76D: dout <= 8'b11111111; // 1901 : 255 - 0xff
      11'h76E: dout <= 8'b11111111; // 1902 : 255 - 0xff
      11'h76F: dout <= 8'b11111111; // 1903 : 255 - 0xff
      11'h770: dout <= 8'b11111111; // 1904 : 255 - 0xff -- Background 0xee
      11'h771: dout <= 8'b01111111; // 1905 : 127 - 0x7f
      11'h772: dout <= 8'b00011111; // 1906 :  31 - 0x1f
      11'h773: dout <= 8'b00001111; // 1907 :  15 - 0xf
      11'h774: dout <= 8'b00001111; // 1908 :  15 - 0xf
      11'h775: dout <= 8'b10011111; // 1909 : 159 - 0x9f
      11'h776: dout <= 8'b10011111; // 1910 : 159 - 0x9f
      11'h777: dout <= 8'b10111111; // 1911 : 191 - 0xbf
      11'h778: dout <= 8'b01111111; // 1912 : 127 - 0x7f -- Background 0xef
      11'h779: dout <= 8'b11111111; // 1913 : 255 - 0xff
      11'h77A: dout <= 8'b11111111; // 1914 : 255 - 0xff
      11'h77B: dout <= 8'b11111111; // 1915 : 255 - 0xff
      11'h77C: dout <= 8'b11111111; // 1916 : 255 - 0xff
      11'h77D: dout <= 8'b11111111; // 1917 : 255 - 0xff
      11'h77E: dout <= 8'b11111111; // 1918 : 255 - 0xff
      11'h77F: dout <= 8'b11001111; // 1919 : 207 - 0xcf
      11'h780: dout <= 8'b00000000; // 1920 :   0 - 0x0 -- Background 0xf0
      11'h781: dout <= 8'b00000000; // 1921 :   0 - 0x0
      11'h782: dout <= 8'b11110000; // 1922 : 240 - 0xf0
      11'h783: dout <= 8'b11111111; // 1923 : 255 - 0xff
      11'h784: dout <= 8'b11111111; // 1924 : 255 - 0xff
      11'h785: dout <= 8'b11111111; // 1925 : 255 - 0xff
      11'h786: dout <= 8'b11111111; // 1926 : 255 - 0xff
      11'h787: dout <= 8'b11111111; // 1927 : 255 - 0xff
      11'h788: dout <= 8'b11111111; // 1928 : 255 - 0xff -- Background 0xf1
      11'h789: dout <= 8'b11111111; // 1929 : 255 - 0xff
      11'h78A: dout <= 8'b11111111; // 1930 : 255 - 0xff
      11'h78B: dout <= 8'b11110001; // 1931 : 241 - 0xf1
      11'h78C: dout <= 8'b11000100; // 1932 : 196 - 0xc4
      11'h78D: dout <= 8'b11101110; // 1933 : 238 - 0xee
      11'h78E: dout <= 8'b11000100; // 1934 : 196 - 0xc4
      11'h78F: dout <= 8'b10000011; // 1935 : 131 - 0x83
      11'h790: dout <= 8'b11000111; // 1936 : 199 - 0xc7 -- Background 0xf2
      11'h791: dout <= 8'b11111001; // 1937 : 249 - 0xf9
      11'h792: dout <= 8'b11110000; // 1938 : 240 - 0xf0
      11'h793: dout <= 8'b11110000; // 1939 : 240 - 0xf0
      11'h794: dout <= 8'b10110001; // 1940 : 177 - 0xb1
      11'h795: dout <= 8'b11011111; // 1941 : 223 - 0xdf
      11'h796: dout <= 8'b11101111; // 1942 : 239 - 0xef
      11'h797: dout <= 8'b10000111; // 1943 : 135 - 0x87
      11'h798: dout <= 8'b00000000; // 1944 :   0 - 0x0 -- Background 0xf3
      11'h799: dout <= 8'b00000000; // 1945 :   0 - 0x0
      11'h79A: dout <= 8'b00000111; // 1946 :   7 - 0x7
      11'h79B: dout <= 8'b11111111; // 1947 : 255 - 0xff
      11'h79C: dout <= 8'b11111111; // 1948 : 255 - 0xff
      11'h79D: dout <= 8'b11111111; // 1949 : 255 - 0xff
      11'h79E: dout <= 8'b11111111; // 1950 : 255 - 0xff
      11'h79F: dout <= 8'b11111111; // 1951 : 255 - 0xff
      11'h7A0: dout <= 8'b11111111; // 1952 : 255 - 0xff -- Background 0xf4
      11'h7A1: dout <= 8'b11111111; // 1953 : 255 - 0xff
      11'h7A2: dout <= 8'b11111111; // 1954 : 255 - 0xff
      11'h7A3: dout <= 8'b11000111; // 1955 : 199 - 0xc7
      11'h7A4: dout <= 8'b01000101; // 1956 :  69 - 0x45
      11'h7A5: dout <= 8'b11101110; // 1957 : 238 - 0xee
      11'h7A6: dout <= 8'b01000100; // 1958 :  68 - 0x44
      11'h7A7: dout <= 8'b11100001; // 1959 : 225 - 0xe1
      11'h7A8: dout <= 8'b11111111; // 1960 : 255 - 0xff -- Background 0xf5
      11'h7A9: dout <= 8'b11001111; // 1961 : 207 - 0xcf
      11'h7AA: dout <= 8'b10000111; // 1962 : 135 - 0x87
      11'h7AB: dout <= 8'b10000111; // 1963 : 135 - 0x87
      11'h7AC: dout <= 8'b11001110; // 1964 : 206 - 0xce
      11'h7AD: dout <= 8'b11111101; // 1965 : 253 - 0xfd
      11'h7AE: dout <= 8'b11111011; // 1966 : 251 - 0xfb
      11'h7AF: dout <= 8'b11110000; // 1967 : 240 - 0xf0
      11'h7B0: dout <= 8'b00000000; // 1968 :   0 - 0x0 -- Background 0xf6
      11'h7B1: dout <= 8'b00000000; // 1969 :   0 - 0x0
      11'h7B2: dout <= 8'b00000000; // 1970 :   0 - 0x0
      11'h7B3: dout <= 8'b00000000; // 1971 :   0 - 0x0
      11'h7B4: dout <= 8'b00000000; // 1972 :   0 - 0x0
      11'h7B5: dout <= 8'b00000001; // 1973 :   1 - 0x1
      11'h7B6: dout <= 8'b00000111; // 1974 :   7 - 0x7
      11'h7B7: dout <= 8'b00001111; // 1975 :  15 - 0xf
      11'h7B8: dout <= 8'b00111111; // 1976 :  63 - 0x3f -- Background 0xf7
      11'h7B9: dout <= 8'b11111111; // 1977 : 255 - 0xff
      11'h7BA: dout <= 8'b11111111; // 1978 : 255 - 0xff
      11'h7BB: dout <= 8'b11111111; // 1979 : 255 - 0xff
      11'h7BC: dout <= 8'b11111111; // 1980 : 255 - 0xff
      11'h7BD: dout <= 8'b11111111; // 1981 : 255 - 0xff
      11'h7BE: dout <= 8'b11111111; // 1982 : 255 - 0xff
      11'h7BF: dout <= 8'b11111111; // 1983 : 255 - 0xff
      11'h7C0: dout <= 8'b11111111; // 1984 : 255 - 0xff -- Background 0xf8
      11'h7C1: dout <= 8'b11111111; // 1985 : 255 - 0xff
      11'h7C2: dout <= 8'b11111101; // 1986 : 253 - 0xfd
      11'h7C3: dout <= 8'b11111000; // 1987 : 248 - 0xf8
      11'h7C4: dout <= 8'b11111111; // 1988 : 255 - 0xff
      11'h7C5: dout <= 8'b11111111; // 1989 : 255 - 0xff
      11'h7C6: dout <= 8'b11111110; // 1990 : 254 - 0xfe
      11'h7C7: dout <= 8'b11111111; // 1991 : 255 - 0xff
      11'h7C8: dout <= 8'b11111111; // 1992 : 255 - 0xff -- Background 0xf9
      11'h7C9: dout <= 8'b11111111; // 1993 : 255 - 0xff
      11'h7CA: dout <= 8'b11111111; // 1994 : 255 - 0xff
      11'h7CB: dout <= 8'b11111111; // 1995 : 255 - 0xff
      11'h7CC: dout <= 8'b11111111; // 1996 : 255 - 0xff
      11'h7CD: dout <= 8'b11111111; // 1997 : 255 - 0xff
      11'h7CE: dout <= 8'b11111111; // 1998 : 255 - 0xff
      11'h7CF: dout <= 8'b11111000; // 1999 : 248 - 0xf8
      11'h7D0: dout <= 8'b00000000; // 2000 :   0 - 0x0 -- Background 0xfa
      11'h7D1: dout <= 8'b00000000; // 2001 :   0 - 0x0
      11'h7D2: dout <= 8'b00000000; // 2002 :   0 - 0x0
      11'h7D3: dout <= 8'b00000000; // 2003 :   0 - 0x0
      11'h7D4: dout <= 8'b00000000; // 2004 :   0 - 0x0
      11'h7D5: dout <= 8'b00000000; // 2005 :   0 - 0x0
      11'h7D6: dout <= 8'b11000000; // 2006 : 192 - 0xc0
      11'h7D7: dout <= 8'b11110000; // 2007 : 240 - 0xf0
      11'h7D8: dout <= 8'b11111100; // 2008 : 252 - 0xfc -- Background 0xfb
      11'h7D9: dout <= 8'b11111110; // 2009 : 254 - 0xfe
      11'h7DA: dout <= 8'b11101100; // 2010 : 236 - 0xec
      11'h7DB: dout <= 8'b11100000; // 2011 : 224 - 0xe0
      11'h7DC: dout <= 8'b11000000; // 2012 : 192 - 0xc0
      11'h7DD: dout <= 8'b11000000; // 2013 : 192 - 0xc0
      11'h7DE: dout <= 8'b10000000; // 2014 : 128 - 0x80
      11'h7DF: dout <= 8'b10000000; // 2015 : 128 - 0x80
      11'h7E0: dout <= 8'b01110000; // 2016 : 112 - 0x70 -- Background 0xfc
      11'h7E1: dout <= 8'b11111100; // 2017 : 252 - 0xfc
      11'h7E2: dout <= 8'b11111100; // 2018 : 252 - 0xfc
      11'h7E3: dout <= 8'b11111100; // 2019 : 252 - 0xfc
      11'h7E4: dout <= 8'b11111100; // 2020 : 252 - 0xfc
      11'h7E5: dout <= 8'b11111100; // 2021 : 252 - 0xfc
      11'h7E6: dout <= 8'b11111110; // 2022 : 254 - 0xfe
      11'h7E7: dout <= 8'b11111110; // 2023 : 254 - 0xfe
      11'h7E8: dout <= 8'b11111110; // 2024 : 254 - 0xfe -- Background 0xfd
      11'h7E9: dout <= 8'b11111100; // 2025 : 252 - 0xfc
      11'h7EA: dout <= 8'b11111100; // 2026 : 252 - 0xfc
      11'h7EB: dout <= 8'b11111000; // 2027 : 248 - 0xf8
      11'h7EC: dout <= 8'b11110000; // 2028 : 240 - 0xf0
      11'h7ED: dout <= 8'b11100000; // 2029 : 224 - 0xe0
      11'h7EE: dout <= 8'b10000000; // 2030 : 128 - 0x80
      11'h7EF: dout <= 8'b00000000; // 2031 :   0 - 0x0
      11'h7F0: dout <= 8'b00000000; // 2032 :   0 - 0x0 -- Background 0xfe
      11'h7F1: dout <= 8'b00000000; // 2033 :   0 - 0x0
      11'h7F2: dout <= 8'b00000000; // 2034 :   0 - 0x0
      11'h7F3: dout <= 8'b00000000; // 2035 :   0 - 0x0
      11'h7F4: dout <= 8'b00000000; // 2036 :   0 - 0x0
      11'h7F5: dout <= 8'b00000000; // 2037 :   0 - 0x0
      11'h7F6: dout <= 8'b00000000; // 2038 :   0 - 0x0
      11'h7F7: dout <= 8'b00000000; // 2039 :   0 - 0x0
      11'h7F8: dout <= 8'b00000000; // 2040 :   0 - 0x0 -- Background 0xff
      11'h7F9: dout <= 8'b00000000; // 2041 :   0 - 0x0
      11'h7FA: dout <= 8'b00000000; // 2042 :   0 - 0x0
      11'h7FB: dout <= 8'b00000000; // 2043 :   0 - 0x0
      11'h7FC: dout <= 8'b00000000; // 2044 :   0 - 0x0
      11'h7FD: dout <= 8'b00000000; // 2045 :   0 - 0x0
      11'h7FE: dout <= 8'b00000000; // 2046 :   0 - 0x0
      11'h7FF: dout <= 8'b00000000; // 2047 :   0 - 0x0
    endcase
  end

endmodule
