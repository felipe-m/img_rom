--- Autcmatically generated VHDL ROM from a NES memory file----
---   SPRITEs MEMORY (OAM)
-- https://wiki.nesdev.com/w/index.php/PPU_OAM


---  Original memory dump file name: lawnmower_oam_00.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_OAM_LAWN_00 is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(8-1 downto 0);  --256 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_OAM_LAWN_00;

architecture BEHAVIORAL of ROM_OAM_LAWN_00 is
  signal addr_int  : natural range 0 to 2**8-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
    "00100000", --    0 -  0x0  :   32 - 0x20 -- Sprite 0x0
    "10101011", --    1 -  0x1  :  171 - 0xab
    "00000000", --    2 -  0x2  :    0 - 0x0
    "00000000", --    3 -  0x3  :    0 - 0x0
    "01111111", --    4 -  0x4  :  127 - 0x7f -- Sprite 0x1
    "11001001", --    5 -  0x5  :  201 - 0xc9
    "00000011", --    6 -  0x6  :    3 - 0x3
    "01101000", --    7 -  0x7  :  104 - 0x68
    "01111111", --    8 -  0x8  :  127 - 0x7f -- Sprite 0x2
    "11001010", --    9 -  0x9  :  202 - 0xca
    "00000011", --   10 -  0xa  :    3 - 0x3
    "01110000", --   11 -  0xb  :  112 - 0x70
    "01111111", --   12 -  0xc  :  127 - 0x7f -- Sprite 0x3
    "11001011", --   13 -  0xd  :  203 - 0xcb
    "00000011", --   14 -  0xe  :    3 - 0x3
    "01111000", --   15 -  0xf  :  120 - 0x78
    "10000111", --   16 - 0x10  :  135 - 0x87 -- Sprite 0x4
    "11001100", --   17 - 0x11  :  204 - 0xcc
    "00000011", --   18 - 0x12  :    3 - 0x3
    "01110000", --   19 - 0x13  :  112 - 0x70
    "10000111", --   20 - 0x14  :  135 - 0x87 -- Sprite 0x5
    "11001101", --   21 - 0x15  :  205 - 0xcd
    "00000011", --   22 - 0x16  :    3 - 0x3
    "01111000", --   23 - 0x17  :  120 - 0x78
    "01111111", --   24 - 0x18  :  127 - 0x7f -- Sprite 0x6
    "10110100", --   25 - 0x19  :  180 - 0xb4
    "00000010", --   26 - 0x1a  :    2 - 0x2
    "01110000", --   27 - 0x1b  :  112 - 0x70
    "01111111", --   28 - 0x1c  :  127 - 0x7f -- Sprite 0x7
    "10110101", --   29 - 0x1d  :  181 - 0xb5
    "00000010", --   30 - 0x1e  :    2 - 0x2
    "01111000", --   31 - 0x1f  :  120 - 0x78
    "10000111", --   32 - 0x20  :  135 - 0x87 -- Sprite 0x8
    "10110110", --   33 - 0x21  :  182 - 0xb6
    "00000010", --   34 - 0x22  :    2 - 0x2
    "01110000", --   35 - 0x23  :  112 - 0x70
    "10000111", --   36 - 0x24  :  135 - 0x87 -- Sprite 0x9
    "10110111", --   37 - 0x25  :  183 - 0xb7
    "00000010", --   38 - 0x26  :    2 - 0x2
    "01111000", --   39 - 0x27  :  120 - 0x78
    "01111111", --   40 - 0x28  :  127 - 0x7f -- Sprite 0xa
    "10101100", --   41 - 0x29  :  172 - 0xac
    "00000010", --   42 - 0x2a  :    2 - 0x2
    "01110000", --   43 - 0x2b  :  112 - 0x70
    "10000011", --   44 - 0x2c  :  131 - 0x83 -- Sprite 0xb
    "10101100", --   45 - 0x2d  :  172 - 0xac
    "00000001", --   46 - 0x2e  :    1 - 0x1
    "01101000", --   47 - 0x2f  :  104 - 0x68
    "11111111", --   48 - 0x30  :  255 - 0xff -- Sprite 0xc
    "11111111", --   49 - 0x31  :  255 - 0xff
    "11100011", --   50 - 0x32  :  227 - 0xe3
    "11111111", --   51 - 0x33  :  255 - 0xff
    "11111111", --   52 - 0x34  :  255 - 0xff -- Sprite 0xd
    "11111111", --   53 - 0x35  :  255 - 0xff
    "11100011", --   54 - 0x36  :  227 - 0xe3
    "11111111", --   55 - 0x37  :  255 - 0xff
    "11111111", --   56 - 0x38  :  255 - 0xff -- Sprite 0xe
    "11111111", --   57 - 0x39  :  255 - 0xff
    "11100011", --   58 - 0x3a  :  227 - 0xe3
    "11111111", --   59 - 0x3b  :  255 - 0xff
    "11111111", --   60 - 0x3c  :  255 - 0xff -- Sprite 0xf
    "11111111", --   61 - 0x3d  :  255 - 0xff
    "11100011", --   62 - 0x3e  :  227 - 0xe3
    "11111111", --   63 - 0x3f  :  255 - 0xff
    "11111111", --   64 - 0x40  :  255 - 0xff -- Sprite 0x10
    "11111111", --   65 - 0x41  :  255 - 0xff
    "11100011", --   66 - 0x42  :  227 - 0xe3
    "11111111", --   67 - 0x43  :  255 - 0xff
    "11111111", --   68 - 0x44  :  255 - 0xff -- Sprite 0x11
    "11111111", --   69 - 0x45  :  255 - 0xff
    "11100011", --   70 - 0x46  :  227 - 0xe3
    "11111111", --   71 - 0x47  :  255 - 0xff
    "11111111", --   72 - 0x48  :  255 - 0xff -- Sprite 0x12
    "11111111", --   73 - 0x49  :  255 - 0xff
    "11100011", --   74 - 0x4a  :  227 - 0xe3
    "11111111", --   75 - 0x4b  :  255 - 0xff
    "11111111", --   76 - 0x4c  :  255 - 0xff -- Sprite 0x13
    "11111111", --   77 - 0x4d  :  255 - 0xff
    "11100011", --   78 - 0x4e  :  227 - 0xe3
    "11111111", --   79 - 0x4f  :  255 - 0xff
    "11111111", --   80 - 0x50  :  255 - 0xff -- Sprite 0x14
    "11111111", --   81 - 0x51  :  255 - 0xff
    "11100011", --   82 - 0x52  :  227 - 0xe3
    "11111111", --   83 - 0x53  :  255 - 0xff
    "11111111", --   84 - 0x54  :  255 - 0xff -- Sprite 0x15
    "11111111", --   85 - 0x55  :  255 - 0xff
    "11100011", --   86 - 0x56  :  227 - 0xe3
    "11111111", --   87 - 0x57  :  255 - 0xff
    "11111111", --   88 - 0x58  :  255 - 0xff -- Sprite 0x16
    "11111111", --   89 - 0x59  :  255 - 0xff
    "11100011", --   90 - 0x5a  :  227 - 0xe3
    "11111111", --   91 - 0x5b  :  255 - 0xff
    "11111111", --   92 - 0x5c  :  255 - 0xff -- Sprite 0x17
    "11111111", --   93 - 0x5d  :  255 - 0xff
    "11100011", --   94 - 0x5e  :  227 - 0xe3
    "11111111", --   95 - 0x5f  :  255 - 0xff
    "11111111", --   96 - 0x60  :  255 - 0xff -- Sprite 0x18
    "11111111", --   97 - 0x61  :  255 - 0xff
    "11100011", --   98 - 0x62  :  227 - 0xe3
    "11111111", --   99 - 0x63  :  255 - 0xff
    "11111111", --  100 - 0x64  :  255 - 0xff -- Sprite 0x19
    "11111111", --  101 - 0x65  :  255 - 0xff
    "11100011", --  102 - 0x66  :  227 - 0xe3
    "11111111", --  103 - 0x67  :  255 - 0xff
    "11111111", --  104 - 0x68  :  255 - 0xff -- Sprite 0x1a
    "11111111", --  105 - 0x69  :  255 - 0xff
    "11100011", --  106 - 0x6a  :  227 - 0xe3
    "11111111", --  107 - 0x6b  :  255 - 0xff
    "11111111", --  108 - 0x6c  :  255 - 0xff -- Sprite 0x1b
    "11111111", --  109 - 0x6d  :  255 - 0xff
    "11100011", --  110 - 0x6e  :  227 - 0xe3
    "11111111", --  111 - 0x6f  :  255 - 0xff
    "11111111", --  112 - 0x70  :  255 - 0xff -- Sprite 0x1c
    "11111111", --  113 - 0x71  :  255 - 0xff
    "11100011", --  114 - 0x72  :  227 - 0xe3
    "11111111", --  115 - 0x73  :  255 - 0xff
    "11111111", --  116 - 0x74  :  255 - 0xff -- Sprite 0x1d
    "11111111", --  117 - 0x75  :  255 - 0xff
    "11100011", --  118 - 0x76  :  227 - 0xe3
    "11111111", --  119 - 0x77  :  255 - 0xff
    "11111111", --  120 - 0x78  :  255 - 0xff -- Sprite 0x1e
    "11111111", --  121 - 0x79  :  255 - 0xff
    "11100011", --  122 - 0x7a  :  227 - 0xe3
    "11111111", --  123 - 0x7b  :  255 - 0xff
    "11111111", --  124 - 0x7c  :  255 - 0xff -- Sprite 0x1f
    "11111111", --  125 - 0x7d  :  255 - 0xff
    "11100011", --  126 - 0x7e  :  227 - 0xe3
    "11111111", --  127 - 0x7f  :  255 - 0xff
    "11111111", --  128 - 0x80  :  255 - 0xff -- Sprite 0x20
    "11111111", --  129 - 0x81  :  255 - 0xff
    "11100011", --  130 - 0x82  :  227 - 0xe3
    "11111111", --  131 - 0x83  :  255 - 0xff
    "11111111", --  132 - 0x84  :  255 - 0xff -- Sprite 0x21
    "11111111", --  133 - 0x85  :  255 - 0xff
    "11100011", --  134 - 0x86  :  227 - 0xe3
    "11111111", --  135 - 0x87  :  255 - 0xff
    "11111111", --  136 - 0x88  :  255 - 0xff -- Sprite 0x22
    "11111111", --  137 - 0x89  :  255 - 0xff
    "11100011", --  138 - 0x8a  :  227 - 0xe3
    "11111111", --  139 - 0x8b  :  255 - 0xff
    "11111111", --  140 - 0x8c  :  255 - 0xff -- Sprite 0x23
    "11111111", --  141 - 0x8d  :  255 - 0xff
    "11100011", --  142 - 0x8e  :  227 - 0xe3
    "11111111", --  143 - 0x8f  :  255 - 0xff
    "11111111", --  144 - 0x90  :  255 - 0xff -- Sprite 0x24
    "11111111", --  145 - 0x91  :  255 - 0xff
    "11100011", --  146 - 0x92  :  227 - 0xe3
    "11111111", --  147 - 0x93  :  255 - 0xff
    "11111111", --  148 - 0x94  :  255 - 0xff -- Sprite 0x25
    "11111111", --  149 - 0x95  :  255 - 0xff
    "11100011", --  150 - 0x96  :  227 - 0xe3
    "11111111", --  151 - 0x97  :  255 - 0xff
    "11111111", --  152 - 0x98  :  255 - 0xff -- Sprite 0x26
    "11111111", --  153 - 0x99  :  255 - 0xff
    "11100011", --  154 - 0x9a  :  227 - 0xe3
    "11111111", --  155 - 0x9b  :  255 - 0xff
    "11111111", --  156 - 0x9c  :  255 - 0xff -- Sprite 0x27
    "11111111", --  157 - 0x9d  :  255 - 0xff
    "11100011", --  158 - 0x9e  :  227 - 0xe3
    "11111111", --  159 - 0x9f  :  255 - 0xff
    "11111111", --  160 - 0xa0  :  255 - 0xff -- Sprite 0x28
    "11111111", --  161 - 0xa1  :  255 - 0xff
    "11100011", --  162 - 0xa2  :  227 - 0xe3
    "11111111", --  163 - 0xa3  :  255 - 0xff
    "11111111", --  164 - 0xa4  :  255 - 0xff -- Sprite 0x29
    "11111111", --  165 - 0xa5  :  255 - 0xff
    "11100011", --  166 - 0xa6  :  227 - 0xe3
    "11111111", --  167 - 0xa7  :  255 - 0xff
    "11111111", --  168 - 0xa8  :  255 - 0xff -- Sprite 0x2a
    "11111111", --  169 - 0xa9  :  255 - 0xff
    "11100011", --  170 - 0xaa  :  227 - 0xe3
    "11111111", --  171 - 0xab  :  255 - 0xff
    "11111111", --  172 - 0xac  :  255 - 0xff -- Sprite 0x2b
    "11111111", --  173 - 0xad  :  255 - 0xff
    "11100011", --  174 - 0xae  :  227 - 0xe3
    "11111111", --  175 - 0xaf  :  255 - 0xff
    "11111111", --  176 - 0xb0  :  255 - 0xff -- Sprite 0x2c
    "11111111", --  177 - 0xb1  :  255 - 0xff
    "11100011", --  178 - 0xb2  :  227 - 0xe3
    "11111111", --  179 - 0xb3  :  255 - 0xff
    "11111111", --  180 - 0xb4  :  255 - 0xff -- Sprite 0x2d
    "11111111", --  181 - 0xb5  :  255 - 0xff
    "11100011", --  182 - 0xb6  :  227 - 0xe3
    "11111111", --  183 - 0xb7  :  255 - 0xff
    "11111111", --  184 - 0xb8  :  255 - 0xff -- Sprite 0x2e
    "11111111", --  185 - 0xb9  :  255 - 0xff
    "11100011", --  186 - 0xba  :  227 - 0xe3
    "11111111", --  187 - 0xbb  :  255 - 0xff
    "11111111", --  188 - 0xbc  :  255 - 0xff -- Sprite 0x2f
    "11111111", --  189 - 0xbd  :  255 - 0xff
    "11100011", --  190 - 0xbe  :  227 - 0xe3
    "11111111", --  191 - 0xbf  :  255 - 0xff
    "11111111", --  192 - 0xc0  :  255 - 0xff -- Sprite 0x30
    "11111111", --  193 - 0xc1  :  255 - 0xff
    "11100011", --  194 - 0xc2  :  227 - 0xe3
    "11111111", --  195 - 0xc3  :  255 - 0xff
    "11111111", --  196 - 0xc4  :  255 - 0xff -- Sprite 0x31
    "11111111", --  197 - 0xc5  :  255 - 0xff
    "11100011", --  198 - 0xc6  :  227 - 0xe3
    "11111111", --  199 - 0xc7  :  255 - 0xff
    "11111111", --  200 - 0xc8  :  255 - 0xff -- Sprite 0x32
    "11111111", --  201 - 0xc9  :  255 - 0xff
    "11100011", --  202 - 0xca  :  227 - 0xe3
    "11111111", --  203 - 0xcb  :  255 - 0xff
    "11111111", --  204 - 0xcc  :  255 - 0xff -- Sprite 0x33
    "11111111", --  205 - 0xcd  :  255 - 0xff
    "11100011", --  206 - 0xce  :  227 - 0xe3
    "11111111", --  207 - 0xcf  :  255 - 0xff
    "11111111", --  208 - 0xd0  :  255 - 0xff -- Sprite 0x34
    "11111111", --  209 - 0xd1  :  255 - 0xff
    "11100011", --  210 - 0xd2  :  227 - 0xe3
    "11111111", --  211 - 0xd3  :  255 - 0xff
    "11111111", --  212 - 0xd4  :  255 - 0xff -- Sprite 0x35
    "11111111", --  213 - 0xd5  :  255 - 0xff
    "11100011", --  214 - 0xd6  :  227 - 0xe3
    "11111111", --  215 - 0xd7  :  255 - 0xff
    "11111111", --  216 - 0xd8  :  255 - 0xff -- Sprite 0x36
    "11111111", --  217 - 0xd9  :  255 - 0xff
    "11100011", --  218 - 0xda  :  227 - 0xe3
    "11111111", --  219 - 0xdb  :  255 - 0xff
    "11111111", --  220 - 0xdc  :  255 - 0xff -- Sprite 0x37
    "11111111", --  221 - 0xdd  :  255 - 0xff
    "11100011", --  222 - 0xde  :  227 - 0xe3
    "11111111", --  223 - 0xdf  :  255 - 0xff
    "00010101", --  224 - 0xe0  :   21 - 0x15 -- Sprite 0x38
    "11111000", --  225 - 0xe1  :  248 - 0xf8
    "00000000", --  226 - 0xe2  :    0 - 0x0
    "01101011", --  227 - 0xe3  :  107 - 0x6b
    "00010101", --  228 - 0xe4  :   21 - 0x15 -- Sprite 0x39
    "11111000", --  229 - 0xe5  :  248 - 0xf8
    "00000000", --  230 - 0xe6  :    0 - 0x0
    "01110011", --  231 - 0xe7  :  115 - 0x73
    "00010101", --  232 - 0xe8  :   21 - 0x15 -- Sprite 0x3a
    "11111000", --  233 - 0xe9  :  248 - 0xf8
    "00000000", --  234 - 0xea  :    0 - 0x0
    "01111011", --  235 - 0xeb  :  123 - 0x7b
    "00010101", --  236 - 0xec  :   21 - 0x15 -- Sprite 0x3b
    "11110100", --  237 - 0xed  :  244 - 0xf4
    "00000000", --  238 - 0xee  :    0 - 0x0
    "10000011", --  239 - 0xef  :  131 - 0x83
    "11101111", --  240 - 0xf0  :  239 - 0xef -- Sprite 0x3c
    "11111000", --  241 - 0xf1  :  248 - 0xf8
    "00000000", --  242 - 0xf2  :    0 - 0x0
    "10001011", --  243 - 0xf3  :  139 - 0x8b
    "11101111", --  244 - 0xf4  :  239 - 0xef -- Sprite 0x3d
    "11111000", --  245 - 0xf5  :  248 - 0xf8
    "00000000", --  246 - 0xf6  :    0 - 0x0
    "10010011", --  247 - 0xf7  :  147 - 0x93
    "11101111", --  248 - 0xf8  :  239 - 0xef -- Sprite 0x3e
    "11111000", --  249 - 0xf9  :  248 - 0xf8
    "00000000", --  250 - 0xfa  :    0 - 0x0
    "10011011", --  251 - 0xfb  :  155 - 0x9b
    "11101111", --  252 - 0xfc  :  239 - 0xef -- Sprite 0x3f
    "11111000", --  253 - 0xfd  :  248 - 0xf8
    "00000000", --  254 - 0xfe  :    0 - 0x0
    "10100011"  --  255 - 0xff  :  163 - 0xa3
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
