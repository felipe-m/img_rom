//- Autcmatically generated verilog ROM from a NES memory file----
//-   PATTERN TABLE
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


//-  Original memory dump file name: lawnmower_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_PTABLE_LAWN
  (
     input     clk,   // clock
     input      [13-1:0] addr,  //8192 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Pattern Table 0---------
      13'h0: dout <= 8'b11111111; //    0 : 255 - 0xff -- Sprite 0x0
      13'h1: dout <= 8'b11111111; //    1 : 255 - 0xff
      13'h2: dout <= 8'b11111111; //    2 : 255 - 0xff
      13'h3: dout <= 8'b11111111; //    3 : 255 - 0xff
      13'h4: dout <= 8'b11111111; //    4 : 255 - 0xff
      13'h5: dout <= 8'b11111111; //    5 : 255 - 0xff
      13'h6: dout <= 8'b11111111; //    6 : 255 - 0xff
      13'h7: dout <= 8'b11111111; //    7 : 255 - 0xff
      13'h8: dout <= 8'b00000000; //    8 :   0 - 0x0
      13'h9: dout <= 8'b00000000; //    9 :   0 - 0x0
      13'hA: dout <= 8'b00000000; //   10 :   0 - 0x0
      13'hB: dout <= 8'b00000000; //   11 :   0 - 0x0
      13'hC: dout <= 8'b00000000; //   12 :   0 - 0x0
      13'hD: dout <= 8'b00000000; //   13 :   0 - 0x0
      13'hE: dout <= 8'b00000000; //   14 :   0 - 0x0
      13'hF: dout <= 8'b00000000; //   15 :   0 - 0x0
      13'h10: dout <= 8'b11111111; //   16 : 255 - 0xff -- Sprite 0x1
      13'h11: dout <= 8'b11111111; //   17 : 255 - 0xff
      13'h12: dout <= 8'b11111111; //   18 : 255 - 0xff
      13'h13: dout <= 8'b11111111; //   19 : 255 - 0xff
      13'h14: dout <= 8'b11111111; //   20 : 255 - 0xff
      13'h15: dout <= 8'b11111111; //   21 : 255 - 0xff
      13'h16: dout <= 8'b11111100; //   22 : 252 - 0xfc
      13'h17: dout <= 8'b11111100; //   23 : 252 - 0xfc
      13'h18: dout <= 8'b00000000; //   24 :   0 - 0x0
      13'h19: dout <= 8'b00000000; //   25 :   0 - 0x0
      13'h1A: dout <= 8'b00000000; //   26 :   0 - 0x0
      13'h1B: dout <= 8'b00000000; //   27 :   0 - 0x0
      13'h1C: dout <= 8'b00000000; //   28 :   0 - 0x0
      13'h1D: dout <= 8'b00000111; //   29 :   7 - 0x7
      13'h1E: dout <= 8'b00000111; //   30 :   7 - 0x7
      13'h1F: dout <= 8'b00000110; //   31 :   6 - 0x6
      13'h20: dout <= 8'b11111111; //   32 : 255 - 0xff -- Sprite 0x2
      13'h21: dout <= 8'b11111111; //   33 : 255 - 0xff
      13'h22: dout <= 8'b11111111; //   34 : 255 - 0xff
      13'h23: dout <= 8'b11111111; //   35 : 255 - 0xff
      13'h24: dout <= 8'b11111111; //   36 : 255 - 0xff
      13'h25: dout <= 8'b11111111; //   37 : 255 - 0xff
      13'h26: dout <= 8'b00000000; //   38 :   0 - 0x0
      13'h27: dout <= 8'b00000000; //   39 :   0 - 0x0
      13'h28: dout <= 8'b00000000; //   40 :   0 - 0x0
      13'h29: dout <= 8'b00000000; //   41 :   0 - 0x0
      13'h2A: dout <= 8'b00000000; //   42 :   0 - 0x0
      13'h2B: dout <= 8'b00000000; //   43 :   0 - 0x0
      13'h2C: dout <= 8'b00000000; //   44 :   0 - 0x0
      13'h2D: dout <= 8'b11111111; //   45 : 255 - 0xff
      13'h2E: dout <= 8'b11111111; //   46 : 255 - 0xff
      13'h2F: dout <= 8'b00000000; //   47 :   0 - 0x0
      13'h30: dout <= 8'b11111111; //   48 : 255 - 0xff -- Sprite 0x3
      13'h31: dout <= 8'b11111111; //   49 : 255 - 0xff
      13'h32: dout <= 8'b11111111; //   50 : 255 - 0xff
      13'h33: dout <= 8'b11111111; //   51 : 255 - 0xff
      13'h34: dout <= 8'b11111111; //   52 : 255 - 0xff
      13'h35: dout <= 8'b11111111; //   53 : 255 - 0xff
      13'h36: dout <= 8'b00011111; //   54 :  31 - 0x1f
      13'h37: dout <= 8'b01000111; //   55 :  71 - 0x47
      13'h38: dout <= 8'b00000000; //   56 :   0 - 0x0
      13'h39: dout <= 8'b00000000; //   57 :   0 - 0x0
      13'h3A: dout <= 8'b00000000; //   58 :   0 - 0x0
      13'h3B: dout <= 8'b00000000; //   59 :   0 - 0x0
      13'h3C: dout <= 8'b00000000; //   60 :   0 - 0x0
      13'h3D: dout <= 8'b11100000; //   61 : 224 - 0xe0
      13'h3E: dout <= 8'b11100000; //   62 : 224 - 0xe0
      13'h3F: dout <= 8'b01100000; //   63 :  96 - 0x60
      13'h40: dout <= 8'b11111111; //   64 : 255 - 0xff -- Sprite 0x4
      13'h41: dout <= 8'b11111111; //   65 : 255 - 0xff
      13'h42: dout <= 8'b11111111; //   66 : 255 - 0xff
      13'h43: dout <= 8'b11111111; //   67 : 255 - 0xff
      13'h44: dout <= 8'b11111111; //   68 : 255 - 0xff
      13'h45: dout <= 8'b11111111; //   69 : 255 - 0xff
      13'h46: dout <= 8'b11100000; //   70 : 224 - 0xe0
      13'h47: dout <= 8'b10000000; //   71 : 128 - 0x80
      13'h48: dout <= 8'b00000000; //   72 :   0 - 0x0
      13'h49: dout <= 8'b00000000; //   73 :   0 - 0x0
      13'h4A: dout <= 8'b00000000; //   74 :   0 - 0x0
      13'h4B: dout <= 8'b00000000; //   75 :   0 - 0x0
      13'h4C: dout <= 8'b00000000; //   76 :   0 - 0x0
      13'h4D: dout <= 8'b00011111; //   77 :  31 - 0x1f
      13'h4E: dout <= 8'b01111111; //   78 : 127 - 0x7f
      13'h4F: dout <= 8'b11110000; //   79 : 240 - 0xf0
      13'h50: dout <= 8'b11111111; //   80 : 255 - 0xff -- Sprite 0x5
      13'h51: dout <= 8'b11111111; //   81 : 255 - 0xff
      13'h52: dout <= 8'b11111111; //   82 : 255 - 0xff
      13'h53: dout <= 8'b11111111; //   83 : 255 - 0xff
      13'h54: dout <= 8'b11111111; //   84 : 255 - 0xff
      13'h55: dout <= 8'b11110111; //   85 : 247 - 0xf7
      13'h56: dout <= 8'b00000001; //   86 :   1 - 0x1
      13'h57: dout <= 8'b00000100; //   87 :   4 - 0x4
      13'h58: dout <= 8'b00000000; //   88 :   0 - 0x0
      13'h59: dout <= 8'b00000000; //   89 :   0 - 0x0
      13'h5A: dout <= 8'b00000000; //   90 :   0 - 0x0
      13'h5B: dout <= 8'b00000000; //   91 :   0 - 0x0
      13'h5C: dout <= 8'b00000000; //   92 :   0 - 0x0
      13'h5D: dout <= 8'b11111000; //   93 : 248 - 0xf8
      13'h5E: dout <= 8'b11111110; //   94 : 254 - 0xfe
      13'h5F: dout <= 8'b00001111; //   95 :  15 - 0xf
      13'h60: dout <= 8'b11111111; //   96 : 255 - 0xff -- Sprite 0x6
      13'h61: dout <= 8'b11111111; //   97 : 255 - 0xff
      13'h62: dout <= 8'b11111111; //   98 : 255 - 0xff
      13'h63: dout <= 8'b11111111; //   99 : 255 - 0xff
      13'h64: dout <= 8'b11111111; //  100 : 255 - 0xff
      13'h65: dout <= 8'b11011111; //  101 : 223 - 0xdf
      13'h66: dout <= 8'b00011100; //  102 :  28 - 0x1c
      13'h67: dout <= 8'b01000100; //  103 :  68 - 0x44
      13'h68: dout <= 8'b00000000; //  104 :   0 - 0x0
      13'h69: dout <= 8'b00000000; //  105 :   0 - 0x0
      13'h6A: dout <= 8'b00000000; //  106 :   0 - 0x0
      13'h6B: dout <= 8'b00000000; //  107 :   0 - 0x0
      13'h6C: dout <= 8'b00000000; //  108 :   0 - 0x0
      13'h6D: dout <= 8'b11100111; //  109 : 231 - 0xe7
      13'h6E: dout <= 8'b11100111; //  110 : 231 - 0xe7
      13'h6F: dout <= 8'b01100110; //  111 : 102 - 0x66
      13'h70: dout <= 8'b11111111; //  112 : 255 - 0xff -- Sprite 0x7
      13'h71: dout <= 8'b11111111; //  113 : 255 - 0xff
      13'h72: dout <= 8'b11111111; //  114 : 255 - 0xff
      13'h73: dout <= 8'b11111111; //  115 : 255 - 0xff
      13'h74: dout <= 8'b11111111; //  116 : 255 - 0xff
      13'h75: dout <= 8'b10111111; //  117 : 191 - 0xbf
      13'h76: dout <= 8'b00111100; //  118 :  60 - 0x3c
      13'h77: dout <= 8'b01001100; //  119 :  76 - 0x4c
      13'h78: dout <= 8'b00000000; //  120 :   0 - 0x0
      13'h79: dout <= 8'b00000000; //  121 :   0 - 0x0
      13'h7A: dout <= 8'b00000000; //  122 :   0 - 0x0
      13'h7B: dout <= 8'b00000000; //  123 :   0 - 0x0
      13'h7C: dout <= 8'b00000000; //  124 :   0 - 0x0
      13'h7D: dout <= 8'b11000111; //  125 : 199 - 0xc7
      13'h7E: dout <= 8'b11000111; //  126 : 199 - 0xc7
      13'h7F: dout <= 8'b01100110; //  127 : 102 - 0x66
      13'h80: dout <= 8'b11111100; //  128 : 252 - 0xfc -- Sprite 0x8
      13'h81: dout <= 8'b11111100; //  129 : 252 - 0xfc
      13'h82: dout <= 8'b11111100; //  130 : 252 - 0xfc
      13'h83: dout <= 8'b11111100; //  131 : 252 - 0xfc
      13'h84: dout <= 8'b11111100; //  132 : 252 - 0xfc
      13'h85: dout <= 8'b11111100; //  133 : 252 - 0xfc
      13'h86: dout <= 8'b11111100; //  134 : 252 - 0xfc
      13'h87: dout <= 8'b11111100; //  135 : 252 - 0xfc
      13'h88: dout <= 8'b00000110; //  136 :   6 - 0x6
      13'h89: dout <= 8'b00000110; //  137 :   6 - 0x6
      13'h8A: dout <= 8'b00000110; //  138 :   6 - 0x6
      13'h8B: dout <= 8'b00000110; //  139 :   6 - 0x6
      13'h8C: dout <= 8'b00000110; //  140 :   6 - 0x6
      13'h8D: dout <= 8'b00000110; //  141 :   6 - 0x6
      13'h8E: dout <= 8'b00000110; //  142 :   6 - 0x6
      13'h8F: dout <= 8'b00000110; //  143 :   6 - 0x6
      13'h90: dout <= 8'b00010000; //  144 :  16 - 0x10 -- Sprite 0x9
      13'h91: dout <= 8'b00111000; //  145 :  56 - 0x38
      13'h92: dout <= 8'b01111100; //  146 : 124 - 0x7c
      13'h93: dout <= 8'b11111000; //  147 : 248 - 0xf8
      13'h94: dout <= 8'b01110000; //  148 : 112 - 0x70
      13'h95: dout <= 8'b00100010; //  149 :  34 - 0x22
      13'h96: dout <= 8'b00000101; //  150 :   5 - 0x5
      13'h97: dout <= 8'b00000010; //  151 :   2 - 0x2
      13'h98: dout <= 8'b11111111; //  152 : 255 - 0xff
      13'h99: dout <= 8'b11111111; //  153 : 255 - 0xff
      13'h9A: dout <= 8'b11111111; //  154 : 255 - 0xff
      13'h9B: dout <= 8'b11111111; //  155 : 255 - 0xff
      13'h9C: dout <= 8'b11111111; //  156 : 255 - 0xff
      13'h9D: dout <= 8'b11111111; //  157 : 255 - 0xff
      13'h9E: dout <= 8'b11111111; //  158 : 255 - 0xff
      13'h9F: dout <= 8'b11111111; //  159 : 255 - 0xff
      13'hA0: dout <= 8'b01000111; //  160 :  71 - 0x47 -- Sprite 0xa
      13'hA1: dout <= 8'b01000111; //  161 :  71 - 0x47
      13'hA2: dout <= 8'b01000111; //  162 :  71 - 0x47
      13'hA3: dout <= 8'b01000111; //  163 :  71 - 0x47
      13'hA4: dout <= 8'b01000111; //  164 :  71 - 0x47
      13'hA5: dout <= 8'b01000111; //  165 :  71 - 0x47
      13'hA6: dout <= 8'b01000111; //  166 :  71 - 0x47
      13'hA7: dout <= 8'b01000111; //  167 :  71 - 0x47
      13'hA8: dout <= 8'b01100000; //  168 :  96 - 0x60
      13'hA9: dout <= 8'b01100000; //  169 :  96 - 0x60
      13'hAA: dout <= 8'b01100000; //  170 :  96 - 0x60
      13'hAB: dout <= 8'b01100000; //  171 :  96 - 0x60
      13'hAC: dout <= 8'b01100000; //  172 :  96 - 0x60
      13'hAD: dout <= 8'b01100000; //  173 :  96 - 0x60
      13'hAE: dout <= 8'b01100000; //  174 :  96 - 0x60
      13'hAF: dout <= 8'b01100000; //  175 :  96 - 0x60
      13'hB0: dout <= 8'b11111111; //  176 : 255 - 0xff -- Sprite 0xb
      13'hB1: dout <= 8'b11111110; //  177 : 254 - 0xfe
      13'hB2: dout <= 8'b11111110; //  178 : 254 - 0xfe
      13'hB3: dout <= 8'b11111100; //  179 : 252 - 0xfc
      13'hB4: dout <= 8'b11111100; //  180 : 252 - 0xfc
      13'hB5: dout <= 8'b11111100; //  181 : 252 - 0xfc
      13'hB6: dout <= 8'b11111100; //  182 : 252 - 0xfc
      13'hB7: dout <= 8'b11111100; //  183 : 252 - 0xfc
      13'hB8: dout <= 8'b00000001; //  184 :   1 - 0x1
      13'hB9: dout <= 8'b00000011; //  185 :   3 - 0x3
      13'hBA: dout <= 8'b00000011; //  186 :   3 - 0x3
      13'hBB: dout <= 8'b00000111; //  187 :   7 - 0x7
      13'hBC: dout <= 8'b00000110; //  188 :   6 - 0x6
      13'hBD: dout <= 8'b00000110; //  189 :   6 - 0x6
      13'hBE: dout <= 8'b00000110; //  190 :   6 - 0x6
      13'hBF: dout <= 8'b00000110; //  191 :   6 - 0x6
      13'hC0: dout <= 8'b00000000; //  192 :   0 - 0x0 -- Sprite 0xc
      13'hC1: dout <= 8'b00001000; //  193 :   8 - 0x8
      13'hC2: dout <= 8'b00011100; //  194 :  28 - 0x1c
      13'hC3: dout <= 8'b00111000; //  195 :  56 - 0x38
      13'hC4: dout <= 8'b01110000; //  196 : 112 - 0x70
      13'hC5: dout <= 8'b00100010; //  197 :  34 - 0x22
      13'hC6: dout <= 8'b00000101; //  198 :   5 - 0x5
      13'hC7: dout <= 8'b00000010; //  199 :   2 - 0x2
      13'hC8: dout <= 8'b11000111; //  200 : 199 - 0xc7
      13'hC9: dout <= 8'b10011111; //  201 : 159 - 0x9f
      13'hCA: dout <= 8'b00111111; //  202 :  63 - 0x3f
      13'hCB: dout <= 8'b01111111; //  203 : 127 - 0x7f
      13'hCC: dout <= 8'b01111111; //  204 : 127 - 0x7f
      13'hCD: dout <= 8'b11111111; //  205 : 255 - 0xff
      13'hCE: dout <= 8'b11111111; //  206 : 255 - 0xff
      13'hCF: dout <= 8'b11111111; //  207 : 255 - 0xff
      13'hD0: dout <= 8'b00000010; //  208 :   2 - 0x2 -- Sprite 0xd
      13'hD1: dout <= 8'b00110001; //  209 :  49 - 0x31
      13'hD2: dout <= 8'b01111000; //  210 : 120 - 0x78
      13'hD3: dout <= 8'b11111000; //  211 : 248 - 0xf8
      13'hD4: dout <= 8'b01110000; //  212 : 112 - 0x70
      13'hD5: dout <= 8'b00100010; //  213 :  34 - 0x22
      13'hD6: dout <= 8'b00000101; //  214 :   5 - 0x5
      13'hD7: dout <= 8'b00000010; //  215 :   2 - 0x2
      13'hD8: dout <= 8'b11100011; //  216 : 227 - 0xe3
      13'hD9: dout <= 8'b11111001; //  217 : 249 - 0xf9
      13'hDA: dout <= 8'b11111100; //  218 : 252 - 0xfc
      13'hDB: dout <= 8'b11111110; //  219 : 254 - 0xfe
      13'hDC: dout <= 8'b11111110; //  220 : 254 - 0xfe
      13'hDD: dout <= 8'b11111111; //  221 : 255 - 0xff
      13'hDE: dout <= 8'b11111111; //  222 : 255 - 0xff
      13'hDF: dout <= 8'b11111111; //  223 : 255 - 0xff
      13'hE0: dout <= 8'b01111100; //  224 : 124 - 0x7c -- Sprite 0xe
      13'hE1: dout <= 8'b00111100; //  225 :  60 - 0x3c
      13'hE2: dout <= 8'b10011100; //  226 : 156 - 0x9c
      13'hE3: dout <= 8'b10001100; //  227 : 140 - 0x8c
      13'hE4: dout <= 8'b01001100; //  228 :  76 - 0x4c
      13'hE5: dout <= 8'b01000100; //  229 :  68 - 0x44
      13'hE6: dout <= 8'b01000100; //  230 :  68 - 0x44
      13'hE7: dout <= 8'b01000100; //  231 :  68 - 0x44
      13'hE8: dout <= 8'b10000110; //  232 : 134 - 0x86
      13'hE9: dout <= 8'b11000110; //  233 : 198 - 0xc6
      13'hEA: dout <= 8'b11000110; //  234 : 198 - 0xc6
      13'hEB: dout <= 8'b11100110; //  235 : 230 - 0xe6
      13'hEC: dout <= 8'b01100110; //  236 : 102 - 0x66
      13'hED: dout <= 8'b01100110; //  237 : 102 - 0x66
      13'hEE: dout <= 8'b01100110; //  238 : 102 - 0x66
      13'hEF: dout <= 8'b01100110; //  239 : 102 - 0x66
      13'hF0: dout <= 8'b01000100; //  240 :  68 - 0x44 -- Sprite 0xf
      13'hF1: dout <= 8'b01000100; //  241 :  68 - 0x44
      13'hF2: dout <= 8'b01000100; //  242 :  68 - 0x44
      13'hF3: dout <= 8'b01000100; //  243 :  68 - 0x44
      13'hF4: dout <= 8'b01000100; //  244 :  68 - 0x44
      13'hF5: dout <= 8'b01000100; //  245 :  68 - 0x44
      13'hF6: dout <= 8'b01000100; //  246 :  68 - 0x44
      13'hF7: dout <= 8'b01000100; //  247 :  68 - 0x44
      13'hF8: dout <= 8'b01100110; //  248 : 102 - 0x66
      13'hF9: dout <= 8'b01100110; //  249 : 102 - 0x66
      13'hFA: dout <= 8'b01100110; //  250 : 102 - 0x66
      13'hFB: dout <= 8'b01100110; //  251 : 102 - 0x66
      13'hFC: dout <= 8'b01100110; //  252 : 102 - 0x66
      13'hFD: dout <= 8'b01100110; //  253 : 102 - 0x66
      13'hFE: dout <= 8'b01100110; //  254 : 102 - 0x66
      13'hFF: dout <= 8'b01100110; //  255 : 102 - 0x66
      13'h100: dout <= 8'b01001100; //  256 :  76 - 0x4c -- Sprite 0x10
      13'h101: dout <= 8'b00100100; //  257 :  36 - 0x24
      13'h102: dout <= 8'b00100100; //  258 :  36 - 0x24
      13'h103: dout <= 8'b10010100; //  259 : 148 - 0x94
      13'h104: dout <= 8'b00010000; //  260 :  16 - 0x10
      13'h105: dout <= 8'b00001000; //  261 :   8 - 0x8
      13'h106: dout <= 8'b00001000; //  262 :   8 - 0x8
      13'h107: dout <= 8'b00000100; //  263 :   4 - 0x4
      13'h108: dout <= 8'b01100110; //  264 : 102 - 0x66
      13'h109: dout <= 8'b00110110; //  265 :  54 - 0x36
      13'h10A: dout <= 8'b10110110; //  266 : 182 - 0xb6
      13'h10B: dout <= 8'b10011110; //  267 : 158 - 0x9e
      13'h10C: dout <= 8'b11011110; //  268 : 222 - 0xde
      13'h10D: dout <= 8'b11001110; //  269 : 206 - 0xce
      13'h10E: dout <= 8'b11101110; //  270 : 238 - 0xee
      13'h10F: dout <= 8'b11100110; //  271 : 230 - 0xe6
      13'h110: dout <= 8'b00000000; //  272 :   0 - 0x0 -- Sprite 0x11
      13'h111: dout <= 8'b00111100; //  273 :  60 - 0x3c
      13'h112: dout <= 8'b01000000; //  274 :  64 - 0x40
      13'h113: dout <= 8'b01000100; //  275 :  68 - 0x44
      13'h114: dout <= 8'b01000100; //  276 :  68 - 0x44
      13'h115: dout <= 8'b01000100; //  277 :  68 - 0x44
      13'h116: dout <= 8'b01000100; //  278 :  68 - 0x44
      13'h117: dout <= 8'b01000100; //  279 :  68 - 0x44
      13'h118: dout <= 8'b10000001; //  280 : 129 - 0x81
      13'h119: dout <= 8'b00111100; //  281 :  60 - 0x3c
      13'h11A: dout <= 8'b01111110; //  282 : 126 - 0x7e
      13'h11B: dout <= 8'b01100110; //  283 : 102 - 0x66
      13'h11C: dout <= 8'b01100110; //  284 : 102 - 0x66
      13'h11D: dout <= 8'b01100110; //  285 : 102 - 0x66
      13'h11E: dout <= 8'b01100110; //  286 : 102 - 0x66
      13'h11F: dout <= 8'b01100110; //  287 : 102 - 0x66
      13'h120: dout <= 8'b00000100; //  288 :   4 - 0x4 -- Sprite 0x12
      13'h121: dout <= 8'b00010010; //  289 :  18 - 0x12
      13'h122: dout <= 8'b00110010; //  290 :  50 - 0x32
      13'h123: dout <= 8'b01111000; //  291 : 120 - 0x78
      13'h124: dout <= 8'b11111000; //  292 : 248 - 0xf8
      13'h125: dout <= 8'b01110000; //  293 : 112 - 0x70
      13'h126: dout <= 8'b00100100; //  294 :  36 - 0x24
      13'h127: dout <= 8'b00000000; //  295 :   0 - 0x0
      13'h128: dout <= 8'b11110110; //  296 : 246 - 0xf6
      13'h129: dout <= 8'b11110010; //  297 : 242 - 0xf2
      13'h12A: dout <= 8'b11111010; //  298 : 250 - 0xfa
      13'h12B: dout <= 8'b11111000; //  299 : 248 - 0xf8
      13'h12C: dout <= 8'b11111100; //  300 : 252 - 0xfc
      13'h12D: dout <= 8'b11111100; //  301 : 252 - 0xfc
      13'h12E: dout <= 8'b11111110; //  302 : 254 - 0xfe
      13'h12F: dout <= 8'b11111110; //  303 : 254 - 0xfe
      13'h130: dout <= 8'b01000100; //  304 :  68 - 0x44 -- Sprite 0x13
      13'h131: dout <= 8'b01000100; //  305 :  68 - 0x44
      13'h132: dout <= 8'b01000100; //  306 :  68 - 0x44
      13'h133: dout <= 8'b01000100; //  307 :  68 - 0x44
      13'h134: dout <= 8'b01000100; //  308 :  68 - 0x44
      13'h135: dout <= 8'b01000100; //  309 :  68 - 0x44
      13'h136: dout <= 8'b01000100; //  310 :  68 - 0x44
      13'h137: dout <= 8'b01011100; //  311 :  92 - 0x5c
      13'h138: dout <= 8'b01100110; //  312 : 102 - 0x66
      13'h139: dout <= 8'b01100110; //  313 : 102 - 0x66
      13'h13A: dout <= 8'b01100110; //  314 : 102 - 0x66
      13'h13B: dout <= 8'b01100110; //  315 : 102 - 0x66
      13'h13C: dout <= 8'b01100110; //  316 : 102 - 0x66
      13'h13D: dout <= 8'b01100110; //  317 : 102 - 0x66
      13'h13E: dout <= 8'b01100110; //  318 : 102 - 0x66
      13'h13F: dout <= 8'b01111110; //  319 : 126 - 0x7e
      13'h140: dout <= 8'b00010000; //  320 :  16 - 0x10 -- Sprite 0x14
      13'h141: dout <= 8'b00111000; //  321 :  56 - 0x38
      13'h142: dout <= 8'b00111100; //  322 :  60 - 0x3c
      13'h143: dout <= 8'b00111000; //  323 :  56 - 0x38
      13'h144: dout <= 8'b00010000; //  324 :  16 - 0x10
      13'h145: dout <= 8'b00000010; //  325 :   2 - 0x2
      13'h146: dout <= 8'b01000101; //  326 :  69 - 0x45
      13'h147: dout <= 8'b01000010; //  327 :  66 - 0x42
      13'h148: dout <= 8'b11111111; //  328 : 255 - 0xff
      13'h149: dout <= 8'b01111111; //  329 : 127 - 0x7f
      13'h14A: dout <= 8'b01111111; //  330 : 127 - 0x7f
      13'h14B: dout <= 8'b00111111; //  331 :  63 - 0x3f
      13'h14C: dout <= 8'b00111111; //  332 :  63 - 0x3f
      13'h14D: dout <= 8'b00011111; //  333 :  31 - 0x1f
      13'h14E: dout <= 8'b01011111; //  334 :  95 - 0x5f
      13'h14F: dout <= 8'b01001111; //  335 :  79 - 0x4f
      13'h150: dout <= 8'b01000100; //  336 :  68 - 0x44 -- Sprite 0x15
      13'h151: dout <= 8'b01000100; //  337 :  68 - 0x44
      13'h152: dout <= 8'b01000100; //  338 :  68 - 0x44
      13'h153: dout <= 8'b01000100; //  339 :  68 - 0x44
      13'h154: dout <= 8'b01000100; //  340 :  68 - 0x44
      13'h155: dout <= 8'b01011100; //  341 :  92 - 0x5c
      13'h156: dout <= 8'b01000000; //  342 :  64 - 0x40
      13'h157: dout <= 8'b00000000; //  343 :   0 - 0x0
      13'h158: dout <= 8'b01100110; //  344 : 102 - 0x66
      13'h159: dout <= 8'b01100110; //  345 : 102 - 0x66
      13'h15A: dout <= 8'b01100110; //  346 : 102 - 0x66
      13'h15B: dout <= 8'b01100110; //  347 : 102 - 0x66
      13'h15C: dout <= 8'b01100110; //  348 : 102 - 0x66
      13'h15D: dout <= 8'b01111110; //  349 : 126 - 0x7e
      13'h15E: dout <= 8'b01111110; //  350 : 126 - 0x7e
      13'h15F: dout <= 8'b00000000; //  351 :   0 - 0x0
      13'h160: dout <= 8'b01000000; //  352 :  64 - 0x40 -- Sprite 0x16
      13'h161: dout <= 8'b01000000; //  353 :  64 - 0x40
      13'h162: dout <= 8'b00000000; //  354 :   0 - 0x0
      13'h163: dout <= 8'b00000000; //  355 :   0 - 0x0
      13'h164: dout <= 8'b00011000; //  356 :  24 - 0x18
      13'h165: dout <= 8'b00111000; //  357 :  56 - 0x38
      13'h166: dout <= 8'b00010000; //  358 :  16 - 0x10
      13'h167: dout <= 8'b00000000; //  359 :   0 - 0x0
      13'h168: dout <= 8'b01111110; //  360 : 126 - 0x7e
      13'h169: dout <= 8'b01100110; //  361 : 102 - 0x66
      13'h16A: dout <= 8'b01000010; //  362 :  66 - 0x42
      13'h16B: dout <= 8'b00011000; //  363 :  24 - 0x18
      13'h16C: dout <= 8'b00111100; //  364 :  60 - 0x3c
      13'h16D: dout <= 8'b01111110; //  365 : 126 - 0x7e
      13'h16E: dout <= 8'b11111111; //  366 : 255 - 0xff
      13'h16F: dout <= 8'b11111111; //  367 : 255 - 0xff
      13'h170: dout <= 8'b01000000; //  368 :  64 - 0x40 -- Sprite 0x17
      13'h171: dout <= 8'b01000000; //  369 :  64 - 0x40
      13'h172: dout <= 8'b01000000; //  370 :  64 - 0x40
      13'h173: dout <= 8'b01000000; //  371 :  64 - 0x40
      13'h174: dout <= 8'b01010000; //  372 :  80 - 0x50
      13'h175: dout <= 8'b01010000; //  373 :  80 - 0x50
      13'h176: dout <= 8'b01001000; //  374 :  72 - 0x48
      13'h177: dout <= 8'b01001000; //  375 :  72 - 0x48
      13'h178: dout <= 8'b01101111; //  376 : 111 - 0x6f
      13'h179: dout <= 8'b01100111; //  377 : 103 - 0x67
      13'h17A: dout <= 8'b01110111; //  378 : 119 - 0x77
      13'h17B: dout <= 8'b01110011; //  379 : 115 - 0x73
      13'h17C: dout <= 8'b01111011; //  380 : 123 - 0x7b
      13'h17D: dout <= 8'b01111001; //  381 : 121 - 0x79
      13'h17E: dout <= 8'b01101101; //  382 : 109 - 0x6d
      13'h17F: dout <= 8'b01101100; //  383 : 108 - 0x6c
      13'h180: dout <= 8'b01000111; //  384 :  71 - 0x47 -- Sprite 0x18
      13'h181: dout <= 8'b01000111; //  385 :  71 - 0x47
      13'h182: dout <= 8'b01000111; //  386 :  71 - 0x47
      13'h183: dout <= 8'b01000111; //  387 :  71 - 0x47
      13'h184: dout <= 8'b01000111; //  388 :  71 - 0x47
      13'h185: dout <= 8'b01011111; //  389 :  95 - 0x5f
      13'h186: dout <= 8'b00000000; //  390 :   0 - 0x0
      13'h187: dout <= 8'b00000000; //  391 :   0 - 0x0
      13'h188: dout <= 8'b01100000; //  392 :  96 - 0x60
      13'h189: dout <= 8'b01100000; //  393 :  96 - 0x60
      13'h18A: dout <= 8'b01100000; //  394 :  96 - 0x60
      13'h18B: dout <= 8'b01100000; //  395 :  96 - 0x60
      13'h18C: dout <= 8'b01100000; //  396 :  96 - 0x60
      13'h18D: dout <= 8'b01111111; //  397 : 127 - 0x7f
      13'h18E: dout <= 8'b01111111; //  398 : 127 - 0x7f
      13'h18F: dout <= 8'b00000000; //  399 :   0 - 0x0
      13'h190: dout <= 8'b11111100; //  400 : 252 - 0xfc -- Sprite 0x19
      13'h191: dout <= 8'b11111100; //  401 : 252 - 0xfc
      13'h192: dout <= 8'b11111100; //  402 : 252 - 0xfc
      13'h193: dout <= 8'b11111100; //  403 : 252 - 0xfc
      13'h194: dout <= 8'b11111100; //  404 : 252 - 0xfc
      13'h195: dout <= 8'b11011100; //  405 : 220 - 0xdc
      13'h196: dout <= 8'b00011100; //  406 :  28 - 0x1c
      13'h197: dout <= 8'b01000100; //  407 :  68 - 0x44
      13'h198: dout <= 8'b00000110; //  408 :   6 - 0x6
      13'h199: dout <= 8'b00000110; //  409 :   6 - 0x6
      13'h19A: dout <= 8'b00000110; //  410 :   6 - 0x6
      13'h19B: dout <= 8'b00000110; //  411 :   6 - 0x6
      13'h19C: dout <= 8'b00000110; //  412 :   6 - 0x6
      13'h19D: dout <= 8'b11100110; //  413 : 230 - 0xe6
      13'h19E: dout <= 8'b11100110; //  414 : 230 - 0xe6
      13'h19F: dout <= 8'b01100110; //  415 : 102 - 0x66
      13'h1A0: dout <= 8'b00010000; //  416 :  16 - 0x10 -- Sprite 0x1a
      13'h1A1: dout <= 8'b00111000; //  417 :  56 - 0x38
      13'h1A2: dout <= 8'b01111100; //  418 : 124 - 0x7c
      13'h1A3: dout <= 8'b11100000; //  419 : 224 - 0xe0
      13'h1A4: dout <= 8'b01000000; //  420 :  64 - 0x40
      13'h1A5: dout <= 8'b00000000; //  421 :   0 - 0x0
      13'h1A6: dout <= 8'b00010000; //  422 :  16 - 0x10
      13'h1A7: dout <= 8'b00100000; //  423 :  32 - 0x20
      13'h1A8: dout <= 8'b11111111; //  424 : 255 - 0xff
      13'h1A9: dout <= 8'b11111111; //  425 : 255 - 0xff
      13'h1AA: dout <= 8'b11111111; //  426 : 255 - 0xff
      13'h1AB: dout <= 8'b11111111; //  427 : 255 - 0xff
      13'h1AC: dout <= 8'b11100111; //  428 : 231 - 0xe7
      13'h1AD: dout <= 8'b11000011; //  429 : 195 - 0xc3
      13'h1AE: dout <= 8'b10011001; //  430 : 153 - 0x99
      13'h1AF: dout <= 8'b00111100; //  431 :  60 - 0x3c
      13'h1B0: dout <= 8'b00000000; //  432 :   0 - 0x0 -- Sprite 0x1b
      13'h1B1: dout <= 8'b01111100; //  433 : 124 - 0x7c
      13'h1B2: dout <= 8'b01000000; //  434 :  64 - 0x40
      13'h1B3: dout <= 8'b01000100; //  435 :  68 - 0x44
      13'h1B4: dout <= 8'b01000100; //  436 :  68 - 0x44
      13'h1B5: dout <= 8'b01000100; //  437 :  68 - 0x44
      13'h1B6: dout <= 8'b01000100; //  438 :  68 - 0x44
      13'h1B7: dout <= 8'b01000100; //  439 :  68 - 0x44
      13'h1B8: dout <= 8'b00000000; //  440 :   0 - 0x0
      13'h1B9: dout <= 8'b01111110; //  441 : 126 - 0x7e
      13'h1BA: dout <= 8'b01111110; //  442 : 126 - 0x7e
      13'h1BB: dout <= 8'b01100110; //  443 : 102 - 0x66
      13'h1BC: dout <= 8'b01100110; //  444 : 102 - 0x66
      13'h1BD: dout <= 8'b01100110; //  445 : 102 - 0x66
      13'h1BE: dout <= 8'b01100110; //  446 : 102 - 0x66
      13'h1BF: dout <= 8'b01100110; //  447 : 102 - 0x66
      13'h1C0: dout <= 8'b00010000; //  448 :  16 - 0x10 -- Sprite 0x1c
      13'h1C1: dout <= 8'b00111000; //  449 :  56 - 0x38
      13'h1C2: dout <= 8'b01110001; //  450 : 113 - 0x71
      13'h1C3: dout <= 8'b11100010; //  451 : 226 - 0xe2
      13'h1C4: dout <= 8'b01000100; //  452 :  68 - 0x44
      13'h1C5: dout <= 8'b00001000; //  453 :   8 - 0x8
      13'h1C6: dout <= 8'b00010000; //  454 :  16 - 0x10
      13'h1C7: dout <= 8'b00100000; //  455 :  32 - 0x20
      13'h1C8: dout <= 8'b11111110; //  456 : 254 - 0xfe
      13'h1C9: dout <= 8'b11111100; //  457 : 252 - 0xfc
      13'h1CA: dout <= 8'b11111001; //  458 : 249 - 0xf9
      13'h1CB: dout <= 8'b11110011; //  459 : 243 - 0xf3
      13'h1CC: dout <= 8'b11100111; //  460 : 231 - 0xe7
      13'h1CD: dout <= 8'b11001110; //  461 : 206 - 0xce
      13'h1CE: dout <= 8'b10011100; //  462 : 156 - 0x9c
      13'h1CF: dout <= 8'b00111000; //  463 :  56 - 0x38
      13'h1D0: dout <= 8'b01000000; //  464 :  64 - 0x40 -- Sprite 0x1d
      13'h1D1: dout <= 8'b10000100; //  465 : 132 - 0x84
      13'h1D2: dout <= 8'b00000010; //  466 :   2 - 0x2
      13'h1D3: dout <= 8'b00000111; //  467 :   7 - 0x7
      13'h1D4: dout <= 8'b00001111; //  468 :  15 - 0xf
      13'h1D5: dout <= 8'b00011111; //  469 :  31 - 0x1f
      13'h1D6: dout <= 8'b00111111; //  470 :  63 - 0x3f
      13'h1D7: dout <= 8'b01111111; //  471 : 127 - 0x7f
      13'h1D8: dout <= 8'b01111110; //  472 : 126 - 0x7e
      13'h1D9: dout <= 8'b11100111; //  473 : 231 - 0xe7
      13'h1DA: dout <= 8'b11000011; //  474 : 195 - 0xc3
      13'h1DB: dout <= 8'b10000001; //  475 : 129 - 0x81
      13'h1DC: dout <= 8'b00000000; //  476 :   0 - 0x0
      13'h1DD: dout <= 8'b00000000; //  477 :   0 - 0x0
      13'h1DE: dout <= 8'b00000000; //  478 :   0 - 0x0
      13'h1DF: dout <= 8'b00000000; //  479 :   0 - 0x0
      13'h1E0: dout <= 8'b00010000; //  480 :  16 - 0x10 -- Sprite 0x1e
      13'h1E1: dout <= 8'b00011000; //  481 :  24 - 0x18
      13'h1E2: dout <= 8'b00001100; //  482 :  12 - 0xc
      13'h1E3: dout <= 8'b00000110; //  483 :   6 - 0x6
      13'h1E4: dout <= 8'b10000000; //  484 : 128 - 0x80
      13'h1E5: dout <= 8'b11000000; //  485 : 192 - 0xc0
      13'h1E6: dout <= 8'b11100000; //  486 : 224 - 0xe0
      13'h1E7: dout <= 8'b11110000; //  487 : 240 - 0xf0
      13'h1E8: dout <= 8'b01111111; //  488 : 127 - 0x7f
      13'h1E9: dout <= 8'b00111111; //  489 :  63 - 0x3f
      13'h1EA: dout <= 8'b10011111; //  490 : 159 - 0x9f
      13'h1EB: dout <= 8'b11001111; //  491 : 207 - 0xcf
      13'h1EC: dout <= 8'b11100111; //  492 : 231 - 0xe7
      13'h1ED: dout <= 8'b01110011; //  493 : 115 - 0x73
      13'h1EE: dout <= 8'b00111001; //  494 :  57 - 0x39
      13'h1EF: dout <= 8'b00011100; //  495 :  28 - 0x1c
      13'h1F0: dout <= 8'b11111100; //  496 : 252 - 0xfc -- Sprite 0x1f
      13'h1F1: dout <= 8'b11111101; //  497 : 253 - 0xfd
      13'h1F2: dout <= 8'b11111100; //  498 : 252 - 0xfc
      13'h1F3: dout <= 8'b11111110; //  499 : 254 - 0xfe
      13'h1F4: dout <= 8'b11111110; //  500 : 254 - 0xfe
      13'h1F5: dout <= 8'b11111111; //  501 : 255 - 0xff
      13'h1F6: dout <= 8'b11111111; //  502 : 255 - 0xff
      13'h1F7: dout <= 8'b11111111; //  503 : 255 - 0xff
      13'h1F8: dout <= 8'b00000110; //  504 :   6 - 0x6
      13'h1F9: dout <= 8'b00000111; //  505 :   7 - 0x7
      13'h1FA: dout <= 8'b00000111; //  506 :   7 - 0x7
      13'h1FB: dout <= 8'b00000000; //  507 :   0 - 0x0
      13'h1FC: dout <= 8'b00000000; //  508 :   0 - 0x0
      13'h1FD: dout <= 8'b00000000; //  509 :   0 - 0x0
      13'h1FE: dout <= 8'b00000000; //  510 :   0 - 0x0
      13'h1FF: dout <= 8'b00000000; //  511 :   0 - 0x0
      13'h200: dout <= 8'b00000000; //  512 :   0 - 0x0 -- Sprite 0x20
      13'h201: dout <= 8'b11111111; //  513 : 255 - 0xff
      13'h202: dout <= 8'b00000000; //  514 :   0 - 0x0
      13'h203: dout <= 8'b00000000; //  515 :   0 - 0x0
      13'h204: dout <= 8'b00000000; //  516 :   0 - 0x0
      13'h205: dout <= 8'b11111111; //  517 : 255 - 0xff
      13'h206: dout <= 8'b11111111; //  518 : 255 - 0xff
      13'h207: dout <= 8'b11111111; //  519 : 255 - 0xff
      13'h208: dout <= 8'b00000000; //  520 :   0 - 0x0
      13'h209: dout <= 8'b11111111; //  521 : 255 - 0xff
      13'h20A: dout <= 8'b11111111; //  522 : 255 - 0xff
      13'h20B: dout <= 8'b00000000; //  523 :   0 - 0x0
      13'h20C: dout <= 8'b00000000; //  524 :   0 - 0x0
      13'h20D: dout <= 8'b00000000; //  525 :   0 - 0x0
      13'h20E: dout <= 8'b00000000; //  526 :   0 - 0x0
      13'h20F: dout <= 8'b00000000; //  527 :   0 - 0x0
      13'h210: dout <= 8'b01000100; //  528 :  68 - 0x44 -- Sprite 0x21
      13'h211: dout <= 8'b11000101; //  529 : 197 - 0xc5
      13'h212: dout <= 8'b00000000; //  530 :   0 - 0x0
      13'h213: dout <= 8'b00000110; //  531 :   6 - 0x6
      13'h214: dout <= 8'b00000110; //  532 :   6 - 0x6
      13'h215: dout <= 8'b11111111; //  533 : 255 - 0xff
      13'h216: dout <= 8'b11111111; //  534 : 255 - 0xff
      13'h217: dout <= 8'b11111111; //  535 : 255 - 0xff
      13'h218: dout <= 8'b01100110; //  536 : 102 - 0x66
      13'h219: dout <= 8'b11100111; //  537 : 231 - 0xe7
      13'h21A: dout <= 8'b11100111; //  538 : 231 - 0xe7
      13'h21B: dout <= 8'b00000000; //  539 :   0 - 0x0
      13'h21C: dout <= 8'b00000000; //  540 :   0 - 0x0
      13'h21D: dout <= 8'b00000000; //  541 :   0 - 0x0
      13'h21E: dout <= 8'b00000000; //  542 :   0 - 0x0
      13'h21F: dout <= 8'b00000000; //  543 :   0 - 0x0
      13'h220: dout <= 8'b01000000; //  544 :  64 - 0x40 -- Sprite 0x22
      13'h221: dout <= 8'b10000001; //  545 : 129 - 0x81
      13'h222: dout <= 8'b00000011; //  546 :   3 - 0x3
      13'h223: dout <= 8'b00000111; //  547 :   7 - 0x7
      13'h224: dout <= 8'b00001111; //  548 :  15 - 0xf
      13'h225: dout <= 8'b11111111; //  549 : 255 - 0xff
      13'h226: dout <= 8'b11111111; //  550 : 255 - 0xff
      13'h227: dout <= 8'b11111111; //  551 : 255 - 0xff
      13'h228: dout <= 8'b01110000; //  552 : 112 - 0x70
      13'h229: dout <= 8'b11100000; //  553 : 224 - 0xe0
      13'h22A: dout <= 8'b11000000; //  554 : 192 - 0xc0
      13'h22B: dout <= 8'b00000000; //  555 :   0 - 0x0
      13'h22C: dout <= 8'b00000000; //  556 :   0 - 0x0
      13'h22D: dout <= 8'b00000000; //  557 :   0 - 0x0
      13'h22E: dout <= 8'b00000000; //  558 :   0 - 0x0
      13'h22F: dout <= 8'b00000000; //  559 :   0 - 0x0
      13'h230: dout <= 8'b11111000; //  560 : 248 - 0xf8 -- Sprite 0x23
      13'h231: dout <= 8'b11111100; //  561 : 252 - 0xfc
      13'h232: dout <= 8'b11111110; //  562 : 254 - 0xfe
      13'h233: dout <= 8'b11111110; //  563 : 254 - 0xfe
      13'h234: dout <= 8'b11111111; //  564 : 255 - 0xff
      13'h235: dout <= 8'b11111111; //  565 : 255 - 0xff
      13'h236: dout <= 8'b11111111; //  566 : 255 - 0xff
      13'h237: dout <= 8'b11111111; //  567 : 255 - 0xff
      13'h238: dout <= 8'b00001110; //  568 :  14 - 0xe
      13'h239: dout <= 8'b00000111; //  569 :   7 - 0x7
      13'h23A: dout <= 8'b00000011; //  570 :   3 - 0x3
      13'h23B: dout <= 8'b00000000; //  571 :   0 - 0x0
      13'h23C: dout <= 8'b00000000; //  572 :   0 - 0x0
      13'h23D: dout <= 8'b00000000; //  573 :   0 - 0x0
      13'h23E: dout <= 8'b00000000; //  574 :   0 - 0x0
      13'h23F: dout <= 8'b00000000; //  575 :   0 - 0x0
      13'h240: dout <= 8'b01000111; //  576 :  71 - 0x47 -- Sprite 0x24
      13'h241: dout <= 8'b11000111; //  577 : 199 - 0xc7
      13'h242: dout <= 8'b00000111; //  578 :   7 - 0x7
      13'h243: dout <= 8'b00000111; //  579 :   7 - 0x7
      13'h244: dout <= 8'b00000111; //  580 :   7 - 0x7
      13'h245: dout <= 8'b11111111; //  581 : 255 - 0xff
      13'h246: dout <= 8'b11111111; //  582 : 255 - 0xff
      13'h247: dout <= 8'b11111111; //  583 : 255 - 0xff
      13'h248: dout <= 8'b01100000; //  584 :  96 - 0x60
      13'h249: dout <= 8'b11100000; //  585 : 224 - 0xe0
      13'h24A: dout <= 8'b11100000; //  586 : 224 - 0xe0
      13'h24B: dout <= 8'b00000000; //  587 :   0 - 0x0
      13'h24C: dout <= 8'b00000000; //  588 :   0 - 0x0
      13'h24D: dout <= 8'b00000000; //  589 :   0 - 0x0
      13'h24E: dout <= 8'b00000000; //  590 :   0 - 0x0
      13'h24F: dout <= 8'b00000000; //  591 :   0 - 0x0
      13'h250: dout <= 8'b11111111; //  592 : 255 - 0xff -- Sprite 0x25
      13'h251: dout <= 8'b11111111; //  593 : 255 - 0xff
      13'h252: dout <= 8'b11111111; //  594 : 255 - 0xff
      13'h253: dout <= 8'b11111111; //  595 : 255 - 0xff
      13'h254: dout <= 8'b11111111; //  596 : 255 - 0xff
      13'h255: dout <= 8'b11111111; //  597 : 255 - 0xff
      13'h256: dout <= 8'b00011111; //  598 :  31 - 0x1f
      13'h257: dout <= 8'b00001111; //  599 :  15 - 0xf
      13'h258: dout <= 8'b00000000; //  600 :   0 - 0x0
      13'h259: dout <= 8'b00000000; //  601 :   0 - 0x0
      13'h25A: dout <= 8'b00000000; //  602 :   0 - 0x0
      13'h25B: dout <= 8'b00000000; //  603 :   0 - 0x0
      13'h25C: dout <= 8'b00000000; //  604 :   0 - 0x0
      13'h25D: dout <= 8'b11000000; //  605 : 192 - 0xc0
      13'h25E: dout <= 8'b11100000; //  606 : 224 - 0xe0
      13'h25F: dout <= 8'b01110000; //  607 : 112 - 0x70
      13'h260: dout <= 8'b11111111; //  608 : 255 - 0xff -- Sprite 0x26
      13'h261: dout <= 8'b11111111; //  609 : 255 - 0xff
      13'h262: dout <= 8'b11111111; //  610 : 255 - 0xff
      13'h263: dout <= 8'b11111111; //  611 : 255 - 0xff
      13'h264: dout <= 8'b11111111; //  612 : 255 - 0xff
      13'h265: dout <= 8'b11111111; //  613 : 255 - 0xff
      13'h266: dout <= 8'b11111100; //  614 : 252 - 0xfc
      13'h267: dout <= 8'b11111000; //  615 : 248 - 0xf8
      13'h268: dout <= 8'b00000000; //  616 :   0 - 0x0
      13'h269: dout <= 8'b00000000; //  617 :   0 - 0x0
      13'h26A: dout <= 8'b00000000; //  618 :   0 - 0x0
      13'h26B: dout <= 8'b00000000; //  619 :   0 - 0x0
      13'h26C: dout <= 8'b00000000; //  620 :   0 - 0x0
      13'h26D: dout <= 8'b00000011; //  621 :   3 - 0x3
      13'h26E: dout <= 8'b00000111; //  622 :   7 - 0x7
      13'h26F: dout <= 8'b00001110; //  623 :  14 - 0xe
      13'h270: dout <= 8'b00100111; //  624 :  39 - 0x27 -- Sprite 0x27
      13'h271: dout <= 8'b00010011; //  625 :  19 - 0x13
      13'h272: dout <= 8'b00001001; //  626 :   9 - 0x9
      13'h273: dout <= 8'b11000100; //  627 : 196 - 0xc4
      13'h274: dout <= 8'b01100010; //  628 :  98 - 0x62
      13'h275: dout <= 8'b00100001; //  629 :  33 - 0x21
      13'h276: dout <= 8'b00000000; //  630 :   0 - 0x0
      13'h277: dout <= 8'b00000000; //  631 :   0 - 0x0
      13'h278: dout <= 8'b00111000; //  632 :  56 - 0x38
      13'h279: dout <= 8'b10011100; //  633 : 156 - 0x9c
      13'h27A: dout <= 8'b11001110; //  634 : 206 - 0xce
      13'h27B: dout <= 8'b11100111; //  635 : 231 - 0xe7
      13'h27C: dout <= 8'b11110011; //  636 : 243 - 0xf3
      13'h27D: dout <= 8'b11111001; //  637 : 249 - 0xf9
      13'h27E: dout <= 8'b11111100; //  638 : 252 - 0xfc
      13'h27F: dout <= 8'b11111110; //  639 : 254 - 0xfe
      13'h280: dout <= 8'b11111111; //  640 : 255 - 0xff -- Sprite 0x28
      13'h281: dout <= 8'b11111111; //  641 : 255 - 0xff
      13'h282: dout <= 8'b11111111; //  642 : 255 - 0xff
      13'h283: dout <= 8'b11111111; //  643 : 255 - 0xff
      13'h284: dout <= 8'b01111111; //  644 : 127 - 0x7f
      13'h285: dout <= 8'b00111110; //  645 :  62 - 0x3e
      13'h286: dout <= 8'b10011100; //  646 : 156 - 0x9c
      13'h287: dout <= 8'b01001000; //  647 :  72 - 0x48
      13'h288: dout <= 8'b00000000; //  648 :   0 - 0x0
      13'h289: dout <= 8'b00000000; //  649 :   0 - 0x0
      13'h28A: dout <= 8'b00000000; //  650 :   0 - 0x0
      13'h28B: dout <= 8'b00000000; //  651 :   0 - 0x0
      13'h28C: dout <= 8'b10000001; //  652 : 129 - 0x81
      13'h28D: dout <= 8'b11000011; //  653 : 195 - 0xc3
      13'h28E: dout <= 8'b11100111; //  654 : 231 - 0xe7
      13'h28F: dout <= 8'b01111110; //  655 : 126 - 0x7e
      13'h290: dout <= 8'b11110000; //  656 : 240 - 0xf0 -- Sprite 0x29
      13'h291: dout <= 8'b11100000; //  657 : 224 - 0xe0
      13'h292: dout <= 8'b11000000; //  658 : 192 - 0xc0
      13'h293: dout <= 8'b10000000; //  659 : 128 - 0x80
      13'h294: dout <= 8'b00000000; //  660 :   0 - 0x0
      13'h295: dout <= 8'b00000010; //  661 :   2 - 0x2
      13'h296: dout <= 8'b00000101; //  662 :   5 - 0x5
      13'h297: dout <= 8'b00000010; //  663 :   2 - 0x2
      13'h298: dout <= 8'b00011100; //  664 :  28 - 0x1c
      13'h299: dout <= 8'b00111001; //  665 :  57 - 0x39
      13'h29A: dout <= 8'b01110011; //  666 : 115 - 0x73
      13'h29B: dout <= 8'b11100111; //  667 : 231 - 0xe7
      13'h29C: dout <= 8'b11001111; //  668 : 207 - 0xcf
      13'h29D: dout <= 8'b10011111; //  669 : 159 - 0x9f
      13'h29E: dout <= 8'b00111111; //  670 :  63 - 0x3f
      13'h29F: dout <= 8'b01111111; //  671 : 127 - 0x7f
      13'h2A0: dout <= 8'b01000111; //  672 :  71 - 0x47 -- Sprite 0x2a
      13'h2A1: dout <= 8'b01000110; //  673 :  70 - 0x46
      13'h2A2: dout <= 8'b01000110; //  674 :  70 - 0x46
      13'h2A3: dout <= 8'b01000100; //  675 :  68 - 0x44
      13'h2A4: dout <= 8'b01000100; //  676 :  68 - 0x44
      13'h2A5: dout <= 8'b01000100; //  677 :  68 - 0x44
      13'h2A6: dout <= 8'b01000100; //  678 :  68 - 0x44
      13'h2A7: dout <= 8'b01000100; //  679 :  68 - 0x44
      13'h2A8: dout <= 8'b01100001; //  680 :  97 - 0x61
      13'h2A9: dout <= 8'b01100011; //  681 :  99 - 0x63
      13'h2AA: dout <= 8'b01100011; //  682 :  99 - 0x63
      13'h2AB: dout <= 8'b01100111; //  683 : 103 - 0x67
      13'h2AC: dout <= 8'b01100110; //  684 : 102 - 0x66
      13'h2AD: dout <= 8'b01100110; //  685 : 102 - 0x66
      13'h2AE: dout <= 8'b01100110; //  686 : 102 - 0x66
      13'h2AF: dout <= 8'b01100110; //  687 : 102 - 0x66
      13'h2B0: dout <= 8'b01111111; //  688 : 127 - 0x7f -- Sprite 0x2b
      13'h2B1: dout <= 8'b00111111; //  689 :  63 - 0x3f
      13'h2B2: dout <= 8'b10011111; //  690 : 159 - 0x9f
      13'h2B3: dout <= 8'b10001111; //  691 : 143 - 0x8f
      13'h2B4: dout <= 8'b01001111; //  692 :  79 - 0x4f
      13'h2B5: dout <= 8'b01000111; //  693 :  71 - 0x47
      13'h2B6: dout <= 8'b01000111; //  694 :  71 - 0x47
      13'h2B7: dout <= 8'b01000111; //  695 :  71 - 0x47
      13'h2B8: dout <= 8'b10000000; //  696 : 128 - 0x80
      13'h2B9: dout <= 8'b11000000; //  697 : 192 - 0xc0
      13'h2BA: dout <= 8'b11000000; //  698 : 192 - 0xc0
      13'h2BB: dout <= 8'b11100000; //  699 : 224 - 0xe0
      13'h2BC: dout <= 8'b01100000; //  700 :  96 - 0x60
      13'h2BD: dout <= 8'b01100000; //  701 :  96 - 0x60
      13'h2BE: dout <= 8'b01100000; //  702 :  96 - 0x60
      13'h2BF: dout <= 8'b01100000; //  703 :  96 - 0x60
      13'h2C0: dout <= 8'b00100000; //  704 :  32 - 0x20 -- Sprite 0x2c
      13'h2C1: dout <= 8'b00010000; //  705 :  16 - 0x10
      13'h2C2: dout <= 8'b00000000; //  706 :   0 - 0x0
      13'h2C3: dout <= 8'b11000000; //  707 : 192 - 0xc0
      13'h2C4: dout <= 8'b01100000; //  708 :  96 - 0x60
      13'h2C5: dout <= 8'b00100010; //  709 :  34 - 0x22
      13'h2C6: dout <= 8'b00000101; //  710 :   5 - 0x5
      13'h2C7: dout <= 8'b00000010; //  711 :   2 - 0x2
      13'h2C8: dout <= 8'b00111100; //  712 :  60 - 0x3c
      13'h2C9: dout <= 8'b10011001; //  713 : 153 - 0x99
      13'h2CA: dout <= 8'b11000011; //  714 : 195 - 0xc3
      13'h2CB: dout <= 8'b11100111; //  715 : 231 - 0xe7
      13'h2CC: dout <= 8'b11111111; //  716 : 255 - 0xff
      13'h2CD: dout <= 8'b11111111; //  717 : 255 - 0xff
      13'h2CE: dout <= 8'b11111111; //  718 : 255 - 0xff
      13'h2CF: dout <= 8'b11111111; //  719 : 255 - 0xff
      13'h2D0: dout <= 8'b00000000; //  720 :   0 - 0x0 -- Sprite 0x2d
      13'h2D1: dout <= 8'b01111111; //  721 : 127 - 0x7f
      13'h2D2: dout <= 8'b01000000; //  722 :  64 - 0x40
      13'h2D3: dout <= 8'b01000000; //  723 :  64 - 0x40
      13'h2D4: dout <= 8'b01000000; //  724 :  64 - 0x40
      13'h2D5: dout <= 8'b01000111; //  725 :  71 - 0x47
      13'h2D6: dout <= 8'b01000111; //  726 :  71 - 0x47
      13'h2D7: dout <= 8'b01000111; //  727 :  71 - 0x47
      13'h2D8: dout <= 8'b00000000; //  728 :   0 - 0x0
      13'h2D9: dout <= 8'b01111111; //  729 : 127 - 0x7f
      13'h2DA: dout <= 8'b01111111; //  730 : 127 - 0x7f
      13'h2DB: dout <= 8'b01100000; //  731 :  96 - 0x60
      13'h2DC: dout <= 8'b01100000; //  732 :  96 - 0x60
      13'h2DD: dout <= 8'b01100000; //  733 :  96 - 0x60
      13'h2DE: dout <= 8'b01100000; //  734 :  96 - 0x60
      13'h2DF: dout <= 8'b01100000; //  735 :  96 - 0x60
      13'h2E0: dout <= 8'b01000100; //  736 :  68 - 0x44 -- Sprite 0x2e
      13'h2E1: dout <= 8'b11000100; //  737 : 196 - 0xc4
      13'h2E2: dout <= 8'b00000100; //  738 :   4 - 0x4
      13'h2E3: dout <= 8'b00000100; //  739 :   4 - 0x4
      13'h2E4: dout <= 8'b00000100; //  740 :   4 - 0x4
      13'h2E5: dout <= 8'b11111100; //  741 : 252 - 0xfc
      13'h2E6: dout <= 8'b11111100; //  742 : 252 - 0xfc
      13'h2E7: dout <= 8'b11111100; //  743 : 252 - 0xfc
      13'h2E8: dout <= 8'b01100110; //  744 : 102 - 0x66
      13'h2E9: dout <= 8'b11100110; //  745 : 230 - 0xe6
      13'h2EA: dout <= 8'b11100110; //  746 : 230 - 0xe6
      13'h2EB: dout <= 8'b00000110; //  747 :   6 - 0x6
      13'h2EC: dout <= 8'b00000110; //  748 :   6 - 0x6
      13'h2ED: dout <= 8'b00000110; //  749 :   6 - 0x6
      13'h2EE: dout <= 8'b00000110; //  750 :   6 - 0x6
      13'h2EF: dout <= 8'b00000110; //  751 :   6 - 0x6
      13'h2F0: dout <= 8'b00000001; //  752 :   1 - 0x1 -- Sprite 0x2f
      13'h2F1: dout <= 8'b01111100; //  753 : 124 - 0x7c
      13'h2F2: dout <= 8'b01000000; //  754 :  64 - 0x40
      13'h2F3: dout <= 8'b01000100; //  755 :  68 - 0x44
      13'h2F4: dout <= 8'b01000100; //  756 :  68 - 0x44
      13'h2F5: dout <= 8'b01000100; //  757 :  68 - 0x44
      13'h2F6: dout <= 8'b01000100; //  758 :  68 - 0x44
      13'h2F7: dout <= 8'b01000100; //  759 :  68 - 0x44
      13'h2F8: dout <= 8'b00000001; //  760 :   1 - 0x1
      13'h2F9: dout <= 8'b01111100; //  761 : 124 - 0x7c
      13'h2FA: dout <= 8'b01111110; //  762 : 126 - 0x7e
      13'h2FB: dout <= 8'b01100110; //  763 : 102 - 0x66
      13'h2FC: dout <= 8'b01100110; //  764 : 102 - 0x66
      13'h2FD: dout <= 8'b01100110; //  765 : 102 - 0x66
      13'h2FE: dout <= 8'b01100110; //  766 : 102 - 0x66
      13'h2FF: dout <= 8'b01100110; //  767 : 102 - 0x66
      13'h300: dout <= 8'b00010000; //  768 :  16 - 0x10 -- Sprite 0x30
      13'h301: dout <= 8'b00111000; //  769 :  56 - 0x38
      13'h302: dout <= 8'b00111100; //  770 :  60 - 0x3c
      13'h303: dout <= 8'b00011000; //  771 :  24 - 0x18
      13'h304: dout <= 8'b00000000; //  772 :   0 - 0x0
      13'h305: dout <= 8'b01000010; //  773 :  66 - 0x42
      13'h306: dout <= 8'b01000100; //  774 :  68 - 0x44
      13'h307: dout <= 8'b01001000; //  775 :  72 - 0x48
      13'h308: dout <= 8'b11111111; //  776 : 255 - 0xff
      13'h309: dout <= 8'b11111111; //  777 : 255 - 0xff
      13'h30A: dout <= 8'b01111110; //  778 : 126 - 0x7e
      13'h30B: dout <= 8'b00111100; //  779 :  60 - 0x3c
      13'h30C: dout <= 8'b00011000; //  780 :  24 - 0x18
      13'h30D: dout <= 8'b01000010; //  781 :  66 - 0x42
      13'h30E: dout <= 8'b01100110; //  782 : 102 - 0x66
      13'h30F: dout <= 8'b01111110; //  783 : 126 - 0x7e
      13'h310: dout <= 8'b01000111; //  784 :  71 - 0x47 -- Sprite 0x31
      13'h311: dout <= 8'b01011111; //  785 :  95 - 0x5f
      13'h312: dout <= 8'b00000000; //  786 :   0 - 0x0
      13'h313: dout <= 8'b00000000; //  787 :   0 - 0x0
      13'h314: dout <= 8'b01110000; //  788 : 112 - 0x70
      13'h315: dout <= 8'b00100010; //  789 :  34 - 0x22
      13'h316: dout <= 8'b00000101; //  790 :   5 - 0x5
      13'h317: dout <= 8'b00000010; //  791 :   2 - 0x2
      13'h318: dout <= 8'b01100000; //  792 :  96 - 0x60
      13'h319: dout <= 8'b01111111; //  793 : 127 - 0x7f
      13'h31A: dout <= 8'b01111111; //  794 : 127 - 0x7f
      13'h31B: dout <= 8'b00000000; //  795 :   0 - 0x0
      13'h31C: dout <= 8'b11111111; //  796 : 255 - 0xff
      13'h31D: dout <= 8'b11111111; //  797 : 255 - 0xff
      13'h31E: dout <= 8'b11111111; //  798 : 255 - 0xff
      13'h31F: dout <= 8'b11111111; //  799 : 255 - 0xff
      13'h320: dout <= 8'b11111111; //  800 : 255 - 0xff -- Sprite 0x32
      13'h321: dout <= 8'b11111111; //  801 : 255 - 0xff
      13'h322: dout <= 8'b00000000; //  802 :   0 - 0x0
      13'h323: dout <= 8'b00000000; //  803 :   0 - 0x0
      13'h324: dout <= 8'b01110000; //  804 : 112 - 0x70
      13'h325: dout <= 8'b00100010; //  805 :  34 - 0x22
      13'h326: dout <= 8'b00000101; //  806 :   5 - 0x5
      13'h327: dout <= 8'b00000010; //  807 :   2 - 0x2
      13'h328: dout <= 8'b00000000; //  808 :   0 - 0x0
      13'h329: dout <= 8'b11111111; //  809 : 255 - 0xff
      13'h32A: dout <= 8'b11111111; //  810 : 255 - 0xff
      13'h32B: dout <= 8'b00000000; //  811 :   0 - 0x0
      13'h32C: dout <= 8'b11111111; //  812 : 255 - 0xff
      13'h32D: dout <= 8'b11111111; //  813 : 255 - 0xff
      13'h32E: dout <= 8'b11111111; //  814 : 255 - 0xff
      13'h32F: dout <= 8'b11111111; //  815 : 255 - 0xff
      13'h330: dout <= 8'b11111111; //  816 : 255 - 0xff -- Sprite 0x33
      13'h331: dout <= 8'b11011111; //  817 : 223 - 0xdf
      13'h332: dout <= 8'b00011111; //  818 :  31 - 0x1f
      13'h333: dout <= 8'b01000111; //  819 :  71 - 0x47
      13'h334: dout <= 8'b01000111; //  820 :  71 - 0x47
      13'h335: dout <= 8'b01000111; //  821 :  71 - 0x47
      13'h336: dout <= 8'b01000111; //  822 :  71 - 0x47
      13'h337: dout <= 8'b01000111; //  823 :  71 - 0x47
      13'h338: dout <= 8'b00000000; //  824 :   0 - 0x0
      13'h339: dout <= 8'b11100000; //  825 : 224 - 0xe0
      13'h33A: dout <= 8'b11100000; //  826 : 224 - 0xe0
      13'h33B: dout <= 8'b01100000; //  827 :  96 - 0x60
      13'h33C: dout <= 8'b01100000; //  828 :  96 - 0x60
      13'h33D: dout <= 8'b01100000; //  829 :  96 - 0x60
      13'h33E: dout <= 8'b01100000; //  830 :  96 - 0x60
      13'h33F: dout <= 8'b01100000; //  831 :  96 - 0x60
      13'h340: dout <= 8'b01000100; //  832 :  68 - 0x44 -- Sprite 0x34
      13'h341: dout <= 8'b01000100; //  833 :  68 - 0x44
      13'h342: dout <= 8'b01000100; //  834 :  68 - 0x44
      13'h343: dout <= 8'b01000100; //  835 :  68 - 0x44
      13'h344: dout <= 8'b01000100; //  836 :  68 - 0x44
      13'h345: dout <= 8'b01000100; //  837 :  68 - 0x44
      13'h346: dout <= 8'b01000100; //  838 :  68 - 0x44
      13'h347: dout <= 8'b01000100; //  839 :  68 - 0x44
      13'h348: dout <= 8'b01111110; //  840 : 126 - 0x7e
      13'h349: dout <= 8'b01100110; //  841 : 102 - 0x66
      13'h34A: dout <= 8'b01100110; //  842 : 102 - 0x66
      13'h34B: dout <= 8'b01100110; //  843 : 102 - 0x66
      13'h34C: dout <= 8'b01100110; //  844 : 102 - 0x66
      13'h34D: dout <= 8'b01100110; //  845 : 102 - 0x66
      13'h34E: dout <= 8'b01100110; //  846 : 102 - 0x66
      13'h34F: dout <= 8'b01100110; //  847 : 102 - 0x66
      13'h350: dout <= 8'b00010000; //  848 :  16 - 0x10 -- Sprite 0x35
      13'h351: dout <= 8'b00111000; //  849 :  56 - 0x38
      13'h352: dout <= 8'b01111100; //  850 : 124 - 0x7c
      13'h353: dout <= 8'b11111000; //  851 : 248 - 0xf8
      13'h354: dout <= 8'b00000000; //  852 :   0 - 0x0
      13'h355: dout <= 8'b01111111; //  853 : 127 - 0x7f
      13'h356: dout <= 8'b01000000; //  854 :  64 - 0x40
      13'h357: dout <= 8'b01000000; //  855 :  64 - 0x40
      13'h358: dout <= 8'b11111111; //  856 : 255 - 0xff
      13'h359: dout <= 8'b11111111; //  857 : 255 - 0xff
      13'h35A: dout <= 8'b11111111; //  858 : 255 - 0xff
      13'h35B: dout <= 8'b11111111; //  859 : 255 - 0xff
      13'h35C: dout <= 8'b00000000; //  860 :   0 - 0x0
      13'h35D: dout <= 8'b01111111; //  861 : 127 - 0x7f
      13'h35E: dout <= 8'b01111111; //  862 : 127 - 0x7f
      13'h35F: dout <= 8'b01100000; //  863 :  96 - 0x60
      13'h360: dout <= 8'b00010000; //  864 :  16 - 0x10 -- Sprite 0x36
      13'h361: dout <= 8'b00111000; //  865 :  56 - 0x38
      13'h362: dout <= 8'b01111100; //  866 : 124 - 0x7c
      13'h363: dout <= 8'b11111000; //  867 : 248 - 0xf8
      13'h364: dout <= 8'b00000000; //  868 :   0 - 0x0
      13'h365: dout <= 8'b11111111; //  869 : 255 - 0xff
      13'h366: dout <= 8'b00000000; //  870 :   0 - 0x0
      13'h367: dout <= 8'b00000000; //  871 :   0 - 0x0
      13'h368: dout <= 8'b11111111; //  872 : 255 - 0xff
      13'h369: dout <= 8'b11111111; //  873 : 255 - 0xff
      13'h36A: dout <= 8'b11111111; //  874 : 255 - 0xff
      13'h36B: dout <= 8'b11111111; //  875 : 255 - 0xff
      13'h36C: dout <= 8'b00000000; //  876 :   0 - 0x0
      13'h36D: dout <= 8'b11111111; //  877 : 255 - 0xff
      13'h36E: dout <= 8'b11111111; //  878 : 255 - 0xff
      13'h36F: dout <= 8'b00000000; //  879 :   0 - 0x0
      13'h370: dout <= 8'b01000111; //  880 :  71 - 0x47 -- Sprite 0x37
      13'h371: dout <= 8'b01000111; //  881 :  71 - 0x47
      13'h372: dout <= 8'b01000111; //  882 :  71 - 0x47
      13'h373: dout <= 8'b01000111; //  883 :  71 - 0x47
      13'h374: dout <= 8'b01000111; //  884 :  71 - 0x47
      13'h375: dout <= 8'b11000111; //  885 : 199 - 0xc7
      13'h376: dout <= 8'b00000111; //  886 :   7 - 0x7
      13'h377: dout <= 8'b00000111; //  887 :   7 - 0x7
      13'h378: dout <= 8'b01100000; //  888 :  96 - 0x60
      13'h379: dout <= 8'b01100000; //  889 :  96 - 0x60
      13'h37A: dout <= 8'b01100000; //  890 :  96 - 0x60
      13'h37B: dout <= 8'b01100000; //  891 :  96 - 0x60
      13'h37C: dout <= 8'b01100000; //  892 :  96 - 0x60
      13'h37D: dout <= 8'b11100000; //  893 : 224 - 0xe0
      13'h37E: dout <= 8'b11100000; //  894 : 224 - 0xe0
      13'h37F: dout <= 8'b00000000; //  895 :   0 - 0x0
      13'h380: dout <= 8'b01000100; //  896 :  68 - 0x44 -- Sprite 0x38
      13'h381: dout <= 8'b01000100; //  897 :  68 - 0x44
      13'h382: dout <= 8'b01000100; //  898 :  68 - 0x44
      13'h383: dout <= 8'b01000100; //  899 :  68 - 0x44
      13'h384: dout <= 8'b01000100; //  900 :  68 - 0x44
      13'h385: dout <= 8'b01011000; //  901 :  88 - 0x58
      13'h386: dout <= 8'b00000000; //  902 :   0 - 0x0
      13'h387: dout <= 8'b00000000; //  903 :   0 - 0x0
      13'h388: dout <= 8'b01100110; //  904 : 102 - 0x66
      13'h389: dout <= 8'b01100110; //  905 : 102 - 0x66
      13'h38A: dout <= 8'b01100110; //  906 : 102 - 0x66
      13'h38B: dout <= 8'b01100110; //  907 : 102 - 0x66
      13'h38C: dout <= 8'b01100110; //  908 : 102 - 0x66
      13'h38D: dout <= 8'b01111110; //  909 : 126 - 0x7e
      13'h38E: dout <= 8'b01111100; //  910 : 124 - 0x7c
      13'h38F: dout <= 8'b00000001; //  911 :   1 - 0x1
      13'h390: dout <= 8'b00010000; //  912 :  16 - 0x10 -- Sprite 0x39
      13'h391: dout <= 8'b00111000; //  913 :  56 - 0x38
      13'h392: dout <= 8'b01111100; //  914 : 124 - 0x7c
      13'h393: dout <= 8'b11111000; //  915 : 248 - 0xf8
      13'h394: dout <= 8'b01110000; //  916 : 112 - 0x70
      13'h395: dout <= 8'b00100010; //  917 :  34 - 0x22
      13'h396: dout <= 8'b00000100; //  918 :   4 - 0x4
      13'h397: dout <= 8'b00000000; //  919 :   0 - 0x0
      13'h398: dout <= 8'b11111111; //  920 : 255 - 0xff
      13'h399: dout <= 8'b11111111; //  921 : 255 - 0xff
      13'h39A: dout <= 8'b11111111; //  922 : 255 - 0xff
      13'h39B: dout <= 8'b11111111; //  923 : 255 - 0xff
      13'h39C: dout <= 8'b11111111; //  924 : 255 - 0xff
      13'h39D: dout <= 8'b11111111; //  925 : 255 - 0xff
      13'h39E: dout <= 8'b11111111; //  926 : 255 - 0xff
      13'h39F: dout <= 8'b11111110; //  927 : 254 - 0xfe
      13'h3A0: dout <= 8'b01000100; //  928 :  68 - 0x44 -- Sprite 0x3a
      13'h3A1: dout <= 8'b01000100; //  929 :  68 - 0x44
      13'h3A2: dout <= 8'b01000100; //  930 :  68 - 0x44
      13'h3A3: dout <= 8'b01000100; //  931 :  68 - 0x44
      13'h3A4: dout <= 8'b01000100; //  932 :  68 - 0x44
      13'h3A5: dout <= 8'b01011000; //  933 :  88 - 0x58
      13'h3A6: dout <= 8'b00000000; //  934 :   0 - 0x0
      13'h3A7: dout <= 8'b00000000; //  935 :   0 - 0x0
      13'h3A8: dout <= 8'b01100110; //  936 : 102 - 0x66
      13'h3A9: dout <= 8'b01100110; //  937 : 102 - 0x66
      13'h3AA: dout <= 8'b01100110; //  938 : 102 - 0x66
      13'h3AB: dout <= 8'b01100110; //  939 : 102 - 0x66
      13'h3AC: dout <= 8'b01100110; //  940 : 102 - 0x66
      13'h3AD: dout <= 8'b01111110; //  941 : 126 - 0x7e
      13'h3AE: dout <= 8'b00111100; //  942 :  60 - 0x3c
      13'h3AF: dout <= 8'b10000001; //  943 : 129 - 0x81
      13'h3B0: dout <= 8'b01000000; //  944 :  64 - 0x40 -- Sprite 0x3b
      13'h3B1: dout <= 8'b01000111; //  945 :  71 - 0x47
      13'h3B2: dout <= 8'b01000111; //  946 :  71 - 0x47
      13'h3B3: dout <= 8'b01000111; //  947 :  71 - 0x47
      13'h3B4: dout <= 8'b01000111; //  948 :  71 - 0x47
      13'h3B5: dout <= 8'b01011111; //  949 :  95 - 0x5f
      13'h3B6: dout <= 8'b00000000; //  950 :   0 - 0x0
      13'h3B7: dout <= 8'b00000000; //  951 :   0 - 0x0
      13'h3B8: dout <= 8'b01100000; //  952 :  96 - 0x60
      13'h3B9: dout <= 8'b01100000; //  953 :  96 - 0x60
      13'h3BA: dout <= 8'b01100000; //  954 :  96 - 0x60
      13'h3BB: dout <= 8'b01100000; //  955 :  96 - 0x60
      13'h3BC: dout <= 8'b01100000; //  956 :  96 - 0x60
      13'h3BD: dout <= 8'b01111111; //  957 : 127 - 0x7f
      13'h3BE: dout <= 8'b01111111; //  958 : 127 - 0x7f
      13'h3BF: dout <= 8'b00000000; //  959 :   0 - 0x0
      13'h3C0: dout <= 8'b00000000; //  960 :   0 - 0x0 -- Sprite 0x3c
      13'h3C1: dout <= 8'b11111111; //  961 : 255 - 0xff
      13'h3C2: dout <= 8'b11111111; //  962 : 255 - 0xff
      13'h3C3: dout <= 8'b11111111; //  963 : 255 - 0xff
      13'h3C4: dout <= 8'b11111111; //  964 : 255 - 0xff
      13'h3C5: dout <= 8'b11111111; //  965 : 255 - 0xff
      13'h3C6: dout <= 8'b00000000; //  966 :   0 - 0x0
      13'h3C7: dout <= 8'b00000000; //  967 :   0 - 0x0
      13'h3C8: dout <= 8'b00000000; //  968 :   0 - 0x0
      13'h3C9: dout <= 8'b00000000; //  969 :   0 - 0x0
      13'h3CA: dout <= 8'b00000000; //  970 :   0 - 0x0
      13'h3CB: dout <= 8'b00000000; //  971 :   0 - 0x0
      13'h3CC: dout <= 8'b00000000; //  972 :   0 - 0x0
      13'h3CD: dout <= 8'b11111111; //  973 : 255 - 0xff
      13'h3CE: dout <= 8'b11111111; //  974 : 255 - 0xff
      13'h3CF: dout <= 8'b00000000; //  975 :   0 - 0x0
      13'h3D0: dout <= 8'b00000111; //  976 :   7 - 0x7 -- Sprite 0x3d
      13'h3D1: dout <= 8'b11111111; //  977 : 255 - 0xff
      13'h3D2: dout <= 8'b11111111; //  978 : 255 - 0xff
      13'h3D3: dout <= 8'b11111111; //  979 : 255 - 0xff
      13'h3D4: dout <= 8'b11111111; //  980 : 255 - 0xff
      13'h3D5: dout <= 8'b11111111; //  981 : 255 - 0xff
      13'h3D6: dout <= 8'b00000000; //  982 :   0 - 0x0
      13'h3D7: dout <= 8'b00000000; //  983 :   0 - 0x0
      13'h3D8: dout <= 8'b00000000; //  984 :   0 - 0x0
      13'h3D9: dout <= 8'b00000000; //  985 :   0 - 0x0
      13'h3DA: dout <= 8'b00000000; //  986 :   0 - 0x0
      13'h3DB: dout <= 8'b00000000; //  987 :   0 - 0x0
      13'h3DC: dout <= 8'b00000000; //  988 :   0 - 0x0
      13'h3DD: dout <= 8'b11111111; //  989 : 255 - 0xff
      13'h3DE: dout <= 8'b11111111; //  990 : 255 - 0xff
      13'h3DF: dout <= 8'b00000000; //  991 :   0 - 0x0
      13'h3E0: dout <= 8'b00010000; //  992 :  16 - 0x10 -- Sprite 0x3e
      13'h3E1: dout <= 8'b00111000; //  993 :  56 - 0x38
      13'h3E2: dout <= 8'b01110001; //  994 : 113 - 0x71
      13'h3E3: dout <= 8'b11100010; //  995 : 226 - 0xe2
      13'h3E4: dout <= 8'b01100010; //  996 :  98 - 0x62
      13'h3E5: dout <= 8'b00100001; //  997 :  33 - 0x21
      13'h3E6: dout <= 8'b00000000; //  998 :   0 - 0x0
      13'h3E7: dout <= 8'b00000000; //  999 :   0 - 0x0
      13'h3E8: dout <= 8'b11111110; // 1000 : 254 - 0xfe
      13'h3E9: dout <= 8'b11111100; // 1001 : 252 - 0xfc
      13'h3EA: dout <= 8'b11111001; // 1002 : 249 - 0xf9
      13'h3EB: dout <= 8'b11110011; // 1003 : 243 - 0xf3
      13'h3EC: dout <= 8'b11110011; // 1004 : 243 - 0xf3
      13'h3ED: dout <= 8'b11111001; // 1005 : 249 - 0xf9
      13'h3EE: dout <= 8'b11111100; // 1006 : 252 - 0xfc
      13'h3EF: dout <= 8'b11111110; // 1007 : 254 - 0xfe
      13'h3F0: dout <= 8'b10000111; // 1008 : 135 - 0x87 -- Sprite 0x3f
      13'h3F1: dout <= 8'b10000111; // 1009 : 135 - 0x87
      13'h3F2: dout <= 8'b00000111; // 1010 :   7 - 0x7
      13'h3F3: dout <= 8'b00001111; // 1011 :  15 - 0xf
      13'h3F4: dout <= 8'b00001111; // 1012 :  15 - 0xf
      13'h3F5: dout <= 8'b00011111; // 1013 :  31 - 0x1f
      13'h3F6: dout <= 8'b10011111; // 1014 : 159 - 0x9f
      13'h3F7: dout <= 8'b10001111; // 1015 : 143 - 0x8f
      13'h3F8: dout <= 8'b11100000; // 1016 : 224 - 0xe0
      13'h3F9: dout <= 8'b11000000; // 1017 : 192 - 0xc0
      13'h3FA: dout <= 8'b11000000; // 1018 : 192 - 0xc0
      13'h3FB: dout <= 8'b10000000; // 1019 : 128 - 0x80
      13'h3FC: dout <= 8'b10000000; // 1020 : 128 - 0x80
      13'h3FD: dout <= 8'b11000000; // 1021 : 192 - 0xc0
      13'h3FE: dout <= 8'b11000000; // 1022 : 192 - 0xc0
      13'h3FF: dout <= 8'b11100000; // 1023 : 224 - 0xe0
      13'h400: dout <= 8'b01000100; // 1024 :  68 - 0x44 -- Sprite 0x40
      13'h401: dout <= 8'b01000100; // 1025 :  68 - 0x44
      13'h402: dout <= 8'b01000100; // 1026 :  68 - 0x44
      13'h403: dout <= 8'b01000100; // 1027 :  68 - 0x44
      13'h404: dout <= 8'b01000100; // 1028 :  68 - 0x44
      13'h405: dout <= 8'b01000110; // 1029 :  70 - 0x46
      13'h406: dout <= 8'b01000110; // 1030 :  70 - 0x46
      13'h407: dout <= 8'b01000111; // 1031 :  71 - 0x47
      13'h408: dout <= 8'b01100110; // 1032 : 102 - 0x66
      13'h409: dout <= 8'b01100110; // 1033 : 102 - 0x66
      13'h40A: dout <= 8'b01100110; // 1034 : 102 - 0x66
      13'h40B: dout <= 8'b01100110; // 1035 : 102 - 0x66
      13'h40C: dout <= 8'b01100111; // 1036 : 103 - 0x67
      13'h40D: dout <= 8'b01100011; // 1037 :  99 - 0x63
      13'h40E: dout <= 8'b01100011; // 1038 :  99 - 0x63
      13'h40F: dout <= 8'b01100001; // 1039 :  97 - 0x61
      13'h410: dout <= 8'b00010000; // 1040 :  16 - 0x10 -- Sprite 0x41
      13'h411: dout <= 8'b00111000; // 1041 :  56 - 0x38
      13'h412: dout <= 8'b01111100; // 1042 : 124 - 0x7c
      13'h413: dout <= 8'b01111000; // 1043 : 120 - 0x78
      13'h414: dout <= 8'b00110000; // 1044 :  48 - 0x30
      13'h415: dout <= 8'b00000010; // 1045 :   2 - 0x2
      13'h416: dout <= 8'b00000101; // 1046 :   5 - 0x5
      13'h417: dout <= 8'b00000010; // 1047 :   2 - 0x2
      13'h418: dout <= 8'b11111111; // 1048 : 255 - 0xff
      13'h419: dout <= 8'b11111111; // 1049 : 255 - 0xff
      13'h41A: dout <= 8'b11111111; // 1050 : 255 - 0xff
      13'h41B: dout <= 8'b01111111; // 1051 : 127 - 0x7f
      13'h41C: dout <= 8'b01111111; // 1052 : 127 - 0x7f
      13'h41D: dout <= 8'b00111111; // 1053 :  63 - 0x3f
      13'h41E: dout <= 8'b10011111; // 1054 : 159 - 0x9f
      13'h41F: dout <= 8'b11000111; // 1055 : 199 - 0xc7
      13'h420: dout <= 8'b00010000; // 1056 :  16 - 0x10 -- Sprite 0x42
      13'h421: dout <= 8'b00111000; // 1057 :  56 - 0x38
      13'h422: dout <= 8'b01111100; // 1058 : 124 - 0x7c
      13'h423: dout <= 8'b11111000; // 1059 : 248 - 0xf8
      13'h424: dout <= 8'b01110000; // 1060 : 112 - 0x70
      13'h425: dout <= 8'b00100000; // 1061 :  32 - 0x20
      13'h426: dout <= 8'b00000001; // 1062 :   1 - 0x1
      13'h427: dout <= 8'b00000010; // 1063 :   2 - 0x2
      13'h428: dout <= 8'b11111111; // 1064 : 255 - 0xff
      13'h429: dout <= 8'b11111111; // 1065 : 255 - 0xff
      13'h42A: dout <= 8'b11111111; // 1066 : 255 - 0xff
      13'h42B: dout <= 8'b11111110; // 1067 : 254 - 0xfe
      13'h42C: dout <= 8'b11111110; // 1068 : 254 - 0xfe
      13'h42D: dout <= 8'b11111100; // 1069 : 252 - 0xfc
      13'h42E: dout <= 8'b11111001; // 1070 : 249 - 0xf9
      13'h42F: dout <= 8'b11100011; // 1071 : 227 - 0xe3
      13'h430: dout <= 8'b01000100; // 1072 :  68 - 0x44 -- Sprite 0x43
      13'h431: dout <= 8'b01000100; // 1073 :  68 - 0x44
      13'h432: dout <= 8'b01000100; // 1074 :  68 - 0x44
      13'h433: dout <= 8'b01000100; // 1075 :  68 - 0x44
      13'h434: dout <= 8'b10000100; // 1076 : 132 - 0x84
      13'h435: dout <= 8'b10000100; // 1077 : 132 - 0x84
      13'h436: dout <= 8'b00000100; // 1078 :   4 - 0x4
      13'h437: dout <= 8'b00001100; // 1079 :  12 - 0xc
      13'h438: dout <= 8'b01100110; // 1080 : 102 - 0x66
      13'h439: dout <= 8'b01100110; // 1081 : 102 - 0x66
      13'h43A: dout <= 8'b01100110; // 1082 : 102 - 0x66
      13'h43B: dout <= 8'b01100110; // 1083 : 102 - 0x66
      13'h43C: dout <= 8'b11100110; // 1084 : 230 - 0xe6
      13'h43D: dout <= 8'b11000110; // 1085 : 198 - 0xc6
      13'h43E: dout <= 8'b11000110; // 1086 : 198 - 0xc6
      13'h43F: dout <= 8'b10000110; // 1087 : 134 - 0x86
      13'h440: dout <= 8'b00010000; // 1088 :  16 - 0x10 -- Sprite 0x44
      13'h441: dout <= 8'b00111000; // 1089 :  56 - 0x38
      13'h442: dout <= 8'b01111100; // 1090 : 124 - 0x7c
      13'h443: dout <= 8'b11111000; // 1091 : 248 - 0xf8
      13'h444: dout <= 8'b01110000; // 1092 : 112 - 0x70
      13'h445: dout <= 8'b00100010; // 1093 :  34 - 0x22
      13'h446: dout <= 8'b00000101; // 1094 :   5 - 0x5
      13'h447: dout <= 8'b00000010; // 1095 :   2 - 0x2
      13'h448: dout <= 8'b11111110; // 1096 : 254 - 0xfe
      13'h449: dout <= 8'b11111111; // 1097 : 255 - 0xff
      13'h44A: dout <= 8'b11111111; // 1098 : 255 - 0xff
      13'h44B: dout <= 8'b11111111; // 1099 : 255 - 0xff
      13'h44C: dout <= 8'b11111111; // 1100 : 255 - 0xff
      13'h44D: dout <= 8'b11111111; // 1101 : 255 - 0xff
      13'h44E: dout <= 8'b11111111; // 1102 : 255 - 0xff
      13'h44F: dout <= 8'b11111111; // 1103 : 255 - 0xff
      13'h450: dout <= 8'b01001111; // 1104 :  79 - 0x4f -- Sprite 0x45
      13'h451: dout <= 8'b01000111; // 1105 :  71 - 0x47
      13'h452: dout <= 8'b01000111; // 1106 :  71 - 0x47
      13'h453: dout <= 8'b01000111; // 1107 :  71 - 0x47
      13'h454: dout <= 8'b01000111; // 1108 :  71 - 0x47
      13'h455: dout <= 8'b01000111; // 1109 :  71 - 0x47
      13'h456: dout <= 8'b01000111; // 1110 :  71 - 0x47
      13'h457: dout <= 8'b01000111; // 1111 :  71 - 0x47
      13'h458: dout <= 8'b01100000; // 1112 :  96 - 0x60
      13'h459: dout <= 8'b01100000; // 1113 :  96 - 0x60
      13'h45A: dout <= 8'b01100000; // 1114 :  96 - 0x60
      13'h45B: dout <= 8'b01100000; // 1115 :  96 - 0x60
      13'h45C: dout <= 8'b01100000; // 1116 :  96 - 0x60
      13'h45D: dout <= 8'b01100000; // 1117 :  96 - 0x60
      13'h45E: dout <= 8'b01100000; // 1118 :  96 - 0x60
      13'h45F: dout <= 8'b01100000; // 1119 :  96 - 0x60
      13'h460: dout <= 8'b10100000; // 1120 : 160 - 0xa0 -- Sprite 0x46
      13'h461: dout <= 8'b10011111; // 1121 : 159 - 0x9f
      13'h462: dout <= 8'b11000000; // 1122 : 192 - 0xc0
      13'h463: dout <= 8'b11100000; // 1123 : 224 - 0xe0
      13'h464: dout <= 8'b11111000; // 1124 : 248 - 0xf8
      13'h465: dout <= 8'b11111111; // 1125 : 255 - 0xff
      13'h466: dout <= 8'b11111111; // 1126 : 255 - 0xff
      13'h467: dout <= 8'b11111111; // 1127 : 255 - 0xff
      13'h468: dout <= 8'b11110000; // 1128 : 240 - 0xf0
      13'h469: dout <= 8'b01111111; // 1129 : 127 - 0x7f
      13'h46A: dout <= 8'b00011111; // 1130 :  31 - 0x1f
      13'h46B: dout <= 8'b00000000; // 1131 :   0 - 0x0
      13'h46C: dout <= 8'b00000000; // 1132 :   0 - 0x0
      13'h46D: dout <= 8'b00000000; // 1133 :   0 - 0x0
      13'h46E: dout <= 8'b00000000; // 1134 :   0 - 0x0
      13'h46F: dout <= 8'b00000000; // 1135 :   0 - 0x0
      13'h470: dout <= 8'b00001100; // 1136 :  12 - 0xc -- Sprite 0x47
      13'h471: dout <= 8'b11110000; // 1137 : 240 - 0xf0
      13'h472: dout <= 8'b00000000; // 1138 :   0 - 0x0
      13'h473: dout <= 8'b00000000; // 1139 :   0 - 0x0
      13'h474: dout <= 8'b00000001; // 1140 :   1 - 0x1
      13'h475: dout <= 8'b11111111; // 1141 : 255 - 0xff
      13'h476: dout <= 8'b11111111; // 1142 : 255 - 0xff
      13'h477: dout <= 8'b11111111; // 1143 : 255 - 0xff
      13'h478: dout <= 8'b00001111; // 1144 :  15 - 0xf
      13'h479: dout <= 8'b11111110; // 1145 : 254 - 0xfe
      13'h47A: dout <= 8'b11111000; // 1146 : 248 - 0xf8
      13'h47B: dout <= 8'b00000000; // 1147 :   0 - 0x0
      13'h47C: dout <= 8'b00000000; // 1148 :   0 - 0x0
      13'h47D: dout <= 8'b00000000; // 1149 :   0 - 0x0
      13'h47E: dout <= 8'b00000000; // 1150 :   0 - 0x0
      13'h47F: dout <= 8'b00000000; // 1151 :   0 - 0x0
      13'h480: dout <= 8'b00001100; // 1152 :  12 - 0xc -- Sprite 0x48
      13'h481: dout <= 8'b00011101; // 1153 :  29 - 0x1d
      13'h482: dout <= 8'b00111000; // 1154 :  56 - 0x38
      13'h483: dout <= 8'b01111110; // 1155 : 126 - 0x7e
      13'h484: dout <= 8'b11111110; // 1156 : 254 - 0xfe
      13'h485: dout <= 8'b11111111; // 1157 : 255 - 0xff
      13'h486: dout <= 8'b11111111; // 1158 : 255 - 0xff
      13'h487: dout <= 8'b11111111; // 1159 : 255 - 0xff
      13'h488: dout <= 8'b00000110; // 1160 :   6 - 0x6
      13'h489: dout <= 8'b00000111; // 1161 :   7 - 0x7
      13'h48A: dout <= 8'b00000111; // 1162 :   7 - 0x7
      13'h48B: dout <= 8'b00000000; // 1163 :   0 - 0x0
      13'h48C: dout <= 8'b00000000; // 1164 :   0 - 0x0
      13'h48D: dout <= 8'b00000000; // 1165 :   0 - 0x0
      13'h48E: dout <= 8'b00000000; // 1166 :   0 - 0x0
      13'h48F: dout <= 8'b00000000; // 1167 :   0 - 0x0
      13'h490: dout <= 8'b11111111; // 1168 : 255 - 0xff -- Sprite 0x49
      13'h491: dout <= 8'b11111111; // 1169 : 255 - 0xff
      13'h492: dout <= 8'b11111111; // 1170 : 255 - 0xff
      13'h493: dout <= 8'b11111111; // 1171 : 255 - 0xff
      13'h494: dout <= 8'b11111111; // 1172 : 255 - 0xff
      13'h495: dout <= 8'b11111111; // 1173 : 255 - 0xff
      13'h496: dout <= 8'b11111111; // 1174 : 255 - 0xff
      13'h497: dout <= 8'b11111111; // 1175 : 255 - 0xff
      13'h498: dout <= 8'b00000000; // 1176 :   0 - 0x0
      13'h499: dout <= 8'b00000000; // 1177 :   0 - 0x0
      13'h49A: dout <= 8'b00000000; // 1178 :   0 - 0x0
      13'h49B: dout <= 8'b00000000; // 1179 :   0 - 0x0
      13'h49C: dout <= 8'b00000000; // 1180 :   0 - 0x0
      13'h49D: dout <= 8'b00000000; // 1181 :   0 - 0x0
      13'h49E: dout <= 8'b00000000; // 1182 :   0 - 0x0
      13'h49F: dout <= 8'b00000000; // 1183 :   0 - 0x0
      13'h4A0: dout <= 8'b11111111; // 1184 : 255 - 0xff -- Sprite 0x4a
      13'h4A1: dout <= 8'b11101111; // 1185 : 239 - 0xef
      13'h4A2: dout <= 8'b11111101; // 1186 : 253 - 0xfd
      13'h4A3: dout <= 8'b11111111; // 1187 : 255 - 0xff
      13'h4A4: dout <= 8'b11111111; // 1188 : 255 - 0xff
      13'h4A5: dout <= 8'b11101111; // 1189 : 239 - 0xef
      13'h4A6: dout <= 8'b11111110; // 1190 : 254 - 0xfe
      13'h4A7: dout <= 8'b11111111; // 1191 : 255 - 0xff
      13'h4A8: dout <= 8'b00000000; // 1192 :   0 - 0x0
      13'h4A9: dout <= 8'b01110110; // 1193 : 118 - 0x76
      13'h4AA: dout <= 8'b01010111; // 1194 :  87 - 0x57
      13'h4AB: dout <= 8'b01010101; // 1195 :  85 - 0x55
      13'h4AC: dout <= 8'b01010101; // 1196 :  85 - 0x55
      13'h4AD: dout <= 8'b01110101; // 1197 : 117 - 0x75
      13'h4AE: dout <= 8'b01000111; // 1198 :  71 - 0x47
      13'h4AF: dout <= 8'b00000000; // 1199 :   0 - 0x0
      13'h4B0: dout <= 8'b11111111; // 1200 : 255 - 0xff -- Sprite 0x4b
      13'h4B1: dout <= 8'b11101010; // 1201 : 234 - 0xea
      13'h4B2: dout <= 8'b11111111; // 1202 : 255 - 0xff
      13'h4B3: dout <= 8'b10101111; // 1203 : 175 - 0xaf
      13'h4B4: dout <= 8'b11111111; // 1204 : 255 - 0xff
      13'h4B5: dout <= 8'b11111111; // 1205 : 255 - 0xff
      13'h4B6: dout <= 8'b11111010; // 1206 : 250 - 0xfa
      13'h4B7: dout <= 8'b11111111; // 1207 : 255 - 0xff
      13'h4B8: dout <= 8'b00000000; // 1208 :   0 - 0x0
      13'h4B9: dout <= 8'b01110111; // 1209 : 119 - 0x77
      13'h4BA: dout <= 8'b00010101; // 1210 :  21 - 0x15
      13'h4BB: dout <= 8'b01110101; // 1211 : 117 - 0x75
      13'h4BC: dout <= 8'b01000101; // 1212 :  69 - 0x45
      13'h4BD: dout <= 8'b01000101; // 1213 :  69 - 0x45
      13'h4BE: dout <= 8'b01110111; // 1214 : 119 - 0x77
      13'h4BF: dout <= 8'b00000000; // 1215 :   0 - 0x0
      13'h4C0: dout <= 8'b11111111; // 1216 : 255 - 0xff -- Sprite 0x4c
      13'h4C1: dout <= 8'b11111111; // 1217 : 255 - 0xff
      13'h4C2: dout <= 8'b11111111; // 1218 : 255 - 0xff
      13'h4C3: dout <= 8'b11111111; // 1219 : 255 - 0xff
      13'h4C4: dout <= 8'b11111111; // 1220 : 255 - 0xff
      13'h4C5: dout <= 8'b11111111; // 1221 : 255 - 0xff
      13'h4C6: dout <= 8'b11111110; // 1222 : 254 - 0xfe
      13'h4C7: dout <= 8'b11111111; // 1223 : 255 - 0xff
      13'h4C8: dout <= 8'b00000000; // 1224 :   0 - 0x0
      13'h4C9: dout <= 8'b00100100; // 1225 :  36 - 0x24
      13'h4CA: dout <= 8'b01101100; // 1226 : 108 - 0x6c
      13'h4CB: dout <= 8'b00100100; // 1227 :  36 - 0x24
      13'h4CC: dout <= 8'b00100100; // 1228 :  36 - 0x24
      13'h4CD: dout <= 8'b00100100; // 1229 :  36 - 0x24
      13'h4CE: dout <= 8'b00100101; // 1230 :  37 - 0x25
      13'h4CF: dout <= 8'b00000000; // 1231 :   0 - 0x0
      13'h4D0: dout <= 8'b11111111; // 1232 : 255 - 0xff -- Sprite 0x4d
      13'h4D1: dout <= 8'b10111111; // 1233 : 191 - 0xbf
      13'h4D2: dout <= 8'b11111110; // 1234 : 254 - 0xfe
      13'h4D3: dout <= 8'b10101111; // 1235 : 175 - 0xaf
      13'h4D4: dout <= 8'b11111111; // 1236 : 255 - 0xff
      13'h4D5: dout <= 8'b11111111; // 1237 : 255 - 0xff
      13'h4D6: dout <= 8'b11101111; // 1238 : 239 - 0xef
      13'h4D7: dout <= 8'b11111111; // 1239 : 255 - 0xff
      13'h4D8: dout <= 8'b00000000; // 1240 :   0 - 0x0
      13'h4D9: dout <= 8'b01110100; // 1241 : 116 - 0x74
      13'h4DA: dout <= 8'b01000111; // 1242 :  71 - 0x47
      13'h4DB: dout <= 8'b01110101; // 1243 : 117 - 0x75
      13'h4DC: dout <= 8'b00010101; // 1244 :  21 - 0x15
      13'h4DD: dout <= 8'b00010101; // 1245 :  21 - 0x15
      13'h4DE: dout <= 8'b01110101; // 1246 : 117 - 0x75
      13'h4DF: dout <= 8'b00000000; // 1247 :   0 - 0x0
      13'h4E0: dout <= 8'b11111111; // 1248 : 255 - 0xff -- Sprite 0x4e
      13'h4E1: dout <= 8'b11111111; // 1249 : 255 - 0xff
      13'h4E2: dout <= 8'b11111011; // 1250 : 251 - 0xfb
      13'h4E3: dout <= 8'b11111111; // 1251 : 255 - 0xff
      13'h4E4: dout <= 8'b11111111; // 1252 : 255 - 0xff
      13'h4E5: dout <= 8'b11111111; // 1253 : 255 - 0xff
      13'h4E6: dout <= 8'b11111110; // 1254 : 254 - 0xfe
      13'h4E7: dout <= 8'b11111111; // 1255 : 255 - 0xff
      13'h4E8: dout <= 8'b00000000; // 1256 :   0 - 0x0
      13'h4E9: dout <= 8'b01000000; // 1257 :  64 - 0x40
      13'h4EA: dout <= 8'b00011101; // 1258 :  29 - 0x1d
      13'h4EB: dout <= 8'b01010101; // 1259 :  85 - 0x55
      13'h4EC: dout <= 8'b01010001; // 1260 :  81 - 0x51
      13'h4ED: dout <= 8'b01010001; // 1261 :  81 - 0x51
      13'h4EE: dout <= 8'b01010001; // 1262 :  81 - 0x51
      13'h4EF: dout <= 8'b00000000; // 1263 :   0 - 0x0
      13'h4F0: dout <= 8'b11111111; // 1264 : 255 - 0xff -- Sprite 0x4f
      13'h4F1: dout <= 8'b11111111; // 1265 : 255 - 0xff
      13'h4F2: dout <= 8'b11110111; // 1266 : 247 - 0xf7
      13'h4F3: dout <= 8'b11111110; // 1267 : 254 - 0xfe
      13'h4F4: dout <= 8'b11111011; // 1268 : 251 - 0xfb
      13'h4F5: dout <= 8'b11111111; // 1269 : 255 - 0xff
      13'h4F6: dout <= 8'b11101111; // 1270 : 239 - 0xef
      13'h4F7: dout <= 8'b11111101; // 1271 : 253 - 0xfd
      13'h4F8: dout <= 8'b00000000; // 1272 :   0 - 0x0
      13'h4F9: dout <= 8'b00000000; // 1273 :   0 - 0x0
      13'h4FA: dout <= 8'b01001000; // 1274 :  72 - 0x48
      13'h4FB: dout <= 8'b01000001; // 1275 :  65 - 0x41
      13'h4FC: dout <= 8'b01000100; // 1276 :  68 - 0x44
      13'h4FD: dout <= 8'b01000000; // 1277 :  64 - 0x40
      13'h4FE: dout <= 8'b11010000; // 1278 : 208 - 0xd0
      13'h4FF: dout <= 8'b00000010; // 1279 :   2 - 0x2
      13'h500: dout <= 8'b11111111; // 1280 : 255 - 0xff -- Sprite 0x50
      13'h501: dout <= 8'b11111111; // 1281 : 255 - 0xff
      13'h502: dout <= 8'b00000011; // 1282 :   3 - 0x3
      13'h503: dout <= 8'b00000001; // 1283 :   1 - 0x1
      13'h504: dout <= 8'b11101110; // 1284 : 238 - 0xee
      13'h505: dout <= 8'b00000000; // 1285 :   0 - 0x0
      13'h506: dout <= 8'b11101110; // 1286 : 238 - 0xee
      13'h507: dout <= 8'b11101110; // 1287 : 238 - 0xee
      13'h508: dout <= 8'b00000000; // 1288 :   0 - 0x0
      13'h509: dout <= 8'b00000000; // 1289 :   0 - 0x0
      13'h50A: dout <= 8'b11111100; // 1290 : 252 - 0xfc
      13'h50B: dout <= 8'b11111110; // 1291 : 254 - 0xfe
      13'h50C: dout <= 8'b11101110; // 1292 : 238 - 0xee
      13'h50D: dout <= 8'b11101110; // 1293 : 238 - 0xee
      13'h50E: dout <= 8'b11101110; // 1294 : 238 - 0xee
      13'h50F: dout <= 8'b11101110; // 1295 : 238 - 0xee
      13'h510: dout <= 8'b11111111; // 1296 : 255 - 0xff -- Sprite 0x51
      13'h511: dout <= 8'b11111111; // 1297 : 255 - 0xff
      13'h512: dout <= 8'b00000011; // 1298 :   3 - 0x3
      13'h513: dout <= 8'b00000001; // 1299 :   1 - 0x1
      13'h514: dout <= 8'b11101110; // 1300 : 238 - 0xee
      13'h515: dout <= 8'b00000000; // 1301 :   0 - 0x0
      13'h516: dout <= 8'b11101110; // 1302 : 238 - 0xee
      13'h517: dout <= 8'b11101110; // 1303 : 238 - 0xee
      13'h518: dout <= 8'b00000000; // 1304 :   0 - 0x0
      13'h519: dout <= 8'b00000000; // 1305 :   0 - 0x0
      13'h51A: dout <= 8'b11111100; // 1306 : 252 - 0xfc
      13'h51B: dout <= 8'b11111110; // 1307 : 254 - 0xfe
      13'h51C: dout <= 8'b11101110; // 1308 : 238 - 0xee
      13'h51D: dout <= 8'b11101110; // 1309 : 238 - 0xee
      13'h51E: dout <= 8'b11101110; // 1310 : 238 - 0xee
      13'h51F: dout <= 8'b11101110; // 1311 : 238 - 0xee
      13'h520: dout <= 8'b11111111; // 1312 : 255 - 0xff -- Sprite 0x52
      13'h521: dout <= 8'b11111111; // 1313 : 255 - 0xff
      13'h522: dout <= 8'b00000001; // 1314 :   1 - 0x1
      13'h523: dout <= 8'b00000000; // 1315 :   0 - 0x0
      13'h524: dout <= 8'b11100000; // 1316 : 224 - 0xe0
      13'h525: dout <= 8'b00001111; // 1317 :  15 - 0xf
      13'h526: dout <= 8'b11111111; // 1318 : 255 - 0xff
      13'h527: dout <= 8'b11111011; // 1319 : 251 - 0xfb
      13'h528: dout <= 8'b00000000; // 1320 :   0 - 0x0
      13'h529: dout <= 8'b00000000; // 1321 :   0 - 0x0
      13'h52A: dout <= 8'b11111110; // 1322 : 254 - 0xfe
      13'h52B: dout <= 8'b11111110; // 1323 : 254 - 0xfe
      13'h52C: dout <= 8'b11100000; // 1324 : 224 - 0xe0
      13'h52D: dout <= 8'b11100000; // 1325 : 224 - 0xe0
      13'h52E: dout <= 8'b11111000; // 1326 : 248 - 0xf8
      13'h52F: dout <= 8'b11111000; // 1327 : 248 - 0xf8
      13'h530: dout <= 8'b11111111; // 1328 : 255 - 0xff -- Sprite 0x53
      13'h531: dout <= 8'b11111111; // 1329 : 255 - 0xff
      13'h532: dout <= 8'b10000011; // 1330 : 131 - 0x83
      13'h533: dout <= 8'b00000001; // 1331 :   1 - 0x1
      13'h534: dout <= 8'b11101110; // 1332 : 238 - 0xee
      13'h535: dout <= 8'b00000000; // 1333 :   0 - 0x0
      13'h536: dout <= 8'b11111111; // 1334 : 255 - 0xff
      13'h537: dout <= 8'b11111111; // 1335 : 255 - 0xff
      13'h538: dout <= 8'b00000000; // 1336 :   0 - 0x0
      13'h539: dout <= 8'b00000000; // 1337 :   0 - 0x0
      13'h53A: dout <= 8'b01111100; // 1338 : 124 - 0x7c
      13'h53B: dout <= 8'b11111110; // 1339 : 254 - 0xfe
      13'h53C: dout <= 8'b11101110; // 1340 : 238 - 0xee
      13'h53D: dout <= 8'b11100000; // 1341 : 224 - 0xe0
      13'h53E: dout <= 8'b11111100; // 1342 : 252 - 0xfc
      13'h53F: dout <= 8'b01111110; // 1343 : 126 - 0x7e
      13'h540: dout <= 8'b11111111; // 1344 : 255 - 0xff -- Sprite 0x54
      13'h541: dout <= 8'b11111111; // 1345 : 255 - 0xff
      13'h542: dout <= 8'b00000001; // 1346 :   1 - 0x1
      13'h543: dout <= 8'b00000000; // 1347 :   0 - 0x0
      13'h544: dout <= 8'b10111000; // 1348 : 184 - 0xb8
      13'h545: dout <= 8'b11000011; // 1349 : 195 - 0xc3
      13'h546: dout <= 8'b11111011; // 1350 : 251 - 0xfb
      13'h547: dout <= 8'b11111011; // 1351 : 251 - 0xfb
      13'h548: dout <= 8'b00000000; // 1352 :   0 - 0x0
      13'h549: dout <= 8'b00000000; // 1353 :   0 - 0x0
      13'h54A: dout <= 8'b11111110; // 1354 : 254 - 0xfe
      13'h54B: dout <= 8'b11111110; // 1355 : 254 - 0xfe
      13'h54C: dout <= 8'b00111000; // 1356 :  56 - 0x38
      13'h54D: dout <= 8'b00111000; // 1357 :  56 - 0x38
      13'h54E: dout <= 8'b00111000; // 1358 :  56 - 0x38
      13'h54F: dout <= 8'b00111000; // 1359 :  56 - 0x38
      13'h550: dout <= 8'b11111111; // 1360 : 255 - 0xff -- Sprite 0x55
      13'h551: dout <= 8'b11111111; // 1361 : 255 - 0xff
      13'h552: dout <= 8'b10000011; // 1362 : 131 - 0x83
      13'h553: dout <= 8'b00000001; // 1363 :   1 - 0x1
      13'h554: dout <= 8'b11101110; // 1364 : 238 - 0xee
      13'h555: dout <= 8'b00000000; // 1365 :   0 - 0x0
      13'h556: dout <= 8'b11101110; // 1366 : 238 - 0xee
      13'h557: dout <= 8'b11101110; // 1367 : 238 - 0xee
      13'h558: dout <= 8'b00000000; // 1368 :   0 - 0x0
      13'h559: dout <= 8'b00000000; // 1369 :   0 - 0x0
      13'h55A: dout <= 8'b01111100; // 1370 : 124 - 0x7c
      13'h55B: dout <= 8'b11111110; // 1371 : 254 - 0xfe
      13'h55C: dout <= 8'b11101110; // 1372 : 238 - 0xee
      13'h55D: dout <= 8'b11101110; // 1373 : 238 - 0xee
      13'h55E: dout <= 8'b11101110; // 1374 : 238 - 0xee
      13'h55F: dout <= 8'b11101110; // 1375 : 238 - 0xee
      13'h560: dout <= 8'b11111111; // 1376 : 255 - 0xff -- Sprite 0x56
      13'h561: dout <= 8'b11111111; // 1377 : 255 - 0xff
      13'h562: dout <= 8'b00011111; // 1378 :  31 - 0x1f
      13'h563: dout <= 8'b00001111; // 1379 :  15 - 0xf
      13'h564: dout <= 8'b11101111; // 1380 : 239 - 0xef
      13'h565: dout <= 8'b00001111; // 1381 :  15 - 0xf
      13'h566: dout <= 8'b11101111; // 1382 : 239 - 0xef
      13'h567: dout <= 8'b11101111; // 1383 : 239 - 0xef
      13'h568: dout <= 8'b00000000; // 1384 :   0 - 0x0
      13'h569: dout <= 8'b00000000; // 1385 :   0 - 0x0
      13'h56A: dout <= 8'b11100000; // 1386 : 224 - 0xe0
      13'h56B: dout <= 8'b11100000; // 1387 : 224 - 0xe0
      13'h56C: dout <= 8'b11100000; // 1388 : 224 - 0xe0
      13'h56D: dout <= 8'b11100000; // 1389 : 224 - 0xe0
      13'h56E: dout <= 8'b11100000; // 1390 : 224 - 0xe0
      13'h56F: dout <= 8'b11100000; // 1391 : 224 - 0xe0
      13'h570: dout <= 8'b11111111; // 1392 : 255 - 0xff -- Sprite 0x57
      13'h571: dout <= 8'b11111111; // 1393 : 255 - 0xff
      13'h572: dout <= 8'b00010001; // 1394 :  17 - 0x11
      13'h573: dout <= 8'b00000000; // 1395 :   0 - 0x0
      13'h574: dout <= 8'b11101110; // 1396 : 238 - 0xee
      13'h575: dout <= 8'b00000000; // 1397 :   0 - 0x0
      13'h576: dout <= 8'b11101110; // 1398 : 238 - 0xee
      13'h577: dout <= 8'b11101110; // 1399 : 238 - 0xee
      13'h578: dout <= 8'b00000000; // 1400 :   0 - 0x0
      13'h579: dout <= 8'b00000000; // 1401 :   0 - 0x0
      13'h57A: dout <= 8'b11101110; // 1402 : 238 - 0xee
      13'h57B: dout <= 8'b11101110; // 1403 : 238 - 0xee
      13'h57C: dout <= 8'b11101110; // 1404 : 238 - 0xee
      13'h57D: dout <= 8'b11101110; // 1405 : 238 - 0xee
      13'h57E: dout <= 8'b11101110; // 1406 : 238 - 0xee
      13'h57F: dout <= 8'b11101110; // 1407 : 238 - 0xee
      13'h580: dout <= 8'b11111111; // 1408 : 255 - 0xff -- Sprite 0x58
      13'h581: dout <= 8'b11111111; // 1409 : 255 - 0xff
      13'h582: dout <= 8'b01110001; // 1410 : 113 - 0x71
      13'h583: dout <= 8'b00110000; // 1411 :  48 - 0x30
      13'h584: dout <= 8'b11111110; // 1412 : 254 - 0xfe
      13'h585: dout <= 8'b00000000; // 1413 :   0 - 0x0
      13'h586: dout <= 8'b11111110; // 1414 : 254 - 0xfe
      13'h587: dout <= 8'b11101110; // 1415 : 238 - 0xee
      13'h588: dout <= 8'b00000000; // 1416 :   0 - 0x0
      13'h589: dout <= 8'b00000000; // 1417 :   0 - 0x0
      13'h58A: dout <= 8'b10001110; // 1418 : 142 - 0x8e
      13'h58B: dout <= 8'b11001110; // 1419 : 206 - 0xce
      13'h58C: dout <= 8'b11101110; // 1420 : 238 - 0xee
      13'h58D: dout <= 8'b11111110; // 1421 : 254 - 0xfe
      13'h58E: dout <= 8'b11111110; // 1422 : 254 - 0xfe
      13'h58F: dout <= 8'b11101110; // 1423 : 238 - 0xee
      13'h590: dout <= 8'b11111111; // 1424 : 255 - 0xff -- Sprite 0x59
      13'h591: dout <= 8'b11111111; // 1425 : 255 - 0xff
      13'h592: dout <= 8'b00000011; // 1426 :   3 - 0x3
      13'h593: dout <= 8'b00000001; // 1427 :   1 - 0x1
      13'h594: dout <= 8'b11101110; // 1428 : 238 - 0xee
      13'h595: dout <= 8'b00000000; // 1429 :   0 - 0x0
      13'h596: dout <= 8'b11101110; // 1430 : 238 - 0xee
      13'h597: dout <= 8'b11101110; // 1431 : 238 - 0xee
      13'h598: dout <= 8'b00000000; // 1432 :   0 - 0x0
      13'h599: dout <= 8'b00000000; // 1433 :   0 - 0x0
      13'h59A: dout <= 8'b11111100; // 1434 : 252 - 0xfc
      13'h59B: dout <= 8'b11111110; // 1435 : 254 - 0xfe
      13'h59C: dout <= 8'b11101110; // 1436 : 238 - 0xee
      13'h59D: dout <= 8'b11101110; // 1437 : 238 - 0xee
      13'h59E: dout <= 8'b11101110; // 1438 : 238 - 0xee
      13'h59F: dout <= 8'b11101110; // 1439 : 238 - 0xee
      13'h5A0: dout <= 8'b11111111; // 1440 : 255 - 0xff -- Sprite 0x5a
      13'h5A1: dout <= 8'b11111111; // 1441 : 255 - 0xff
      13'h5A2: dout <= 8'b10000011; // 1442 : 131 - 0x83
      13'h5A3: dout <= 8'b00000001; // 1443 :   1 - 0x1
      13'h5A4: dout <= 8'b11101110; // 1444 : 238 - 0xee
      13'h5A5: dout <= 8'b00000000; // 1445 :   0 - 0x0
      13'h5A6: dout <= 8'b11101110; // 1446 : 238 - 0xee
      13'h5A7: dout <= 8'b11101110; // 1447 : 238 - 0xee
      13'h5A8: dout <= 8'b00000000; // 1448 :   0 - 0x0
      13'h5A9: dout <= 8'b00000000; // 1449 :   0 - 0x0
      13'h5AA: dout <= 8'b01111100; // 1450 : 124 - 0x7c
      13'h5AB: dout <= 8'b11111110; // 1451 : 254 - 0xfe
      13'h5AC: dout <= 8'b11101110; // 1452 : 238 - 0xee
      13'h5AD: dout <= 8'b11101110; // 1453 : 238 - 0xee
      13'h5AE: dout <= 8'b11101110; // 1454 : 238 - 0xee
      13'h5AF: dout <= 8'b11101110; // 1455 : 238 - 0xee
      13'h5B0: dout <= 8'b11111111; // 1456 : 255 - 0xff -- Sprite 0x5b
      13'h5B1: dout <= 8'b11111111; // 1457 : 255 - 0xff
      13'h5B2: dout <= 8'b00000001; // 1458 :   1 - 0x1
      13'h5B3: dout <= 8'b00000000; // 1459 :   0 - 0x0
      13'h5B4: dout <= 8'b11100000; // 1460 : 224 - 0xe0
      13'h5B5: dout <= 8'b00001111; // 1461 :  15 - 0xf
      13'h5B6: dout <= 8'b11111111; // 1462 : 255 - 0xff
      13'h5B7: dout <= 8'b11111011; // 1463 : 251 - 0xfb
      13'h5B8: dout <= 8'b00000000; // 1464 :   0 - 0x0
      13'h5B9: dout <= 8'b00000000; // 1465 :   0 - 0x0
      13'h5BA: dout <= 8'b11111110; // 1466 : 254 - 0xfe
      13'h5BB: dout <= 8'b11111110; // 1467 : 254 - 0xfe
      13'h5BC: dout <= 8'b11100000; // 1468 : 224 - 0xe0
      13'h5BD: dout <= 8'b11100000; // 1469 : 224 - 0xe0
      13'h5BE: dout <= 8'b11111000; // 1470 : 248 - 0xf8
      13'h5BF: dout <= 8'b11111000; // 1471 : 248 - 0xf8
      13'h5C0: dout <= 8'b11111111; // 1472 : 255 - 0xff -- Sprite 0x5c
      13'h5C1: dout <= 8'b11111111; // 1473 : 255 - 0xff
      13'h5C2: dout <= 8'b11111111; // 1474 : 255 - 0xff
      13'h5C3: dout <= 8'b11111111; // 1475 : 255 - 0xff
      13'h5C4: dout <= 8'b11111111; // 1476 : 255 - 0xff
      13'h5C5: dout <= 8'b11111111; // 1477 : 255 - 0xff
      13'h5C6: dout <= 8'b11111111; // 1478 : 255 - 0xff
      13'h5C7: dout <= 8'b11011101; // 1479 : 221 - 0xdd
      13'h5C8: dout <= 8'b00000000; // 1480 :   0 - 0x0
      13'h5C9: dout <= 8'b00000000; // 1481 :   0 - 0x0
      13'h5CA: dout <= 8'b00000000; // 1482 :   0 - 0x0
      13'h5CB: dout <= 8'b00000000; // 1483 :   0 - 0x0
      13'h5CC: dout <= 8'b00000000; // 1484 :   0 - 0x0
      13'h5CD: dout <= 8'b00000000; // 1485 :   0 - 0x0
      13'h5CE: dout <= 8'b11001100; // 1486 : 204 - 0xcc
      13'h5CF: dout <= 8'b11001100; // 1487 : 204 - 0xcc
      13'h5D0: dout <= 8'b11111111; // 1488 : 255 - 0xff -- Sprite 0x5d
      13'h5D1: dout <= 8'b11111111; // 1489 : 255 - 0xff
      13'h5D2: dout <= 8'b00000001; // 1490 :   1 - 0x1
      13'h5D3: dout <= 8'b00000000; // 1491 :   0 - 0x0
      13'h5D4: dout <= 8'b11100000; // 1492 : 224 - 0xe0
      13'h5D5: dout <= 8'b00001111; // 1493 :  15 - 0xf
      13'h5D6: dout <= 8'b11111111; // 1494 : 255 - 0xff
      13'h5D7: dout <= 8'b11111011; // 1495 : 251 - 0xfb
      13'h5D8: dout <= 8'b00000000; // 1496 :   0 - 0x0
      13'h5D9: dout <= 8'b00000000; // 1497 :   0 - 0x0
      13'h5DA: dout <= 8'b11111110; // 1498 : 254 - 0xfe
      13'h5DB: dout <= 8'b11111110; // 1499 : 254 - 0xfe
      13'h5DC: dout <= 8'b11100000; // 1500 : 224 - 0xe0
      13'h5DD: dout <= 8'b11100000; // 1501 : 224 - 0xe0
      13'h5DE: dout <= 8'b11111000; // 1502 : 248 - 0xf8
      13'h5DF: dout <= 8'b11111000; // 1503 : 248 - 0xf8
      13'h5E0: dout <= 8'b11111111; // 1504 : 255 - 0xff -- Sprite 0x5e
      13'h5E1: dout <= 8'b11111111; // 1505 : 255 - 0xff
      13'h5E2: dout <= 8'b00010001; // 1506 :  17 - 0x11
      13'h5E3: dout <= 8'b00000000; // 1507 :   0 - 0x0
      13'h5E4: dout <= 8'b11101110; // 1508 : 238 - 0xee
      13'h5E5: dout <= 8'b00000000; // 1509 :   0 - 0x0
      13'h5E6: dout <= 8'b11101110; // 1510 : 238 - 0xee
      13'h5E7: dout <= 8'b11101110; // 1511 : 238 - 0xee
      13'h5E8: dout <= 8'b00000000; // 1512 :   0 - 0x0
      13'h5E9: dout <= 8'b00000000; // 1513 :   0 - 0x0
      13'h5EA: dout <= 8'b11101110; // 1514 : 238 - 0xee
      13'h5EB: dout <= 8'b11101110; // 1515 : 238 - 0xee
      13'h5EC: dout <= 8'b11101110; // 1516 : 238 - 0xee
      13'h5ED: dout <= 8'b11101110; // 1517 : 238 - 0xee
      13'h5EE: dout <= 8'b11101110; // 1518 : 238 - 0xee
      13'h5EF: dout <= 8'b11101110; // 1519 : 238 - 0xee
      13'h5F0: dout <= 8'b10111101; // 1520 : 189 - 0xbd -- Sprite 0x5f
      13'h5F1: dout <= 8'b11111111; // 1521 : 255 - 0xff
      13'h5F2: dout <= 8'b11111111; // 1522 : 255 - 0xff
      13'h5F3: dout <= 8'b11111111; // 1523 : 255 - 0xff
      13'h5F4: dout <= 8'b11111111; // 1524 : 255 - 0xff
      13'h5F5: dout <= 8'b11111111; // 1525 : 255 - 0xff
      13'h5F6: dout <= 8'b11111111; // 1526 : 255 - 0xff
      13'h5F7: dout <= 8'b11111111; // 1527 : 255 - 0xff
      13'h5F8: dout <= 8'b01111110; // 1528 : 126 - 0x7e
      13'h5F9: dout <= 8'b01111110; // 1529 : 126 - 0x7e
      13'h5FA: dout <= 8'b01111110; // 1530 : 126 - 0x7e
      13'h5FB: dout <= 8'b01111110; // 1531 : 126 - 0x7e
      13'h5FC: dout <= 8'b01111110; // 1532 : 126 - 0x7e
      13'h5FD: dout <= 8'b01111110; // 1533 : 126 - 0x7e
      13'h5FE: dout <= 8'b01111110; // 1534 : 126 - 0x7e
      13'h5FF: dout <= 8'b01111110; // 1535 : 126 - 0x7e
      13'h600: dout <= 8'b11101110; // 1536 : 238 - 0xee -- Sprite 0x60
      13'h601: dout <= 8'b00000000; // 1537 :   0 - 0x0
      13'h602: dout <= 8'b11111110; // 1538 : 254 - 0xfe
      13'h603: dout <= 8'b00000000; // 1539 :   0 - 0x0
      13'h604: dout <= 8'b00000001; // 1540 :   1 - 0x1
      13'h605: dout <= 8'b00001111; // 1541 :  15 - 0xf
      13'h606: dout <= 8'b10001111; // 1542 : 143 - 0x8f
      13'h607: dout <= 8'b11111111; // 1543 : 255 - 0xff
      13'h608: dout <= 8'b11101110; // 1544 : 238 - 0xee
      13'h609: dout <= 8'b11101110; // 1545 : 238 - 0xee
      13'h60A: dout <= 8'b11111110; // 1546 : 254 - 0xfe
      13'h60B: dout <= 8'b11111100; // 1547 : 252 - 0xfc
      13'h60C: dout <= 8'b11100000; // 1548 : 224 - 0xe0
      13'h60D: dout <= 8'b11100000; // 1549 : 224 - 0xe0
      13'h60E: dout <= 8'b00000000; // 1550 :   0 - 0x0
      13'h60F: dout <= 8'b00000000; // 1551 :   0 - 0x0
      13'h610: dout <= 8'b11101110; // 1552 : 238 - 0xee -- Sprite 0x61
      13'h611: dout <= 8'b00000000; // 1553 :   0 - 0x0
      13'h612: dout <= 8'b11111100; // 1554 : 252 - 0xfc
      13'h613: dout <= 8'b00000001; // 1555 :   1 - 0x1
      13'h614: dout <= 8'b00000001; // 1556 :   1 - 0x1
      13'h615: dout <= 8'b00000000; // 1557 :   0 - 0x0
      13'h616: dout <= 8'b10001000; // 1558 : 136 - 0x88
      13'h617: dout <= 8'b11111111; // 1559 : 255 - 0xff
      13'h618: dout <= 8'b11101110; // 1560 : 238 - 0xee
      13'h619: dout <= 8'b11101110; // 1561 : 238 - 0xee
      13'h61A: dout <= 8'b11111100; // 1562 : 252 - 0xfc
      13'h61B: dout <= 8'b11111100; // 1563 : 252 - 0xfc
      13'h61C: dout <= 8'b11101110; // 1564 : 238 - 0xee
      13'h61D: dout <= 8'b11101110; // 1565 : 238 - 0xee
      13'h61E: dout <= 8'b00000000; // 1566 :   0 - 0x0
      13'h61F: dout <= 8'b00000000; // 1567 :   0 - 0x0
      13'h620: dout <= 8'b11100011; // 1568 : 227 - 0xe3 -- Sprite 0x62
      13'h621: dout <= 8'b00001111; // 1569 :  15 - 0xf
      13'h622: dout <= 8'b11101111; // 1570 : 239 - 0xef
      13'h623: dout <= 8'b00001111; // 1571 :  15 - 0xf
      13'h624: dout <= 8'b00000001; // 1572 :   1 - 0x1
      13'h625: dout <= 8'b00000000; // 1573 :   0 - 0x0
      13'h626: dout <= 8'b10000000; // 1574 : 128 - 0x80
      13'h627: dout <= 8'b11111111; // 1575 : 255 - 0xff
      13'h628: dout <= 8'b11100000; // 1576 : 224 - 0xe0
      13'h629: dout <= 8'b11100000; // 1577 : 224 - 0xe0
      13'h62A: dout <= 8'b11100000; // 1578 : 224 - 0xe0
      13'h62B: dout <= 8'b11100000; // 1579 : 224 - 0xe0
      13'h62C: dout <= 8'b11111110; // 1580 : 254 - 0xfe
      13'h62D: dout <= 8'b11111110; // 1581 : 254 - 0xfe
      13'h62E: dout <= 8'b00000000; // 1582 :   0 - 0x0
      13'h62F: dout <= 8'b00000000; // 1583 :   0 - 0x0
      13'h630: dout <= 8'b11001110; // 1584 : 206 - 0xce -- Sprite 0x63
      13'h631: dout <= 8'b11110000; // 1585 : 240 - 0xf0
      13'h632: dout <= 8'b11111110; // 1586 : 254 - 0xfe
      13'h633: dout <= 8'b00010000; // 1587 :  16 - 0x10
      13'h634: dout <= 8'b00000000; // 1588 :   0 - 0x0
      13'h635: dout <= 8'b10000000; // 1589 : 128 - 0x80
      13'h636: dout <= 8'b11000001; // 1590 : 193 - 0xc1
      13'h637: dout <= 8'b11111111; // 1591 : 255 - 0xff
      13'h638: dout <= 8'b00001110; // 1592 :  14 - 0xe
      13'h639: dout <= 8'b00001110; // 1593 :  14 - 0xe
      13'h63A: dout <= 8'b00001110; // 1594 :  14 - 0xe
      13'h63B: dout <= 8'b11101110; // 1595 : 238 - 0xee
      13'h63C: dout <= 8'b11111110; // 1596 : 254 - 0xfe
      13'h63D: dout <= 8'b01111100; // 1597 : 124 - 0x7c
      13'h63E: dout <= 8'b00000000; // 1598 :   0 - 0x0
      13'h63F: dout <= 8'b00000000; // 1599 :   0 - 0x0
      13'h640: dout <= 8'b11111011; // 1600 : 251 - 0xfb -- Sprite 0x64
      13'h641: dout <= 8'b11000011; // 1601 : 195 - 0xc3
      13'h642: dout <= 8'b11111011; // 1602 : 251 - 0xfb
      13'h643: dout <= 8'b11000011; // 1603 : 195 - 0xc3
      13'h644: dout <= 8'b11000011; // 1604 : 195 - 0xc3
      13'h645: dout <= 8'b11000011; // 1605 : 195 - 0xc3
      13'h646: dout <= 8'b11100011; // 1606 : 227 - 0xe3
      13'h647: dout <= 8'b11111111; // 1607 : 255 - 0xff
      13'h648: dout <= 8'b00111000; // 1608 :  56 - 0x38
      13'h649: dout <= 8'b00111000; // 1609 :  56 - 0x38
      13'h64A: dout <= 8'b00111000; // 1610 :  56 - 0x38
      13'h64B: dout <= 8'b00111000; // 1611 :  56 - 0x38
      13'h64C: dout <= 8'b00111000; // 1612 :  56 - 0x38
      13'h64D: dout <= 8'b00111000; // 1613 :  56 - 0x38
      13'h64E: dout <= 8'b00000000; // 1614 :   0 - 0x0
      13'h64F: dout <= 8'b00000000; // 1615 :   0 - 0x0
      13'h650: dout <= 8'b11101110; // 1616 : 238 - 0xee -- Sprite 0x65
      13'h651: dout <= 8'b00000000; // 1617 :   0 - 0x0
      13'h652: dout <= 8'b11111110; // 1618 : 254 - 0xfe
      13'h653: dout <= 8'b00000000; // 1619 :   0 - 0x0
      13'h654: dout <= 8'b00000000; // 1620 :   0 - 0x0
      13'h655: dout <= 8'b00000000; // 1621 :   0 - 0x0
      13'h656: dout <= 8'b10001000; // 1622 : 136 - 0x88
      13'h657: dout <= 8'b11111111; // 1623 : 255 - 0xff
      13'h658: dout <= 8'b11101110; // 1624 : 238 - 0xee
      13'h659: dout <= 8'b11101110; // 1625 : 238 - 0xee
      13'h65A: dout <= 8'b11111110; // 1626 : 254 - 0xfe
      13'h65B: dout <= 8'b11111110; // 1627 : 254 - 0xfe
      13'h65C: dout <= 8'b11101110; // 1628 : 238 - 0xee
      13'h65D: dout <= 8'b11101110; // 1629 : 238 - 0xee
      13'h65E: dout <= 8'b00000000; // 1630 :   0 - 0x0
      13'h65F: dout <= 8'b00000000; // 1631 :   0 - 0x0
      13'h660: dout <= 8'b11101111; // 1632 : 239 - 0xef -- Sprite 0x66
      13'h661: dout <= 8'b00001111; // 1633 :  15 - 0xf
      13'h662: dout <= 8'b11101111; // 1634 : 239 - 0xef
      13'h663: dout <= 8'b00000001; // 1635 :   1 - 0x1
      13'h664: dout <= 8'b00000000; // 1636 :   0 - 0x0
      13'h665: dout <= 8'b00000000; // 1637 :   0 - 0x0
      13'h666: dout <= 8'b10000000; // 1638 : 128 - 0x80
      13'h667: dout <= 8'b11111111; // 1639 : 255 - 0xff
      13'h668: dout <= 8'b11100000; // 1640 : 224 - 0xe0
      13'h669: dout <= 8'b11100000; // 1641 : 224 - 0xe0
      13'h66A: dout <= 8'b11100000; // 1642 : 224 - 0xe0
      13'h66B: dout <= 8'b11101110; // 1643 : 238 - 0xee
      13'h66C: dout <= 8'b11111110; // 1644 : 254 - 0xfe
      13'h66D: dout <= 8'b11111110; // 1645 : 254 - 0xfe
      13'h66E: dout <= 8'b00000000; // 1646 :   0 - 0x0
      13'h66F: dout <= 8'b00000000; // 1647 :   0 - 0x0
      13'h670: dout <= 8'b11101110; // 1648 : 238 - 0xee -- Sprite 0x67
      13'h671: dout <= 8'b00000000; // 1649 :   0 - 0x0
      13'h672: dout <= 8'b11111110; // 1650 : 254 - 0xfe
      13'h673: dout <= 8'b00000000; // 1651 :   0 - 0x0
      13'h674: dout <= 8'b00000000; // 1652 :   0 - 0x0
      13'h675: dout <= 8'b00001000; // 1653 :   8 - 0x8
      13'h676: dout <= 8'b10011100; // 1654 : 156 - 0x9c
      13'h677: dout <= 8'b11111111; // 1655 : 255 - 0xff
      13'h678: dout <= 8'b11101110; // 1656 : 238 - 0xee
      13'h679: dout <= 8'b11101110; // 1657 : 238 - 0xee
      13'h67A: dout <= 8'b11111110; // 1658 : 254 - 0xfe
      13'h67B: dout <= 8'b11111110; // 1659 : 254 - 0xfe
      13'h67C: dout <= 8'b11101110; // 1660 : 238 - 0xee
      13'h67D: dout <= 8'b11000110; // 1661 : 198 - 0xc6
      13'h67E: dout <= 8'b00000000; // 1662 :   0 - 0x0
      13'h67F: dout <= 8'b00000000; // 1663 :   0 - 0x0
      13'h680: dout <= 8'b11101110; // 1664 : 238 - 0xee -- Sprite 0x68
      13'h681: dout <= 8'b00000000; // 1665 :   0 - 0x0
      13'h682: dout <= 8'b11101110; // 1666 : 238 - 0xee
      13'h683: dout <= 8'b00000000; // 1667 :   0 - 0x0
      13'h684: dout <= 8'b00000000; // 1668 :   0 - 0x0
      13'h685: dout <= 8'b00000000; // 1669 :   0 - 0x0
      13'h686: dout <= 8'b10001000; // 1670 : 136 - 0x88
      13'h687: dout <= 8'b11111111; // 1671 : 255 - 0xff
      13'h688: dout <= 8'b11101110; // 1672 : 238 - 0xee
      13'h689: dout <= 8'b11101110; // 1673 : 238 - 0xee
      13'h68A: dout <= 8'b11101110; // 1674 : 238 - 0xee
      13'h68B: dout <= 8'b11101110; // 1675 : 238 - 0xee
      13'h68C: dout <= 8'b11101110; // 1676 : 238 - 0xee
      13'h68D: dout <= 8'b11101110; // 1677 : 238 - 0xee
      13'h68E: dout <= 8'b00000000; // 1678 :   0 - 0x0
      13'h68F: dout <= 8'b00000000; // 1679 :   0 - 0x0
      13'h690: dout <= 8'b11101110; // 1680 : 238 - 0xee -- Sprite 0x69
      13'h691: dout <= 8'b00000000; // 1681 :   0 - 0x0
      13'h692: dout <= 8'b11101110; // 1682 : 238 - 0xee
      13'h693: dout <= 8'b00000000; // 1683 :   0 - 0x0
      13'h694: dout <= 8'b00000000; // 1684 :   0 - 0x0
      13'h695: dout <= 8'b00000000; // 1685 :   0 - 0x0
      13'h696: dout <= 8'b10000001; // 1686 : 129 - 0x81
      13'h697: dout <= 8'b11111111; // 1687 : 255 - 0xff
      13'h698: dout <= 8'b11101110; // 1688 : 238 - 0xee
      13'h699: dout <= 8'b11101110; // 1689 : 238 - 0xee
      13'h69A: dout <= 8'b11101110; // 1690 : 238 - 0xee
      13'h69B: dout <= 8'b11101110; // 1691 : 238 - 0xee
      13'h69C: dout <= 8'b11111110; // 1692 : 254 - 0xfe
      13'h69D: dout <= 8'b11111100; // 1693 : 252 - 0xfc
      13'h69E: dout <= 8'b00000000; // 1694 :   0 - 0x0
      13'h69F: dout <= 8'b00000000; // 1695 :   0 - 0x0
      13'h6A0: dout <= 8'b11101110; // 1696 : 238 - 0xee -- Sprite 0x6a
      13'h6A1: dout <= 8'b00000000; // 1697 :   0 - 0x0
      13'h6A2: dout <= 8'b11101110; // 1698 : 238 - 0xee
      13'h6A3: dout <= 8'b00000000; // 1699 :   0 - 0x0
      13'h6A4: dout <= 8'b00000000; // 1700 :   0 - 0x0
      13'h6A5: dout <= 8'b10000000; // 1701 : 128 - 0x80
      13'h6A6: dout <= 8'b11000001; // 1702 : 193 - 0xc1
      13'h6A7: dout <= 8'b11111111; // 1703 : 255 - 0xff
      13'h6A8: dout <= 8'b11101110; // 1704 : 238 - 0xee
      13'h6A9: dout <= 8'b11101110; // 1705 : 238 - 0xee
      13'h6AA: dout <= 8'b11101110; // 1706 : 238 - 0xee
      13'h6AB: dout <= 8'b11101110; // 1707 : 238 - 0xee
      13'h6AC: dout <= 8'b11111110; // 1708 : 254 - 0xfe
      13'h6AD: dout <= 8'b01111100; // 1709 : 124 - 0x7c
      13'h6AE: dout <= 8'b00000000; // 1710 :   0 - 0x0
      13'h6AF: dout <= 8'b00000000; // 1711 :   0 - 0x0
      13'h6B0: dout <= 8'b11100011; // 1712 : 227 - 0xe3 -- Sprite 0x6b
      13'h6B1: dout <= 8'b00001111; // 1713 :  15 - 0xf
      13'h6B2: dout <= 8'b11101111; // 1714 : 239 - 0xef
      13'h6B3: dout <= 8'b00001111; // 1715 :  15 - 0xf
      13'h6B4: dout <= 8'b00000001; // 1716 :   1 - 0x1
      13'h6B5: dout <= 8'b00000000; // 1717 :   0 - 0x0
      13'h6B6: dout <= 8'b10000000; // 1718 : 128 - 0x80
      13'h6B7: dout <= 8'b11111111; // 1719 : 255 - 0xff
      13'h6B8: dout <= 8'b11100000; // 1720 : 224 - 0xe0
      13'h6B9: dout <= 8'b11100000; // 1721 : 224 - 0xe0
      13'h6BA: dout <= 8'b11100000; // 1722 : 224 - 0xe0
      13'h6BB: dout <= 8'b11100000; // 1723 : 224 - 0xe0
      13'h6BC: dout <= 8'b11111110; // 1724 : 254 - 0xfe
      13'h6BD: dout <= 8'b11111110; // 1725 : 254 - 0xfe
      13'h6BE: dout <= 8'b00000000; // 1726 :   0 - 0x0
      13'h6BF: dout <= 8'b00000000; // 1727 :   0 - 0x0
      13'h6C0: dout <= 8'b10011001; // 1728 : 153 - 0x99 -- Sprite 0x6c
      13'h6C1: dout <= 8'b11100011; // 1729 : 227 - 0xe3
      13'h6C2: dout <= 8'b11110011; // 1730 : 243 - 0xf3
      13'h6C3: dout <= 8'b11000111; // 1731 : 199 - 0xc7
      13'h6C4: dout <= 8'b10000001; // 1732 : 129 - 0x81
      13'h6C5: dout <= 8'b10001000; // 1733 : 136 - 0x88
      13'h6C6: dout <= 8'b11001100; // 1734 : 204 - 0xcc
      13'h6C7: dout <= 8'b11111111; // 1735 : 255 - 0xff
      13'h6C8: dout <= 8'b00011000; // 1736 :  24 - 0x18
      13'h6C9: dout <= 8'b00011000; // 1737 :  24 - 0x18
      13'h6CA: dout <= 8'b00110000; // 1738 :  48 - 0x30
      13'h6CB: dout <= 8'b00110000; // 1739 :  48 - 0x30
      13'h6CC: dout <= 8'b01100110; // 1740 : 102 - 0x66
      13'h6CD: dout <= 8'b01100110; // 1741 : 102 - 0x66
      13'h6CE: dout <= 8'b00000000; // 1742 :   0 - 0x0
      13'h6CF: dout <= 8'b00000000; // 1743 :   0 - 0x0
      13'h6D0: dout <= 8'b11100011; // 1744 : 227 - 0xe3 -- Sprite 0x6d
      13'h6D1: dout <= 8'b00001111; // 1745 :  15 - 0xf
      13'h6D2: dout <= 8'b11101111; // 1746 : 239 - 0xef
      13'h6D3: dout <= 8'b00001111; // 1747 :  15 - 0xf
      13'h6D4: dout <= 8'b00001111; // 1748 :  15 - 0xf
      13'h6D5: dout <= 8'b00001111; // 1749 :  15 - 0xf
      13'h6D6: dout <= 8'b10001111; // 1750 : 143 - 0x8f
      13'h6D7: dout <= 8'b11111111; // 1751 : 255 - 0xff
      13'h6D8: dout <= 8'b11100000; // 1752 : 224 - 0xe0
      13'h6D9: dout <= 8'b11100000; // 1753 : 224 - 0xe0
      13'h6DA: dout <= 8'b11100000; // 1754 : 224 - 0xe0
      13'h6DB: dout <= 8'b11100000; // 1755 : 224 - 0xe0
      13'h6DC: dout <= 8'b11100000; // 1756 : 224 - 0xe0
      13'h6DD: dout <= 8'b11100000; // 1757 : 224 - 0xe0
      13'h6DE: dout <= 8'b00000000; // 1758 :   0 - 0x0
      13'h6DF: dout <= 8'b00000000; // 1759 :   0 - 0x0
      13'h6E0: dout <= 8'b11101110; // 1760 : 238 - 0xee -- Sprite 0x6e
      13'h6E1: dout <= 8'b00000000; // 1761 :   0 - 0x0
      13'h6E2: dout <= 8'b11101110; // 1762 : 238 - 0xee
      13'h6E3: dout <= 8'b00000000; // 1763 :   0 - 0x0
      13'h6E4: dout <= 8'b00000000; // 1764 :   0 - 0x0
      13'h6E5: dout <= 8'b10000000; // 1765 : 128 - 0x80
      13'h6E6: dout <= 8'b11000001; // 1766 : 193 - 0xc1
      13'h6E7: dout <= 8'b11111111; // 1767 : 255 - 0xff
      13'h6E8: dout <= 8'b11101110; // 1768 : 238 - 0xee
      13'h6E9: dout <= 8'b11101110; // 1769 : 238 - 0xee
      13'h6EA: dout <= 8'b11101110; // 1770 : 238 - 0xee
      13'h6EB: dout <= 8'b11101110; // 1771 : 238 - 0xee
      13'h6EC: dout <= 8'b11111110; // 1772 : 254 - 0xfe
      13'h6ED: dout <= 8'b01111100; // 1773 : 124 - 0x7c
      13'h6EE: dout <= 8'b00000000; // 1774 :   0 - 0x0
      13'h6EF: dout <= 8'b00000000; // 1775 :   0 - 0x0
      13'h6F0: dout <= 8'b11111111; // 1776 : 255 - 0xff -- Sprite 0x6f
      13'h6F1: dout <= 8'b11111111; // 1777 : 255 - 0xff
      13'h6F2: dout <= 8'b11111111; // 1778 : 255 - 0xff
      13'h6F3: dout <= 8'b10111101; // 1779 : 189 - 0xbd
      13'h6F4: dout <= 8'b11111111; // 1780 : 255 - 0xff
      13'h6F5: dout <= 8'b11011011; // 1781 : 219 - 0xdb
      13'h6F6: dout <= 8'b11111111; // 1782 : 255 - 0xff
      13'h6F7: dout <= 8'b11111111; // 1783 : 255 - 0xff
      13'h6F8: dout <= 8'b01111110; // 1784 : 126 - 0x7e
      13'h6F9: dout <= 8'b01111110; // 1785 : 126 - 0x7e
      13'h6FA: dout <= 8'b01111110; // 1786 : 126 - 0x7e
      13'h6FB: dout <= 8'b01111110; // 1787 : 126 - 0x7e
      13'h6FC: dout <= 8'b00111100; // 1788 :  60 - 0x3c
      13'h6FD: dout <= 8'b00111100; // 1789 :  60 - 0x3c
      13'h6FE: dout <= 8'b00000000; // 1790 :   0 - 0x0
      13'h6FF: dout <= 8'b00000000; // 1791 :   0 - 0x0
      13'h700: dout <= 8'b11111011; // 1792 : 251 - 0xfb -- Sprite 0x70
      13'h701: dout <= 8'b11101111; // 1793 : 239 - 0xef
      13'h702: dout <= 8'b11011111; // 1794 : 223 - 0xdf
      13'h703: dout <= 8'b11111111; // 1795 : 255 - 0xff
      13'h704: dout <= 8'b10111111; // 1796 : 191 - 0xbf
      13'h705: dout <= 8'b10111111; // 1797 : 191 - 0xbf
      13'h706: dout <= 8'b11111110; // 1798 : 254 - 0xfe
      13'h707: dout <= 8'b11111111; // 1799 : 255 - 0xff
      13'h708: dout <= 8'b00000111; // 1800 :   7 - 0x7
      13'h709: dout <= 8'b00011111; // 1801 :  31 - 0x1f
      13'h70A: dout <= 8'b00111111; // 1802 :  63 - 0x3f
      13'h70B: dout <= 8'b00111111; // 1803 :  63 - 0x3f
      13'h70C: dout <= 8'b01111111; // 1804 : 127 - 0x7f
      13'h70D: dout <= 8'b01111111; // 1805 : 127 - 0x7f
      13'h70E: dout <= 8'b01111111; // 1806 : 127 - 0x7f
      13'h70F: dout <= 8'b01111110; // 1807 : 126 - 0x7e
      13'h710: dout <= 8'b11011111; // 1808 : 223 - 0xdf -- Sprite 0x71
      13'h711: dout <= 8'b11110111; // 1809 : 247 - 0xf7
      13'h712: dout <= 8'b11111011; // 1810 : 251 - 0xfb
      13'h713: dout <= 8'b11111111; // 1811 : 255 - 0xff
      13'h714: dout <= 8'b11111101; // 1812 : 253 - 0xfd
      13'h715: dout <= 8'b11111101; // 1813 : 253 - 0xfd
      13'h716: dout <= 8'b01111111; // 1814 : 127 - 0x7f
      13'h717: dout <= 8'b11111111; // 1815 : 255 - 0xff
      13'h718: dout <= 8'b11100000; // 1816 : 224 - 0xe0
      13'h719: dout <= 8'b11111000; // 1817 : 248 - 0xf8
      13'h71A: dout <= 8'b11111100; // 1818 : 252 - 0xfc
      13'h71B: dout <= 8'b11111100; // 1819 : 252 - 0xfc
      13'h71C: dout <= 8'b11111110; // 1820 : 254 - 0xfe
      13'h71D: dout <= 8'b11111110; // 1821 : 254 - 0xfe
      13'h71E: dout <= 8'b11111110; // 1822 : 254 - 0xfe
      13'h71F: dout <= 8'b01111110; // 1823 : 126 - 0x7e
      13'h720: dout <= 8'b11111111; // 1824 : 255 - 0xff -- Sprite 0x72
      13'h721: dout <= 8'b11111111; // 1825 : 255 - 0xff
      13'h722: dout <= 8'b11111111; // 1826 : 255 - 0xff
      13'h723: dout <= 8'b11111111; // 1827 : 255 - 0xff
      13'h724: dout <= 8'b11111111; // 1828 : 255 - 0xff
      13'h725: dout <= 8'b11111111; // 1829 : 255 - 0xff
      13'h726: dout <= 8'b11111111; // 1830 : 255 - 0xff
      13'h727: dout <= 8'b11111111; // 1831 : 255 - 0xff
      13'h728: dout <= 8'b01111110; // 1832 : 126 - 0x7e
      13'h729: dout <= 8'b01111110; // 1833 : 126 - 0x7e
      13'h72A: dout <= 8'b01111110; // 1834 : 126 - 0x7e
      13'h72B: dout <= 8'b01111110; // 1835 : 126 - 0x7e
      13'h72C: dout <= 8'b01111110; // 1836 : 126 - 0x7e
      13'h72D: dout <= 8'b01111110; // 1837 : 126 - 0x7e
      13'h72E: dout <= 8'b01111110; // 1838 : 126 - 0x7e
      13'h72F: dout <= 8'b01111110; // 1839 : 126 - 0x7e
      13'h730: dout <= 8'b11111111; // 1840 : 255 - 0xff -- Sprite 0x73
      13'h731: dout <= 8'b11111110; // 1841 : 254 - 0xfe
      13'h732: dout <= 8'b10111111; // 1842 : 191 - 0xbf
      13'h733: dout <= 8'b10111111; // 1843 : 191 - 0xbf
      13'h734: dout <= 8'b11111111; // 1844 : 255 - 0xff
      13'h735: dout <= 8'b11011111; // 1845 : 223 - 0xdf
      13'h736: dout <= 8'b11101111; // 1846 : 239 - 0xef
      13'h737: dout <= 8'b11111011; // 1847 : 251 - 0xfb
      13'h738: dout <= 8'b01111110; // 1848 : 126 - 0x7e
      13'h739: dout <= 8'b01111111; // 1849 : 127 - 0x7f
      13'h73A: dout <= 8'b01111111; // 1850 : 127 - 0x7f
      13'h73B: dout <= 8'b01111111; // 1851 : 127 - 0x7f
      13'h73C: dout <= 8'b00111111; // 1852 :  63 - 0x3f
      13'h73D: dout <= 8'b00111111; // 1853 :  63 - 0x3f
      13'h73E: dout <= 8'b00011111; // 1854 :  31 - 0x1f
      13'h73F: dout <= 8'b00000111; // 1855 :   7 - 0x7
      13'h740: dout <= 8'b11111111; // 1856 : 255 - 0xff -- Sprite 0x74
      13'h741: dout <= 8'b01111111; // 1857 : 127 - 0x7f
      13'h742: dout <= 8'b11111101; // 1858 : 253 - 0xfd
      13'h743: dout <= 8'b11111101; // 1859 : 253 - 0xfd
      13'h744: dout <= 8'b11111111; // 1860 : 255 - 0xff
      13'h745: dout <= 8'b11111011; // 1861 : 251 - 0xfb
      13'h746: dout <= 8'b11110111; // 1862 : 247 - 0xf7
      13'h747: dout <= 8'b11011111; // 1863 : 223 - 0xdf
      13'h748: dout <= 8'b01111110; // 1864 : 126 - 0x7e
      13'h749: dout <= 8'b11111110; // 1865 : 254 - 0xfe
      13'h74A: dout <= 8'b11111110; // 1866 : 254 - 0xfe
      13'h74B: dout <= 8'b11111110; // 1867 : 254 - 0xfe
      13'h74C: dout <= 8'b11111100; // 1868 : 252 - 0xfc
      13'h74D: dout <= 8'b11111100; // 1869 : 252 - 0xfc
      13'h74E: dout <= 8'b11111000; // 1870 : 248 - 0xf8
      13'h74F: dout <= 8'b11100000; // 1871 : 224 - 0xe0
      13'h750: dout <= 8'b11111111; // 1872 : 255 - 0xff -- Sprite 0x75
      13'h751: dout <= 8'b11111111; // 1873 : 255 - 0xff
      13'h752: dout <= 8'b11111111; // 1874 : 255 - 0xff
      13'h753: dout <= 8'b11111111; // 1875 : 255 - 0xff
      13'h754: dout <= 8'b11111111; // 1876 : 255 - 0xff
      13'h755: dout <= 8'b11111111; // 1877 : 255 - 0xff
      13'h756: dout <= 8'b11111111; // 1878 : 255 - 0xff
      13'h757: dout <= 8'b11111111; // 1879 : 255 - 0xff
      13'h758: dout <= 8'b01111111; // 1880 : 127 - 0x7f
      13'h759: dout <= 8'b01111111; // 1881 : 127 - 0x7f
      13'h75A: dout <= 8'b01111111; // 1882 : 127 - 0x7f
      13'h75B: dout <= 8'b01111111; // 1883 : 127 - 0x7f
      13'h75C: dout <= 8'b01111111; // 1884 : 127 - 0x7f
      13'h75D: dout <= 8'b01111111; // 1885 : 127 - 0x7f
      13'h75E: dout <= 8'b00000111; // 1886 :   7 - 0x7
      13'h75F: dout <= 8'b00000111; // 1887 :   7 - 0x7
      13'h760: dout <= 8'b11111111; // 1888 : 255 - 0xff -- Sprite 0x76
      13'h761: dout <= 8'b11111111; // 1889 : 255 - 0xff
      13'h762: dout <= 8'b11111111; // 1890 : 255 - 0xff
      13'h763: dout <= 8'b11111111; // 1891 : 255 - 0xff
      13'h764: dout <= 8'b11111111; // 1892 : 255 - 0xff
      13'h765: dout <= 8'b11111111; // 1893 : 255 - 0xff
      13'h766: dout <= 8'b11111111; // 1894 : 255 - 0xff
      13'h767: dout <= 8'b11111111; // 1895 : 255 - 0xff
      13'h768: dout <= 8'b11111110; // 1896 : 254 - 0xfe
      13'h769: dout <= 8'b11111110; // 1897 : 254 - 0xfe
      13'h76A: dout <= 8'b11111110; // 1898 : 254 - 0xfe
      13'h76B: dout <= 8'b11111110; // 1899 : 254 - 0xfe
      13'h76C: dout <= 8'b11111110; // 1900 : 254 - 0xfe
      13'h76D: dout <= 8'b11111110; // 1901 : 254 - 0xfe
      13'h76E: dout <= 8'b11100000; // 1902 : 224 - 0xe0
      13'h76F: dout <= 8'b11100000; // 1903 : 224 - 0xe0
      13'h770: dout <= 8'b11111111; // 1904 : 255 - 0xff -- Sprite 0x77
      13'h771: dout <= 8'b11111111; // 1905 : 255 - 0xff
      13'h772: dout <= 8'b11111111; // 1906 : 255 - 0xff
      13'h773: dout <= 8'b11111111; // 1907 : 255 - 0xff
      13'h774: dout <= 8'b11111111; // 1908 : 255 - 0xff
      13'h775: dout <= 8'b11111111; // 1909 : 255 - 0xff
      13'h776: dout <= 8'b11111111; // 1910 : 255 - 0xff
      13'h777: dout <= 8'b11111111; // 1911 : 255 - 0xff
      13'h778: dout <= 8'b00000111; // 1912 :   7 - 0x7
      13'h779: dout <= 8'b00000111; // 1913 :   7 - 0x7
      13'h77A: dout <= 8'b00000111; // 1914 :   7 - 0x7
      13'h77B: dout <= 8'b00000111; // 1915 :   7 - 0x7
      13'h77C: dout <= 8'b00000111; // 1916 :   7 - 0x7
      13'h77D: dout <= 8'b00000111; // 1917 :   7 - 0x7
      13'h77E: dout <= 8'b00000111; // 1918 :   7 - 0x7
      13'h77F: dout <= 8'b00000111; // 1919 :   7 - 0x7
      13'h780: dout <= 8'b11111111; // 1920 : 255 - 0xff -- Sprite 0x78
      13'h781: dout <= 8'b11111111; // 1921 : 255 - 0xff
      13'h782: dout <= 8'b11111111; // 1922 : 255 - 0xff
      13'h783: dout <= 8'b11111111; // 1923 : 255 - 0xff
      13'h784: dout <= 8'b11111111; // 1924 : 255 - 0xff
      13'h785: dout <= 8'b11111111; // 1925 : 255 - 0xff
      13'h786: dout <= 8'b11111111; // 1926 : 255 - 0xff
      13'h787: dout <= 8'b11111111; // 1927 : 255 - 0xff
      13'h788: dout <= 8'b11100000; // 1928 : 224 - 0xe0
      13'h789: dout <= 8'b11100000; // 1929 : 224 - 0xe0
      13'h78A: dout <= 8'b11100000; // 1930 : 224 - 0xe0
      13'h78B: dout <= 8'b11100000; // 1931 : 224 - 0xe0
      13'h78C: dout <= 8'b11100000; // 1932 : 224 - 0xe0
      13'h78D: dout <= 8'b11100000; // 1933 : 224 - 0xe0
      13'h78E: dout <= 8'b11100000; // 1934 : 224 - 0xe0
      13'h78F: dout <= 8'b11100000; // 1935 : 224 - 0xe0
      13'h790: dout <= 8'b11111111; // 1936 : 255 - 0xff -- Sprite 0x79
      13'h791: dout <= 8'b11111111; // 1937 : 255 - 0xff
      13'h792: dout <= 8'b11111111; // 1938 : 255 - 0xff
      13'h793: dout <= 8'b11111111; // 1939 : 255 - 0xff
      13'h794: dout <= 8'b11111111; // 1940 : 255 - 0xff
      13'h795: dout <= 8'b11111111; // 1941 : 255 - 0xff
      13'h796: dout <= 8'b11111111; // 1942 : 255 - 0xff
      13'h797: dout <= 8'b11111111; // 1943 : 255 - 0xff
      13'h798: dout <= 8'b01111111; // 1944 : 127 - 0x7f
      13'h799: dout <= 8'b01111111; // 1945 : 127 - 0x7f
      13'h79A: dout <= 8'b01111111; // 1946 : 127 - 0x7f
      13'h79B: dout <= 8'b01111111; // 1947 : 127 - 0x7f
      13'h79C: dout <= 8'b01111111; // 1948 : 127 - 0x7f
      13'h79D: dout <= 8'b01111111; // 1949 : 127 - 0x7f
      13'h79E: dout <= 8'b01111110; // 1950 : 126 - 0x7e
      13'h79F: dout <= 8'b01111110; // 1951 : 126 - 0x7e
      13'h7A0: dout <= 8'b11111111; // 1952 : 255 - 0xff -- Sprite 0x7a
      13'h7A1: dout <= 8'b11111111; // 1953 : 255 - 0xff
      13'h7A2: dout <= 8'b11111111; // 1954 : 255 - 0xff
      13'h7A3: dout <= 8'b11111111; // 1955 : 255 - 0xff
      13'h7A4: dout <= 8'b11111111; // 1956 : 255 - 0xff
      13'h7A5: dout <= 8'b11111111; // 1957 : 255 - 0xff
      13'h7A6: dout <= 8'b11111111; // 1958 : 255 - 0xff
      13'h7A7: dout <= 8'b11111111; // 1959 : 255 - 0xff
      13'h7A8: dout <= 8'b11111110; // 1960 : 254 - 0xfe
      13'h7A9: dout <= 8'b11111110; // 1961 : 254 - 0xfe
      13'h7AA: dout <= 8'b11111110; // 1962 : 254 - 0xfe
      13'h7AB: dout <= 8'b11111110; // 1963 : 254 - 0xfe
      13'h7AC: dout <= 8'b11111110; // 1964 : 254 - 0xfe
      13'h7AD: dout <= 8'b11111110; // 1965 : 254 - 0xfe
      13'h7AE: dout <= 8'b00000000; // 1966 :   0 - 0x0
      13'h7AF: dout <= 8'b00000000; // 1967 :   0 - 0x0
      13'h7B0: dout <= 8'b11111111; // 1968 : 255 - 0xff -- Sprite 0x7b
      13'h7B1: dout <= 8'b11111111; // 1969 : 255 - 0xff
      13'h7B2: dout <= 8'b11111111; // 1970 : 255 - 0xff
      13'h7B3: dout <= 8'b11111111; // 1971 : 255 - 0xff
      13'h7B4: dout <= 8'b11111111; // 1972 : 255 - 0xff
      13'h7B5: dout <= 8'b11111111; // 1973 : 255 - 0xff
      13'h7B6: dout <= 8'b11111111; // 1974 : 255 - 0xff
      13'h7B7: dout <= 8'b11111111; // 1975 : 255 - 0xff
      13'h7B8: dout <= 8'b01111110; // 1976 : 126 - 0x7e
      13'h7B9: dout <= 8'b01111111; // 1977 : 127 - 0x7f
      13'h7BA: dout <= 8'b01111111; // 1978 : 127 - 0x7f
      13'h7BB: dout <= 8'b01111111; // 1979 : 127 - 0x7f
      13'h7BC: dout <= 8'b01111111; // 1980 : 127 - 0x7f
      13'h7BD: dout <= 8'b01111111; // 1981 : 127 - 0x7f
      13'h7BE: dout <= 8'b01111111; // 1982 : 127 - 0x7f
      13'h7BF: dout <= 8'b01111110; // 1983 : 126 - 0x7e
      13'h7C0: dout <= 8'b11111111; // 1984 : 255 - 0xff -- Sprite 0x7c
      13'h7C1: dout <= 8'b11111111; // 1985 : 255 - 0xff
      13'h7C2: dout <= 8'b11111111; // 1986 : 255 - 0xff
      13'h7C3: dout <= 8'b11111111; // 1987 : 255 - 0xff
      13'h7C4: dout <= 8'b11111111; // 1988 : 255 - 0xff
      13'h7C5: dout <= 8'b11111111; // 1989 : 255 - 0xff
      13'h7C6: dout <= 8'b11111111; // 1990 : 255 - 0xff
      13'h7C7: dout <= 8'b11111111; // 1991 : 255 - 0xff
      13'h7C8: dout <= 8'b00000000; // 1992 :   0 - 0x0
      13'h7C9: dout <= 8'b11110000; // 1993 : 240 - 0xf0
      13'h7CA: dout <= 8'b11110000; // 1994 : 240 - 0xf0
      13'h7CB: dout <= 8'b11110000; // 1995 : 240 - 0xf0
      13'h7CC: dout <= 8'b11110000; // 1996 : 240 - 0xf0
      13'h7CD: dout <= 8'b11110000; // 1997 : 240 - 0xf0
      13'h7CE: dout <= 8'b11110000; // 1998 : 240 - 0xf0
      13'h7CF: dout <= 8'b00000000; // 1999 :   0 - 0x0
      13'h7D0: dout <= 8'b11111111; // 2000 : 255 - 0xff -- Sprite 0x7d
      13'h7D1: dout <= 8'b11111111; // 2001 : 255 - 0xff
      13'h7D2: dout <= 8'b11111111; // 2002 : 255 - 0xff
      13'h7D3: dout <= 8'b11111111; // 2003 : 255 - 0xff
      13'h7D4: dout <= 8'b11111111; // 2004 : 255 - 0xff
      13'h7D5: dout <= 8'b11111111; // 2005 : 255 - 0xff
      13'h7D6: dout <= 8'b11111111; // 2006 : 255 - 0xff
      13'h7D7: dout <= 8'b11111111; // 2007 : 255 - 0xff
      13'h7D8: dout <= 8'b01111110; // 2008 : 126 - 0x7e
      13'h7D9: dout <= 8'b01111110; // 2009 : 126 - 0x7e
      13'h7DA: dout <= 8'b01111111; // 2010 : 127 - 0x7f
      13'h7DB: dout <= 8'b01111111; // 2011 : 127 - 0x7f
      13'h7DC: dout <= 8'b01111111; // 2012 : 127 - 0x7f
      13'h7DD: dout <= 8'b01111111; // 2013 : 127 - 0x7f
      13'h7DE: dout <= 8'b01111111; // 2014 : 127 - 0x7f
      13'h7DF: dout <= 8'b01111111; // 2015 : 127 - 0x7f
      13'h7E0: dout <= 8'b11111111; // 2016 : 255 - 0xff -- Sprite 0x7e
      13'h7E1: dout <= 8'b11111111; // 2017 : 255 - 0xff
      13'h7E2: dout <= 8'b11111111; // 2018 : 255 - 0xff
      13'h7E3: dout <= 8'b11111111; // 2019 : 255 - 0xff
      13'h7E4: dout <= 8'b11111111; // 2020 : 255 - 0xff
      13'h7E5: dout <= 8'b11111111; // 2021 : 255 - 0xff
      13'h7E6: dout <= 8'b11111111; // 2022 : 255 - 0xff
      13'h7E7: dout <= 8'b11111111; // 2023 : 255 - 0xff
      13'h7E8: dout <= 8'b00000000; // 2024 :   0 - 0x0
      13'h7E9: dout <= 8'b00000000; // 2025 :   0 - 0x0
      13'h7EA: dout <= 8'b11111110; // 2026 : 254 - 0xfe
      13'h7EB: dout <= 8'b11111110; // 2027 : 254 - 0xfe
      13'h7EC: dout <= 8'b11111110; // 2028 : 254 - 0xfe
      13'h7ED: dout <= 8'b11111110; // 2029 : 254 - 0xfe
      13'h7EE: dout <= 8'b11111110; // 2030 : 254 - 0xfe
      13'h7EF: dout <= 8'b11111110; // 2031 : 254 - 0xfe
      13'h7F0: dout <= 8'b11111111; // 2032 : 255 - 0xff -- Sprite 0x7f
      13'h7F1: dout <= 8'b11111111; // 2033 : 255 - 0xff
      13'h7F2: dout <= 8'b11111111; // 2034 : 255 - 0xff
      13'h7F3: dout <= 8'b11111111; // 2035 : 255 - 0xff
      13'h7F4: dout <= 8'b11111111; // 2036 : 255 - 0xff
      13'h7F5: dout <= 8'b11111111; // 2037 : 255 - 0xff
      13'h7F6: dout <= 8'b11111111; // 2038 : 255 - 0xff
      13'h7F7: dout <= 8'b11111111; // 2039 : 255 - 0xff
      13'h7F8: dout <= 8'b01111110; // 2040 : 126 - 0x7e
      13'h7F9: dout <= 8'b11111110; // 2041 : 254 - 0xfe
      13'h7FA: dout <= 8'b11111110; // 2042 : 254 - 0xfe
      13'h7FB: dout <= 8'b11111110; // 2043 : 254 - 0xfe
      13'h7FC: dout <= 8'b11111110; // 2044 : 254 - 0xfe
      13'h7FD: dout <= 8'b11111110; // 2045 : 254 - 0xfe
      13'h7FE: dout <= 8'b11111110; // 2046 : 254 - 0xfe
      13'h7FF: dout <= 8'b01111110; // 2047 : 126 - 0x7e
      13'h800: dout <= 8'b10111111; // 2048 : 191 - 0xbf -- Sprite 0x80
      13'h801: dout <= 8'b11110111; // 2049 : 247 - 0xf7
      13'h802: dout <= 8'b11111101; // 2050 : 253 - 0xfd
      13'h803: dout <= 8'b11011111; // 2051 : 223 - 0xdf
      13'h804: dout <= 8'b11111011; // 2052 : 251 - 0xfb
      13'h805: dout <= 8'b10111111; // 2053 : 191 - 0xbf
      13'h806: dout <= 8'b11111110; // 2054 : 254 - 0xfe
      13'h807: dout <= 8'b11101111; // 2055 : 239 - 0xef
      13'h808: dout <= 8'b01000000; // 2056 :  64 - 0x40
      13'h809: dout <= 8'b00001000; // 2057 :   8 - 0x8
      13'h80A: dout <= 8'b00000010; // 2058 :   2 - 0x2
      13'h80B: dout <= 8'b00100000; // 2059 :  32 - 0x20
      13'h80C: dout <= 8'b00000100; // 2060 :   4 - 0x4
      13'h80D: dout <= 8'b01000000; // 2061 :  64 - 0x40
      13'h80E: dout <= 8'b00000001; // 2062 :   1 - 0x1
      13'h80F: dout <= 8'b00010000; // 2063 :  16 - 0x10
      13'h810: dout <= 8'b11111111; // 2064 : 255 - 0xff -- Sprite 0x81
      13'h811: dout <= 8'b11101110; // 2065 : 238 - 0xee
      13'h812: dout <= 8'b11111111; // 2066 : 255 - 0xff
      13'h813: dout <= 8'b11011111; // 2067 : 223 - 0xdf
      13'h814: dout <= 8'b01110111; // 2068 : 119 - 0x77
      13'h815: dout <= 8'b11111101; // 2069 : 253 - 0xfd
      13'h816: dout <= 8'b11011111; // 2070 : 223 - 0xdf
      13'h817: dout <= 8'b10111111; // 2071 : 191 - 0xbf
      13'h818: dout <= 8'b00000000; // 2072 :   0 - 0x0
      13'h819: dout <= 8'b00010001; // 2073 :  17 - 0x11
      13'h81A: dout <= 8'b00000000; // 2074 :   0 - 0x0
      13'h81B: dout <= 8'b00100000; // 2075 :  32 - 0x20
      13'h81C: dout <= 8'b10001000; // 2076 : 136 - 0x88
      13'h81D: dout <= 8'b00000010; // 2077 :   2 - 0x2
      13'h81E: dout <= 8'b00100000; // 2078 :  32 - 0x20
      13'h81F: dout <= 8'b01000000; // 2079 :  64 - 0x40
      13'h820: dout <= 8'b11111110; // 2080 : 254 - 0xfe -- Sprite 0x82
      13'h821: dout <= 8'b11101111; // 2081 : 239 - 0xef
      13'h822: dout <= 8'b10111111; // 2082 : 191 - 0xbf
      13'h823: dout <= 8'b11110111; // 2083 : 247 - 0xf7
      13'h824: dout <= 8'b11111101; // 2084 : 253 - 0xfd
      13'h825: dout <= 8'b11011111; // 2085 : 223 - 0xdf
      13'h826: dout <= 8'b11111011; // 2086 : 251 - 0xfb
      13'h827: dout <= 8'b10111111; // 2087 : 191 - 0xbf
      13'h828: dout <= 8'b00000001; // 2088 :   1 - 0x1
      13'h829: dout <= 8'b00010000; // 2089 :  16 - 0x10
      13'h82A: dout <= 8'b01000000; // 2090 :  64 - 0x40
      13'h82B: dout <= 8'b00001000; // 2091 :   8 - 0x8
      13'h82C: dout <= 8'b00000010; // 2092 :   2 - 0x2
      13'h82D: dout <= 8'b00100000; // 2093 :  32 - 0x20
      13'h82E: dout <= 8'b00000100; // 2094 :   4 - 0x4
      13'h82F: dout <= 8'b01000000; // 2095 :  64 - 0x40
      13'h830: dout <= 8'b11101111; // 2096 : 239 - 0xef -- Sprite 0x83
      13'h831: dout <= 8'b11111111; // 2097 : 255 - 0xff
      13'h832: dout <= 8'b10111011; // 2098 : 187 - 0xbb
      13'h833: dout <= 8'b11111111; // 2099 : 255 - 0xff
      13'h834: dout <= 8'b11110111; // 2100 : 247 - 0xf7
      13'h835: dout <= 8'b11011101; // 2101 : 221 - 0xdd
      13'h836: dout <= 8'b01111111; // 2102 : 127 - 0x7f
      13'h837: dout <= 8'b11110111; // 2103 : 247 - 0xf7
      13'h838: dout <= 8'b00010000; // 2104 :  16 - 0x10
      13'h839: dout <= 8'b00000000; // 2105 :   0 - 0x0
      13'h83A: dout <= 8'b01000100; // 2106 :  68 - 0x44
      13'h83B: dout <= 8'b00000000; // 2107 :   0 - 0x0
      13'h83C: dout <= 8'b00001000; // 2108 :   8 - 0x8
      13'h83D: dout <= 8'b00100010; // 2109 :  34 - 0x22
      13'h83E: dout <= 8'b10000000; // 2110 : 128 - 0x80
      13'h83F: dout <= 8'b00001000; // 2111 :   8 - 0x8
      13'h840: dout <= 8'b11111111; // 2112 : 255 - 0xff -- Sprite 0x84
      13'h841: dout <= 8'b11101110; // 2113 : 238 - 0xee
      13'h842: dout <= 8'b11111011; // 2114 : 251 - 0xfb
      13'h843: dout <= 8'b10111111; // 2115 : 191 - 0xbf
      13'h844: dout <= 8'b01111111; // 2116 : 127 - 0x7f
      13'h845: dout <= 8'b11101101; // 2117 : 237 - 0xed
      13'h846: dout <= 8'b11111111; // 2118 : 255 - 0xff
      13'h847: dout <= 8'b10111111; // 2119 : 191 - 0xbf
      13'h848: dout <= 8'b00010100; // 2120 :  20 - 0x14
      13'h849: dout <= 8'b10110101; // 2121 : 181 - 0xb5
      13'h84A: dout <= 8'b01000100; // 2122 :  68 - 0x44
      13'h84B: dout <= 8'b01001010; // 2123 :  74 - 0x4a
      13'h84C: dout <= 8'b10010010; // 2124 : 146 - 0x92
      13'h84D: dout <= 8'b10010010; // 2125 : 146 - 0x92
      13'h84E: dout <= 8'b01000100; // 2126 :  68 - 0x44
      13'h84F: dout <= 8'b01001001; // 2127 :  73 - 0x49
      13'h850: dout <= 8'b11111111; // 2128 : 255 - 0xff -- Sprite 0x85
      13'h851: dout <= 8'b10111111; // 2129 : 191 - 0xbf
      13'h852: dout <= 8'b01111101; // 2130 : 125 - 0x7d
      13'h853: dout <= 8'b11110111; // 2131 : 247 - 0xf7
      13'h854: dout <= 8'b11011011; // 2132 : 219 - 0xdb
      13'h855: dout <= 8'b11111101; // 2133 : 253 - 0xfd
      13'h856: dout <= 8'b01111110; // 2134 : 126 - 0x7e
      13'h857: dout <= 8'b11111011; // 2135 : 251 - 0xfb
      13'h858: dout <= 8'b01000010; // 2136 :  66 - 0x42
      13'h859: dout <= 8'b01001010; // 2137 :  74 - 0x4a
      13'h85A: dout <= 8'b11001010; // 2138 : 202 - 0xca
      13'h85B: dout <= 8'b00101001; // 2139 :  41 - 0x29
      13'h85C: dout <= 8'b10100110; // 2140 : 166 - 0xa6
      13'h85D: dout <= 8'b10010010; // 2141 : 146 - 0x92
      13'h85E: dout <= 8'b10001001; // 2142 : 137 - 0x89
      13'h85F: dout <= 8'b00101101; // 2143 :  45 - 0x2d
      13'h860: dout <= 8'b11111111; // 2144 : 255 - 0xff -- Sprite 0x86
      13'h861: dout <= 8'b11110111; // 2145 : 247 - 0xf7
      13'h862: dout <= 8'b11111111; // 2146 : 255 - 0xff
      13'h863: dout <= 8'b11011101; // 2147 : 221 - 0xdd
      13'h864: dout <= 8'b01111111; // 2148 : 127 - 0x7f
      13'h865: dout <= 8'b11110111; // 2149 : 247 - 0xf7
      13'h866: dout <= 8'b11101111; // 2150 : 239 - 0xef
      13'h867: dout <= 8'b10111101; // 2151 : 189 - 0xbd
      13'h868: dout <= 8'b10001000; // 2152 : 136 - 0x88
      13'h869: dout <= 8'b00101001; // 2153 :  41 - 0x29
      13'h86A: dout <= 8'b10000010; // 2154 : 130 - 0x82
      13'h86B: dout <= 8'b10110110; // 2155 : 182 - 0xb6
      13'h86C: dout <= 8'b10001000; // 2156 : 136 - 0x88
      13'h86D: dout <= 8'b01001001; // 2157 :  73 - 0x49
      13'h86E: dout <= 8'b01010010; // 2158 :  82 - 0x52
      13'h86F: dout <= 8'b01010010; // 2159 :  82 - 0x52
      13'h870: dout <= 8'b01011111; // 2160 :  95 - 0x5f -- Sprite 0x87
      13'h871: dout <= 8'b11111101; // 2161 : 253 - 0xfd
      13'h872: dout <= 8'b11110110; // 2162 : 246 - 0xf6
      13'h873: dout <= 8'b01111111; // 2163 : 127 - 0x7f
      13'h874: dout <= 8'b10011111; // 2164 : 159 - 0x9f
      13'h875: dout <= 8'b11111110; // 2165 : 254 - 0xfe
      13'h876: dout <= 8'b11111111; // 2166 : 255 - 0xff
      13'h877: dout <= 8'b11101111; // 2167 : 239 - 0xef
      13'h878: dout <= 8'b10110010; // 2168 : 178 - 0xb2
      13'h879: dout <= 8'b01001010; // 2169 :  74 - 0x4a
      13'h87A: dout <= 8'b10101001; // 2170 : 169 - 0xa9
      13'h87B: dout <= 8'b10100100; // 2171 : 164 - 0xa4
      13'h87C: dout <= 8'b01100010; // 2172 :  98 - 0x62
      13'h87D: dout <= 8'b01001011; // 2173 :  75 - 0x4b
      13'h87E: dout <= 8'b10010000; // 2174 : 144 - 0x90
      13'h87F: dout <= 8'b10010010; // 2175 : 146 - 0x92
      13'h880: dout <= 8'b11111111; // 2176 : 255 - 0xff -- Sprite 0x88
      13'h881: dout <= 8'b11111111; // 2177 : 255 - 0xff
      13'h882: dout <= 8'b10011111; // 2178 : 159 - 0x9f
      13'h883: dout <= 8'b10110011; // 2179 : 179 - 0xb3
      13'h884: dout <= 8'b11110011; // 2180 : 243 - 0xf3
      13'h885: dout <= 8'b11111111; // 2181 : 255 - 0xff
      13'h886: dout <= 8'b11111111; // 2182 : 255 - 0xff
      13'h887: dout <= 8'b11111111; // 2183 : 255 - 0xff
      13'h888: dout <= 8'b00000000; // 2184 :   0 - 0x0
      13'h889: dout <= 8'b01100000; // 2185 :  96 - 0x60
      13'h88A: dout <= 8'b11111110; // 2186 : 254 - 0xfe
      13'h88B: dout <= 8'b11111111; // 2187 : 255 - 0xff
      13'h88C: dout <= 8'b01111111; // 2188 : 127 - 0x7f
      13'h88D: dout <= 8'b00011111; // 2189 :  31 - 0x1f
      13'h88E: dout <= 8'b00001110; // 2190 :  14 - 0xe
      13'h88F: dout <= 8'b00000000; // 2191 :   0 - 0x0
      13'h890: dout <= 8'b11111111; // 2192 : 255 - 0xff -- Sprite 0x89
      13'h891: dout <= 8'b11001111; // 2193 : 207 - 0xcf
      13'h892: dout <= 8'b11011111; // 2194 : 223 - 0xdf
      13'h893: dout <= 8'b11111111; // 2195 : 255 - 0xff
      13'h894: dout <= 8'b11110011; // 2196 : 243 - 0xf3
      13'h895: dout <= 8'b11110011; // 2197 : 243 - 0xf3
      13'h896: dout <= 8'b11111111; // 2198 : 255 - 0xff
      13'h897: dout <= 8'b11111111; // 2199 : 255 - 0xff
      13'h898: dout <= 8'b00110000; // 2200 :  48 - 0x30
      13'h899: dout <= 8'b01111000; // 2201 : 120 - 0x78
      13'h89A: dout <= 8'b01111000; // 2202 : 120 - 0x78
      13'h89B: dout <= 8'b00111110; // 2203 :  62 - 0x3e
      13'h89C: dout <= 8'b00011111; // 2204 :  31 - 0x1f
      13'h89D: dout <= 8'b00011111; // 2205 :  31 - 0x1f
      13'h89E: dout <= 8'b00011111; // 2206 :  31 - 0x1f
      13'h89F: dout <= 8'b00001110; // 2207 :  14 - 0xe
      13'h8A0: dout <= 8'b10111111; // 2208 : 191 - 0xbf -- Sprite 0x8a
      13'h8A1: dout <= 8'b11110111; // 2209 : 247 - 0xf7
      13'h8A2: dout <= 8'b11111101; // 2210 : 253 - 0xfd
      13'h8A3: dout <= 8'b11111111; // 2211 : 255 - 0xff
      13'h8A4: dout <= 8'b11111011; // 2212 : 251 - 0xfb
      13'h8A5: dout <= 8'b10111111; // 2213 : 191 - 0xbf
      13'h8A6: dout <= 8'b11111110; // 2214 : 254 - 0xfe
      13'h8A7: dout <= 8'b11101111; // 2215 : 239 - 0xef
      13'h8A8: dout <= 8'b01000000; // 2216 :  64 - 0x40
      13'h8A9: dout <= 8'b00001000; // 2217 :   8 - 0x8
      13'h8AA: dout <= 8'b00000010; // 2218 :   2 - 0x2
      13'h8AB: dout <= 8'b00101000; // 2219 :  40 - 0x28
      13'h8AC: dout <= 8'b00010100; // 2220 :  20 - 0x14
      13'h8AD: dout <= 8'b01010100; // 2221 :  84 - 0x54
      13'h8AE: dout <= 8'b00000001; // 2222 :   1 - 0x1
      13'h8AF: dout <= 8'b00010000; // 2223 :  16 - 0x10
      13'h8B0: dout <= 8'b10111111; // 2224 : 191 - 0xbf -- Sprite 0x8b
      13'h8B1: dout <= 8'b11111111; // 2225 : 255 - 0xff
      13'h8B2: dout <= 8'b11101110; // 2226 : 238 - 0xee
      13'h8B3: dout <= 8'b11111111; // 2227 : 255 - 0xff
      13'h8B4: dout <= 8'b11011111; // 2228 : 223 - 0xdf
      13'h8B5: dout <= 8'b01111101; // 2229 : 125 - 0x7d
      13'h8B6: dout <= 8'b11111111; // 2230 : 255 - 0xff
      13'h8B7: dout <= 8'b11011111; // 2231 : 223 - 0xdf
      13'h8B8: dout <= 8'b01000000; // 2232 :  64 - 0x40
      13'h8B9: dout <= 8'b00000000; // 2233 :   0 - 0x0
      13'h8BA: dout <= 8'b10010001; // 2234 : 145 - 0x91
      13'h8BB: dout <= 8'b00010100; // 2235 :  20 - 0x14
      13'h8BC: dout <= 8'b00101000; // 2236 :  40 - 0x28
      13'h8BD: dout <= 8'b10001010; // 2237 : 138 - 0x8a
      13'h8BE: dout <= 8'b01000000; // 2238 :  64 - 0x40
      13'h8BF: dout <= 8'b00100000; // 2239 :  32 - 0x20
      13'h8C0: dout <= 8'b11111111; // 2240 : 255 - 0xff -- Sprite 0x8c
      13'h8C1: dout <= 8'b11111000; // 2241 : 248 - 0xf8
      13'h8C2: dout <= 8'b11100010; // 2242 : 226 - 0xe2
      13'h8C3: dout <= 8'b11010111; // 2243 : 215 - 0xd7
      13'h8C4: dout <= 8'b11001111; // 2244 : 207 - 0xcf
      13'h8C5: dout <= 8'b10011111; // 2245 : 159 - 0x9f
      13'h8C6: dout <= 8'b10111110; // 2246 : 190 - 0xbe
      13'h8C7: dout <= 8'b10011101; // 2247 : 157 - 0x9d
      13'h8C8: dout <= 8'b00000000; // 2248 :   0 - 0x0
      13'h8C9: dout <= 8'b00000111; // 2249 :   7 - 0x7
      13'h8CA: dout <= 8'b00011111; // 2250 :  31 - 0x1f
      13'h8CB: dout <= 8'b00111111; // 2251 :  63 - 0x3f
      13'h8CC: dout <= 8'b00111111; // 2252 :  63 - 0x3f
      13'h8CD: dout <= 8'b01111111; // 2253 : 127 - 0x7f
      13'h8CE: dout <= 8'b01111111; // 2254 : 127 - 0x7f
      13'h8CF: dout <= 8'b01111111; // 2255 : 127 - 0x7f
      13'h8D0: dout <= 8'b11111111; // 2256 : 255 - 0xff -- Sprite 0x8d
      13'h8D1: dout <= 8'b00011111; // 2257 :  31 - 0x1f
      13'h8D2: dout <= 8'b10100111; // 2258 : 167 - 0xa7
      13'h8D3: dout <= 8'b11000011; // 2259 : 195 - 0xc3
      13'h8D4: dout <= 8'b11100011; // 2260 : 227 - 0xe3
      13'h8D5: dout <= 8'b01000001; // 2261 :  65 - 0x41
      13'h8D6: dout <= 8'b10100001; // 2262 : 161 - 0xa1
      13'h8D7: dout <= 8'b00000001; // 2263 :   1 - 0x1
      13'h8D8: dout <= 8'b00000000; // 2264 :   0 - 0x0
      13'h8D9: dout <= 8'b11100000; // 2265 : 224 - 0xe0
      13'h8DA: dout <= 8'b11111000; // 2266 : 248 - 0xf8
      13'h8DB: dout <= 8'b11111000; // 2267 : 248 - 0xf8
      13'h8DC: dout <= 8'b11110000; // 2268 : 240 - 0xf0
      13'h8DD: dout <= 8'b11111000; // 2269 : 248 - 0xf8
      13'h8DE: dout <= 8'b11110100; // 2270 : 244 - 0xf4
      13'h8DF: dout <= 8'b11111000; // 2271 : 248 - 0xf8
      13'h8E0: dout <= 8'b10111110; // 2272 : 190 - 0xbe -- Sprite 0x8e
      13'h8E1: dout <= 8'b11111111; // 2273 : 255 - 0xff
      13'h8E2: dout <= 8'b11011111; // 2274 : 223 - 0xdf
      13'h8E3: dout <= 8'b11111111; // 2275 : 255 - 0xff
      13'h8E4: dout <= 8'b11101111; // 2276 : 239 - 0xef
      13'h8E5: dout <= 8'b11111111; // 2277 : 255 - 0xff
      13'h8E6: dout <= 8'b11110111; // 2278 : 247 - 0xf7
      13'h8E7: dout <= 8'b11111111; // 2279 : 255 - 0xff
      13'h8E8: dout <= 8'b01111111; // 2280 : 127 - 0x7f
      13'h8E9: dout <= 8'b00111111; // 2281 :  63 - 0x3f
      13'h8EA: dout <= 8'b00111111; // 2282 :  63 - 0x3f
      13'h8EB: dout <= 8'b00011111; // 2283 :  31 - 0x1f
      13'h8EC: dout <= 8'b00011111; // 2284 :  31 - 0x1f
      13'h8ED: dout <= 8'b00001111; // 2285 :  15 - 0xf
      13'h8EE: dout <= 8'b00001111; // 2286 :  15 - 0xf
      13'h8EF: dout <= 8'b00000111; // 2287 :   7 - 0x7
      13'h8F0: dout <= 8'b01111101; // 2288 : 125 - 0x7d -- Sprite 0x8f
      13'h8F1: dout <= 8'b11111111; // 2289 : 255 - 0xff
      13'h8F2: dout <= 8'b11111011; // 2290 : 251 - 0xfb
      13'h8F3: dout <= 8'b11111111; // 2291 : 255 - 0xff
      13'h8F4: dout <= 8'b11110111; // 2292 : 247 - 0xf7
      13'h8F5: dout <= 8'b11111111; // 2293 : 255 - 0xff
      13'h8F6: dout <= 8'b11101111; // 2294 : 239 - 0xef
      13'h8F7: dout <= 8'b11111111; // 2295 : 255 - 0xff
      13'h8F8: dout <= 8'b11111110; // 2296 : 254 - 0xfe
      13'h8F9: dout <= 8'b11111100; // 2297 : 252 - 0xfc
      13'h8FA: dout <= 8'b11111100; // 2298 : 252 - 0xfc
      13'h8FB: dout <= 8'b11111000; // 2299 : 248 - 0xf8
      13'h8FC: dout <= 8'b11111000; // 2300 : 248 - 0xf8
      13'h8FD: dout <= 8'b11110000; // 2301 : 240 - 0xf0
      13'h8FE: dout <= 8'b11110000; // 2302 : 240 - 0xf0
      13'h8FF: dout <= 8'b11100000; // 2303 : 224 - 0xe0
      13'h900: dout <= 8'b10111110; // 2304 : 190 - 0xbe -- Sprite 0x90
      13'h901: dout <= 8'b11110111; // 2305 : 247 - 0xf7
      13'h902: dout <= 8'b11111111; // 2306 : 255 - 0xff
      13'h903: dout <= 8'b11011111; // 2307 : 223 - 0xdf
      13'h904: dout <= 8'b11111011; // 2308 : 251 - 0xfb
      13'h905: dout <= 8'b11111110; // 2309 : 254 - 0xfe
      13'h906: dout <= 8'b10111111; // 2310 : 191 - 0xbf
      13'h907: dout <= 8'b11110111; // 2311 : 247 - 0xf7
      13'h908: dout <= 8'b01000001; // 2312 :  65 - 0x41
      13'h909: dout <= 8'b00001000; // 2313 :   8 - 0x8
      13'h90A: dout <= 8'b00000000; // 2314 :   0 - 0x0
      13'h90B: dout <= 8'b00100000; // 2315 :  32 - 0x20
      13'h90C: dout <= 8'b00000100; // 2316 :   4 - 0x4
      13'h90D: dout <= 8'b00000001; // 2317 :   1 - 0x1
      13'h90E: dout <= 8'b01000000; // 2318 :  64 - 0x40
      13'h90F: dout <= 8'b00001000; // 2319 :   8 - 0x8
      13'h910: dout <= 8'b11101110; // 2320 : 238 - 0xee -- Sprite 0x91
      13'h911: dout <= 8'b11111111; // 2321 : 255 - 0xff
      13'h912: dout <= 8'b01111011; // 2322 : 123 - 0x7b
      13'h913: dout <= 8'b11111101; // 2323 : 253 - 0xfd
      13'h914: dout <= 8'b11101111; // 2324 : 239 - 0xef
      13'h915: dout <= 8'b11111111; // 2325 : 255 - 0xff
      13'h916: dout <= 8'b10111101; // 2326 : 189 - 0xbd
      13'h917: dout <= 8'b11111111; // 2327 : 255 - 0xff
      13'h918: dout <= 8'b00010001; // 2328 :  17 - 0x11
      13'h919: dout <= 8'b00000000; // 2329 :   0 - 0x0
      13'h91A: dout <= 8'b10000100; // 2330 : 132 - 0x84
      13'h91B: dout <= 8'b00000010; // 2331 :   2 - 0x2
      13'h91C: dout <= 8'b00010000; // 2332 :  16 - 0x10
      13'h91D: dout <= 8'b00000000; // 2333 :   0 - 0x0
      13'h91E: dout <= 8'b01000010; // 2334 :  66 - 0x42
      13'h91F: dout <= 8'b00000000; // 2335 :   0 - 0x0
      13'h920: dout <= 8'b11111011; // 2336 : 251 - 0xfb -- Sprite 0x92
      13'h921: dout <= 8'b10111111; // 2337 : 191 - 0xbf
      13'h922: dout <= 8'b11101111; // 2338 : 239 - 0xef
      13'h923: dout <= 8'b11111101; // 2339 : 253 - 0xfd
      13'h924: dout <= 8'b11111111; // 2340 : 255 - 0xff
      13'h925: dout <= 8'b10111111; // 2341 : 191 - 0xbf
      13'h926: dout <= 8'b11111011; // 2342 : 251 - 0xfb
      13'h927: dout <= 8'b11011111; // 2343 : 223 - 0xdf
      13'h928: dout <= 8'b00000100; // 2344 :   4 - 0x4
      13'h929: dout <= 8'b01000000; // 2345 :  64 - 0x40
      13'h92A: dout <= 8'b00010000; // 2346 :  16 - 0x10
      13'h92B: dout <= 8'b00000010; // 2347 :   2 - 0x2
      13'h92C: dout <= 8'b00000000; // 2348 :   0 - 0x0
      13'h92D: dout <= 8'b01000000; // 2349 :  64 - 0x40
      13'h92E: dout <= 8'b00000100; // 2350 :   4 - 0x4
      13'h92F: dout <= 8'b00100000; // 2351 :  32 - 0x20
      13'h930: dout <= 8'b10111101; // 2352 : 189 - 0xbd -- Sprite 0x93
      13'h931: dout <= 8'b11111111; // 2353 : 255 - 0xff
      13'h932: dout <= 8'b01110111; // 2354 : 119 - 0x77
      13'h933: dout <= 8'b11111110; // 2355 : 254 - 0xfe
      13'h934: dout <= 8'b11011111; // 2356 : 223 - 0xdf
      13'h935: dout <= 8'b11111011; // 2357 : 251 - 0xfb
      13'h936: dout <= 8'b11101111; // 2358 : 239 - 0xef
      13'h937: dout <= 8'b01111111; // 2359 : 127 - 0x7f
      13'h938: dout <= 8'b01000010; // 2360 :  66 - 0x42
      13'h939: dout <= 8'b00000000; // 2361 :   0 - 0x0
      13'h93A: dout <= 8'b10001000; // 2362 : 136 - 0x88
      13'h93B: dout <= 8'b00000001; // 2363 :   1 - 0x1
      13'h93C: dout <= 8'b00100000; // 2364 :  32 - 0x20
      13'h93D: dout <= 8'b00000100; // 2365 :   4 - 0x4
      13'h93E: dout <= 8'b00010000; // 2366 :  16 - 0x10
      13'h93F: dout <= 8'b10000000; // 2367 : 128 - 0x80
      13'h940: dout <= 8'b01111111; // 2368 : 127 - 0x7f -- Sprite 0x94
      13'h941: dout <= 8'b11110111; // 2369 : 247 - 0xf7
      13'h942: dout <= 8'b11011101; // 2370 : 221 - 0xdd
      13'h943: dout <= 8'b01111011; // 2371 : 123 - 0x7b
      13'h944: dout <= 8'b11111111; // 2372 : 255 - 0xff
      13'h945: dout <= 8'b11101110; // 2373 : 238 - 0xee
      13'h946: dout <= 8'b10111011; // 2374 : 187 - 0xbb
      13'h947: dout <= 8'b11111101; // 2375 : 253 - 0xfd
      13'h948: dout <= 8'b11001000; // 2376 : 200 - 0xc8
      13'h949: dout <= 8'b00101010; // 2377 :  42 - 0x2a
      13'h94A: dout <= 8'b10100010; // 2378 : 162 - 0xa2
      13'h94B: dout <= 8'b10010100; // 2379 : 148 - 0x94
      13'h94C: dout <= 8'b10010001; // 2380 : 145 - 0x91
      13'h94D: dout <= 8'b01010101; // 2381 :  85 - 0x55
      13'h94E: dout <= 8'b01000100; // 2382 :  68 - 0x44
      13'h94F: dout <= 8'b00010010; // 2383 :  18 - 0x12
      13'h950: dout <= 8'b11010111; // 2384 : 215 - 0xd7 -- Sprite 0x95
      13'h951: dout <= 8'b01111111; // 2385 : 127 - 0x7f
      13'h952: dout <= 8'b11111101; // 2386 : 253 - 0xfd
      13'h953: dout <= 8'b11101110; // 2387 : 238 - 0xee
      13'h954: dout <= 8'b11110111; // 2388 : 247 - 0xf7
      13'h955: dout <= 8'b10111011; // 2389 : 187 - 0xbb
      13'h956: dout <= 8'b11101111; // 2390 : 239 - 0xef
      13'h957: dout <= 8'b11110111; // 2391 : 247 - 0xf7
      13'h958: dout <= 8'b10101010; // 2392 : 170 - 0xaa
      13'h959: dout <= 8'b10100010; // 2393 : 162 - 0xa2
      13'h95A: dout <= 8'b00010010; // 2394 :  18 - 0x12
      13'h95B: dout <= 8'b01010011; // 2395 :  83 - 0x53
      13'h95C: dout <= 8'b01001100; // 2396 :  76 - 0x4c
      13'h95D: dout <= 8'b01010101; // 2397 :  85 - 0x55
      13'h95E: dout <= 8'b10010001; // 2398 : 145 - 0x91
      13'h95F: dout <= 8'b01001000; // 2399 :  72 - 0x48
      13'h960: dout <= 8'b10111111; // 2400 : 191 - 0xbf -- Sprite 0x96
      13'h961: dout <= 8'b11101110; // 2401 : 238 - 0xee
      13'h962: dout <= 8'b11011011; // 2402 : 219 - 0xdb
      13'h963: dout <= 8'b11111111; // 2403 : 255 - 0xff
      13'h964: dout <= 8'b01110111; // 2404 : 119 - 0x77
      13'h965: dout <= 8'b11011101; // 2405 : 221 - 0xdd
      13'h966: dout <= 8'b11101111; // 2406 : 239 - 0xef
      13'h967: dout <= 8'b11111011; // 2407 : 251 - 0xfb
      13'h968: dout <= 8'b01010001; // 2408 :  81 - 0x51
      13'h969: dout <= 8'b00010101; // 2409 :  21 - 0x15
      13'h96A: dout <= 8'b10100100; // 2410 : 164 - 0xa4
      13'h96B: dout <= 8'b10001100; // 2411 : 140 - 0x8c
      13'h96C: dout <= 8'b10101010; // 2412 : 170 - 0xaa
      13'h96D: dout <= 8'b00100010; // 2413 :  34 - 0x22
      13'h96E: dout <= 8'b10010000; // 2414 : 144 - 0x90
      13'h96F: dout <= 8'b01000110; // 2415 :  70 - 0x46
      13'h970: dout <= 8'b11111101; // 2416 : 253 - 0xfd -- Sprite 0x97
      13'h971: dout <= 8'b11101110; // 2417 : 238 - 0xee
      13'h972: dout <= 8'b11111011; // 2418 : 251 - 0xfb
      13'h973: dout <= 8'b11111101; // 2419 : 253 - 0xfd
      13'h974: dout <= 8'b11110101; // 2420 : 245 - 0xf5
      13'h975: dout <= 8'b11011111; // 2421 : 223 - 0xdf
      13'h976: dout <= 8'b01111111; // 2422 : 127 - 0x7f
      13'h977: dout <= 8'b10111011; // 2423 : 187 - 0xbb
      13'h978: dout <= 8'b00010011; // 2424 :  19 - 0x13
      13'h979: dout <= 8'b01010101; // 2425 :  85 - 0x55
      13'h97A: dout <= 8'b01100100; // 2426 : 100 - 0x64
      13'h97B: dout <= 8'b00010010; // 2427 :  18 - 0x12
      13'h97C: dout <= 8'b10101010; // 2428 : 170 - 0xaa
      13'h97D: dout <= 8'b10101000; // 2429 : 168 - 0xa8
      13'h97E: dout <= 8'b10000100; // 2430 : 132 - 0x84
      13'h97F: dout <= 8'b11010100; // 2431 : 212 - 0xd4
      13'h980: dout <= 8'b11111111; // 2432 : 255 - 0xff -- Sprite 0x98
      13'h981: dout <= 8'b11001111; // 2433 : 207 - 0xcf
      13'h982: dout <= 8'b11011111; // 2434 : 223 - 0xdf
      13'h983: dout <= 8'b11111111; // 2435 : 255 - 0xff
      13'h984: dout <= 8'b11110011; // 2436 : 243 - 0xf3
      13'h985: dout <= 8'b11110011; // 2437 : 243 - 0xf3
      13'h986: dout <= 8'b11111111; // 2438 : 255 - 0xff
      13'h987: dout <= 8'b11111111; // 2439 : 255 - 0xff
      13'h988: dout <= 8'b00110000; // 2440 :  48 - 0x30
      13'h989: dout <= 8'b01111000; // 2441 : 120 - 0x78
      13'h98A: dout <= 8'b01111000; // 2442 : 120 - 0x78
      13'h98B: dout <= 8'b00111110; // 2443 :  62 - 0x3e
      13'h98C: dout <= 8'b00011111; // 2444 :  31 - 0x1f
      13'h98D: dout <= 8'b00011111; // 2445 :  31 - 0x1f
      13'h98E: dout <= 8'b00011111; // 2446 :  31 - 0x1f
      13'h98F: dout <= 8'b00001110; // 2447 :  14 - 0xe
      13'h990: dout <= 8'b11111111; // 2448 : 255 - 0xff -- Sprite 0x99
      13'h991: dout <= 8'b11111111; // 2449 : 255 - 0xff
      13'h992: dout <= 8'b10011111; // 2450 : 159 - 0x9f
      13'h993: dout <= 8'b10110011; // 2451 : 179 - 0xb3
      13'h994: dout <= 8'b11110011; // 2452 : 243 - 0xf3
      13'h995: dout <= 8'b11111111; // 2453 : 255 - 0xff
      13'h996: dout <= 8'b11111111; // 2454 : 255 - 0xff
      13'h997: dout <= 8'b11111111; // 2455 : 255 - 0xff
      13'h998: dout <= 8'b00000000; // 2456 :   0 - 0x0
      13'h999: dout <= 8'b01100000; // 2457 :  96 - 0x60
      13'h99A: dout <= 8'b11111110; // 2458 : 254 - 0xfe
      13'h99B: dout <= 8'b11111111; // 2459 : 255 - 0xff
      13'h99C: dout <= 8'b01111111; // 2460 : 127 - 0x7f
      13'h99D: dout <= 8'b00011111; // 2461 :  31 - 0x1f
      13'h99E: dout <= 8'b00001110; // 2462 :  14 - 0xe
      13'h99F: dout <= 8'b00000000; // 2463 :   0 - 0x0
      13'h9A0: dout <= 8'b10111111; // 2464 : 191 - 0xbf -- Sprite 0x9a
      13'h9A1: dout <= 8'b11110111; // 2465 : 247 - 0xf7
      13'h9A2: dout <= 8'b11111111; // 2466 : 255 - 0xff
      13'h9A3: dout <= 8'b11011111; // 2467 : 223 - 0xdf
      13'h9A4: dout <= 8'b11111011; // 2468 : 251 - 0xfb
      13'h9A5: dout <= 8'b11111111; // 2469 : 255 - 0xff
      13'h9A6: dout <= 8'b10111111; // 2470 : 191 - 0xbf
      13'h9A7: dout <= 8'b11110111; // 2471 : 247 - 0xf7
      13'h9A8: dout <= 8'b01000000; // 2472 :  64 - 0x40
      13'h9A9: dout <= 8'b00001100; // 2473 :  12 - 0xc
      13'h9AA: dout <= 8'b00000000; // 2474 :   0 - 0x0
      13'h9AB: dout <= 8'b00101000; // 2475 :  40 - 0x28
      13'h9AC: dout <= 8'b00101100; // 2476 :  44 - 0x2c
      13'h9AD: dout <= 8'b00010001; // 2477 :  17 - 0x11
      13'h9AE: dout <= 8'b01000000; // 2478 :  64 - 0x40
      13'h9AF: dout <= 8'b00001000; // 2479 :   8 - 0x8
      13'h9B0: dout <= 8'b11011111; // 2480 : 223 - 0xdf -- Sprite 0x9b
      13'h9B1: dout <= 8'b11111111; // 2481 : 255 - 0xff
      13'h9B2: dout <= 8'b01111011; // 2482 : 123 - 0x7b
      13'h9B3: dout <= 8'b11111111; // 2483 : 255 - 0xff
      13'h9B4: dout <= 8'b11101111; // 2484 : 239 - 0xef
      13'h9B5: dout <= 8'b11111101; // 2485 : 253 - 0xfd
      13'h9B6: dout <= 8'b10111111; // 2486 : 191 - 0xbf
      13'h9B7: dout <= 8'b11111111; // 2487 : 255 - 0xff
      13'h9B8: dout <= 8'b00100000; // 2488 :  32 - 0x20
      13'h9B9: dout <= 8'b00000000; // 2489 :   0 - 0x0
      13'h9BA: dout <= 8'b10010100; // 2490 : 148 - 0x94
      13'h9BB: dout <= 8'b01001000; // 2491 :  72 - 0x48
      13'h9BC: dout <= 8'b00011000; // 2492 :  24 - 0x18
      13'h9BD: dout <= 8'b00000110; // 2493 :   6 - 0x6
      13'h9BE: dout <= 8'b01000000; // 2494 :  64 - 0x40
      13'h9BF: dout <= 8'b00000000; // 2495 :   0 - 0x0
      13'h9C0: dout <= 8'b10111010; // 2496 : 186 - 0xba -- Sprite 0x9c
      13'h9C1: dout <= 8'b10011100; // 2497 : 156 - 0x9c
      13'h9C2: dout <= 8'b10101010; // 2498 : 170 - 0xaa
      13'h9C3: dout <= 8'b11000000; // 2499 : 192 - 0xc0
      13'h9C4: dout <= 8'b11000000; // 2500 : 192 - 0xc0
      13'h9C5: dout <= 8'b11100000; // 2501 : 224 - 0xe0
      13'h9C6: dout <= 8'b11111000; // 2502 : 248 - 0xf8
      13'h9C7: dout <= 8'b11111111; // 2503 : 255 - 0xff
      13'h9C8: dout <= 8'b01111111; // 2504 : 127 - 0x7f
      13'h9C9: dout <= 8'b01111111; // 2505 : 127 - 0x7f
      13'h9CA: dout <= 8'b01111111; // 2506 : 127 - 0x7f
      13'h9CB: dout <= 8'b00111111; // 2507 :  63 - 0x3f
      13'h9CC: dout <= 8'b00110101; // 2508 :  53 - 0x35
      13'h9CD: dout <= 8'b00000010; // 2509 :   2 - 0x2
      13'h9CE: dout <= 8'b00000000; // 2510 :   0 - 0x0
      13'h9CF: dout <= 8'b00000000; // 2511 :   0 - 0x0
      13'h9D0: dout <= 8'b00000001; // 2512 :   1 - 0x1 -- Sprite 0x9d
      13'h9D1: dout <= 8'b00000001; // 2513 :   1 - 0x1
      13'h9D2: dout <= 8'b00000001; // 2514 :   1 - 0x1
      13'h9D3: dout <= 8'b00000011; // 2515 :   3 - 0x3
      13'h9D4: dout <= 8'b00000011; // 2516 :   3 - 0x3
      13'h9D5: dout <= 8'b00000111; // 2517 :   7 - 0x7
      13'h9D6: dout <= 8'b00011111; // 2518 :  31 - 0x1f
      13'h9D7: dout <= 8'b11111111; // 2519 : 255 - 0xff
      13'h9D8: dout <= 8'b11110100; // 2520 : 244 - 0xf4
      13'h9D9: dout <= 8'b11111000; // 2521 : 248 - 0xf8
      13'h9DA: dout <= 8'b11110000; // 2522 : 240 - 0xf0
      13'h9DB: dout <= 8'b11101000; // 2523 : 232 - 0xe8
      13'h9DC: dout <= 8'b01010000; // 2524 :  80 - 0x50
      13'h9DD: dout <= 8'b10000000; // 2525 : 128 - 0x80
      13'h9DE: dout <= 8'b00000000; // 2526 :   0 - 0x0
      13'h9DF: dout <= 8'b00000000; // 2527 :   0 - 0x0
      13'h9E0: dout <= 8'b01111101; // 2528 : 125 - 0x7d -- Sprite 0x9e
      13'h9E1: dout <= 8'b11111111; // 2529 : 255 - 0xff
      13'h9E2: dout <= 8'b11111011; // 2530 : 251 - 0xfb
      13'h9E3: dout <= 8'b11111111; // 2531 : 255 - 0xff
      13'h9E4: dout <= 8'b11111111; // 2532 : 255 - 0xff
      13'h9E5: dout <= 8'b11111011; // 2533 : 251 - 0xfb
      13'h9E6: dout <= 8'b11111111; // 2534 : 255 - 0xff
      13'h9E7: dout <= 8'b01111101; // 2535 : 125 - 0x7d
      13'h9E8: dout <= 8'b11111110; // 2536 : 254 - 0xfe
      13'h9E9: dout <= 8'b11111100; // 2537 : 252 - 0xfc
      13'h9EA: dout <= 8'b11111100; // 2538 : 252 - 0xfc
      13'h9EB: dout <= 8'b11111000; // 2539 : 248 - 0xf8
      13'h9EC: dout <= 8'b11111000; // 2540 : 248 - 0xf8
      13'h9ED: dout <= 8'b11111100; // 2541 : 252 - 0xfc
      13'h9EE: dout <= 8'b11111100; // 2542 : 252 - 0xfc
      13'h9EF: dout <= 8'b11111110; // 2543 : 254 - 0xfe
      13'h9F0: dout <= 8'b11111111; // 2544 : 255 - 0xff -- Sprite 0x9f
      13'h9F1: dout <= 8'b11111111; // 2545 : 255 - 0xff
      13'h9F2: dout <= 8'b10111101; // 2546 : 189 - 0xbd
      13'h9F3: dout <= 8'b11111111; // 2547 : 255 - 0xff
      13'h9F4: dout <= 8'b11111111; // 2548 : 255 - 0xff
      13'h9F5: dout <= 8'b11111111; // 2549 : 255 - 0xff
      13'h9F6: dout <= 8'b11111111; // 2550 : 255 - 0xff
      13'h9F7: dout <= 8'b10111101; // 2551 : 189 - 0xbd
      13'h9F8: dout <= 8'b00000000; // 2552 :   0 - 0x0
      13'h9F9: dout <= 8'b00000000; // 2553 :   0 - 0x0
      13'h9FA: dout <= 8'b01111110; // 2554 : 126 - 0x7e
      13'h9FB: dout <= 8'b01111110; // 2555 : 126 - 0x7e
      13'h9FC: dout <= 8'b01111110; // 2556 : 126 - 0x7e
      13'h9FD: dout <= 8'b01111110; // 2557 : 126 - 0x7e
      13'h9FE: dout <= 8'b01111110; // 2558 : 126 - 0x7e
      13'h9FF: dout <= 8'b01111110; // 2559 : 126 - 0x7e
      13'hA00: dout <= 8'b11101111; // 2560 : 239 - 0xef -- Sprite 0xa0
      13'hA01: dout <= 8'b11000111; // 2561 : 199 - 0xc7
      13'hA02: dout <= 8'b10000011; // 2562 : 131 - 0x83
      13'hA03: dout <= 8'b00000111; // 2563 :   7 - 0x7
      13'hA04: dout <= 8'b10001111; // 2564 : 143 - 0x8f
      13'hA05: dout <= 8'b11011101; // 2565 : 221 - 0xdd
      13'hA06: dout <= 8'b11111010; // 2566 : 250 - 0xfa
      13'hA07: dout <= 8'b11111101; // 2567 : 253 - 0xfd
      13'hA08: dout <= 8'b00010000; // 2568 :  16 - 0x10
      13'hA09: dout <= 8'b00111000; // 2569 :  56 - 0x38
      13'hA0A: dout <= 8'b01111100; // 2570 : 124 - 0x7c
      13'hA0B: dout <= 8'b11111000; // 2571 : 248 - 0xf8
      13'hA0C: dout <= 8'b01110000; // 2572 : 112 - 0x70
      13'hA0D: dout <= 8'b00100010; // 2573 :  34 - 0x22
      13'hA0E: dout <= 8'b00000101; // 2574 :   5 - 0x5
      13'hA0F: dout <= 8'b00000010; // 2575 :   2 - 0x2
      13'hA10: dout <= 8'b11101111; // 2576 : 239 - 0xef -- Sprite 0xa1
      13'hA11: dout <= 8'b11000111; // 2577 : 199 - 0xc7
      13'hA12: dout <= 8'b10000011; // 2578 : 131 - 0x83
      13'hA13: dout <= 8'b00011111; // 2579 :  31 - 0x1f
      13'hA14: dout <= 8'b10010000; // 2580 : 144 - 0x90
      13'hA15: dout <= 8'b11010100; // 2581 : 212 - 0xd4
      13'hA16: dout <= 8'b11110011; // 2582 : 243 - 0xf3
      13'hA17: dout <= 8'b11110010; // 2583 : 242 - 0xf2
      13'hA18: dout <= 8'b00010000; // 2584 :  16 - 0x10
      13'hA19: dout <= 8'b00111000; // 2585 :  56 - 0x38
      13'hA1A: dout <= 8'b01111100; // 2586 : 124 - 0x7c
      13'hA1B: dout <= 8'b11100000; // 2587 : 224 - 0xe0
      13'hA1C: dout <= 8'b01100000; // 2588 :  96 - 0x60
      13'hA1D: dout <= 8'b00100000; // 2589 :  32 - 0x20
      13'hA1E: dout <= 8'b00000000; // 2590 :   0 - 0x0
      13'hA1F: dout <= 8'b00000000; // 2591 :   0 - 0x0
      13'hA20: dout <= 8'b11101111; // 2592 : 239 - 0xef -- Sprite 0xa2
      13'hA21: dout <= 8'b11000111; // 2593 : 199 - 0xc7
      13'hA22: dout <= 8'b10000011; // 2594 : 131 - 0x83
      13'hA23: dout <= 8'b11111111; // 2595 : 255 - 0xff
      13'hA24: dout <= 8'b00000000; // 2596 :   0 - 0x0
      13'hA25: dout <= 8'b00000000; // 2597 :   0 - 0x0
      13'hA26: dout <= 8'b01010101; // 2598 :  85 - 0x55
      13'hA27: dout <= 8'b00000000; // 2599 :   0 - 0x0
      13'hA28: dout <= 8'b00010000; // 2600 :  16 - 0x10
      13'hA29: dout <= 8'b00111000; // 2601 :  56 - 0x38
      13'hA2A: dout <= 8'b01111100; // 2602 : 124 - 0x7c
      13'hA2B: dout <= 8'b00000000; // 2603 :   0 - 0x0
      13'hA2C: dout <= 8'b00000000; // 2604 :   0 - 0x0
      13'hA2D: dout <= 8'b00000000; // 2605 :   0 - 0x0
      13'hA2E: dout <= 8'b00000000; // 2606 :   0 - 0x0
      13'hA2F: dout <= 8'b00000000; // 2607 :   0 - 0x0
      13'hA30: dout <= 8'b11110000; // 2608 : 240 - 0xf0 -- Sprite 0xa3
      13'hA31: dout <= 8'b11010010; // 2609 : 210 - 0xd2
      13'hA32: dout <= 8'b10010000; // 2610 : 144 - 0x90
      13'hA33: dout <= 8'b00010010; // 2611 :  18 - 0x12
      13'hA34: dout <= 8'b10010000; // 2612 : 144 - 0x90
      13'hA35: dout <= 8'b11010010; // 2613 : 210 - 0xd2
      13'hA36: dout <= 8'b11110000; // 2614 : 240 - 0xf0
      13'hA37: dout <= 8'b11110010; // 2615 : 242 - 0xf2
      13'hA38: dout <= 8'b00000000; // 2616 :   0 - 0x0
      13'hA39: dout <= 8'b00100000; // 2617 :  32 - 0x20
      13'hA3A: dout <= 8'b01100000; // 2618 :  96 - 0x60
      13'hA3B: dout <= 8'b11100000; // 2619 : 224 - 0xe0
      13'hA3C: dout <= 8'b01100000; // 2620 :  96 - 0x60
      13'hA3D: dout <= 8'b00100000; // 2621 :  32 - 0x20
      13'hA3E: dout <= 8'b00000000; // 2622 :   0 - 0x0
      13'hA3F: dout <= 8'b00000000; // 2623 :   0 - 0x0
      13'hA40: dout <= 8'b11110000; // 2624 : 240 - 0xf0 -- Sprite 0xa4
      13'hA41: dout <= 8'b11010011; // 2625 : 211 - 0xd3
      13'hA42: dout <= 8'b10010100; // 2626 : 148 - 0x94
      13'hA43: dout <= 8'b00011000; // 2627 :  24 - 0x18
      13'hA44: dout <= 8'b10011111; // 2628 : 159 - 0x9f
      13'hA45: dout <= 8'b11011101; // 2629 : 221 - 0xdd
      13'hA46: dout <= 8'b11111010; // 2630 : 250 - 0xfa
      13'hA47: dout <= 8'b11111101; // 2631 : 253 - 0xfd
      13'hA48: dout <= 8'b00000000; // 2632 :   0 - 0x0
      13'hA49: dout <= 8'b00100000; // 2633 :  32 - 0x20
      13'hA4A: dout <= 8'b01100011; // 2634 :  99 - 0x63
      13'hA4B: dout <= 8'b11100111; // 2635 : 231 - 0xe7
      13'hA4C: dout <= 8'b01100000; // 2636 :  96 - 0x60
      13'hA4D: dout <= 8'b00100010; // 2637 :  34 - 0x22
      13'hA4E: dout <= 8'b00000101; // 2638 :   5 - 0x5
      13'hA4F: dout <= 8'b00000010; // 2639 :   2 - 0x2
      13'hA50: dout <= 8'b00000000; // 2640 :   0 - 0x0 -- Sprite 0xa5
      13'hA51: dout <= 8'b11111111; // 2641 : 255 - 0xff
      13'hA52: dout <= 8'b00000000; // 2642 :   0 - 0x0
      13'hA53: dout <= 8'b00000000; // 2643 :   0 - 0x0
      13'hA54: dout <= 8'b11111111; // 2644 : 255 - 0xff
      13'hA55: dout <= 8'b11011101; // 2645 : 221 - 0xdd
      13'hA56: dout <= 8'b11111010; // 2646 : 250 - 0xfa
      13'hA57: dout <= 8'b11111101; // 2647 : 253 - 0xfd
      13'hA58: dout <= 8'b00000000; // 2648 :   0 - 0x0
      13'hA59: dout <= 8'b00000000; // 2649 :   0 - 0x0
      13'hA5A: dout <= 8'b11111111; // 2650 : 255 - 0xff
      13'hA5B: dout <= 8'b11111111; // 2651 : 255 - 0xff
      13'hA5C: dout <= 8'b00000000; // 2652 :   0 - 0x0
      13'hA5D: dout <= 8'b00100010; // 2653 :  34 - 0x22
      13'hA5E: dout <= 8'b00000101; // 2654 :   5 - 0x5
      13'hA5F: dout <= 8'b00000010; // 2655 :   2 - 0x2
      13'hA60: dout <= 8'b11101111; // 2656 : 239 - 0xef -- Sprite 0xa6
      13'hA61: dout <= 8'b11000111; // 2657 : 199 - 0xc7
      13'hA62: dout <= 8'b10000011; // 2658 : 131 - 0x83
      13'hA63: dout <= 8'b11111111; // 2659 : 255 - 0xff
      13'hA64: dout <= 8'b00011111; // 2660 :  31 - 0x1f
      13'hA65: dout <= 8'b00101101; // 2661 :  45 - 0x2d
      13'hA66: dout <= 8'b01001010; // 2662 :  74 - 0x4a
      13'hA67: dout <= 8'b01001101; // 2663 :  77 - 0x4d
      13'hA68: dout <= 8'b00010000; // 2664 :  16 - 0x10
      13'hA69: dout <= 8'b00111000; // 2665 :  56 - 0x38
      13'hA6A: dout <= 8'b01111100; // 2666 : 124 - 0x7c
      13'hA6B: dout <= 8'b00000000; // 2667 :   0 - 0x0
      13'hA6C: dout <= 8'b00000000; // 2668 :   0 - 0x0
      13'hA6D: dout <= 8'b00010010; // 2669 :  18 - 0x12
      13'hA6E: dout <= 8'b00110101; // 2670 :  53 - 0x35
      13'hA6F: dout <= 8'b00110010; // 2671 :  50 - 0x32
      13'hA70: dout <= 8'b01001111; // 2672 :  79 - 0x4f -- Sprite 0xa7
      13'hA71: dout <= 8'b01001111; // 2673 :  79 - 0x4f
      13'hA72: dout <= 8'b01001011; // 2674 :  75 - 0x4b
      13'hA73: dout <= 8'b01001111; // 2675 :  79 - 0x4f
      13'hA74: dout <= 8'b01001111; // 2676 :  79 - 0x4f
      13'hA75: dout <= 8'b01001101; // 2677 :  77 - 0x4d
      13'hA76: dout <= 8'b01001010; // 2678 :  74 - 0x4a
      13'hA77: dout <= 8'b01001101; // 2679 :  77 - 0x4d
      13'hA78: dout <= 8'b00110000; // 2680 :  48 - 0x30
      13'hA79: dout <= 8'b00110000; // 2681 :  48 - 0x30
      13'hA7A: dout <= 8'b00110100; // 2682 :  52 - 0x34
      13'hA7B: dout <= 8'b00110000; // 2683 :  48 - 0x30
      13'hA7C: dout <= 8'b00110000; // 2684 :  48 - 0x30
      13'hA7D: dout <= 8'b00110010; // 2685 :  50 - 0x32
      13'hA7E: dout <= 8'b00110101; // 2686 :  53 - 0x35
      13'hA7F: dout <= 8'b00110010; // 2687 :  50 - 0x32
      13'hA80: dout <= 8'b01001111; // 2688 :  79 - 0x4f -- Sprite 0xa8
      13'hA81: dout <= 8'b11001111; // 2689 : 207 - 0xcf
      13'hA82: dout <= 8'b00001011; // 2690 :  11 - 0xb
      13'hA83: dout <= 8'b00001111; // 2691 :  15 - 0xf
      13'hA84: dout <= 8'b11111111; // 2692 : 255 - 0xff
      13'hA85: dout <= 8'b11011101; // 2693 : 221 - 0xdd
      13'hA86: dout <= 8'b11111010; // 2694 : 250 - 0xfa
      13'hA87: dout <= 8'b11111101; // 2695 : 253 - 0xfd
      13'hA88: dout <= 8'b00110000; // 2696 :  48 - 0x30
      13'hA89: dout <= 8'b00110000; // 2697 :  48 - 0x30
      13'hA8A: dout <= 8'b11110100; // 2698 : 244 - 0xf4
      13'hA8B: dout <= 8'b11110000; // 2699 : 240 - 0xf0
      13'hA8C: dout <= 8'b00000000; // 2700 :   0 - 0x0
      13'hA8D: dout <= 8'b00100010; // 2701 :  34 - 0x22
      13'hA8E: dout <= 8'b00000101; // 2702 :   5 - 0x5
      13'hA8F: dout <= 8'b00000010; // 2703 :   2 - 0x2
      13'hA90: dout <= 8'b11111111; // 2704 : 255 - 0xff -- Sprite 0xa9
      13'hA91: dout <= 8'b11111111; // 2705 : 255 - 0xff
      13'hA92: dout <= 8'b11111111; // 2706 : 255 - 0xff
      13'hA93: dout <= 8'b11111111; // 2707 : 255 - 0xff
      13'hA94: dout <= 8'b11111111; // 2708 : 255 - 0xff
      13'hA95: dout <= 8'b11111111; // 2709 : 255 - 0xff
      13'hA96: dout <= 8'b11111111; // 2710 : 255 - 0xff
      13'hA97: dout <= 8'b11111111; // 2711 : 255 - 0xff
      13'hA98: dout <= 8'b00000000; // 2712 :   0 - 0x0
      13'hA99: dout <= 8'b00000000; // 2713 :   0 - 0x0
      13'hA9A: dout <= 8'b00000000; // 2714 :   0 - 0x0
      13'hA9B: dout <= 8'b00000000; // 2715 :   0 - 0x0
      13'hA9C: dout <= 8'b00000000; // 2716 :   0 - 0x0
      13'hA9D: dout <= 8'b00000000; // 2717 :   0 - 0x0
      13'hA9E: dout <= 8'b00000000; // 2718 :   0 - 0x0
      13'hA9F: dout <= 8'b00000000; // 2719 :   0 - 0x0
      13'hAA0: dout <= 8'b11111111; // 2720 : 255 - 0xff -- Sprite 0xaa
      13'hAA1: dout <= 8'b11111111; // 2721 : 255 - 0xff
      13'hAA2: dout <= 8'b10101111; // 2722 : 175 - 0xaf
      13'hAA3: dout <= 8'b01010111; // 2723 :  87 - 0x57
      13'hAA4: dout <= 8'b10001111; // 2724 : 143 - 0x8f
      13'hAA5: dout <= 8'b11011101; // 2725 : 221 - 0xdd
      13'hAA6: dout <= 8'b11111010; // 2726 : 250 - 0xfa
      13'hAA7: dout <= 8'b11111101; // 2727 : 253 - 0xfd
      13'hAA8: dout <= 8'b00000000; // 2728 :   0 - 0x0
      13'hAA9: dout <= 8'b00000000; // 2729 :   0 - 0x0
      13'hAAA: dout <= 8'b01010000; // 2730 :  80 - 0x50
      13'hAAB: dout <= 8'b10101000; // 2731 : 168 - 0xa8
      13'hAAC: dout <= 8'b01110000; // 2732 : 112 - 0x70
      13'hAAD: dout <= 8'b00100010; // 2733 :  34 - 0x22
      13'hAAE: dout <= 8'b00000101; // 2734 :   5 - 0x5
      13'hAAF: dout <= 8'b00000010; // 2735 :   2 - 0x2
      13'hAB0: dout <= 8'b11111111; // 2736 : 255 - 0xff -- Sprite 0xab
      13'hAB1: dout <= 8'b00000000; // 2737 :   0 - 0x0
      13'hAB2: dout <= 8'b00000000; // 2738 :   0 - 0x0
      13'hAB3: dout <= 8'b00000000; // 2739 :   0 - 0x0
      13'hAB4: dout <= 8'b00000000; // 2740 :   0 - 0x0
      13'hAB5: dout <= 8'b00000000; // 2741 :   0 - 0x0
      13'hAB6: dout <= 8'b00000000; // 2742 :   0 - 0x0
      13'hAB7: dout <= 8'b00000000; // 2743 :   0 - 0x0
      13'hAB8: dout <= 8'b00000000; // 2744 :   0 - 0x0
      13'hAB9: dout <= 8'b00000000; // 2745 :   0 - 0x0
      13'hABA: dout <= 8'b00000000; // 2746 :   0 - 0x0
      13'hABB: dout <= 8'b00000000; // 2747 :   0 - 0x0
      13'hABC: dout <= 8'b00000000; // 2748 :   0 - 0x0
      13'hABD: dout <= 8'b00000000; // 2749 :   0 - 0x0
      13'hABE: dout <= 8'b00000000; // 2750 :   0 - 0x0
      13'hABF: dout <= 8'b00000000; // 2751 :   0 - 0x0
      13'hAC0: dout <= 8'b00000000; // 2752 :   0 - 0x0 -- Sprite 0xac
      13'hAC1: dout <= 8'b00000000; // 2753 :   0 - 0x0
      13'hAC2: dout <= 8'b00000000; // 2754 :   0 - 0x0
      13'hAC3: dout <= 8'b00000000; // 2755 :   0 - 0x0
      13'hAC4: dout <= 8'b00000000; // 2756 :   0 - 0x0
      13'hAC5: dout <= 8'b00000000; // 2757 :   0 - 0x0
      13'hAC6: dout <= 8'b00000000; // 2758 :   0 - 0x0
      13'hAC7: dout <= 8'b00000000; // 2759 :   0 - 0x0
      13'hAC8: dout <= 8'b00000000; // 2760 :   0 - 0x0
      13'hAC9: dout <= 8'b00000000; // 2761 :   0 - 0x0
      13'hACA: dout <= 8'b00000000; // 2762 :   0 - 0x0
      13'hACB: dout <= 8'b00000000; // 2763 :   0 - 0x0
      13'hACC: dout <= 8'b00000000; // 2764 :   0 - 0x0
      13'hACD: dout <= 8'b00000000; // 2765 :   0 - 0x0
      13'hACE: dout <= 8'b00000000; // 2766 :   0 - 0x0
      13'hACF: dout <= 8'b00000000; // 2767 :   0 - 0x0
      13'hAD0: dout <= 8'b00000000; // 2768 :   0 - 0x0 -- Sprite 0xad
      13'hAD1: dout <= 8'b11111111; // 2769 : 255 - 0xff
      13'hAD2: dout <= 8'b00000000; // 2770 :   0 - 0x0
      13'hAD3: dout <= 8'b11111111; // 2771 : 255 - 0xff
      13'hAD4: dout <= 8'b11111111; // 2772 : 255 - 0xff
      13'hAD5: dout <= 8'b11111111; // 2773 : 255 - 0xff
      13'hAD6: dout <= 8'b11111111; // 2774 : 255 - 0xff
      13'hAD7: dout <= 8'b11111111; // 2775 : 255 - 0xff
      13'hAD8: dout <= 8'b00000000; // 2776 :   0 - 0x0
      13'hAD9: dout <= 8'b00000000; // 2777 :   0 - 0x0
      13'hADA: dout <= 8'b11111111; // 2778 : 255 - 0xff
      13'hADB: dout <= 8'b00000000; // 2779 :   0 - 0x0
      13'hADC: dout <= 8'b00000000; // 2780 :   0 - 0x0
      13'hADD: dout <= 8'b00000000; // 2781 :   0 - 0x0
      13'hADE: dout <= 8'b00000000; // 2782 :   0 - 0x0
      13'hADF: dout <= 8'b00000000; // 2783 :   0 - 0x0
      13'hAE0: dout <= 8'b11111111; // 2784 : 255 - 0xff -- Sprite 0xae
      13'hAE1: dout <= 8'b11111111; // 2785 : 255 - 0xff
      13'hAE2: dout <= 8'b11111111; // 2786 : 255 - 0xff
      13'hAE3: dout <= 8'b11111111; // 2787 : 255 - 0xff
      13'hAE4: dout <= 8'b11111111; // 2788 : 255 - 0xff
      13'hAE5: dout <= 8'b00000000; // 2789 :   0 - 0x0
      13'hAE6: dout <= 8'b11111111; // 2790 : 255 - 0xff
      13'hAE7: dout <= 8'b00000000; // 2791 :   0 - 0x0
      13'hAE8: dout <= 8'b00000000; // 2792 :   0 - 0x0
      13'hAE9: dout <= 8'b00000000; // 2793 :   0 - 0x0
      13'hAEA: dout <= 8'b00000000; // 2794 :   0 - 0x0
      13'hAEB: dout <= 8'b00000000; // 2795 :   0 - 0x0
      13'hAEC: dout <= 8'b00000000; // 2796 :   0 - 0x0
      13'hAED: dout <= 8'b11111111; // 2797 : 255 - 0xff
      13'hAEE: dout <= 8'b00000000; // 2798 :   0 - 0x0
      13'hAEF: dout <= 8'b00000000; // 2799 :   0 - 0x0
      13'hAF0: dout <= 8'b11111111; // 2800 : 255 - 0xff -- Sprite 0xaf
      13'hAF1: dout <= 8'b11111111; // 2801 : 255 - 0xff
      13'hAF2: dout <= 8'b11111111; // 2802 : 255 - 0xff
      13'hAF3: dout <= 8'b11111111; // 2803 : 255 - 0xff
      13'hAF4: dout <= 8'b11111111; // 2804 : 255 - 0xff
      13'hAF5: dout <= 8'b11111111; // 2805 : 255 - 0xff
      13'hAF6: dout <= 8'b11111111; // 2806 : 255 - 0xff
      13'hAF7: dout <= 8'b11111111; // 2807 : 255 - 0xff
      13'hAF8: dout <= 8'b00000000; // 2808 :   0 - 0x0
      13'hAF9: dout <= 8'b00000000; // 2809 :   0 - 0x0
      13'hAFA: dout <= 8'b00000000; // 2810 :   0 - 0x0
      13'hAFB: dout <= 8'b00000000; // 2811 :   0 - 0x0
      13'hAFC: dout <= 8'b00000000; // 2812 :   0 - 0x0
      13'hAFD: dout <= 8'b00000000; // 2813 :   0 - 0x0
      13'hAFE: dout <= 8'b00000000; // 2814 :   0 - 0x0
      13'hAFF: dout <= 8'b00000000; // 2815 :   0 - 0x0
      13'hB00: dout <= 8'b00000000; // 2816 :   0 - 0x0 -- Sprite 0xb0
      13'hB01: dout <= 8'b00011111; // 2817 :  31 - 0x1f
      13'hB02: dout <= 8'b00010000; // 2818 :  16 - 0x10
      13'hB03: dout <= 8'b00010000; // 2819 :  16 - 0x10
      13'hB04: dout <= 8'b00010000; // 2820 :  16 - 0x10
      13'hB05: dout <= 8'b00010000; // 2821 :  16 - 0x10
      13'hB06: dout <= 8'b00010000; // 2822 :  16 - 0x10
      13'hB07: dout <= 8'b00010000; // 2823 :  16 - 0x10
      13'hB08: dout <= 8'b00000000; // 2824 :   0 - 0x0
      13'hB09: dout <= 8'b00011111; // 2825 :  31 - 0x1f
      13'hB0A: dout <= 8'b00011111; // 2826 :  31 - 0x1f
      13'hB0B: dout <= 8'b00011111; // 2827 :  31 - 0x1f
      13'hB0C: dout <= 8'b00011111; // 2828 :  31 - 0x1f
      13'hB0D: dout <= 8'b00011111; // 2829 :  31 - 0x1f
      13'hB0E: dout <= 8'b00011111; // 2830 :  31 - 0x1f
      13'hB0F: dout <= 8'b00011111; // 2831 :  31 - 0x1f
      13'hB10: dout <= 8'b00000000; // 2832 :   0 - 0x0 -- Sprite 0xb1
      13'hB11: dout <= 8'b11111000; // 2833 : 248 - 0xf8
      13'hB12: dout <= 8'b00001000; // 2834 :   8 - 0x8
      13'hB13: dout <= 8'b00001000; // 2835 :   8 - 0x8
      13'hB14: dout <= 8'b00001000; // 2836 :   8 - 0x8
      13'hB15: dout <= 8'b00001000; // 2837 :   8 - 0x8
      13'hB16: dout <= 8'b00001000; // 2838 :   8 - 0x8
      13'hB17: dout <= 8'b00001000; // 2839 :   8 - 0x8
      13'hB18: dout <= 8'b00000000; // 2840 :   0 - 0x0
      13'hB19: dout <= 8'b11110000; // 2841 : 240 - 0xf0
      13'hB1A: dout <= 8'b11110000; // 2842 : 240 - 0xf0
      13'hB1B: dout <= 8'b11110000; // 2843 : 240 - 0xf0
      13'hB1C: dout <= 8'b11110000; // 2844 : 240 - 0xf0
      13'hB1D: dout <= 8'b11110000; // 2845 : 240 - 0xf0
      13'hB1E: dout <= 8'b11110000; // 2846 : 240 - 0xf0
      13'hB1F: dout <= 8'b11110000; // 2847 : 240 - 0xf0
      13'hB20: dout <= 8'b00010000; // 2848 :  16 - 0x10 -- Sprite 0xb2
      13'hB21: dout <= 8'b00010000; // 2849 :  16 - 0x10
      13'hB22: dout <= 8'b00010000; // 2850 :  16 - 0x10
      13'hB23: dout <= 8'b00010000; // 2851 :  16 - 0x10
      13'hB24: dout <= 8'b00011111; // 2852 :  31 - 0x1f
      13'hB25: dout <= 8'b00011111; // 2853 :  31 - 0x1f
      13'hB26: dout <= 8'b00001111; // 2854 :  15 - 0xf
      13'hB27: dout <= 8'b00000000; // 2855 :   0 - 0x0
      13'hB28: dout <= 8'b00011111; // 2856 :  31 - 0x1f
      13'hB29: dout <= 8'b00011111; // 2857 :  31 - 0x1f
      13'hB2A: dout <= 8'b00011111; // 2858 :  31 - 0x1f
      13'hB2B: dout <= 8'b00011111; // 2859 :  31 - 0x1f
      13'hB2C: dout <= 8'b00000000; // 2860 :   0 - 0x0
      13'hB2D: dout <= 8'b00000000; // 2861 :   0 - 0x0
      13'hB2E: dout <= 8'b00000000; // 2862 :   0 - 0x0
      13'hB2F: dout <= 8'b00000000; // 2863 :   0 - 0x0
      13'hB30: dout <= 8'b00001000; // 2864 :   8 - 0x8 -- Sprite 0xb3
      13'hB31: dout <= 8'b00001000; // 2865 :   8 - 0x8
      13'hB32: dout <= 8'b00001000; // 2866 :   8 - 0x8
      13'hB33: dout <= 8'b00001000; // 2867 :   8 - 0x8
      13'hB34: dout <= 8'b11111000; // 2868 : 248 - 0xf8
      13'hB35: dout <= 8'b11111000; // 2869 : 248 - 0xf8
      13'hB36: dout <= 8'b11110000; // 2870 : 240 - 0xf0
      13'hB37: dout <= 8'b00000000; // 2871 :   0 - 0x0
      13'hB38: dout <= 8'b11110000; // 2872 : 240 - 0xf0
      13'hB39: dout <= 8'b11110000; // 2873 : 240 - 0xf0
      13'hB3A: dout <= 8'b11110000; // 2874 : 240 - 0xf0
      13'hB3B: dout <= 8'b11110000; // 2875 : 240 - 0xf0
      13'hB3C: dout <= 8'b00000000; // 2876 :   0 - 0x0
      13'hB3D: dout <= 8'b00000000; // 2877 :   0 - 0x0
      13'hB3E: dout <= 8'b00000000; // 2878 :   0 - 0x0
      13'hB3F: dout <= 8'b00000000; // 2879 :   0 - 0x0
      13'hB40: dout <= 8'b00000000; // 2880 :   0 - 0x0 -- Sprite 0xb4
      13'hB41: dout <= 8'b00000000; // 2881 :   0 - 0x0
      13'hB42: dout <= 8'b00111111; // 2882 :  63 - 0x3f
      13'hB43: dout <= 8'b01100000; // 2883 :  96 - 0x60
      13'hB44: dout <= 8'b01100000; // 2884 :  96 - 0x60
      13'hB45: dout <= 8'b01100000; // 2885 :  96 - 0x60
      13'hB46: dout <= 8'b01100000; // 2886 :  96 - 0x60
      13'hB47: dout <= 8'b01100000; // 2887 :  96 - 0x60
      13'hB48: dout <= 8'b00000000; // 2888 :   0 - 0x0
      13'hB49: dout <= 8'b00000000; // 2889 :   0 - 0x0
      13'hB4A: dout <= 8'b00111111; // 2890 :  63 - 0x3f
      13'hB4B: dout <= 8'b01111111; // 2891 : 127 - 0x7f
      13'hB4C: dout <= 8'b01111111; // 2892 : 127 - 0x7f
      13'hB4D: dout <= 8'b01111111; // 2893 : 127 - 0x7f
      13'hB4E: dout <= 8'b01111111; // 2894 : 127 - 0x7f
      13'hB4F: dout <= 8'b01111111; // 2895 : 127 - 0x7f
      13'hB50: dout <= 8'b00000000; // 2896 :   0 - 0x0 -- Sprite 0xb5
      13'hB51: dout <= 8'b00000000; // 2897 :   0 - 0x0
      13'hB52: dout <= 8'b11111100; // 2898 : 252 - 0xfc
      13'hB53: dout <= 8'b00000110; // 2899 :   6 - 0x6
      13'hB54: dout <= 8'b00000110; // 2900 :   6 - 0x6
      13'hB55: dout <= 8'b00000110; // 2901 :   6 - 0x6
      13'hB56: dout <= 8'b00000110; // 2902 :   6 - 0x6
      13'hB57: dout <= 8'b00000110; // 2903 :   6 - 0x6
      13'hB58: dout <= 8'b00000000; // 2904 :   0 - 0x0
      13'hB59: dout <= 8'b00000000; // 2905 :   0 - 0x0
      13'hB5A: dout <= 8'b11111000; // 2906 : 248 - 0xf8
      13'hB5B: dout <= 8'b11111000; // 2907 : 248 - 0xf8
      13'hB5C: dout <= 8'b11111000; // 2908 : 248 - 0xf8
      13'hB5D: dout <= 8'b11111000; // 2909 : 248 - 0xf8
      13'hB5E: dout <= 8'b11111000; // 2910 : 248 - 0xf8
      13'hB5F: dout <= 8'b11111000; // 2911 : 248 - 0xf8
      13'hB60: dout <= 8'b01100000; // 2912 :  96 - 0x60 -- Sprite 0xb6
      13'hB61: dout <= 8'b01100000; // 2913 :  96 - 0x60
      13'hB62: dout <= 8'b01100000; // 2914 :  96 - 0x60
      13'hB63: dout <= 8'b01111111; // 2915 : 127 - 0x7f
      13'hB64: dout <= 8'b01111111; // 2916 : 127 - 0x7f
      13'hB65: dout <= 8'b00111111; // 2917 :  63 - 0x3f
      13'hB66: dout <= 8'b00000000; // 2918 :   0 - 0x0
      13'hB67: dout <= 8'b00000000; // 2919 :   0 - 0x0
      13'hB68: dout <= 8'b01111111; // 2920 : 127 - 0x7f
      13'hB69: dout <= 8'b01111111; // 2921 : 127 - 0x7f
      13'hB6A: dout <= 8'b01111111; // 2922 : 127 - 0x7f
      13'hB6B: dout <= 8'b01000000; // 2923 :  64 - 0x40
      13'hB6C: dout <= 8'b00000000; // 2924 :   0 - 0x0
      13'hB6D: dout <= 8'b00000000; // 2925 :   0 - 0x0
      13'hB6E: dout <= 8'b00000000; // 2926 :   0 - 0x0
      13'hB6F: dout <= 8'b00000000; // 2927 :   0 - 0x0
      13'hB70: dout <= 8'b00000110; // 2928 :   6 - 0x6 -- Sprite 0xb7
      13'hB71: dout <= 8'b00000110; // 2929 :   6 - 0x6
      13'hB72: dout <= 8'b00000110; // 2930 :   6 - 0x6
      13'hB73: dout <= 8'b11111110; // 2931 : 254 - 0xfe
      13'hB74: dout <= 8'b11111110; // 2932 : 254 - 0xfe
      13'hB75: dout <= 8'b11111100; // 2933 : 252 - 0xfc
      13'hB76: dout <= 8'b00000000; // 2934 :   0 - 0x0
      13'hB77: dout <= 8'b00000000; // 2935 :   0 - 0x0
      13'hB78: dout <= 8'b11111000; // 2936 : 248 - 0xf8
      13'hB79: dout <= 8'b11111000; // 2937 : 248 - 0xf8
      13'hB7A: dout <= 8'b11111000; // 2938 : 248 - 0xf8
      13'hB7B: dout <= 8'b00000000; // 2939 :   0 - 0x0
      13'hB7C: dout <= 8'b00000000; // 2940 :   0 - 0x0
      13'hB7D: dout <= 8'b00000000; // 2941 :   0 - 0x0
      13'hB7E: dout <= 8'b00000000; // 2942 :   0 - 0x0
      13'hB7F: dout <= 8'b00000000; // 2943 :   0 - 0x0
      13'hB80: dout <= 8'b01100000; // 2944 :  96 - 0x60 -- Sprite 0xb8
      13'hB81: dout <= 8'b11110011; // 2945 : 243 - 0xf3
      13'hB82: dout <= 8'b11000111; // 2946 : 199 - 0xc7
      13'hB83: dout <= 8'b10000110; // 2947 : 134 - 0x86
      13'hB84: dout <= 8'b00000100; // 2948 :   4 - 0x4
      13'hB85: dout <= 8'b00000100; // 2949 :   4 - 0x4
      13'hB86: dout <= 8'b00000111; // 2950 :   7 - 0x7
      13'hB87: dout <= 8'b00000111; // 2951 :   7 - 0x7
      13'hB88: dout <= 8'b00000000; // 2952 :   0 - 0x0
      13'hB89: dout <= 8'b00000011; // 2953 :   3 - 0x3
      13'hB8A: dout <= 8'b00000111; // 2954 :   7 - 0x7
      13'hB8B: dout <= 8'b00000111; // 2955 :   7 - 0x7
      13'hB8C: dout <= 8'b00000111; // 2956 :   7 - 0x7
      13'hB8D: dout <= 8'b00000011; // 2957 :   3 - 0x3
      13'hB8E: dout <= 8'b00000000; // 2958 :   0 - 0x0
      13'hB8F: dout <= 8'b00000000; // 2959 :   0 - 0x0
      13'hB90: dout <= 8'b00000110; // 2960 :   6 - 0x6 -- Sprite 0xb9
      13'hB91: dout <= 8'b10001111; // 2961 : 143 - 0x8f
      13'hB92: dout <= 8'b11000101; // 2962 : 197 - 0xc5
      13'hB93: dout <= 8'b00100011; // 2963 :  35 - 0x23
      13'hB94: dout <= 8'b00101110; // 2964 :  46 - 0x2e
      13'hB95: dout <= 8'b01100000; // 2965 :  96 - 0x60
      13'hB96: dout <= 8'b11100001; // 2966 : 225 - 0xe1
      13'hB97: dout <= 8'b11100001; // 2967 : 225 - 0xe1
      13'hB98: dout <= 8'b00000000; // 2968 :   0 - 0x0
      13'hB99: dout <= 8'b11000001; // 2969 : 193 - 0xc1
      13'hB9A: dout <= 8'b11100010; // 2970 : 226 - 0xe2
      13'hB9B: dout <= 8'b11001100; // 2971 : 204 - 0xcc
      13'hB9C: dout <= 8'b11000000; // 2972 : 192 - 0xc0
      13'hB9D: dout <= 8'b10000000; // 2973 : 128 - 0x80
      13'hB9E: dout <= 8'b00000001; // 2974 :   1 - 0x1
      13'hB9F: dout <= 8'b00000010; // 2975 :   2 - 0x2
      13'hBA0: dout <= 8'b11001000; // 2976 : 200 - 0xc8 -- Sprite 0xba
      13'hBA1: dout <= 8'b11111000; // 2977 : 248 - 0xf8
      13'hBA2: dout <= 8'b10110000; // 2978 : 176 - 0xb0
      13'hBA3: dout <= 8'b00010000; // 2979 :  16 - 0x10
      13'hBA4: dout <= 8'b00110000; // 2980 :  48 - 0x30
      13'hBA5: dout <= 8'b11001000; // 2981 : 200 - 0xc8
      13'hBA6: dout <= 8'b11111000; // 2982 : 248 - 0xf8
      13'hBA7: dout <= 8'b10000000; // 2983 : 128 - 0x80
      13'hBA8: dout <= 8'b11110000; // 2984 : 240 - 0xf0
      13'hBA9: dout <= 8'b00000000; // 2985 :   0 - 0x0
      13'hBAA: dout <= 8'b00100000; // 2986 :  32 - 0x20
      13'hBAB: dout <= 8'b00100000; // 2987 :  32 - 0x20
      13'hBAC: dout <= 8'b00000000; // 2988 :   0 - 0x0
      13'hBAD: dout <= 8'b11110000; // 2989 : 240 - 0xf0
      13'hBAE: dout <= 8'b00000000; // 2990 :   0 - 0x0
      13'hBAF: dout <= 8'b00000000; // 2991 :   0 - 0x0
      13'hBB0: dout <= 8'b00000011; // 2992 :   3 - 0x3 -- Sprite 0xbb
      13'hBB1: dout <= 8'b00000000; // 2993 :   0 - 0x0
      13'hBB2: dout <= 8'b00000000; // 2994 :   0 - 0x0
      13'hBB3: dout <= 8'b01100000; // 2995 :  96 - 0x60
      13'hBB4: dout <= 8'b11110000; // 2996 : 240 - 0xf0
      13'hBB5: dout <= 8'b11010000; // 2997 : 208 - 0xd0
      13'hBB6: dout <= 8'b10010000; // 2998 : 144 - 0x90
      13'hBB7: dout <= 8'b01100000; // 2999 :  96 - 0x60
      13'hBB8: dout <= 8'b00000000; // 3000 :   0 - 0x0
      13'hBB9: dout <= 8'b00000000; // 3001 :   0 - 0x0
      13'hBBA: dout <= 8'b00000000; // 3002 :   0 - 0x0
      13'hBBB: dout <= 8'b00000000; // 3003 :   0 - 0x0
      13'hBBC: dout <= 8'b00000000; // 3004 :   0 - 0x0
      13'hBBD: dout <= 8'b01100000; // 3005 :  96 - 0x60
      13'hBBE: dout <= 8'b01100000; // 3006 :  96 - 0x60
      13'hBBF: dout <= 8'b00000000; // 3007 :   0 - 0x0
      13'hBC0: dout <= 8'b11000011; // 3008 : 195 - 0xc3 -- Sprite 0xbc
      13'hBC1: dout <= 8'b00001110; // 3009 :  14 - 0xe
      13'hBC2: dout <= 8'b00000000; // 3010 :   0 - 0x0
      13'hBC3: dout <= 8'b00000110; // 3011 :   6 - 0x6
      13'hBC4: dout <= 8'b00001111; // 3012 :  15 - 0xf
      13'hBC5: dout <= 8'b00001101; // 3013 :  13 - 0xd
      13'hBC6: dout <= 8'b00001001; // 3014 :   9 - 0x9
      13'hBC7: dout <= 8'b00000110; // 3015 :   6 - 0x6
      13'hBC8: dout <= 8'b00001100; // 3016 :  12 - 0xc
      13'hBC9: dout <= 8'b00000000; // 3017 :   0 - 0x0
      13'hBCA: dout <= 8'b00000000; // 3018 :   0 - 0x0
      13'hBCB: dout <= 8'b00000000; // 3019 :   0 - 0x0
      13'hBCC: dout <= 8'b00000000; // 3020 :   0 - 0x0
      13'hBCD: dout <= 8'b00000110; // 3021 :   6 - 0x6
      13'hBCE: dout <= 8'b00000110; // 3022 :   6 - 0x6
      13'hBCF: dout <= 8'b00000000; // 3023 :   0 - 0x0
      13'hBD0: dout <= 8'b11100000; // 3024 : 224 - 0xe0 -- Sprite 0xbd
      13'hBD1: dout <= 8'b01100011; // 3025 :  99 - 0x63
      13'hBD2: dout <= 8'b11100111; // 3026 : 231 - 0xe7
      13'hBD3: dout <= 8'b11100110; // 3027 : 230 - 0xe6
      13'hBD4: dout <= 8'b00000100; // 3028 :   4 - 0x4
      13'hBD5: dout <= 8'b00000100; // 3029 :   4 - 0x4
      13'hBD6: dout <= 8'b00000111; // 3030 :   7 - 0x7
      13'hBD7: dout <= 8'b00000111; // 3031 :   7 - 0x7
      13'hBD8: dout <= 8'b00000000; // 3032 :   0 - 0x0
      13'hBD9: dout <= 8'b10000011; // 3033 : 131 - 0x83
      13'hBDA: dout <= 8'b00000111; // 3034 :   7 - 0x7
      13'hBDB: dout <= 8'b00000111; // 3035 :   7 - 0x7
      13'hBDC: dout <= 8'b00000111; // 3036 :   7 - 0x7
      13'hBDD: dout <= 8'b00000011; // 3037 :   3 - 0x3
      13'hBDE: dout <= 8'b00000000; // 3038 :   0 - 0x0
      13'hBDF: dout <= 8'b00000000; // 3039 :   0 - 0x0
      13'hBE0: dout <= 8'b00000111; // 3040 :   7 - 0x7 -- Sprite 0xbe
      13'hBE1: dout <= 8'b10000011; // 3041 : 131 - 0x83
      13'hBE2: dout <= 8'b11000111; // 3042 : 199 - 0xc7
      13'hBE3: dout <= 8'b00100111; // 3043 :  39 - 0x27
      13'hBE4: dout <= 8'b00100000; // 3044 :  32 - 0x20
      13'hBE5: dout <= 8'b01100000; // 3045 :  96 - 0x60
      13'hBE6: dout <= 8'b11100000; // 3046 : 224 - 0xe0
      13'hBE7: dout <= 8'b11100000; // 3047 : 224 - 0xe0
      13'hBE8: dout <= 8'b00000000; // 3048 :   0 - 0x0
      13'hBE9: dout <= 8'b11000100; // 3049 : 196 - 0xc4
      13'hBEA: dout <= 8'b11100000; // 3050 : 224 - 0xe0
      13'hBEB: dout <= 8'b11000000; // 3051 : 192 - 0xc0
      13'hBEC: dout <= 8'b11000000; // 3052 : 192 - 0xc0
      13'hBED: dout <= 8'b10000000; // 3053 : 128 - 0x80
      13'hBEE: dout <= 8'b00000000; // 3054 :   0 - 0x0
      13'hBEF: dout <= 8'b00000000; // 3055 :   0 - 0x0
      13'hBF0: dout <= 8'b00000011; // 3056 :   3 - 0x3 -- Sprite 0xbf
      13'hBF1: dout <= 8'b00000000; // 3057 :   0 - 0x0
      13'hBF2: dout <= 8'b00001100; // 3058 :  12 - 0xc
      13'hBF3: dout <= 8'b00001100; // 3059 :  12 - 0xc
      13'hBF4: dout <= 8'b11100100; // 3060 : 228 - 0xe4
      13'hBF5: dout <= 8'b01101100; // 3061 : 108 - 0x6c
      13'hBF6: dout <= 8'b11101101; // 3062 : 237 - 0xed
      13'hBF7: dout <= 8'b11100111; // 3063 : 231 - 0xe7
      13'hBF8: dout <= 8'b00000000; // 3064 :   0 - 0x0
      13'hBF9: dout <= 8'b00000000; // 3065 :   0 - 0x0
      13'hBFA: dout <= 8'b00000000; // 3066 :   0 - 0x0
      13'hBFB: dout <= 8'b00000000; // 3067 :   0 - 0x0
      13'hBFC: dout <= 8'b00001000; // 3068 :   8 - 0x8
      13'hBFD: dout <= 8'b10001000; // 3069 : 136 - 0x88
      13'hBFE: dout <= 8'b00001011; // 3070 :  11 - 0xb
      13'hBFF: dout <= 8'b00001000; // 3071 :   8 - 0x8
      13'hC00: dout <= 8'b11000000; // 3072 : 192 - 0xc0 -- Sprite 0xc0
      13'hC01: dout <= 8'b00000000; // 3073 :   0 - 0x0
      13'hC02: dout <= 8'b00110000; // 3074 :  48 - 0x30
      13'hC03: dout <= 8'b00110000; // 3075 :  48 - 0x30
      13'hC04: dout <= 8'b00010111; // 3076 :  23 - 0x17
      13'hC05: dout <= 8'b00110011; // 3077 :  51 - 0x33
      13'hC06: dout <= 8'b01110111; // 3078 : 119 - 0x77
      13'hC07: dout <= 8'b11010111; // 3079 : 215 - 0xd7
      13'hC08: dout <= 8'b00000000; // 3080 :   0 - 0x0
      13'hC09: dout <= 8'b00000000; // 3081 :   0 - 0x0
      13'hC0A: dout <= 8'b00000000; // 3082 :   0 - 0x0
      13'hC0B: dout <= 8'b00000000; // 3083 :   0 - 0x0
      13'hC0C: dout <= 8'b00100000; // 3084 :  32 - 0x20
      13'hC0D: dout <= 8'b00100100; // 3085 :  36 - 0x24
      13'hC0E: dout <= 8'b10100000; // 3086 : 160 - 0xa0
      13'hC0F: dout <= 8'b00100000; // 3087 :  32 - 0x20
      13'hC10: dout <= 8'b00001100; // 3088 :  12 - 0xc -- Sprite 0xc1
      13'hC11: dout <= 8'b00000000; // 3089 :   0 - 0x0
      13'hC12: dout <= 8'b00000000; // 3090 :   0 - 0x0
      13'hC13: dout <= 8'b00000000; // 3091 :   0 - 0x0
      13'hC14: dout <= 8'b00000000; // 3092 :   0 - 0x0
      13'hC15: dout <= 8'b00000000; // 3093 :   0 - 0x0
      13'hC16: dout <= 8'b00000000; // 3094 :   0 - 0x0
      13'hC17: dout <= 8'b00000000; // 3095 :   0 - 0x0
      13'hC18: dout <= 8'b00000000; // 3096 :   0 - 0x0
      13'hC19: dout <= 8'b00000000; // 3097 :   0 - 0x0
      13'hC1A: dout <= 8'b00000000; // 3098 :   0 - 0x0
      13'hC1B: dout <= 8'b00000000; // 3099 :   0 - 0x0
      13'hC1C: dout <= 8'b00000000; // 3100 :   0 - 0x0
      13'hC1D: dout <= 8'b00000000; // 3101 :   0 - 0x0
      13'hC1E: dout <= 8'b00000000; // 3102 :   0 - 0x0
      13'hC1F: dout <= 8'b00000000; // 3103 :   0 - 0x0
      13'hC20: dout <= 8'b00110000; // 3104 :  48 - 0x30 -- Sprite 0xc2
      13'hC21: dout <= 8'b00000000; // 3105 :   0 - 0x0
      13'hC22: dout <= 8'b00000000; // 3106 :   0 - 0x0
      13'hC23: dout <= 8'b00000000; // 3107 :   0 - 0x0
      13'hC24: dout <= 8'b00000000; // 3108 :   0 - 0x0
      13'hC25: dout <= 8'b00000000; // 3109 :   0 - 0x0
      13'hC26: dout <= 8'b00000000; // 3110 :   0 - 0x0
      13'hC27: dout <= 8'b00000000; // 3111 :   0 - 0x0
      13'hC28: dout <= 8'b00000000; // 3112 :   0 - 0x0
      13'hC29: dout <= 8'b00000000; // 3113 :   0 - 0x0
      13'hC2A: dout <= 8'b00000000; // 3114 :   0 - 0x0
      13'hC2B: dout <= 8'b00000000; // 3115 :   0 - 0x0
      13'hC2C: dout <= 8'b00000000; // 3116 :   0 - 0x0
      13'hC2D: dout <= 8'b00000000; // 3117 :   0 - 0x0
      13'hC2E: dout <= 8'b00000000; // 3118 :   0 - 0x0
      13'hC2F: dout <= 8'b00000000; // 3119 :   0 - 0x0
      13'hC30: dout <= 8'b00000000; // 3120 :   0 - 0x0 -- Sprite 0xc3
      13'hC31: dout <= 8'b00000000; // 3121 :   0 - 0x0
      13'hC32: dout <= 8'b00000100; // 3122 :   4 - 0x4
      13'hC33: dout <= 8'b00001101; // 3123 :  13 - 0xd
      13'hC34: dout <= 8'b00001111; // 3124 :  15 - 0xf
      13'hC35: dout <= 8'b00001100; // 3125 :  12 - 0xc
      13'hC36: dout <= 8'b00001100; // 3126 :  12 - 0xc
      13'hC37: dout <= 8'b00000100; // 3127 :   4 - 0x4
      13'hC38: dout <= 8'b00000000; // 3128 :   0 - 0x0
      13'hC39: dout <= 8'b00000000; // 3129 :   0 - 0x0
      13'hC3A: dout <= 8'b00001000; // 3130 :   8 - 0x8
      13'hC3B: dout <= 8'b00001011; // 3131 :  11 - 0xb
      13'hC3C: dout <= 8'b00001000; // 3132 :   8 - 0x8
      13'hC3D: dout <= 8'b00001000; // 3133 :   8 - 0x8
      13'hC3E: dout <= 8'b00001000; // 3134 :   8 - 0x8
      13'hC3F: dout <= 8'b00001000; // 3135 :   8 - 0x8
      13'hC40: dout <= 8'b00000000; // 3136 :   0 - 0x0 -- Sprite 0xc4
      13'hC41: dout <= 8'b00000000; // 3137 :   0 - 0x0
      13'hC42: dout <= 8'b00010000; // 3138 :  16 - 0x10
      13'hC43: dout <= 8'b01110000; // 3139 : 112 - 0x70
      13'hC44: dout <= 8'b11110000; // 3140 : 240 - 0xf0
      13'hC45: dout <= 8'b00110000; // 3141 :  48 - 0x30
      13'hC46: dout <= 8'b00110000; // 3142 :  48 - 0x30
      13'hC47: dout <= 8'b00010000; // 3143 :  16 - 0x10
      13'hC48: dout <= 8'b00000000; // 3144 :   0 - 0x0
      13'hC49: dout <= 8'b00000000; // 3145 :   0 - 0x0
      13'hC4A: dout <= 8'b00100000; // 3146 :  32 - 0x20
      13'hC4B: dout <= 8'b10100000; // 3147 : 160 - 0xa0
      13'hC4C: dout <= 8'b00100000; // 3148 :  32 - 0x20
      13'hC4D: dout <= 8'b00100000; // 3149 :  32 - 0x20
      13'hC4E: dout <= 8'b00100000; // 3150 :  32 - 0x20
      13'hC4F: dout <= 8'b00100000; // 3151 :  32 - 0x20
      13'hC50: dout <= 8'b11100100; // 3152 : 228 - 0xe4 -- Sprite 0xc5
      13'hC51: dout <= 8'b00100100; // 3153 :  36 - 0x24
      13'hC52: dout <= 8'b11101111; // 3154 : 239 - 0xef
      13'hC53: dout <= 8'b11100111; // 3155 : 231 - 0xe7
      13'hC54: dout <= 8'b00000110; // 3156 :   6 - 0x6
      13'hC55: dout <= 8'b00000100; // 3157 :   4 - 0x4
      13'hC56: dout <= 8'b00000100; // 3158 :   4 - 0x4
      13'hC57: dout <= 8'b00000111; // 3159 :   7 - 0x7
      13'hC58: dout <= 8'b00001000; // 3160 :   8 - 0x8
      13'hC59: dout <= 8'b11001000; // 3161 : 200 - 0xc8
      13'hC5A: dout <= 8'b00000011; // 3162 :   3 - 0x3
      13'hC5B: dout <= 8'b00000111; // 3163 :   7 - 0x7
      13'hC5C: dout <= 8'b00000111; // 3164 :   7 - 0x7
      13'hC5D: dout <= 8'b00000111; // 3165 :   7 - 0x7
      13'hC5E: dout <= 8'b00000011; // 3166 :   3 - 0x3
      13'hC5F: dout <= 8'b00000000; // 3167 :   0 - 0x0
      13'hC60: dout <= 8'b00010111; // 3168 :  23 - 0x17 -- Sprite 0xc6
      13'hC61: dout <= 8'b00010001; // 3169 :  17 - 0x11
      13'hC62: dout <= 8'b10110111; // 3170 : 183 - 0xb7
      13'hC63: dout <= 8'b11000111; // 3171 : 199 - 0xc7
      13'hC64: dout <= 8'b00100000; // 3172 :  32 - 0x20
      13'hC65: dout <= 8'b00100000; // 3173 :  32 - 0x20
      13'hC66: dout <= 8'b01100000; // 3174 :  96 - 0x60
      13'hC67: dout <= 8'b11100000; // 3175 : 224 - 0xe0
      13'hC68: dout <= 8'b00100000; // 3176 :  32 - 0x20
      13'hC69: dout <= 8'b00100110; // 3177 :  38 - 0x26
      13'hC6A: dout <= 8'b11000000; // 3178 : 192 - 0xc0
      13'hC6B: dout <= 8'b11100000; // 3179 : 224 - 0xe0
      13'hC6C: dout <= 8'b11000000; // 3180 : 192 - 0xc0
      13'hC6D: dout <= 8'b11000000; // 3181 : 192 - 0xc0
      13'hC6E: dout <= 8'b10000000; // 3182 : 128 - 0x80
      13'hC6F: dout <= 8'b00000000; // 3183 :   0 - 0x0
      13'hC70: dout <= 8'b00000111; // 3184 :   7 - 0x7 -- Sprite 0xc7
      13'hC71: dout <= 8'b00000011; // 3185 :   3 - 0x3
      13'hC72: dout <= 8'b00000000; // 3186 :   0 - 0x0
      13'hC73: dout <= 8'b00000000; // 3187 :   0 - 0x0
      13'hC74: dout <= 8'b11100000; // 3188 : 224 - 0xe0
      13'hC75: dout <= 8'b00100000; // 3189 :  32 - 0x20
      13'hC76: dout <= 8'b11100000; // 3190 : 224 - 0xe0
      13'hC77: dout <= 8'b11100000; // 3191 : 224 - 0xe0
      13'hC78: dout <= 8'b00000000; // 3192 :   0 - 0x0
      13'hC79: dout <= 8'b00000000; // 3193 :   0 - 0x0
      13'hC7A: dout <= 8'b00000000; // 3194 :   0 - 0x0
      13'hC7B: dout <= 8'b00000000; // 3195 :   0 - 0x0
      13'hC7C: dout <= 8'b00000000; // 3196 :   0 - 0x0
      13'hC7D: dout <= 8'b11000000; // 3197 : 192 - 0xc0
      13'hC7E: dout <= 8'b00000000; // 3198 :   0 - 0x0
      13'hC7F: dout <= 8'b00000000; // 3199 :   0 - 0x0
      13'hC80: dout <= 8'b11100000; // 3200 : 224 - 0xe0 -- Sprite 0xc8
      13'hC81: dout <= 8'b11000000; // 3201 : 192 - 0xc0
      13'hC82: dout <= 8'b00000000; // 3202 :   0 - 0x0
      13'hC83: dout <= 8'b00000000; // 3203 :   0 - 0x0
      13'hC84: dout <= 8'b00000111; // 3204 :   7 - 0x7
      13'hC85: dout <= 8'b00000001; // 3205 :   1 - 0x1
      13'hC86: dout <= 8'b00000111; // 3206 :   7 - 0x7
      13'hC87: dout <= 8'b00000111; // 3207 :   7 - 0x7
      13'hC88: dout <= 8'b00000000; // 3208 :   0 - 0x0
      13'hC89: dout <= 8'b00000000; // 3209 :   0 - 0x0
      13'hC8A: dout <= 8'b00000000; // 3210 :   0 - 0x0
      13'hC8B: dout <= 8'b00000000; // 3211 :   0 - 0x0
      13'hC8C: dout <= 8'b00000000; // 3212 :   0 - 0x0
      13'hC8D: dout <= 8'b00000110; // 3213 :   6 - 0x6
      13'hC8E: dout <= 8'b00000000; // 3214 :   0 - 0x0
      13'hC8F: dout <= 8'b00000000; // 3215 :   0 - 0x0
      13'hC90: dout <= 8'b00010011; // 3216 :  19 - 0x13 -- Sprite 0xc9
      13'hC91: dout <= 8'b00011111; // 3217 :  31 - 0x1f
      13'hC92: dout <= 8'b00001101; // 3218 :  13 - 0xd
      13'hC93: dout <= 8'b00000100; // 3219 :   4 - 0x4
      13'hC94: dout <= 8'b00001100; // 3220 :  12 - 0xc
      13'hC95: dout <= 8'b00010011; // 3221 :  19 - 0x13
      13'hC96: dout <= 8'b00011111; // 3222 :  31 - 0x1f
      13'hC97: dout <= 8'b00000001; // 3223 :   1 - 0x1
      13'hC98: dout <= 8'b00001111; // 3224 :  15 - 0xf
      13'hC99: dout <= 8'b00000000; // 3225 :   0 - 0x0
      13'hC9A: dout <= 8'b00001000; // 3226 :   8 - 0x8
      13'hC9B: dout <= 8'b00001000; // 3227 :   8 - 0x8
      13'hC9C: dout <= 8'b00000000; // 3228 :   0 - 0x0
      13'hC9D: dout <= 8'b00001111; // 3229 :  15 - 0xf
      13'hC9E: dout <= 8'b00000000; // 3230 :   0 - 0x0
      13'hC9F: dout <= 8'b00000000; // 3231 :   0 - 0x0
      13'hCA0: dout <= 8'b01100000; // 3232 :  96 - 0x60 -- Sprite 0xca
      13'hCA1: dout <= 8'b11110011; // 3233 : 243 - 0xf3
      13'hCA2: dout <= 8'b10100111; // 3234 : 167 - 0xa7
      13'hCA3: dout <= 8'b11000110; // 3235 : 198 - 0xc6
      13'hCA4: dout <= 8'b01110100; // 3236 : 116 - 0x74
      13'hCA5: dout <= 8'b00000100; // 3237 :   4 - 0x4
      13'hCA6: dout <= 8'b10000111; // 3238 : 135 - 0x87
      13'hCA7: dout <= 8'b10000111; // 3239 : 135 - 0x87
      13'hCA8: dout <= 8'b00000000; // 3240 :   0 - 0x0
      13'hCA9: dout <= 8'b10000011; // 3241 : 131 - 0x83
      13'hCAA: dout <= 8'b01000111; // 3242 :  71 - 0x47
      13'hCAB: dout <= 8'b00110111; // 3243 :  55 - 0x37
      13'hCAC: dout <= 8'b00000111; // 3244 :   7 - 0x7
      13'hCAD: dout <= 8'b00000011; // 3245 :   3 - 0x3
      13'hCAE: dout <= 8'b10000000; // 3246 : 128 - 0x80
      13'hCAF: dout <= 8'b01000000; // 3247 :  64 - 0x40
      13'hCB0: dout <= 8'b00000110; // 3248 :   6 - 0x6 -- Sprite 0xcb
      13'hCB1: dout <= 8'b10001111; // 3249 : 143 - 0x8f
      13'hCB2: dout <= 8'b11000011; // 3250 : 195 - 0xc3
      13'hCB3: dout <= 8'b00100001; // 3251 :  33 - 0x21
      13'hCB4: dout <= 8'b00100000; // 3252 :  32 - 0x20
      13'hCB5: dout <= 8'b01100000; // 3253 :  96 - 0x60
      13'hCB6: dout <= 8'b11100000; // 3254 : 224 - 0xe0
      13'hCB7: dout <= 8'b11100000; // 3255 : 224 - 0xe0
      13'hCB8: dout <= 8'b00000000; // 3256 :   0 - 0x0
      13'hCB9: dout <= 8'b11000000; // 3257 : 192 - 0xc0
      13'hCBA: dout <= 8'b11100000; // 3258 : 224 - 0xe0
      13'hCBB: dout <= 8'b11000000; // 3259 : 192 - 0xc0
      13'hCBC: dout <= 8'b11000000; // 3260 : 192 - 0xc0
      13'hCBD: dout <= 8'b10000000; // 3261 : 128 - 0x80
      13'hCBE: dout <= 8'b00000000; // 3262 :   0 - 0x0
      13'hCBF: dout <= 8'b00000000; // 3263 :   0 - 0x0
      13'hCC0: dout <= 8'b11000011; // 3264 : 195 - 0xc3 -- Sprite 0xcc
      13'hCC1: dout <= 8'b01110000; // 3265 : 112 - 0x70
      13'hCC2: dout <= 8'b00000000; // 3266 :   0 - 0x0
      13'hCC3: dout <= 8'b01100000; // 3267 :  96 - 0x60
      13'hCC4: dout <= 8'b11110000; // 3268 : 240 - 0xf0
      13'hCC5: dout <= 8'b11010000; // 3269 : 208 - 0xd0
      13'hCC6: dout <= 8'b10010000; // 3270 : 144 - 0x90
      13'hCC7: dout <= 8'b01100000; // 3271 :  96 - 0x60
      13'hCC8: dout <= 8'b00110000; // 3272 :  48 - 0x30
      13'hCC9: dout <= 8'b00000000; // 3273 :   0 - 0x0
      13'hCCA: dout <= 8'b00000000; // 3274 :   0 - 0x0
      13'hCCB: dout <= 8'b00000000; // 3275 :   0 - 0x0
      13'hCCC: dout <= 8'b00000000; // 3276 :   0 - 0x0
      13'hCCD: dout <= 8'b01100000; // 3277 :  96 - 0x60
      13'hCCE: dout <= 8'b01100000; // 3278 :  96 - 0x60
      13'hCCF: dout <= 8'b00000000; // 3279 :   0 - 0x0
      13'hCD0: dout <= 8'b11000000; // 3280 : 192 - 0xc0 -- Sprite 0xcd
      13'hCD1: dout <= 8'b00000000; // 3281 :   0 - 0x0
      13'hCD2: dout <= 8'b00000000; // 3282 :   0 - 0x0
      13'hCD3: dout <= 8'b00000110; // 3283 :   6 - 0x6
      13'hCD4: dout <= 8'b00001111; // 3284 :  15 - 0xf
      13'hCD5: dout <= 8'b00001101; // 3285 :  13 - 0xd
      13'hCD6: dout <= 8'b00001001; // 3286 :   9 - 0x9
      13'hCD7: dout <= 8'b00000110; // 3287 :   6 - 0x6
      13'hCD8: dout <= 8'b00000000; // 3288 :   0 - 0x0
      13'hCD9: dout <= 8'b00000000; // 3289 :   0 - 0x0
      13'hCDA: dout <= 8'b00000000; // 3290 :   0 - 0x0
      13'hCDB: dout <= 8'b00000000; // 3291 :   0 - 0x0
      13'hCDC: dout <= 8'b00000000; // 3292 :   0 - 0x0
      13'hCDD: dout <= 8'b00000110; // 3293 :   6 - 0x6
      13'hCDE: dout <= 8'b00000110; // 3294 :   6 - 0x6
      13'hCDF: dout <= 8'b00000000; // 3295 :   0 - 0x0
      13'hCE0: dout <= 8'b11111100; // 3296 : 252 - 0xfc -- Sprite 0xce
      13'hCE1: dout <= 8'b11000000; // 3297 : 192 - 0xc0
      13'hCE2: dout <= 8'b11010001; // 3298 : 209 - 0xd1
      13'hCE3: dout <= 8'b11000010; // 3299 : 194 - 0xc2
      13'hCE4: dout <= 8'b10011110; // 3300 : 158 - 0x9e
      13'hCE5: dout <= 8'b10111111; // 3301 : 191 - 0xbf
      13'hCE6: dout <= 8'b10110000; // 3302 : 176 - 0xb0
      13'hCE7: dout <= 8'b10110011; // 3303 : 179 - 0xb3
      13'hCE8: dout <= 8'b00000000; // 3304 :   0 - 0x0
      13'hCE9: dout <= 8'b00000001; // 3305 :   1 - 0x1
      13'hCEA: dout <= 8'b00011011; // 3306 :  27 - 0x1b
      13'hCEB: dout <= 8'b00010011; // 3307 :  19 - 0x13
      13'hCEC: dout <= 8'b00011111; // 3308 :  31 - 0x1f
      13'hCED: dout <= 8'b00111111; // 3309 :  63 - 0x3f
      13'hCEE: dout <= 8'b00111111; // 3310 :  63 - 0x3f
      13'hCEF: dout <= 8'b00111111; // 3311 :  63 - 0x3f
      13'hCF0: dout <= 8'b00000111; // 3312 :   7 - 0x7 -- Sprite 0xcf
      13'hCF1: dout <= 8'b11110011; // 3313 : 243 - 0xf3
      13'hCF2: dout <= 8'b00001011; // 3314 :  11 - 0xb
      13'hCF3: dout <= 8'b01111011; // 3315 : 123 - 0x7b
      13'hCF4: dout <= 8'b01111011; // 3316 : 123 - 0x7b
      13'hCF5: dout <= 8'b11111001; // 3317 : 249 - 0xf9
      13'hCF6: dout <= 8'b00001101; // 3318 :  13 - 0xd
      13'hCF7: dout <= 8'b11101101; // 3319 : 237 - 0xed
      13'hCF8: dout <= 8'b00000000; // 3320 :   0 - 0x0
      13'hCF9: dout <= 8'b11111000; // 3321 : 248 - 0xf8
      13'hCFA: dout <= 8'b00001000; // 3322 :   8 - 0x8
      13'hCFB: dout <= 8'b00001000; // 3323 :   8 - 0x8
      13'hCFC: dout <= 8'b00001000; // 3324 :   8 - 0x8
      13'hCFD: dout <= 8'b11111000; // 3325 : 248 - 0xf8
      13'hCFE: dout <= 8'b11110000; // 3326 : 240 - 0xf0
      13'hCFF: dout <= 8'b11010000; // 3327 : 208 - 0xd0
      13'hD00: dout <= 8'b11111111; // 3328 : 255 - 0xff -- Sprite 0xd0
      13'hD01: dout <= 8'b11111111; // 3329 : 255 - 0xff
      13'hD02: dout <= 8'b11111111; // 3330 : 255 - 0xff
      13'hD03: dout <= 8'b11111111; // 3331 : 255 - 0xff
      13'hD04: dout <= 8'b11101110; // 3332 : 238 - 0xee
      13'hD05: dout <= 8'b11101110; // 3333 : 238 - 0xee
      13'hD06: dout <= 8'b11101110; // 3334 : 238 - 0xee
      13'hD07: dout <= 8'b11101110; // 3335 : 238 - 0xee
      13'hD08: dout <= 8'b00000000; // 3336 :   0 - 0x0
      13'hD09: dout <= 8'b00000000; // 3337 :   0 - 0x0
      13'hD0A: dout <= 8'b01111100; // 3338 : 124 - 0x7c
      13'hD0B: dout <= 8'b11111110; // 3339 : 254 - 0xfe
      13'hD0C: dout <= 8'b11101110; // 3340 : 238 - 0xee
      13'hD0D: dout <= 8'b11101110; // 3341 : 238 - 0xee
      13'hD0E: dout <= 8'b11101110; // 3342 : 238 - 0xee
      13'hD0F: dout <= 8'b11101110; // 3343 : 238 - 0xee
      13'hD10: dout <= 8'b11111111; // 3344 : 255 - 0xff -- Sprite 0xd1
      13'hD11: dout <= 8'b11111111; // 3345 : 255 - 0xff
      13'hD12: dout <= 8'b11111111; // 3346 : 255 - 0xff
      13'hD13: dout <= 8'b11111011; // 3347 : 251 - 0xfb
      13'hD14: dout <= 8'b11111011; // 3348 : 251 - 0xfb
      13'hD15: dout <= 8'b11111011; // 3349 : 251 - 0xfb
      13'hD16: dout <= 8'b11111011; // 3350 : 251 - 0xfb
      13'hD17: dout <= 8'b11111011; // 3351 : 251 - 0xfb
      13'hD18: dout <= 8'b00000000; // 3352 :   0 - 0x0
      13'hD19: dout <= 8'b00000000; // 3353 :   0 - 0x0
      13'hD1A: dout <= 8'b00111000; // 3354 :  56 - 0x38
      13'hD1B: dout <= 8'b01111000; // 3355 : 120 - 0x78
      13'hD1C: dout <= 8'b01111000; // 3356 : 120 - 0x78
      13'hD1D: dout <= 8'b00111000; // 3357 :  56 - 0x38
      13'hD1E: dout <= 8'b00111000; // 3358 :  56 - 0x38
      13'hD1F: dout <= 8'b00111000; // 3359 :  56 - 0x38
      13'hD20: dout <= 8'b11111111; // 3360 : 255 - 0xff -- Sprite 0xd2
      13'hD21: dout <= 8'b11111111; // 3361 : 255 - 0xff
      13'hD22: dout <= 8'b11111111; // 3362 : 255 - 0xff
      13'hD23: dout <= 8'b11111111; // 3363 : 255 - 0xff
      13'hD24: dout <= 8'b11101110; // 3364 : 238 - 0xee
      13'hD25: dout <= 8'b10001110; // 3365 : 142 - 0x8e
      13'hD26: dout <= 8'b11111110; // 3366 : 254 - 0xfe
      13'hD27: dout <= 8'b11111110; // 3367 : 254 - 0xfe
      13'hD28: dout <= 8'b00000000; // 3368 :   0 - 0x0
      13'hD29: dout <= 8'b00000000; // 3369 :   0 - 0x0
      13'hD2A: dout <= 8'b01111100; // 3370 : 124 - 0x7c
      13'hD2B: dout <= 8'b11111110; // 3371 : 254 - 0xfe
      13'hD2C: dout <= 8'b11101110; // 3372 : 238 - 0xee
      13'hD2D: dout <= 8'b00001110; // 3373 :  14 - 0xe
      13'hD2E: dout <= 8'b00001110; // 3374 :  14 - 0xe
      13'hD2F: dout <= 8'b01111110; // 3375 : 126 - 0x7e
      13'hD30: dout <= 8'b11111111; // 3376 : 255 - 0xff -- Sprite 0xd3
      13'hD31: dout <= 8'b11111111; // 3377 : 255 - 0xff
      13'hD32: dout <= 8'b11111111; // 3378 : 255 - 0xff
      13'hD33: dout <= 8'b11111111; // 3379 : 255 - 0xff
      13'hD34: dout <= 8'b11101110; // 3380 : 238 - 0xee
      13'hD35: dout <= 8'b10001110; // 3381 : 142 - 0x8e
      13'hD36: dout <= 8'b11111100; // 3382 : 252 - 0xfc
      13'hD37: dout <= 8'b11111101; // 3383 : 253 - 0xfd
      13'hD38: dout <= 8'b00000000; // 3384 :   0 - 0x0
      13'hD39: dout <= 8'b00000000; // 3385 :   0 - 0x0
      13'hD3A: dout <= 8'b01111100; // 3386 : 124 - 0x7c
      13'hD3B: dout <= 8'b11111110; // 3387 : 254 - 0xfe
      13'hD3C: dout <= 8'b11101110; // 3388 : 238 - 0xee
      13'hD3D: dout <= 8'b00001110; // 3389 :  14 - 0xe
      13'hD3E: dout <= 8'b00111100; // 3390 :  60 - 0x3c
      13'hD3F: dout <= 8'b00111100; // 3391 :  60 - 0x3c
      13'hD40: dout <= 8'b11111111; // 3392 : 255 - 0xff -- Sprite 0xd4
      13'hD41: dout <= 8'b11111111; // 3393 : 255 - 0xff
      13'hD42: dout <= 8'b11111111; // 3394 : 255 - 0xff
      13'hD43: dout <= 8'b11111110; // 3395 : 254 - 0xfe
      13'hD44: dout <= 8'b11101110; // 3396 : 238 - 0xee
      13'hD45: dout <= 8'b11101110; // 3397 : 238 - 0xee
      13'hD46: dout <= 8'b11101110; // 3398 : 238 - 0xee
      13'hD47: dout <= 8'b11101110; // 3399 : 238 - 0xee
      13'hD48: dout <= 8'b00000000; // 3400 :   0 - 0x0
      13'hD49: dout <= 8'b00000000; // 3401 :   0 - 0x0
      13'hD4A: dout <= 8'b00111110; // 3402 :  62 - 0x3e
      13'hD4B: dout <= 8'b01111110; // 3403 : 126 - 0x7e
      13'hD4C: dout <= 8'b11101110; // 3404 : 238 - 0xee
      13'hD4D: dout <= 8'b11101110; // 3405 : 238 - 0xee
      13'hD4E: dout <= 8'b11101110; // 3406 : 238 - 0xee
      13'hD4F: dout <= 8'b11101110; // 3407 : 238 - 0xee
      13'hD50: dout <= 8'b11111111; // 3408 : 255 - 0xff -- Sprite 0xd5
      13'hD51: dout <= 8'b11111111; // 3409 : 255 - 0xff
      13'hD52: dout <= 8'b11111111; // 3410 : 255 - 0xff
      13'hD53: dout <= 8'b11111101; // 3411 : 253 - 0xfd
      13'hD54: dout <= 8'b11100001; // 3412 : 225 - 0xe1
      13'hD55: dout <= 8'b11101111; // 3413 : 239 - 0xef
      13'hD56: dout <= 8'b11111111; // 3414 : 255 - 0xff
      13'hD57: dout <= 8'b11111111; // 3415 : 255 - 0xff
      13'hD58: dout <= 8'b00000000; // 3416 :   0 - 0x0
      13'hD59: dout <= 8'b00000000; // 3417 :   0 - 0x0
      13'hD5A: dout <= 8'b11111100; // 3418 : 252 - 0xfc
      13'hD5B: dout <= 8'b11111100; // 3419 : 252 - 0xfc
      13'hD5C: dout <= 8'b11100000; // 3420 : 224 - 0xe0
      13'hD5D: dout <= 8'b11100000; // 3421 : 224 - 0xe0
      13'hD5E: dout <= 8'b11111100; // 3422 : 252 - 0xfc
      13'hD5F: dout <= 8'b11111110; // 3423 : 254 - 0xfe
      13'hD60: dout <= 8'b11111111; // 3424 : 255 - 0xff -- Sprite 0xd6
      13'hD61: dout <= 8'b11111111; // 3425 : 255 - 0xff
      13'hD62: dout <= 8'b11111111; // 3426 : 255 - 0xff
      13'hD63: dout <= 8'b11111101; // 3427 : 253 - 0xfd
      13'hD64: dout <= 8'b11100001; // 3428 : 225 - 0xe1
      13'hD65: dout <= 8'b11101111; // 3429 : 239 - 0xef
      13'hD66: dout <= 8'b11111111; // 3430 : 255 - 0xff
      13'hD67: dout <= 8'b11111111; // 3431 : 255 - 0xff
      13'hD68: dout <= 8'b00000000; // 3432 :   0 - 0x0
      13'hD69: dout <= 8'b00000000; // 3433 :   0 - 0x0
      13'hD6A: dout <= 8'b01111100; // 3434 : 124 - 0x7c
      13'hD6B: dout <= 8'b11111100; // 3435 : 252 - 0xfc
      13'hD6C: dout <= 8'b11100000; // 3436 : 224 - 0xe0
      13'hD6D: dout <= 8'b11100000; // 3437 : 224 - 0xe0
      13'hD6E: dout <= 8'b11111100; // 3438 : 252 - 0xfc
      13'hD6F: dout <= 8'b11111110; // 3439 : 254 - 0xfe
      13'hD70: dout <= 8'b11111111; // 3440 : 255 - 0xff -- Sprite 0xd7
      13'hD71: dout <= 8'b11111111; // 3441 : 255 - 0xff
      13'hD72: dout <= 8'b11111111; // 3442 : 255 - 0xff
      13'hD73: dout <= 8'b11111110; // 3443 : 254 - 0xfe
      13'hD74: dout <= 8'b11101110; // 3444 : 238 - 0xee
      13'hD75: dout <= 8'b10001110; // 3445 : 142 - 0x8e
      13'hD76: dout <= 8'b11111110; // 3446 : 254 - 0xfe
      13'hD77: dout <= 8'b11111100; // 3447 : 252 - 0xfc
      13'hD78: dout <= 8'b00000000; // 3448 :   0 - 0x0
      13'hD79: dout <= 8'b00000000; // 3449 :   0 - 0x0
      13'hD7A: dout <= 8'b11111110; // 3450 : 254 - 0xfe
      13'hD7B: dout <= 8'b11111110; // 3451 : 254 - 0xfe
      13'hD7C: dout <= 8'b11101110; // 3452 : 238 - 0xee
      13'hD7D: dout <= 8'b00001110; // 3453 :  14 - 0xe
      13'hD7E: dout <= 8'b00001110; // 3454 :  14 - 0xe
      13'hD7F: dout <= 8'b00011100; // 3455 :  28 - 0x1c
      13'hD80: dout <= 8'b11111111; // 3456 : 255 - 0xff -- Sprite 0xd8
      13'hD81: dout <= 8'b11111111; // 3457 : 255 - 0xff
      13'hD82: dout <= 8'b11111111; // 3458 : 255 - 0xff
      13'hD83: dout <= 8'b11111111; // 3459 : 255 - 0xff
      13'hD84: dout <= 8'b11101110; // 3460 : 238 - 0xee
      13'hD85: dout <= 8'b11101110; // 3461 : 238 - 0xee
      13'hD86: dout <= 8'b11111100; // 3462 : 252 - 0xfc
      13'hD87: dout <= 8'b11111111; // 3463 : 255 - 0xff
      13'hD88: dout <= 8'b00000000; // 3464 :   0 - 0x0
      13'hD89: dout <= 8'b00000000; // 3465 :   0 - 0x0
      13'hD8A: dout <= 8'b01111100; // 3466 : 124 - 0x7c
      13'hD8B: dout <= 8'b11111110; // 3467 : 254 - 0xfe
      13'hD8C: dout <= 8'b11101110; // 3468 : 238 - 0xee
      13'hD8D: dout <= 8'b11101110; // 3469 : 238 - 0xee
      13'hD8E: dout <= 8'b01111100; // 3470 : 124 - 0x7c
      13'hD8F: dout <= 8'b11111110; // 3471 : 254 - 0xfe
      13'hD90: dout <= 8'b11111111; // 3472 : 255 - 0xff -- Sprite 0xd9
      13'hD91: dout <= 8'b11111111; // 3473 : 255 - 0xff
      13'hD92: dout <= 8'b11111111; // 3474 : 255 - 0xff
      13'hD93: dout <= 8'b11111111; // 3475 : 255 - 0xff
      13'hD94: dout <= 8'b11101110; // 3476 : 238 - 0xee
      13'hD95: dout <= 8'b11101110; // 3477 : 238 - 0xee
      13'hD96: dout <= 8'b11101110; // 3478 : 238 - 0xee
      13'hD97: dout <= 8'b11101110; // 3479 : 238 - 0xee
      13'hD98: dout <= 8'b00000000; // 3480 :   0 - 0x0
      13'hD99: dout <= 8'b00000000; // 3481 :   0 - 0x0
      13'hD9A: dout <= 8'b01111100; // 3482 : 124 - 0x7c
      13'hD9B: dout <= 8'b11111110; // 3483 : 254 - 0xfe
      13'hD9C: dout <= 8'b11101110; // 3484 : 238 - 0xee
      13'hD9D: dout <= 8'b11101110; // 3485 : 238 - 0xee
      13'hD9E: dout <= 8'b11101110; // 3486 : 238 - 0xee
      13'hD9F: dout <= 8'b11101110; // 3487 : 238 - 0xee
      13'hDA0: dout <= 8'b00000000; // 3488 :   0 - 0x0 -- Sprite 0xda
      13'hDA1: dout <= 8'b00000000; // 3489 :   0 - 0x0
      13'hDA2: dout <= 8'b00000000; // 3490 :   0 - 0x0
      13'hDA3: dout <= 8'b10000000; // 3491 : 128 - 0x80
      13'hDA4: dout <= 8'b00000000; // 3492 :   0 - 0x0
      13'hDA5: dout <= 8'b00000000; // 3493 :   0 - 0x0
      13'hDA6: dout <= 8'b00000100; // 3494 :   4 - 0x4
      13'hDA7: dout <= 8'b00000000; // 3495 :   0 - 0x0
      13'hDA8: dout <= 8'b00000000; // 3496 :   0 - 0x0
      13'hDA9: dout <= 8'b00100000; // 3497 :  32 - 0x20
      13'hDAA: dout <= 8'b00000000; // 3498 :   0 - 0x0
      13'hDAB: dout <= 8'b00000010; // 3499 :   2 - 0x2
      13'hDAC: dout <= 8'b00000000; // 3500 :   0 - 0x0
      13'hDAD: dout <= 8'b00100000; // 3501 :  32 - 0x20
      13'hDAE: dout <= 8'b00000000; // 3502 :   0 - 0x0
      13'hDAF: dout <= 8'b00000000; // 3503 :   0 - 0x0
      13'hDB0: dout <= 8'b00000000; // 3504 :   0 - 0x0 -- Sprite 0xdb
      13'hDB1: dout <= 8'b00000100; // 3505 :   4 - 0x4
      13'hDB2: dout <= 8'b00000000; // 3506 :   0 - 0x0
      13'hDB3: dout <= 8'b00010001; // 3507 :  17 - 0x11
      13'hDB4: dout <= 8'b00000000; // 3508 :   0 - 0x0
      13'hDB5: dout <= 8'b00000000; // 3509 :   0 - 0x0
      13'hDB6: dout <= 8'b00000000; // 3510 :   0 - 0x0
      13'hDB7: dout <= 8'b00100000; // 3511 :  32 - 0x20
      13'hDB8: dout <= 8'b00100000; // 3512 :  32 - 0x20
      13'hDB9: dout <= 8'b00000000; // 3513 :   0 - 0x0
      13'hDBA: dout <= 8'b00000000; // 3514 :   0 - 0x0
      13'hDBB: dout <= 8'b00000000; // 3515 :   0 - 0x0
      13'hDBC: dout <= 8'b10000000; // 3516 : 128 - 0x80
      13'hDBD: dout <= 8'b00000000; // 3517 :   0 - 0x0
      13'hDBE: dout <= 8'b00000100; // 3518 :   4 - 0x4
      13'hDBF: dout <= 8'b00000000; // 3519 :   0 - 0x0
      13'hDC0: dout <= 8'b00000000; // 3520 :   0 - 0x0 -- Sprite 0xdc
      13'hDC1: dout <= 8'b00000000; // 3521 :   0 - 0x0
      13'hDC2: dout <= 8'b00000000; // 3522 :   0 - 0x0
      13'hDC3: dout <= 8'b00100000; // 3523 :  32 - 0x20
      13'hDC4: dout <= 8'b00000000; // 3524 :   0 - 0x0
      13'hDC5: dout <= 8'b00000000; // 3525 :   0 - 0x0
      13'hDC6: dout <= 8'b00000000; // 3526 :   0 - 0x0
      13'hDC7: dout <= 8'b00000100; // 3527 :   4 - 0x4
      13'hDC8: dout <= 8'b00000000; // 3528 :   0 - 0x0
      13'hDC9: dout <= 8'b00001000; // 3529 :   8 - 0x8
      13'hDCA: dout <= 8'b00000000; // 3530 :   0 - 0x0
      13'hDCB: dout <= 8'b00000000; // 3531 :   0 - 0x0
      13'hDCC: dout <= 8'b00000010; // 3532 :   2 - 0x2
      13'hDCD: dout <= 8'b00000000; // 3533 :   0 - 0x0
      13'hDCE: dout <= 8'b01000000; // 3534 :  64 - 0x40
      13'hDCF: dout <= 8'b00000000; // 3535 :   0 - 0x0
      13'hDD0: dout <= 8'b00000000; // 3536 :   0 - 0x0 -- Sprite 0xdd
      13'hDD1: dout <= 8'b00000000; // 3537 :   0 - 0x0
      13'hDD2: dout <= 8'b00010001; // 3538 :  17 - 0x11
      13'hDD3: dout <= 8'b00000000; // 3539 :   0 - 0x0
      13'hDD4: dout <= 8'b00000000; // 3540 :   0 - 0x0
      13'hDD5: dout <= 8'b10000000; // 3541 : 128 - 0x80
      13'hDD6: dout <= 8'b00000000; // 3542 :   0 - 0x0
      13'hDD7: dout <= 8'b00000000; // 3543 :   0 - 0x0
      13'hDD8: dout <= 8'b00000000; // 3544 :   0 - 0x0
      13'hDD9: dout <= 8'b01000000; // 3545 :  64 - 0x40
      13'hDDA: dout <= 8'b00000000; // 3546 :   0 - 0x0
      13'hDDB: dout <= 8'b00000000; // 3547 :   0 - 0x0
      13'hDDC: dout <= 8'b00000000; // 3548 :   0 - 0x0
      13'hDDD: dout <= 8'b00000000; // 3549 :   0 - 0x0
      13'hDDE: dout <= 8'b00000010; // 3550 :   2 - 0x2
      13'hDDF: dout <= 8'b00100000; // 3551 :  32 - 0x20
      13'hDE0: dout <= 8'b10110011; // 3552 : 179 - 0xb3 -- Sprite 0xde
      13'hDE1: dout <= 8'b10110011; // 3553 : 179 - 0xb3
      13'hDE2: dout <= 8'b10110011; // 3554 : 179 - 0xb3
      13'hDE3: dout <= 8'b10110011; // 3555 : 179 - 0xb3
      13'hDE4: dout <= 8'b10110000; // 3556 : 176 - 0xb0
      13'hDE5: dout <= 8'b10101111; // 3557 : 175 - 0xaf
      13'hDE6: dout <= 8'b10011111; // 3558 : 159 - 0x9f
      13'hDE7: dout <= 8'b11000000; // 3559 : 192 - 0xc0
      13'hDE8: dout <= 8'b00111110; // 3560 :  62 - 0x3e
      13'hDE9: dout <= 8'b00111111; // 3561 :  63 - 0x3f
      13'hDEA: dout <= 8'b00111110; // 3562 :  62 - 0x3e
      13'hDEB: dout <= 8'b00111100; // 3563 :  60 - 0x3c
      13'hDEC: dout <= 8'b00111111; // 3564 :  63 - 0x3f
      13'hDED: dout <= 8'b00110000; // 3565 :  48 - 0x30
      13'hDEE: dout <= 8'b00000000; // 3566 :   0 - 0x0
      13'hDEF: dout <= 8'b00000000; // 3567 :   0 - 0x0
      13'hDF0: dout <= 8'b11101101; // 3568 : 237 - 0xed -- Sprite 0xdf
      13'hDF1: dout <= 8'b11001101; // 3569 : 205 - 0xcd
      13'hDF2: dout <= 8'b11001101; // 3570 : 205 - 0xcd
      13'hDF3: dout <= 8'b00001101; // 3571 :  13 - 0xd
      13'hDF4: dout <= 8'b00001101; // 3572 :  13 - 0xd
      13'hDF5: dout <= 8'b11111101; // 3573 : 253 - 0xfd
      13'hDF6: dout <= 8'b11111101; // 3574 : 253 - 0xfd
      13'hDF7: dout <= 8'b00000011; // 3575 :   3 - 0x3
      13'hDF8: dout <= 8'b00010000; // 3576 :  16 - 0x10
      13'hDF9: dout <= 8'b10110000; // 3577 : 176 - 0xb0
      13'hDFA: dout <= 8'b00110000; // 3578 :  48 - 0x30
      13'hDFB: dout <= 8'b11110000; // 3579 : 240 - 0xf0
      13'hDFC: dout <= 8'b11110000; // 3580 : 240 - 0xf0
      13'hDFD: dout <= 8'b00000000; // 3581 :   0 - 0x0
      13'hDFE: dout <= 8'b00000000; // 3582 :   0 - 0x0
      13'hDFF: dout <= 8'b00000000; // 3583 :   0 - 0x0
      13'hE00: dout <= 8'b11101110; // 3584 : 238 - 0xee -- Sprite 0xe0
      13'hE01: dout <= 8'b11101110; // 3585 : 238 - 0xee
      13'hE02: dout <= 8'b11101110; // 3586 : 238 - 0xee
      13'hE03: dout <= 8'b11101110; // 3587 : 238 - 0xee
      13'hE04: dout <= 8'b11111110; // 3588 : 254 - 0xfe
      13'hE05: dout <= 8'b11111100; // 3589 : 252 - 0xfc
      13'hE06: dout <= 8'b11000001; // 3590 : 193 - 0xc1
      13'hE07: dout <= 8'b11111111; // 3591 : 255 - 0xff
      13'hE08: dout <= 8'b11101110; // 3592 : 238 - 0xee
      13'hE09: dout <= 8'b11101110; // 3593 : 238 - 0xee
      13'hE0A: dout <= 8'b11101110; // 3594 : 238 - 0xee
      13'hE0B: dout <= 8'b11101110; // 3595 : 238 - 0xee
      13'hE0C: dout <= 8'b11111110; // 3596 : 254 - 0xfe
      13'hE0D: dout <= 8'b01111100; // 3597 : 124 - 0x7c
      13'hE0E: dout <= 8'b00000000; // 3598 :   0 - 0x0
      13'hE0F: dout <= 8'b00000000; // 3599 :   0 - 0x0
      13'hE10: dout <= 8'b11111011; // 3600 : 251 - 0xfb -- Sprite 0xe1
      13'hE11: dout <= 8'b11111011; // 3601 : 251 - 0xfb
      13'hE12: dout <= 8'b11111011; // 3602 : 251 - 0xfb
      13'hE13: dout <= 8'b11111011; // 3603 : 251 - 0xfb
      13'hE14: dout <= 8'b11111111; // 3604 : 255 - 0xff
      13'hE15: dout <= 8'b11111101; // 3605 : 253 - 0xfd
      13'hE16: dout <= 8'b11000001; // 3606 : 193 - 0xc1
      13'hE17: dout <= 8'b11111111; // 3607 : 255 - 0xff
      13'hE18: dout <= 8'b00111000; // 3608 :  56 - 0x38
      13'hE19: dout <= 8'b00111000; // 3609 :  56 - 0x38
      13'hE1A: dout <= 8'b00111000; // 3610 :  56 - 0x38
      13'hE1B: dout <= 8'b00111000; // 3611 :  56 - 0x38
      13'hE1C: dout <= 8'b01111100; // 3612 : 124 - 0x7c
      13'hE1D: dout <= 8'b01111100; // 3613 : 124 - 0x7c
      13'hE1E: dout <= 8'b00000000; // 3614 :   0 - 0x0
      13'hE1F: dout <= 8'b00000000; // 3615 :   0 - 0x0
      13'hE20: dout <= 8'b11111100; // 3616 : 252 - 0xfc -- Sprite 0xe2
      13'hE21: dout <= 8'b11100001; // 3617 : 225 - 0xe1
      13'hE22: dout <= 8'b11101111; // 3618 : 239 - 0xef
      13'hE23: dout <= 8'b11101111; // 3619 : 239 - 0xef
      13'hE24: dout <= 8'b11111111; // 3620 : 255 - 0xff
      13'hE25: dout <= 8'b11111110; // 3621 : 254 - 0xfe
      13'hE26: dout <= 8'b10000000; // 3622 : 128 - 0x80
      13'hE27: dout <= 8'b11111111; // 3623 : 255 - 0xff
      13'hE28: dout <= 8'b11111100; // 3624 : 252 - 0xfc
      13'hE29: dout <= 8'b11100000; // 3625 : 224 - 0xe0
      13'hE2A: dout <= 8'b11100000; // 3626 : 224 - 0xe0
      13'hE2B: dout <= 8'b11100000; // 3627 : 224 - 0xe0
      13'hE2C: dout <= 8'b11111110; // 3628 : 254 - 0xfe
      13'hE2D: dout <= 8'b11111110; // 3629 : 254 - 0xfe
      13'hE2E: dout <= 8'b00000000; // 3630 :   0 - 0x0
      13'hE2F: dout <= 8'b00000000; // 3631 :   0 - 0x0
      13'hE30: dout <= 8'b11101110; // 3632 : 238 - 0xee -- Sprite 0xe3
      13'hE31: dout <= 8'b11111110; // 3633 : 254 - 0xfe
      13'hE32: dout <= 8'b11111110; // 3634 : 254 - 0xfe
      13'hE33: dout <= 8'b11111110; // 3635 : 254 - 0xfe
      13'hE34: dout <= 8'b11111110; // 3636 : 254 - 0xfe
      13'hE35: dout <= 8'b11111100; // 3637 : 252 - 0xfc
      13'hE36: dout <= 8'b11000001; // 3638 : 193 - 0xc1
      13'hE37: dout <= 8'b11111111; // 3639 : 255 - 0xff
      13'hE38: dout <= 8'b00001110; // 3640 :  14 - 0xe
      13'hE39: dout <= 8'b00001110; // 3641 :  14 - 0xe
      13'hE3A: dout <= 8'b00001110; // 3642 :  14 - 0xe
      13'hE3B: dout <= 8'b11101110; // 3643 : 238 - 0xee
      13'hE3C: dout <= 8'b11111110; // 3644 : 254 - 0xfe
      13'hE3D: dout <= 8'b01111100; // 3645 : 124 - 0x7c
      13'hE3E: dout <= 8'b00000000; // 3646 :   0 - 0x0
      13'hE3F: dout <= 8'b00000000; // 3647 :   0 - 0x0
      13'hE40: dout <= 8'b11101110; // 3648 : 238 - 0xee -- Sprite 0xe4
      13'hE41: dout <= 8'b11101110; // 3649 : 238 - 0xee
      13'hE42: dout <= 8'b11111110; // 3650 : 254 - 0xfe
      13'hE43: dout <= 8'b11111110; // 3651 : 254 - 0xfe
      13'hE44: dout <= 8'b10001110; // 3652 : 142 - 0x8e
      13'hE45: dout <= 8'b11111110; // 3653 : 254 - 0xfe
      13'hE46: dout <= 8'b11111000; // 3654 : 248 - 0xf8
      13'hE47: dout <= 8'b11111111; // 3655 : 255 - 0xff
      13'hE48: dout <= 8'b11101110; // 3656 : 238 - 0xee
      13'hE49: dout <= 8'b11101110; // 3657 : 238 - 0xee
      13'hE4A: dout <= 8'b11111110; // 3658 : 254 - 0xfe
      13'hE4B: dout <= 8'b11111110; // 3659 : 254 - 0xfe
      13'hE4C: dout <= 8'b00001110; // 3660 :  14 - 0xe
      13'hE4D: dout <= 8'b00001110; // 3661 :  14 - 0xe
      13'hE4E: dout <= 8'b00000000; // 3662 :   0 - 0x0
      13'hE4F: dout <= 8'b00000000; // 3663 :   0 - 0x0
      13'hE50: dout <= 8'b10001110; // 3664 : 142 - 0x8e -- Sprite 0xe5
      13'hE51: dout <= 8'b11111110; // 3665 : 254 - 0xfe
      13'hE52: dout <= 8'b11111110; // 3666 : 254 - 0xfe
      13'hE53: dout <= 8'b11111110; // 3667 : 254 - 0xfe
      13'hE54: dout <= 8'b11111110; // 3668 : 254 - 0xfe
      13'hE55: dout <= 8'b11111100; // 3669 : 252 - 0xfc
      13'hE56: dout <= 8'b11000001; // 3670 : 193 - 0xc1
      13'hE57: dout <= 8'b11111111; // 3671 : 255 - 0xff
      13'hE58: dout <= 8'b00001110; // 3672 :  14 - 0xe
      13'hE59: dout <= 8'b00001110; // 3673 :  14 - 0xe
      13'hE5A: dout <= 8'b00001110; // 3674 :  14 - 0xe
      13'hE5B: dout <= 8'b11101110; // 3675 : 238 - 0xee
      13'hE5C: dout <= 8'b11111110; // 3676 : 254 - 0xfe
      13'hE5D: dout <= 8'b01111100; // 3677 : 124 - 0x7c
      13'hE5E: dout <= 8'b00000000; // 3678 :   0 - 0x0
      13'hE5F: dout <= 8'b00000000; // 3679 :   0 - 0x0
      13'hE60: dout <= 8'b11101110; // 3680 : 238 - 0xee -- Sprite 0xe6
      13'hE61: dout <= 8'b11101110; // 3681 : 238 - 0xee
      13'hE62: dout <= 8'b11101110; // 3682 : 238 - 0xee
      13'hE63: dout <= 8'b11101110; // 3683 : 238 - 0xee
      13'hE64: dout <= 8'b11111110; // 3684 : 254 - 0xfe
      13'hE65: dout <= 8'b11111100; // 3685 : 252 - 0xfc
      13'hE66: dout <= 8'b11000001; // 3686 : 193 - 0xc1
      13'hE67: dout <= 8'b11111111; // 3687 : 255 - 0xff
      13'hE68: dout <= 8'b11101110; // 3688 : 238 - 0xee
      13'hE69: dout <= 8'b11101110; // 3689 : 238 - 0xee
      13'hE6A: dout <= 8'b11101110; // 3690 : 238 - 0xee
      13'hE6B: dout <= 8'b11101110; // 3691 : 238 - 0xee
      13'hE6C: dout <= 8'b11111110; // 3692 : 254 - 0xfe
      13'hE6D: dout <= 8'b01111100; // 3693 : 124 - 0x7c
      13'hE6E: dout <= 8'b00000000; // 3694 :   0 - 0x0
      13'hE6F: dout <= 8'b00000000; // 3695 :   0 - 0x0
      13'hE70: dout <= 8'b11111101; // 3696 : 253 - 0xfd -- Sprite 0xe7
      13'hE71: dout <= 8'b11111101; // 3697 : 253 - 0xfd
      13'hE72: dout <= 8'b11111001; // 3698 : 249 - 0xf9
      13'hE73: dout <= 8'b11111011; // 3699 : 251 - 0xfb
      13'hE74: dout <= 8'b11111011; // 3700 : 251 - 0xfb
      13'hE75: dout <= 8'b11111011; // 3701 : 251 - 0xfb
      13'hE76: dout <= 8'b11100011; // 3702 : 227 - 0xe3
      13'hE77: dout <= 8'b11111111; // 3703 : 255 - 0xff
      13'hE78: dout <= 8'b00011100; // 3704 :  28 - 0x1c
      13'hE79: dout <= 8'b00011100; // 3705 :  28 - 0x1c
      13'hE7A: dout <= 8'b00111000; // 3706 :  56 - 0x38
      13'hE7B: dout <= 8'b00111000; // 3707 :  56 - 0x38
      13'hE7C: dout <= 8'b00111000; // 3708 :  56 - 0x38
      13'hE7D: dout <= 8'b00111000; // 3709 :  56 - 0x38
      13'hE7E: dout <= 8'b00000000; // 3710 :   0 - 0x0
      13'hE7F: dout <= 8'b00000000; // 3711 :   0 - 0x0
      13'hE80: dout <= 8'b11101110; // 3712 : 238 - 0xee -- Sprite 0xe8
      13'hE81: dout <= 8'b11101110; // 3713 : 238 - 0xee
      13'hE82: dout <= 8'b11101110; // 3714 : 238 - 0xee
      13'hE83: dout <= 8'b11101110; // 3715 : 238 - 0xee
      13'hE84: dout <= 8'b11111110; // 3716 : 254 - 0xfe
      13'hE85: dout <= 8'b11111100; // 3717 : 252 - 0xfc
      13'hE86: dout <= 8'b11000001; // 3718 : 193 - 0xc1
      13'hE87: dout <= 8'b11111111; // 3719 : 255 - 0xff
      13'hE88: dout <= 8'b11101110; // 3720 : 238 - 0xee
      13'hE89: dout <= 8'b11101110; // 3721 : 238 - 0xee
      13'hE8A: dout <= 8'b11101110; // 3722 : 238 - 0xee
      13'hE8B: dout <= 8'b11101110; // 3723 : 238 - 0xee
      13'hE8C: dout <= 8'b11111110; // 3724 : 254 - 0xfe
      13'hE8D: dout <= 8'b01111100; // 3725 : 124 - 0x7c
      13'hE8E: dout <= 8'b00000000; // 3726 :   0 - 0x0
      13'hE8F: dout <= 8'b00000000; // 3727 :   0 - 0x0
      13'hE90: dout <= 8'b11111110; // 3728 : 254 - 0xfe -- Sprite 0xe9
      13'hE91: dout <= 8'b11111110; // 3729 : 254 - 0xfe
      13'hE92: dout <= 8'b11001110; // 3730 : 206 - 0xce
      13'hE93: dout <= 8'b11111110; // 3731 : 254 - 0xfe
      13'hE94: dout <= 8'b11111110; // 3732 : 254 - 0xfe
      13'hE95: dout <= 8'b11111100; // 3733 : 252 - 0xfc
      13'hE96: dout <= 8'b11000001; // 3734 : 193 - 0xc1
      13'hE97: dout <= 8'b11111111; // 3735 : 255 - 0xff
      13'hE98: dout <= 8'b11111110; // 3736 : 254 - 0xfe
      13'hE99: dout <= 8'b01111110; // 3737 : 126 - 0x7e
      13'hE9A: dout <= 8'b00001110; // 3738 :  14 - 0xe
      13'hE9B: dout <= 8'b00001110; // 3739 :  14 - 0xe
      13'hE9C: dout <= 8'b01111110; // 3740 : 126 - 0x7e
      13'hE9D: dout <= 8'b01111100; // 3741 : 124 - 0x7c
      13'hE9E: dout <= 8'b00000000; // 3742 :   0 - 0x0
      13'hE9F: dout <= 8'b00000000; // 3743 :   0 - 0x0
      13'hEA0: dout <= 8'b00000000; // 3744 :   0 - 0x0 -- Sprite 0xea
      13'hEA1: dout <= 8'b01110000; // 3745 : 112 - 0x70
      13'hEA2: dout <= 8'b00111000; // 3746 :  56 - 0x38
      13'hEA3: dout <= 8'b00000000; // 3747 :   0 - 0x0
      13'hEA4: dout <= 8'b00000010; // 3748 :   2 - 0x2
      13'hEA5: dout <= 8'b00000111; // 3749 :   7 - 0x7
      13'hEA6: dout <= 8'b00000011; // 3750 :   3 - 0x3
      13'hEA7: dout <= 8'b00000000; // 3751 :   0 - 0x0
      13'hEA8: dout <= 8'b00000000; // 3752 :   0 - 0x0
      13'hEA9: dout <= 8'b01110000; // 3753 : 112 - 0x70
      13'hEAA: dout <= 8'b00111000; // 3754 :  56 - 0x38
      13'hEAB: dout <= 8'b00000000; // 3755 :   0 - 0x0
      13'hEAC: dout <= 8'b00000010; // 3756 :   2 - 0x2
      13'hEAD: dout <= 8'b00000111; // 3757 :   7 - 0x7
      13'hEAE: dout <= 8'b00000011; // 3758 :   3 - 0x3
      13'hEAF: dout <= 8'b00000000; // 3759 :   0 - 0x0
      13'hEB0: dout <= 8'b00000000; // 3760 :   0 - 0x0 -- Sprite 0xeb
      13'hEB1: dout <= 8'b00001100; // 3761 :  12 - 0xc
      13'hEB2: dout <= 8'b00000110; // 3762 :   6 - 0x6
      13'hEB3: dout <= 8'b00000110; // 3763 :   6 - 0x6
      13'hEB4: dout <= 8'b01100000; // 3764 :  96 - 0x60
      13'hEB5: dout <= 8'b01110000; // 3765 : 112 - 0x70
      13'hEB6: dout <= 8'b00110000; // 3766 :  48 - 0x30
      13'hEB7: dout <= 8'b00000000; // 3767 :   0 - 0x0
      13'hEB8: dout <= 8'b00000000; // 3768 :   0 - 0x0
      13'hEB9: dout <= 8'b00001100; // 3769 :  12 - 0xc
      13'hEBA: dout <= 8'b00000110; // 3770 :   6 - 0x6
      13'hEBB: dout <= 8'b00000110; // 3771 :   6 - 0x6
      13'hEBC: dout <= 8'b01100000; // 3772 :  96 - 0x60
      13'hEBD: dout <= 8'b01110000; // 3773 : 112 - 0x70
      13'hEBE: dout <= 8'b00110000; // 3774 :  48 - 0x30
      13'hEBF: dout <= 8'b00000000; // 3775 :   0 - 0x0
      13'hEC0: dout <= 8'b00000000; // 3776 :   0 - 0x0 -- Sprite 0xec
      13'hEC1: dout <= 8'b11000000; // 3777 : 192 - 0xc0
      13'hEC2: dout <= 8'b11100000; // 3778 : 224 - 0xe0
      13'hEC3: dout <= 8'b01100000; // 3779 :  96 - 0x60
      13'hEC4: dout <= 8'b00000000; // 3780 :   0 - 0x0
      13'hEC5: dout <= 8'b00001100; // 3781 :  12 - 0xc
      13'hEC6: dout <= 8'b00001110; // 3782 :  14 - 0xe
      13'hEC7: dout <= 8'b00000110; // 3783 :   6 - 0x6
      13'hEC8: dout <= 8'b00000000; // 3784 :   0 - 0x0
      13'hEC9: dout <= 8'b11000000; // 3785 : 192 - 0xc0
      13'hECA: dout <= 8'b11100000; // 3786 : 224 - 0xe0
      13'hECB: dout <= 8'b01100000; // 3787 :  96 - 0x60
      13'hECC: dout <= 8'b00000000; // 3788 :   0 - 0x0
      13'hECD: dout <= 8'b00001100; // 3789 :  12 - 0xc
      13'hECE: dout <= 8'b00001110; // 3790 :  14 - 0xe
      13'hECF: dout <= 8'b00000110; // 3791 :   6 - 0x6
      13'hED0: dout <= 8'b01100000; // 3792 :  96 - 0x60 -- Sprite 0xed
      13'hED1: dout <= 8'b01110000; // 3793 : 112 - 0x70
      13'hED2: dout <= 8'b00110000; // 3794 :  48 - 0x30
      13'hED3: dout <= 8'b00000000; // 3795 :   0 - 0x0
      13'hED4: dout <= 8'b00000000; // 3796 :   0 - 0x0
      13'hED5: dout <= 8'b00001100; // 3797 :  12 - 0xc
      13'hED6: dout <= 8'b00001110; // 3798 :  14 - 0xe
      13'hED7: dout <= 8'b00000110; // 3799 :   6 - 0x6
      13'hED8: dout <= 8'b01100000; // 3800 :  96 - 0x60
      13'hED9: dout <= 8'b01110000; // 3801 : 112 - 0x70
      13'hEDA: dout <= 8'b00110000; // 3802 :  48 - 0x30
      13'hEDB: dout <= 8'b00000000; // 3803 :   0 - 0x0
      13'hEDC: dout <= 8'b00000000; // 3804 :   0 - 0x0
      13'hEDD: dout <= 8'b00001100; // 3805 :  12 - 0xc
      13'hEDE: dout <= 8'b00001110; // 3806 :  14 - 0xe
      13'hEDF: dout <= 8'b00000110; // 3807 :   6 - 0x6
      13'hEE0: dout <= 8'b11111111; // 3808 : 255 - 0xff -- Sprite 0xee
      13'hEE1: dout <= 8'b11111111; // 3809 : 255 - 0xff
      13'hEE2: dout <= 8'b10111101; // 3810 : 189 - 0xbd
      13'hEE3: dout <= 8'b11111111; // 3811 : 255 - 0xff
      13'hEE4: dout <= 8'b11111111; // 3812 : 255 - 0xff
      13'hEE5: dout <= 8'b11111011; // 3813 : 251 - 0xfb
      13'hEE6: dout <= 8'b11111111; // 3814 : 255 - 0xff
      13'hEE7: dout <= 8'b11111111; // 3815 : 255 - 0xff
      13'hEE8: dout <= 8'b00000000; // 3816 :   0 - 0x0
      13'hEE9: dout <= 8'b00000000; // 3817 :   0 - 0x0
      13'hEEA: dout <= 8'b01000010; // 3818 :  66 - 0x42
      13'hEEB: dout <= 8'b00000000; // 3819 :   0 - 0x0
      13'hEEC: dout <= 8'b00000000; // 3820 :   0 - 0x0
      13'hEED: dout <= 8'b00000100; // 3821 :   4 - 0x4
      13'hEEE: dout <= 8'b00000000; // 3822 :   0 - 0x0
      13'hEEF: dout <= 8'b00000000; // 3823 :   0 - 0x0
      13'hEF0: dout <= 8'b11111111; // 3824 : 255 - 0xff -- Sprite 0xef
      13'hEF1: dout <= 8'b11111111; // 3825 : 255 - 0xff
      13'hEF2: dout <= 8'b11111011; // 3826 : 251 - 0xfb
      13'hEF3: dout <= 8'b11111111; // 3827 : 255 - 0xff
      13'hEF4: dout <= 8'b11011111; // 3828 : 223 - 0xdf
      13'hEF5: dout <= 8'b11111111; // 3829 : 255 - 0xff
      13'hEF6: dout <= 8'b11111111; // 3830 : 255 - 0xff
      13'hEF7: dout <= 8'b11111111; // 3831 : 255 - 0xff
      13'hEF8: dout <= 8'b00000000; // 3832 :   0 - 0x0
      13'hEF9: dout <= 8'b00000000; // 3833 :   0 - 0x0
      13'hEFA: dout <= 8'b00000100; // 3834 :   4 - 0x4
      13'hEFB: dout <= 8'b00000000; // 3835 :   0 - 0x0
      13'hEFC: dout <= 8'b00100000; // 3836 :  32 - 0x20
      13'hEFD: dout <= 8'b00000000; // 3837 :   0 - 0x0
      13'hEFE: dout <= 8'b00000000; // 3838 :   0 - 0x0
      13'hEFF: dout <= 8'b00000000; // 3839 :   0 - 0x0
      13'hF00: dout <= 8'b00000000; // 3840 :   0 - 0x0 -- Sprite 0xf0
      13'hF01: dout <= 8'b00000000; // 3841 :   0 - 0x0
      13'hF02: dout <= 8'b00000000; // 3842 :   0 - 0x0
      13'hF03: dout <= 8'b00000000; // 3843 :   0 - 0x0
      13'hF04: dout <= 8'b00000000; // 3844 :   0 - 0x0
      13'hF05: dout <= 8'b00000000; // 3845 :   0 - 0x0
      13'hF06: dout <= 8'b00000000; // 3846 :   0 - 0x0
      13'hF07: dout <= 8'b00000000; // 3847 :   0 - 0x0
      13'hF08: dout <= 8'b00000000; // 3848 :   0 - 0x0
      13'hF09: dout <= 8'b00000000; // 3849 :   0 - 0x0
      13'hF0A: dout <= 8'b00000000; // 3850 :   0 - 0x0
      13'hF0B: dout <= 8'b00000000; // 3851 :   0 - 0x0
      13'hF0C: dout <= 8'b00000000; // 3852 :   0 - 0x0
      13'hF0D: dout <= 8'b00000000; // 3853 :   0 - 0x0
      13'hF0E: dout <= 8'b00000000; // 3854 :   0 - 0x0
      13'hF0F: dout <= 8'b00000000; // 3855 :   0 - 0x0
      13'hF10: dout <= 8'b00000000; // 3856 :   0 - 0x0 -- Sprite 0xf1
      13'hF11: dout <= 8'b10000000; // 3857 : 128 - 0x80
      13'hF12: dout <= 8'b00000000; // 3858 :   0 - 0x0
      13'hF13: dout <= 8'b00000000; // 3859 :   0 - 0x0
      13'hF14: dout <= 8'b00000000; // 3860 :   0 - 0x0
      13'hF15: dout <= 8'b00000000; // 3861 :   0 - 0x0
      13'hF16: dout <= 8'b00000000; // 3862 :   0 - 0x0
      13'hF17: dout <= 8'b00000000; // 3863 :   0 - 0x0
      13'hF18: dout <= 8'b10000000; // 3864 : 128 - 0x80
      13'hF19: dout <= 8'b10000000; // 3865 : 128 - 0x80
      13'hF1A: dout <= 8'b10000000; // 3866 : 128 - 0x80
      13'hF1B: dout <= 8'b10000000; // 3867 : 128 - 0x80
      13'hF1C: dout <= 8'b00000000; // 3868 :   0 - 0x0
      13'hF1D: dout <= 8'b00000000; // 3869 :   0 - 0x0
      13'hF1E: dout <= 8'b00000000; // 3870 :   0 - 0x0
      13'hF1F: dout <= 8'b00000000; // 3871 :   0 - 0x0
      13'hF20: dout <= 8'b00000000; // 3872 :   0 - 0x0 -- Sprite 0xf2
      13'hF21: dout <= 8'b11000000; // 3873 : 192 - 0xc0
      13'hF22: dout <= 8'b00000000; // 3874 :   0 - 0x0
      13'hF23: dout <= 8'b00000000; // 3875 :   0 - 0x0
      13'hF24: dout <= 8'b00000000; // 3876 :   0 - 0x0
      13'hF25: dout <= 8'b00000000; // 3877 :   0 - 0x0
      13'hF26: dout <= 8'b00000000; // 3878 :   0 - 0x0
      13'hF27: dout <= 8'b00000000; // 3879 :   0 - 0x0
      13'hF28: dout <= 8'b11000000; // 3880 : 192 - 0xc0
      13'hF29: dout <= 8'b11000000; // 3881 : 192 - 0xc0
      13'hF2A: dout <= 8'b11000000; // 3882 : 192 - 0xc0
      13'hF2B: dout <= 8'b11000000; // 3883 : 192 - 0xc0
      13'hF2C: dout <= 8'b00000000; // 3884 :   0 - 0x0
      13'hF2D: dout <= 8'b00000000; // 3885 :   0 - 0x0
      13'hF2E: dout <= 8'b00000000; // 3886 :   0 - 0x0
      13'hF2F: dout <= 8'b00000000; // 3887 :   0 - 0x0
      13'hF30: dout <= 8'b00000000; // 3888 :   0 - 0x0 -- Sprite 0xf3
      13'hF31: dout <= 8'b11100000; // 3889 : 224 - 0xe0
      13'hF32: dout <= 8'b00000000; // 3890 :   0 - 0x0
      13'hF33: dout <= 8'b00000000; // 3891 :   0 - 0x0
      13'hF34: dout <= 8'b00000000; // 3892 :   0 - 0x0
      13'hF35: dout <= 8'b00000000; // 3893 :   0 - 0x0
      13'hF36: dout <= 8'b00000000; // 3894 :   0 - 0x0
      13'hF37: dout <= 8'b00000000; // 3895 :   0 - 0x0
      13'hF38: dout <= 8'b11100000; // 3896 : 224 - 0xe0
      13'hF39: dout <= 8'b11100000; // 3897 : 224 - 0xe0
      13'hF3A: dout <= 8'b11100000; // 3898 : 224 - 0xe0
      13'hF3B: dout <= 8'b11100000; // 3899 : 224 - 0xe0
      13'hF3C: dout <= 8'b00000000; // 3900 :   0 - 0x0
      13'hF3D: dout <= 8'b00000000; // 3901 :   0 - 0x0
      13'hF3E: dout <= 8'b00000000; // 3902 :   0 - 0x0
      13'hF3F: dout <= 8'b00000000; // 3903 :   0 - 0x0
      13'hF40: dout <= 8'b00000000; // 3904 :   0 - 0x0 -- Sprite 0xf4
      13'hF41: dout <= 8'b11110000; // 3905 : 240 - 0xf0
      13'hF42: dout <= 8'b00000000; // 3906 :   0 - 0x0
      13'hF43: dout <= 8'b00000000; // 3907 :   0 - 0x0
      13'hF44: dout <= 8'b00000000; // 3908 :   0 - 0x0
      13'hF45: dout <= 8'b00000000; // 3909 :   0 - 0x0
      13'hF46: dout <= 8'b00000000; // 3910 :   0 - 0x0
      13'hF47: dout <= 8'b00000000; // 3911 :   0 - 0x0
      13'hF48: dout <= 8'b11110000; // 3912 : 240 - 0xf0
      13'hF49: dout <= 8'b11110000; // 3913 : 240 - 0xf0
      13'hF4A: dout <= 8'b11110000; // 3914 : 240 - 0xf0
      13'hF4B: dout <= 8'b11110000; // 3915 : 240 - 0xf0
      13'hF4C: dout <= 8'b00000000; // 3916 :   0 - 0x0
      13'hF4D: dout <= 8'b00000000; // 3917 :   0 - 0x0
      13'hF4E: dout <= 8'b00000000; // 3918 :   0 - 0x0
      13'hF4F: dout <= 8'b00000000; // 3919 :   0 - 0x0
      13'hF50: dout <= 8'b00000000; // 3920 :   0 - 0x0 -- Sprite 0xf5
      13'hF51: dout <= 8'b11111000; // 3921 : 248 - 0xf8
      13'hF52: dout <= 8'b00000000; // 3922 :   0 - 0x0
      13'hF53: dout <= 8'b00000000; // 3923 :   0 - 0x0
      13'hF54: dout <= 8'b00000000; // 3924 :   0 - 0x0
      13'hF55: dout <= 8'b00000000; // 3925 :   0 - 0x0
      13'hF56: dout <= 8'b00000000; // 3926 :   0 - 0x0
      13'hF57: dout <= 8'b00000000; // 3927 :   0 - 0x0
      13'hF58: dout <= 8'b11111000; // 3928 : 248 - 0xf8
      13'hF59: dout <= 8'b11111000; // 3929 : 248 - 0xf8
      13'hF5A: dout <= 8'b11111000; // 3930 : 248 - 0xf8
      13'hF5B: dout <= 8'b11111000; // 3931 : 248 - 0xf8
      13'hF5C: dout <= 8'b00000000; // 3932 :   0 - 0x0
      13'hF5D: dout <= 8'b00000000; // 3933 :   0 - 0x0
      13'hF5E: dout <= 8'b00000000; // 3934 :   0 - 0x0
      13'hF5F: dout <= 8'b00000000; // 3935 :   0 - 0x0
      13'hF60: dout <= 8'b00000000; // 3936 :   0 - 0x0 -- Sprite 0xf6
      13'hF61: dout <= 8'b11111100; // 3937 : 252 - 0xfc
      13'hF62: dout <= 8'b00000000; // 3938 :   0 - 0x0
      13'hF63: dout <= 8'b00000000; // 3939 :   0 - 0x0
      13'hF64: dout <= 8'b00000000; // 3940 :   0 - 0x0
      13'hF65: dout <= 8'b00000000; // 3941 :   0 - 0x0
      13'hF66: dout <= 8'b00000000; // 3942 :   0 - 0x0
      13'hF67: dout <= 8'b00000000; // 3943 :   0 - 0x0
      13'hF68: dout <= 8'b11111100; // 3944 : 252 - 0xfc
      13'hF69: dout <= 8'b11111100; // 3945 : 252 - 0xfc
      13'hF6A: dout <= 8'b11111100; // 3946 : 252 - 0xfc
      13'hF6B: dout <= 8'b11111100; // 3947 : 252 - 0xfc
      13'hF6C: dout <= 8'b00000000; // 3948 :   0 - 0x0
      13'hF6D: dout <= 8'b00000000; // 3949 :   0 - 0x0
      13'hF6E: dout <= 8'b00000000; // 3950 :   0 - 0x0
      13'hF6F: dout <= 8'b00000000; // 3951 :   0 - 0x0
      13'hF70: dout <= 8'b00000000; // 3952 :   0 - 0x0 -- Sprite 0xf7
      13'hF71: dout <= 8'b11111110; // 3953 : 254 - 0xfe
      13'hF72: dout <= 8'b00000000; // 3954 :   0 - 0x0
      13'hF73: dout <= 8'b00000000; // 3955 :   0 - 0x0
      13'hF74: dout <= 8'b00000000; // 3956 :   0 - 0x0
      13'hF75: dout <= 8'b00000000; // 3957 :   0 - 0x0
      13'hF76: dout <= 8'b00000000; // 3958 :   0 - 0x0
      13'hF77: dout <= 8'b00000000; // 3959 :   0 - 0x0
      13'hF78: dout <= 8'b11111110; // 3960 : 254 - 0xfe
      13'hF79: dout <= 8'b11111110; // 3961 : 254 - 0xfe
      13'hF7A: dout <= 8'b11111110; // 3962 : 254 - 0xfe
      13'hF7B: dout <= 8'b11111110; // 3963 : 254 - 0xfe
      13'hF7C: dout <= 8'b00000000; // 3964 :   0 - 0x0
      13'hF7D: dout <= 8'b00000000; // 3965 :   0 - 0x0
      13'hF7E: dout <= 8'b00000000; // 3966 :   0 - 0x0
      13'hF7F: dout <= 8'b00000000; // 3967 :   0 - 0x0
      13'hF80: dout <= 8'b00000000; // 3968 :   0 - 0x0 -- Sprite 0xf8
      13'hF81: dout <= 8'b11111111; // 3969 : 255 - 0xff
      13'hF82: dout <= 8'b00000000; // 3970 :   0 - 0x0
      13'hF83: dout <= 8'b00000000; // 3971 :   0 - 0x0
      13'hF84: dout <= 8'b00000000; // 3972 :   0 - 0x0
      13'hF85: dout <= 8'b00000000; // 3973 :   0 - 0x0
      13'hF86: dout <= 8'b00000000; // 3974 :   0 - 0x0
      13'hF87: dout <= 8'b00000000; // 3975 :   0 - 0x0
      13'hF88: dout <= 8'b11111111; // 3976 : 255 - 0xff
      13'hF89: dout <= 8'b11111111; // 3977 : 255 - 0xff
      13'hF8A: dout <= 8'b11111111; // 3978 : 255 - 0xff
      13'hF8B: dout <= 8'b11111111; // 3979 : 255 - 0xff
      13'hF8C: dout <= 8'b00000000; // 3980 :   0 - 0x0
      13'hF8D: dout <= 8'b00000000; // 3981 :   0 - 0x0
      13'hF8E: dout <= 8'b00000000; // 3982 :   0 - 0x0
      13'hF8F: dout <= 8'b00000000; // 3983 :   0 - 0x0
      13'hF90: dout <= 8'b11111111; // 3984 : 255 - 0xff -- Sprite 0xf9
      13'hF91: dout <= 8'b11111111; // 3985 : 255 - 0xff
      13'hF92: dout <= 8'b11111111; // 3986 : 255 - 0xff
      13'hF93: dout <= 8'b11111111; // 3987 : 255 - 0xff
      13'hF94: dout <= 8'b10000000; // 3988 : 128 - 0x80
      13'hF95: dout <= 8'b10000000; // 3989 : 128 - 0x80
      13'hF96: dout <= 8'b11000000; // 3990 : 192 - 0xc0
      13'hF97: dout <= 8'b11000000; // 3991 : 192 - 0xc0
      13'hF98: dout <= 8'b00000000; // 3992 :   0 - 0x0
      13'hF99: dout <= 8'b00000000; // 3993 :   0 - 0x0
      13'hF9A: dout <= 8'b00000000; // 3994 :   0 - 0x0
      13'hF9B: dout <= 8'b00000000; // 3995 :   0 - 0x0
      13'hF9C: dout <= 8'b01111111; // 3996 : 127 - 0x7f
      13'hF9D: dout <= 8'b01000000; // 3997 :  64 - 0x40
      13'hF9E: dout <= 8'b01000000; // 3998 :  64 - 0x40
      13'hF9F: dout <= 8'b01000000; // 3999 :  64 - 0x40
      13'hFA0: dout <= 8'b11111111; // 4000 : 255 - 0xff -- Sprite 0xfa
      13'hFA1: dout <= 8'b11111111; // 4001 : 255 - 0xff
      13'hFA2: dout <= 8'b11111111; // 4002 : 255 - 0xff
      13'hFA3: dout <= 8'b11111111; // 4003 : 255 - 0xff
      13'hFA4: dout <= 8'b00000000; // 4004 :   0 - 0x0
      13'hFA5: dout <= 8'b00000000; // 4005 :   0 - 0x0
      13'hFA6: dout <= 8'b00000000; // 4006 :   0 - 0x0
      13'hFA7: dout <= 8'b00000000; // 4007 :   0 - 0x0
      13'hFA8: dout <= 8'b00000000; // 4008 :   0 - 0x0
      13'hFA9: dout <= 8'b00000000; // 4009 :   0 - 0x0
      13'hFAA: dout <= 8'b00000000; // 4010 :   0 - 0x0
      13'hFAB: dout <= 8'b00000000; // 4011 :   0 - 0x0
      13'hFAC: dout <= 8'b11111111; // 4012 : 255 - 0xff
      13'hFAD: dout <= 8'b00000000; // 4013 :   0 - 0x0
      13'hFAE: dout <= 8'b00000000; // 4014 :   0 - 0x0
      13'hFAF: dout <= 8'b00000000; // 4015 :   0 - 0x0
      13'hFB0: dout <= 8'b11111111; // 4016 : 255 - 0xff -- Sprite 0xfb
      13'hFB1: dout <= 8'b11111111; // 4017 : 255 - 0xff
      13'hFB2: dout <= 8'b11111111; // 4018 : 255 - 0xff
      13'hFB3: dout <= 8'b11111111; // 4019 : 255 - 0xff
      13'hFB4: dout <= 8'b00000001; // 4020 :   1 - 0x1
      13'hFB5: dout <= 8'b00000000; // 4021 :   0 - 0x0
      13'hFB6: dout <= 8'b00000010; // 4022 :   2 - 0x2
      13'hFB7: dout <= 8'b00000010; // 4023 :   2 - 0x2
      13'hFB8: dout <= 8'b00000000; // 4024 :   0 - 0x0
      13'hFB9: dout <= 8'b00000000; // 4025 :   0 - 0x0
      13'hFBA: dout <= 8'b00000000; // 4026 :   0 - 0x0
      13'hFBB: dout <= 8'b00000000; // 4027 :   0 - 0x0
      13'hFBC: dout <= 8'b11111110; // 4028 : 254 - 0xfe
      13'hFBD: dout <= 8'b00000010; // 4029 :   2 - 0x2
      13'hFBE: dout <= 8'b00000010; // 4030 :   2 - 0x2
      13'hFBF: dout <= 8'b00000010; // 4031 :   2 - 0x2
      13'hFC0: dout <= 8'b11000000; // 4032 : 192 - 0xc0 -- Sprite 0xfc
      13'hFC1: dout <= 8'b11000000; // 4033 : 192 - 0xc0
      13'hFC2: dout <= 8'b10000000; // 4034 : 128 - 0x80
      13'hFC3: dout <= 8'b10000000; // 4035 : 128 - 0x80
      13'hFC4: dout <= 8'b11000000; // 4036 : 192 - 0xc0
      13'hFC5: dout <= 8'b11111111; // 4037 : 255 - 0xff
      13'hFC6: dout <= 8'b11111111; // 4038 : 255 - 0xff
      13'hFC7: dout <= 8'b11111111; // 4039 : 255 - 0xff
      13'hFC8: dout <= 8'b01000000; // 4040 :  64 - 0x40
      13'hFC9: dout <= 8'b01000000; // 4041 :  64 - 0x40
      13'hFCA: dout <= 8'b01000000; // 4042 :  64 - 0x40
      13'hFCB: dout <= 8'b01111111; // 4043 : 127 - 0x7f
      13'hFCC: dout <= 8'b00000000; // 4044 :   0 - 0x0
      13'hFCD: dout <= 8'b00000000; // 4045 :   0 - 0x0
      13'hFCE: dout <= 8'b00000000; // 4046 :   0 - 0x0
      13'hFCF: dout <= 8'b00000000; // 4047 :   0 - 0x0
      13'hFD0: dout <= 8'b00000000; // 4048 :   0 - 0x0 -- Sprite 0xfd
      13'hFD1: dout <= 8'b00000000; // 4049 :   0 - 0x0
      13'hFD2: dout <= 8'b00000000; // 4050 :   0 - 0x0
      13'hFD3: dout <= 8'b00000000; // 4051 :   0 - 0x0
      13'hFD4: dout <= 8'b00000000; // 4052 :   0 - 0x0
      13'hFD5: dout <= 8'b11111111; // 4053 : 255 - 0xff
      13'hFD6: dout <= 8'b11111111; // 4054 : 255 - 0xff
      13'hFD7: dout <= 8'b11111111; // 4055 : 255 - 0xff
      13'hFD8: dout <= 8'b00000000; // 4056 :   0 - 0x0
      13'hFD9: dout <= 8'b00000000; // 4057 :   0 - 0x0
      13'hFDA: dout <= 8'b00000000; // 4058 :   0 - 0x0
      13'hFDB: dout <= 8'b11111111; // 4059 : 255 - 0xff
      13'hFDC: dout <= 8'b00000000; // 4060 :   0 - 0x0
      13'hFDD: dout <= 8'b00000000; // 4061 :   0 - 0x0
      13'hFDE: dout <= 8'b00000000; // 4062 :   0 - 0x0
      13'hFDF: dout <= 8'b00000000; // 4063 :   0 - 0x0
      13'hFE0: dout <= 8'b00000010; // 4064 :   2 - 0x2 -- Sprite 0xfe
      13'hFE1: dout <= 8'b00000010; // 4065 :   2 - 0x2
      13'hFE2: dout <= 8'b00000000; // 4066 :   0 - 0x0
      13'hFE3: dout <= 8'b00000000; // 4067 :   0 - 0x0
      13'hFE4: dout <= 8'b00000000; // 4068 :   0 - 0x0
      13'hFE5: dout <= 8'b11111111; // 4069 : 255 - 0xff
      13'hFE6: dout <= 8'b11111111; // 4070 : 255 - 0xff
      13'hFE7: dout <= 8'b11111111; // 4071 : 255 - 0xff
      13'hFE8: dout <= 8'b00000010; // 4072 :   2 - 0x2
      13'hFE9: dout <= 8'b00000010; // 4073 :   2 - 0x2
      13'hFEA: dout <= 8'b00000010; // 4074 :   2 - 0x2
      13'hFEB: dout <= 8'b11111110; // 4075 : 254 - 0xfe
      13'hFEC: dout <= 8'b00000000; // 4076 :   0 - 0x0
      13'hFED: dout <= 8'b00000000; // 4077 :   0 - 0x0
      13'hFEE: dout <= 8'b00000000; // 4078 :   0 - 0x0
      13'hFEF: dout <= 8'b00000000; // 4079 :   0 - 0x0
      13'hFF0: dout <= 8'b11111111; // 4080 : 255 - 0xff -- Sprite 0xff
      13'hFF1: dout <= 8'b11111111; // 4081 : 255 - 0xff
      13'hFF2: dout <= 8'b11111111; // 4082 : 255 - 0xff
      13'hFF3: dout <= 8'b11111111; // 4083 : 255 - 0xff
      13'hFF4: dout <= 8'b11111111; // 4084 : 255 - 0xff
      13'hFF5: dout <= 8'b11111111; // 4085 : 255 - 0xff
      13'hFF6: dout <= 8'b11111111; // 4086 : 255 - 0xff
      13'hFF7: dout <= 8'b11111111; // 4087 : 255 - 0xff
      13'hFF8: dout <= 8'b00000000; // 4088 :   0 - 0x0
      13'hFF9: dout <= 8'b00000000; // 4089 :   0 - 0x0
      13'hFFA: dout <= 8'b00000000; // 4090 :   0 - 0x0
      13'hFFB: dout <= 8'b00000000; // 4091 :   0 - 0x0
      13'hFFC: dout <= 8'b00000000; // 4092 :   0 - 0x0
      13'hFFD: dout <= 8'b00000000; // 4093 :   0 - 0x0
      13'hFFE: dout <= 8'b00000000; // 4094 :   0 - 0x0
      13'hFFF: dout <= 8'b00000000; // 4095 :   0 - 0x0
          // Pattern Table 1---------
      13'h1000: dout <= 8'b00000000; // 4096 :   0 - 0x0 -- Background 0x0
      13'h1001: dout <= 8'b00000000; // 4097 :   0 - 0x0
      13'h1002: dout <= 8'b00000000; // 4098 :   0 - 0x0
      13'h1003: dout <= 8'b00000000; // 4099 :   0 - 0x0
      13'h1004: dout <= 8'b00000000; // 4100 :   0 - 0x0
      13'h1005: dout <= 8'b00000000; // 4101 :   0 - 0x0
      13'h1006: dout <= 8'b00000000; // 4102 :   0 - 0x0
      13'h1007: dout <= 8'b00000000; // 4103 :   0 - 0x0
      13'h1008: dout <= 8'b00000101; // 4104 :   5 - 0x5
      13'h1009: dout <= 8'b01010101; // 4105 :  85 - 0x55
      13'h100A: dout <= 8'b01010101; // 4106 :  85 - 0x55
      13'h100B: dout <= 8'b01010000; // 4107 :  80 - 0x50
      13'h100C: dout <= 8'b00000000; // 4108 :   0 - 0x0
      13'h100D: dout <= 8'b00000000; // 4109 :   0 - 0x0
      13'h100E: dout <= 8'b00000000; // 4110 :   0 - 0x0
      13'h100F: dout <= 8'b00000000; // 4111 :   0 - 0x0
      13'h1010: dout <= 8'b00000101; // 4112 :   5 - 0x5 -- Background 0x1
      13'h1011: dout <= 8'b01010101; // 4113 :  85 - 0x55
      13'h1012: dout <= 8'b01010101; // 4114 :  85 - 0x55
      13'h1013: dout <= 8'b01010000; // 4115 :  80 - 0x50
      13'h1014: dout <= 8'b00000000; // 4116 :   0 - 0x0
      13'h1015: dout <= 8'b00000000; // 4117 :   0 - 0x0
      13'h1016: dout <= 8'b00000000; // 4118 :   0 - 0x0
      13'h1017: dout <= 8'b00000000; // 4119 :   0 - 0x0
      13'h1018: dout <= 8'b00000101; // 4120 :   5 - 0x5
      13'h1019: dout <= 8'b01010101; // 4121 :  85 - 0x55
      13'h101A: dout <= 8'b01010101; // 4122 :  85 - 0x55
      13'h101B: dout <= 8'b01010000; // 4123 :  80 - 0x50
      13'h101C: dout <= 8'b00000000; // 4124 :   0 - 0x0
      13'h101D: dout <= 8'b00000000; // 4125 :   0 - 0x0
      13'h101E: dout <= 8'b00000000; // 4126 :   0 - 0x0
      13'h101F: dout <= 8'b00000000; // 4127 :   0 - 0x0
      13'h1020: dout <= 8'b00000101; // 4128 :   5 - 0x5 -- Background 0x2
      13'h1021: dout <= 8'b01010000; // 4129 :  80 - 0x50
      13'h1022: dout <= 8'b00000101; // 4130 :   5 - 0x5
      13'h1023: dout <= 8'b01010000; // 4131 :  80 - 0x50
      13'h1024: dout <= 8'b00000000; // 4132 :   0 - 0x0
      13'h1025: dout <= 8'b00000000; // 4133 :   0 - 0x0
      13'h1026: dout <= 8'b00000000; // 4134 :   0 - 0x0
      13'h1027: dout <= 8'b00000000; // 4135 :   0 - 0x0
      13'h1028: dout <= 8'b00000101; // 4136 :   5 - 0x5
      13'h1029: dout <= 8'b01010000; // 4137 :  80 - 0x50
      13'h102A: dout <= 8'b00000101; // 4138 :   5 - 0x5
      13'h102B: dout <= 8'b01010000; // 4139 :  80 - 0x50
      13'h102C: dout <= 8'b00000000; // 4140 :   0 - 0x0
      13'h102D: dout <= 8'b00000000; // 4141 :   0 - 0x0
      13'h102E: dout <= 8'b00000000; // 4142 :   0 - 0x0
      13'h102F: dout <= 8'b00000000; // 4143 :   0 - 0x0
      13'h1030: dout <= 8'b00000101; // 4144 :   5 - 0x5 -- Background 0x3
      13'h1031: dout <= 8'b01010000; // 4145 :  80 - 0x50
      13'h1032: dout <= 8'b00000101; // 4146 :   5 - 0x5
      13'h1033: dout <= 8'b01010000; // 4147 :  80 - 0x50
      13'h1034: dout <= 8'b00000000; // 4148 :   0 - 0x0
      13'h1035: dout <= 8'b00000000; // 4149 :   0 - 0x0
      13'h1036: dout <= 8'b00000000; // 4150 :   0 - 0x0
      13'h1037: dout <= 8'b00000000; // 4151 :   0 - 0x0
      13'h1038: dout <= 8'b00000101; // 4152 :   5 - 0x5
      13'h1039: dout <= 8'b01010101; // 4153 :  85 - 0x55
      13'h103A: dout <= 8'b01010101; // 4154 :  85 - 0x55
      13'h103B: dout <= 8'b01010000; // 4155 :  80 - 0x50
      13'h103C: dout <= 8'b00000000; // 4156 :   0 - 0x0
      13'h103D: dout <= 8'b00000000; // 4157 :   0 - 0x0
      13'h103E: dout <= 8'b00000000; // 4158 :   0 - 0x0
      13'h103F: dout <= 8'b00000000; // 4159 :   0 - 0x0
      13'h1040: dout <= 8'b00000101; // 4160 :   5 - 0x5 -- Background 0x4
      13'h1041: dout <= 8'b01010101; // 4161 :  85 - 0x55
      13'h1042: dout <= 8'b01010101; // 4162 :  85 - 0x55
      13'h1043: dout <= 8'b01010000; // 4163 :  80 - 0x50
      13'h1044: dout <= 8'b00000000; // 4164 :   0 - 0x0
      13'h1045: dout <= 8'b00000000; // 4165 :   0 - 0x0
      13'h1046: dout <= 8'b00000000; // 4166 :   0 - 0x0
      13'h1047: dout <= 8'b00000000; // 4167 :   0 - 0x0
      13'h1048: dout <= 8'b00000101; // 4168 :   5 - 0x5
      13'h1049: dout <= 8'b01010101; // 4169 :  85 - 0x55
      13'h104A: dout <= 8'b01010101; // 4170 :  85 - 0x55
      13'h104B: dout <= 8'b01010000; // 4171 :  80 - 0x50
      13'h104C: dout <= 8'b00000000; // 4172 :   0 - 0x0
      13'h104D: dout <= 8'b00000000; // 4173 :   0 - 0x0
      13'h104E: dout <= 8'b00000000; // 4174 :   0 - 0x0
      13'h104F: dout <= 8'b00000000; // 4175 :   0 - 0x0
      13'h1050: dout <= 8'b00000000; // 4176 :   0 - 0x0 -- Background 0x5
      13'h1051: dout <= 8'b00000000; // 4177 :   0 - 0x0
      13'h1052: dout <= 8'b00000000; // 4178 :   0 - 0x0
      13'h1053: dout <= 8'b00000000; // 4179 :   0 - 0x0
      13'h1054: dout <= 8'b00000000; // 4180 :   0 - 0x0
      13'h1055: dout <= 8'b00000000; // 4181 :   0 - 0x0
      13'h1056: dout <= 8'b00000000; // 4182 :   0 - 0x0
      13'h1057: dout <= 8'b00000000; // 4183 :   0 - 0x0
      13'h1058: dout <= 8'b00001110; // 4184 :  14 - 0xe
      13'h1059: dout <= 8'b00000111; // 4185 :   7 - 0x7
      13'h105A: dout <= 8'b00001000; // 4186 :   8 - 0x8
      13'h105B: dout <= 8'b01100000; // 4187 :  96 - 0x60
      13'h105C: dout <= 8'b00000000; // 4188 :   0 - 0x0
      13'h105D: dout <= 8'b00001010; // 4189 :  10 - 0xa
      13'h105E: dout <= 8'b00000001; // 4190 :   1 - 0x1
      13'h105F: dout <= 8'b00010101; // 4191 :  21 - 0x15
      13'h1060: dout <= 8'b01010101; // 4192 :  85 - 0x55 -- Background 0x6
      13'h1061: dout <= 8'b01010101; // 4193 :  85 - 0x55
      13'h1062: dout <= 8'b01010100; // 4194 :  84 - 0x54
      13'h1063: dout <= 8'b00000000; // 4195 :   0 - 0x0
      13'h1064: dout <= 8'b00000000; // 4196 :   0 - 0x0
      13'h1065: dout <= 8'b00000000; // 4197 :   0 - 0x0
      13'h1066: dout <= 8'b00000000; // 4198 :   0 - 0x0
      13'h1067: dout <= 8'b00010101; // 4199 :  21 - 0x15
      13'h1068: dout <= 8'b01010101; // 4200 :  85 - 0x55
      13'h1069: dout <= 8'b01010101; // 4201 :  85 - 0x55
      13'h106A: dout <= 8'b01010100; // 4202 :  84 - 0x54
      13'h106B: dout <= 8'b00000000; // 4203 :   0 - 0x0
      13'h106C: dout <= 8'b00000000; // 4204 :   0 - 0x0
      13'h106D: dout <= 8'b00000000; // 4205 :   0 - 0x0
      13'h106E: dout <= 8'b00000000; // 4206 :   0 - 0x0
      13'h106F: dout <= 8'b00010110; // 4207 :  22 - 0x16
      13'h1070: dout <= 8'b10101010; // 4208 : 170 - 0xaa -- Background 0x7
      13'h1071: dout <= 8'b10011010; // 4209 : 154 - 0x9a
      13'h1072: dout <= 8'b10010100; // 4210 : 148 - 0x94
      13'h1073: dout <= 8'b00000000; // 4211 :   0 - 0x0
      13'h1074: dout <= 8'b00000000; // 4212 :   0 - 0x0
      13'h1075: dout <= 8'b00000000; // 4213 :   0 - 0x0
      13'h1076: dout <= 8'b00000000; // 4214 :   0 - 0x0
      13'h1077: dout <= 8'b00010110; // 4215 :  22 - 0x16
      13'h1078: dout <= 8'b01010101; // 4216 :  85 - 0x55
      13'h1079: dout <= 8'b01010101; // 4217 :  85 - 0x55
      13'h107A: dout <= 8'b10010100; // 4218 : 148 - 0x94
      13'h107B: dout <= 8'b00000000; // 4219 :   0 - 0x0
      13'h107C: dout <= 8'b00000000; // 4220 :   0 - 0x0
      13'h107D: dout <= 8'b00000000; // 4221 :   0 - 0x0
      13'h107E: dout <= 8'b00000000; // 4222 :   0 - 0x0
      13'h107F: dout <= 8'b00010110; // 4223 :  22 - 0x16
      13'h1080: dout <= 8'b01010000; // 4224 :  80 - 0x50 -- Background 0x8
      13'h1081: dout <= 8'b00000101; // 4225 :   5 - 0x5
      13'h1082: dout <= 8'b10010100; // 4226 : 148 - 0x94
      13'h1083: dout <= 8'b00000000; // 4227 :   0 - 0x0
      13'h1084: dout <= 8'b00000000; // 4228 :   0 - 0x0
      13'h1085: dout <= 8'b00000000; // 4229 :   0 - 0x0
      13'h1086: dout <= 8'b00000000; // 4230 :   0 - 0x0
      13'h1087: dout <= 8'b00010101; // 4231 :  21 - 0x15
      13'h1088: dout <= 8'b01010000; // 4232 :  80 - 0x50
      13'h1089: dout <= 8'b00000101; // 4233 :   5 - 0x5
      13'h108A: dout <= 8'b01010100; // 4234 :  84 - 0x54
      13'h108B: dout <= 8'b00000000; // 4235 :   0 - 0x0
      13'h108C: dout <= 8'b00000000; // 4236 :   0 - 0x0
      13'h108D: dout <= 8'b00000000; // 4237 :   0 - 0x0
      13'h108E: dout <= 8'b00000000; // 4238 :   0 - 0x0
      13'h108F: dout <= 8'b00010110; // 4239 :  22 - 0x16
      13'h1090: dout <= 8'b01010000; // 4240 :  80 - 0x50 -- Background 0x9
      13'h1091: dout <= 8'b00000101; // 4241 :   5 - 0x5
      13'h1092: dout <= 8'b10010100; // 4242 : 148 - 0x94
      13'h1093: dout <= 8'b00000000; // 4243 :   0 - 0x0
      13'h1094: dout <= 8'b00000000; // 4244 :   0 - 0x0
      13'h1095: dout <= 8'b00000000; // 4245 :   0 - 0x0
      13'h1096: dout <= 8'b00000000; // 4246 :   0 - 0x0
      13'h1097: dout <= 8'b00010110; // 4247 :  22 - 0x16
      13'h1098: dout <= 8'b01010101; // 4248 :  85 - 0x55
      13'h1099: dout <= 8'b01010101; // 4249 :  85 - 0x55
      13'h109A: dout <= 8'b10010100; // 4250 : 148 - 0x94
      13'h109B: dout <= 8'b00000000; // 4251 :   0 - 0x0
      13'h109C: dout <= 8'b00000000; // 4252 :   0 - 0x0
      13'h109D: dout <= 8'b00000000; // 4253 :   0 - 0x0
      13'h109E: dout <= 8'b00000000; // 4254 :   0 - 0x0
      13'h109F: dout <= 8'b00010110; // 4255 :  22 - 0x16
      13'h10A0: dout <= 8'b10100110; // 4256 : 166 - 0xa6 -- Background 0xa
      13'h10A1: dout <= 8'b10101010; // 4257 : 170 - 0xaa
      13'h10A2: dout <= 8'b10010100; // 4258 : 148 - 0x94
      13'h10A3: dout <= 8'b00000000; // 4259 :   0 - 0x0
      13'h10A4: dout <= 8'b00000000; // 4260 :   0 - 0x0
      13'h10A5: dout <= 8'b00000000; // 4261 :   0 - 0x0
      13'h10A6: dout <= 8'b00000000; // 4262 :   0 - 0x0
      13'h10A7: dout <= 8'b00010101; // 4263 :  21 - 0x15
      13'h10A8: dout <= 8'b01010101; // 4264 :  85 - 0x55
      13'h10A9: dout <= 8'b01010101; // 4265 :  85 - 0x55
      13'h10AA: dout <= 8'b01010100; // 4266 :  84 - 0x54
      13'h10AB: dout <= 8'b00000000; // 4267 :   0 - 0x0
      13'h10AC: dout <= 8'b00000000; // 4268 :   0 - 0x0
      13'h10AD: dout <= 8'b00000000; // 4269 :   0 - 0x0
      13'h10AE: dout <= 8'b00000000; // 4270 :   0 - 0x0
      13'h10AF: dout <= 8'b00010101; // 4271 :  21 - 0x15
      13'h10B0: dout <= 8'b01010101; // 4272 :  85 - 0x55 -- Background 0xb
      13'h10B1: dout <= 8'b01010101; // 4273 :  85 - 0x55
      13'h10B2: dout <= 8'b01010100; // 4274 :  84 - 0x54
      13'h10B3: dout <= 8'b00000000; // 4275 :   0 - 0x0
      13'h10B4: dout <= 8'b00000000; // 4276 :   0 - 0x0
      13'h10B5: dout <= 8'b00000000; // 4277 :   0 - 0x0
      13'h10B6: dout <= 8'b00000000; // 4278 :   0 - 0x0
      13'h10B7: dout <= 8'b00001110; // 4279 :  14 - 0xe
      13'h10B8: dout <= 8'b00000111; // 4280 :   7 - 0x7
      13'h10B9: dout <= 8'b00001000; // 4281 :   8 - 0x8
      13'h10BA: dout <= 8'b01110100; // 4282 : 116 - 0x74
      13'h10BB: dout <= 8'b00000000; // 4283 :   0 - 0x0
      13'h10BC: dout <= 8'b11011100; // 4284 : 220 - 0xdc
      13'h10BD: dout <= 8'b00000000; // 4285 :   0 - 0x0
      13'h10BE: dout <= 8'b00010101; // 4286 :  21 - 0x15
      13'h10BF: dout <= 8'b01010101; // 4287 :  85 - 0x55
      13'h10C0: dout <= 8'b01010101; // 4288 :  85 - 0x55 -- Background 0xc
      13'h10C1: dout <= 8'b01010100; // 4289 :  84 - 0x54
      13'h10C2: dout <= 8'b00000000; // 4290 :   0 - 0x0
      13'h10C3: dout <= 8'b00000000; // 4291 :   0 - 0x0
      13'h10C4: dout <= 8'b00000000; // 4292 :   0 - 0x0
      13'h10C5: dout <= 8'b00000000; // 4293 :   0 - 0x0
      13'h10C6: dout <= 8'b00011010; // 4294 :  26 - 0x1a
      13'h10C7: dout <= 8'b10011101; // 4295 : 157 - 0x9d
      13'h10C8: dout <= 8'b01110110; // 4296 : 118 - 0x76
      13'h10C9: dout <= 8'b10100100; // 4297 : 164 - 0xa4
      13'h10CA: dout <= 8'b00000000; // 4298 :   0 - 0x0
      13'h10CB: dout <= 8'b00000000; // 4299 :   0 - 0x0
      13'h10CC: dout <= 8'b00000000; // 4300 :   0 - 0x0
      13'h10CD: dout <= 8'b00000000; // 4301 :   0 - 0x0
      13'h10CE: dout <= 8'b00010101; // 4302 :  21 - 0x15
      13'h10CF: dout <= 8'b01010101; // 4303 :  85 - 0x55
      13'h10D0: dout <= 8'b01010101; // 4304 :  85 - 0x55 -- Background 0xd
      13'h10D1: dout <= 8'b01010100; // 4305 :  84 - 0x54
      13'h10D2: dout <= 8'b00000000; // 4306 :   0 - 0x0
      13'h10D3: dout <= 8'b00000000; // 4307 :   0 - 0x0
      13'h10D4: dout <= 8'b00000000; // 4308 :   0 - 0x0
      13'h10D5: dout <= 8'b00000000; // 4309 :   0 - 0x0
      13'h10D6: dout <= 8'b00010111; // 4310 :  23 - 0x17
      13'h10D7: dout <= 8'b01010101; // 4311 :  85 - 0x55
      13'h10D8: dout <= 8'b01010101; // 4312 :  85 - 0x55
      13'h10D9: dout <= 8'b11010100; // 4313 : 212 - 0xd4
      13'h10DA: dout <= 8'b00000000; // 4314 :   0 - 0x0
      13'h10DB: dout <= 8'b00000000; // 4315 :   0 - 0x0
      13'h10DC: dout <= 8'b00000000; // 4316 :   0 - 0x0
      13'h10DD: dout <= 8'b00000000; // 4317 :   0 - 0x0
      13'h10DE: dout <= 8'b00010101; // 4318 :  21 - 0x15
      13'h10DF: dout <= 8'b01010000; // 4319 :  80 - 0x50
      13'h10E0: dout <= 8'b00000101; // 4320 :   5 - 0x5 -- Background 0xe
      13'h10E1: dout <= 8'b01010100; // 4321 :  84 - 0x54
      13'h10E2: dout <= 8'b00000000; // 4322 :   0 - 0x0
      13'h10E3: dout <= 8'b00000000; // 4323 :   0 - 0x0
      13'h10E4: dout <= 8'b00000000; // 4324 :   0 - 0x0
      13'h10E5: dout <= 8'b00000000; // 4325 :   0 - 0x0
      13'h10E6: dout <= 8'b00010101; // 4326 :  21 - 0x15
      13'h10E7: dout <= 8'b01010000; // 4327 :  80 - 0x50
      13'h10E8: dout <= 8'b00000101; // 4328 :   5 - 0x5
      13'h10E9: dout <= 8'b01010100; // 4329 :  84 - 0x54
      13'h10EA: dout <= 8'b00000000; // 4330 :   0 - 0x0
      13'h10EB: dout <= 8'b00000000; // 4331 :   0 - 0x0
      13'h10EC: dout <= 8'b00000000; // 4332 :   0 - 0x0
      13'h10ED: dout <= 8'b00000000; // 4333 :   0 - 0x0
      13'h10EE: dout <= 8'b00010101; // 4334 :  21 - 0x15
      13'h10EF: dout <= 8'b01010000; // 4335 :  80 - 0x50
      13'h10F0: dout <= 8'b00000101; // 4336 :   5 - 0x5 -- Background 0xf
      13'h10F1: dout <= 8'b01010100; // 4337 :  84 - 0x54
      13'h10F2: dout <= 8'b00000000; // 4338 :   0 - 0x0
      13'h10F3: dout <= 8'b00000000; // 4339 :   0 - 0x0
      13'h10F4: dout <= 8'b00000000; // 4340 :   0 - 0x0
      13'h10F5: dout <= 8'b00000000; // 4341 :   0 - 0x0
      13'h10F6: dout <= 8'b00010111; // 4342 :  23 - 0x17
      13'h10F7: dout <= 8'b01010101; // 4343 :  85 - 0x55
      13'h10F8: dout <= 8'b01010101; // 4344 :  85 - 0x55
      13'h10F9: dout <= 8'b11010100; // 4345 : 212 - 0xd4
      13'h10FA: dout <= 8'b00000000; // 4346 :   0 - 0x0
      13'h10FB: dout <= 8'b00000000; // 4347 :   0 - 0x0
      13'h10FC: dout <= 8'b00000000; // 4348 :   0 - 0x0
      13'h10FD: dout <= 8'b00000000; // 4349 :   0 - 0x0
      13'h10FE: dout <= 8'b00010101; // 4350 :  21 - 0x15
      13'h10FF: dout <= 8'b01010101; // 4351 :  85 - 0x55
      13'h1100: dout <= 8'b01010101; // 4352 :  85 - 0x55 -- Background 0x10
      13'h1101: dout <= 8'b01010100; // 4353 :  84 - 0x54
      13'h1102: dout <= 8'b00000000; // 4354 :   0 - 0x0
      13'h1103: dout <= 8'b00000000; // 4355 :   0 - 0x0
      13'h1104: dout <= 8'b00000000; // 4356 :   0 - 0x0
      13'h1105: dout <= 8'b00000000; // 4357 :   0 - 0x0
      13'h1106: dout <= 8'b00011010; // 4358 :  26 - 0x1a
      13'h1107: dout <= 8'b10011101; // 4359 : 157 - 0x9d
      13'h1108: dout <= 8'b01110110; // 4360 : 118 - 0x76
      13'h1109: dout <= 8'b10100100; // 4361 : 164 - 0xa4
      13'h110A: dout <= 8'b00000000; // 4362 :   0 - 0x0
      13'h110B: dout <= 8'b00000000; // 4363 :   0 - 0x0
      13'h110C: dout <= 8'b00000000; // 4364 :   0 - 0x0
      13'h110D: dout <= 8'b00000000; // 4365 :   0 - 0x0
      13'h110E: dout <= 8'b00010101; // 4366 :  21 - 0x15
      13'h110F: dout <= 8'b01010101; // 4367 :  85 - 0x55
      13'h1110: dout <= 8'b01010101; // 4368 :  85 - 0x55 -- Background 0x11
      13'h1111: dout <= 8'b01010100; // 4369 :  84 - 0x54
      13'h1112: dout <= 8'b00000000; // 4370 :   0 - 0x0
      13'h1113: dout <= 8'b00000000; // 4371 :   0 - 0x0
      13'h1114: dout <= 8'b00000000; // 4372 :   0 - 0x0
      13'h1115: dout <= 8'b00000000; // 4373 :   0 - 0x0
      13'h1116: dout <= 8'b00001110; // 4374 :  14 - 0xe
      13'h1117: dout <= 8'b00000111; // 4375 :   7 - 0x7
      13'h1118: dout <= 8'b00001000; // 4376 :   8 - 0x8
      13'h1119: dout <= 8'b01111010; // 4377 : 122 - 0x7a
      13'h111A: dout <= 8'b00000000; // 4378 :   0 - 0x0
      13'h111B: dout <= 8'b11010001; // 4379 : 209 - 0xd1
      13'h111C: dout <= 8'b00000000; // 4380 :   0 - 0x0
      13'h111D: dout <= 8'b00010101; // 4381 :  21 - 0x15
      13'h111E: dout <= 8'b01010101; // 4382 :  85 - 0x55
      13'h111F: dout <= 8'b01010101; // 4383 :  85 - 0x55
      13'h1120: dout <= 8'b01010101; // 4384 :  85 - 0x55 -- Background 0x12
      13'h1121: dout <= 8'b01010101; // 4385 :  85 - 0x55
      13'h1122: dout <= 8'b01000000; // 4386 :  64 - 0x40
      13'h1123: dout <= 8'b00000000; // 4387 :   0 - 0x0
      13'h1124: dout <= 8'b00000000; // 4388 :   0 - 0x0
      13'h1125: dout <= 8'b00010101; // 4389 :  21 - 0x15
      13'h1126: dout <= 8'b01010101; // 4390 :  85 - 0x55
      13'h1127: dout <= 8'b01010101; // 4391 :  85 - 0x55
      13'h1128: dout <= 8'b01010101; // 4392 :  85 - 0x55
      13'h1129: dout <= 8'b01010101; // 4393 :  85 - 0x55
      13'h112A: dout <= 8'b01000000; // 4394 :  64 - 0x40
      13'h112B: dout <= 8'b00000000; // 4395 :   0 - 0x0
      13'h112C: dout <= 8'b00000000; // 4396 :   0 - 0x0
      13'h112D: dout <= 8'b00010110; // 4397 :  22 - 0x16
      13'h112E: dout <= 8'b10100101; // 4398 : 165 - 0xa5
      13'h112F: dout <= 8'b01010101; // 4399 :  85 - 0x55
      13'h1130: dout <= 8'b01010101; // 4400 :  85 - 0x55 -- Background 0x13
      13'h1131: dout <= 8'b10101001; // 4401 : 169 - 0xa9
      13'h1132: dout <= 8'b01000000; // 4402 :  64 - 0x40
      13'h1133: dout <= 8'b00000000; // 4403 :   0 - 0x0
      13'h1134: dout <= 8'b00000000; // 4404 :   0 - 0x0
      13'h1135: dout <= 8'b00010110; // 4405 :  22 - 0x16
      13'h1136: dout <= 8'b01010101; // 4406 :  85 - 0x55
      13'h1137: dout <= 8'b01101010; // 4407 : 106 - 0x6a
      13'h1138: dout <= 8'b10010101; // 4408 : 149 - 0x95
      13'h1139: dout <= 8'b01011001; // 4409 :  89 - 0x59
      13'h113A: dout <= 8'b01000000; // 4410 :  64 - 0x40
      13'h113B: dout <= 8'b00000000; // 4411 :   0 - 0x0
      13'h113C: dout <= 8'b00000000; // 4412 :   0 - 0x0
      13'h113D: dout <= 8'b00010110; // 4413 :  22 - 0x16
      13'h113E: dout <= 8'b01000000; // 4414 :  64 - 0x40
      13'h113F: dout <= 8'b01010101; // 4415 :  85 - 0x55
      13'h1140: dout <= 8'b01010101; // 4416 :  85 - 0x55 -- Background 0x14
      13'h1141: dout <= 8'b01011001; // 4417 :  89 - 0x59
      13'h1142: dout <= 8'b01000000; // 4418 :  64 - 0x40
      13'h1143: dout <= 8'b00000000; // 4419 :   0 - 0x0
      13'h1144: dout <= 8'b00000000; // 4420 :   0 - 0x0
      13'h1145: dout <= 8'b00010101; // 4421 :  21 - 0x15
      13'h1146: dout <= 8'b01000000; // 4422 :  64 - 0x40
      13'h1147: dout <= 8'b01010101; // 4423 :  85 - 0x55
      13'h1148: dout <= 8'b01010101; // 4424 :  85 - 0x55
      13'h1149: dout <= 8'b01010101; // 4425 :  85 - 0x55
      13'h114A: dout <= 8'b01000000; // 4426 :  64 - 0x40
      13'h114B: dout <= 8'b00000000; // 4427 :   0 - 0x0
      13'h114C: dout <= 8'b00000000; // 4428 :   0 - 0x0
      13'h114D: dout <= 8'b00010110; // 4429 :  22 - 0x16
      13'h114E: dout <= 8'b01000000; // 4430 :  64 - 0x40
      13'h114F: dout <= 8'b01010101; // 4431 :  85 - 0x55
      13'h1150: dout <= 8'b01010101; // 4432 :  85 - 0x55 -- Background 0x15
      13'h1151: dout <= 8'b01011001; // 4433 :  89 - 0x59
      13'h1152: dout <= 8'b01000000; // 4434 :  64 - 0x40
      13'h1153: dout <= 8'b00000000; // 4435 :   0 - 0x0
      13'h1154: dout <= 8'b00000000; // 4436 :   0 - 0x0
      13'h1155: dout <= 8'b00010110; // 4437 :  22 - 0x16
      13'h1156: dout <= 8'b01010101; // 4438 :  85 - 0x55
      13'h1157: dout <= 8'b01101010; // 4439 : 106 - 0x6a
      13'h1158: dout <= 8'b10010101; // 4440 : 149 - 0x95
      13'h1159: dout <= 8'b01011001; // 4441 :  89 - 0x59
      13'h115A: dout <= 8'b01000000; // 4442 :  64 - 0x40
      13'h115B: dout <= 8'b00000000; // 4443 :   0 - 0x0
      13'h115C: dout <= 8'b00000000; // 4444 :   0 - 0x0
      13'h115D: dout <= 8'b00010110; // 4445 :  22 - 0x16
      13'h115E: dout <= 8'b10100101; // 4446 : 165 - 0xa5
      13'h115F: dout <= 8'b01010101; // 4447 :  85 - 0x55
      13'h1160: dout <= 8'b01010101; // 4448 :  85 - 0x55 -- Background 0x16
      13'h1161: dout <= 8'b10101001; // 4449 : 169 - 0xa9
      13'h1162: dout <= 8'b01000000; // 4450 :  64 - 0x40
      13'h1163: dout <= 8'b00000000; // 4451 :   0 - 0x0
      13'h1164: dout <= 8'b00000000; // 4452 :   0 - 0x0
      13'h1165: dout <= 8'b00010101; // 4453 :  21 - 0x15
      13'h1166: dout <= 8'b01010101; // 4454 :  85 - 0x55
      13'h1167: dout <= 8'b01010101; // 4455 :  85 - 0x55
      13'h1168: dout <= 8'b01010101; // 4456 :  85 - 0x55
      13'h1169: dout <= 8'b01010101; // 4457 :  85 - 0x55
      13'h116A: dout <= 8'b01000000; // 4458 :  64 - 0x40
      13'h116B: dout <= 8'b00000000; // 4459 :   0 - 0x0
      13'h116C: dout <= 8'b00000000; // 4460 :   0 - 0x0
      13'h116D: dout <= 8'b00010101; // 4461 :  21 - 0x15
      13'h116E: dout <= 8'b01010101; // 4462 :  85 - 0x55
      13'h116F: dout <= 8'b01010101; // 4463 :  85 - 0x55
      13'h1170: dout <= 8'b01010101; // 4464 :  85 - 0x55 -- Background 0x17
      13'h1171: dout <= 8'b01010101; // 4465 :  85 - 0x55
      13'h1172: dout <= 8'b01000000; // 4466 :  64 - 0x40
      13'h1173: dout <= 8'b00000000; // 4467 :   0 - 0x0
      13'h1174: dout <= 8'b00000000; // 4468 :   0 - 0x0
      13'h1175: dout <= 8'b00010100; // 4469 :  20 - 0x14
      13'h1176: dout <= 8'b00000110; // 4470 :   6 - 0x6
      13'h1177: dout <= 8'b00001000; // 4471 :   8 - 0x8
      13'h1178: dout <= 8'b10110111; // 4472 : 183 - 0xb7
      13'h1179: dout <= 8'b00000000; // 4473 :   0 - 0x0
      13'h117A: dout <= 8'b10001011; // 4474 : 139 - 0x8b
      13'h117B: dout <= 8'b00000000; // 4475 :   0 - 0x0
      13'h117C: dout <= 8'b00010101; // 4476 :  21 - 0x15
      13'h117D: dout <= 8'b01010101; // 4477 :  85 - 0x55
      13'h117E: dout <= 8'b01010101; // 4478 :  85 - 0x55
      13'h117F: dout <= 8'b01010101; // 4479 :  85 - 0x55
      13'h1180: dout <= 8'b01010101; // 4480 :  85 - 0x55 -- Background 0x18
      13'h1181: dout <= 8'b01000000; // 4481 :  64 - 0x40
      13'h1182: dout <= 8'b00000000; // 4482 :   0 - 0x0
      13'h1183: dout <= 8'b00000000; // 4483 :   0 - 0x0
      13'h1184: dout <= 8'b00011010; // 4484 :  26 - 0x1a
      13'h1185: dout <= 8'b01010111; // 4485 :  87 - 0x57
      13'h1186: dout <= 8'b01010101; // 4486 :  85 - 0x55
      13'h1187: dout <= 8'b01011101; // 4487 :  93 - 0x5d
      13'h1188: dout <= 8'b01011010; // 4488 :  90 - 0x5a
      13'h1189: dout <= 8'b01000000; // 4489 :  64 - 0x40
      13'h118A: dout <= 8'b00000000; // 4490 :   0 - 0x0
      13'h118B: dout <= 8'b00000000; // 4491 :   0 - 0x0
      13'h118C: dout <= 8'b00011010; // 4492 :  26 - 0x1a
      13'h118D: dout <= 8'b01010111; // 4493 :  87 - 0x57
      13'h118E: dout <= 8'b01010101; // 4494 :  85 - 0x55
      13'h118F: dout <= 8'b01011101; // 4495 :  93 - 0x5d
      13'h1190: dout <= 8'b01011010; // 4496 :  90 - 0x5a -- Background 0x19
      13'h1191: dout <= 8'b01000000; // 4497 :  64 - 0x40
      13'h1192: dout <= 8'b00000000; // 4498 :   0 - 0x0
      13'h1193: dout <= 8'b00000000; // 4499 :   0 - 0x0
      13'h1194: dout <= 8'b00010101; // 4500 :  21 - 0x15
      13'h1195: dout <= 8'b01010111; // 4501 :  87 - 0x57
      13'h1196: dout <= 8'b01011010; // 4502 :  90 - 0x5a
      13'h1197: dout <= 8'b01011101; // 4503 :  93 - 0x5d
      13'h1198: dout <= 8'b01010101; // 4504 :  85 - 0x55
      13'h1199: dout <= 8'b01000000; // 4505 :  64 - 0x40
      13'h119A: dout <= 8'b00000000; // 4506 :   0 - 0x0
      13'h119B: dout <= 8'b00000000; // 4507 :   0 - 0x0
      13'h119C: dout <= 8'b00010000; // 4508 :  16 - 0x10
      13'h119D: dout <= 8'b00010101; // 4509 :  21 - 0x15
      13'h119E: dout <= 8'b01011010; // 4510 :  90 - 0x5a
      13'h119F: dout <= 8'b01010101; // 4511 :  85 - 0x55
      13'h11A0: dout <= 8'b01010101; // 4512 :  85 - 0x55 -- Background 0x1a
      13'h11A1: dout <= 8'b01000000; // 4513 :  64 - 0x40
      13'h11A2: dout <= 8'b00000000; // 4514 :   0 - 0x0
      13'h11A3: dout <= 8'b00000000; // 4515 :   0 - 0x0
      13'h11A4: dout <= 8'b00010000; // 4516 :  16 - 0x10
      13'h11A5: dout <= 8'b00010101; // 4517 :  21 - 0x15
      13'h11A6: dout <= 8'b01011010; // 4518 :  90 - 0x5a
      13'h11A7: dout <= 8'b01010101; // 4519 :  85 - 0x55
      13'h11A8: dout <= 8'b01010101; // 4520 :  85 - 0x55
      13'h11A9: dout <= 8'b01000000; // 4521 :  64 - 0x40
      13'h11AA: dout <= 8'b00000000; // 4522 :   0 - 0x0
      13'h11AB: dout <= 8'b00000000; // 4523 :   0 - 0x0
      13'h11AC: dout <= 8'b00010000; // 4524 :  16 - 0x10
      13'h11AD: dout <= 8'b00010101; // 4525 :  21 - 0x15
      13'h11AE: dout <= 8'b01011010; // 4526 :  90 - 0x5a
      13'h11AF: dout <= 8'b01010101; // 4527 :  85 - 0x55
      13'h11B0: dout <= 8'b01010101; // 4528 :  85 - 0x55 -- Background 0x1b
      13'h11B1: dout <= 8'b01000000; // 4529 :  64 - 0x40
      13'h11B2: dout <= 8'b00000000; // 4530 :   0 - 0x0
      13'h11B3: dout <= 8'b00000000; // 4531 :   0 - 0x0
      13'h11B4: dout <= 8'b00010101; // 4532 :  21 - 0x15
      13'h11B5: dout <= 8'b01010111; // 4533 :  87 - 0x57
      13'h11B6: dout <= 8'b01011010; // 4534 :  90 - 0x5a
      13'h11B7: dout <= 8'b01011101; // 4535 :  93 - 0x5d
      13'h11B8: dout <= 8'b01010101; // 4536 :  85 - 0x55
      13'h11B9: dout <= 8'b01000000; // 4537 :  64 - 0x40
      13'h11BA: dout <= 8'b00000000; // 4538 :   0 - 0x0
      13'h11BB: dout <= 8'b00000000; // 4539 :   0 - 0x0
      13'h11BC: dout <= 8'b00011010; // 4540 :  26 - 0x1a
      13'h11BD: dout <= 8'b01010111; // 4541 :  87 - 0x57
      13'h11BE: dout <= 8'b01010101; // 4542 :  85 - 0x55
      13'h11BF: dout <= 8'b01011101; // 4543 :  93 - 0x5d
      13'h11C0: dout <= 8'b01011010; // 4544 :  90 - 0x5a -- Background 0x1c
      13'h11C1: dout <= 8'b01000000; // 4545 :  64 - 0x40
      13'h11C2: dout <= 8'b00000000; // 4546 :   0 - 0x0
      13'h11C3: dout <= 8'b00000000; // 4547 :   0 - 0x0
      13'h11C4: dout <= 8'b00011010; // 4548 :  26 - 0x1a
      13'h11C5: dout <= 8'b01010111; // 4549 :  87 - 0x57
      13'h11C6: dout <= 8'b01010101; // 4550 :  85 - 0x55
      13'h11C7: dout <= 8'b01011101; // 4551 :  93 - 0x5d
      13'h11C8: dout <= 8'b01011010; // 4552 :  90 - 0x5a
      13'h11C9: dout <= 8'b01000000; // 4553 :  64 - 0x40
      13'h11CA: dout <= 8'b00000000; // 4554 :   0 - 0x0
      13'h11CB: dout <= 8'b00000000; // 4555 :   0 - 0x0
      13'h11CC: dout <= 8'b00010101; // 4556 :  21 - 0x15
      13'h11CD: dout <= 8'b01010101; // 4557 :  85 - 0x55
      13'h11CE: dout <= 8'b01010101; // 4558 :  85 - 0x55
      13'h11CF: dout <= 8'b01010101; // 4559 :  85 - 0x55
      13'h11D0: dout <= 8'b01010101; // 4560 :  85 - 0x55 -- Background 0x1d
      13'h11D1: dout <= 8'b01000000; // 4561 :  64 - 0x40
      13'h11D2: dout <= 8'b00000000; // 4562 :   0 - 0x0
      13'h11D3: dout <= 8'b00000000; // 4563 :   0 - 0x0
      13'h11D4: dout <= 8'b00010100; // 4564 :  20 - 0x14
      13'h11D5: dout <= 8'b00000011; // 4565 :   3 - 0x3
      13'h11D6: dout <= 8'b00001000; // 4566 :   8 - 0x8
      13'h11D7: dout <= 8'b10101101; // 4567 : 173 - 0xad
      13'h11D8: dout <= 8'b00000000; // 4568 :   0 - 0x0
      13'h11D9: dout <= 8'b10010011; // 4569 : 147 - 0x93
      13'h11DA: dout <= 8'b00000000; // 4570 :   0 - 0x0
      13'h11DB: dout <= 8'b00010101; // 4571 :  21 - 0x15
      13'h11DC: dout <= 8'b01010101; // 4572 :  85 - 0x55
      13'h11DD: dout <= 8'b01010101; // 4573 :  85 - 0x55
      13'h11DE: dout <= 8'b01010101; // 4574 :  85 - 0x55
      13'h11DF: dout <= 8'b01010101; // 4575 :  85 - 0x55
      13'h11E0: dout <= 8'b01010101; // 4576 :  85 - 0x55 -- Background 0x1e
      13'h11E1: dout <= 8'b01010000; // 4577 :  80 - 0x50
      13'h11E2: dout <= 8'b00000000; // 4578 :   0 - 0x0
      13'h11E3: dout <= 8'b00010101; // 4579 :  21 - 0x15
      13'h11E4: dout <= 8'b01110101; // 4580 : 117 - 0x75
      13'h11E5: dout <= 8'b01010101; // 4581 :  85 - 0x55
      13'h11E6: dout <= 8'b01010111; // 4582 :  87 - 0x57
      13'h11E7: dout <= 8'b01010101; // 4583 :  85 - 0x55
      13'h11E8: dout <= 8'b01010111; // 4584 :  87 - 0x57
      13'h11E9: dout <= 8'b01010000; // 4585 :  80 - 0x50
      13'h11EA: dout <= 8'b00000000; // 4586 :   0 - 0x0
      13'h11EB: dout <= 8'b00011101; // 4587 :  29 - 0x1d
      13'h11EC: dout <= 8'b01010101; // 4588 :  85 - 0x55
      13'h11ED: dout <= 8'b01110101; // 4589 : 117 - 0x75
      13'h11EE: dout <= 8'b01010101; // 4590 :  85 - 0x55
      13'h11EF: dout <= 8'b01011101; // 4591 :  93 - 0x5d
      13'h11F0: dout <= 8'b01010101; // 4592 :  85 - 0x55 -- Background 0x1f
      13'h11F1: dout <= 8'b01010000; // 4593 :  80 - 0x50
      13'h11F2: dout <= 8'b00000000; // 4594 :   0 - 0x0
      13'h11F3: dout <= 8'b00010101; // 4595 :  21 - 0x15
      13'h11F4: dout <= 8'b01010111; // 4596 :  87 - 0x57
      13'h11F5: dout <= 8'b01010101; // 4597 :  85 - 0x55
      13'h11F6: dout <= 8'b01010101; // 4598 :  85 - 0x55
      13'h11F7: dout <= 8'b01010101; // 4599 :  85 - 0x55
      13'h11F8: dout <= 8'b01110101; // 4600 : 117 - 0x75
      13'h11F9: dout <= 8'b01010000; // 4601 :  80 - 0x50
      13'h11FA: dout <= 8'b00000000; // 4602 :   0 - 0x0
      13'h11FB: dout <= 8'b00010101; // 4603 :  21 - 0x15
      13'h11FC: dout <= 8'b01010101; // 4604 :  85 - 0x55
      13'h11FD: dout <= 8'b01010101; // 4605 :  85 - 0x55
      13'h11FE: dout <= 8'b00000001; // 4606 :   1 - 0x1
      13'h11FF: dout <= 8'b01010101; // 4607 :  85 - 0x55
      13'h1200: dout <= 8'b01010101; // 4608 :  85 - 0x55 -- Background 0x20
      13'h1201: dout <= 8'b11010000; // 4609 : 208 - 0xd0
      13'h1202: dout <= 8'b00000000; // 4610 :   0 - 0x0
      13'h1203: dout <= 8'b00010111; // 4611 :  23 - 0x17
      13'h1204: dout <= 8'b01010101; // 4612 :  85 - 0x55
      13'h1205: dout <= 8'b01010101; // 4613 :  85 - 0x55
      13'h1206: dout <= 8'b00000001; // 4614 :   1 - 0x1
      13'h1207: dout <= 8'b01010111; // 4615 :  87 - 0x57
      13'h1208: dout <= 8'b01010101; // 4616 :  85 - 0x55
      13'h1209: dout <= 8'b01010000; // 4617 :  80 - 0x50
      13'h120A: dout <= 8'b00000000; // 4618 :   0 - 0x0
      13'h120B: dout <= 8'b00010101; // 4619 :  21 - 0x15
      13'h120C: dout <= 8'b01011101; // 4620 :  93 - 0x5d
      13'h120D: dout <= 8'b01010101; // 4621 :  85 - 0x55
      13'h120E: dout <= 8'b00000001; // 4622 :   1 - 0x1
      13'h120F: dout <= 8'b01010101; // 4623 :  85 - 0x55
      13'h1210: dout <= 8'b01010101; // 4624 :  85 - 0x55 -- Background 0x21
      13'h1211: dout <= 8'b01010000; // 4625 :  80 - 0x50
      13'h1212: dout <= 8'b00000000; // 4626 :   0 - 0x0
      13'h1213: dout <= 8'b00010101; // 4627 :  21 - 0x15
      13'h1214: dout <= 8'b01010101; // 4628 :  85 - 0x55
      13'h1215: dout <= 8'b01110101; // 4629 : 117 - 0x75
      13'h1216: dout <= 8'b01010101; // 4630 :  85 - 0x55
      13'h1217: dout <= 8'b01010101; // 4631 :  85 - 0x55
      13'h1218: dout <= 8'b01110101; // 4632 : 117 - 0x75
      13'h1219: dout <= 8'b01010000; // 4633 :  80 - 0x50
      13'h121A: dout <= 8'b00000000; // 4634 :   0 - 0x0
      13'h121B: dout <= 8'b00011101; // 4635 :  29 - 0x1d
      13'h121C: dout <= 8'b01010101; // 4636 :  85 - 0x55
      13'h121D: dout <= 8'b01010101; // 4637 :  85 - 0x55
      13'h121E: dout <= 8'b01010101; // 4638 :  85 - 0x55
      13'h121F: dout <= 8'b01110101; // 4639 : 117 - 0x75
      13'h1220: dout <= 8'b01010101; // 4640 :  85 - 0x55 -- Background 0x22
      13'h1221: dout <= 8'b01010000; // 4641 :  80 - 0x50
      13'h1222: dout <= 8'b00000000; // 4642 :   0 - 0x0
      13'h1223: dout <= 8'b00010101; // 4643 :  21 - 0x15
      13'h1224: dout <= 8'b01110101; // 4644 : 117 - 0x75
      13'h1225: dout <= 8'b01010101; // 4645 :  85 - 0x55
      13'h1226: dout <= 8'b11010101; // 4646 : 213 - 0xd5
      13'h1227: dout <= 8'b01010101; // 4647 :  85 - 0x55
      13'h1228: dout <= 8'b01010111; // 4648 :  87 - 0x57
      13'h1229: dout <= 8'b01010000; // 4649 :  80 - 0x50
      13'h122A: dout <= 8'b00000000; // 4650 :   0 - 0x0
      13'h122B: dout <= 8'b00010101; // 4651 :  21 - 0x15
      13'h122C: dout <= 8'b01010101; // 4652 :  85 - 0x55
      13'h122D: dout <= 8'b01010101; // 4653 :  85 - 0x55
      13'h122E: dout <= 8'b01010101; // 4654 :  85 - 0x55
      13'h122F: dout <= 8'b01010101; // 4655 :  85 - 0x55
      13'h1230: dout <= 8'b01010101; // 4656 :  85 - 0x55 -- Background 0x23
      13'h1231: dout <= 8'b01010000; // 4657 :  80 - 0x50
      13'h1232: dout <= 8'b00000000; // 4658 :   0 - 0x0
      13'h1233: dout <= 8'b00011001; // 4659 :  25 - 0x19
      13'h1234: dout <= 8'b00001101; // 4660 :  13 - 0xd
      13'h1235: dout <= 8'b00001000; // 4661 :   8 - 0x8
      13'h1236: dout <= 8'b11110111; // 4662 : 247 - 0xf7
      13'h1237: dout <= 8'b00000000; // 4663 :   0 - 0x0
      13'h1238: dout <= 8'b01100111; // 4664 : 103 - 0x67
      13'h1239: dout <= 8'b00000000; // 4665 :   0 - 0x0
      13'h123A: dout <= 8'b00010101; // 4666 :  21 - 0x15
      13'h123B: dout <= 8'b01010101; // 4667 :  85 - 0x55
      13'h123C: dout <= 8'b01010101; // 4668 :  85 - 0x55
      13'h123D: dout <= 8'b01010101; // 4669 :  85 - 0x55
      13'h123E: dout <= 8'b01010101; // 4670 :  85 - 0x55
      13'h123F: dout <= 8'b01010101; // 4671 :  85 - 0x55
      13'h1240: dout <= 8'b01010000; // 4672 :  80 - 0x50 -- Background 0x24
      13'h1241: dout <= 8'b00000000; // 4673 :   0 - 0x0
      13'h1242: dout <= 8'b00011010; // 4674 :  26 - 0x1a
      13'h1243: dout <= 8'b10101001; // 4675 : 169 - 0xa9
      13'h1244: dout <= 8'b10101010; // 4676 : 170 - 0xaa
      13'h1245: dout <= 8'b10011001; // 4677 : 153 - 0x99
      13'h1246: dout <= 8'b01011001; // 4678 :  89 - 0x59
      13'h1247: dout <= 8'b10101010; // 4679 : 170 - 0xaa
      13'h1248: dout <= 8'b10010000; // 4680 : 144 - 0x90
      13'h1249: dout <= 8'b00000000; // 4681 :   0 - 0x0
      13'h124A: dout <= 8'b00011001; // 4682 :  25 - 0x19
      13'h124B: dout <= 8'b01011001; // 4683 :  89 - 0x59
      13'h124C: dout <= 8'b10010101; // 4684 : 149 - 0x95
      13'h124D: dout <= 8'b10011001; // 4685 : 153 - 0x99
      13'h124E: dout <= 8'b01011001; // 4686 :  89 - 0x59
      13'h124F: dout <= 8'b10010101; // 4687 : 149 - 0x95
      13'h1250: dout <= 8'b10010000; // 4688 : 144 - 0x90 -- Background 0x25
      13'h1251: dout <= 8'b00000000; // 4689 :   0 - 0x0
      13'h1252: dout <= 8'b00010101; // 4690 :  21 - 0x15
      13'h1253: dout <= 8'b01011001; // 4691 :  89 - 0x59
      13'h1254: dout <= 8'b10010101; // 4692 : 149 - 0x95
      13'h1255: dout <= 8'b10011001; // 4693 : 153 - 0x99
      13'h1256: dout <= 8'b01011001; // 4694 :  89 - 0x59
      13'h1257: dout <= 8'b10010101; // 4695 : 149 - 0x95
      13'h1258: dout <= 8'b01010000; // 4696 :  80 - 0x50
      13'h1259: dout <= 8'b00000000; // 4697 :   0 - 0x0
      13'h125A: dout <= 8'b00010000; // 4698 :  16 - 0x10
      13'h125B: dout <= 8'b00010101; // 4699 :  21 - 0x15
      13'h125C: dout <= 8'b10010101; // 4700 : 149 - 0x95
      13'h125D: dout <= 8'b10011010; // 4701 : 154 - 0x9a
      13'h125E: dout <= 8'b10101001; // 4702 : 169 - 0xa9
      13'h125F: dout <= 8'b01010101; // 4703 :  85 - 0x55
      13'h1260: dout <= 8'b01010000; // 4704 :  80 - 0x50 -- Background 0x26
      13'h1261: dout <= 8'b00000000; // 4705 :   0 - 0x0
      13'h1262: dout <= 8'b00010000; // 4706 :  16 - 0x10
      13'h1263: dout <= 8'b00010101; // 4707 :  21 - 0x15
      13'h1264: dout <= 8'b01010101; // 4708 :  85 - 0x55
      13'h1265: dout <= 8'b01010101; // 4709 :  85 - 0x55
      13'h1266: dout <= 8'b01010101; // 4710 :  85 - 0x55
      13'h1267: dout <= 8'b01010101; // 4711 :  85 - 0x55
      13'h1268: dout <= 8'b01010000; // 4712 :  80 - 0x50
      13'h1269: dout <= 8'b00000000; // 4713 :   0 - 0x0
      13'h126A: dout <= 8'b00010000; // 4714 :  16 - 0x10
      13'h126B: dout <= 8'b00010101; // 4715 :  21 - 0x15
      13'h126C: dout <= 8'b10101010; // 4716 : 170 - 0xaa
      13'h126D: dout <= 8'b10011001; // 4717 : 153 - 0x99
      13'h126E: dout <= 8'b01011001; // 4718 :  89 - 0x59
      13'h126F: dout <= 8'b01010101; // 4719 :  85 - 0x55
      13'h1270: dout <= 8'b01010000; // 4720 :  80 - 0x50 -- Background 0x27
      13'h1271: dout <= 8'b00000000; // 4721 :   0 - 0x0
      13'h1272: dout <= 8'b00010101; // 4722 :  21 - 0x15
      13'h1273: dout <= 8'b01011001; // 4723 :  89 - 0x59
      13'h1274: dout <= 8'b10010101; // 4724 : 149 - 0x95
      13'h1275: dout <= 8'b10011001; // 4725 : 153 - 0x99
      13'h1276: dout <= 8'b01011001; // 4726 :  89 - 0x59
      13'h1277: dout <= 8'b10010101; // 4727 : 149 - 0x95
      13'h1278: dout <= 8'b01010000; // 4728 :  80 - 0x50
      13'h1279: dout <= 8'b00000000; // 4729 :   0 - 0x0
      13'h127A: dout <= 8'b00011001; // 4730 :  25 - 0x19
      13'h127B: dout <= 8'b01011001; // 4731 :  89 - 0x59
      13'h127C: dout <= 8'b10010101; // 4732 : 149 - 0x95
      13'h127D: dout <= 8'b10011001; // 4733 : 153 - 0x99
      13'h127E: dout <= 8'b01011001; // 4734 :  89 - 0x59
      13'h127F: dout <= 8'b10010101; // 4735 : 149 - 0x95
      13'h1280: dout <= 8'b10010000; // 4736 : 144 - 0x90 -- Background 0x28
      13'h1281: dout <= 8'b00000000; // 4737 :   0 - 0x0
      13'h1282: dout <= 8'b00011010; // 4738 :  26 - 0x1a
      13'h1283: dout <= 8'b10101001; // 4739 : 169 - 0xa9
      13'h1284: dout <= 8'b10010101; // 4740 : 149 - 0x95
      13'h1285: dout <= 8'b10011010; // 4741 : 154 - 0x9a
      13'h1286: dout <= 8'b10101001; // 4742 : 169 - 0xa9
      13'h1287: dout <= 8'b10101010; // 4743 : 170 - 0xaa
      13'h1288: dout <= 8'b10010000; // 4744 : 144 - 0x90
      13'h1289: dout <= 8'b00000000; // 4745 :   0 - 0x0
      13'h128A: dout <= 8'b00010101; // 4746 :  21 - 0x15
      13'h128B: dout <= 8'b01010101; // 4747 :  85 - 0x55
      13'h128C: dout <= 8'b01010101; // 4748 :  85 - 0x55
      13'h128D: dout <= 8'b01010101; // 4749 :  85 - 0x55
      13'h128E: dout <= 8'b01010101; // 4750 :  85 - 0x55
      13'h128F: dout <= 8'b01010101; // 4751 :  85 - 0x55
      13'h1290: dout <= 8'b01010000; // 4752 :  80 - 0x50 -- Background 0x29
      13'h1291: dout <= 8'b00000000; // 4753 :   0 - 0x0
      13'h1292: dout <= 8'b00011001; // 4754 :  25 - 0x19
      13'h1293: dout <= 8'b00000011; // 4755 :   3 - 0x3
      13'h1294: dout <= 8'b00001000; // 4756 :   8 - 0x8
      13'h1295: dout <= 8'b10111110; // 4757 : 190 - 0xbe
      13'h1296: dout <= 8'b00000000; // 4758 :   0 - 0x0
      13'h1297: dout <= 8'b10000110; // 4759 : 134 - 0x86
      13'h1298: dout <= 8'b00000000; // 4760 :   0 - 0x0
      13'h1299: dout <= 8'b00010101; // 4761 :  21 - 0x15
      13'h129A: dout <= 8'b01010111; // 4762 :  87 - 0x57
      13'h129B: dout <= 8'b01010101; // 4763 :  85 - 0x55
      13'h129C: dout <= 8'b01010101; // 4764 :  85 - 0x55
      13'h129D: dout <= 8'b01010111; // 4765 :  87 - 0x57
      13'h129E: dout <= 8'b01010101; // 4766 :  85 - 0x55
      13'h129F: dout <= 8'b01010000; // 4767 :  80 - 0x50
      13'h12A0: dout <= 8'b00000000; // 4768 :   0 - 0x0 -- Background 0x2a
      13'h12A1: dout <= 8'b00010101; // 4769 :  21 - 0x15
      13'h12A2: dout <= 8'b01010111; // 4770 :  87 - 0x57
      13'h12A3: dout <= 8'b01101010; // 4771 : 106 - 0x6a
      13'h12A4: dout <= 8'b01010110; // 4772 :  86 - 0x56
      13'h12A5: dout <= 8'b10100111; // 4773 : 167 - 0xa7
      13'h12A6: dout <= 8'b01010101; // 4774 :  85 - 0x55
      13'h12A7: dout <= 8'b01010000; // 4775 :  80 - 0x50
      13'h12A8: dout <= 8'b00000000; // 4776 :   0 - 0x0
      13'h12A9: dout <= 8'b00010101; // 4777 :  21 - 0x15
      13'h12AA: dout <= 8'b01010111; // 4778 :  87 - 0x57
      13'h12AB: dout <= 8'b01101010; // 4779 : 106 - 0x6a
      13'h12AC: dout <= 8'b01010110; // 4780 :  86 - 0x56
      13'h12AD: dout <= 8'b10100111; // 4781 : 167 - 0xa7
      13'h12AE: dout <= 8'b01010101; // 4782 :  85 - 0x55
      13'h12AF: dout <= 8'b01010000; // 4783 :  80 - 0x50
      13'h12B0: dout <= 8'b00000000; // 4784 :   0 - 0x0 -- Background 0x2b
      13'h12B1: dout <= 8'b00010101; // 4785 :  21 - 0x15
      13'h12B2: dout <= 8'b01010111; // 4786 :  87 - 0x57
      13'h12B3: dout <= 8'b01010101; // 4787 :  85 - 0x55
      13'h12B4: dout <= 8'b01110101; // 4788 : 117 - 0x75
      13'h12B5: dout <= 8'b01010111; // 4789 :  87 - 0x57
      13'h12B6: dout <= 8'b01010101; // 4790 :  85 - 0x55
      13'h12B7: dout <= 8'b01010000; // 4791 :  80 - 0x50
      13'h12B8: dout <= 8'b00000000; // 4792 :   0 - 0x0
      13'h12B9: dout <= 8'b00010000; // 4793 :  16 - 0x10
      13'h12BA: dout <= 8'b00010101; // 4794 :  21 - 0x15
      13'h12BB: dout <= 8'b01010101; // 4795 :  85 - 0x55
      13'h12BC: dout <= 8'b01110101; // 4796 : 117 - 0x75
      13'h12BD: dout <= 8'b01010101; // 4797 :  85 - 0x55
      13'h12BE: dout <= 8'b01010101; // 4798 :  85 - 0x55
      13'h12BF: dout <= 8'b01010000; // 4799 :  80 - 0x50
      13'h12C0: dout <= 8'b00000000; // 4800 :   0 - 0x0 -- Background 0x2c
      13'h12C1: dout <= 8'b00010000; // 4801 :  16 - 0x10
      13'h12C2: dout <= 8'b00010101; // 4802 :  21 - 0x15
      13'h12C3: dout <= 8'b01010101; // 4803 :  85 - 0x55
      13'h12C4: dout <= 8'b01110101; // 4804 : 117 - 0x75
      13'h12C5: dout <= 8'b01010101; // 4805 :  85 - 0x55
      13'h12C6: dout <= 8'b01010101; // 4806 :  85 - 0x55
      13'h12C7: dout <= 8'b01010000; // 4807 :  80 - 0x50
      13'h12C8: dout <= 8'b00000000; // 4808 :   0 - 0x0
      13'h12C9: dout <= 8'b00010000; // 4809 :  16 - 0x10
      13'h12CA: dout <= 8'b00010101; // 4810 :  21 - 0x15
      13'h12CB: dout <= 8'b01010101; // 4811 :  85 - 0x55
      13'h12CC: dout <= 8'b01110101; // 4812 : 117 - 0x75
      13'h12CD: dout <= 8'b01010101; // 4813 :  85 - 0x55
      13'h12CE: dout <= 8'b01010101; // 4814 :  85 - 0x55
      13'h12CF: dout <= 8'b01010000; // 4815 :  80 - 0x50
      13'h12D0: dout <= 8'b00000000; // 4816 :   0 - 0x0 -- Background 0x2d
      13'h12D1: dout <= 8'b00010101; // 4817 :  21 - 0x15
      13'h12D2: dout <= 8'b01010111; // 4818 :  87 - 0x57
      13'h12D3: dout <= 8'b01010101; // 4819 :  85 - 0x55
      13'h12D4: dout <= 8'b01110101; // 4820 : 117 - 0x75
      13'h12D5: dout <= 8'b01010111; // 4821 :  87 - 0x57
      13'h12D6: dout <= 8'b01010101; // 4822 :  85 - 0x55
      13'h12D7: dout <= 8'b01010000; // 4823 :  80 - 0x50
      13'h12D8: dout <= 8'b00000000; // 4824 :   0 - 0x0
      13'h12D9: dout <= 8'b00010101; // 4825 :  21 - 0x15
      13'h12DA: dout <= 8'b01010111; // 4826 :  87 - 0x57
      13'h12DB: dout <= 8'b01101010; // 4827 : 106 - 0x6a
      13'h12DC: dout <= 8'b01010110; // 4828 :  86 - 0x56
      13'h12DD: dout <= 8'b10100111; // 4829 : 167 - 0xa7
      13'h12DE: dout <= 8'b01010101; // 4830 :  85 - 0x55
      13'h12DF: dout <= 8'b01010000; // 4831 :  80 - 0x50
      13'h12E0: dout <= 8'b00000000; // 4832 :   0 - 0x0 -- Background 0x2e
      13'h12E1: dout <= 8'b00010101; // 4833 :  21 - 0x15
      13'h12E2: dout <= 8'b01010111; // 4834 :  87 - 0x57
      13'h12E3: dout <= 8'b01101010; // 4835 : 106 - 0x6a
      13'h12E4: dout <= 8'b01010110; // 4836 :  86 - 0x56
      13'h12E5: dout <= 8'b10100111; // 4837 : 167 - 0xa7
      13'h12E6: dout <= 8'b01010101; // 4838 :  85 - 0x55
      13'h12E7: dout <= 8'b01010000; // 4839 :  80 - 0x50
      13'h12E8: dout <= 8'b00000000; // 4840 :   0 - 0x0
      13'h12E9: dout <= 8'b00010101; // 4841 :  21 - 0x15
      13'h12EA: dout <= 8'b01010111; // 4842 :  87 - 0x57
      13'h12EB: dout <= 8'b01010101; // 4843 :  85 - 0x55
      13'h12EC: dout <= 8'b01010101; // 4844 :  85 - 0x55
      13'h12ED: dout <= 8'b01010111; // 4845 :  87 - 0x57
      13'h12EE: dout <= 8'b01010101; // 4846 :  85 - 0x55
      13'h12EF: dout <= 8'b01010000; // 4847 :  80 - 0x50
      13'h12F0: dout <= 8'b00000000; // 4848 :   0 - 0x0 -- Background 0x2f
      13'h12F1: dout <= 8'b00011001; // 4849 :  25 - 0x19
      13'h12F2: dout <= 8'b00000011; // 4850 :   3 - 0x3
      13'h12F3: dout <= 8'b00001000; // 4851 :   8 - 0x8
      13'h12F4: dout <= 8'b11011101; // 4852 : 221 - 0xdd
      13'h12F5: dout <= 8'b00000000; // 4853 :   0 - 0x0
      13'h12F6: dout <= 8'b01110011; // 4854 : 115 - 0x73
      13'h12F7: dout <= 8'b00000000; // 4855 :   0 - 0x0
      13'h12F8: dout <= 8'b00010101; // 4856 :  21 - 0x15
      13'h12F9: dout <= 8'b01010101; // 4857 :  85 - 0x55
      13'h12FA: dout <= 8'b01010101; // 4858 :  85 - 0x55
      13'h12FB: dout <= 8'b01010101; // 4859 :  85 - 0x55
      13'h12FC: dout <= 8'b01010101; // 4860 :  85 - 0x55
      13'h12FD: dout <= 8'b01010101; // 4861 :  85 - 0x55
      13'h12FE: dout <= 8'b01010101; // 4862 :  85 - 0x55
      13'h12FF: dout <= 8'b01010100; // 4863 :  84 - 0x54
      13'h1300: dout <= 8'b00011001; // 4864 :  25 - 0x19 -- Background 0x30
      13'h1301: dout <= 8'b01100101; // 4865 : 101 - 0x65
      13'h1302: dout <= 8'b10010110; // 4866 : 150 - 0x96
      13'h1303: dout <= 8'b10100101; // 4867 : 165 - 0xa5
      13'h1304: dout <= 8'b01011010; // 4868 :  90 - 0x5a
      13'h1305: dout <= 8'b10010110; // 4869 : 150 - 0x96
      13'h1306: dout <= 8'b01011001; // 4870 :  89 - 0x59
      13'h1307: dout <= 8'b01100100; // 4871 : 100 - 0x64
      13'h1308: dout <= 8'b00011001; // 4872 :  25 - 0x19
      13'h1309: dout <= 8'b01100101; // 4873 : 101 - 0x65
      13'h130A: dout <= 8'b10010101; // 4874 : 149 - 0x95
      13'h130B: dout <= 8'b01010101; // 4875 :  85 - 0x55
      13'h130C: dout <= 8'b01010101; // 4876 :  85 - 0x55
      13'h130D: dout <= 8'b01010110; // 4877 :  86 - 0x56
      13'h130E: dout <= 8'b01011001; // 4878 :  89 - 0x59
      13'h130F: dout <= 8'b01100100; // 4879 : 100 - 0x64
      13'h1310: dout <= 8'b00011001; // 4880 :  25 - 0x19 -- Background 0x31
      13'h1311: dout <= 8'b01100101; // 4881 : 101 - 0x65
      13'h1312: dout <= 8'b10010110; // 4882 : 150 - 0x96
      13'h1313: dout <= 8'b10100101; // 4883 : 165 - 0xa5
      13'h1314: dout <= 8'b01011010; // 4884 :  90 - 0x5a
      13'h1315: dout <= 8'b10010110; // 4885 : 150 - 0x96
      13'h1316: dout <= 8'b01011001; // 4886 :  89 - 0x59
      13'h1317: dout <= 8'b01100100; // 4887 : 100 - 0x64
      13'h1318: dout <= 8'b00010101; // 4888 :  21 - 0x15
      13'h1319: dout <= 8'b01010101; // 4889 :  85 - 0x55
      13'h131A: dout <= 8'b01010101; // 4890 :  85 - 0x55
      13'h131B: dout <= 8'b01010000; // 4891 :  80 - 0x50
      13'h131C: dout <= 8'b00000101; // 4892 :   5 - 0x5
      13'h131D: dout <= 8'b01010101; // 4893 :  85 - 0x55
      13'h131E: dout <= 8'b01010101; // 4894 :  85 - 0x55
      13'h131F: dout <= 8'b01010100; // 4895 :  84 - 0x54
      13'h1320: dout <= 8'b00011111; // 4896 :  31 - 0x1f -- Background 0x32
      13'h1321: dout <= 8'b01111101; // 4897 : 125 - 0x7d
      13'h1322: dout <= 8'b11010101; // 4898 : 213 - 0xd5
      13'h1323: dout <= 8'b01010000; // 4899 :  80 - 0x50
      13'h1324: dout <= 8'b00000101; // 4900 :   5 - 0x5
      13'h1325: dout <= 8'b01010111; // 4901 :  87 - 0x57
      13'h1326: dout <= 8'b11111111; // 4902 : 255 - 0xff
      13'h1327: dout <= 8'b01110100; // 4903 : 116 - 0x74
      13'h1328: dout <= 8'b00010101; // 4904 :  21 - 0x15
      13'h1329: dout <= 8'b01010101; // 4905 :  85 - 0x55
      13'h132A: dout <= 8'b01010101; // 4906 :  85 - 0x55
      13'h132B: dout <= 8'b01010000; // 4907 :  80 - 0x50
      13'h132C: dout <= 8'b00000101; // 4908 :   5 - 0x5
      13'h132D: dout <= 8'b01010101; // 4909 :  85 - 0x55
      13'h132E: dout <= 8'b01010101; // 4910 :  85 - 0x55
      13'h132F: dout <= 8'b01010100; // 4911 :  84 - 0x54
      13'h1330: dout <= 8'b00011001; // 4912 :  25 - 0x19 -- Background 0x33
      13'h1331: dout <= 8'b01100101; // 4913 : 101 - 0x65
      13'h1332: dout <= 8'b10010110; // 4914 : 150 - 0x96
      13'h1333: dout <= 8'b10100101; // 4915 : 165 - 0xa5
      13'h1334: dout <= 8'b01011010; // 4916 :  90 - 0x5a
      13'h1335: dout <= 8'b10010110; // 4917 : 150 - 0x96
      13'h1336: dout <= 8'b01011001; // 4918 :  89 - 0x59
      13'h1337: dout <= 8'b01100100; // 4919 : 100 - 0x64
      13'h1338: dout <= 8'b00011001; // 4920 :  25 - 0x19
      13'h1339: dout <= 8'b01100101; // 4921 : 101 - 0x65
      13'h133A: dout <= 8'b10010101; // 4922 : 149 - 0x95
      13'h133B: dout <= 8'b01010101; // 4923 :  85 - 0x55
      13'h133C: dout <= 8'b01010101; // 4924 :  85 - 0x55
      13'h133D: dout <= 8'b01010110; // 4925 :  86 - 0x56
      13'h133E: dout <= 8'b01011001; // 4926 :  89 - 0x59
      13'h133F: dout <= 8'b01100100; // 4927 : 100 - 0x64
      13'h1340: dout <= 8'b00011001; // 4928 :  25 - 0x19 -- Background 0x34
      13'h1341: dout <= 8'b01100101; // 4929 : 101 - 0x65
      13'h1342: dout <= 8'b10010110; // 4930 : 150 - 0x96
      13'h1343: dout <= 8'b10100101; // 4931 : 165 - 0xa5
      13'h1344: dout <= 8'b01011010; // 4932 :  90 - 0x5a
      13'h1345: dout <= 8'b10010110; // 4933 : 150 - 0x96
      13'h1346: dout <= 8'b01011001; // 4934 :  89 - 0x59
      13'h1347: dout <= 8'b01100100; // 4935 : 100 - 0x64
      13'h1348: dout <= 8'b00010101; // 4936 :  21 - 0x15
      13'h1349: dout <= 8'b01010101; // 4937 :  85 - 0x55
      13'h134A: dout <= 8'b01010101; // 4938 :  85 - 0x55
      13'h134B: dout <= 8'b01010101; // 4939 :  85 - 0x55
      13'h134C: dout <= 8'b01010101; // 4940 :  85 - 0x55
      13'h134D: dout <= 8'b01010101; // 4941 :  85 - 0x55
      13'h134E: dout <= 8'b01010101; // 4942 :  85 - 0x55
      13'h134F: dout <= 8'b01010100; // 4943 :  84 - 0x54
      13'h1350: dout <= 8'b00011110; // 4944 :  30 - 0x1e -- Background 0x35
      13'h1351: dout <= 8'b00001111; // 4945 :  15 - 0xf
      13'h1352: dout <= 8'b00001000; // 4946 :   8 - 0x8
      13'h1353: dout <= 8'b11110111; // 4947 : 247 - 0xf7
      13'h1354: dout <= 8'b00000000; // 4948 :   0 - 0x0
      13'h1355: dout <= 8'b01100111; // 4949 : 103 - 0x67
      13'h1356: dout <= 8'b00000000; // 4950 :   0 - 0x0
      13'h1357: dout <= 8'b00010101; // 4951 :  21 - 0x15
      13'h1358: dout <= 8'b01010101; // 4952 :  85 - 0x55
      13'h1359: dout <= 8'b01010101; // 4953 :  85 - 0x55
      13'h135A: dout <= 8'b01010101; // 4954 :  85 - 0x55
      13'h135B: dout <= 8'b01010101; // 4955 :  85 - 0x55
      13'h135C: dout <= 8'b01010101; // 4956 :  85 - 0x55
      13'h135D: dout <= 8'b01010101; // 4957 :  85 - 0x55
      13'h135E: dout <= 8'b01010100; // 4958 :  84 - 0x54
      13'h135F: dout <= 8'b00010111; // 4959 :  23 - 0x17
      13'h1360: dout <= 8'b01110101; // 4960 : 117 - 0x75 -- Background 0x36
      13'h1361: dout <= 8'b01010110; // 4961 :  86 - 0x56
      13'h1362: dout <= 8'b10100101; // 4962 : 165 - 0xa5
      13'h1363: dout <= 8'b01011010; // 4963 :  90 - 0x5a
      13'h1364: dout <= 8'b10010101; // 4964 : 149 - 0x95
      13'h1365: dout <= 8'b01011101; // 4965 :  93 - 0x5d
      13'h1366: dout <= 8'b11010100; // 4966 : 212 - 0xd4
      13'h1367: dout <= 8'b00010101; // 4967 :  21 - 0x15
      13'h1368: dout <= 8'b01010101; // 4968 :  85 - 0x55
      13'h1369: dout <= 8'b01110110; // 4969 : 118 - 0x76
      13'h136A: dout <= 8'b10100101; // 4970 : 165 - 0xa5
      13'h136B: dout <= 8'b01011010; // 4971 :  90 - 0x5a
      13'h136C: dout <= 8'b10011101; // 4972 : 157 - 0x9d
      13'h136D: dout <= 8'b01010101; // 4973 :  85 - 0x55
      13'h136E: dout <= 8'b01010100; // 4974 :  84 - 0x54
      13'h136F: dout <= 8'b00010111; // 4975 :  23 - 0x17
      13'h1370: dout <= 8'b01010101; // 4976 :  85 - 0x55 -- Background 0x37
      13'h1371: dout <= 8'b01110101; // 4977 : 117 - 0x75
      13'h1372: dout <= 8'b01010101; // 4978 :  85 - 0x55
      13'h1373: dout <= 8'b01010101; // 4979 :  85 - 0x55
      13'h1374: dout <= 8'b01011101; // 4980 :  93 - 0x5d
      13'h1375: dout <= 8'b01010101; // 4981 :  85 - 0x55
      13'h1376: dout <= 8'b11010100; // 4982 : 212 - 0xd4
      13'h1377: dout <= 8'b00010101; // 4983 :  21 - 0x15
      13'h1378: dout <= 8'b01101010; // 4984 : 106 - 0x6a
      13'h1379: dout <= 8'b01110101; // 4985 : 117 - 0x75
      13'h137A: dout <= 8'b01010000; // 4986 :  80 - 0x50
      13'h137B: dout <= 8'b00000101; // 4987 :   5 - 0x5
      13'h137C: dout <= 8'b01011101; // 4988 :  93 - 0x5d
      13'h137D: dout <= 8'b10101001; // 4989 : 169 - 0xa9
      13'h137E: dout <= 8'b01010100; // 4990 :  84 - 0x54
      13'h137F: dout <= 8'b00010101; // 4991 :  21 - 0x15
      13'h1380: dout <= 8'b01101110; // 4992 : 110 - 0x6e -- Background 0x38
      13'h1381: dout <= 8'b01110101; // 4993 : 117 - 0x75
      13'h1382: dout <= 8'b01010000; // 4994 :  80 - 0x50
      13'h1383: dout <= 8'b00000101; // 4995 :   5 - 0x5
      13'h1384: dout <= 8'b01011101; // 4996 :  93 - 0x5d
      13'h1385: dout <= 8'b10111001; // 4997 : 185 - 0xb9
      13'h1386: dout <= 8'b01010100; // 4998 :  84 - 0x54
      13'h1387: dout <= 8'b00010101; // 4999 :  21 - 0x15
      13'h1388: dout <= 8'b01101010; // 5000 : 106 - 0x6a
      13'h1389: dout <= 8'b01110101; // 5001 : 117 - 0x75
      13'h138A: dout <= 8'b01010000; // 5002 :  80 - 0x50
      13'h138B: dout <= 8'b00000101; // 5003 :   5 - 0x5
      13'h138C: dout <= 8'b01011101; // 5004 :  93 - 0x5d
      13'h138D: dout <= 8'b10101001; // 5005 : 169 - 0xa9
      13'h138E: dout <= 8'b01010100; // 5006 :  84 - 0x54
      13'h138F: dout <= 8'b00010111; // 5007 :  23 - 0x17
      13'h1390: dout <= 8'b01010101; // 5008 :  85 - 0x55 -- Background 0x39
      13'h1391: dout <= 8'b01110101; // 5009 : 117 - 0x75
      13'h1392: dout <= 8'b01010101; // 5010 :  85 - 0x55
      13'h1393: dout <= 8'b01010101; // 5011 :  85 - 0x55
      13'h1394: dout <= 8'b01011101; // 5012 :  93 - 0x5d
      13'h1395: dout <= 8'b01010101; // 5013 :  85 - 0x55
      13'h1396: dout <= 8'b11010100; // 5014 : 212 - 0xd4
      13'h1397: dout <= 8'b00010101; // 5015 :  21 - 0x15
      13'h1398: dout <= 8'b01010101; // 5016 :  85 - 0x55
      13'h1399: dout <= 8'b01110101; // 5017 : 117 - 0x75
      13'h139A: dout <= 8'b10101010; // 5018 : 170 - 0xaa
      13'h139B: dout <= 8'b10101010; // 5019 : 170 - 0xaa
      13'h139C: dout <= 8'b01011101; // 5020 :  93 - 0x5d
      13'h139D: dout <= 8'b01010101; // 5021 :  85 - 0x55
      13'h139E: dout <= 8'b01010100; // 5022 :  84 - 0x54
      13'h139F: dout <= 8'b00010111; // 5023 :  23 - 0x17
      13'h13A0: dout <= 8'b01110101; // 5024 : 117 - 0x75 -- Background 0x3a
      13'h13A1: dout <= 8'b01010101; // 5025 :  85 - 0x55
      13'h13A2: dout <= 8'b01101010; // 5026 : 106 - 0x6a
      13'h13A3: dout <= 8'b10101001; // 5027 : 169 - 0xa9
      13'h13A4: dout <= 8'b01010101; // 5028 :  85 - 0x55
      13'h13A5: dout <= 8'b01011101; // 5029 :  93 - 0x5d
      13'h13A6: dout <= 8'b11010100; // 5030 : 212 - 0xd4
      13'h13A7: dout <= 8'b00010101; // 5031 :  21 - 0x15
      13'h13A8: dout <= 8'b01010101; // 5032 :  85 - 0x55
      13'h13A9: dout <= 8'b01010101; // 5033 :  85 - 0x55
      13'h13AA: dout <= 8'b01010101; // 5034 :  85 - 0x55
      13'h13AB: dout <= 8'b01010101; // 5035 :  85 - 0x55
      13'h13AC: dout <= 8'b01010101; // 5036 :  85 - 0x55
      13'h13AD: dout <= 8'b01010101; // 5037 :  85 - 0x55
      13'h13AE: dout <= 8'b01010100; // 5038 :  84 - 0x54
      13'h13AF: dout <= 8'b00011110; // 5039 :  30 - 0x1e
      13'h13B0: dout <= 8'b00001111; // 5040 :  15 - 0xf -- Background 0x3b
      13'h13B1: dout <= 8'b00001000; // 5041 :   8 - 0x8
      13'h13B2: dout <= 8'b11111000; // 5042 : 248 - 0xf8
      13'h13B3: dout <= 8'b00000000; // 5043 :   0 - 0x0
      13'h13B4: dout <= 8'b01100111; // 5044 : 103 - 0x67
      13'h13B5: dout <= 8'b00000000; // 5045 :   0 - 0x0
      13'h13B6: dout <= 8'b00000000; // 5046 :   0 - 0x0
      13'h13B7: dout <= 8'b00000000; // 5047 :   0 - 0x0
      13'h13B8: dout <= 8'b00000000; // 5048 :   0 - 0x0
      13'h13B9: dout <= 8'b00000000; // 5049 :   0 - 0x0
      13'h13BA: dout <= 8'b00000000; // 5050 :   0 - 0x0
      13'h13BB: dout <= 8'b00000000; // 5051 :   0 - 0x0
      13'h13BC: dout <= 8'b00000000; // 5052 :   0 - 0x0
      13'h13BD: dout <= 8'b00000000; // 5053 :   0 - 0x0
      13'h13BE: dout <= 8'b00000000; // 5054 :   0 - 0x0
      13'h13BF: dout <= 8'b00000000; // 5055 :   0 - 0x0
      13'h13C0: dout <= 8'b00000000; // 5056 :   0 - 0x0 -- Background 0x3c
      13'h13C1: dout <= 8'b00000000; // 5057 :   0 - 0x0
      13'h13C2: dout <= 8'b00000000; // 5058 :   0 - 0x0
      13'h13C3: dout <= 8'b00000000; // 5059 :   0 - 0x0
      13'h13C4: dout <= 8'b00000000; // 5060 :   0 - 0x0
      13'h13C5: dout <= 8'b00000000; // 5061 :   0 - 0x0
      13'h13C6: dout <= 8'b00000000; // 5062 :   0 - 0x0
      13'h13C7: dout <= 8'b00000000; // 5063 :   0 - 0x0
      13'h13C8: dout <= 8'b00000000; // 5064 :   0 - 0x0
      13'h13C9: dout <= 8'b00000000; // 5065 :   0 - 0x0
      13'h13CA: dout <= 8'b00000000; // 5066 :   0 - 0x0
      13'h13CB: dout <= 8'b00000000; // 5067 :   0 - 0x0
      13'h13CC: dout <= 8'b00000000; // 5068 :   0 - 0x0
      13'h13CD: dout <= 8'b00000000; // 5069 :   0 - 0x0
      13'h13CE: dout <= 8'b00000000; // 5070 :   0 - 0x0
      13'h13CF: dout <= 8'b00000000; // 5071 :   0 - 0x0
      13'h13D0: dout <= 8'b00000000; // 5072 :   0 - 0x0 -- Background 0x3d
      13'h13D1: dout <= 8'b00000000; // 5073 :   0 - 0x0
      13'h13D2: dout <= 8'b00000000; // 5074 :   0 - 0x0
      13'h13D3: dout <= 8'b00000000; // 5075 :   0 - 0x0
      13'h13D4: dout <= 8'b00000000; // 5076 :   0 - 0x0
      13'h13D5: dout <= 8'b00000000; // 5077 :   0 - 0x0
      13'h13D6: dout <= 8'b00000000; // 5078 :   0 - 0x0
      13'h13D7: dout <= 8'b00000000; // 5079 :   0 - 0x0
      13'h13D8: dout <= 8'b00000000; // 5080 :   0 - 0x0
      13'h13D9: dout <= 8'b00000000; // 5081 :   0 - 0x0
      13'h13DA: dout <= 8'b00000000; // 5082 :   0 - 0x0
      13'h13DB: dout <= 8'b00000000; // 5083 :   0 - 0x0
      13'h13DC: dout <= 8'b00000000; // 5084 :   0 - 0x0
      13'h13DD: dout <= 8'b00000000; // 5085 :   0 - 0x0
      13'h13DE: dout <= 8'b00000000; // 5086 :   0 - 0x0
      13'h13DF: dout <= 8'b00000000; // 5087 :   0 - 0x0
      13'h13E0: dout <= 8'b00000000; // 5088 :   0 - 0x0 -- Background 0x3e
      13'h13E1: dout <= 8'b00000000; // 5089 :   0 - 0x0
      13'h13E2: dout <= 8'b00000000; // 5090 :   0 - 0x0
      13'h13E3: dout <= 8'b00000000; // 5091 :   0 - 0x0
      13'h13E4: dout <= 8'b00000000; // 5092 :   0 - 0x0
      13'h13E5: dout <= 8'b00000000; // 5093 :   0 - 0x0
      13'h13E6: dout <= 8'b00000000; // 5094 :   0 - 0x0
      13'h13E7: dout <= 8'b00000000; // 5095 :   0 - 0x0
      13'h13E8: dout <= 8'b00000000; // 5096 :   0 - 0x0
      13'h13E9: dout <= 8'b00000000; // 5097 :   0 - 0x0
      13'h13EA: dout <= 8'b00000000; // 5098 :   0 - 0x0
      13'h13EB: dout <= 8'b00000000; // 5099 :   0 - 0x0
      13'h13EC: dout <= 8'b00000000; // 5100 :   0 - 0x0
      13'h13ED: dout <= 8'b00000000; // 5101 :   0 - 0x0
      13'h13EE: dout <= 8'b00000000; // 5102 :   0 - 0x0
      13'h13EF: dout <= 8'b00000000; // 5103 :   0 - 0x0
      13'h13F0: dout <= 8'b00000000; // 5104 :   0 - 0x0 -- Background 0x3f
      13'h13F1: dout <= 8'b00000000; // 5105 :   0 - 0x0
      13'h13F2: dout <= 8'b00000000; // 5106 :   0 - 0x0
      13'h13F3: dout <= 8'b00000000; // 5107 :   0 - 0x0
      13'h13F4: dout <= 8'b00000000; // 5108 :   0 - 0x0
      13'h13F5: dout <= 8'b00000000; // 5109 :   0 - 0x0
      13'h13F6: dout <= 8'b00000000; // 5110 :   0 - 0x0
      13'h13F7: dout <= 8'b00000000; // 5111 :   0 - 0x0
      13'h13F8: dout <= 8'b00000000; // 5112 :   0 - 0x0
      13'h13F9: dout <= 8'b00000000; // 5113 :   0 - 0x0
      13'h13FA: dout <= 8'b00000000; // 5114 :   0 - 0x0
      13'h13FB: dout <= 8'b00000000; // 5115 :   0 - 0x0
      13'h13FC: dout <= 8'b00000000; // 5116 :   0 - 0x0
      13'h13FD: dout <= 8'b00000000; // 5117 :   0 - 0x0
      13'h13FE: dout <= 8'b00000000; // 5118 :   0 - 0x0
      13'h13FF: dout <= 8'b00000000; // 5119 :   0 - 0x0
      13'h1400: dout <= 8'b00000000; // 5120 :   0 - 0x0 -- Background 0x40
      13'h1401: dout <= 8'b00000000; // 5121 :   0 - 0x0
      13'h1402: dout <= 8'b00000000; // 5122 :   0 - 0x0
      13'h1403: dout <= 8'b00000000; // 5123 :   0 - 0x0
      13'h1404: dout <= 8'b00000000; // 5124 :   0 - 0x0
      13'h1405: dout <= 8'b00000000; // 5125 :   0 - 0x0
      13'h1406: dout <= 8'b00000000; // 5126 :   0 - 0x0
      13'h1407: dout <= 8'b00000000; // 5127 :   0 - 0x0
      13'h1408: dout <= 8'b00000000; // 5128 :   0 - 0x0
      13'h1409: dout <= 8'b00000000; // 5129 :   0 - 0x0
      13'h140A: dout <= 8'b00000000; // 5130 :   0 - 0x0
      13'h140B: dout <= 8'b00000000; // 5131 :   0 - 0x0
      13'h140C: dout <= 8'b00000000; // 5132 :   0 - 0x0
      13'h140D: dout <= 8'b00000000; // 5133 :   0 - 0x0
      13'h140E: dout <= 8'b00000000; // 5134 :   0 - 0x0
      13'h140F: dout <= 8'b00000000; // 5135 :   0 - 0x0
      13'h1410: dout <= 8'b00000000; // 5136 :   0 - 0x0 -- Background 0x41
      13'h1411: dout <= 8'b00000000; // 5137 :   0 - 0x0
      13'h1412: dout <= 8'b00000000; // 5138 :   0 - 0x0
      13'h1413: dout <= 8'b00000000; // 5139 :   0 - 0x0
      13'h1414: dout <= 8'b00000000; // 5140 :   0 - 0x0
      13'h1415: dout <= 8'b00000000; // 5141 :   0 - 0x0
      13'h1416: dout <= 8'b00000000; // 5142 :   0 - 0x0
      13'h1417: dout <= 8'b00000000; // 5143 :   0 - 0x0
      13'h1418: dout <= 8'b00000000; // 5144 :   0 - 0x0
      13'h1419: dout <= 8'b00000000; // 5145 :   0 - 0x0
      13'h141A: dout <= 8'b00000000; // 5146 :   0 - 0x0
      13'h141B: dout <= 8'b00000000; // 5147 :   0 - 0x0
      13'h141C: dout <= 8'b00000000; // 5148 :   0 - 0x0
      13'h141D: dout <= 8'b00000000; // 5149 :   0 - 0x0
      13'h141E: dout <= 8'b00000000; // 5150 :   0 - 0x0
      13'h141F: dout <= 8'b00000000; // 5151 :   0 - 0x0
      13'h1420: dout <= 8'b00000000; // 5152 :   0 - 0x0 -- Background 0x42
      13'h1421: dout <= 8'b00000000; // 5153 :   0 - 0x0
      13'h1422: dout <= 8'b00000000; // 5154 :   0 - 0x0
      13'h1423: dout <= 8'b00000000; // 5155 :   0 - 0x0
      13'h1424: dout <= 8'b00000000; // 5156 :   0 - 0x0
      13'h1425: dout <= 8'b00000000; // 5157 :   0 - 0x0
      13'h1426: dout <= 8'b00000000; // 5158 :   0 - 0x0
      13'h1427: dout <= 8'b00000000; // 5159 :   0 - 0x0
      13'h1428: dout <= 8'b00000000; // 5160 :   0 - 0x0
      13'h1429: dout <= 8'b00000000; // 5161 :   0 - 0x0
      13'h142A: dout <= 8'b00000000; // 5162 :   0 - 0x0
      13'h142B: dout <= 8'b00000000; // 5163 :   0 - 0x0
      13'h142C: dout <= 8'b00000000; // 5164 :   0 - 0x0
      13'h142D: dout <= 8'b00000000; // 5165 :   0 - 0x0
      13'h142E: dout <= 8'b00000000; // 5166 :   0 - 0x0
      13'h142F: dout <= 8'b00000000; // 5167 :   0 - 0x0
      13'h1430: dout <= 8'b00000000; // 5168 :   0 - 0x0 -- Background 0x43
      13'h1431: dout <= 8'b00000000; // 5169 :   0 - 0x0
      13'h1432: dout <= 8'b00000000; // 5170 :   0 - 0x0
      13'h1433: dout <= 8'b00000000; // 5171 :   0 - 0x0
      13'h1434: dout <= 8'b00000000; // 5172 :   0 - 0x0
      13'h1435: dout <= 8'b00000000; // 5173 :   0 - 0x0
      13'h1436: dout <= 8'b00000000; // 5174 :   0 - 0x0
      13'h1437: dout <= 8'b00000000; // 5175 :   0 - 0x0
      13'h1438: dout <= 8'b00000000; // 5176 :   0 - 0x0
      13'h1439: dout <= 8'b00000000; // 5177 :   0 - 0x0
      13'h143A: dout <= 8'b00000000; // 5178 :   0 - 0x0
      13'h143B: dout <= 8'b00000000; // 5179 :   0 - 0x0
      13'h143C: dout <= 8'b00000000; // 5180 :   0 - 0x0
      13'h143D: dout <= 8'b00000000; // 5181 :   0 - 0x0
      13'h143E: dout <= 8'b00000000; // 5182 :   0 - 0x0
      13'h143F: dout <= 8'b00000000; // 5183 :   0 - 0x0
      13'h1440: dout <= 8'b00000000; // 5184 :   0 - 0x0 -- Background 0x44
      13'h1441: dout <= 8'b00000000; // 5185 :   0 - 0x0
      13'h1442: dout <= 8'b00000000; // 5186 :   0 - 0x0
      13'h1443: dout <= 8'b00000000; // 5187 :   0 - 0x0
      13'h1444: dout <= 8'b00000000; // 5188 :   0 - 0x0
      13'h1445: dout <= 8'b00000000; // 5189 :   0 - 0x0
      13'h1446: dout <= 8'b00000000; // 5190 :   0 - 0x0
      13'h1447: dout <= 8'b00000000; // 5191 :   0 - 0x0
      13'h1448: dout <= 8'b00000000; // 5192 :   0 - 0x0
      13'h1449: dout <= 8'b00000000; // 5193 :   0 - 0x0
      13'h144A: dout <= 8'b00000000; // 5194 :   0 - 0x0
      13'h144B: dout <= 8'b00000000; // 5195 :   0 - 0x0
      13'h144C: dout <= 8'b00000000; // 5196 :   0 - 0x0
      13'h144D: dout <= 8'b00000000; // 5197 :   0 - 0x0
      13'h144E: dout <= 8'b00000000; // 5198 :   0 - 0x0
      13'h144F: dout <= 8'b00000000; // 5199 :   0 - 0x0
      13'h1450: dout <= 8'b00000000; // 5200 :   0 - 0x0 -- Background 0x45
      13'h1451: dout <= 8'b00000000; // 5201 :   0 - 0x0
      13'h1452: dout <= 8'b00000000; // 5202 :   0 - 0x0
      13'h1453: dout <= 8'b00000000; // 5203 :   0 - 0x0
      13'h1454: dout <= 8'b00000000; // 5204 :   0 - 0x0
      13'h1455: dout <= 8'b00000000; // 5205 :   0 - 0x0
      13'h1456: dout <= 8'b00000000; // 5206 :   0 - 0x0
      13'h1457: dout <= 8'b00000000; // 5207 :   0 - 0x0
      13'h1458: dout <= 8'b00000000; // 5208 :   0 - 0x0
      13'h1459: dout <= 8'b00000000; // 5209 :   0 - 0x0
      13'h145A: dout <= 8'b00000000; // 5210 :   0 - 0x0
      13'h145B: dout <= 8'b00000000; // 5211 :   0 - 0x0
      13'h145C: dout <= 8'b00000000; // 5212 :   0 - 0x0
      13'h145D: dout <= 8'b00000000; // 5213 :   0 - 0x0
      13'h145E: dout <= 8'b00000000; // 5214 :   0 - 0x0
      13'h145F: dout <= 8'b00000000; // 5215 :   0 - 0x0
      13'h1460: dout <= 8'b00000000; // 5216 :   0 - 0x0 -- Background 0x46
      13'h1461: dout <= 8'b00000000; // 5217 :   0 - 0x0
      13'h1462: dout <= 8'b00000000; // 5218 :   0 - 0x0
      13'h1463: dout <= 8'b00000000; // 5219 :   0 - 0x0
      13'h1464: dout <= 8'b00000000; // 5220 :   0 - 0x0
      13'h1465: dout <= 8'b00000000; // 5221 :   0 - 0x0
      13'h1466: dout <= 8'b00000000; // 5222 :   0 - 0x0
      13'h1467: dout <= 8'b00000000; // 5223 :   0 - 0x0
      13'h1468: dout <= 8'b00000000; // 5224 :   0 - 0x0
      13'h1469: dout <= 8'b00000000; // 5225 :   0 - 0x0
      13'h146A: dout <= 8'b00000000; // 5226 :   0 - 0x0
      13'h146B: dout <= 8'b00000000; // 5227 :   0 - 0x0
      13'h146C: dout <= 8'b00000000; // 5228 :   0 - 0x0
      13'h146D: dout <= 8'b00000000; // 5229 :   0 - 0x0
      13'h146E: dout <= 8'b00000000; // 5230 :   0 - 0x0
      13'h146F: dout <= 8'b00000000; // 5231 :   0 - 0x0
      13'h1470: dout <= 8'b00000000; // 5232 :   0 - 0x0 -- Background 0x47
      13'h1471: dout <= 8'b00000000; // 5233 :   0 - 0x0
      13'h1472: dout <= 8'b00000000; // 5234 :   0 - 0x0
      13'h1473: dout <= 8'b00000000; // 5235 :   0 - 0x0
      13'h1474: dout <= 8'b00000000; // 5236 :   0 - 0x0
      13'h1475: dout <= 8'b00000000; // 5237 :   0 - 0x0
      13'h1476: dout <= 8'b00000000; // 5238 :   0 - 0x0
      13'h1477: dout <= 8'b00000000; // 5239 :   0 - 0x0
      13'h1478: dout <= 8'b00000000; // 5240 :   0 - 0x0
      13'h1479: dout <= 8'b00000000; // 5241 :   0 - 0x0
      13'h147A: dout <= 8'b00000000; // 5242 :   0 - 0x0
      13'h147B: dout <= 8'b00000000; // 5243 :   0 - 0x0
      13'h147C: dout <= 8'b00000000; // 5244 :   0 - 0x0
      13'h147D: dout <= 8'b00000000; // 5245 :   0 - 0x0
      13'h147E: dout <= 8'b00000000; // 5246 :   0 - 0x0
      13'h147F: dout <= 8'b00000000; // 5247 :   0 - 0x0
      13'h1480: dout <= 8'b00000000; // 5248 :   0 - 0x0 -- Background 0x48
      13'h1481: dout <= 8'b00000000; // 5249 :   0 - 0x0
      13'h1482: dout <= 8'b00000000; // 5250 :   0 - 0x0
      13'h1483: dout <= 8'b00000000; // 5251 :   0 - 0x0
      13'h1484: dout <= 8'b00000000; // 5252 :   0 - 0x0
      13'h1485: dout <= 8'b00000000; // 5253 :   0 - 0x0
      13'h1486: dout <= 8'b00000000; // 5254 :   0 - 0x0
      13'h1487: dout <= 8'b00000000; // 5255 :   0 - 0x0
      13'h1488: dout <= 8'b00000000; // 5256 :   0 - 0x0
      13'h1489: dout <= 8'b00000000; // 5257 :   0 - 0x0
      13'h148A: dout <= 8'b00000000; // 5258 :   0 - 0x0
      13'h148B: dout <= 8'b00000000; // 5259 :   0 - 0x0
      13'h148C: dout <= 8'b00000000; // 5260 :   0 - 0x0
      13'h148D: dout <= 8'b00000000; // 5261 :   0 - 0x0
      13'h148E: dout <= 8'b00000000; // 5262 :   0 - 0x0
      13'h148F: dout <= 8'b00000000; // 5263 :   0 - 0x0
      13'h1490: dout <= 8'b00000000; // 5264 :   0 - 0x0 -- Background 0x49
      13'h1491: dout <= 8'b00000000; // 5265 :   0 - 0x0
      13'h1492: dout <= 8'b00000000; // 5266 :   0 - 0x0
      13'h1493: dout <= 8'b00000000; // 5267 :   0 - 0x0
      13'h1494: dout <= 8'b00000000; // 5268 :   0 - 0x0
      13'h1495: dout <= 8'b00000000; // 5269 :   0 - 0x0
      13'h1496: dout <= 8'b00000000; // 5270 :   0 - 0x0
      13'h1497: dout <= 8'b00000000; // 5271 :   0 - 0x0
      13'h1498: dout <= 8'b00000000; // 5272 :   0 - 0x0
      13'h1499: dout <= 8'b00000000; // 5273 :   0 - 0x0
      13'h149A: dout <= 8'b00000000; // 5274 :   0 - 0x0
      13'h149B: dout <= 8'b00000000; // 5275 :   0 - 0x0
      13'h149C: dout <= 8'b00000000; // 5276 :   0 - 0x0
      13'h149D: dout <= 8'b00000000; // 5277 :   0 - 0x0
      13'h149E: dout <= 8'b00000000; // 5278 :   0 - 0x0
      13'h149F: dout <= 8'b00000000; // 5279 :   0 - 0x0
      13'h14A0: dout <= 8'b00000000; // 5280 :   0 - 0x0 -- Background 0x4a
      13'h14A1: dout <= 8'b00000000; // 5281 :   0 - 0x0
      13'h14A2: dout <= 8'b00000000; // 5282 :   0 - 0x0
      13'h14A3: dout <= 8'b00000000; // 5283 :   0 - 0x0
      13'h14A4: dout <= 8'b00000000; // 5284 :   0 - 0x0
      13'h14A5: dout <= 8'b00000000; // 5285 :   0 - 0x0
      13'h14A6: dout <= 8'b00000000; // 5286 :   0 - 0x0
      13'h14A7: dout <= 8'b00000000; // 5287 :   0 - 0x0
      13'h14A8: dout <= 8'b00000000; // 5288 :   0 - 0x0
      13'h14A9: dout <= 8'b00000000; // 5289 :   0 - 0x0
      13'h14AA: dout <= 8'b00000000; // 5290 :   0 - 0x0
      13'h14AB: dout <= 8'b00000000; // 5291 :   0 - 0x0
      13'h14AC: dout <= 8'b00000000; // 5292 :   0 - 0x0
      13'h14AD: dout <= 8'b00000000; // 5293 :   0 - 0x0
      13'h14AE: dout <= 8'b00000000; // 5294 :   0 - 0x0
      13'h14AF: dout <= 8'b00000000; // 5295 :   0 - 0x0
      13'h14B0: dout <= 8'b00000000; // 5296 :   0 - 0x0 -- Background 0x4b
      13'h14B1: dout <= 8'b00000000; // 5297 :   0 - 0x0
      13'h14B2: dout <= 8'b00000000; // 5298 :   0 - 0x0
      13'h14B3: dout <= 8'b00000000; // 5299 :   0 - 0x0
      13'h14B4: dout <= 8'b00000000; // 5300 :   0 - 0x0
      13'h14B5: dout <= 8'b00000000; // 5301 :   0 - 0x0
      13'h14B6: dout <= 8'b00000000; // 5302 :   0 - 0x0
      13'h14B7: dout <= 8'b00000000; // 5303 :   0 - 0x0
      13'h14B8: dout <= 8'b00000000; // 5304 :   0 - 0x0
      13'h14B9: dout <= 8'b00000000; // 5305 :   0 - 0x0
      13'h14BA: dout <= 8'b00000000; // 5306 :   0 - 0x0
      13'h14BB: dout <= 8'b00000000; // 5307 :   0 - 0x0
      13'h14BC: dout <= 8'b00000000; // 5308 :   0 - 0x0
      13'h14BD: dout <= 8'b00000000; // 5309 :   0 - 0x0
      13'h14BE: dout <= 8'b00000000; // 5310 :   0 - 0x0
      13'h14BF: dout <= 8'b00000000; // 5311 :   0 - 0x0
      13'h14C0: dout <= 8'b00000000; // 5312 :   0 - 0x0 -- Background 0x4c
      13'h14C1: dout <= 8'b00000000; // 5313 :   0 - 0x0
      13'h14C2: dout <= 8'b00000000; // 5314 :   0 - 0x0
      13'h14C3: dout <= 8'b00000000; // 5315 :   0 - 0x0
      13'h14C4: dout <= 8'b00000000; // 5316 :   0 - 0x0
      13'h14C5: dout <= 8'b00000000; // 5317 :   0 - 0x0
      13'h14C6: dout <= 8'b00000000; // 5318 :   0 - 0x0
      13'h14C7: dout <= 8'b00000000; // 5319 :   0 - 0x0
      13'h14C8: dout <= 8'b00000000; // 5320 :   0 - 0x0
      13'h14C9: dout <= 8'b00000000; // 5321 :   0 - 0x0
      13'h14CA: dout <= 8'b00000000; // 5322 :   0 - 0x0
      13'h14CB: dout <= 8'b00000000; // 5323 :   0 - 0x0
      13'h14CC: dout <= 8'b00000000; // 5324 :   0 - 0x0
      13'h14CD: dout <= 8'b00000000; // 5325 :   0 - 0x0
      13'h14CE: dout <= 8'b00000000; // 5326 :   0 - 0x0
      13'h14CF: dout <= 8'b00000000; // 5327 :   0 - 0x0
      13'h14D0: dout <= 8'b00000000; // 5328 :   0 - 0x0 -- Background 0x4d
      13'h14D1: dout <= 8'b00000000; // 5329 :   0 - 0x0
      13'h14D2: dout <= 8'b00000000; // 5330 :   0 - 0x0
      13'h14D3: dout <= 8'b00000000; // 5331 :   0 - 0x0
      13'h14D4: dout <= 8'b00000000; // 5332 :   0 - 0x0
      13'h14D5: dout <= 8'b00000000; // 5333 :   0 - 0x0
      13'h14D6: dout <= 8'b00000000; // 5334 :   0 - 0x0
      13'h14D7: dout <= 8'b00000000; // 5335 :   0 - 0x0
      13'h14D8: dout <= 8'b00000000; // 5336 :   0 - 0x0
      13'h14D9: dout <= 8'b00000000; // 5337 :   0 - 0x0
      13'h14DA: dout <= 8'b00000000; // 5338 :   0 - 0x0
      13'h14DB: dout <= 8'b00000000; // 5339 :   0 - 0x0
      13'h14DC: dout <= 8'b00000000; // 5340 :   0 - 0x0
      13'h14DD: dout <= 8'b00000000; // 5341 :   0 - 0x0
      13'h14DE: dout <= 8'b00000000; // 5342 :   0 - 0x0
      13'h14DF: dout <= 8'b00000000; // 5343 :   0 - 0x0
      13'h14E0: dout <= 8'b00000000; // 5344 :   0 - 0x0 -- Background 0x4e
      13'h14E1: dout <= 8'b00000000; // 5345 :   0 - 0x0
      13'h14E2: dout <= 8'b00000000; // 5346 :   0 - 0x0
      13'h14E3: dout <= 8'b00000000; // 5347 :   0 - 0x0
      13'h14E4: dout <= 8'b00000000; // 5348 :   0 - 0x0
      13'h14E5: dout <= 8'b00000000; // 5349 :   0 - 0x0
      13'h14E6: dout <= 8'b00000000; // 5350 :   0 - 0x0
      13'h14E7: dout <= 8'b00000000; // 5351 :   0 - 0x0
      13'h14E8: dout <= 8'b00000000; // 5352 :   0 - 0x0
      13'h14E9: dout <= 8'b00000000; // 5353 :   0 - 0x0
      13'h14EA: dout <= 8'b00000000; // 5354 :   0 - 0x0
      13'h14EB: dout <= 8'b00000000; // 5355 :   0 - 0x0
      13'h14EC: dout <= 8'b00000000; // 5356 :   0 - 0x0
      13'h14ED: dout <= 8'b00000000; // 5357 :   0 - 0x0
      13'h14EE: dout <= 8'b00000000; // 5358 :   0 - 0x0
      13'h14EF: dout <= 8'b00000000; // 5359 :   0 - 0x0
      13'h14F0: dout <= 8'b00000000; // 5360 :   0 - 0x0 -- Background 0x4f
      13'h14F1: dout <= 8'b00000000; // 5361 :   0 - 0x0
      13'h14F2: dout <= 8'b00000000; // 5362 :   0 - 0x0
      13'h14F3: dout <= 8'b00000000; // 5363 :   0 - 0x0
      13'h14F4: dout <= 8'b00000000; // 5364 :   0 - 0x0
      13'h14F5: dout <= 8'b00000000; // 5365 :   0 - 0x0
      13'h14F6: dout <= 8'b00000000; // 5366 :   0 - 0x0
      13'h14F7: dout <= 8'b00000000; // 5367 :   0 - 0x0
      13'h14F8: dout <= 8'b00000000; // 5368 :   0 - 0x0
      13'h14F9: dout <= 8'b00000000; // 5369 :   0 - 0x0
      13'h14FA: dout <= 8'b00000000; // 5370 :   0 - 0x0
      13'h14FB: dout <= 8'b00000000; // 5371 :   0 - 0x0
      13'h14FC: dout <= 8'b00000000; // 5372 :   0 - 0x0
      13'h14FD: dout <= 8'b00000000; // 5373 :   0 - 0x0
      13'h14FE: dout <= 8'b00000000; // 5374 :   0 - 0x0
      13'h14FF: dout <= 8'b00000000; // 5375 :   0 - 0x0
      13'h1500: dout <= 8'b00000000; // 5376 :   0 - 0x0 -- Background 0x50
      13'h1501: dout <= 8'b00000000; // 5377 :   0 - 0x0
      13'h1502: dout <= 8'b00000000; // 5378 :   0 - 0x0
      13'h1503: dout <= 8'b00000000; // 5379 :   0 - 0x0
      13'h1504: dout <= 8'b00000000; // 5380 :   0 - 0x0
      13'h1505: dout <= 8'b00000000; // 5381 :   0 - 0x0
      13'h1506: dout <= 8'b00000000; // 5382 :   0 - 0x0
      13'h1507: dout <= 8'b00000000; // 5383 :   0 - 0x0
      13'h1508: dout <= 8'b00000000; // 5384 :   0 - 0x0
      13'h1509: dout <= 8'b00000000; // 5385 :   0 - 0x0
      13'h150A: dout <= 8'b00000000; // 5386 :   0 - 0x0
      13'h150B: dout <= 8'b00000000; // 5387 :   0 - 0x0
      13'h150C: dout <= 8'b00000000; // 5388 :   0 - 0x0
      13'h150D: dout <= 8'b00000000; // 5389 :   0 - 0x0
      13'h150E: dout <= 8'b00000000; // 5390 :   0 - 0x0
      13'h150F: dout <= 8'b00000000; // 5391 :   0 - 0x0
      13'h1510: dout <= 8'b00000000; // 5392 :   0 - 0x0 -- Background 0x51
      13'h1511: dout <= 8'b00000000; // 5393 :   0 - 0x0
      13'h1512: dout <= 8'b00000000; // 5394 :   0 - 0x0
      13'h1513: dout <= 8'b00000000; // 5395 :   0 - 0x0
      13'h1514: dout <= 8'b00000000; // 5396 :   0 - 0x0
      13'h1515: dout <= 8'b00000000; // 5397 :   0 - 0x0
      13'h1516: dout <= 8'b00000000; // 5398 :   0 - 0x0
      13'h1517: dout <= 8'b00000000; // 5399 :   0 - 0x0
      13'h1518: dout <= 8'b00000000; // 5400 :   0 - 0x0
      13'h1519: dout <= 8'b00000000; // 5401 :   0 - 0x0
      13'h151A: dout <= 8'b00000000; // 5402 :   0 - 0x0
      13'h151B: dout <= 8'b00000000; // 5403 :   0 - 0x0
      13'h151C: dout <= 8'b00000000; // 5404 :   0 - 0x0
      13'h151D: dout <= 8'b00000000; // 5405 :   0 - 0x0
      13'h151E: dout <= 8'b00000000; // 5406 :   0 - 0x0
      13'h151F: dout <= 8'b00000000; // 5407 :   0 - 0x0
      13'h1520: dout <= 8'b00000000; // 5408 :   0 - 0x0 -- Background 0x52
      13'h1521: dout <= 8'b00000000; // 5409 :   0 - 0x0
      13'h1522: dout <= 8'b00000000; // 5410 :   0 - 0x0
      13'h1523: dout <= 8'b00000000; // 5411 :   0 - 0x0
      13'h1524: dout <= 8'b00000000; // 5412 :   0 - 0x0
      13'h1525: dout <= 8'b00000000; // 5413 :   0 - 0x0
      13'h1526: dout <= 8'b00000000; // 5414 :   0 - 0x0
      13'h1527: dout <= 8'b00000000; // 5415 :   0 - 0x0
      13'h1528: dout <= 8'b00000000; // 5416 :   0 - 0x0
      13'h1529: dout <= 8'b00000000; // 5417 :   0 - 0x0
      13'h152A: dout <= 8'b00000000; // 5418 :   0 - 0x0
      13'h152B: dout <= 8'b00000000; // 5419 :   0 - 0x0
      13'h152C: dout <= 8'b00000000; // 5420 :   0 - 0x0
      13'h152D: dout <= 8'b00000000; // 5421 :   0 - 0x0
      13'h152E: dout <= 8'b00000000; // 5422 :   0 - 0x0
      13'h152F: dout <= 8'b00000000; // 5423 :   0 - 0x0
      13'h1530: dout <= 8'b00000000; // 5424 :   0 - 0x0 -- Background 0x53
      13'h1531: dout <= 8'b00000000; // 5425 :   0 - 0x0
      13'h1532: dout <= 8'b00000000; // 5426 :   0 - 0x0
      13'h1533: dout <= 8'b00000000; // 5427 :   0 - 0x0
      13'h1534: dout <= 8'b00000000; // 5428 :   0 - 0x0
      13'h1535: dout <= 8'b00000000; // 5429 :   0 - 0x0
      13'h1536: dout <= 8'b00000000; // 5430 :   0 - 0x0
      13'h1537: dout <= 8'b00000000; // 5431 :   0 - 0x0
      13'h1538: dout <= 8'b00000000; // 5432 :   0 - 0x0
      13'h1539: dout <= 8'b00000000; // 5433 :   0 - 0x0
      13'h153A: dout <= 8'b00000000; // 5434 :   0 - 0x0
      13'h153B: dout <= 8'b00000000; // 5435 :   0 - 0x0
      13'h153C: dout <= 8'b00000000; // 5436 :   0 - 0x0
      13'h153D: dout <= 8'b00000000; // 5437 :   0 - 0x0
      13'h153E: dout <= 8'b00000000; // 5438 :   0 - 0x0
      13'h153F: dout <= 8'b00000000; // 5439 :   0 - 0x0
      13'h1540: dout <= 8'b00000000; // 5440 :   0 - 0x0 -- Background 0x54
      13'h1541: dout <= 8'b00000000; // 5441 :   0 - 0x0
      13'h1542: dout <= 8'b00000000; // 5442 :   0 - 0x0
      13'h1543: dout <= 8'b00000000; // 5443 :   0 - 0x0
      13'h1544: dout <= 8'b00000000; // 5444 :   0 - 0x0
      13'h1545: dout <= 8'b00000000; // 5445 :   0 - 0x0
      13'h1546: dout <= 8'b00000000; // 5446 :   0 - 0x0
      13'h1547: dout <= 8'b00000000; // 5447 :   0 - 0x0
      13'h1548: dout <= 8'b00000000; // 5448 :   0 - 0x0
      13'h1549: dout <= 8'b00000000; // 5449 :   0 - 0x0
      13'h154A: dout <= 8'b00000000; // 5450 :   0 - 0x0
      13'h154B: dout <= 8'b00000000; // 5451 :   0 - 0x0
      13'h154C: dout <= 8'b00000000; // 5452 :   0 - 0x0
      13'h154D: dout <= 8'b00000000; // 5453 :   0 - 0x0
      13'h154E: dout <= 8'b00000000; // 5454 :   0 - 0x0
      13'h154F: dout <= 8'b00000000; // 5455 :   0 - 0x0
      13'h1550: dout <= 8'b00000000; // 5456 :   0 - 0x0 -- Background 0x55
      13'h1551: dout <= 8'b00000000; // 5457 :   0 - 0x0
      13'h1552: dout <= 8'b00000000; // 5458 :   0 - 0x0
      13'h1553: dout <= 8'b00000000; // 5459 :   0 - 0x0
      13'h1554: dout <= 8'b00000000; // 5460 :   0 - 0x0
      13'h1555: dout <= 8'b00000000; // 5461 :   0 - 0x0
      13'h1556: dout <= 8'b00000000; // 5462 :   0 - 0x0
      13'h1557: dout <= 8'b00000000; // 5463 :   0 - 0x0
      13'h1558: dout <= 8'b00000000; // 5464 :   0 - 0x0
      13'h1559: dout <= 8'b00000000; // 5465 :   0 - 0x0
      13'h155A: dout <= 8'b00000000; // 5466 :   0 - 0x0
      13'h155B: dout <= 8'b00000000; // 5467 :   0 - 0x0
      13'h155C: dout <= 8'b00000000; // 5468 :   0 - 0x0
      13'h155D: dout <= 8'b00000000; // 5469 :   0 - 0x0
      13'h155E: dout <= 8'b00000000; // 5470 :   0 - 0x0
      13'h155F: dout <= 8'b00000000; // 5471 :   0 - 0x0
      13'h1560: dout <= 8'b00000000; // 5472 :   0 - 0x0 -- Background 0x56
      13'h1561: dout <= 8'b00000000; // 5473 :   0 - 0x0
      13'h1562: dout <= 8'b00000000; // 5474 :   0 - 0x0
      13'h1563: dout <= 8'b00000000; // 5475 :   0 - 0x0
      13'h1564: dout <= 8'b00000000; // 5476 :   0 - 0x0
      13'h1565: dout <= 8'b00000000; // 5477 :   0 - 0x0
      13'h1566: dout <= 8'b00000000; // 5478 :   0 - 0x0
      13'h1567: dout <= 8'b00000000; // 5479 :   0 - 0x0
      13'h1568: dout <= 8'b00000000; // 5480 :   0 - 0x0
      13'h1569: dout <= 8'b00000000; // 5481 :   0 - 0x0
      13'h156A: dout <= 8'b00000000; // 5482 :   0 - 0x0
      13'h156B: dout <= 8'b00000000; // 5483 :   0 - 0x0
      13'h156C: dout <= 8'b00000000; // 5484 :   0 - 0x0
      13'h156D: dout <= 8'b00000000; // 5485 :   0 - 0x0
      13'h156E: dout <= 8'b00000000; // 5486 :   0 - 0x0
      13'h156F: dout <= 8'b00000000; // 5487 :   0 - 0x0
      13'h1570: dout <= 8'b00000000; // 5488 :   0 - 0x0 -- Background 0x57
      13'h1571: dout <= 8'b00000000; // 5489 :   0 - 0x0
      13'h1572: dout <= 8'b00000000; // 5490 :   0 - 0x0
      13'h1573: dout <= 8'b00000000; // 5491 :   0 - 0x0
      13'h1574: dout <= 8'b00000000; // 5492 :   0 - 0x0
      13'h1575: dout <= 8'b00000000; // 5493 :   0 - 0x0
      13'h1576: dout <= 8'b00000000; // 5494 :   0 - 0x0
      13'h1577: dout <= 8'b00000000; // 5495 :   0 - 0x0
      13'h1578: dout <= 8'b00000000; // 5496 :   0 - 0x0
      13'h1579: dout <= 8'b00000000; // 5497 :   0 - 0x0
      13'h157A: dout <= 8'b00000000; // 5498 :   0 - 0x0
      13'h157B: dout <= 8'b00000000; // 5499 :   0 - 0x0
      13'h157C: dout <= 8'b00000000; // 5500 :   0 - 0x0
      13'h157D: dout <= 8'b00000000; // 5501 :   0 - 0x0
      13'h157E: dout <= 8'b00000000; // 5502 :   0 - 0x0
      13'h157F: dout <= 8'b00000000; // 5503 :   0 - 0x0
      13'h1580: dout <= 8'b00000000; // 5504 :   0 - 0x0 -- Background 0x58
      13'h1581: dout <= 8'b00000000; // 5505 :   0 - 0x0
      13'h1582: dout <= 8'b00000000; // 5506 :   0 - 0x0
      13'h1583: dout <= 8'b00000000; // 5507 :   0 - 0x0
      13'h1584: dout <= 8'b00000000; // 5508 :   0 - 0x0
      13'h1585: dout <= 8'b00000000; // 5509 :   0 - 0x0
      13'h1586: dout <= 8'b00000000; // 5510 :   0 - 0x0
      13'h1587: dout <= 8'b00000000; // 5511 :   0 - 0x0
      13'h1588: dout <= 8'b00000000; // 5512 :   0 - 0x0
      13'h1589: dout <= 8'b00000000; // 5513 :   0 - 0x0
      13'h158A: dout <= 8'b00000000; // 5514 :   0 - 0x0
      13'h158B: dout <= 8'b00000000; // 5515 :   0 - 0x0
      13'h158C: dout <= 8'b00000000; // 5516 :   0 - 0x0
      13'h158D: dout <= 8'b00000000; // 5517 :   0 - 0x0
      13'h158E: dout <= 8'b00000000; // 5518 :   0 - 0x0
      13'h158F: dout <= 8'b00000000; // 5519 :   0 - 0x0
      13'h1590: dout <= 8'b00000000; // 5520 :   0 - 0x0 -- Background 0x59
      13'h1591: dout <= 8'b00000000; // 5521 :   0 - 0x0
      13'h1592: dout <= 8'b00000000; // 5522 :   0 - 0x0
      13'h1593: dout <= 8'b00000000; // 5523 :   0 - 0x0
      13'h1594: dout <= 8'b00000000; // 5524 :   0 - 0x0
      13'h1595: dout <= 8'b00000000; // 5525 :   0 - 0x0
      13'h1596: dout <= 8'b00000000; // 5526 :   0 - 0x0
      13'h1597: dout <= 8'b00000000; // 5527 :   0 - 0x0
      13'h1598: dout <= 8'b00000000; // 5528 :   0 - 0x0
      13'h1599: dout <= 8'b00000000; // 5529 :   0 - 0x0
      13'h159A: dout <= 8'b00000000; // 5530 :   0 - 0x0
      13'h159B: dout <= 8'b00000000; // 5531 :   0 - 0x0
      13'h159C: dout <= 8'b00000000; // 5532 :   0 - 0x0
      13'h159D: dout <= 8'b00000000; // 5533 :   0 - 0x0
      13'h159E: dout <= 8'b00000000; // 5534 :   0 - 0x0
      13'h159F: dout <= 8'b00000000; // 5535 :   0 - 0x0
      13'h15A0: dout <= 8'b00000000; // 5536 :   0 - 0x0 -- Background 0x5a
      13'h15A1: dout <= 8'b00000000; // 5537 :   0 - 0x0
      13'h15A2: dout <= 8'b00000000; // 5538 :   0 - 0x0
      13'h15A3: dout <= 8'b00000000; // 5539 :   0 - 0x0
      13'h15A4: dout <= 8'b00000000; // 5540 :   0 - 0x0
      13'h15A5: dout <= 8'b00000000; // 5541 :   0 - 0x0
      13'h15A6: dout <= 8'b00000000; // 5542 :   0 - 0x0
      13'h15A7: dout <= 8'b00000000; // 5543 :   0 - 0x0
      13'h15A8: dout <= 8'b00000000; // 5544 :   0 - 0x0
      13'h15A9: dout <= 8'b00000000; // 5545 :   0 - 0x0
      13'h15AA: dout <= 8'b00000000; // 5546 :   0 - 0x0
      13'h15AB: dout <= 8'b00000000; // 5547 :   0 - 0x0
      13'h15AC: dout <= 8'b00000000; // 5548 :   0 - 0x0
      13'h15AD: dout <= 8'b00000000; // 5549 :   0 - 0x0
      13'h15AE: dout <= 8'b00000000; // 5550 :   0 - 0x0
      13'h15AF: dout <= 8'b00000000; // 5551 :   0 - 0x0
      13'h15B0: dout <= 8'b00000000; // 5552 :   0 - 0x0 -- Background 0x5b
      13'h15B1: dout <= 8'b00000000; // 5553 :   0 - 0x0
      13'h15B2: dout <= 8'b00000000; // 5554 :   0 - 0x0
      13'h15B3: dout <= 8'b00000000; // 5555 :   0 - 0x0
      13'h15B4: dout <= 8'b00000000; // 5556 :   0 - 0x0
      13'h15B5: dout <= 8'b00000000; // 5557 :   0 - 0x0
      13'h15B6: dout <= 8'b00000000; // 5558 :   0 - 0x0
      13'h15B7: dout <= 8'b00000000; // 5559 :   0 - 0x0
      13'h15B8: dout <= 8'b00000000; // 5560 :   0 - 0x0
      13'h15B9: dout <= 8'b00000000; // 5561 :   0 - 0x0
      13'h15BA: dout <= 8'b00000000; // 5562 :   0 - 0x0
      13'h15BB: dout <= 8'b00000000; // 5563 :   0 - 0x0
      13'h15BC: dout <= 8'b00000000; // 5564 :   0 - 0x0
      13'h15BD: dout <= 8'b00000000; // 5565 :   0 - 0x0
      13'h15BE: dout <= 8'b00000000; // 5566 :   0 - 0x0
      13'h15BF: dout <= 8'b00000000; // 5567 :   0 - 0x0
      13'h15C0: dout <= 8'b00000000; // 5568 :   0 - 0x0 -- Background 0x5c
      13'h15C1: dout <= 8'b00000000; // 5569 :   0 - 0x0
      13'h15C2: dout <= 8'b00000000; // 5570 :   0 - 0x0
      13'h15C3: dout <= 8'b00000000; // 5571 :   0 - 0x0
      13'h15C4: dout <= 8'b00000000; // 5572 :   0 - 0x0
      13'h15C5: dout <= 8'b00000000; // 5573 :   0 - 0x0
      13'h15C6: dout <= 8'b00000000; // 5574 :   0 - 0x0
      13'h15C7: dout <= 8'b00000000; // 5575 :   0 - 0x0
      13'h15C8: dout <= 8'b00000000; // 5576 :   0 - 0x0
      13'h15C9: dout <= 8'b00000000; // 5577 :   0 - 0x0
      13'h15CA: dout <= 8'b00000000; // 5578 :   0 - 0x0
      13'h15CB: dout <= 8'b00000000; // 5579 :   0 - 0x0
      13'h15CC: dout <= 8'b00000000; // 5580 :   0 - 0x0
      13'h15CD: dout <= 8'b00000000; // 5581 :   0 - 0x0
      13'h15CE: dout <= 8'b00000000; // 5582 :   0 - 0x0
      13'h15CF: dout <= 8'b00000000; // 5583 :   0 - 0x0
      13'h15D0: dout <= 8'b00000000; // 5584 :   0 - 0x0 -- Background 0x5d
      13'h15D1: dout <= 8'b00000000; // 5585 :   0 - 0x0
      13'h15D2: dout <= 8'b00000000; // 5586 :   0 - 0x0
      13'h15D3: dout <= 8'b00000000; // 5587 :   0 - 0x0
      13'h15D4: dout <= 8'b00000000; // 5588 :   0 - 0x0
      13'h15D5: dout <= 8'b00000000; // 5589 :   0 - 0x0
      13'h15D6: dout <= 8'b00000000; // 5590 :   0 - 0x0
      13'h15D7: dout <= 8'b00000000; // 5591 :   0 - 0x0
      13'h15D8: dout <= 8'b00000000; // 5592 :   0 - 0x0
      13'h15D9: dout <= 8'b00000000; // 5593 :   0 - 0x0
      13'h15DA: dout <= 8'b00000000; // 5594 :   0 - 0x0
      13'h15DB: dout <= 8'b00000000; // 5595 :   0 - 0x0
      13'h15DC: dout <= 8'b00000000; // 5596 :   0 - 0x0
      13'h15DD: dout <= 8'b00000000; // 5597 :   0 - 0x0
      13'h15DE: dout <= 8'b00000000; // 5598 :   0 - 0x0
      13'h15DF: dout <= 8'b00000000; // 5599 :   0 - 0x0
      13'h15E0: dout <= 8'b00000000; // 5600 :   0 - 0x0 -- Background 0x5e
      13'h15E1: dout <= 8'b00000000; // 5601 :   0 - 0x0
      13'h15E2: dout <= 8'b00000000; // 5602 :   0 - 0x0
      13'h15E3: dout <= 8'b00000000; // 5603 :   0 - 0x0
      13'h15E4: dout <= 8'b00000000; // 5604 :   0 - 0x0
      13'h15E5: dout <= 8'b00000000; // 5605 :   0 - 0x0
      13'h15E6: dout <= 8'b00000000; // 5606 :   0 - 0x0
      13'h15E7: dout <= 8'b00000000; // 5607 :   0 - 0x0
      13'h15E8: dout <= 8'b00000000; // 5608 :   0 - 0x0
      13'h15E9: dout <= 8'b00000000; // 5609 :   0 - 0x0
      13'h15EA: dout <= 8'b00000000; // 5610 :   0 - 0x0
      13'h15EB: dout <= 8'b00000000; // 5611 :   0 - 0x0
      13'h15EC: dout <= 8'b00000000; // 5612 :   0 - 0x0
      13'h15ED: dout <= 8'b00000000; // 5613 :   0 - 0x0
      13'h15EE: dout <= 8'b00000000; // 5614 :   0 - 0x0
      13'h15EF: dout <= 8'b00000000; // 5615 :   0 - 0x0
      13'h15F0: dout <= 8'b00000000; // 5616 :   0 - 0x0 -- Background 0x5f
      13'h15F1: dout <= 8'b00000000; // 5617 :   0 - 0x0
      13'h15F2: dout <= 8'b00000000; // 5618 :   0 - 0x0
      13'h15F3: dout <= 8'b00000000; // 5619 :   0 - 0x0
      13'h15F4: dout <= 8'b00000000; // 5620 :   0 - 0x0
      13'h15F5: dout <= 8'b00000000; // 5621 :   0 - 0x0
      13'h15F6: dout <= 8'b00000000; // 5622 :   0 - 0x0
      13'h15F7: dout <= 8'b00000000; // 5623 :   0 - 0x0
      13'h15F8: dout <= 8'b00000000; // 5624 :   0 - 0x0
      13'h15F9: dout <= 8'b00000000; // 5625 :   0 - 0x0
      13'h15FA: dout <= 8'b00000000; // 5626 :   0 - 0x0
      13'h15FB: dout <= 8'b00000000; // 5627 :   0 - 0x0
      13'h15FC: dout <= 8'b00000000; // 5628 :   0 - 0x0
      13'h15FD: dout <= 8'b00000000; // 5629 :   0 - 0x0
      13'h15FE: dout <= 8'b00000000; // 5630 :   0 - 0x0
      13'h15FF: dout <= 8'b00000000; // 5631 :   0 - 0x0
      13'h1600: dout <= 8'b00000000; // 5632 :   0 - 0x0 -- Background 0x60
      13'h1601: dout <= 8'b00000000; // 5633 :   0 - 0x0
      13'h1602: dout <= 8'b00000000; // 5634 :   0 - 0x0
      13'h1603: dout <= 8'b00000000; // 5635 :   0 - 0x0
      13'h1604: dout <= 8'b00000000; // 5636 :   0 - 0x0
      13'h1605: dout <= 8'b00000000; // 5637 :   0 - 0x0
      13'h1606: dout <= 8'b00000000; // 5638 :   0 - 0x0
      13'h1607: dout <= 8'b00000000; // 5639 :   0 - 0x0
      13'h1608: dout <= 8'b00000000; // 5640 :   0 - 0x0
      13'h1609: dout <= 8'b00000000; // 5641 :   0 - 0x0
      13'h160A: dout <= 8'b00000000; // 5642 :   0 - 0x0
      13'h160B: dout <= 8'b00000000; // 5643 :   0 - 0x0
      13'h160C: dout <= 8'b00000000; // 5644 :   0 - 0x0
      13'h160D: dout <= 8'b00000000; // 5645 :   0 - 0x0
      13'h160E: dout <= 8'b00000000; // 5646 :   0 - 0x0
      13'h160F: dout <= 8'b00000000; // 5647 :   0 - 0x0
      13'h1610: dout <= 8'b00000000; // 5648 :   0 - 0x0 -- Background 0x61
      13'h1611: dout <= 8'b00000000; // 5649 :   0 - 0x0
      13'h1612: dout <= 8'b00000000; // 5650 :   0 - 0x0
      13'h1613: dout <= 8'b00000000; // 5651 :   0 - 0x0
      13'h1614: dout <= 8'b00000000; // 5652 :   0 - 0x0
      13'h1615: dout <= 8'b00000000; // 5653 :   0 - 0x0
      13'h1616: dout <= 8'b00000000; // 5654 :   0 - 0x0
      13'h1617: dout <= 8'b00000000; // 5655 :   0 - 0x0
      13'h1618: dout <= 8'b00000000; // 5656 :   0 - 0x0
      13'h1619: dout <= 8'b00000000; // 5657 :   0 - 0x0
      13'h161A: dout <= 8'b00000000; // 5658 :   0 - 0x0
      13'h161B: dout <= 8'b00000000; // 5659 :   0 - 0x0
      13'h161C: dout <= 8'b00000000; // 5660 :   0 - 0x0
      13'h161D: dout <= 8'b00000000; // 5661 :   0 - 0x0
      13'h161E: dout <= 8'b00000000; // 5662 :   0 - 0x0
      13'h161F: dout <= 8'b00000000; // 5663 :   0 - 0x0
      13'h1620: dout <= 8'b00000000; // 5664 :   0 - 0x0 -- Background 0x62
      13'h1621: dout <= 8'b00000000; // 5665 :   0 - 0x0
      13'h1622: dout <= 8'b00000000; // 5666 :   0 - 0x0
      13'h1623: dout <= 8'b00000000; // 5667 :   0 - 0x0
      13'h1624: dout <= 8'b00000000; // 5668 :   0 - 0x0
      13'h1625: dout <= 8'b00000000; // 5669 :   0 - 0x0
      13'h1626: dout <= 8'b00000000; // 5670 :   0 - 0x0
      13'h1627: dout <= 8'b00000000; // 5671 :   0 - 0x0
      13'h1628: dout <= 8'b00000000; // 5672 :   0 - 0x0
      13'h1629: dout <= 8'b00000000; // 5673 :   0 - 0x0
      13'h162A: dout <= 8'b00000000; // 5674 :   0 - 0x0
      13'h162B: dout <= 8'b00000000; // 5675 :   0 - 0x0
      13'h162C: dout <= 8'b00000000; // 5676 :   0 - 0x0
      13'h162D: dout <= 8'b00000000; // 5677 :   0 - 0x0
      13'h162E: dout <= 8'b00000000; // 5678 :   0 - 0x0
      13'h162F: dout <= 8'b00000000; // 5679 :   0 - 0x0
      13'h1630: dout <= 8'b00000000; // 5680 :   0 - 0x0 -- Background 0x63
      13'h1631: dout <= 8'b00000000; // 5681 :   0 - 0x0
      13'h1632: dout <= 8'b00000000; // 5682 :   0 - 0x0
      13'h1633: dout <= 8'b00000000; // 5683 :   0 - 0x0
      13'h1634: dout <= 8'b00000000; // 5684 :   0 - 0x0
      13'h1635: dout <= 8'b00000000; // 5685 :   0 - 0x0
      13'h1636: dout <= 8'b00000000; // 5686 :   0 - 0x0
      13'h1637: dout <= 8'b00000000; // 5687 :   0 - 0x0
      13'h1638: dout <= 8'b00000000; // 5688 :   0 - 0x0
      13'h1639: dout <= 8'b00000000; // 5689 :   0 - 0x0
      13'h163A: dout <= 8'b00000000; // 5690 :   0 - 0x0
      13'h163B: dout <= 8'b00000000; // 5691 :   0 - 0x0
      13'h163C: dout <= 8'b00000000; // 5692 :   0 - 0x0
      13'h163D: dout <= 8'b00000000; // 5693 :   0 - 0x0
      13'h163E: dout <= 8'b00000000; // 5694 :   0 - 0x0
      13'h163F: dout <= 8'b00000000; // 5695 :   0 - 0x0
      13'h1640: dout <= 8'b00000000; // 5696 :   0 - 0x0 -- Background 0x64
      13'h1641: dout <= 8'b00000000; // 5697 :   0 - 0x0
      13'h1642: dout <= 8'b00000000; // 5698 :   0 - 0x0
      13'h1643: dout <= 8'b00000000; // 5699 :   0 - 0x0
      13'h1644: dout <= 8'b00000000; // 5700 :   0 - 0x0
      13'h1645: dout <= 8'b00000000; // 5701 :   0 - 0x0
      13'h1646: dout <= 8'b00000000; // 5702 :   0 - 0x0
      13'h1647: dout <= 8'b00000000; // 5703 :   0 - 0x0
      13'h1648: dout <= 8'b00000000; // 5704 :   0 - 0x0
      13'h1649: dout <= 8'b00000000; // 5705 :   0 - 0x0
      13'h164A: dout <= 8'b00000000; // 5706 :   0 - 0x0
      13'h164B: dout <= 8'b00000000; // 5707 :   0 - 0x0
      13'h164C: dout <= 8'b00000000; // 5708 :   0 - 0x0
      13'h164D: dout <= 8'b00000000; // 5709 :   0 - 0x0
      13'h164E: dout <= 8'b00000000; // 5710 :   0 - 0x0
      13'h164F: dout <= 8'b00000000; // 5711 :   0 - 0x0
      13'h1650: dout <= 8'b00000000; // 5712 :   0 - 0x0 -- Background 0x65
      13'h1651: dout <= 8'b00000000; // 5713 :   0 - 0x0
      13'h1652: dout <= 8'b00000000; // 5714 :   0 - 0x0
      13'h1653: dout <= 8'b00000000; // 5715 :   0 - 0x0
      13'h1654: dout <= 8'b00000000; // 5716 :   0 - 0x0
      13'h1655: dout <= 8'b00000000; // 5717 :   0 - 0x0
      13'h1656: dout <= 8'b00000000; // 5718 :   0 - 0x0
      13'h1657: dout <= 8'b00000000; // 5719 :   0 - 0x0
      13'h1658: dout <= 8'b00000000; // 5720 :   0 - 0x0
      13'h1659: dout <= 8'b00000000; // 5721 :   0 - 0x0
      13'h165A: dout <= 8'b00000000; // 5722 :   0 - 0x0
      13'h165B: dout <= 8'b00000000; // 5723 :   0 - 0x0
      13'h165C: dout <= 8'b00000000; // 5724 :   0 - 0x0
      13'h165D: dout <= 8'b00000000; // 5725 :   0 - 0x0
      13'h165E: dout <= 8'b00000000; // 5726 :   0 - 0x0
      13'h165F: dout <= 8'b00000000; // 5727 :   0 - 0x0
      13'h1660: dout <= 8'b00000000; // 5728 :   0 - 0x0 -- Background 0x66
      13'h1661: dout <= 8'b00000000; // 5729 :   0 - 0x0
      13'h1662: dout <= 8'b00000000; // 5730 :   0 - 0x0
      13'h1663: dout <= 8'b00000000; // 5731 :   0 - 0x0
      13'h1664: dout <= 8'b00000000; // 5732 :   0 - 0x0
      13'h1665: dout <= 8'b00000000; // 5733 :   0 - 0x0
      13'h1666: dout <= 8'b00000000; // 5734 :   0 - 0x0
      13'h1667: dout <= 8'b00000000; // 5735 :   0 - 0x0
      13'h1668: dout <= 8'b00000000; // 5736 :   0 - 0x0
      13'h1669: dout <= 8'b00000000; // 5737 :   0 - 0x0
      13'h166A: dout <= 8'b00000000; // 5738 :   0 - 0x0
      13'h166B: dout <= 8'b00000000; // 5739 :   0 - 0x0
      13'h166C: dout <= 8'b00000000; // 5740 :   0 - 0x0
      13'h166D: dout <= 8'b00000000; // 5741 :   0 - 0x0
      13'h166E: dout <= 8'b00000000; // 5742 :   0 - 0x0
      13'h166F: dout <= 8'b00000000; // 5743 :   0 - 0x0
      13'h1670: dout <= 8'b00000000; // 5744 :   0 - 0x0 -- Background 0x67
      13'h1671: dout <= 8'b00000000; // 5745 :   0 - 0x0
      13'h1672: dout <= 8'b00000000; // 5746 :   0 - 0x0
      13'h1673: dout <= 8'b00000000; // 5747 :   0 - 0x0
      13'h1674: dout <= 8'b00000000; // 5748 :   0 - 0x0
      13'h1675: dout <= 8'b00000000; // 5749 :   0 - 0x0
      13'h1676: dout <= 8'b00000000; // 5750 :   0 - 0x0
      13'h1677: dout <= 8'b00000000; // 5751 :   0 - 0x0
      13'h1678: dout <= 8'b00000000; // 5752 :   0 - 0x0
      13'h1679: dout <= 8'b00000000; // 5753 :   0 - 0x0
      13'h167A: dout <= 8'b00000000; // 5754 :   0 - 0x0
      13'h167B: dout <= 8'b00000000; // 5755 :   0 - 0x0
      13'h167C: dout <= 8'b00000000; // 5756 :   0 - 0x0
      13'h167D: dout <= 8'b00000000; // 5757 :   0 - 0x0
      13'h167E: dout <= 8'b00000000; // 5758 :   0 - 0x0
      13'h167F: dout <= 8'b00000000; // 5759 :   0 - 0x0
      13'h1680: dout <= 8'b00000000; // 5760 :   0 - 0x0 -- Background 0x68
      13'h1681: dout <= 8'b00000000; // 5761 :   0 - 0x0
      13'h1682: dout <= 8'b00000000; // 5762 :   0 - 0x0
      13'h1683: dout <= 8'b00000000; // 5763 :   0 - 0x0
      13'h1684: dout <= 8'b00000000; // 5764 :   0 - 0x0
      13'h1685: dout <= 8'b00000000; // 5765 :   0 - 0x0
      13'h1686: dout <= 8'b00000000; // 5766 :   0 - 0x0
      13'h1687: dout <= 8'b00000000; // 5767 :   0 - 0x0
      13'h1688: dout <= 8'b00000000; // 5768 :   0 - 0x0
      13'h1689: dout <= 8'b00000000; // 5769 :   0 - 0x0
      13'h168A: dout <= 8'b00000000; // 5770 :   0 - 0x0
      13'h168B: dout <= 8'b00000000; // 5771 :   0 - 0x0
      13'h168C: dout <= 8'b00000000; // 5772 :   0 - 0x0
      13'h168D: dout <= 8'b00000000; // 5773 :   0 - 0x0
      13'h168E: dout <= 8'b00000000; // 5774 :   0 - 0x0
      13'h168F: dout <= 8'b00000000; // 5775 :   0 - 0x0
      13'h1690: dout <= 8'b00000000; // 5776 :   0 - 0x0 -- Background 0x69
      13'h1691: dout <= 8'b00000000; // 5777 :   0 - 0x0
      13'h1692: dout <= 8'b00000000; // 5778 :   0 - 0x0
      13'h1693: dout <= 8'b00000000; // 5779 :   0 - 0x0
      13'h1694: dout <= 8'b00000000; // 5780 :   0 - 0x0
      13'h1695: dout <= 8'b00000000; // 5781 :   0 - 0x0
      13'h1696: dout <= 8'b00000000; // 5782 :   0 - 0x0
      13'h1697: dout <= 8'b00000000; // 5783 :   0 - 0x0
      13'h1698: dout <= 8'b00000000; // 5784 :   0 - 0x0
      13'h1699: dout <= 8'b00000000; // 5785 :   0 - 0x0
      13'h169A: dout <= 8'b00000000; // 5786 :   0 - 0x0
      13'h169B: dout <= 8'b00000000; // 5787 :   0 - 0x0
      13'h169C: dout <= 8'b00000000; // 5788 :   0 - 0x0
      13'h169D: dout <= 8'b00000000; // 5789 :   0 - 0x0
      13'h169E: dout <= 8'b00000000; // 5790 :   0 - 0x0
      13'h169F: dout <= 8'b00000000; // 5791 :   0 - 0x0
      13'h16A0: dout <= 8'b00000000; // 5792 :   0 - 0x0 -- Background 0x6a
      13'h16A1: dout <= 8'b00000000; // 5793 :   0 - 0x0
      13'h16A2: dout <= 8'b00000000; // 5794 :   0 - 0x0
      13'h16A3: dout <= 8'b00000000; // 5795 :   0 - 0x0
      13'h16A4: dout <= 8'b00000000; // 5796 :   0 - 0x0
      13'h16A5: dout <= 8'b00000000; // 5797 :   0 - 0x0
      13'h16A6: dout <= 8'b00000000; // 5798 :   0 - 0x0
      13'h16A7: dout <= 8'b00000000; // 5799 :   0 - 0x0
      13'h16A8: dout <= 8'b00000000; // 5800 :   0 - 0x0
      13'h16A9: dout <= 8'b00000000; // 5801 :   0 - 0x0
      13'h16AA: dout <= 8'b00000000; // 5802 :   0 - 0x0
      13'h16AB: dout <= 8'b00000000; // 5803 :   0 - 0x0
      13'h16AC: dout <= 8'b00000000; // 5804 :   0 - 0x0
      13'h16AD: dout <= 8'b00000000; // 5805 :   0 - 0x0
      13'h16AE: dout <= 8'b00000000; // 5806 :   0 - 0x0
      13'h16AF: dout <= 8'b00000000; // 5807 :   0 - 0x0
      13'h16B0: dout <= 8'b00000000; // 5808 :   0 - 0x0 -- Background 0x6b
      13'h16B1: dout <= 8'b00000000; // 5809 :   0 - 0x0
      13'h16B2: dout <= 8'b00000000; // 5810 :   0 - 0x0
      13'h16B3: dout <= 8'b00000000; // 5811 :   0 - 0x0
      13'h16B4: dout <= 8'b00000000; // 5812 :   0 - 0x0
      13'h16B5: dout <= 8'b00000000; // 5813 :   0 - 0x0
      13'h16B6: dout <= 8'b00000000; // 5814 :   0 - 0x0
      13'h16B7: dout <= 8'b00000000; // 5815 :   0 - 0x0
      13'h16B8: dout <= 8'b00000000; // 5816 :   0 - 0x0
      13'h16B9: dout <= 8'b00000000; // 5817 :   0 - 0x0
      13'h16BA: dout <= 8'b00000000; // 5818 :   0 - 0x0
      13'h16BB: dout <= 8'b00000000; // 5819 :   0 - 0x0
      13'h16BC: dout <= 8'b00000000; // 5820 :   0 - 0x0
      13'h16BD: dout <= 8'b00000000; // 5821 :   0 - 0x0
      13'h16BE: dout <= 8'b00000000; // 5822 :   0 - 0x0
      13'h16BF: dout <= 8'b00000000; // 5823 :   0 - 0x0
      13'h16C0: dout <= 8'b00000000; // 5824 :   0 - 0x0 -- Background 0x6c
      13'h16C1: dout <= 8'b00000000; // 5825 :   0 - 0x0
      13'h16C2: dout <= 8'b00000000; // 5826 :   0 - 0x0
      13'h16C3: dout <= 8'b00000000; // 5827 :   0 - 0x0
      13'h16C4: dout <= 8'b00000000; // 5828 :   0 - 0x0
      13'h16C5: dout <= 8'b00000000; // 5829 :   0 - 0x0
      13'h16C6: dout <= 8'b00000000; // 5830 :   0 - 0x0
      13'h16C7: dout <= 8'b00000000; // 5831 :   0 - 0x0
      13'h16C8: dout <= 8'b00000000; // 5832 :   0 - 0x0
      13'h16C9: dout <= 8'b00000000; // 5833 :   0 - 0x0
      13'h16CA: dout <= 8'b00000000; // 5834 :   0 - 0x0
      13'h16CB: dout <= 8'b00000000; // 5835 :   0 - 0x0
      13'h16CC: dout <= 8'b00000000; // 5836 :   0 - 0x0
      13'h16CD: dout <= 8'b00000000; // 5837 :   0 - 0x0
      13'h16CE: dout <= 8'b00000000; // 5838 :   0 - 0x0
      13'h16CF: dout <= 8'b00000000; // 5839 :   0 - 0x0
      13'h16D0: dout <= 8'b00000000; // 5840 :   0 - 0x0 -- Background 0x6d
      13'h16D1: dout <= 8'b00000000; // 5841 :   0 - 0x0
      13'h16D2: dout <= 8'b00000000; // 5842 :   0 - 0x0
      13'h16D3: dout <= 8'b00000000; // 5843 :   0 - 0x0
      13'h16D4: dout <= 8'b00000000; // 5844 :   0 - 0x0
      13'h16D5: dout <= 8'b00000000; // 5845 :   0 - 0x0
      13'h16D6: dout <= 8'b00000000; // 5846 :   0 - 0x0
      13'h16D7: dout <= 8'b00000000; // 5847 :   0 - 0x0
      13'h16D8: dout <= 8'b00000000; // 5848 :   0 - 0x0
      13'h16D9: dout <= 8'b00000000; // 5849 :   0 - 0x0
      13'h16DA: dout <= 8'b00000000; // 5850 :   0 - 0x0
      13'h16DB: dout <= 8'b00000000; // 5851 :   0 - 0x0
      13'h16DC: dout <= 8'b00000000; // 5852 :   0 - 0x0
      13'h16DD: dout <= 8'b00000000; // 5853 :   0 - 0x0
      13'h16DE: dout <= 8'b00000000; // 5854 :   0 - 0x0
      13'h16DF: dout <= 8'b00000000; // 5855 :   0 - 0x0
      13'h16E0: dout <= 8'b00000000; // 5856 :   0 - 0x0 -- Background 0x6e
      13'h16E1: dout <= 8'b00000000; // 5857 :   0 - 0x0
      13'h16E2: dout <= 8'b00000000; // 5858 :   0 - 0x0
      13'h16E3: dout <= 8'b00000000; // 5859 :   0 - 0x0
      13'h16E4: dout <= 8'b00000000; // 5860 :   0 - 0x0
      13'h16E5: dout <= 8'b00000000; // 5861 :   0 - 0x0
      13'h16E6: dout <= 8'b00000000; // 5862 :   0 - 0x0
      13'h16E7: dout <= 8'b00000000; // 5863 :   0 - 0x0
      13'h16E8: dout <= 8'b00000000; // 5864 :   0 - 0x0
      13'h16E9: dout <= 8'b00000000; // 5865 :   0 - 0x0
      13'h16EA: dout <= 8'b00000000; // 5866 :   0 - 0x0
      13'h16EB: dout <= 8'b00000000; // 5867 :   0 - 0x0
      13'h16EC: dout <= 8'b00000000; // 5868 :   0 - 0x0
      13'h16ED: dout <= 8'b00000000; // 5869 :   0 - 0x0
      13'h16EE: dout <= 8'b00000000; // 5870 :   0 - 0x0
      13'h16EF: dout <= 8'b00000000; // 5871 :   0 - 0x0
      13'h16F0: dout <= 8'b00000000; // 5872 :   0 - 0x0 -- Background 0x6f
      13'h16F1: dout <= 8'b00000000; // 5873 :   0 - 0x0
      13'h16F2: dout <= 8'b00000000; // 5874 :   0 - 0x0
      13'h16F3: dout <= 8'b00000000; // 5875 :   0 - 0x0
      13'h16F4: dout <= 8'b00000000; // 5876 :   0 - 0x0
      13'h16F5: dout <= 8'b00000000; // 5877 :   0 - 0x0
      13'h16F6: dout <= 8'b00000000; // 5878 :   0 - 0x0
      13'h16F7: dout <= 8'b00000000; // 5879 :   0 - 0x0
      13'h16F8: dout <= 8'b00000000; // 5880 :   0 - 0x0
      13'h16F9: dout <= 8'b00000000; // 5881 :   0 - 0x0
      13'h16FA: dout <= 8'b00000000; // 5882 :   0 - 0x0
      13'h16FB: dout <= 8'b00000000; // 5883 :   0 - 0x0
      13'h16FC: dout <= 8'b00000000; // 5884 :   0 - 0x0
      13'h16FD: dout <= 8'b00000000; // 5885 :   0 - 0x0
      13'h16FE: dout <= 8'b00000000; // 5886 :   0 - 0x0
      13'h16FF: dout <= 8'b00000000; // 5887 :   0 - 0x0
      13'h1700: dout <= 8'b00000000; // 5888 :   0 - 0x0 -- Background 0x70
      13'h1701: dout <= 8'b00000000; // 5889 :   0 - 0x0
      13'h1702: dout <= 8'b00000000; // 5890 :   0 - 0x0
      13'h1703: dout <= 8'b00000000; // 5891 :   0 - 0x0
      13'h1704: dout <= 8'b00000000; // 5892 :   0 - 0x0
      13'h1705: dout <= 8'b00000000; // 5893 :   0 - 0x0
      13'h1706: dout <= 8'b00000000; // 5894 :   0 - 0x0
      13'h1707: dout <= 8'b00000000; // 5895 :   0 - 0x0
      13'h1708: dout <= 8'b00000000; // 5896 :   0 - 0x0
      13'h1709: dout <= 8'b00000000; // 5897 :   0 - 0x0
      13'h170A: dout <= 8'b00000000; // 5898 :   0 - 0x0
      13'h170B: dout <= 8'b00000000; // 5899 :   0 - 0x0
      13'h170C: dout <= 8'b00000000; // 5900 :   0 - 0x0
      13'h170D: dout <= 8'b00000000; // 5901 :   0 - 0x0
      13'h170E: dout <= 8'b00000000; // 5902 :   0 - 0x0
      13'h170F: dout <= 8'b00000000; // 5903 :   0 - 0x0
      13'h1710: dout <= 8'b00000000; // 5904 :   0 - 0x0 -- Background 0x71
      13'h1711: dout <= 8'b00000000; // 5905 :   0 - 0x0
      13'h1712: dout <= 8'b00000000; // 5906 :   0 - 0x0
      13'h1713: dout <= 8'b00000000; // 5907 :   0 - 0x0
      13'h1714: dout <= 8'b00000000; // 5908 :   0 - 0x0
      13'h1715: dout <= 8'b00000000; // 5909 :   0 - 0x0
      13'h1716: dout <= 8'b00000000; // 5910 :   0 - 0x0
      13'h1717: dout <= 8'b00000000; // 5911 :   0 - 0x0
      13'h1718: dout <= 8'b00000000; // 5912 :   0 - 0x0
      13'h1719: dout <= 8'b00000000; // 5913 :   0 - 0x0
      13'h171A: dout <= 8'b00000000; // 5914 :   0 - 0x0
      13'h171B: dout <= 8'b00000000; // 5915 :   0 - 0x0
      13'h171C: dout <= 8'b00000000; // 5916 :   0 - 0x0
      13'h171D: dout <= 8'b00000000; // 5917 :   0 - 0x0
      13'h171E: dout <= 8'b00000000; // 5918 :   0 - 0x0
      13'h171F: dout <= 8'b00000000; // 5919 :   0 - 0x0
      13'h1720: dout <= 8'b00000000; // 5920 :   0 - 0x0 -- Background 0x72
      13'h1721: dout <= 8'b00000000; // 5921 :   0 - 0x0
      13'h1722: dout <= 8'b00000000; // 5922 :   0 - 0x0
      13'h1723: dout <= 8'b00000000; // 5923 :   0 - 0x0
      13'h1724: dout <= 8'b00000000; // 5924 :   0 - 0x0
      13'h1725: dout <= 8'b00000000; // 5925 :   0 - 0x0
      13'h1726: dout <= 8'b00000000; // 5926 :   0 - 0x0
      13'h1727: dout <= 8'b00000000; // 5927 :   0 - 0x0
      13'h1728: dout <= 8'b00000000; // 5928 :   0 - 0x0
      13'h1729: dout <= 8'b00000000; // 5929 :   0 - 0x0
      13'h172A: dout <= 8'b00000000; // 5930 :   0 - 0x0
      13'h172B: dout <= 8'b00000000; // 5931 :   0 - 0x0
      13'h172C: dout <= 8'b00000000; // 5932 :   0 - 0x0
      13'h172D: dout <= 8'b00000000; // 5933 :   0 - 0x0
      13'h172E: dout <= 8'b00000000; // 5934 :   0 - 0x0
      13'h172F: dout <= 8'b00000000; // 5935 :   0 - 0x0
      13'h1730: dout <= 8'b00000000; // 5936 :   0 - 0x0 -- Background 0x73
      13'h1731: dout <= 8'b00000000; // 5937 :   0 - 0x0
      13'h1732: dout <= 8'b00000000; // 5938 :   0 - 0x0
      13'h1733: dout <= 8'b00000000; // 5939 :   0 - 0x0
      13'h1734: dout <= 8'b00000000; // 5940 :   0 - 0x0
      13'h1735: dout <= 8'b00000000; // 5941 :   0 - 0x0
      13'h1736: dout <= 8'b00000000; // 5942 :   0 - 0x0
      13'h1737: dout <= 8'b00000000; // 5943 :   0 - 0x0
      13'h1738: dout <= 8'b00000000; // 5944 :   0 - 0x0
      13'h1739: dout <= 8'b00000000; // 5945 :   0 - 0x0
      13'h173A: dout <= 8'b00000000; // 5946 :   0 - 0x0
      13'h173B: dout <= 8'b00000000; // 5947 :   0 - 0x0
      13'h173C: dout <= 8'b00000000; // 5948 :   0 - 0x0
      13'h173D: dout <= 8'b00000000; // 5949 :   0 - 0x0
      13'h173E: dout <= 8'b00000000; // 5950 :   0 - 0x0
      13'h173F: dout <= 8'b00000000; // 5951 :   0 - 0x0
      13'h1740: dout <= 8'b00000000; // 5952 :   0 - 0x0 -- Background 0x74
      13'h1741: dout <= 8'b00000000; // 5953 :   0 - 0x0
      13'h1742: dout <= 8'b00000000; // 5954 :   0 - 0x0
      13'h1743: dout <= 8'b00000000; // 5955 :   0 - 0x0
      13'h1744: dout <= 8'b00000000; // 5956 :   0 - 0x0
      13'h1745: dout <= 8'b00000000; // 5957 :   0 - 0x0
      13'h1746: dout <= 8'b00000000; // 5958 :   0 - 0x0
      13'h1747: dout <= 8'b00000000; // 5959 :   0 - 0x0
      13'h1748: dout <= 8'b00000000; // 5960 :   0 - 0x0
      13'h1749: dout <= 8'b00000000; // 5961 :   0 - 0x0
      13'h174A: dout <= 8'b00000000; // 5962 :   0 - 0x0
      13'h174B: dout <= 8'b00000000; // 5963 :   0 - 0x0
      13'h174C: dout <= 8'b00000000; // 5964 :   0 - 0x0
      13'h174D: dout <= 8'b00000000; // 5965 :   0 - 0x0
      13'h174E: dout <= 8'b00000000; // 5966 :   0 - 0x0
      13'h174F: dout <= 8'b00000000; // 5967 :   0 - 0x0
      13'h1750: dout <= 8'b00000000; // 5968 :   0 - 0x0 -- Background 0x75
      13'h1751: dout <= 8'b00000000; // 5969 :   0 - 0x0
      13'h1752: dout <= 8'b00000000; // 5970 :   0 - 0x0
      13'h1753: dout <= 8'b00000000; // 5971 :   0 - 0x0
      13'h1754: dout <= 8'b00000000; // 5972 :   0 - 0x0
      13'h1755: dout <= 8'b00000000; // 5973 :   0 - 0x0
      13'h1756: dout <= 8'b00000000; // 5974 :   0 - 0x0
      13'h1757: dout <= 8'b00000000; // 5975 :   0 - 0x0
      13'h1758: dout <= 8'b00000000; // 5976 :   0 - 0x0
      13'h1759: dout <= 8'b00000000; // 5977 :   0 - 0x0
      13'h175A: dout <= 8'b00000000; // 5978 :   0 - 0x0
      13'h175B: dout <= 8'b00000000; // 5979 :   0 - 0x0
      13'h175C: dout <= 8'b00000000; // 5980 :   0 - 0x0
      13'h175D: dout <= 8'b00000000; // 5981 :   0 - 0x0
      13'h175E: dout <= 8'b00000000; // 5982 :   0 - 0x0
      13'h175F: dout <= 8'b00000000; // 5983 :   0 - 0x0
      13'h1760: dout <= 8'b00000000; // 5984 :   0 - 0x0 -- Background 0x76
      13'h1761: dout <= 8'b00000000; // 5985 :   0 - 0x0
      13'h1762: dout <= 8'b00000000; // 5986 :   0 - 0x0
      13'h1763: dout <= 8'b00000000; // 5987 :   0 - 0x0
      13'h1764: dout <= 8'b00000000; // 5988 :   0 - 0x0
      13'h1765: dout <= 8'b00000000; // 5989 :   0 - 0x0
      13'h1766: dout <= 8'b00000000; // 5990 :   0 - 0x0
      13'h1767: dout <= 8'b00000000; // 5991 :   0 - 0x0
      13'h1768: dout <= 8'b00000000; // 5992 :   0 - 0x0
      13'h1769: dout <= 8'b00000000; // 5993 :   0 - 0x0
      13'h176A: dout <= 8'b00000000; // 5994 :   0 - 0x0
      13'h176B: dout <= 8'b00000000; // 5995 :   0 - 0x0
      13'h176C: dout <= 8'b00000000; // 5996 :   0 - 0x0
      13'h176D: dout <= 8'b00000000; // 5997 :   0 - 0x0
      13'h176E: dout <= 8'b00000000; // 5998 :   0 - 0x0
      13'h176F: dout <= 8'b00000000; // 5999 :   0 - 0x0
      13'h1770: dout <= 8'b00000000; // 6000 :   0 - 0x0 -- Background 0x77
      13'h1771: dout <= 8'b00000000; // 6001 :   0 - 0x0
      13'h1772: dout <= 8'b00000000; // 6002 :   0 - 0x0
      13'h1773: dout <= 8'b00000000; // 6003 :   0 - 0x0
      13'h1774: dout <= 8'b00000000; // 6004 :   0 - 0x0
      13'h1775: dout <= 8'b00000000; // 6005 :   0 - 0x0
      13'h1776: dout <= 8'b00000000; // 6006 :   0 - 0x0
      13'h1777: dout <= 8'b00000000; // 6007 :   0 - 0x0
      13'h1778: dout <= 8'b00000000; // 6008 :   0 - 0x0
      13'h1779: dout <= 8'b00000000; // 6009 :   0 - 0x0
      13'h177A: dout <= 8'b00000000; // 6010 :   0 - 0x0
      13'h177B: dout <= 8'b00000000; // 6011 :   0 - 0x0
      13'h177C: dout <= 8'b00000000; // 6012 :   0 - 0x0
      13'h177D: dout <= 8'b00000000; // 6013 :   0 - 0x0
      13'h177E: dout <= 8'b00000000; // 6014 :   0 - 0x0
      13'h177F: dout <= 8'b00000000; // 6015 :   0 - 0x0
      13'h1780: dout <= 8'b00000000; // 6016 :   0 - 0x0 -- Background 0x78
      13'h1781: dout <= 8'b00000000; // 6017 :   0 - 0x0
      13'h1782: dout <= 8'b00000000; // 6018 :   0 - 0x0
      13'h1783: dout <= 8'b00000000; // 6019 :   0 - 0x0
      13'h1784: dout <= 8'b00000000; // 6020 :   0 - 0x0
      13'h1785: dout <= 8'b00000000; // 6021 :   0 - 0x0
      13'h1786: dout <= 8'b00000000; // 6022 :   0 - 0x0
      13'h1787: dout <= 8'b00000000; // 6023 :   0 - 0x0
      13'h1788: dout <= 8'b00000000; // 6024 :   0 - 0x0
      13'h1789: dout <= 8'b00000000; // 6025 :   0 - 0x0
      13'h178A: dout <= 8'b00000000; // 6026 :   0 - 0x0
      13'h178B: dout <= 8'b00000000; // 6027 :   0 - 0x0
      13'h178C: dout <= 8'b00000000; // 6028 :   0 - 0x0
      13'h178D: dout <= 8'b00000000; // 6029 :   0 - 0x0
      13'h178E: dout <= 8'b00000000; // 6030 :   0 - 0x0
      13'h178F: dout <= 8'b00000000; // 6031 :   0 - 0x0
      13'h1790: dout <= 8'b00000000; // 6032 :   0 - 0x0 -- Background 0x79
      13'h1791: dout <= 8'b00000000; // 6033 :   0 - 0x0
      13'h1792: dout <= 8'b00000000; // 6034 :   0 - 0x0
      13'h1793: dout <= 8'b00000000; // 6035 :   0 - 0x0
      13'h1794: dout <= 8'b00000000; // 6036 :   0 - 0x0
      13'h1795: dout <= 8'b00000000; // 6037 :   0 - 0x0
      13'h1796: dout <= 8'b00000000; // 6038 :   0 - 0x0
      13'h1797: dout <= 8'b00000000; // 6039 :   0 - 0x0
      13'h1798: dout <= 8'b00000000; // 6040 :   0 - 0x0
      13'h1799: dout <= 8'b00000000; // 6041 :   0 - 0x0
      13'h179A: dout <= 8'b00000000; // 6042 :   0 - 0x0
      13'h179B: dout <= 8'b00000000; // 6043 :   0 - 0x0
      13'h179C: dout <= 8'b00000000; // 6044 :   0 - 0x0
      13'h179D: dout <= 8'b00000000; // 6045 :   0 - 0x0
      13'h179E: dout <= 8'b00000000; // 6046 :   0 - 0x0
      13'h179F: dout <= 8'b00000000; // 6047 :   0 - 0x0
      13'h17A0: dout <= 8'b00000000; // 6048 :   0 - 0x0 -- Background 0x7a
      13'h17A1: dout <= 8'b00000000; // 6049 :   0 - 0x0
      13'h17A2: dout <= 8'b00000000; // 6050 :   0 - 0x0
      13'h17A3: dout <= 8'b00000000; // 6051 :   0 - 0x0
      13'h17A4: dout <= 8'b00000000; // 6052 :   0 - 0x0
      13'h17A5: dout <= 8'b00000000; // 6053 :   0 - 0x0
      13'h17A6: dout <= 8'b00000000; // 6054 :   0 - 0x0
      13'h17A7: dout <= 8'b00000000; // 6055 :   0 - 0x0
      13'h17A8: dout <= 8'b00000000; // 6056 :   0 - 0x0
      13'h17A9: dout <= 8'b00000000; // 6057 :   0 - 0x0
      13'h17AA: dout <= 8'b00000000; // 6058 :   0 - 0x0
      13'h17AB: dout <= 8'b00000000; // 6059 :   0 - 0x0
      13'h17AC: dout <= 8'b00000000; // 6060 :   0 - 0x0
      13'h17AD: dout <= 8'b00000000; // 6061 :   0 - 0x0
      13'h17AE: dout <= 8'b00000000; // 6062 :   0 - 0x0
      13'h17AF: dout <= 8'b00000000; // 6063 :   0 - 0x0
      13'h17B0: dout <= 8'b00000000; // 6064 :   0 - 0x0 -- Background 0x7b
      13'h17B1: dout <= 8'b00000000; // 6065 :   0 - 0x0
      13'h17B2: dout <= 8'b00000000; // 6066 :   0 - 0x0
      13'h17B3: dout <= 8'b00000000; // 6067 :   0 - 0x0
      13'h17B4: dout <= 8'b00000000; // 6068 :   0 - 0x0
      13'h17B5: dout <= 8'b00000000; // 6069 :   0 - 0x0
      13'h17B6: dout <= 8'b00000000; // 6070 :   0 - 0x0
      13'h17B7: dout <= 8'b00000000; // 6071 :   0 - 0x0
      13'h17B8: dout <= 8'b00000000; // 6072 :   0 - 0x0
      13'h17B9: dout <= 8'b00000000; // 6073 :   0 - 0x0
      13'h17BA: dout <= 8'b00000000; // 6074 :   0 - 0x0
      13'h17BB: dout <= 8'b00000000; // 6075 :   0 - 0x0
      13'h17BC: dout <= 8'b00000000; // 6076 :   0 - 0x0
      13'h17BD: dout <= 8'b00000000; // 6077 :   0 - 0x0
      13'h17BE: dout <= 8'b00000000; // 6078 :   0 - 0x0
      13'h17BF: dout <= 8'b00000000; // 6079 :   0 - 0x0
      13'h17C0: dout <= 8'b00000000; // 6080 :   0 - 0x0 -- Background 0x7c
      13'h17C1: dout <= 8'b00000000; // 6081 :   0 - 0x0
      13'h17C2: dout <= 8'b00000000; // 6082 :   0 - 0x0
      13'h17C3: dout <= 8'b00000000; // 6083 :   0 - 0x0
      13'h17C4: dout <= 8'b00000000; // 6084 :   0 - 0x0
      13'h17C5: dout <= 8'b00000000; // 6085 :   0 - 0x0
      13'h17C6: dout <= 8'b00000000; // 6086 :   0 - 0x0
      13'h17C7: dout <= 8'b00000000; // 6087 :   0 - 0x0
      13'h17C8: dout <= 8'b00000000; // 6088 :   0 - 0x0
      13'h17C9: dout <= 8'b00000000; // 6089 :   0 - 0x0
      13'h17CA: dout <= 8'b00000000; // 6090 :   0 - 0x0
      13'h17CB: dout <= 8'b00000000; // 6091 :   0 - 0x0
      13'h17CC: dout <= 8'b00000000; // 6092 :   0 - 0x0
      13'h17CD: dout <= 8'b00000000; // 6093 :   0 - 0x0
      13'h17CE: dout <= 8'b00000000; // 6094 :   0 - 0x0
      13'h17CF: dout <= 8'b00000000; // 6095 :   0 - 0x0
      13'h17D0: dout <= 8'b00000000; // 6096 :   0 - 0x0 -- Background 0x7d
      13'h17D1: dout <= 8'b00000000; // 6097 :   0 - 0x0
      13'h17D2: dout <= 8'b00000000; // 6098 :   0 - 0x0
      13'h17D3: dout <= 8'b00000000; // 6099 :   0 - 0x0
      13'h17D4: dout <= 8'b00000000; // 6100 :   0 - 0x0
      13'h17D5: dout <= 8'b00000000; // 6101 :   0 - 0x0
      13'h17D6: dout <= 8'b00000000; // 6102 :   0 - 0x0
      13'h17D7: dout <= 8'b00000000; // 6103 :   0 - 0x0
      13'h17D8: dout <= 8'b00000000; // 6104 :   0 - 0x0
      13'h17D9: dout <= 8'b00000000; // 6105 :   0 - 0x0
      13'h17DA: dout <= 8'b00000000; // 6106 :   0 - 0x0
      13'h17DB: dout <= 8'b00000000; // 6107 :   0 - 0x0
      13'h17DC: dout <= 8'b00000000; // 6108 :   0 - 0x0
      13'h17DD: dout <= 8'b00000000; // 6109 :   0 - 0x0
      13'h17DE: dout <= 8'b00000000; // 6110 :   0 - 0x0
      13'h17DF: dout <= 8'b00000000; // 6111 :   0 - 0x0
      13'h17E0: dout <= 8'b00000000; // 6112 :   0 - 0x0 -- Background 0x7e
      13'h17E1: dout <= 8'b00000000; // 6113 :   0 - 0x0
      13'h17E2: dout <= 8'b00000000; // 6114 :   0 - 0x0
      13'h17E3: dout <= 8'b00000000; // 6115 :   0 - 0x0
      13'h17E4: dout <= 8'b00000000; // 6116 :   0 - 0x0
      13'h17E5: dout <= 8'b00000000; // 6117 :   0 - 0x0
      13'h17E6: dout <= 8'b00000000; // 6118 :   0 - 0x0
      13'h17E7: dout <= 8'b00000000; // 6119 :   0 - 0x0
      13'h17E8: dout <= 8'b00000000; // 6120 :   0 - 0x0
      13'h17E9: dout <= 8'b00000000; // 6121 :   0 - 0x0
      13'h17EA: dout <= 8'b00000000; // 6122 :   0 - 0x0
      13'h17EB: dout <= 8'b00000000; // 6123 :   0 - 0x0
      13'h17EC: dout <= 8'b00000000; // 6124 :   0 - 0x0
      13'h17ED: dout <= 8'b00000000; // 6125 :   0 - 0x0
      13'h17EE: dout <= 8'b00000000; // 6126 :   0 - 0x0
      13'h17EF: dout <= 8'b00000000; // 6127 :   0 - 0x0
      13'h17F0: dout <= 8'b00000000; // 6128 :   0 - 0x0 -- Background 0x7f
      13'h17F1: dout <= 8'b00000000; // 6129 :   0 - 0x0
      13'h17F2: dout <= 8'b00000000; // 6130 :   0 - 0x0
      13'h17F3: dout <= 8'b00000000; // 6131 :   0 - 0x0
      13'h17F4: dout <= 8'b00000000; // 6132 :   0 - 0x0
      13'h17F5: dout <= 8'b00000000; // 6133 :   0 - 0x0
      13'h17F6: dout <= 8'b00000000; // 6134 :   0 - 0x0
      13'h17F7: dout <= 8'b00000000; // 6135 :   0 - 0x0
      13'h17F8: dout <= 8'b00000000; // 6136 :   0 - 0x0
      13'h17F9: dout <= 8'b00000000; // 6137 :   0 - 0x0
      13'h17FA: dout <= 8'b00000000; // 6138 :   0 - 0x0
      13'h17FB: dout <= 8'b00000000; // 6139 :   0 - 0x0
      13'h17FC: dout <= 8'b00000000; // 6140 :   0 - 0x0
      13'h17FD: dout <= 8'b00000000; // 6141 :   0 - 0x0
      13'h17FE: dout <= 8'b00000000; // 6142 :   0 - 0x0
      13'h17FF: dout <= 8'b00000000; // 6143 :   0 - 0x0
      13'h1800: dout <= 8'b10111111; // 6144 : 191 - 0xbf -- Background 0x80
      13'h1801: dout <= 8'b11110111; // 6145 : 247 - 0xf7
      13'h1802: dout <= 8'b11111101; // 6146 : 253 - 0xfd
      13'h1803: dout <= 8'b11011111; // 6147 : 223 - 0xdf
      13'h1804: dout <= 8'b11111011; // 6148 : 251 - 0xfb
      13'h1805: dout <= 8'b10111111; // 6149 : 191 - 0xbf
      13'h1806: dout <= 8'b11111110; // 6150 : 254 - 0xfe
      13'h1807: dout <= 8'b11101111; // 6151 : 239 - 0xef
      13'h1808: dout <= 8'b01000000; // 6152 :  64 - 0x40
      13'h1809: dout <= 8'b00001000; // 6153 :   8 - 0x8
      13'h180A: dout <= 8'b00000010; // 6154 :   2 - 0x2
      13'h180B: dout <= 8'b00100000; // 6155 :  32 - 0x20
      13'h180C: dout <= 8'b00000100; // 6156 :   4 - 0x4
      13'h180D: dout <= 8'b01000000; // 6157 :  64 - 0x40
      13'h180E: dout <= 8'b00000001; // 6158 :   1 - 0x1
      13'h180F: dout <= 8'b00010000; // 6159 :  16 - 0x10
      13'h1810: dout <= 8'b11111111; // 6160 : 255 - 0xff -- Background 0x81
      13'h1811: dout <= 8'b11101110; // 6161 : 238 - 0xee
      13'h1812: dout <= 8'b11111111; // 6162 : 255 - 0xff
      13'h1813: dout <= 8'b11011111; // 6163 : 223 - 0xdf
      13'h1814: dout <= 8'b01110111; // 6164 : 119 - 0x77
      13'h1815: dout <= 8'b11111101; // 6165 : 253 - 0xfd
      13'h1816: dout <= 8'b11011111; // 6166 : 223 - 0xdf
      13'h1817: dout <= 8'b10111111; // 6167 : 191 - 0xbf
      13'h1818: dout <= 8'b00000000; // 6168 :   0 - 0x0
      13'h1819: dout <= 8'b00010001; // 6169 :  17 - 0x11
      13'h181A: dout <= 8'b00000000; // 6170 :   0 - 0x0
      13'h181B: dout <= 8'b00100000; // 6171 :  32 - 0x20
      13'h181C: dout <= 8'b10001000; // 6172 : 136 - 0x88
      13'h181D: dout <= 8'b00000010; // 6173 :   2 - 0x2
      13'h181E: dout <= 8'b00100000; // 6174 :  32 - 0x20
      13'h181F: dout <= 8'b01000000; // 6175 :  64 - 0x40
      13'h1820: dout <= 8'b11111110; // 6176 : 254 - 0xfe -- Background 0x82
      13'h1821: dout <= 8'b11101111; // 6177 : 239 - 0xef
      13'h1822: dout <= 8'b10111111; // 6178 : 191 - 0xbf
      13'h1823: dout <= 8'b11110111; // 6179 : 247 - 0xf7
      13'h1824: dout <= 8'b11111101; // 6180 : 253 - 0xfd
      13'h1825: dout <= 8'b11011111; // 6181 : 223 - 0xdf
      13'h1826: dout <= 8'b11111011; // 6182 : 251 - 0xfb
      13'h1827: dout <= 8'b10111111; // 6183 : 191 - 0xbf
      13'h1828: dout <= 8'b00000001; // 6184 :   1 - 0x1
      13'h1829: dout <= 8'b00010000; // 6185 :  16 - 0x10
      13'h182A: dout <= 8'b01000000; // 6186 :  64 - 0x40
      13'h182B: dout <= 8'b00001000; // 6187 :   8 - 0x8
      13'h182C: dout <= 8'b00000010; // 6188 :   2 - 0x2
      13'h182D: dout <= 8'b00100000; // 6189 :  32 - 0x20
      13'h182E: dout <= 8'b00000100; // 6190 :   4 - 0x4
      13'h182F: dout <= 8'b01000000; // 6191 :  64 - 0x40
      13'h1830: dout <= 8'b11101111; // 6192 : 239 - 0xef -- Background 0x83
      13'h1831: dout <= 8'b11111111; // 6193 : 255 - 0xff
      13'h1832: dout <= 8'b10111011; // 6194 : 187 - 0xbb
      13'h1833: dout <= 8'b11111111; // 6195 : 255 - 0xff
      13'h1834: dout <= 8'b11110111; // 6196 : 247 - 0xf7
      13'h1835: dout <= 8'b11011101; // 6197 : 221 - 0xdd
      13'h1836: dout <= 8'b01111111; // 6198 : 127 - 0x7f
      13'h1837: dout <= 8'b11110111; // 6199 : 247 - 0xf7
      13'h1838: dout <= 8'b00010000; // 6200 :  16 - 0x10
      13'h1839: dout <= 8'b00000000; // 6201 :   0 - 0x0
      13'h183A: dout <= 8'b01000100; // 6202 :  68 - 0x44
      13'h183B: dout <= 8'b00000000; // 6203 :   0 - 0x0
      13'h183C: dout <= 8'b00001000; // 6204 :   8 - 0x8
      13'h183D: dout <= 8'b00100010; // 6205 :  34 - 0x22
      13'h183E: dout <= 8'b10000000; // 6206 : 128 - 0x80
      13'h183F: dout <= 8'b00001000; // 6207 :   8 - 0x8
      13'h1840: dout <= 8'b11111111; // 6208 : 255 - 0xff -- Background 0x84
      13'h1841: dout <= 8'b11101110; // 6209 : 238 - 0xee
      13'h1842: dout <= 8'b11111011; // 6210 : 251 - 0xfb
      13'h1843: dout <= 8'b10111111; // 6211 : 191 - 0xbf
      13'h1844: dout <= 8'b01111111; // 6212 : 127 - 0x7f
      13'h1845: dout <= 8'b11101101; // 6213 : 237 - 0xed
      13'h1846: dout <= 8'b11111111; // 6214 : 255 - 0xff
      13'h1847: dout <= 8'b10111111; // 6215 : 191 - 0xbf
      13'h1848: dout <= 8'b00010100; // 6216 :  20 - 0x14
      13'h1849: dout <= 8'b10110101; // 6217 : 181 - 0xb5
      13'h184A: dout <= 8'b01000100; // 6218 :  68 - 0x44
      13'h184B: dout <= 8'b01001010; // 6219 :  74 - 0x4a
      13'h184C: dout <= 8'b10010010; // 6220 : 146 - 0x92
      13'h184D: dout <= 8'b10010010; // 6221 : 146 - 0x92
      13'h184E: dout <= 8'b01000100; // 6222 :  68 - 0x44
      13'h184F: dout <= 8'b01001001; // 6223 :  73 - 0x49
      13'h1850: dout <= 8'b11111111; // 6224 : 255 - 0xff -- Background 0x85
      13'h1851: dout <= 8'b10111111; // 6225 : 191 - 0xbf
      13'h1852: dout <= 8'b01111101; // 6226 : 125 - 0x7d
      13'h1853: dout <= 8'b11110111; // 6227 : 247 - 0xf7
      13'h1854: dout <= 8'b11011011; // 6228 : 219 - 0xdb
      13'h1855: dout <= 8'b11111101; // 6229 : 253 - 0xfd
      13'h1856: dout <= 8'b01111110; // 6230 : 126 - 0x7e
      13'h1857: dout <= 8'b11111011; // 6231 : 251 - 0xfb
      13'h1858: dout <= 8'b01000010; // 6232 :  66 - 0x42
      13'h1859: dout <= 8'b01001010; // 6233 :  74 - 0x4a
      13'h185A: dout <= 8'b11001010; // 6234 : 202 - 0xca
      13'h185B: dout <= 8'b00101001; // 6235 :  41 - 0x29
      13'h185C: dout <= 8'b10100110; // 6236 : 166 - 0xa6
      13'h185D: dout <= 8'b10010010; // 6237 : 146 - 0x92
      13'h185E: dout <= 8'b10001001; // 6238 : 137 - 0x89
      13'h185F: dout <= 8'b00101101; // 6239 :  45 - 0x2d
      13'h1860: dout <= 8'b11111111; // 6240 : 255 - 0xff -- Background 0x86
      13'h1861: dout <= 8'b11110111; // 6241 : 247 - 0xf7
      13'h1862: dout <= 8'b11111111; // 6242 : 255 - 0xff
      13'h1863: dout <= 8'b11011101; // 6243 : 221 - 0xdd
      13'h1864: dout <= 8'b01111111; // 6244 : 127 - 0x7f
      13'h1865: dout <= 8'b11110111; // 6245 : 247 - 0xf7
      13'h1866: dout <= 8'b11101111; // 6246 : 239 - 0xef
      13'h1867: dout <= 8'b10111101; // 6247 : 189 - 0xbd
      13'h1868: dout <= 8'b10001000; // 6248 : 136 - 0x88
      13'h1869: dout <= 8'b00101001; // 6249 :  41 - 0x29
      13'h186A: dout <= 8'b10000010; // 6250 : 130 - 0x82
      13'h186B: dout <= 8'b10110110; // 6251 : 182 - 0xb6
      13'h186C: dout <= 8'b10001000; // 6252 : 136 - 0x88
      13'h186D: dout <= 8'b01001001; // 6253 :  73 - 0x49
      13'h186E: dout <= 8'b01010010; // 6254 :  82 - 0x52
      13'h186F: dout <= 8'b01010010; // 6255 :  82 - 0x52
      13'h1870: dout <= 8'b01011111; // 6256 :  95 - 0x5f -- Background 0x87
      13'h1871: dout <= 8'b11111101; // 6257 : 253 - 0xfd
      13'h1872: dout <= 8'b11110110; // 6258 : 246 - 0xf6
      13'h1873: dout <= 8'b01111111; // 6259 : 127 - 0x7f
      13'h1874: dout <= 8'b10011111; // 6260 : 159 - 0x9f
      13'h1875: dout <= 8'b11111110; // 6261 : 254 - 0xfe
      13'h1876: dout <= 8'b11111111; // 6262 : 255 - 0xff
      13'h1877: dout <= 8'b11101111; // 6263 : 239 - 0xef
      13'h1878: dout <= 8'b10110010; // 6264 : 178 - 0xb2
      13'h1879: dout <= 8'b01001010; // 6265 :  74 - 0x4a
      13'h187A: dout <= 8'b10101001; // 6266 : 169 - 0xa9
      13'h187B: dout <= 8'b10100100; // 6267 : 164 - 0xa4
      13'h187C: dout <= 8'b01100010; // 6268 :  98 - 0x62
      13'h187D: dout <= 8'b01001011; // 6269 :  75 - 0x4b
      13'h187E: dout <= 8'b10010000; // 6270 : 144 - 0x90
      13'h187F: dout <= 8'b10010010; // 6271 : 146 - 0x92
      13'h1880: dout <= 8'b11111111; // 6272 : 255 - 0xff -- Background 0x88
      13'h1881: dout <= 8'b10011111; // 6273 : 159 - 0x9f
      13'h1882: dout <= 8'b10111111; // 6274 : 191 - 0xbf
      13'h1883: dout <= 8'b11111111; // 6275 : 255 - 0xff
      13'h1884: dout <= 8'b11110011; // 6276 : 243 - 0xf3
      13'h1885: dout <= 8'b11110011; // 6277 : 243 - 0xf3
      13'h1886: dout <= 8'b11111111; // 6278 : 255 - 0xff
      13'h1887: dout <= 8'b11111111; // 6279 : 255 - 0xff
      13'h1888: dout <= 8'b01100000; // 6280 :  96 - 0x60
      13'h1889: dout <= 8'b11110000; // 6281 : 240 - 0xf0
      13'h188A: dout <= 8'b11110000; // 6282 : 240 - 0xf0
      13'h188B: dout <= 8'b01101110; // 6283 : 110 - 0x6e
      13'h188C: dout <= 8'b00011111; // 6284 :  31 - 0x1f
      13'h188D: dout <= 8'b00011111; // 6285 :  31 - 0x1f
      13'h188E: dout <= 8'b00011111; // 6286 :  31 - 0x1f
      13'h188F: dout <= 8'b00001110; // 6287 :  14 - 0xe
      13'h1890: dout <= 8'b11111111; // 6288 : 255 - 0xff -- Background 0x89
      13'h1891: dout <= 8'b10011111; // 6289 : 159 - 0x9f
      13'h1892: dout <= 8'b10111111; // 6290 : 191 - 0xbf
      13'h1893: dout <= 8'b11110011; // 6291 : 243 - 0xf3
      13'h1894: dout <= 8'b11110011; // 6292 : 243 - 0xf3
      13'h1895: dout <= 8'b11111111; // 6293 : 255 - 0xff
      13'h1896: dout <= 8'b11111111; // 6294 : 255 - 0xff
      13'h1897: dout <= 8'b11111111; // 6295 : 255 - 0xff
      13'h1898: dout <= 8'b01100000; // 6296 :  96 - 0x60
      13'h1899: dout <= 8'b11110000; // 6297 : 240 - 0xf0
      13'h189A: dout <= 8'b11111110; // 6298 : 254 - 0xfe
      13'h189B: dout <= 8'b01111111; // 6299 : 127 - 0x7f
      13'h189C: dout <= 8'b00011111; // 6300 :  31 - 0x1f
      13'h189D: dout <= 8'b00011111; // 6301 :  31 - 0x1f
      13'h189E: dout <= 8'b00001110; // 6302 :  14 - 0xe
      13'h189F: dout <= 8'b00000000; // 6303 :   0 - 0x0
      13'h18A0: dout <= 8'b10111111; // 6304 : 191 - 0xbf -- Background 0x8a
      13'h18A1: dout <= 8'b11110111; // 6305 : 247 - 0xf7
      13'h18A2: dout <= 8'b11111101; // 6306 : 253 - 0xfd
      13'h18A3: dout <= 8'b11111111; // 6307 : 255 - 0xff
      13'h18A4: dout <= 8'b11111011; // 6308 : 251 - 0xfb
      13'h18A5: dout <= 8'b10111111; // 6309 : 191 - 0xbf
      13'h18A6: dout <= 8'b11111110; // 6310 : 254 - 0xfe
      13'h18A7: dout <= 8'b11101111; // 6311 : 239 - 0xef
      13'h18A8: dout <= 8'b01000000; // 6312 :  64 - 0x40
      13'h18A9: dout <= 8'b00001000; // 6313 :   8 - 0x8
      13'h18AA: dout <= 8'b00000010; // 6314 :   2 - 0x2
      13'h18AB: dout <= 8'b00101000; // 6315 :  40 - 0x28
      13'h18AC: dout <= 8'b00010100; // 6316 :  20 - 0x14
      13'h18AD: dout <= 8'b01010100; // 6317 :  84 - 0x54
      13'h18AE: dout <= 8'b00000001; // 6318 :   1 - 0x1
      13'h18AF: dout <= 8'b00010000; // 6319 :  16 - 0x10
      13'h18B0: dout <= 8'b10111111; // 6320 : 191 - 0xbf -- Background 0x8b
      13'h18B1: dout <= 8'b11111111; // 6321 : 255 - 0xff
      13'h18B2: dout <= 8'b11101110; // 6322 : 238 - 0xee
      13'h18B3: dout <= 8'b11111111; // 6323 : 255 - 0xff
      13'h18B4: dout <= 8'b11011111; // 6324 : 223 - 0xdf
      13'h18B5: dout <= 8'b01111101; // 6325 : 125 - 0x7d
      13'h18B6: dout <= 8'b11111111; // 6326 : 255 - 0xff
      13'h18B7: dout <= 8'b11011111; // 6327 : 223 - 0xdf
      13'h18B8: dout <= 8'b01000000; // 6328 :  64 - 0x40
      13'h18B9: dout <= 8'b00000000; // 6329 :   0 - 0x0
      13'h18BA: dout <= 8'b10010001; // 6330 : 145 - 0x91
      13'h18BB: dout <= 8'b00010100; // 6331 :  20 - 0x14
      13'h18BC: dout <= 8'b00101000; // 6332 :  40 - 0x28
      13'h18BD: dout <= 8'b10001010; // 6333 : 138 - 0x8a
      13'h18BE: dout <= 8'b01000000; // 6334 :  64 - 0x40
      13'h18BF: dout <= 8'b00100000; // 6335 :  32 - 0x20
      13'h18C0: dout <= 8'b11111111; // 6336 : 255 - 0xff -- Background 0x8c
      13'h18C1: dout <= 8'b11111000; // 6337 : 248 - 0xf8
      13'h18C2: dout <= 8'b11100010; // 6338 : 226 - 0xe2
      13'h18C3: dout <= 8'b11010111; // 6339 : 215 - 0xd7
      13'h18C4: dout <= 8'b11001111; // 6340 : 207 - 0xcf
      13'h18C5: dout <= 8'b10011111; // 6341 : 159 - 0x9f
      13'h18C6: dout <= 8'b10111110; // 6342 : 190 - 0xbe
      13'h18C7: dout <= 8'b10011101; // 6343 : 157 - 0x9d
      13'h18C8: dout <= 8'b00000000; // 6344 :   0 - 0x0
      13'h18C9: dout <= 8'b00000111; // 6345 :   7 - 0x7
      13'h18CA: dout <= 8'b00011111; // 6346 :  31 - 0x1f
      13'h18CB: dout <= 8'b00111111; // 6347 :  63 - 0x3f
      13'h18CC: dout <= 8'b00111111; // 6348 :  63 - 0x3f
      13'h18CD: dout <= 8'b01111111; // 6349 : 127 - 0x7f
      13'h18CE: dout <= 8'b01111111; // 6350 : 127 - 0x7f
      13'h18CF: dout <= 8'b01111111; // 6351 : 127 - 0x7f
      13'h18D0: dout <= 8'b11111111; // 6352 : 255 - 0xff -- Background 0x8d
      13'h18D1: dout <= 8'b00011111; // 6353 :  31 - 0x1f
      13'h18D2: dout <= 8'b10100111; // 6354 : 167 - 0xa7
      13'h18D3: dout <= 8'b11000011; // 6355 : 195 - 0xc3
      13'h18D4: dout <= 8'b11100011; // 6356 : 227 - 0xe3
      13'h18D5: dout <= 8'b01000001; // 6357 :  65 - 0x41
      13'h18D6: dout <= 8'b10100001; // 6358 : 161 - 0xa1
      13'h18D7: dout <= 8'b00000001; // 6359 :   1 - 0x1
      13'h18D8: dout <= 8'b00000000; // 6360 :   0 - 0x0
      13'h18D9: dout <= 8'b11100000; // 6361 : 224 - 0xe0
      13'h18DA: dout <= 8'b11111000; // 6362 : 248 - 0xf8
      13'h18DB: dout <= 8'b11111000; // 6363 : 248 - 0xf8
      13'h18DC: dout <= 8'b11110000; // 6364 : 240 - 0xf0
      13'h18DD: dout <= 8'b11111000; // 6365 : 248 - 0xf8
      13'h18DE: dout <= 8'b11110100; // 6366 : 244 - 0xf4
      13'h18DF: dout <= 8'b11111000; // 6367 : 248 - 0xf8
      13'h18E0: dout <= 8'b10111110; // 6368 : 190 - 0xbe -- Background 0x8e
      13'h18E1: dout <= 8'b11111111; // 6369 : 255 - 0xff
      13'h18E2: dout <= 8'b11011111; // 6370 : 223 - 0xdf
      13'h18E3: dout <= 8'b11111111; // 6371 : 255 - 0xff
      13'h18E4: dout <= 8'b11101111; // 6372 : 239 - 0xef
      13'h18E5: dout <= 8'b11111111; // 6373 : 255 - 0xff
      13'h18E6: dout <= 8'b11110111; // 6374 : 247 - 0xf7
      13'h18E7: dout <= 8'b11111111; // 6375 : 255 - 0xff
      13'h18E8: dout <= 8'b01111111; // 6376 : 127 - 0x7f
      13'h18E9: dout <= 8'b00111111; // 6377 :  63 - 0x3f
      13'h18EA: dout <= 8'b00111111; // 6378 :  63 - 0x3f
      13'h18EB: dout <= 8'b00011111; // 6379 :  31 - 0x1f
      13'h18EC: dout <= 8'b00011111; // 6380 :  31 - 0x1f
      13'h18ED: dout <= 8'b00001111; // 6381 :  15 - 0xf
      13'h18EE: dout <= 8'b00001111; // 6382 :  15 - 0xf
      13'h18EF: dout <= 8'b00000111; // 6383 :   7 - 0x7
      13'h18F0: dout <= 8'b01111101; // 6384 : 125 - 0x7d -- Background 0x8f
      13'h18F1: dout <= 8'b11111111; // 6385 : 255 - 0xff
      13'h18F2: dout <= 8'b11111011; // 6386 : 251 - 0xfb
      13'h18F3: dout <= 8'b11111111; // 6387 : 255 - 0xff
      13'h18F4: dout <= 8'b11110111; // 6388 : 247 - 0xf7
      13'h18F5: dout <= 8'b11111111; // 6389 : 255 - 0xff
      13'h18F6: dout <= 8'b11101111; // 6390 : 239 - 0xef
      13'h18F7: dout <= 8'b11111111; // 6391 : 255 - 0xff
      13'h18F8: dout <= 8'b11111110; // 6392 : 254 - 0xfe
      13'h18F9: dout <= 8'b11111100; // 6393 : 252 - 0xfc
      13'h18FA: dout <= 8'b11111100; // 6394 : 252 - 0xfc
      13'h18FB: dout <= 8'b11111000; // 6395 : 248 - 0xf8
      13'h18FC: dout <= 8'b11111000; // 6396 : 248 - 0xf8
      13'h18FD: dout <= 8'b11110000; // 6397 : 240 - 0xf0
      13'h18FE: dout <= 8'b11110000; // 6398 : 240 - 0xf0
      13'h18FF: dout <= 8'b11100000; // 6399 : 224 - 0xe0
      13'h1900: dout <= 8'b10111110; // 6400 : 190 - 0xbe -- Background 0x90
      13'h1901: dout <= 8'b11110111; // 6401 : 247 - 0xf7
      13'h1902: dout <= 8'b11111111; // 6402 : 255 - 0xff
      13'h1903: dout <= 8'b11011111; // 6403 : 223 - 0xdf
      13'h1904: dout <= 8'b11111011; // 6404 : 251 - 0xfb
      13'h1905: dout <= 8'b11111110; // 6405 : 254 - 0xfe
      13'h1906: dout <= 8'b10111111; // 6406 : 191 - 0xbf
      13'h1907: dout <= 8'b11110111; // 6407 : 247 - 0xf7
      13'h1908: dout <= 8'b01000001; // 6408 :  65 - 0x41
      13'h1909: dout <= 8'b00001000; // 6409 :   8 - 0x8
      13'h190A: dout <= 8'b00000000; // 6410 :   0 - 0x0
      13'h190B: dout <= 8'b00100000; // 6411 :  32 - 0x20
      13'h190C: dout <= 8'b00000100; // 6412 :   4 - 0x4
      13'h190D: dout <= 8'b00000001; // 6413 :   1 - 0x1
      13'h190E: dout <= 8'b01000000; // 6414 :  64 - 0x40
      13'h190F: dout <= 8'b00001000; // 6415 :   8 - 0x8
      13'h1910: dout <= 8'b11101110; // 6416 : 238 - 0xee -- Background 0x91
      13'h1911: dout <= 8'b11111111; // 6417 : 255 - 0xff
      13'h1912: dout <= 8'b01111011; // 6418 : 123 - 0x7b
      13'h1913: dout <= 8'b11111101; // 6419 : 253 - 0xfd
      13'h1914: dout <= 8'b11101111; // 6420 : 239 - 0xef
      13'h1915: dout <= 8'b11111111; // 6421 : 255 - 0xff
      13'h1916: dout <= 8'b10111101; // 6422 : 189 - 0xbd
      13'h1917: dout <= 8'b11111111; // 6423 : 255 - 0xff
      13'h1918: dout <= 8'b00010001; // 6424 :  17 - 0x11
      13'h1919: dout <= 8'b00000000; // 6425 :   0 - 0x0
      13'h191A: dout <= 8'b10000100; // 6426 : 132 - 0x84
      13'h191B: dout <= 8'b00000010; // 6427 :   2 - 0x2
      13'h191C: dout <= 8'b00010000; // 6428 :  16 - 0x10
      13'h191D: dout <= 8'b00000000; // 6429 :   0 - 0x0
      13'h191E: dout <= 8'b01000010; // 6430 :  66 - 0x42
      13'h191F: dout <= 8'b00000000; // 6431 :   0 - 0x0
      13'h1920: dout <= 8'b11111011; // 6432 : 251 - 0xfb -- Background 0x92
      13'h1921: dout <= 8'b10111111; // 6433 : 191 - 0xbf
      13'h1922: dout <= 8'b11101111; // 6434 : 239 - 0xef
      13'h1923: dout <= 8'b11111101; // 6435 : 253 - 0xfd
      13'h1924: dout <= 8'b11111111; // 6436 : 255 - 0xff
      13'h1925: dout <= 8'b10111111; // 6437 : 191 - 0xbf
      13'h1926: dout <= 8'b11111011; // 6438 : 251 - 0xfb
      13'h1927: dout <= 8'b11011111; // 6439 : 223 - 0xdf
      13'h1928: dout <= 8'b00000100; // 6440 :   4 - 0x4
      13'h1929: dout <= 8'b01000000; // 6441 :  64 - 0x40
      13'h192A: dout <= 8'b00010000; // 6442 :  16 - 0x10
      13'h192B: dout <= 8'b00000010; // 6443 :   2 - 0x2
      13'h192C: dout <= 8'b00000000; // 6444 :   0 - 0x0
      13'h192D: dout <= 8'b01000000; // 6445 :  64 - 0x40
      13'h192E: dout <= 8'b00000100; // 6446 :   4 - 0x4
      13'h192F: dout <= 8'b00100000; // 6447 :  32 - 0x20
      13'h1930: dout <= 8'b10111101; // 6448 : 189 - 0xbd -- Background 0x93
      13'h1931: dout <= 8'b11111111; // 6449 : 255 - 0xff
      13'h1932: dout <= 8'b01110111; // 6450 : 119 - 0x77
      13'h1933: dout <= 8'b11111110; // 6451 : 254 - 0xfe
      13'h1934: dout <= 8'b11011111; // 6452 : 223 - 0xdf
      13'h1935: dout <= 8'b11111011; // 6453 : 251 - 0xfb
      13'h1936: dout <= 8'b11101111; // 6454 : 239 - 0xef
      13'h1937: dout <= 8'b01111111; // 6455 : 127 - 0x7f
      13'h1938: dout <= 8'b01000010; // 6456 :  66 - 0x42
      13'h1939: dout <= 8'b00000000; // 6457 :   0 - 0x0
      13'h193A: dout <= 8'b10001000; // 6458 : 136 - 0x88
      13'h193B: dout <= 8'b00000001; // 6459 :   1 - 0x1
      13'h193C: dout <= 8'b00100000; // 6460 :  32 - 0x20
      13'h193D: dout <= 8'b00000100; // 6461 :   4 - 0x4
      13'h193E: dout <= 8'b00010000; // 6462 :  16 - 0x10
      13'h193F: dout <= 8'b10000000; // 6463 : 128 - 0x80
      13'h1940: dout <= 8'b01111111; // 6464 : 127 - 0x7f -- Background 0x94
      13'h1941: dout <= 8'b11110111; // 6465 : 247 - 0xf7
      13'h1942: dout <= 8'b11011101; // 6466 : 221 - 0xdd
      13'h1943: dout <= 8'b01111011; // 6467 : 123 - 0x7b
      13'h1944: dout <= 8'b11111111; // 6468 : 255 - 0xff
      13'h1945: dout <= 8'b11101110; // 6469 : 238 - 0xee
      13'h1946: dout <= 8'b10111011; // 6470 : 187 - 0xbb
      13'h1947: dout <= 8'b11111101; // 6471 : 253 - 0xfd
      13'h1948: dout <= 8'b11001000; // 6472 : 200 - 0xc8
      13'h1949: dout <= 8'b00101010; // 6473 :  42 - 0x2a
      13'h194A: dout <= 8'b10100010; // 6474 : 162 - 0xa2
      13'h194B: dout <= 8'b10010100; // 6475 : 148 - 0x94
      13'h194C: dout <= 8'b10010001; // 6476 : 145 - 0x91
      13'h194D: dout <= 8'b01010101; // 6477 :  85 - 0x55
      13'h194E: dout <= 8'b01000100; // 6478 :  68 - 0x44
      13'h194F: dout <= 8'b00010010; // 6479 :  18 - 0x12
      13'h1950: dout <= 8'b11010111; // 6480 : 215 - 0xd7 -- Background 0x95
      13'h1951: dout <= 8'b01111111; // 6481 : 127 - 0x7f
      13'h1952: dout <= 8'b11111101; // 6482 : 253 - 0xfd
      13'h1953: dout <= 8'b11101110; // 6483 : 238 - 0xee
      13'h1954: dout <= 8'b11110111; // 6484 : 247 - 0xf7
      13'h1955: dout <= 8'b10111011; // 6485 : 187 - 0xbb
      13'h1956: dout <= 8'b11101111; // 6486 : 239 - 0xef
      13'h1957: dout <= 8'b11110111; // 6487 : 247 - 0xf7
      13'h1958: dout <= 8'b10101010; // 6488 : 170 - 0xaa
      13'h1959: dout <= 8'b10100010; // 6489 : 162 - 0xa2
      13'h195A: dout <= 8'b00010010; // 6490 :  18 - 0x12
      13'h195B: dout <= 8'b01010011; // 6491 :  83 - 0x53
      13'h195C: dout <= 8'b01001100; // 6492 :  76 - 0x4c
      13'h195D: dout <= 8'b01010101; // 6493 :  85 - 0x55
      13'h195E: dout <= 8'b10010001; // 6494 : 145 - 0x91
      13'h195F: dout <= 8'b01001000; // 6495 :  72 - 0x48
      13'h1960: dout <= 8'b10111111; // 6496 : 191 - 0xbf -- Background 0x96
      13'h1961: dout <= 8'b11101110; // 6497 : 238 - 0xee
      13'h1962: dout <= 8'b11011011; // 6498 : 219 - 0xdb
      13'h1963: dout <= 8'b11111111; // 6499 : 255 - 0xff
      13'h1964: dout <= 8'b01110111; // 6500 : 119 - 0x77
      13'h1965: dout <= 8'b11011101; // 6501 : 221 - 0xdd
      13'h1966: dout <= 8'b11101111; // 6502 : 239 - 0xef
      13'h1967: dout <= 8'b11111011; // 6503 : 251 - 0xfb
      13'h1968: dout <= 8'b01010001; // 6504 :  81 - 0x51
      13'h1969: dout <= 8'b00010101; // 6505 :  21 - 0x15
      13'h196A: dout <= 8'b10100100; // 6506 : 164 - 0xa4
      13'h196B: dout <= 8'b10001100; // 6507 : 140 - 0x8c
      13'h196C: dout <= 8'b10101010; // 6508 : 170 - 0xaa
      13'h196D: dout <= 8'b00100010; // 6509 :  34 - 0x22
      13'h196E: dout <= 8'b10010000; // 6510 : 144 - 0x90
      13'h196F: dout <= 8'b01000110; // 6511 :  70 - 0x46
      13'h1970: dout <= 8'b11111101; // 6512 : 253 - 0xfd -- Background 0x97
      13'h1971: dout <= 8'b11101110; // 6513 : 238 - 0xee
      13'h1972: dout <= 8'b11111011; // 6514 : 251 - 0xfb
      13'h1973: dout <= 8'b11111101; // 6515 : 253 - 0xfd
      13'h1974: dout <= 8'b11110101; // 6516 : 245 - 0xf5
      13'h1975: dout <= 8'b11011111; // 6517 : 223 - 0xdf
      13'h1976: dout <= 8'b01111111; // 6518 : 127 - 0x7f
      13'h1977: dout <= 8'b10111011; // 6519 : 187 - 0xbb
      13'h1978: dout <= 8'b00010011; // 6520 :  19 - 0x13
      13'h1979: dout <= 8'b01010101; // 6521 :  85 - 0x55
      13'h197A: dout <= 8'b01100100; // 6522 : 100 - 0x64
      13'h197B: dout <= 8'b00010010; // 6523 :  18 - 0x12
      13'h197C: dout <= 8'b10101010; // 6524 : 170 - 0xaa
      13'h197D: dout <= 8'b10101000; // 6525 : 168 - 0xa8
      13'h197E: dout <= 8'b10000100; // 6526 : 132 - 0x84
      13'h197F: dout <= 8'b11010100; // 6527 : 212 - 0xd4
      13'h1980: dout <= 8'b11111111; // 6528 : 255 - 0xff -- Background 0x98
      13'h1981: dout <= 8'b10011111; // 6529 : 159 - 0x9f
      13'h1982: dout <= 8'b10111111; // 6530 : 191 - 0xbf
      13'h1983: dout <= 8'b11110011; // 6531 : 243 - 0xf3
      13'h1984: dout <= 8'b11110011; // 6532 : 243 - 0xf3
      13'h1985: dout <= 8'b11111111; // 6533 : 255 - 0xff
      13'h1986: dout <= 8'b11111111; // 6534 : 255 - 0xff
      13'h1987: dout <= 8'b11111111; // 6535 : 255 - 0xff
      13'h1988: dout <= 8'b01100000; // 6536 :  96 - 0x60
      13'h1989: dout <= 8'b11110000; // 6537 : 240 - 0xf0
      13'h198A: dout <= 8'b11111110; // 6538 : 254 - 0xfe
      13'h198B: dout <= 8'b01111111; // 6539 : 127 - 0x7f
      13'h198C: dout <= 8'b00011111; // 6540 :  31 - 0x1f
      13'h198D: dout <= 8'b00011111; // 6541 :  31 - 0x1f
      13'h198E: dout <= 8'b00001110; // 6542 :  14 - 0xe
      13'h198F: dout <= 8'b00000000; // 6543 :   0 - 0x0
      13'h1990: dout <= 8'b11111111; // 6544 : 255 - 0xff -- Background 0x99
      13'h1991: dout <= 8'b10011111; // 6545 : 159 - 0x9f
      13'h1992: dout <= 8'b10111111; // 6546 : 191 - 0xbf
      13'h1993: dout <= 8'b11111111; // 6547 : 255 - 0xff
      13'h1994: dout <= 8'b11110011; // 6548 : 243 - 0xf3
      13'h1995: dout <= 8'b11110011; // 6549 : 243 - 0xf3
      13'h1996: dout <= 8'b11111111; // 6550 : 255 - 0xff
      13'h1997: dout <= 8'b11111111; // 6551 : 255 - 0xff
      13'h1998: dout <= 8'b01100000; // 6552 :  96 - 0x60
      13'h1999: dout <= 8'b11110000; // 6553 : 240 - 0xf0
      13'h199A: dout <= 8'b11110000; // 6554 : 240 - 0xf0
      13'h199B: dout <= 8'b01101110; // 6555 : 110 - 0x6e
      13'h199C: dout <= 8'b00011111; // 6556 :  31 - 0x1f
      13'h199D: dout <= 8'b00011111; // 6557 :  31 - 0x1f
      13'h199E: dout <= 8'b00011111; // 6558 :  31 - 0x1f
      13'h199F: dout <= 8'b00001110; // 6559 :  14 - 0xe
      13'h19A0: dout <= 8'b10111111; // 6560 : 191 - 0xbf -- Background 0x9a
      13'h19A1: dout <= 8'b11110111; // 6561 : 247 - 0xf7
      13'h19A2: dout <= 8'b11111111; // 6562 : 255 - 0xff
      13'h19A3: dout <= 8'b11011111; // 6563 : 223 - 0xdf
      13'h19A4: dout <= 8'b11111011; // 6564 : 251 - 0xfb
      13'h19A5: dout <= 8'b11111111; // 6565 : 255 - 0xff
      13'h19A6: dout <= 8'b10111111; // 6566 : 191 - 0xbf
      13'h19A7: dout <= 8'b11110111; // 6567 : 247 - 0xf7
      13'h19A8: dout <= 8'b01000000; // 6568 :  64 - 0x40
      13'h19A9: dout <= 8'b00001100; // 6569 :  12 - 0xc
      13'h19AA: dout <= 8'b00000000; // 6570 :   0 - 0x0
      13'h19AB: dout <= 8'b00101000; // 6571 :  40 - 0x28
      13'h19AC: dout <= 8'b00101100; // 6572 :  44 - 0x2c
      13'h19AD: dout <= 8'b00010001; // 6573 :  17 - 0x11
      13'h19AE: dout <= 8'b01000000; // 6574 :  64 - 0x40
      13'h19AF: dout <= 8'b00001000; // 6575 :   8 - 0x8
      13'h19B0: dout <= 8'b11011111; // 6576 : 223 - 0xdf -- Background 0x9b
      13'h19B1: dout <= 8'b11111111; // 6577 : 255 - 0xff
      13'h19B2: dout <= 8'b01111011; // 6578 : 123 - 0x7b
      13'h19B3: dout <= 8'b11111111; // 6579 : 255 - 0xff
      13'h19B4: dout <= 8'b11101111; // 6580 : 239 - 0xef
      13'h19B5: dout <= 8'b11111101; // 6581 : 253 - 0xfd
      13'h19B6: dout <= 8'b10111111; // 6582 : 191 - 0xbf
      13'h19B7: dout <= 8'b11111111; // 6583 : 255 - 0xff
      13'h19B8: dout <= 8'b00100000; // 6584 :  32 - 0x20
      13'h19B9: dout <= 8'b00000000; // 6585 :   0 - 0x0
      13'h19BA: dout <= 8'b10010100; // 6586 : 148 - 0x94
      13'h19BB: dout <= 8'b01001000; // 6587 :  72 - 0x48
      13'h19BC: dout <= 8'b00011000; // 6588 :  24 - 0x18
      13'h19BD: dout <= 8'b00000110; // 6589 :   6 - 0x6
      13'h19BE: dout <= 8'b01000000; // 6590 :  64 - 0x40
      13'h19BF: dout <= 8'b00000000; // 6591 :   0 - 0x0
      13'h19C0: dout <= 8'b10111010; // 6592 : 186 - 0xba -- Background 0x9c
      13'h19C1: dout <= 8'b10011100; // 6593 : 156 - 0x9c
      13'h19C2: dout <= 8'b10101010; // 6594 : 170 - 0xaa
      13'h19C3: dout <= 8'b11000000; // 6595 : 192 - 0xc0
      13'h19C4: dout <= 8'b11000000; // 6596 : 192 - 0xc0
      13'h19C5: dout <= 8'b11100000; // 6597 : 224 - 0xe0
      13'h19C6: dout <= 8'b11111000; // 6598 : 248 - 0xf8
      13'h19C7: dout <= 8'b11111111; // 6599 : 255 - 0xff
      13'h19C8: dout <= 8'b01111111; // 6600 : 127 - 0x7f
      13'h19C9: dout <= 8'b01111111; // 6601 : 127 - 0x7f
      13'h19CA: dout <= 8'b01111111; // 6602 : 127 - 0x7f
      13'h19CB: dout <= 8'b00111111; // 6603 :  63 - 0x3f
      13'h19CC: dout <= 8'b00110101; // 6604 :  53 - 0x35
      13'h19CD: dout <= 8'b00000010; // 6605 :   2 - 0x2
      13'h19CE: dout <= 8'b00000000; // 6606 :   0 - 0x0
      13'h19CF: dout <= 8'b00000000; // 6607 :   0 - 0x0
      13'h19D0: dout <= 8'b00000001; // 6608 :   1 - 0x1 -- Background 0x9d
      13'h19D1: dout <= 8'b00000001; // 6609 :   1 - 0x1
      13'h19D2: dout <= 8'b00000001; // 6610 :   1 - 0x1
      13'h19D3: dout <= 8'b00000011; // 6611 :   3 - 0x3
      13'h19D4: dout <= 8'b00000011; // 6612 :   3 - 0x3
      13'h19D5: dout <= 8'b00000111; // 6613 :   7 - 0x7
      13'h19D6: dout <= 8'b00011111; // 6614 :  31 - 0x1f
      13'h19D7: dout <= 8'b11111111; // 6615 : 255 - 0xff
      13'h19D8: dout <= 8'b11110100; // 6616 : 244 - 0xf4
      13'h19D9: dout <= 8'b11111000; // 6617 : 248 - 0xf8
      13'h19DA: dout <= 8'b11110000; // 6618 : 240 - 0xf0
      13'h19DB: dout <= 8'b11101000; // 6619 : 232 - 0xe8
      13'h19DC: dout <= 8'b01010000; // 6620 :  80 - 0x50
      13'h19DD: dout <= 8'b10000000; // 6621 : 128 - 0x80
      13'h19DE: dout <= 8'b00000000; // 6622 :   0 - 0x0
      13'h19DF: dout <= 8'b00000000; // 6623 :   0 - 0x0
      13'h19E0: dout <= 8'b01111101; // 6624 : 125 - 0x7d -- Background 0x9e
      13'h19E1: dout <= 8'b11111111; // 6625 : 255 - 0xff
      13'h19E2: dout <= 8'b11111011; // 6626 : 251 - 0xfb
      13'h19E3: dout <= 8'b11111111; // 6627 : 255 - 0xff
      13'h19E4: dout <= 8'b11111111; // 6628 : 255 - 0xff
      13'h19E5: dout <= 8'b11111011; // 6629 : 251 - 0xfb
      13'h19E6: dout <= 8'b11111111; // 6630 : 255 - 0xff
      13'h19E7: dout <= 8'b01111101; // 6631 : 125 - 0x7d
      13'h19E8: dout <= 8'b11111110; // 6632 : 254 - 0xfe
      13'h19E9: dout <= 8'b11111100; // 6633 : 252 - 0xfc
      13'h19EA: dout <= 8'b11111100; // 6634 : 252 - 0xfc
      13'h19EB: dout <= 8'b11111000; // 6635 : 248 - 0xf8
      13'h19EC: dout <= 8'b11111000; // 6636 : 248 - 0xf8
      13'h19ED: dout <= 8'b11111100; // 6637 : 252 - 0xfc
      13'h19EE: dout <= 8'b11111100; // 6638 : 252 - 0xfc
      13'h19EF: dout <= 8'b11111110; // 6639 : 254 - 0xfe
      13'h19F0: dout <= 8'b11111111; // 6640 : 255 - 0xff -- Background 0x9f
      13'h19F1: dout <= 8'b11111111; // 6641 : 255 - 0xff
      13'h19F2: dout <= 8'b10111101; // 6642 : 189 - 0xbd
      13'h19F3: dout <= 8'b11111111; // 6643 : 255 - 0xff
      13'h19F4: dout <= 8'b11111111; // 6644 : 255 - 0xff
      13'h19F5: dout <= 8'b11111111; // 6645 : 255 - 0xff
      13'h19F6: dout <= 8'b11111111; // 6646 : 255 - 0xff
      13'h19F7: dout <= 8'b10111101; // 6647 : 189 - 0xbd
      13'h19F8: dout <= 8'b00000000; // 6648 :   0 - 0x0
      13'h19F9: dout <= 8'b00000000; // 6649 :   0 - 0x0
      13'h19FA: dout <= 8'b01111110; // 6650 : 126 - 0x7e
      13'h19FB: dout <= 8'b01111110; // 6651 : 126 - 0x7e
      13'h19FC: dout <= 8'b01111110; // 6652 : 126 - 0x7e
      13'h19FD: dout <= 8'b01111110; // 6653 : 126 - 0x7e
      13'h19FE: dout <= 8'b01111110; // 6654 : 126 - 0x7e
      13'h19FF: dout <= 8'b01111110; // 6655 : 126 - 0x7e
      13'h1A00: dout <= 8'b11101111; // 6656 : 239 - 0xef -- Background 0xa0
      13'h1A01: dout <= 8'b11000111; // 6657 : 199 - 0xc7
      13'h1A02: dout <= 8'b10000011; // 6658 : 131 - 0x83
      13'h1A03: dout <= 8'b00000111; // 6659 :   7 - 0x7
      13'h1A04: dout <= 8'b10001111; // 6660 : 143 - 0x8f
      13'h1A05: dout <= 8'b11011101; // 6661 : 221 - 0xdd
      13'h1A06: dout <= 8'b11111010; // 6662 : 250 - 0xfa
      13'h1A07: dout <= 8'b11111101; // 6663 : 253 - 0xfd
      13'h1A08: dout <= 8'b00010000; // 6664 :  16 - 0x10
      13'h1A09: dout <= 8'b00111000; // 6665 :  56 - 0x38
      13'h1A0A: dout <= 8'b01111100; // 6666 : 124 - 0x7c
      13'h1A0B: dout <= 8'b11111000; // 6667 : 248 - 0xf8
      13'h1A0C: dout <= 8'b01110000; // 6668 : 112 - 0x70
      13'h1A0D: dout <= 8'b00100010; // 6669 :  34 - 0x22
      13'h1A0E: dout <= 8'b00000101; // 6670 :   5 - 0x5
      13'h1A0F: dout <= 8'b00000010; // 6671 :   2 - 0x2
      13'h1A10: dout <= 8'b11101111; // 6672 : 239 - 0xef -- Background 0xa1
      13'h1A11: dout <= 8'b11000111; // 6673 : 199 - 0xc7
      13'h1A12: dout <= 8'b10000011; // 6674 : 131 - 0x83
      13'h1A13: dout <= 8'b00011111; // 6675 :  31 - 0x1f
      13'h1A14: dout <= 8'b10010000; // 6676 : 144 - 0x90
      13'h1A15: dout <= 8'b11010100; // 6677 : 212 - 0xd4
      13'h1A16: dout <= 8'b11110011; // 6678 : 243 - 0xf3
      13'h1A17: dout <= 8'b11110010; // 6679 : 242 - 0xf2
      13'h1A18: dout <= 8'b00010000; // 6680 :  16 - 0x10
      13'h1A19: dout <= 8'b00111000; // 6681 :  56 - 0x38
      13'h1A1A: dout <= 8'b01111100; // 6682 : 124 - 0x7c
      13'h1A1B: dout <= 8'b11100000; // 6683 : 224 - 0xe0
      13'h1A1C: dout <= 8'b01100000; // 6684 :  96 - 0x60
      13'h1A1D: dout <= 8'b00100000; // 6685 :  32 - 0x20
      13'h1A1E: dout <= 8'b00000000; // 6686 :   0 - 0x0
      13'h1A1F: dout <= 8'b00000000; // 6687 :   0 - 0x0
      13'h1A20: dout <= 8'b11101111; // 6688 : 239 - 0xef -- Background 0xa2
      13'h1A21: dout <= 8'b11000111; // 6689 : 199 - 0xc7
      13'h1A22: dout <= 8'b10000011; // 6690 : 131 - 0x83
      13'h1A23: dout <= 8'b11111111; // 6691 : 255 - 0xff
      13'h1A24: dout <= 8'b00000000; // 6692 :   0 - 0x0
      13'h1A25: dout <= 8'b00000000; // 6693 :   0 - 0x0
      13'h1A26: dout <= 8'b01010101; // 6694 :  85 - 0x55
      13'h1A27: dout <= 8'b00000000; // 6695 :   0 - 0x0
      13'h1A28: dout <= 8'b00010000; // 6696 :  16 - 0x10
      13'h1A29: dout <= 8'b00111000; // 6697 :  56 - 0x38
      13'h1A2A: dout <= 8'b01111100; // 6698 : 124 - 0x7c
      13'h1A2B: dout <= 8'b00000000; // 6699 :   0 - 0x0
      13'h1A2C: dout <= 8'b00000000; // 6700 :   0 - 0x0
      13'h1A2D: dout <= 8'b00000000; // 6701 :   0 - 0x0
      13'h1A2E: dout <= 8'b00000000; // 6702 :   0 - 0x0
      13'h1A2F: dout <= 8'b00000000; // 6703 :   0 - 0x0
      13'h1A30: dout <= 8'b11110000; // 6704 : 240 - 0xf0 -- Background 0xa3
      13'h1A31: dout <= 8'b11010010; // 6705 : 210 - 0xd2
      13'h1A32: dout <= 8'b10010000; // 6706 : 144 - 0x90
      13'h1A33: dout <= 8'b00010010; // 6707 :  18 - 0x12
      13'h1A34: dout <= 8'b10010000; // 6708 : 144 - 0x90
      13'h1A35: dout <= 8'b11010010; // 6709 : 210 - 0xd2
      13'h1A36: dout <= 8'b11110000; // 6710 : 240 - 0xf0
      13'h1A37: dout <= 8'b11110010; // 6711 : 242 - 0xf2
      13'h1A38: dout <= 8'b00000000; // 6712 :   0 - 0x0
      13'h1A39: dout <= 8'b00100000; // 6713 :  32 - 0x20
      13'h1A3A: dout <= 8'b01100000; // 6714 :  96 - 0x60
      13'h1A3B: dout <= 8'b11100000; // 6715 : 224 - 0xe0
      13'h1A3C: dout <= 8'b01100000; // 6716 :  96 - 0x60
      13'h1A3D: dout <= 8'b00100000; // 6717 :  32 - 0x20
      13'h1A3E: dout <= 8'b00000000; // 6718 :   0 - 0x0
      13'h1A3F: dout <= 8'b00000000; // 6719 :   0 - 0x0
      13'h1A40: dout <= 8'b11110000; // 6720 : 240 - 0xf0 -- Background 0xa4
      13'h1A41: dout <= 8'b11010011; // 6721 : 211 - 0xd3
      13'h1A42: dout <= 8'b10010100; // 6722 : 148 - 0x94
      13'h1A43: dout <= 8'b00011000; // 6723 :  24 - 0x18
      13'h1A44: dout <= 8'b10011111; // 6724 : 159 - 0x9f
      13'h1A45: dout <= 8'b11011101; // 6725 : 221 - 0xdd
      13'h1A46: dout <= 8'b11111010; // 6726 : 250 - 0xfa
      13'h1A47: dout <= 8'b11111101; // 6727 : 253 - 0xfd
      13'h1A48: dout <= 8'b00000000; // 6728 :   0 - 0x0
      13'h1A49: dout <= 8'b00100000; // 6729 :  32 - 0x20
      13'h1A4A: dout <= 8'b01100011; // 6730 :  99 - 0x63
      13'h1A4B: dout <= 8'b11100111; // 6731 : 231 - 0xe7
      13'h1A4C: dout <= 8'b01100000; // 6732 :  96 - 0x60
      13'h1A4D: dout <= 8'b00100010; // 6733 :  34 - 0x22
      13'h1A4E: dout <= 8'b00000101; // 6734 :   5 - 0x5
      13'h1A4F: dout <= 8'b00000010; // 6735 :   2 - 0x2
      13'h1A50: dout <= 8'b00000000; // 6736 :   0 - 0x0 -- Background 0xa5
      13'h1A51: dout <= 8'b11111111; // 6737 : 255 - 0xff
      13'h1A52: dout <= 8'b00000000; // 6738 :   0 - 0x0
      13'h1A53: dout <= 8'b00000000; // 6739 :   0 - 0x0
      13'h1A54: dout <= 8'b11111111; // 6740 : 255 - 0xff
      13'h1A55: dout <= 8'b11011101; // 6741 : 221 - 0xdd
      13'h1A56: dout <= 8'b11111010; // 6742 : 250 - 0xfa
      13'h1A57: dout <= 8'b11111101; // 6743 : 253 - 0xfd
      13'h1A58: dout <= 8'b00000000; // 6744 :   0 - 0x0
      13'h1A59: dout <= 8'b00000000; // 6745 :   0 - 0x0
      13'h1A5A: dout <= 8'b11111111; // 6746 : 255 - 0xff
      13'h1A5B: dout <= 8'b11111111; // 6747 : 255 - 0xff
      13'h1A5C: dout <= 8'b00000000; // 6748 :   0 - 0x0
      13'h1A5D: dout <= 8'b00100010; // 6749 :  34 - 0x22
      13'h1A5E: dout <= 8'b00000101; // 6750 :   5 - 0x5
      13'h1A5F: dout <= 8'b00000010; // 6751 :   2 - 0x2
      13'h1A60: dout <= 8'b11101111; // 6752 : 239 - 0xef -- Background 0xa6
      13'h1A61: dout <= 8'b11000111; // 6753 : 199 - 0xc7
      13'h1A62: dout <= 8'b10000011; // 6754 : 131 - 0x83
      13'h1A63: dout <= 8'b11111111; // 6755 : 255 - 0xff
      13'h1A64: dout <= 8'b00011111; // 6756 :  31 - 0x1f
      13'h1A65: dout <= 8'b00101101; // 6757 :  45 - 0x2d
      13'h1A66: dout <= 8'b01001010; // 6758 :  74 - 0x4a
      13'h1A67: dout <= 8'b01001101; // 6759 :  77 - 0x4d
      13'h1A68: dout <= 8'b00010000; // 6760 :  16 - 0x10
      13'h1A69: dout <= 8'b00111000; // 6761 :  56 - 0x38
      13'h1A6A: dout <= 8'b01111100; // 6762 : 124 - 0x7c
      13'h1A6B: dout <= 8'b00000000; // 6763 :   0 - 0x0
      13'h1A6C: dout <= 8'b00000000; // 6764 :   0 - 0x0
      13'h1A6D: dout <= 8'b00010010; // 6765 :  18 - 0x12
      13'h1A6E: dout <= 8'b00110101; // 6766 :  53 - 0x35
      13'h1A6F: dout <= 8'b00110010; // 6767 :  50 - 0x32
      13'h1A70: dout <= 8'b01001111; // 6768 :  79 - 0x4f -- Background 0xa7
      13'h1A71: dout <= 8'b01001111; // 6769 :  79 - 0x4f
      13'h1A72: dout <= 8'b01001011; // 6770 :  75 - 0x4b
      13'h1A73: dout <= 8'b01001111; // 6771 :  79 - 0x4f
      13'h1A74: dout <= 8'b01001111; // 6772 :  79 - 0x4f
      13'h1A75: dout <= 8'b01001101; // 6773 :  77 - 0x4d
      13'h1A76: dout <= 8'b01001010; // 6774 :  74 - 0x4a
      13'h1A77: dout <= 8'b01001101; // 6775 :  77 - 0x4d
      13'h1A78: dout <= 8'b00110000; // 6776 :  48 - 0x30
      13'h1A79: dout <= 8'b00110000; // 6777 :  48 - 0x30
      13'h1A7A: dout <= 8'b00110100; // 6778 :  52 - 0x34
      13'h1A7B: dout <= 8'b00110000; // 6779 :  48 - 0x30
      13'h1A7C: dout <= 8'b00110000; // 6780 :  48 - 0x30
      13'h1A7D: dout <= 8'b00110010; // 6781 :  50 - 0x32
      13'h1A7E: dout <= 8'b00110101; // 6782 :  53 - 0x35
      13'h1A7F: dout <= 8'b00110010; // 6783 :  50 - 0x32
      13'h1A80: dout <= 8'b01001111; // 6784 :  79 - 0x4f -- Background 0xa8
      13'h1A81: dout <= 8'b11001111; // 6785 : 207 - 0xcf
      13'h1A82: dout <= 8'b00001011; // 6786 :  11 - 0xb
      13'h1A83: dout <= 8'b00001111; // 6787 :  15 - 0xf
      13'h1A84: dout <= 8'b11111111; // 6788 : 255 - 0xff
      13'h1A85: dout <= 8'b11011101; // 6789 : 221 - 0xdd
      13'h1A86: dout <= 8'b11111010; // 6790 : 250 - 0xfa
      13'h1A87: dout <= 8'b11111101; // 6791 : 253 - 0xfd
      13'h1A88: dout <= 8'b00110000; // 6792 :  48 - 0x30
      13'h1A89: dout <= 8'b00110000; // 6793 :  48 - 0x30
      13'h1A8A: dout <= 8'b11110100; // 6794 : 244 - 0xf4
      13'h1A8B: dout <= 8'b11110000; // 6795 : 240 - 0xf0
      13'h1A8C: dout <= 8'b00000000; // 6796 :   0 - 0x0
      13'h1A8D: dout <= 8'b00100010; // 6797 :  34 - 0x22
      13'h1A8E: dout <= 8'b00000101; // 6798 :   5 - 0x5
      13'h1A8F: dout <= 8'b00000010; // 6799 :   2 - 0x2
      13'h1A90: dout <= 8'b11111111; // 6800 : 255 - 0xff -- Background 0xa9
      13'h1A91: dout <= 8'b11111111; // 6801 : 255 - 0xff
      13'h1A92: dout <= 8'b11111111; // 6802 : 255 - 0xff
      13'h1A93: dout <= 8'b11111111; // 6803 : 255 - 0xff
      13'h1A94: dout <= 8'b11111111; // 6804 : 255 - 0xff
      13'h1A95: dout <= 8'b11111111; // 6805 : 255 - 0xff
      13'h1A96: dout <= 8'b11111111; // 6806 : 255 - 0xff
      13'h1A97: dout <= 8'b11111111; // 6807 : 255 - 0xff
      13'h1A98: dout <= 8'b00000000; // 6808 :   0 - 0x0
      13'h1A99: dout <= 8'b00000000; // 6809 :   0 - 0x0
      13'h1A9A: dout <= 8'b00000000; // 6810 :   0 - 0x0
      13'h1A9B: dout <= 8'b00000000; // 6811 :   0 - 0x0
      13'h1A9C: dout <= 8'b00000000; // 6812 :   0 - 0x0
      13'h1A9D: dout <= 8'b00000000; // 6813 :   0 - 0x0
      13'h1A9E: dout <= 8'b00000000; // 6814 :   0 - 0x0
      13'h1A9F: dout <= 8'b00000000; // 6815 :   0 - 0x0
      13'h1AA0: dout <= 8'b11111111; // 6816 : 255 - 0xff -- Background 0xaa
      13'h1AA1: dout <= 8'b11111111; // 6817 : 255 - 0xff
      13'h1AA2: dout <= 8'b10101111; // 6818 : 175 - 0xaf
      13'h1AA3: dout <= 8'b01010111; // 6819 :  87 - 0x57
      13'h1AA4: dout <= 8'b10001111; // 6820 : 143 - 0x8f
      13'h1AA5: dout <= 8'b11011101; // 6821 : 221 - 0xdd
      13'h1AA6: dout <= 8'b11111010; // 6822 : 250 - 0xfa
      13'h1AA7: dout <= 8'b11111101; // 6823 : 253 - 0xfd
      13'h1AA8: dout <= 8'b00000000; // 6824 :   0 - 0x0
      13'h1AA9: dout <= 8'b00000000; // 6825 :   0 - 0x0
      13'h1AAA: dout <= 8'b01010000; // 6826 :  80 - 0x50
      13'h1AAB: dout <= 8'b10101000; // 6827 : 168 - 0xa8
      13'h1AAC: dout <= 8'b01110000; // 6828 : 112 - 0x70
      13'h1AAD: dout <= 8'b00100010; // 6829 :  34 - 0x22
      13'h1AAE: dout <= 8'b00000101; // 6830 :   5 - 0x5
      13'h1AAF: dout <= 8'b00000010; // 6831 :   2 - 0x2
      13'h1AB0: dout <= 8'b11111111; // 6832 : 255 - 0xff -- Background 0xab
      13'h1AB1: dout <= 8'b00000000; // 6833 :   0 - 0x0
      13'h1AB2: dout <= 8'b00000000; // 6834 :   0 - 0x0
      13'h1AB3: dout <= 8'b00000000; // 6835 :   0 - 0x0
      13'h1AB4: dout <= 8'b00000000; // 6836 :   0 - 0x0
      13'h1AB5: dout <= 8'b00000000; // 6837 :   0 - 0x0
      13'h1AB6: dout <= 8'b00000000; // 6838 :   0 - 0x0
      13'h1AB7: dout <= 8'b00000000; // 6839 :   0 - 0x0
      13'h1AB8: dout <= 8'b00000000; // 6840 :   0 - 0x0
      13'h1AB9: dout <= 8'b00000000; // 6841 :   0 - 0x0
      13'h1ABA: dout <= 8'b00000000; // 6842 :   0 - 0x0
      13'h1ABB: dout <= 8'b00000000; // 6843 :   0 - 0x0
      13'h1ABC: dout <= 8'b00000000; // 6844 :   0 - 0x0
      13'h1ABD: dout <= 8'b00000000; // 6845 :   0 - 0x0
      13'h1ABE: dout <= 8'b00000000; // 6846 :   0 - 0x0
      13'h1ABF: dout <= 8'b00000000; // 6847 :   0 - 0x0
      13'h1AC0: dout <= 8'b00000000; // 6848 :   0 - 0x0 -- Background 0xac
      13'h1AC1: dout <= 8'b00000000; // 6849 :   0 - 0x0
      13'h1AC2: dout <= 8'b00000000; // 6850 :   0 - 0x0
      13'h1AC3: dout <= 8'b00000000; // 6851 :   0 - 0x0
      13'h1AC4: dout <= 8'b00000000; // 6852 :   0 - 0x0
      13'h1AC5: dout <= 8'b00000000; // 6853 :   0 - 0x0
      13'h1AC6: dout <= 8'b00000000; // 6854 :   0 - 0x0
      13'h1AC7: dout <= 8'b00000000; // 6855 :   0 - 0x0
      13'h1AC8: dout <= 8'b00000000; // 6856 :   0 - 0x0
      13'h1AC9: dout <= 8'b00000000; // 6857 :   0 - 0x0
      13'h1ACA: dout <= 8'b00000000; // 6858 :   0 - 0x0
      13'h1ACB: dout <= 8'b00000000; // 6859 :   0 - 0x0
      13'h1ACC: dout <= 8'b00000000; // 6860 :   0 - 0x0
      13'h1ACD: dout <= 8'b00000000; // 6861 :   0 - 0x0
      13'h1ACE: dout <= 8'b00000000; // 6862 :   0 - 0x0
      13'h1ACF: dout <= 8'b00000000; // 6863 :   0 - 0x0
      13'h1AD0: dout <= 8'b00000000; // 6864 :   0 - 0x0 -- Background 0xad
      13'h1AD1: dout <= 8'b11111111; // 6865 : 255 - 0xff
      13'h1AD2: dout <= 8'b00000000; // 6866 :   0 - 0x0
      13'h1AD3: dout <= 8'b11111111; // 6867 : 255 - 0xff
      13'h1AD4: dout <= 8'b11111111; // 6868 : 255 - 0xff
      13'h1AD5: dout <= 8'b11111111; // 6869 : 255 - 0xff
      13'h1AD6: dout <= 8'b11111111; // 6870 : 255 - 0xff
      13'h1AD7: dout <= 8'b11111111; // 6871 : 255 - 0xff
      13'h1AD8: dout <= 8'b00000000; // 6872 :   0 - 0x0
      13'h1AD9: dout <= 8'b00000000; // 6873 :   0 - 0x0
      13'h1ADA: dout <= 8'b11111111; // 6874 : 255 - 0xff
      13'h1ADB: dout <= 8'b00000000; // 6875 :   0 - 0x0
      13'h1ADC: dout <= 8'b00000000; // 6876 :   0 - 0x0
      13'h1ADD: dout <= 8'b00000000; // 6877 :   0 - 0x0
      13'h1ADE: dout <= 8'b00000000; // 6878 :   0 - 0x0
      13'h1ADF: dout <= 8'b00000000; // 6879 :   0 - 0x0
      13'h1AE0: dout <= 8'b11111111; // 6880 : 255 - 0xff -- Background 0xae
      13'h1AE1: dout <= 8'b11111111; // 6881 : 255 - 0xff
      13'h1AE2: dout <= 8'b11111111; // 6882 : 255 - 0xff
      13'h1AE3: dout <= 8'b11111111; // 6883 : 255 - 0xff
      13'h1AE4: dout <= 8'b11111111; // 6884 : 255 - 0xff
      13'h1AE5: dout <= 8'b00000000; // 6885 :   0 - 0x0
      13'h1AE6: dout <= 8'b11111111; // 6886 : 255 - 0xff
      13'h1AE7: dout <= 8'b00000000; // 6887 :   0 - 0x0
      13'h1AE8: dout <= 8'b00000000; // 6888 :   0 - 0x0
      13'h1AE9: dout <= 8'b00000000; // 6889 :   0 - 0x0
      13'h1AEA: dout <= 8'b00000000; // 6890 :   0 - 0x0
      13'h1AEB: dout <= 8'b00000000; // 6891 :   0 - 0x0
      13'h1AEC: dout <= 8'b00000000; // 6892 :   0 - 0x0
      13'h1AED: dout <= 8'b11111111; // 6893 : 255 - 0xff
      13'h1AEE: dout <= 8'b00000000; // 6894 :   0 - 0x0
      13'h1AEF: dout <= 8'b00000000; // 6895 :   0 - 0x0
      13'h1AF0: dout <= 8'b11111111; // 6896 : 255 - 0xff -- Background 0xaf
      13'h1AF1: dout <= 8'b11111111; // 6897 : 255 - 0xff
      13'h1AF2: dout <= 8'b11111111; // 6898 : 255 - 0xff
      13'h1AF3: dout <= 8'b11111111; // 6899 : 255 - 0xff
      13'h1AF4: dout <= 8'b11111111; // 6900 : 255 - 0xff
      13'h1AF5: dout <= 8'b11111111; // 6901 : 255 - 0xff
      13'h1AF6: dout <= 8'b11111111; // 6902 : 255 - 0xff
      13'h1AF7: dout <= 8'b11111111; // 6903 : 255 - 0xff
      13'h1AF8: dout <= 8'b00000000; // 6904 :   0 - 0x0
      13'h1AF9: dout <= 8'b00000000; // 6905 :   0 - 0x0
      13'h1AFA: dout <= 8'b00000000; // 6906 :   0 - 0x0
      13'h1AFB: dout <= 8'b00000000; // 6907 :   0 - 0x0
      13'h1AFC: dout <= 8'b00000000; // 6908 :   0 - 0x0
      13'h1AFD: dout <= 8'b00000000; // 6909 :   0 - 0x0
      13'h1AFE: dout <= 8'b00000000; // 6910 :   0 - 0x0
      13'h1AFF: dout <= 8'b00000000; // 6911 :   0 - 0x0
      13'h1B00: dout <= 8'b00000000; // 6912 :   0 - 0x0 -- Background 0xb0
      13'h1B01: dout <= 8'b00000000; // 6913 :   0 - 0x0
      13'h1B02: dout <= 8'b00011111; // 6914 :  31 - 0x1f
      13'h1B03: dout <= 8'b00010000; // 6915 :  16 - 0x10
      13'h1B04: dout <= 8'b00010000; // 6916 :  16 - 0x10
      13'h1B05: dout <= 8'b00010000; // 6917 :  16 - 0x10
      13'h1B06: dout <= 8'b00010000; // 6918 :  16 - 0x10
      13'h1B07: dout <= 8'b00010000; // 6919 :  16 - 0x10
      13'h1B08: dout <= 8'b00000000; // 6920 :   0 - 0x0
      13'h1B09: dout <= 8'b00000000; // 6921 :   0 - 0x0
      13'h1B0A: dout <= 8'b00011111; // 6922 :  31 - 0x1f
      13'h1B0B: dout <= 8'b00011111; // 6923 :  31 - 0x1f
      13'h1B0C: dout <= 8'b00011111; // 6924 :  31 - 0x1f
      13'h1B0D: dout <= 8'b00011111; // 6925 :  31 - 0x1f
      13'h1B0E: dout <= 8'b00011111; // 6926 :  31 - 0x1f
      13'h1B0F: dout <= 8'b00011111; // 6927 :  31 - 0x1f
      13'h1B10: dout <= 8'b00000000; // 6928 :   0 - 0x0 -- Background 0xb1
      13'h1B11: dout <= 8'b00000000; // 6929 :   0 - 0x0
      13'h1B12: dout <= 8'b11111000; // 6930 : 248 - 0xf8
      13'h1B13: dout <= 8'b00001000; // 6931 :   8 - 0x8
      13'h1B14: dout <= 8'b00001000; // 6932 :   8 - 0x8
      13'h1B15: dout <= 8'b00001000; // 6933 :   8 - 0x8
      13'h1B16: dout <= 8'b00001000; // 6934 :   8 - 0x8
      13'h1B17: dout <= 8'b00001000; // 6935 :   8 - 0x8
      13'h1B18: dout <= 8'b00000000; // 6936 :   0 - 0x0
      13'h1B19: dout <= 8'b00000000; // 6937 :   0 - 0x0
      13'h1B1A: dout <= 8'b11110000; // 6938 : 240 - 0xf0
      13'h1B1B: dout <= 8'b11110000; // 6939 : 240 - 0xf0
      13'h1B1C: dout <= 8'b11110000; // 6940 : 240 - 0xf0
      13'h1B1D: dout <= 8'b11110000; // 6941 : 240 - 0xf0
      13'h1B1E: dout <= 8'b11110000; // 6942 : 240 - 0xf0
      13'h1B1F: dout <= 8'b11110000; // 6943 : 240 - 0xf0
      13'h1B20: dout <= 8'b00010000; // 6944 :  16 - 0x10 -- Background 0xb2
      13'h1B21: dout <= 8'b00010000; // 6945 :  16 - 0x10
      13'h1B22: dout <= 8'b00010000; // 6946 :  16 - 0x10
      13'h1B23: dout <= 8'b00010000; // 6947 :  16 - 0x10
      13'h1B24: dout <= 8'b00010000; // 6948 :  16 - 0x10
      13'h1B25: dout <= 8'b00011111; // 6949 :  31 - 0x1f
      13'h1B26: dout <= 8'b00011111; // 6950 :  31 - 0x1f
      13'h1B27: dout <= 8'b00001111; // 6951 :  15 - 0xf
      13'h1B28: dout <= 8'b00011111; // 6952 :  31 - 0x1f
      13'h1B29: dout <= 8'b00011111; // 6953 :  31 - 0x1f
      13'h1B2A: dout <= 8'b00011111; // 6954 :  31 - 0x1f
      13'h1B2B: dout <= 8'b00011111; // 6955 :  31 - 0x1f
      13'h1B2C: dout <= 8'b00011111; // 6956 :  31 - 0x1f
      13'h1B2D: dout <= 8'b00000000; // 6957 :   0 - 0x0
      13'h1B2E: dout <= 8'b00000000; // 6958 :   0 - 0x0
      13'h1B2F: dout <= 8'b00000000; // 6959 :   0 - 0x0
      13'h1B30: dout <= 8'b00001000; // 6960 :   8 - 0x8 -- Background 0xb3
      13'h1B31: dout <= 8'b00001000; // 6961 :   8 - 0x8
      13'h1B32: dout <= 8'b00001000; // 6962 :   8 - 0x8
      13'h1B33: dout <= 8'b00001000; // 6963 :   8 - 0x8
      13'h1B34: dout <= 8'b00001000; // 6964 :   8 - 0x8
      13'h1B35: dout <= 8'b11111000; // 6965 : 248 - 0xf8
      13'h1B36: dout <= 8'b11111000; // 6966 : 248 - 0xf8
      13'h1B37: dout <= 8'b11110000; // 6967 : 240 - 0xf0
      13'h1B38: dout <= 8'b11110000; // 6968 : 240 - 0xf0
      13'h1B39: dout <= 8'b11110000; // 6969 : 240 - 0xf0
      13'h1B3A: dout <= 8'b11110000; // 6970 : 240 - 0xf0
      13'h1B3B: dout <= 8'b11110000; // 6971 : 240 - 0xf0
      13'h1B3C: dout <= 8'b11110000; // 6972 : 240 - 0xf0
      13'h1B3D: dout <= 8'b00000000; // 6973 :   0 - 0x0
      13'h1B3E: dout <= 8'b00000000; // 6974 :   0 - 0x0
      13'h1B3F: dout <= 8'b00000000; // 6975 :   0 - 0x0
      13'h1B40: dout <= 8'b00000000; // 6976 :   0 - 0x0 -- Background 0xb4
      13'h1B41: dout <= 8'b00000000; // 6977 :   0 - 0x0
      13'h1B42: dout <= 8'b00000000; // 6978 :   0 - 0x0
      13'h1B43: dout <= 8'b00111111; // 6979 :  63 - 0x3f
      13'h1B44: dout <= 8'b01100000; // 6980 :  96 - 0x60
      13'h1B45: dout <= 8'b01100000; // 6981 :  96 - 0x60
      13'h1B46: dout <= 8'b01100000; // 6982 :  96 - 0x60
      13'h1B47: dout <= 8'b01100000; // 6983 :  96 - 0x60
      13'h1B48: dout <= 8'b00000000; // 6984 :   0 - 0x0
      13'h1B49: dout <= 8'b00000000; // 6985 :   0 - 0x0
      13'h1B4A: dout <= 8'b00000000; // 6986 :   0 - 0x0
      13'h1B4B: dout <= 8'b00111111; // 6987 :  63 - 0x3f
      13'h1B4C: dout <= 8'b01111111; // 6988 : 127 - 0x7f
      13'h1B4D: dout <= 8'b01111111; // 6989 : 127 - 0x7f
      13'h1B4E: dout <= 8'b01111111; // 6990 : 127 - 0x7f
      13'h1B4F: dout <= 8'b01111111; // 6991 : 127 - 0x7f
      13'h1B50: dout <= 8'b00000000; // 6992 :   0 - 0x0 -- Background 0xb5
      13'h1B51: dout <= 8'b00000000; // 6993 :   0 - 0x0
      13'h1B52: dout <= 8'b00000000; // 6994 :   0 - 0x0
      13'h1B53: dout <= 8'b11111100; // 6995 : 252 - 0xfc
      13'h1B54: dout <= 8'b00000110; // 6996 :   6 - 0x6
      13'h1B55: dout <= 8'b00000110; // 6997 :   6 - 0x6
      13'h1B56: dout <= 8'b00000110; // 6998 :   6 - 0x6
      13'h1B57: dout <= 8'b00000110; // 6999 :   6 - 0x6
      13'h1B58: dout <= 8'b00000000; // 7000 :   0 - 0x0
      13'h1B59: dout <= 8'b00000000; // 7001 :   0 - 0x0
      13'h1B5A: dout <= 8'b00000000; // 7002 :   0 - 0x0
      13'h1B5B: dout <= 8'b11111000; // 7003 : 248 - 0xf8
      13'h1B5C: dout <= 8'b11111000; // 7004 : 248 - 0xf8
      13'h1B5D: dout <= 8'b11111000; // 7005 : 248 - 0xf8
      13'h1B5E: dout <= 8'b11111000; // 7006 : 248 - 0xf8
      13'h1B5F: dout <= 8'b11111000; // 7007 : 248 - 0xf8
      13'h1B60: dout <= 8'b01100000; // 7008 :  96 - 0x60 -- Background 0xb6
      13'h1B61: dout <= 8'b01100000; // 7009 :  96 - 0x60
      13'h1B62: dout <= 8'b01100000; // 7010 :  96 - 0x60
      13'h1B63: dout <= 8'b01100000; // 7011 :  96 - 0x60
      13'h1B64: dout <= 8'b01111111; // 7012 : 127 - 0x7f
      13'h1B65: dout <= 8'b01111111; // 7013 : 127 - 0x7f
      13'h1B66: dout <= 8'b00111111; // 7014 :  63 - 0x3f
      13'h1B67: dout <= 8'b00000000; // 7015 :   0 - 0x0
      13'h1B68: dout <= 8'b01111111; // 7016 : 127 - 0x7f
      13'h1B69: dout <= 8'b01111111; // 7017 : 127 - 0x7f
      13'h1B6A: dout <= 8'b01111111; // 7018 : 127 - 0x7f
      13'h1B6B: dout <= 8'b01111111; // 7019 : 127 - 0x7f
      13'h1B6C: dout <= 8'b01000000; // 7020 :  64 - 0x40
      13'h1B6D: dout <= 8'b00000000; // 7021 :   0 - 0x0
      13'h1B6E: dout <= 8'b00000000; // 7022 :   0 - 0x0
      13'h1B6F: dout <= 8'b00000000; // 7023 :   0 - 0x0
      13'h1B70: dout <= 8'b00000110; // 7024 :   6 - 0x6 -- Background 0xb7
      13'h1B71: dout <= 8'b00000110; // 7025 :   6 - 0x6
      13'h1B72: dout <= 8'b00000110; // 7026 :   6 - 0x6
      13'h1B73: dout <= 8'b00000110; // 7027 :   6 - 0x6
      13'h1B74: dout <= 8'b11111110; // 7028 : 254 - 0xfe
      13'h1B75: dout <= 8'b11111110; // 7029 : 254 - 0xfe
      13'h1B76: dout <= 8'b11111100; // 7030 : 252 - 0xfc
      13'h1B77: dout <= 8'b00000000; // 7031 :   0 - 0x0
      13'h1B78: dout <= 8'b11111000; // 7032 : 248 - 0xf8
      13'h1B79: dout <= 8'b11111000; // 7033 : 248 - 0xf8
      13'h1B7A: dout <= 8'b11111000; // 7034 : 248 - 0xf8
      13'h1B7B: dout <= 8'b11111000; // 7035 : 248 - 0xf8
      13'h1B7C: dout <= 8'b00000000; // 7036 :   0 - 0x0
      13'h1B7D: dout <= 8'b00000000; // 7037 :   0 - 0x0
      13'h1B7E: dout <= 8'b00000000; // 7038 :   0 - 0x0
      13'h1B7F: dout <= 8'b00000000; // 7039 :   0 - 0x0
      13'h1B80: dout <= 8'b01100000; // 7040 :  96 - 0x60 -- Background 0xb8
      13'h1B81: dout <= 8'b11110000; // 7041 : 240 - 0xf0
      13'h1B82: dout <= 8'b11000011; // 7042 : 195 - 0xc3
      13'h1B83: dout <= 8'b10000111; // 7043 : 135 - 0x87
      13'h1B84: dout <= 8'b00000110; // 7044 :   6 - 0x6
      13'h1B85: dout <= 8'b00000100; // 7045 :   4 - 0x4
      13'h1B86: dout <= 8'b00000100; // 7046 :   4 - 0x4
      13'h1B87: dout <= 8'b00000111; // 7047 :   7 - 0x7
      13'h1B88: dout <= 8'b00000000; // 7048 :   0 - 0x0
      13'h1B89: dout <= 8'b00000000; // 7049 :   0 - 0x0
      13'h1B8A: dout <= 8'b00000011; // 7050 :   3 - 0x3
      13'h1B8B: dout <= 8'b00000111; // 7051 :   7 - 0x7
      13'h1B8C: dout <= 8'b00000111; // 7052 :   7 - 0x7
      13'h1B8D: dout <= 8'b00000111; // 7053 :   7 - 0x7
      13'h1B8E: dout <= 8'b00000011; // 7054 :   3 - 0x3
      13'h1B8F: dout <= 8'b00000000; // 7055 :   0 - 0x0
      13'h1B90: dout <= 8'b00000110; // 7056 :   6 - 0x6 -- Background 0xb9
      13'h1B91: dout <= 8'b00001111; // 7057 :  15 - 0xf
      13'h1B92: dout <= 8'b10000111; // 7058 : 135 - 0x87
      13'h1B93: dout <= 8'b11000001; // 7059 : 193 - 0xc1
      13'h1B94: dout <= 8'b00100011; // 7060 :  35 - 0x23
      13'h1B95: dout <= 8'b00101110; // 7061 :  46 - 0x2e
      13'h1B96: dout <= 8'b01100000; // 7062 :  96 - 0x60
      13'h1B97: dout <= 8'b11100001; // 7063 : 225 - 0xe1
      13'h1B98: dout <= 8'b00000000; // 7064 :   0 - 0x0
      13'h1B99: dout <= 8'b00000000; // 7065 :   0 - 0x0
      13'h1B9A: dout <= 8'b11000001; // 7066 : 193 - 0xc1
      13'h1B9B: dout <= 8'b11100010; // 7067 : 226 - 0xe2
      13'h1B9C: dout <= 8'b11001100; // 7068 : 204 - 0xcc
      13'h1B9D: dout <= 8'b11000000; // 7069 : 192 - 0xc0
      13'h1B9E: dout <= 8'b10000000; // 7070 : 128 - 0x80
      13'h1B9F: dout <= 8'b00000001; // 7071 :   1 - 0x1
      13'h1BA0: dout <= 8'b00000000; // 7072 :   0 - 0x0 -- Background 0xba
      13'h1BA1: dout <= 8'b11001000; // 7073 : 200 - 0xc8
      13'h1BA2: dout <= 8'b11111000; // 7074 : 248 - 0xf8
      13'h1BA3: dout <= 8'b10110000; // 7075 : 176 - 0xb0
      13'h1BA4: dout <= 8'b00010000; // 7076 :  16 - 0x10
      13'h1BA5: dout <= 8'b00110000; // 7077 :  48 - 0x30
      13'h1BA6: dout <= 8'b11001000; // 7078 : 200 - 0xc8
      13'h1BA7: dout <= 8'b11111000; // 7079 : 248 - 0xf8
      13'h1BA8: dout <= 8'b00000000; // 7080 :   0 - 0x0
      13'h1BA9: dout <= 8'b11110000; // 7081 : 240 - 0xf0
      13'h1BAA: dout <= 8'b00000000; // 7082 :   0 - 0x0
      13'h1BAB: dout <= 8'b00100000; // 7083 :  32 - 0x20
      13'h1BAC: dout <= 8'b00100000; // 7084 :  32 - 0x20
      13'h1BAD: dout <= 8'b00000000; // 7085 :   0 - 0x0
      13'h1BAE: dout <= 8'b11110000; // 7086 : 240 - 0xf0
      13'h1BAF: dout <= 8'b00000000; // 7087 :   0 - 0x0
      13'h1BB0: dout <= 8'b00000111; // 7088 :   7 - 0x7 -- Background 0xbb
      13'h1BB1: dout <= 8'b00000011; // 7089 :   3 - 0x3
      13'h1BB2: dout <= 8'b00000000; // 7090 :   0 - 0x0
      13'h1BB3: dout <= 8'b01100000; // 7091 :  96 - 0x60
      13'h1BB4: dout <= 8'b11110000; // 7092 : 240 - 0xf0
      13'h1BB5: dout <= 8'b11010000; // 7093 : 208 - 0xd0
      13'h1BB6: dout <= 8'b10010000; // 7094 : 144 - 0x90
      13'h1BB7: dout <= 8'b01100000; // 7095 :  96 - 0x60
      13'h1BB8: dout <= 8'b00000000; // 7096 :   0 - 0x0
      13'h1BB9: dout <= 8'b00000000; // 7097 :   0 - 0x0
      13'h1BBA: dout <= 8'b00000000; // 7098 :   0 - 0x0
      13'h1BBB: dout <= 8'b00000000; // 7099 :   0 - 0x0
      13'h1BBC: dout <= 8'b00000000; // 7100 :   0 - 0x0
      13'h1BBD: dout <= 8'b01100000; // 7101 :  96 - 0x60
      13'h1BBE: dout <= 8'b01100000; // 7102 :  96 - 0x60
      13'h1BBF: dout <= 8'b00000000; // 7103 :   0 - 0x0
      13'h1BC0: dout <= 8'b11100001; // 7104 : 225 - 0xe1 -- Background 0xbc
      13'h1BC1: dout <= 8'b11000011; // 7105 : 195 - 0xc3
      13'h1BC2: dout <= 8'b00001110; // 7106 :  14 - 0xe
      13'h1BC3: dout <= 8'b00000110; // 7107 :   6 - 0x6
      13'h1BC4: dout <= 8'b00001111; // 7108 :  15 - 0xf
      13'h1BC5: dout <= 8'b00001101; // 7109 :  13 - 0xd
      13'h1BC6: dout <= 8'b00001001; // 7110 :   9 - 0x9
      13'h1BC7: dout <= 8'b00000110; // 7111 :   6 - 0x6
      13'h1BC8: dout <= 8'b00000010; // 7112 :   2 - 0x2
      13'h1BC9: dout <= 8'b00001100; // 7113 :  12 - 0xc
      13'h1BCA: dout <= 8'b00000000; // 7114 :   0 - 0x0
      13'h1BCB: dout <= 8'b00000000; // 7115 :   0 - 0x0
      13'h1BCC: dout <= 8'b00000000; // 7116 :   0 - 0x0
      13'h1BCD: dout <= 8'b00000110; // 7117 :   6 - 0x6
      13'h1BCE: dout <= 8'b00000110; // 7118 :   6 - 0x6
      13'h1BCF: dout <= 8'b00000000; // 7119 :   0 - 0x0
      13'h1BD0: dout <= 8'b11100000; // 7120 : 224 - 0xe0 -- Background 0xbd
      13'h1BD1: dout <= 8'b01100000; // 7121 :  96 - 0x60
      13'h1BD2: dout <= 8'b11100011; // 7122 : 227 - 0xe3
      13'h1BD3: dout <= 8'b11100111; // 7123 : 231 - 0xe7
      13'h1BD4: dout <= 8'b00000110; // 7124 :   6 - 0x6
      13'h1BD5: dout <= 8'b00000100; // 7125 :   4 - 0x4
      13'h1BD6: dout <= 8'b00000100; // 7126 :   4 - 0x4
      13'h1BD7: dout <= 8'b00000111; // 7127 :   7 - 0x7
      13'h1BD8: dout <= 8'b00000000; // 7128 :   0 - 0x0
      13'h1BD9: dout <= 8'b10000000; // 7129 : 128 - 0x80
      13'h1BDA: dout <= 8'b00000011; // 7130 :   3 - 0x3
      13'h1BDB: dout <= 8'b00000111; // 7131 :   7 - 0x7
      13'h1BDC: dout <= 8'b00000111; // 7132 :   7 - 0x7
      13'h1BDD: dout <= 8'b00000111; // 7133 :   7 - 0x7
      13'h1BDE: dout <= 8'b00000011; // 7134 :   3 - 0x3
      13'h1BDF: dout <= 8'b00000000; // 7135 :   0 - 0x0
      13'h1BE0: dout <= 8'b00000111; // 7136 :   7 - 0x7 -- Background 0xbe
      13'h1BE1: dout <= 8'b00000011; // 7137 :   3 - 0x3
      13'h1BE2: dout <= 8'b10000111; // 7138 : 135 - 0x87
      13'h1BE3: dout <= 8'b11000111; // 7139 : 199 - 0xc7
      13'h1BE4: dout <= 8'b00100000; // 7140 :  32 - 0x20
      13'h1BE5: dout <= 8'b00100000; // 7141 :  32 - 0x20
      13'h1BE6: dout <= 8'b01100000; // 7142 :  96 - 0x60
      13'h1BE7: dout <= 8'b11100000; // 7143 : 224 - 0xe0
      13'h1BE8: dout <= 8'b00000000; // 7144 :   0 - 0x0
      13'h1BE9: dout <= 8'b00000100; // 7145 :   4 - 0x4
      13'h1BEA: dout <= 8'b11000000; // 7146 : 192 - 0xc0
      13'h1BEB: dout <= 8'b11100000; // 7147 : 224 - 0xe0
      13'h1BEC: dout <= 8'b11000000; // 7148 : 192 - 0xc0
      13'h1BED: dout <= 8'b11000000; // 7149 : 192 - 0xc0
      13'h1BEE: dout <= 8'b10000000; // 7150 : 128 - 0x80
      13'h1BEF: dout <= 8'b00000000; // 7151 :   0 - 0x0
      13'h1BF0: dout <= 8'b00000111; // 7152 :   7 - 0x7 -- Background 0xbf
      13'h1BF1: dout <= 8'b00000011; // 7153 :   3 - 0x3
      13'h1BF2: dout <= 8'b00000000; // 7154 :   0 - 0x0
      13'h1BF3: dout <= 8'b00001100; // 7155 :  12 - 0xc
      13'h1BF4: dout <= 8'b11101100; // 7156 : 236 - 0xec
      13'h1BF5: dout <= 8'b01100100; // 7157 : 100 - 0x64
      13'h1BF6: dout <= 8'b11101100; // 7158 : 236 - 0xec
      13'h1BF7: dout <= 8'b11101101; // 7159 : 237 - 0xed
      13'h1BF8: dout <= 8'b00000000; // 7160 :   0 - 0x0
      13'h1BF9: dout <= 8'b00000000; // 7161 :   0 - 0x0
      13'h1BFA: dout <= 8'b00000000; // 7162 :   0 - 0x0
      13'h1BFB: dout <= 8'b00000000; // 7163 :   0 - 0x0
      13'h1BFC: dout <= 8'b00000000; // 7164 :   0 - 0x0
      13'h1BFD: dout <= 8'b10001000; // 7165 : 136 - 0x88
      13'h1BFE: dout <= 8'b00001000; // 7166 :   8 - 0x8
      13'h1BFF: dout <= 8'b00001011; // 7167 :  11 - 0xb
      13'h1C00: dout <= 8'b11100000; // 7168 : 224 - 0xe0 -- Background 0xc0
      13'h1C01: dout <= 8'b11000000; // 7169 : 192 - 0xc0
      13'h1C02: dout <= 8'b00000000; // 7170 :   0 - 0x0
      13'h1C03: dout <= 8'b00110000; // 7171 :  48 - 0x30
      13'h1C04: dout <= 8'b00110111; // 7172 :  55 - 0x37
      13'h1C05: dout <= 8'b00010011; // 7173 :  19 - 0x13
      13'h1C06: dout <= 8'b00110111; // 7174 :  55 - 0x37
      13'h1C07: dout <= 8'b01110111; // 7175 : 119 - 0x77
      13'h1C08: dout <= 8'b00000000; // 7176 :   0 - 0x0
      13'h1C09: dout <= 8'b00000000; // 7177 :   0 - 0x0
      13'h1C0A: dout <= 8'b00000000; // 7178 :   0 - 0x0
      13'h1C0B: dout <= 8'b00000000; // 7179 :   0 - 0x0
      13'h1C0C: dout <= 8'b00000000; // 7180 :   0 - 0x0
      13'h1C0D: dout <= 8'b00100100; // 7181 :  36 - 0x24
      13'h1C0E: dout <= 8'b00100000; // 7182 :  32 - 0x20
      13'h1C0F: dout <= 8'b10100000; // 7183 : 160 - 0xa0
      13'h1C10: dout <= 8'b00001111; // 7184 :  15 - 0xf -- Background 0xc1
      13'h1C11: dout <= 8'b00001100; // 7185 :  12 - 0xc
      13'h1C12: dout <= 8'b00000000; // 7186 :   0 - 0x0
      13'h1C13: dout <= 8'b00000000; // 7187 :   0 - 0x0
      13'h1C14: dout <= 8'b00000000; // 7188 :   0 - 0x0
      13'h1C15: dout <= 8'b00000000; // 7189 :   0 - 0x0
      13'h1C16: dout <= 8'b00000000; // 7190 :   0 - 0x0
      13'h1C17: dout <= 8'b00000000; // 7191 :   0 - 0x0
      13'h1C18: dout <= 8'b00000000; // 7192 :   0 - 0x0
      13'h1C19: dout <= 8'b00000000; // 7193 :   0 - 0x0
      13'h1C1A: dout <= 8'b00000000; // 7194 :   0 - 0x0
      13'h1C1B: dout <= 8'b00000000; // 7195 :   0 - 0x0
      13'h1C1C: dout <= 8'b00000000; // 7196 :   0 - 0x0
      13'h1C1D: dout <= 8'b00000000; // 7197 :   0 - 0x0
      13'h1C1E: dout <= 8'b00000000; // 7198 :   0 - 0x0
      13'h1C1F: dout <= 8'b00000000; // 7199 :   0 - 0x0
      13'h1C20: dout <= 8'b11110000; // 7200 : 240 - 0xf0 -- Background 0xc2
      13'h1C21: dout <= 8'b00110000; // 7201 :  48 - 0x30
      13'h1C22: dout <= 8'b00000000; // 7202 :   0 - 0x0
      13'h1C23: dout <= 8'b00000000; // 7203 :   0 - 0x0
      13'h1C24: dout <= 8'b00000000; // 7204 :   0 - 0x0
      13'h1C25: dout <= 8'b00000000; // 7205 :   0 - 0x0
      13'h1C26: dout <= 8'b00000000; // 7206 :   0 - 0x0
      13'h1C27: dout <= 8'b00000000; // 7207 :   0 - 0x0
      13'h1C28: dout <= 8'b00000000; // 7208 :   0 - 0x0
      13'h1C29: dout <= 8'b00000000; // 7209 :   0 - 0x0
      13'h1C2A: dout <= 8'b00000000; // 7210 :   0 - 0x0
      13'h1C2B: dout <= 8'b00000000; // 7211 :   0 - 0x0
      13'h1C2C: dout <= 8'b00000000; // 7212 :   0 - 0x0
      13'h1C2D: dout <= 8'b00000000; // 7213 :   0 - 0x0
      13'h1C2E: dout <= 8'b00000000; // 7214 :   0 - 0x0
      13'h1C2F: dout <= 8'b00000000; // 7215 :   0 - 0x0
      13'h1C30: dout <= 8'b00000000; // 7216 :   0 - 0x0 -- Background 0xc3
      13'h1C31: dout <= 8'b00000000; // 7217 :   0 - 0x0
      13'h1C32: dout <= 8'b00000000; // 7218 :   0 - 0x0
      13'h1C33: dout <= 8'b00000100; // 7219 :   4 - 0x4
      13'h1C34: dout <= 8'b00001101; // 7220 :  13 - 0xd
      13'h1C35: dout <= 8'b00001111; // 7221 :  15 - 0xf
      13'h1C36: dout <= 8'b00001100; // 7222 :  12 - 0xc
      13'h1C37: dout <= 8'b00001100; // 7223 :  12 - 0xc
      13'h1C38: dout <= 8'b00000000; // 7224 :   0 - 0x0
      13'h1C39: dout <= 8'b00000000; // 7225 :   0 - 0x0
      13'h1C3A: dout <= 8'b00000000; // 7226 :   0 - 0x0
      13'h1C3B: dout <= 8'b00001000; // 7227 :   8 - 0x8
      13'h1C3C: dout <= 8'b00001011; // 7228 :  11 - 0xb
      13'h1C3D: dout <= 8'b00001000; // 7229 :   8 - 0x8
      13'h1C3E: dout <= 8'b00001000; // 7230 :   8 - 0x8
      13'h1C3F: dout <= 8'b00001000; // 7231 :   8 - 0x8
      13'h1C40: dout <= 8'b00000000; // 7232 :   0 - 0x0 -- Background 0xc4
      13'h1C41: dout <= 8'b00000000; // 7233 :   0 - 0x0
      13'h1C42: dout <= 8'b00000000; // 7234 :   0 - 0x0
      13'h1C43: dout <= 8'b00010000; // 7235 :  16 - 0x10
      13'h1C44: dout <= 8'b01110000; // 7236 : 112 - 0x70
      13'h1C45: dout <= 8'b11110000; // 7237 : 240 - 0xf0
      13'h1C46: dout <= 8'b00110000; // 7238 :  48 - 0x30
      13'h1C47: dout <= 8'b00110000; // 7239 :  48 - 0x30
      13'h1C48: dout <= 8'b00000000; // 7240 :   0 - 0x0
      13'h1C49: dout <= 8'b00000000; // 7241 :   0 - 0x0
      13'h1C4A: dout <= 8'b00000000; // 7242 :   0 - 0x0
      13'h1C4B: dout <= 8'b00100000; // 7243 :  32 - 0x20
      13'h1C4C: dout <= 8'b10100000; // 7244 : 160 - 0xa0
      13'h1C4D: dout <= 8'b00100000; // 7245 :  32 - 0x20
      13'h1C4E: dout <= 8'b00100000; // 7246 :  32 - 0x20
      13'h1C4F: dout <= 8'b00100000; // 7247 :  32 - 0x20
      13'h1C50: dout <= 8'b11100100; // 7248 : 228 - 0xe4 -- Background 0xc5
      13'h1C51: dout <= 8'b00100100; // 7249 :  36 - 0x24
      13'h1C52: dout <= 8'b11100100; // 7250 : 228 - 0xe4
      13'h1C53: dout <= 8'b11101111; // 7251 : 239 - 0xef
      13'h1C54: dout <= 8'b00000111; // 7252 :   7 - 0x7
      13'h1C55: dout <= 8'b00000110; // 7253 :   6 - 0x6
      13'h1C56: dout <= 8'b00000100; // 7254 :   4 - 0x4
      13'h1C57: dout <= 8'b00000100; // 7255 :   4 - 0x4
      13'h1C58: dout <= 8'b00001000; // 7256 :   8 - 0x8
      13'h1C59: dout <= 8'b11001000; // 7257 : 200 - 0xc8
      13'h1C5A: dout <= 8'b00001000; // 7258 :   8 - 0x8
      13'h1C5B: dout <= 8'b00000011; // 7259 :   3 - 0x3
      13'h1C5C: dout <= 8'b00000111; // 7260 :   7 - 0x7
      13'h1C5D: dout <= 8'b00000111; // 7261 :   7 - 0x7
      13'h1C5E: dout <= 8'b00000111; // 7262 :   7 - 0x7
      13'h1C5F: dout <= 8'b00000011; // 7263 :   3 - 0x3
      13'h1C60: dout <= 8'b00010111; // 7264 :  23 - 0x17 -- Background 0xc6
      13'h1C61: dout <= 8'b00010001; // 7265 :  17 - 0x11
      13'h1C62: dout <= 8'b00010111; // 7266 :  23 - 0x17
      13'h1C63: dout <= 8'b10110111; // 7267 : 183 - 0xb7
      13'h1C64: dout <= 8'b11000000; // 7268 : 192 - 0xc0
      13'h1C65: dout <= 8'b00100000; // 7269 :  32 - 0x20
      13'h1C66: dout <= 8'b00100000; // 7270 :  32 - 0x20
      13'h1C67: dout <= 8'b01100000; // 7271 :  96 - 0x60
      13'h1C68: dout <= 8'b00100000; // 7272 :  32 - 0x20
      13'h1C69: dout <= 8'b00100110; // 7273 :  38 - 0x26
      13'h1C6A: dout <= 8'b00100000; // 7274 :  32 - 0x20
      13'h1C6B: dout <= 8'b11000000; // 7275 : 192 - 0xc0
      13'h1C6C: dout <= 8'b11100000; // 7276 : 224 - 0xe0
      13'h1C6D: dout <= 8'b11000000; // 7277 : 192 - 0xc0
      13'h1C6E: dout <= 8'b11000000; // 7278 : 192 - 0xc0
      13'h1C6F: dout <= 8'b10000000; // 7279 : 128 - 0x80
      13'h1C70: dout <= 8'b00000111; // 7280 :   7 - 0x7 -- Background 0xc7
      13'h1C71: dout <= 8'b00000111; // 7281 :   7 - 0x7
      13'h1C72: dout <= 8'b00000011; // 7282 :   3 - 0x3
      13'h1C73: dout <= 8'b00000000; // 7283 :   0 - 0x0
      13'h1C74: dout <= 8'b11100000; // 7284 : 224 - 0xe0
      13'h1C75: dout <= 8'b00100000; // 7285 :  32 - 0x20
      13'h1C76: dout <= 8'b11100000; // 7286 : 224 - 0xe0
      13'h1C77: dout <= 8'b11100000; // 7287 : 224 - 0xe0
      13'h1C78: dout <= 8'b00000000; // 7288 :   0 - 0x0
      13'h1C79: dout <= 8'b00000000; // 7289 :   0 - 0x0
      13'h1C7A: dout <= 8'b00000000; // 7290 :   0 - 0x0
      13'h1C7B: dout <= 8'b00000000; // 7291 :   0 - 0x0
      13'h1C7C: dout <= 8'b00000000; // 7292 :   0 - 0x0
      13'h1C7D: dout <= 8'b11000000; // 7293 : 192 - 0xc0
      13'h1C7E: dout <= 8'b00000000; // 7294 :   0 - 0x0
      13'h1C7F: dout <= 8'b00000000; // 7295 :   0 - 0x0
      13'h1C80: dout <= 8'b11100000; // 7296 : 224 - 0xe0 -- Background 0xc8
      13'h1C81: dout <= 8'b11100000; // 7297 : 224 - 0xe0
      13'h1C82: dout <= 8'b11000000; // 7298 : 192 - 0xc0
      13'h1C83: dout <= 8'b00000000; // 7299 :   0 - 0x0
      13'h1C84: dout <= 8'b00000111; // 7300 :   7 - 0x7
      13'h1C85: dout <= 8'b00000001; // 7301 :   1 - 0x1
      13'h1C86: dout <= 8'b00000111; // 7302 :   7 - 0x7
      13'h1C87: dout <= 8'b00000111; // 7303 :   7 - 0x7
      13'h1C88: dout <= 8'b00000000; // 7304 :   0 - 0x0
      13'h1C89: dout <= 8'b00000000; // 7305 :   0 - 0x0
      13'h1C8A: dout <= 8'b00000000; // 7306 :   0 - 0x0
      13'h1C8B: dout <= 8'b00000000; // 7307 :   0 - 0x0
      13'h1C8C: dout <= 8'b00000000; // 7308 :   0 - 0x0
      13'h1C8D: dout <= 8'b00000110; // 7309 :   6 - 0x6
      13'h1C8E: dout <= 8'b00000000; // 7310 :   0 - 0x0
      13'h1C8F: dout <= 8'b00000000; // 7311 :   0 - 0x0
      13'h1C90: dout <= 8'b00000001; // 7312 :   1 - 0x1 -- Background 0xc9
      13'h1C91: dout <= 8'b00010011; // 7313 :  19 - 0x13
      13'h1C92: dout <= 8'b00011111; // 7314 :  31 - 0x1f
      13'h1C93: dout <= 8'b00001101; // 7315 :  13 - 0xd
      13'h1C94: dout <= 8'b00000100; // 7316 :   4 - 0x4
      13'h1C95: dout <= 8'b00001100; // 7317 :  12 - 0xc
      13'h1C96: dout <= 8'b00010011; // 7318 :  19 - 0x13
      13'h1C97: dout <= 8'b00011111; // 7319 :  31 - 0x1f
      13'h1C98: dout <= 8'b00000000; // 7320 :   0 - 0x0
      13'h1C99: dout <= 8'b00001111; // 7321 :  15 - 0xf
      13'h1C9A: dout <= 8'b00000000; // 7322 :   0 - 0x0
      13'h1C9B: dout <= 8'b00001000; // 7323 :   8 - 0x8
      13'h1C9C: dout <= 8'b00001000; // 7324 :   8 - 0x8
      13'h1C9D: dout <= 8'b00000000; // 7325 :   0 - 0x0
      13'h1C9E: dout <= 8'b00001111; // 7326 :  15 - 0xf
      13'h1C9F: dout <= 8'b00000000; // 7327 :   0 - 0x0
      13'h1CA0: dout <= 8'b01100000; // 7328 :  96 - 0x60 -- Background 0xca
      13'h1CA1: dout <= 8'b01110000; // 7329 : 112 - 0x70
      13'h1CA2: dout <= 8'b10100011; // 7330 : 163 - 0xa3
      13'h1CA3: dout <= 8'b10000111; // 7331 : 135 - 0x87
      13'h1CA4: dout <= 8'b11000110; // 7332 : 198 - 0xc6
      13'h1CA5: dout <= 8'b01110100; // 7333 : 116 - 0x74
      13'h1CA6: dout <= 8'b00000100; // 7334 :   4 - 0x4
      13'h1CA7: dout <= 8'b10000111; // 7335 : 135 - 0x87
      13'h1CA8: dout <= 8'b00000000; // 7336 :   0 - 0x0
      13'h1CA9: dout <= 8'b00000000; // 7337 :   0 - 0x0
      13'h1CAA: dout <= 8'b10000011; // 7338 : 131 - 0x83
      13'h1CAB: dout <= 8'b01000111; // 7339 :  71 - 0x47
      13'h1CAC: dout <= 8'b00110111; // 7340 :  55 - 0x37
      13'h1CAD: dout <= 8'b00000111; // 7341 :   7 - 0x7
      13'h1CAE: dout <= 8'b00000011; // 7342 :   3 - 0x3
      13'h1CAF: dout <= 8'b10000000; // 7343 : 128 - 0x80
      13'h1CB0: dout <= 8'b00000110; // 7344 :   6 - 0x6 -- Background 0xcb
      13'h1CB1: dout <= 8'b00001111; // 7345 :  15 - 0xf
      13'h1CB2: dout <= 8'b10000011; // 7346 : 131 - 0x83
      13'h1CB3: dout <= 8'b11000001; // 7347 : 193 - 0xc1
      13'h1CB4: dout <= 8'b00100000; // 7348 :  32 - 0x20
      13'h1CB5: dout <= 8'b00100000; // 7349 :  32 - 0x20
      13'h1CB6: dout <= 8'b01100000; // 7350 :  96 - 0x60
      13'h1CB7: dout <= 8'b11100000; // 7351 : 224 - 0xe0
      13'h1CB8: dout <= 8'b00000000; // 7352 :   0 - 0x0
      13'h1CB9: dout <= 8'b00000000; // 7353 :   0 - 0x0
      13'h1CBA: dout <= 8'b11000000; // 7354 : 192 - 0xc0
      13'h1CBB: dout <= 8'b11100000; // 7355 : 224 - 0xe0
      13'h1CBC: dout <= 8'b11000000; // 7356 : 192 - 0xc0
      13'h1CBD: dout <= 8'b11000000; // 7357 : 192 - 0xc0
      13'h1CBE: dout <= 8'b10000000; // 7358 : 128 - 0x80
      13'h1CBF: dout <= 8'b00000000; // 7359 :   0 - 0x0
      13'h1CC0: dout <= 8'b10000111; // 7360 : 135 - 0x87 -- Background 0xcc
      13'h1CC1: dout <= 8'b01000011; // 7361 :  67 - 0x43
      13'h1CC2: dout <= 8'b00110000; // 7362 :  48 - 0x30
      13'h1CC3: dout <= 8'b01100000; // 7363 :  96 - 0x60
      13'h1CC4: dout <= 8'b11110000; // 7364 : 240 - 0xf0
      13'h1CC5: dout <= 8'b11010000; // 7365 : 208 - 0xd0
      13'h1CC6: dout <= 8'b10010000; // 7366 : 144 - 0x90
      13'h1CC7: dout <= 8'b01100000; // 7367 :  96 - 0x60
      13'h1CC8: dout <= 8'b01000000; // 7368 :  64 - 0x40
      13'h1CC9: dout <= 8'b00110000; // 7369 :  48 - 0x30
      13'h1CCA: dout <= 8'b00000000; // 7370 :   0 - 0x0
      13'h1CCB: dout <= 8'b00000000; // 7371 :   0 - 0x0
      13'h1CCC: dout <= 8'b00000000; // 7372 :   0 - 0x0
      13'h1CCD: dout <= 8'b01100000; // 7373 :  96 - 0x60
      13'h1CCE: dout <= 8'b01100000; // 7374 :  96 - 0x60
      13'h1CCF: dout <= 8'b00000000; // 7375 :   0 - 0x0
      13'h1CD0: dout <= 8'b11100000; // 7376 : 224 - 0xe0 -- Background 0xcd
      13'h1CD1: dout <= 8'b11000000; // 7377 : 192 - 0xc0
      13'h1CD2: dout <= 8'b00000000; // 7378 :   0 - 0x0
      13'h1CD3: dout <= 8'b00000110; // 7379 :   6 - 0x6
      13'h1CD4: dout <= 8'b00001111; // 7380 :  15 - 0xf
      13'h1CD5: dout <= 8'b00001101; // 7381 :  13 - 0xd
      13'h1CD6: dout <= 8'b00001001; // 7382 :   9 - 0x9
      13'h1CD7: dout <= 8'b00000110; // 7383 :   6 - 0x6
      13'h1CD8: dout <= 8'b00000000; // 7384 :   0 - 0x0
      13'h1CD9: dout <= 8'b00000000; // 7385 :   0 - 0x0
      13'h1CDA: dout <= 8'b00000000; // 7386 :   0 - 0x0
      13'h1CDB: dout <= 8'b00000000; // 7387 :   0 - 0x0
      13'h1CDC: dout <= 8'b00000000; // 7388 :   0 - 0x0
      13'h1CDD: dout <= 8'b00000110; // 7389 :   6 - 0x6
      13'h1CDE: dout <= 8'b00000110; // 7390 :   6 - 0x6
      13'h1CDF: dout <= 8'b00000000; // 7391 :   0 - 0x0
      13'h1CE0: dout <= 8'b11111100; // 7392 : 252 - 0xfc -- Background 0xce
      13'h1CE1: dout <= 8'b11000000; // 7393 : 192 - 0xc0
      13'h1CE2: dout <= 8'b11010001; // 7394 : 209 - 0xd1
      13'h1CE3: dout <= 8'b11000010; // 7395 : 194 - 0xc2
      13'h1CE4: dout <= 8'b10011110; // 7396 : 158 - 0x9e
      13'h1CE5: dout <= 8'b10111111; // 7397 : 191 - 0xbf
      13'h1CE6: dout <= 8'b10110000; // 7398 : 176 - 0xb0
      13'h1CE7: dout <= 8'b10110011; // 7399 : 179 - 0xb3
      13'h1CE8: dout <= 8'b00000000; // 7400 :   0 - 0x0
      13'h1CE9: dout <= 8'b00000001; // 7401 :   1 - 0x1
      13'h1CEA: dout <= 8'b00011011; // 7402 :  27 - 0x1b
      13'h1CEB: dout <= 8'b00010011; // 7403 :  19 - 0x13
      13'h1CEC: dout <= 8'b00011111; // 7404 :  31 - 0x1f
      13'h1CED: dout <= 8'b00111111; // 7405 :  63 - 0x3f
      13'h1CEE: dout <= 8'b00111111; // 7406 :  63 - 0x3f
      13'h1CEF: dout <= 8'b00111111; // 7407 :  63 - 0x3f
      13'h1CF0: dout <= 8'b00000111; // 7408 :   7 - 0x7 -- Background 0xcf
      13'h1CF1: dout <= 8'b11110011; // 7409 : 243 - 0xf3
      13'h1CF2: dout <= 8'b00001011; // 7410 :  11 - 0xb
      13'h1CF3: dout <= 8'b01111011; // 7411 : 123 - 0x7b
      13'h1CF4: dout <= 8'b01111011; // 7412 : 123 - 0x7b
      13'h1CF5: dout <= 8'b11111001; // 7413 : 249 - 0xf9
      13'h1CF6: dout <= 8'b00001101; // 7414 :  13 - 0xd
      13'h1CF7: dout <= 8'b11101101; // 7415 : 237 - 0xed
      13'h1CF8: dout <= 8'b00000000; // 7416 :   0 - 0x0
      13'h1CF9: dout <= 8'b11111000; // 7417 : 248 - 0xf8
      13'h1CFA: dout <= 8'b00001000; // 7418 :   8 - 0x8
      13'h1CFB: dout <= 8'b00001000; // 7419 :   8 - 0x8
      13'h1CFC: dout <= 8'b00001000; // 7420 :   8 - 0x8
      13'h1CFD: dout <= 8'b11111000; // 7421 : 248 - 0xf8
      13'h1CFE: dout <= 8'b11110000; // 7422 : 240 - 0xf0
      13'h1CFF: dout <= 8'b11010000; // 7423 : 208 - 0xd0
      13'h1D00: dout <= 8'b11111111; // 7424 : 255 - 0xff -- Background 0xd0
      13'h1D01: dout <= 8'b11111111; // 7425 : 255 - 0xff
      13'h1D02: dout <= 8'b11111111; // 7426 : 255 - 0xff
      13'h1D03: dout <= 8'b11111111; // 7427 : 255 - 0xff
      13'h1D04: dout <= 8'b11101110; // 7428 : 238 - 0xee
      13'h1D05: dout <= 8'b11101110; // 7429 : 238 - 0xee
      13'h1D06: dout <= 8'b11101110; // 7430 : 238 - 0xee
      13'h1D07: dout <= 8'b11101110; // 7431 : 238 - 0xee
      13'h1D08: dout <= 8'b00000000; // 7432 :   0 - 0x0
      13'h1D09: dout <= 8'b00000000; // 7433 :   0 - 0x0
      13'h1D0A: dout <= 8'b01111100; // 7434 : 124 - 0x7c
      13'h1D0B: dout <= 8'b11111110; // 7435 : 254 - 0xfe
      13'h1D0C: dout <= 8'b11101110; // 7436 : 238 - 0xee
      13'h1D0D: dout <= 8'b11101110; // 7437 : 238 - 0xee
      13'h1D0E: dout <= 8'b11101110; // 7438 : 238 - 0xee
      13'h1D0F: dout <= 8'b11101110; // 7439 : 238 - 0xee
      13'h1D10: dout <= 8'b11111111; // 7440 : 255 - 0xff -- Background 0xd1
      13'h1D11: dout <= 8'b11111111; // 7441 : 255 - 0xff
      13'h1D12: dout <= 8'b11111111; // 7442 : 255 - 0xff
      13'h1D13: dout <= 8'b11111011; // 7443 : 251 - 0xfb
      13'h1D14: dout <= 8'b11111011; // 7444 : 251 - 0xfb
      13'h1D15: dout <= 8'b11111011; // 7445 : 251 - 0xfb
      13'h1D16: dout <= 8'b11111011; // 7446 : 251 - 0xfb
      13'h1D17: dout <= 8'b11111011; // 7447 : 251 - 0xfb
      13'h1D18: dout <= 8'b00000000; // 7448 :   0 - 0x0
      13'h1D19: dout <= 8'b00000000; // 7449 :   0 - 0x0
      13'h1D1A: dout <= 8'b00111000; // 7450 :  56 - 0x38
      13'h1D1B: dout <= 8'b01111000; // 7451 : 120 - 0x78
      13'h1D1C: dout <= 8'b01111000; // 7452 : 120 - 0x78
      13'h1D1D: dout <= 8'b00111000; // 7453 :  56 - 0x38
      13'h1D1E: dout <= 8'b00111000; // 7454 :  56 - 0x38
      13'h1D1F: dout <= 8'b00111000; // 7455 :  56 - 0x38
      13'h1D20: dout <= 8'b11111111; // 7456 : 255 - 0xff -- Background 0xd2
      13'h1D21: dout <= 8'b11111111; // 7457 : 255 - 0xff
      13'h1D22: dout <= 8'b11111111; // 7458 : 255 - 0xff
      13'h1D23: dout <= 8'b11111111; // 7459 : 255 - 0xff
      13'h1D24: dout <= 8'b11101110; // 7460 : 238 - 0xee
      13'h1D25: dout <= 8'b10001110; // 7461 : 142 - 0x8e
      13'h1D26: dout <= 8'b11111110; // 7462 : 254 - 0xfe
      13'h1D27: dout <= 8'b11111110; // 7463 : 254 - 0xfe
      13'h1D28: dout <= 8'b00000000; // 7464 :   0 - 0x0
      13'h1D29: dout <= 8'b00000000; // 7465 :   0 - 0x0
      13'h1D2A: dout <= 8'b01111100; // 7466 : 124 - 0x7c
      13'h1D2B: dout <= 8'b11111110; // 7467 : 254 - 0xfe
      13'h1D2C: dout <= 8'b11101110; // 7468 : 238 - 0xee
      13'h1D2D: dout <= 8'b00001110; // 7469 :  14 - 0xe
      13'h1D2E: dout <= 8'b00001110; // 7470 :  14 - 0xe
      13'h1D2F: dout <= 8'b01111110; // 7471 : 126 - 0x7e
      13'h1D30: dout <= 8'b11111111; // 7472 : 255 - 0xff -- Background 0xd3
      13'h1D31: dout <= 8'b11111111; // 7473 : 255 - 0xff
      13'h1D32: dout <= 8'b11111111; // 7474 : 255 - 0xff
      13'h1D33: dout <= 8'b11111111; // 7475 : 255 - 0xff
      13'h1D34: dout <= 8'b11101110; // 7476 : 238 - 0xee
      13'h1D35: dout <= 8'b10001110; // 7477 : 142 - 0x8e
      13'h1D36: dout <= 8'b11111100; // 7478 : 252 - 0xfc
      13'h1D37: dout <= 8'b11111101; // 7479 : 253 - 0xfd
      13'h1D38: dout <= 8'b00000000; // 7480 :   0 - 0x0
      13'h1D39: dout <= 8'b00000000; // 7481 :   0 - 0x0
      13'h1D3A: dout <= 8'b01111100; // 7482 : 124 - 0x7c
      13'h1D3B: dout <= 8'b11111110; // 7483 : 254 - 0xfe
      13'h1D3C: dout <= 8'b11101110; // 7484 : 238 - 0xee
      13'h1D3D: dout <= 8'b00001110; // 7485 :  14 - 0xe
      13'h1D3E: dout <= 8'b00111100; // 7486 :  60 - 0x3c
      13'h1D3F: dout <= 8'b00111100; // 7487 :  60 - 0x3c
      13'h1D40: dout <= 8'b11111111; // 7488 : 255 - 0xff -- Background 0xd4
      13'h1D41: dout <= 8'b11111111; // 7489 : 255 - 0xff
      13'h1D42: dout <= 8'b11111111; // 7490 : 255 - 0xff
      13'h1D43: dout <= 8'b11111110; // 7491 : 254 - 0xfe
      13'h1D44: dout <= 8'b11101110; // 7492 : 238 - 0xee
      13'h1D45: dout <= 8'b11101110; // 7493 : 238 - 0xee
      13'h1D46: dout <= 8'b11101110; // 7494 : 238 - 0xee
      13'h1D47: dout <= 8'b11101110; // 7495 : 238 - 0xee
      13'h1D48: dout <= 8'b00000000; // 7496 :   0 - 0x0
      13'h1D49: dout <= 8'b00000000; // 7497 :   0 - 0x0
      13'h1D4A: dout <= 8'b00111110; // 7498 :  62 - 0x3e
      13'h1D4B: dout <= 8'b01111110; // 7499 : 126 - 0x7e
      13'h1D4C: dout <= 8'b11101110; // 7500 : 238 - 0xee
      13'h1D4D: dout <= 8'b11101110; // 7501 : 238 - 0xee
      13'h1D4E: dout <= 8'b11101110; // 7502 : 238 - 0xee
      13'h1D4F: dout <= 8'b11101110; // 7503 : 238 - 0xee
      13'h1D50: dout <= 8'b11111111; // 7504 : 255 - 0xff -- Background 0xd5
      13'h1D51: dout <= 8'b11111111; // 7505 : 255 - 0xff
      13'h1D52: dout <= 8'b11111111; // 7506 : 255 - 0xff
      13'h1D53: dout <= 8'b11111101; // 7507 : 253 - 0xfd
      13'h1D54: dout <= 8'b11100001; // 7508 : 225 - 0xe1
      13'h1D55: dout <= 8'b11101111; // 7509 : 239 - 0xef
      13'h1D56: dout <= 8'b11111111; // 7510 : 255 - 0xff
      13'h1D57: dout <= 8'b11111111; // 7511 : 255 - 0xff
      13'h1D58: dout <= 8'b00000000; // 7512 :   0 - 0x0
      13'h1D59: dout <= 8'b00000000; // 7513 :   0 - 0x0
      13'h1D5A: dout <= 8'b11111100; // 7514 : 252 - 0xfc
      13'h1D5B: dout <= 8'b11111100; // 7515 : 252 - 0xfc
      13'h1D5C: dout <= 8'b11100000; // 7516 : 224 - 0xe0
      13'h1D5D: dout <= 8'b11100000; // 7517 : 224 - 0xe0
      13'h1D5E: dout <= 8'b11111100; // 7518 : 252 - 0xfc
      13'h1D5F: dout <= 8'b11111110; // 7519 : 254 - 0xfe
      13'h1D60: dout <= 8'b11111111; // 7520 : 255 - 0xff -- Background 0xd6
      13'h1D61: dout <= 8'b11111111; // 7521 : 255 - 0xff
      13'h1D62: dout <= 8'b11111111; // 7522 : 255 - 0xff
      13'h1D63: dout <= 8'b11111101; // 7523 : 253 - 0xfd
      13'h1D64: dout <= 8'b11100001; // 7524 : 225 - 0xe1
      13'h1D65: dout <= 8'b11101111; // 7525 : 239 - 0xef
      13'h1D66: dout <= 8'b11111111; // 7526 : 255 - 0xff
      13'h1D67: dout <= 8'b11111111; // 7527 : 255 - 0xff
      13'h1D68: dout <= 8'b00000000; // 7528 :   0 - 0x0
      13'h1D69: dout <= 8'b00000000; // 7529 :   0 - 0x0
      13'h1D6A: dout <= 8'b01111100; // 7530 : 124 - 0x7c
      13'h1D6B: dout <= 8'b11111100; // 7531 : 252 - 0xfc
      13'h1D6C: dout <= 8'b11100000; // 7532 : 224 - 0xe0
      13'h1D6D: dout <= 8'b11100000; // 7533 : 224 - 0xe0
      13'h1D6E: dout <= 8'b11111100; // 7534 : 252 - 0xfc
      13'h1D6F: dout <= 8'b11111110; // 7535 : 254 - 0xfe
      13'h1D70: dout <= 8'b11111111; // 7536 : 255 - 0xff -- Background 0xd7
      13'h1D71: dout <= 8'b11111111; // 7537 : 255 - 0xff
      13'h1D72: dout <= 8'b11111111; // 7538 : 255 - 0xff
      13'h1D73: dout <= 8'b11111110; // 7539 : 254 - 0xfe
      13'h1D74: dout <= 8'b11101110; // 7540 : 238 - 0xee
      13'h1D75: dout <= 8'b10001110; // 7541 : 142 - 0x8e
      13'h1D76: dout <= 8'b11111110; // 7542 : 254 - 0xfe
      13'h1D77: dout <= 8'b11111100; // 7543 : 252 - 0xfc
      13'h1D78: dout <= 8'b00000000; // 7544 :   0 - 0x0
      13'h1D79: dout <= 8'b00000000; // 7545 :   0 - 0x0
      13'h1D7A: dout <= 8'b11111110; // 7546 : 254 - 0xfe
      13'h1D7B: dout <= 8'b11111110; // 7547 : 254 - 0xfe
      13'h1D7C: dout <= 8'b11101110; // 7548 : 238 - 0xee
      13'h1D7D: dout <= 8'b00001110; // 7549 :  14 - 0xe
      13'h1D7E: dout <= 8'b00001110; // 7550 :  14 - 0xe
      13'h1D7F: dout <= 8'b00011100; // 7551 :  28 - 0x1c
      13'h1D80: dout <= 8'b11111111; // 7552 : 255 - 0xff -- Background 0xd8
      13'h1D81: dout <= 8'b11111111; // 7553 : 255 - 0xff
      13'h1D82: dout <= 8'b11111111; // 7554 : 255 - 0xff
      13'h1D83: dout <= 8'b11111111; // 7555 : 255 - 0xff
      13'h1D84: dout <= 8'b11101110; // 7556 : 238 - 0xee
      13'h1D85: dout <= 8'b11101110; // 7557 : 238 - 0xee
      13'h1D86: dout <= 8'b11111100; // 7558 : 252 - 0xfc
      13'h1D87: dout <= 8'b11111111; // 7559 : 255 - 0xff
      13'h1D88: dout <= 8'b00000000; // 7560 :   0 - 0x0
      13'h1D89: dout <= 8'b00000000; // 7561 :   0 - 0x0
      13'h1D8A: dout <= 8'b01111100; // 7562 : 124 - 0x7c
      13'h1D8B: dout <= 8'b11111110; // 7563 : 254 - 0xfe
      13'h1D8C: dout <= 8'b11101110; // 7564 : 238 - 0xee
      13'h1D8D: dout <= 8'b11101110; // 7565 : 238 - 0xee
      13'h1D8E: dout <= 8'b01111100; // 7566 : 124 - 0x7c
      13'h1D8F: dout <= 8'b11111110; // 7567 : 254 - 0xfe
      13'h1D90: dout <= 8'b11111111; // 7568 : 255 - 0xff -- Background 0xd9
      13'h1D91: dout <= 8'b11111111; // 7569 : 255 - 0xff
      13'h1D92: dout <= 8'b11111111; // 7570 : 255 - 0xff
      13'h1D93: dout <= 8'b11111111; // 7571 : 255 - 0xff
      13'h1D94: dout <= 8'b11101110; // 7572 : 238 - 0xee
      13'h1D95: dout <= 8'b11101110; // 7573 : 238 - 0xee
      13'h1D96: dout <= 8'b11101110; // 7574 : 238 - 0xee
      13'h1D97: dout <= 8'b11101110; // 7575 : 238 - 0xee
      13'h1D98: dout <= 8'b00000000; // 7576 :   0 - 0x0
      13'h1D99: dout <= 8'b00000000; // 7577 :   0 - 0x0
      13'h1D9A: dout <= 8'b01111100; // 7578 : 124 - 0x7c
      13'h1D9B: dout <= 8'b11111110; // 7579 : 254 - 0xfe
      13'h1D9C: dout <= 8'b11101110; // 7580 : 238 - 0xee
      13'h1D9D: dout <= 8'b11101110; // 7581 : 238 - 0xee
      13'h1D9E: dout <= 8'b11101110; // 7582 : 238 - 0xee
      13'h1D9F: dout <= 8'b11101110; // 7583 : 238 - 0xee
      13'h1DA0: dout <= 8'b00000000; // 7584 :   0 - 0x0 -- Background 0xda
      13'h1DA1: dout <= 8'b00000000; // 7585 :   0 - 0x0
      13'h1DA2: dout <= 8'b00000000; // 7586 :   0 - 0x0
      13'h1DA3: dout <= 8'b10000000; // 7587 : 128 - 0x80
      13'h1DA4: dout <= 8'b00000000; // 7588 :   0 - 0x0
      13'h1DA5: dout <= 8'b00000000; // 7589 :   0 - 0x0
      13'h1DA6: dout <= 8'b00000100; // 7590 :   4 - 0x4
      13'h1DA7: dout <= 8'b00000000; // 7591 :   0 - 0x0
      13'h1DA8: dout <= 8'b00000000; // 7592 :   0 - 0x0
      13'h1DA9: dout <= 8'b00100000; // 7593 :  32 - 0x20
      13'h1DAA: dout <= 8'b00000000; // 7594 :   0 - 0x0
      13'h1DAB: dout <= 8'b00000010; // 7595 :   2 - 0x2
      13'h1DAC: dout <= 8'b00000000; // 7596 :   0 - 0x0
      13'h1DAD: dout <= 8'b00100000; // 7597 :  32 - 0x20
      13'h1DAE: dout <= 8'b00000000; // 7598 :   0 - 0x0
      13'h1DAF: dout <= 8'b00000000; // 7599 :   0 - 0x0
      13'h1DB0: dout <= 8'b00000000; // 7600 :   0 - 0x0 -- Background 0xdb
      13'h1DB1: dout <= 8'b00000100; // 7601 :   4 - 0x4
      13'h1DB2: dout <= 8'b00000000; // 7602 :   0 - 0x0
      13'h1DB3: dout <= 8'b00010001; // 7603 :  17 - 0x11
      13'h1DB4: dout <= 8'b00000000; // 7604 :   0 - 0x0
      13'h1DB5: dout <= 8'b00000000; // 7605 :   0 - 0x0
      13'h1DB6: dout <= 8'b00000000; // 7606 :   0 - 0x0
      13'h1DB7: dout <= 8'b00100000; // 7607 :  32 - 0x20
      13'h1DB8: dout <= 8'b00100000; // 7608 :  32 - 0x20
      13'h1DB9: dout <= 8'b00000000; // 7609 :   0 - 0x0
      13'h1DBA: dout <= 8'b00000000; // 7610 :   0 - 0x0
      13'h1DBB: dout <= 8'b00000000; // 7611 :   0 - 0x0
      13'h1DBC: dout <= 8'b10000000; // 7612 : 128 - 0x80
      13'h1DBD: dout <= 8'b00000000; // 7613 :   0 - 0x0
      13'h1DBE: dout <= 8'b00000100; // 7614 :   4 - 0x4
      13'h1DBF: dout <= 8'b00000000; // 7615 :   0 - 0x0
      13'h1DC0: dout <= 8'b00000000; // 7616 :   0 - 0x0 -- Background 0xdc
      13'h1DC1: dout <= 8'b00000000; // 7617 :   0 - 0x0
      13'h1DC2: dout <= 8'b00000000; // 7618 :   0 - 0x0
      13'h1DC3: dout <= 8'b00100000; // 7619 :  32 - 0x20
      13'h1DC4: dout <= 8'b00000000; // 7620 :   0 - 0x0
      13'h1DC5: dout <= 8'b00000000; // 7621 :   0 - 0x0
      13'h1DC6: dout <= 8'b00000000; // 7622 :   0 - 0x0
      13'h1DC7: dout <= 8'b00000100; // 7623 :   4 - 0x4
      13'h1DC8: dout <= 8'b00000000; // 7624 :   0 - 0x0
      13'h1DC9: dout <= 8'b00001000; // 7625 :   8 - 0x8
      13'h1DCA: dout <= 8'b00000000; // 7626 :   0 - 0x0
      13'h1DCB: dout <= 8'b00000000; // 7627 :   0 - 0x0
      13'h1DCC: dout <= 8'b00000010; // 7628 :   2 - 0x2
      13'h1DCD: dout <= 8'b00000000; // 7629 :   0 - 0x0
      13'h1DCE: dout <= 8'b01000000; // 7630 :  64 - 0x40
      13'h1DCF: dout <= 8'b00000000; // 7631 :   0 - 0x0
      13'h1DD0: dout <= 8'b00000000; // 7632 :   0 - 0x0 -- Background 0xdd
      13'h1DD1: dout <= 8'b00000000; // 7633 :   0 - 0x0
      13'h1DD2: dout <= 8'b00010001; // 7634 :  17 - 0x11
      13'h1DD3: dout <= 8'b00000000; // 7635 :   0 - 0x0
      13'h1DD4: dout <= 8'b00000000; // 7636 :   0 - 0x0
      13'h1DD5: dout <= 8'b10000000; // 7637 : 128 - 0x80
      13'h1DD6: dout <= 8'b00000000; // 7638 :   0 - 0x0
      13'h1DD7: dout <= 8'b00000000; // 7639 :   0 - 0x0
      13'h1DD8: dout <= 8'b00000000; // 7640 :   0 - 0x0
      13'h1DD9: dout <= 8'b01000000; // 7641 :  64 - 0x40
      13'h1DDA: dout <= 8'b00000000; // 7642 :   0 - 0x0
      13'h1DDB: dout <= 8'b00000000; // 7643 :   0 - 0x0
      13'h1DDC: dout <= 8'b00000000; // 7644 :   0 - 0x0
      13'h1DDD: dout <= 8'b00000000; // 7645 :   0 - 0x0
      13'h1DDE: dout <= 8'b00000010; // 7646 :   2 - 0x2
      13'h1DDF: dout <= 8'b00100000; // 7647 :  32 - 0x20
      13'h1DE0: dout <= 8'b10110011; // 7648 : 179 - 0xb3 -- Background 0xde
      13'h1DE1: dout <= 8'b10110011; // 7649 : 179 - 0xb3
      13'h1DE2: dout <= 8'b10110011; // 7650 : 179 - 0xb3
      13'h1DE3: dout <= 8'b10110011; // 7651 : 179 - 0xb3
      13'h1DE4: dout <= 8'b10110000; // 7652 : 176 - 0xb0
      13'h1DE5: dout <= 8'b10101111; // 7653 : 175 - 0xaf
      13'h1DE6: dout <= 8'b10011111; // 7654 : 159 - 0x9f
      13'h1DE7: dout <= 8'b11000000; // 7655 : 192 - 0xc0
      13'h1DE8: dout <= 8'b00111110; // 7656 :  62 - 0x3e
      13'h1DE9: dout <= 8'b00111111; // 7657 :  63 - 0x3f
      13'h1DEA: dout <= 8'b00111110; // 7658 :  62 - 0x3e
      13'h1DEB: dout <= 8'b00111100; // 7659 :  60 - 0x3c
      13'h1DEC: dout <= 8'b00111111; // 7660 :  63 - 0x3f
      13'h1DED: dout <= 8'b00110000; // 7661 :  48 - 0x30
      13'h1DEE: dout <= 8'b00000000; // 7662 :   0 - 0x0
      13'h1DEF: dout <= 8'b00000000; // 7663 :   0 - 0x0
      13'h1DF0: dout <= 8'b11101101; // 7664 : 237 - 0xed -- Background 0xdf
      13'h1DF1: dout <= 8'b11001101; // 7665 : 205 - 0xcd
      13'h1DF2: dout <= 8'b11001101; // 7666 : 205 - 0xcd
      13'h1DF3: dout <= 8'b00001101; // 7667 :  13 - 0xd
      13'h1DF4: dout <= 8'b00001101; // 7668 :  13 - 0xd
      13'h1DF5: dout <= 8'b11111101; // 7669 : 253 - 0xfd
      13'h1DF6: dout <= 8'b11111101; // 7670 : 253 - 0xfd
      13'h1DF7: dout <= 8'b00000011; // 7671 :   3 - 0x3
      13'h1DF8: dout <= 8'b00010000; // 7672 :  16 - 0x10
      13'h1DF9: dout <= 8'b10110000; // 7673 : 176 - 0xb0
      13'h1DFA: dout <= 8'b00110000; // 7674 :  48 - 0x30
      13'h1DFB: dout <= 8'b11110000; // 7675 : 240 - 0xf0
      13'h1DFC: dout <= 8'b11110000; // 7676 : 240 - 0xf0
      13'h1DFD: dout <= 8'b00000000; // 7677 :   0 - 0x0
      13'h1DFE: dout <= 8'b00000000; // 7678 :   0 - 0x0
      13'h1DFF: dout <= 8'b00000000; // 7679 :   0 - 0x0
      13'h1E00: dout <= 8'b11101110; // 7680 : 238 - 0xee -- Background 0xe0
      13'h1E01: dout <= 8'b11101110; // 7681 : 238 - 0xee
      13'h1E02: dout <= 8'b11101110; // 7682 : 238 - 0xee
      13'h1E03: dout <= 8'b11101110; // 7683 : 238 - 0xee
      13'h1E04: dout <= 8'b11111110; // 7684 : 254 - 0xfe
      13'h1E05: dout <= 8'b11111100; // 7685 : 252 - 0xfc
      13'h1E06: dout <= 8'b11000001; // 7686 : 193 - 0xc1
      13'h1E07: dout <= 8'b11111111; // 7687 : 255 - 0xff
      13'h1E08: dout <= 8'b11101110; // 7688 : 238 - 0xee
      13'h1E09: dout <= 8'b11101110; // 7689 : 238 - 0xee
      13'h1E0A: dout <= 8'b11101110; // 7690 : 238 - 0xee
      13'h1E0B: dout <= 8'b11101110; // 7691 : 238 - 0xee
      13'h1E0C: dout <= 8'b11111110; // 7692 : 254 - 0xfe
      13'h1E0D: dout <= 8'b01111100; // 7693 : 124 - 0x7c
      13'h1E0E: dout <= 8'b00000000; // 7694 :   0 - 0x0
      13'h1E0F: dout <= 8'b00000000; // 7695 :   0 - 0x0
      13'h1E10: dout <= 8'b11111011; // 7696 : 251 - 0xfb -- Background 0xe1
      13'h1E11: dout <= 8'b11111011; // 7697 : 251 - 0xfb
      13'h1E12: dout <= 8'b11111011; // 7698 : 251 - 0xfb
      13'h1E13: dout <= 8'b11111011; // 7699 : 251 - 0xfb
      13'h1E14: dout <= 8'b11111111; // 7700 : 255 - 0xff
      13'h1E15: dout <= 8'b11111101; // 7701 : 253 - 0xfd
      13'h1E16: dout <= 8'b11000001; // 7702 : 193 - 0xc1
      13'h1E17: dout <= 8'b11111111; // 7703 : 255 - 0xff
      13'h1E18: dout <= 8'b00111000; // 7704 :  56 - 0x38
      13'h1E19: dout <= 8'b00111000; // 7705 :  56 - 0x38
      13'h1E1A: dout <= 8'b00111000; // 7706 :  56 - 0x38
      13'h1E1B: dout <= 8'b00111000; // 7707 :  56 - 0x38
      13'h1E1C: dout <= 8'b01111100; // 7708 : 124 - 0x7c
      13'h1E1D: dout <= 8'b01111100; // 7709 : 124 - 0x7c
      13'h1E1E: dout <= 8'b00000000; // 7710 :   0 - 0x0
      13'h1E1F: dout <= 8'b00000000; // 7711 :   0 - 0x0
      13'h1E20: dout <= 8'b11111100; // 7712 : 252 - 0xfc -- Background 0xe2
      13'h1E21: dout <= 8'b11100001; // 7713 : 225 - 0xe1
      13'h1E22: dout <= 8'b11101111; // 7714 : 239 - 0xef
      13'h1E23: dout <= 8'b11101111; // 7715 : 239 - 0xef
      13'h1E24: dout <= 8'b11111111; // 7716 : 255 - 0xff
      13'h1E25: dout <= 8'b11111110; // 7717 : 254 - 0xfe
      13'h1E26: dout <= 8'b10000000; // 7718 : 128 - 0x80
      13'h1E27: dout <= 8'b11111111; // 7719 : 255 - 0xff
      13'h1E28: dout <= 8'b11111100; // 7720 : 252 - 0xfc
      13'h1E29: dout <= 8'b11100000; // 7721 : 224 - 0xe0
      13'h1E2A: dout <= 8'b11100000; // 7722 : 224 - 0xe0
      13'h1E2B: dout <= 8'b11100000; // 7723 : 224 - 0xe0
      13'h1E2C: dout <= 8'b11111110; // 7724 : 254 - 0xfe
      13'h1E2D: dout <= 8'b11111110; // 7725 : 254 - 0xfe
      13'h1E2E: dout <= 8'b00000000; // 7726 :   0 - 0x0
      13'h1E2F: dout <= 8'b00000000; // 7727 :   0 - 0x0
      13'h1E30: dout <= 8'b11101110; // 7728 : 238 - 0xee -- Background 0xe3
      13'h1E31: dout <= 8'b11111110; // 7729 : 254 - 0xfe
      13'h1E32: dout <= 8'b11111110; // 7730 : 254 - 0xfe
      13'h1E33: dout <= 8'b11111110; // 7731 : 254 - 0xfe
      13'h1E34: dout <= 8'b11111110; // 7732 : 254 - 0xfe
      13'h1E35: dout <= 8'b11111100; // 7733 : 252 - 0xfc
      13'h1E36: dout <= 8'b11000001; // 7734 : 193 - 0xc1
      13'h1E37: dout <= 8'b11111111; // 7735 : 255 - 0xff
      13'h1E38: dout <= 8'b00001110; // 7736 :  14 - 0xe
      13'h1E39: dout <= 8'b00001110; // 7737 :  14 - 0xe
      13'h1E3A: dout <= 8'b00001110; // 7738 :  14 - 0xe
      13'h1E3B: dout <= 8'b11101110; // 7739 : 238 - 0xee
      13'h1E3C: dout <= 8'b11111110; // 7740 : 254 - 0xfe
      13'h1E3D: dout <= 8'b01111100; // 7741 : 124 - 0x7c
      13'h1E3E: dout <= 8'b00000000; // 7742 :   0 - 0x0
      13'h1E3F: dout <= 8'b00000000; // 7743 :   0 - 0x0
      13'h1E40: dout <= 8'b11101110; // 7744 : 238 - 0xee -- Background 0xe4
      13'h1E41: dout <= 8'b11101110; // 7745 : 238 - 0xee
      13'h1E42: dout <= 8'b11111110; // 7746 : 254 - 0xfe
      13'h1E43: dout <= 8'b11111110; // 7747 : 254 - 0xfe
      13'h1E44: dout <= 8'b10001110; // 7748 : 142 - 0x8e
      13'h1E45: dout <= 8'b11111110; // 7749 : 254 - 0xfe
      13'h1E46: dout <= 8'b11111000; // 7750 : 248 - 0xf8
      13'h1E47: dout <= 8'b11111111; // 7751 : 255 - 0xff
      13'h1E48: dout <= 8'b11101110; // 7752 : 238 - 0xee
      13'h1E49: dout <= 8'b11101110; // 7753 : 238 - 0xee
      13'h1E4A: dout <= 8'b11111110; // 7754 : 254 - 0xfe
      13'h1E4B: dout <= 8'b11111110; // 7755 : 254 - 0xfe
      13'h1E4C: dout <= 8'b00001110; // 7756 :  14 - 0xe
      13'h1E4D: dout <= 8'b00001110; // 7757 :  14 - 0xe
      13'h1E4E: dout <= 8'b00000000; // 7758 :   0 - 0x0
      13'h1E4F: dout <= 8'b00000000; // 7759 :   0 - 0x0
      13'h1E50: dout <= 8'b10001110; // 7760 : 142 - 0x8e -- Background 0xe5
      13'h1E51: dout <= 8'b11111110; // 7761 : 254 - 0xfe
      13'h1E52: dout <= 8'b11111110; // 7762 : 254 - 0xfe
      13'h1E53: dout <= 8'b11111110; // 7763 : 254 - 0xfe
      13'h1E54: dout <= 8'b11111110; // 7764 : 254 - 0xfe
      13'h1E55: dout <= 8'b11111100; // 7765 : 252 - 0xfc
      13'h1E56: dout <= 8'b11000001; // 7766 : 193 - 0xc1
      13'h1E57: dout <= 8'b11111111; // 7767 : 255 - 0xff
      13'h1E58: dout <= 8'b00001110; // 7768 :  14 - 0xe
      13'h1E59: dout <= 8'b00001110; // 7769 :  14 - 0xe
      13'h1E5A: dout <= 8'b00001110; // 7770 :  14 - 0xe
      13'h1E5B: dout <= 8'b11101110; // 7771 : 238 - 0xee
      13'h1E5C: dout <= 8'b11111110; // 7772 : 254 - 0xfe
      13'h1E5D: dout <= 8'b01111100; // 7773 : 124 - 0x7c
      13'h1E5E: dout <= 8'b00000000; // 7774 :   0 - 0x0
      13'h1E5F: dout <= 8'b00000000; // 7775 :   0 - 0x0
      13'h1E60: dout <= 8'b11101110; // 7776 : 238 - 0xee -- Background 0xe6
      13'h1E61: dout <= 8'b11101110; // 7777 : 238 - 0xee
      13'h1E62: dout <= 8'b11101110; // 7778 : 238 - 0xee
      13'h1E63: dout <= 8'b11101110; // 7779 : 238 - 0xee
      13'h1E64: dout <= 8'b11111110; // 7780 : 254 - 0xfe
      13'h1E65: dout <= 8'b11111100; // 7781 : 252 - 0xfc
      13'h1E66: dout <= 8'b11000001; // 7782 : 193 - 0xc1
      13'h1E67: dout <= 8'b11111111; // 7783 : 255 - 0xff
      13'h1E68: dout <= 8'b11101110; // 7784 : 238 - 0xee
      13'h1E69: dout <= 8'b11101110; // 7785 : 238 - 0xee
      13'h1E6A: dout <= 8'b11101110; // 7786 : 238 - 0xee
      13'h1E6B: dout <= 8'b11101110; // 7787 : 238 - 0xee
      13'h1E6C: dout <= 8'b11111110; // 7788 : 254 - 0xfe
      13'h1E6D: dout <= 8'b01111100; // 7789 : 124 - 0x7c
      13'h1E6E: dout <= 8'b00000000; // 7790 :   0 - 0x0
      13'h1E6F: dout <= 8'b00000000; // 7791 :   0 - 0x0
      13'h1E70: dout <= 8'b11111101; // 7792 : 253 - 0xfd -- Background 0xe7
      13'h1E71: dout <= 8'b11111101; // 7793 : 253 - 0xfd
      13'h1E72: dout <= 8'b11111001; // 7794 : 249 - 0xf9
      13'h1E73: dout <= 8'b11111011; // 7795 : 251 - 0xfb
      13'h1E74: dout <= 8'b11111011; // 7796 : 251 - 0xfb
      13'h1E75: dout <= 8'b11111011; // 7797 : 251 - 0xfb
      13'h1E76: dout <= 8'b11100011; // 7798 : 227 - 0xe3
      13'h1E77: dout <= 8'b11111111; // 7799 : 255 - 0xff
      13'h1E78: dout <= 8'b00011100; // 7800 :  28 - 0x1c
      13'h1E79: dout <= 8'b00011100; // 7801 :  28 - 0x1c
      13'h1E7A: dout <= 8'b00111000; // 7802 :  56 - 0x38
      13'h1E7B: dout <= 8'b00111000; // 7803 :  56 - 0x38
      13'h1E7C: dout <= 8'b00111000; // 7804 :  56 - 0x38
      13'h1E7D: dout <= 8'b00111000; // 7805 :  56 - 0x38
      13'h1E7E: dout <= 8'b00000000; // 7806 :   0 - 0x0
      13'h1E7F: dout <= 8'b00000000; // 7807 :   0 - 0x0
      13'h1E80: dout <= 8'b11101110; // 7808 : 238 - 0xee -- Background 0xe8
      13'h1E81: dout <= 8'b11101110; // 7809 : 238 - 0xee
      13'h1E82: dout <= 8'b11101110; // 7810 : 238 - 0xee
      13'h1E83: dout <= 8'b11101110; // 7811 : 238 - 0xee
      13'h1E84: dout <= 8'b11111110; // 7812 : 254 - 0xfe
      13'h1E85: dout <= 8'b11111100; // 7813 : 252 - 0xfc
      13'h1E86: dout <= 8'b11000001; // 7814 : 193 - 0xc1
      13'h1E87: dout <= 8'b11111111; // 7815 : 255 - 0xff
      13'h1E88: dout <= 8'b11101110; // 7816 : 238 - 0xee
      13'h1E89: dout <= 8'b11101110; // 7817 : 238 - 0xee
      13'h1E8A: dout <= 8'b11101110; // 7818 : 238 - 0xee
      13'h1E8B: dout <= 8'b11101110; // 7819 : 238 - 0xee
      13'h1E8C: dout <= 8'b11111110; // 7820 : 254 - 0xfe
      13'h1E8D: dout <= 8'b01111100; // 7821 : 124 - 0x7c
      13'h1E8E: dout <= 8'b00000000; // 7822 :   0 - 0x0
      13'h1E8F: dout <= 8'b00000000; // 7823 :   0 - 0x0
      13'h1E90: dout <= 8'b11111110; // 7824 : 254 - 0xfe -- Background 0xe9
      13'h1E91: dout <= 8'b11111110; // 7825 : 254 - 0xfe
      13'h1E92: dout <= 8'b11001110; // 7826 : 206 - 0xce
      13'h1E93: dout <= 8'b11111110; // 7827 : 254 - 0xfe
      13'h1E94: dout <= 8'b11111110; // 7828 : 254 - 0xfe
      13'h1E95: dout <= 8'b11111100; // 7829 : 252 - 0xfc
      13'h1E96: dout <= 8'b11000001; // 7830 : 193 - 0xc1
      13'h1E97: dout <= 8'b11111111; // 7831 : 255 - 0xff
      13'h1E98: dout <= 8'b11111110; // 7832 : 254 - 0xfe
      13'h1E99: dout <= 8'b01111110; // 7833 : 126 - 0x7e
      13'h1E9A: dout <= 8'b00001110; // 7834 :  14 - 0xe
      13'h1E9B: dout <= 8'b00001110; // 7835 :  14 - 0xe
      13'h1E9C: dout <= 8'b01111110; // 7836 : 126 - 0x7e
      13'h1E9D: dout <= 8'b01111100; // 7837 : 124 - 0x7c
      13'h1E9E: dout <= 8'b00000000; // 7838 :   0 - 0x0
      13'h1E9F: dout <= 8'b00000000; // 7839 :   0 - 0x0
      13'h1EA0: dout <= 8'b00000000; // 7840 :   0 - 0x0 -- Background 0xea
      13'h1EA1: dout <= 8'b01110000; // 7841 : 112 - 0x70
      13'h1EA2: dout <= 8'b00111000; // 7842 :  56 - 0x38
      13'h1EA3: dout <= 8'b00000000; // 7843 :   0 - 0x0
      13'h1EA4: dout <= 8'b00000010; // 7844 :   2 - 0x2
      13'h1EA5: dout <= 8'b00000111; // 7845 :   7 - 0x7
      13'h1EA6: dout <= 8'b00000011; // 7846 :   3 - 0x3
      13'h1EA7: dout <= 8'b00000000; // 7847 :   0 - 0x0
      13'h1EA8: dout <= 8'b00000000; // 7848 :   0 - 0x0
      13'h1EA9: dout <= 8'b01110000; // 7849 : 112 - 0x70
      13'h1EAA: dout <= 8'b00111000; // 7850 :  56 - 0x38
      13'h1EAB: dout <= 8'b00000000; // 7851 :   0 - 0x0
      13'h1EAC: dout <= 8'b00000010; // 7852 :   2 - 0x2
      13'h1EAD: dout <= 8'b00000111; // 7853 :   7 - 0x7
      13'h1EAE: dout <= 8'b00000011; // 7854 :   3 - 0x3
      13'h1EAF: dout <= 8'b00000000; // 7855 :   0 - 0x0
      13'h1EB0: dout <= 8'b00000000; // 7856 :   0 - 0x0 -- Background 0xeb
      13'h1EB1: dout <= 8'b00001100; // 7857 :  12 - 0xc
      13'h1EB2: dout <= 8'b00000110; // 7858 :   6 - 0x6
      13'h1EB3: dout <= 8'b00000110; // 7859 :   6 - 0x6
      13'h1EB4: dout <= 8'b01100000; // 7860 :  96 - 0x60
      13'h1EB5: dout <= 8'b01110000; // 7861 : 112 - 0x70
      13'h1EB6: dout <= 8'b00110000; // 7862 :  48 - 0x30
      13'h1EB7: dout <= 8'b00000000; // 7863 :   0 - 0x0
      13'h1EB8: dout <= 8'b00000000; // 7864 :   0 - 0x0
      13'h1EB9: dout <= 8'b00001100; // 7865 :  12 - 0xc
      13'h1EBA: dout <= 8'b00000110; // 7866 :   6 - 0x6
      13'h1EBB: dout <= 8'b00000110; // 7867 :   6 - 0x6
      13'h1EBC: dout <= 8'b01100000; // 7868 :  96 - 0x60
      13'h1EBD: dout <= 8'b01110000; // 7869 : 112 - 0x70
      13'h1EBE: dout <= 8'b00110000; // 7870 :  48 - 0x30
      13'h1EBF: dout <= 8'b00000000; // 7871 :   0 - 0x0
      13'h1EC0: dout <= 8'b00000000; // 7872 :   0 - 0x0 -- Background 0xec
      13'h1EC1: dout <= 8'b11000000; // 7873 : 192 - 0xc0
      13'h1EC2: dout <= 8'b11100000; // 7874 : 224 - 0xe0
      13'h1EC3: dout <= 8'b01100000; // 7875 :  96 - 0x60
      13'h1EC4: dout <= 8'b00000000; // 7876 :   0 - 0x0
      13'h1EC5: dout <= 8'b00001100; // 7877 :  12 - 0xc
      13'h1EC6: dout <= 8'b00001110; // 7878 :  14 - 0xe
      13'h1EC7: dout <= 8'b00000110; // 7879 :   6 - 0x6
      13'h1EC8: dout <= 8'b00000000; // 7880 :   0 - 0x0
      13'h1EC9: dout <= 8'b11000000; // 7881 : 192 - 0xc0
      13'h1ECA: dout <= 8'b11100000; // 7882 : 224 - 0xe0
      13'h1ECB: dout <= 8'b01100000; // 7883 :  96 - 0x60
      13'h1ECC: dout <= 8'b00000000; // 7884 :   0 - 0x0
      13'h1ECD: dout <= 8'b00001100; // 7885 :  12 - 0xc
      13'h1ECE: dout <= 8'b00001110; // 7886 :  14 - 0xe
      13'h1ECF: dout <= 8'b00000110; // 7887 :   6 - 0x6
      13'h1ED0: dout <= 8'b01100000; // 7888 :  96 - 0x60 -- Background 0xed
      13'h1ED1: dout <= 8'b01110000; // 7889 : 112 - 0x70
      13'h1ED2: dout <= 8'b00110000; // 7890 :  48 - 0x30
      13'h1ED3: dout <= 8'b00000000; // 7891 :   0 - 0x0
      13'h1ED4: dout <= 8'b00000000; // 7892 :   0 - 0x0
      13'h1ED5: dout <= 8'b00001100; // 7893 :  12 - 0xc
      13'h1ED6: dout <= 8'b00001110; // 7894 :  14 - 0xe
      13'h1ED7: dout <= 8'b00000110; // 7895 :   6 - 0x6
      13'h1ED8: dout <= 8'b01100000; // 7896 :  96 - 0x60
      13'h1ED9: dout <= 8'b01110000; // 7897 : 112 - 0x70
      13'h1EDA: dout <= 8'b00110000; // 7898 :  48 - 0x30
      13'h1EDB: dout <= 8'b00000000; // 7899 :   0 - 0x0
      13'h1EDC: dout <= 8'b00000000; // 7900 :   0 - 0x0
      13'h1EDD: dout <= 8'b00001100; // 7901 :  12 - 0xc
      13'h1EDE: dout <= 8'b00001110; // 7902 :  14 - 0xe
      13'h1EDF: dout <= 8'b00000110; // 7903 :   6 - 0x6
      13'h1EE0: dout <= 8'b11111111; // 7904 : 255 - 0xff -- Background 0xee
      13'h1EE1: dout <= 8'b11111111; // 7905 : 255 - 0xff
      13'h1EE2: dout <= 8'b10111101; // 7906 : 189 - 0xbd
      13'h1EE3: dout <= 8'b11111111; // 7907 : 255 - 0xff
      13'h1EE4: dout <= 8'b11111111; // 7908 : 255 - 0xff
      13'h1EE5: dout <= 8'b11111011; // 7909 : 251 - 0xfb
      13'h1EE6: dout <= 8'b11111111; // 7910 : 255 - 0xff
      13'h1EE7: dout <= 8'b11111111; // 7911 : 255 - 0xff
      13'h1EE8: dout <= 8'b00000000; // 7912 :   0 - 0x0
      13'h1EE9: dout <= 8'b00000000; // 7913 :   0 - 0x0
      13'h1EEA: dout <= 8'b01000010; // 7914 :  66 - 0x42
      13'h1EEB: dout <= 8'b00000000; // 7915 :   0 - 0x0
      13'h1EEC: dout <= 8'b00000000; // 7916 :   0 - 0x0
      13'h1EED: dout <= 8'b00000100; // 7917 :   4 - 0x4
      13'h1EEE: dout <= 8'b00000000; // 7918 :   0 - 0x0
      13'h1EEF: dout <= 8'b00000000; // 7919 :   0 - 0x0
      13'h1EF0: dout <= 8'b11111111; // 7920 : 255 - 0xff -- Background 0xef
      13'h1EF1: dout <= 8'b11111111; // 7921 : 255 - 0xff
      13'h1EF2: dout <= 8'b11111011; // 7922 : 251 - 0xfb
      13'h1EF3: dout <= 8'b11111111; // 7923 : 255 - 0xff
      13'h1EF4: dout <= 8'b11011111; // 7924 : 223 - 0xdf
      13'h1EF5: dout <= 8'b11111111; // 7925 : 255 - 0xff
      13'h1EF6: dout <= 8'b11111111; // 7926 : 255 - 0xff
      13'h1EF7: dout <= 8'b11111111; // 7927 : 255 - 0xff
      13'h1EF8: dout <= 8'b00000000; // 7928 :   0 - 0x0
      13'h1EF9: dout <= 8'b00000000; // 7929 :   0 - 0x0
      13'h1EFA: dout <= 8'b00000100; // 7930 :   4 - 0x4
      13'h1EFB: dout <= 8'b00000000; // 7931 :   0 - 0x0
      13'h1EFC: dout <= 8'b00100000; // 7932 :  32 - 0x20
      13'h1EFD: dout <= 8'b00000000; // 7933 :   0 - 0x0
      13'h1EFE: dout <= 8'b00000000; // 7934 :   0 - 0x0
      13'h1EFF: dout <= 8'b00000000; // 7935 :   0 - 0x0
      13'h1F00: dout <= 8'b00000000; // 7936 :   0 - 0x0 -- Background 0xf0
      13'h1F01: dout <= 8'b00000000; // 7937 :   0 - 0x0
      13'h1F02: dout <= 8'b00000000; // 7938 :   0 - 0x0
      13'h1F03: dout <= 8'b00000000; // 7939 :   0 - 0x0
      13'h1F04: dout <= 8'b00000000; // 7940 :   0 - 0x0
      13'h1F05: dout <= 8'b00000000; // 7941 :   0 - 0x0
      13'h1F06: dout <= 8'b00000000; // 7942 :   0 - 0x0
      13'h1F07: dout <= 8'b00000000; // 7943 :   0 - 0x0
      13'h1F08: dout <= 8'b00000000; // 7944 :   0 - 0x0
      13'h1F09: dout <= 8'b00000000; // 7945 :   0 - 0x0
      13'h1F0A: dout <= 8'b00000000; // 7946 :   0 - 0x0
      13'h1F0B: dout <= 8'b00000000; // 7947 :   0 - 0x0
      13'h1F0C: dout <= 8'b00000000; // 7948 :   0 - 0x0
      13'h1F0D: dout <= 8'b00000000; // 7949 :   0 - 0x0
      13'h1F0E: dout <= 8'b00000000; // 7950 :   0 - 0x0
      13'h1F0F: dout <= 8'b00000000; // 7951 :   0 - 0x0
      13'h1F10: dout <= 8'b00000000; // 7952 :   0 - 0x0 -- Background 0xf1
      13'h1F11: dout <= 8'b10000000; // 7953 : 128 - 0x80
      13'h1F12: dout <= 8'b00000000; // 7954 :   0 - 0x0
      13'h1F13: dout <= 8'b00000000; // 7955 :   0 - 0x0
      13'h1F14: dout <= 8'b00000000; // 7956 :   0 - 0x0
      13'h1F15: dout <= 8'b00000000; // 7957 :   0 - 0x0
      13'h1F16: dout <= 8'b00000000; // 7958 :   0 - 0x0
      13'h1F17: dout <= 8'b00000000; // 7959 :   0 - 0x0
      13'h1F18: dout <= 8'b10000000; // 7960 : 128 - 0x80
      13'h1F19: dout <= 8'b10000000; // 7961 : 128 - 0x80
      13'h1F1A: dout <= 8'b10000000; // 7962 : 128 - 0x80
      13'h1F1B: dout <= 8'b10000000; // 7963 : 128 - 0x80
      13'h1F1C: dout <= 8'b00000000; // 7964 :   0 - 0x0
      13'h1F1D: dout <= 8'b00000000; // 7965 :   0 - 0x0
      13'h1F1E: dout <= 8'b00000000; // 7966 :   0 - 0x0
      13'h1F1F: dout <= 8'b00000000; // 7967 :   0 - 0x0
      13'h1F20: dout <= 8'b00000000; // 7968 :   0 - 0x0 -- Background 0xf2
      13'h1F21: dout <= 8'b11000000; // 7969 : 192 - 0xc0
      13'h1F22: dout <= 8'b00000000; // 7970 :   0 - 0x0
      13'h1F23: dout <= 8'b00000000; // 7971 :   0 - 0x0
      13'h1F24: dout <= 8'b00000000; // 7972 :   0 - 0x0
      13'h1F25: dout <= 8'b00000000; // 7973 :   0 - 0x0
      13'h1F26: dout <= 8'b00000000; // 7974 :   0 - 0x0
      13'h1F27: dout <= 8'b00000000; // 7975 :   0 - 0x0
      13'h1F28: dout <= 8'b11000000; // 7976 : 192 - 0xc0
      13'h1F29: dout <= 8'b11000000; // 7977 : 192 - 0xc0
      13'h1F2A: dout <= 8'b11000000; // 7978 : 192 - 0xc0
      13'h1F2B: dout <= 8'b11000000; // 7979 : 192 - 0xc0
      13'h1F2C: dout <= 8'b00000000; // 7980 :   0 - 0x0
      13'h1F2D: dout <= 8'b00000000; // 7981 :   0 - 0x0
      13'h1F2E: dout <= 8'b00000000; // 7982 :   0 - 0x0
      13'h1F2F: dout <= 8'b00000000; // 7983 :   0 - 0x0
      13'h1F30: dout <= 8'b00000000; // 7984 :   0 - 0x0 -- Background 0xf3
      13'h1F31: dout <= 8'b11100000; // 7985 : 224 - 0xe0
      13'h1F32: dout <= 8'b00000000; // 7986 :   0 - 0x0
      13'h1F33: dout <= 8'b00000000; // 7987 :   0 - 0x0
      13'h1F34: dout <= 8'b00000000; // 7988 :   0 - 0x0
      13'h1F35: dout <= 8'b00000000; // 7989 :   0 - 0x0
      13'h1F36: dout <= 8'b00000000; // 7990 :   0 - 0x0
      13'h1F37: dout <= 8'b00000000; // 7991 :   0 - 0x0
      13'h1F38: dout <= 8'b11100000; // 7992 : 224 - 0xe0
      13'h1F39: dout <= 8'b11100000; // 7993 : 224 - 0xe0
      13'h1F3A: dout <= 8'b11100000; // 7994 : 224 - 0xe0
      13'h1F3B: dout <= 8'b11100000; // 7995 : 224 - 0xe0
      13'h1F3C: dout <= 8'b00000000; // 7996 :   0 - 0x0
      13'h1F3D: dout <= 8'b00000000; // 7997 :   0 - 0x0
      13'h1F3E: dout <= 8'b00000000; // 7998 :   0 - 0x0
      13'h1F3F: dout <= 8'b00000000; // 7999 :   0 - 0x0
      13'h1F40: dout <= 8'b00000000; // 8000 :   0 - 0x0 -- Background 0xf4
      13'h1F41: dout <= 8'b11110000; // 8001 : 240 - 0xf0
      13'h1F42: dout <= 8'b00000000; // 8002 :   0 - 0x0
      13'h1F43: dout <= 8'b00000000; // 8003 :   0 - 0x0
      13'h1F44: dout <= 8'b00000000; // 8004 :   0 - 0x0
      13'h1F45: dout <= 8'b00000000; // 8005 :   0 - 0x0
      13'h1F46: dout <= 8'b00000000; // 8006 :   0 - 0x0
      13'h1F47: dout <= 8'b00000000; // 8007 :   0 - 0x0
      13'h1F48: dout <= 8'b11110000; // 8008 : 240 - 0xf0
      13'h1F49: dout <= 8'b11110000; // 8009 : 240 - 0xf0
      13'h1F4A: dout <= 8'b11110000; // 8010 : 240 - 0xf0
      13'h1F4B: dout <= 8'b11110000; // 8011 : 240 - 0xf0
      13'h1F4C: dout <= 8'b00000000; // 8012 :   0 - 0x0
      13'h1F4D: dout <= 8'b00000000; // 8013 :   0 - 0x0
      13'h1F4E: dout <= 8'b00000000; // 8014 :   0 - 0x0
      13'h1F4F: dout <= 8'b00000000; // 8015 :   0 - 0x0
      13'h1F50: dout <= 8'b00000000; // 8016 :   0 - 0x0 -- Background 0xf5
      13'h1F51: dout <= 8'b11111000; // 8017 : 248 - 0xf8
      13'h1F52: dout <= 8'b00000000; // 8018 :   0 - 0x0
      13'h1F53: dout <= 8'b00000000; // 8019 :   0 - 0x0
      13'h1F54: dout <= 8'b00000000; // 8020 :   0 - 0x0
      13'h1F55: dout <= 8'b00000000; // 8021 :   0 - 0x0
      13'h1F56: dout <= 8'b00000000; // 8022 :   0 - 0x0
      13'h1F57: dout <= 8'b00000000; // 8023 :   0 - 0x0
      13'h1F58: dout <= 8'b11111000; // 8024 : 248 - 0xf8
      13'h1F59: dout <= 8'b11111000; // 8025 : 248 - 0xf8
      13'h1F5A: dout <= 8'b11111000; // 8026 : 248 - 0xf8
      13'h1F5B: dout <= 8'b11111000; // 8027 : 248 - 0xf8
      13'h1F5C: dout <= 8'b00000000; // 8028 :   0 - 0x0
      13'h1F5D: dout <= 8'b00000000; // 8029 :   0 - 0x0
      13'h1F5E: dout <= 8'b00000000; // 8030 :   0 - 0x0
      13'h1F5F: dout <= 8'b00000000; // 8031 :   0 - 0x0
      13'h1F60: dout <= 8'b00000000; // 8032 :   0 - 0x0 -- Background 0xf6
      13'h1F61: dout <= 8'b11111100; // 8033 : 252 - 0xfc
      13'h1F62: dout <= 8'b00000000; // 8034 :   0 - 0x0
      13'h1F63: dout <= 8'b00000000; // 8035 :   0 - 0x0
      13'h1F64: dout <= 8'b00000000; // 8036 :   0 - 0x0
      13'h1F65: dout <= 8'b00000000; // 8037 :   0 - 0x0
      13'h1F66: dout <= 8'b00000000; // 8038 :   0 - 0x0
      13'h1F67: dout <= 8'b00000000; // 8039 :   0 - 0x0
      13'h1F68: dout <= 8'b11111100; // 8040 : 252 - 0xfc
      13'h1F69: dout <= 8'b11111100; // 8041 : 252 - 0xfc
      13'h1F6A: dout <= 8'b11111100; // 8042 : 252 - 0xfc
      13'h1F6B: dout <= 8'b11111100; // 8043 : 252 - 0xfc
      13'h1F6C: dout <= 8'b00000000; // 8044 :   0 - 0x0
      13'h1F6D: dout <= 8'b00000000; // 8045 :   0 - 0x0
      13'h1F6E: dout <= 8'b00000000; // 8046 :   0 - 0x0
      13'h1F6F: dout <= 8'b00000000; // 8047 :   0 - 0x0
      13'h1F70: dout <= 8'b00000000; // 8048 :   0 - 0x0 -- Background 0xf7
      13'h1F71: dout <= 8'b11111110; // 8049 : 254 - 0xfe
      13'h1F72: dout <= 8'b00000000; // 8050 :   0 - 0x0
      13'h1F73: dout <= 8'b00000000; // 8051 :   0 - 0x0
      13'h1F74: dout <= 8'b00000000; // 8052 :   0 - 0x0
      13'h1F75: dout <= 8'b00000000; // 8053 :   0 - 0x0
      13'h1F76: dout <= 8'b00000000; // 8054 :   0 - 0x0
      13'h1F77: dout <= 8'b00000000; // 8055 :   0 - 0x0
      13'h1F78: dout <= 8'b11111110; // 8056 : 254 - 0xfe
      13'h1F79: dout <= 8'b11111110; // 8057 : 254 - 0xfe
      13'h1F7A: dout <= 8'b11111110; // 8058 : 254 - 0xfe
      13'h1F7B: dout <= 8'b11111110; // 8059 : 254 - 0xfe
      13'h1F7C: dout <= 8'b00000000; // 8060 :   0 - 0x0
      13'h1F7D: dout <= 8'b00000000; // 8061 :   0 - 0x0
      13'h1F7E: dout <= 8'b00000000; // 8062 :   0 - 0x0
      13'h1F7F: dout <= 8'b00000000; // 8063 :   0 - 0x0
      13'h1F80: dout <= 8'b00000000; // 8064 :   0 - 0x0 -- Background 0xf8
      13'h1F81: dout <= 8'b11111111; // 8065 : 255 - 0xff
      13'h1F82: dout <= 8'b00000000; // 8066 :   0 - 0x0
      13'h1F83: dout <= 8'b00000000; // 8067 :   0 - 0x0
      13'h1F84: dout <= 8'b00000000; // 8068 :   0 - 0x0
      13'h1F85: dout <= 8'b00000000; // 8069 :   0 - 0x0
      13'h1F86: dout <= 8'b00000000; // 8070 :   0 - 0x0
      13'h1F87: dout <= 8'b00000000; // 8071 :   0 - 0x0
      13'h1F88: dout <= 8'b11111111; // 8072 : 255 - 0xff
      13'h1F89: dout <= 8'b11111111; // 8073 : 255 - 0xff
      13'h1F8A: dout <= 8'b11111111; // 8074 : 255 - 0xff
      13'h1F8B: dout <= 8'b11111111; // 8075 : 255 - 0xff
      13'h1F8C: dout <= 8'b00000000; // 8076 :   0 - 0x0
      13'h1F8D: dout <= 8'b00000000; // 8077 :   0 - 0x0
      13'h1F8E: dout <= 8'b00000000; // 8078 :   0 - 0x0
      13'h1F8F: dout <= 8'b00000000; // 8079 :   0 - 0x0
      13'h1F90: dout <= 8'b11111111; // 8080 : 255 - 0xff -- Background 0xf9
      13'h1F91: dout <= 8'b11111111; // 8081 : 255 - 0xff
      13'h1F92: dout <= 8'b11111111; // 8082 : 255 - 0xff
      13'h1F93: dout <= 8'b11111111; // 8083 : 255 - 0xff
      13'h1F94: dout <= 8'b10000000; // 8084 : 128 - 0x80
      13'h1F95: dout <= 8'b10000000; // 8085 : 128 - 0x80
      13'h1F96: dout <= 8'b11000000; // 8086 : 192 - 0xc0
      13'h1F97: dout <= 8'b11000000; // 8087 : 192 - 0xc0
      13'h1F98: dout <= 8'b00000000; // 8088 :   0 - 0x0
      13'h1F99: dout <= 8'b00000000; // 8089 :   0 - 0x0
      13'h1F9A: dout <= 8'b00000000; // 8090 :   0 - 0x0
      13'h1F9B: dout <= 8'b00000000; // 8091 :   0 - 0x0
      13'h1F9C: dout <= 8'b01111111; // 8092 : 127 - 0x7f
      13'h1F9D: dout <= 8'b01000000; // 8093 :  64 - 0x40
      13'h1F9E: dout <= 8'b01000000; // 8094 :  64 - 0x40
      13'h1F9F: dout <= 8'b01000000; // 8095 :  64 - 0x40
      13'h1FA0: dout <= 8'b11111111; // 8096 : 255 - 0xff -- Background 0xfa
      13'h1FA1: dout <= 8'b11111111; // 8097 : 255 - 0xff
      13'h1FA2: dout <= 8'b11111111; // 8098 : 255 - 0xff
      13'h1FA3: dout <= 8'b11111111; // 8099 : 255 - 0xff
      13'h1FA4: dout <= 8'b00000000; // 8100 :   0 - 0x0
      13'h1FA5: dout <= 8'b00000000; // 8101 :   0 - 0x0
      13'h1FA6: dout <= 8'b00000000; // 8102 :   0 - 0x0
      13'h1FA7: dout <= 8'b00000000; // 8103 :   0 - 0x0
      13'h1FA8: dout <= 8'b00000000; // 8104 :   0 - 0x0
      13'h1FA9: dout <= 8'b00000000; // 8105 :   0 - 0x0
      13'h1FAA: dout <= 8'b00000000; // 8106 :   0 - 0x0
      13'h1FAB: dout <= 8'b00000000; // 8107 :   0 - 0x0
      13'h1FAC: dout <= 8'b11111111; // 8108 : 255 - 0xff
      13'h1FAD: dout <= 8'b00000000; // 8109 :   0 - 0x0
      13'h1FAE: dout <= 8'b00000000; // 8110 :   0 - 0x0
      13'h1FAF: dout <= 8'b00000000; // 8111 :   0 - 0x0
      13'h1FB0: dout <= 8'b11111111; // 8112 : 255 - 0xff -- Background 0xfb
      13'h1FB1: dout <= 8'b11111111; // 8113 : 255 - 0xff
      13'h1FB2: dout <= 8'b11111111; // 8114 : 255 - 0xff
      13'h1FB3: dout <= 8'b11111111; // 8115 : 255 - 0xff
      13'h1FB4: dout <= 8'b00000001; // 8116 :   1 - 0x1
      13'h1FB5: dout <= 8'b00000000; // 8117 :   0 - 0x0
      13'h1FB6: dout <= 8'b00000010; // 8118 :   2 - 0x2
      13'h1FB7: dout <= 8'b00000010; // 8119 :   2 - 0x2
      13'h1FB8: dout <= 8'b00000000; // 8120 :   0 - 0x0
      13'h1FB9: dout <= 8'b00000000; // 8121 :   0 - 0x0
      13'h1FBA: dout <= 8'b00000000; // 8122 :   0 - 0x0
      13'h1FBB: dout <= 8'b00000000; // 8123 :   0 - 0x0
      13'h1FBC: dout <= 8'b11111110; // 8124 : 254 - 0xfe
      13'h1FBD: dout <= 8'b00000010; // 8125 :   2 - 0x2
      13'h1FBE: dout <= 8'b00000010; // 8126 :   2 - 0x2
      13'h1FBF: dout <= 8'b00000010; // 8127 :   2 - 0x2
      13'h1FC0: dout <= 8'b11000000; // 8128 : 192 - 0xc0 -- Background 0xfc
      13'h1FC1: dout <= 8'b11000000; // 8129 : 192 - 0xc0
      13'h1FC2: dout <= 8'b10000000; // 8130 : 128 - 0x80
      13'h1FC3: dout <= 8'b10000000; // 8131 : 128 - 0x80
      13'h1FC4: dout <= 8'b11000000; // 8132 : 192 - 0xc0
      13'h1FC5: dout <= 8'b11111111; // 8133 : 255 - 0xff
      13'h1FC6: dout <= 8'b11111111; // 8134 : 255 - 0xff
      13'h1FC7: dout <= 8'b11111111; // 8135 : 255 - 0xff
      13'h1FC8: dout <= 8'b01000000; // 8136 :  64 - 0x40
      13'h1FC9: dout <= 8'b01000000; // 8137 :  64 - 0x40
      13'h1FCA: dout <= 8'b01000000; // 8138 :  64 - 0x40
      13'h1FCB: dout <= 8'b01111111; // 8139 : 127 - 0x7f
      13'h1FCC: dout <= 8'b00000000; // 8140 :   0 - 0x0
      13'h1FCD: dout <= 8'b00000000; // 8141 :   0 - 0x0
      13'h1FCE: dout <= 8'b00000000; // 8142 :   0 - 0x0
      13'h1FCF: dout <= 8'b00000000; // 8143 :   0 - 0x0
      13'h1FD0: dout <= 8'b00000000; // 8144 :   0 - 0x0 -- Background 0xfd
      13'h1FD1: dout <= 8'b00000000; // 8145 :   0 - 0x0
      13'h1FD2: dout <= 8'b00000000; // 8146 :   0 - 0x0
      13'h1FD3: dout <= 8'b00000000; // 8147 :   0 - 0x0
      13'h1FD4: dout <= 8'b00000000; // 8148 :   0 - 0x0
      13'h1FD5: dout <= 8'b11111111; // 8149 : 255 - 0xff
      13'h1FD6: dout <= 8'b11111111; // 8150 : 255 - 0xff
      13'h1FD7: dout <= 8'b11111111; // 8151 : 255 - 0xff
      13'h1FD8: dout <= 8'b00000000; // 8152 :   0 - 0x0
      13'h1FD9: dout <= 8'b00000000; // 8153 :   0 - 0x0
      13'h1FDA: dout <= 8'b00000000; // 8154 :   0 - 0x0
      13'h1FDB: dout <= 8'b11111111; // 8155 : 255 - 0xff
      13'h1FDC: dout <= 8'b00000000; // 8156 :   0 - 0x0
      13'h1FDD: dout <= 8'b00000000; // 8157 :   0 - 0x0
      13'h1FDE: dout <= 8'b00000000; // 8158 :   0 - 0x0
      13'h1FDF: dout <= 8'b00000000; // 8159 :   0 - 0x0
      13'h1FE0: dout <= 8'b00000010; // 8160 :   2 - 0x2 -- Background 0xfe
      13'h1FE1: dout <= 8'b00000010; // 8161 :   2 - 0x2
      13'h1FE2: dout <= 8'b00000000; // 8162 :   0 - 0x0
      13'h1FE3: dout <= 8'b00000000; // 8163 :   0 - 0x0
      13'h1FE4: dout <= 8'b00000000; // 8164 :   0 - 0x0
      13'h1FE5: dout <= 8'b11111111; // 8165 : 255 - 0xff
      13'h1FE6: dout <= 8'b11111111; // 8166 : 255 - 0xff
      13'h1FE7: dout <= 8'b11111111; // 8167 : 255 - 0xff
      13'h1FE8: dout <= 8'b00000010; // 8168 :   2 - 0x2
      13'h1FE9: dout <= 8'b00000010; // 8169 :   2 - 0x2
      13'h1FEA: dout <= 8'b00000010; // 8170 :   2 - 0x2
      13'h1FEB: dout <= 8'b11111110; // 8171 : 254 - 0xfe
      13'h1FEC: dout <= 8'b00000000; // 8172 :   0 - 0x0
      13'h1FED: dout <= 8'b00000000; // 8173 :   0 - 0x0
      13'h1FEE: dout <= 8'b00000000; // 8174 :   0 - 0x0
      13'h1FEF: dout <= 8'b00000000; // 8175 :   0 - 0x0
      13'h1FF0: dout <= 8'b11111111; // 8176 : 255 - 0xff -- Background 0xff
      13'h1FF1: dout <= 8'b11111111; // 8177 : 255 - 0xff
      13'h1FF2: dout <= 8'b11111111; // 8178 : 255 - 0xff
      13'h1FF3: dout <= 8'b11111111; // 8179 : 255 - 0xff
      13'h1FF4: dout <= 8'b11111111; // 8180 : 255 - 0xff
      13'h1FF5: dout <= 8'b11111111; // 8181 : 255 - 0xff
      13'h1FF6: dout <= 8'b11111111; // 8182 : 255 - 0xff
      13'h1FF7: dout <= 8'b11111111; // 8183 : 255 - 0xff
      13'h1FF8: dout <= 8'b00000000; // 8184 :   0 - 0x0
      13'h1FF9: dout <= 8'b00000000; // 8185 :   0 - 0x0
      13'h1FFA: dout <= 8'b00000000; // 8186 :   0 - 0x0
      13'h1FFB: dout <= 8'b00000000; // 8187 :   0 - 0x0
      13'h1FFC: dout <= 8'b00000000; // 8188 :   0 - 0x0
      13'h1FFD: dout <= 8'b00000000; // 8189 :   0 - 0x0
      13'h1FFE: dout <= 8'b00000000; // 8190 :   0 - 0x0
      13'h1FFF: dout <= 8'b00000000; // 8191 :   0 - 0x0
    endcase
  end

endmodule
