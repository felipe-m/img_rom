//-   Sprites Pattern table COLOR PLANE 1
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
//- Autcmatically generated verilog ROM from a NES memory file----


//-  Original memory dump file name: smario_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_PTABLE_SMARIO_SPR_PLN1
  (
     //input     clk,   // clock
     input      [11-1:0] addr,  //2048 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Sprite pattern Table COLOR PLANE 1
      11'h0: dout  = 8'b00000000; //    0 :   0 - 0x0 -- Sprite 0x0
      11'h1: dout  = 8'b00000000; //    1 :   0 - 0x0
      11'h2: dout  = 8'b00000000; //    2 :   0 - 0x0
      11'h3: dout  = 8'b00000000; //    3 :   0 - 0x0
      11'h4: dout  = 8'b00011111; //    4 :  31 - 0x1f
      11'h5: dout  = 8'b00111111; //    5 :  63 - 0x3f
      11'h6: dout  = 8'b00111111; //    6 :  63 - 0x3f
      11'h7: dout  = 8'b01111111; //    7 : 127 - 0x7f
      11'h8: dout  = 8'b00000000; //    8 :   0 - 0x0 -- Sprite 0x1
      11'h9: dout  = 8'b00100000; //    9 :  32 - 0x20
      11'hA: dout  = 8'b01100000; //   10 :  96 - 0x60
      11'hB: dout  = 8'b00000000; //   11 :   0 - 0x0
      11'hC: dout  = 8'b11110000; //   12 : 240 - 0xf0
      11'hD: dout  = 8'b11111100; //   13 : 252 - 0xfc
      11'hE: dout  = 8'b11111110; //   14 : 254 - 0xfe
      11'hF: dout  = 8'b11111110; //   15 : 254 - 0xfe
      11'h10: dout  = 8'b01111111; //   16 : 127 - 0x7f -- Sprite 0x2
      11'h11: dout  = 8'b01111111; //   17 : 127 - 0x7f
      11'h12: dout  = 8'b00011111; //   18 :  31 - 0x1f
      11'h13: dout  = 8'b00000111; //   19 :   7 - 0x7
      11'h14: dout  = 8'b00000000; //   20 :   0 - 0x0
      11'h15: dout  = 8'b00011110; //   21 :  30 - 0x1e
      11'h16: dout  = 8'b00111111; //   22 :  63 - 0x3f
      11'h17: dout  = 8'b01111111; //   23 : 127 - 0x7f
      11'h18: dout  = 8'b11111100; //   24 : 252 - 0xfc -- Sprite 0x3
      11'h19: dout  = 8'b11111100; //   25 : 252 - 0xfc
      11'h1A: dout  = 8'b11111000; //   26 : 248 - 0xf8
      11'h1B: dout  = 8'b11000000; //   27 : 192 - 0xc0
      11'h1C: dout  = 8'b11000010; //   28 : 194 - 0xc2
      11'h1D: dout  = 8'b01100111; //   29 : 103 - 0x67
      11'h1E: dout  = 8'b00101111; //   30 :  47 - 0x2f
      11'h1F: dout  = 8'b00110111; //   31 :  55 - 0x37
      11'h20: dout  = 8'b01111111; //   32 : 127 - 0x7f -- Sprite 0x4
      11'h21: dout  = 8'b01111110; //   33 : 126 - 0x7e
      11'h22: dout  = 8'b11111100; //   34 : 252 - 0xfc
      11'h23: dout  = 8'b11110000; //   35 : 240 - 0xf0
      11'h24: dout  = 8'b11111000; //   36 : 248 - 0xf8
      11'h25: dout  = 8'b11111000; //   37 : 248 - 0xf8
      11'h26: dout  = 8'b11110000; //   38 : 240 - 0xf0
      11'h27: dout  = 8'b01110000; //   39 : 112 - 0x70
      11'h28: dout  = 8'b00110111; //   40 :  55 - 0x37 -- Sprite 0x5
      11'h29: dout  = 8'b00110110; //   41 :  54 - 0x36
      11'h2A: dout  = 8'b01011100; //   42 :  92 - 0x5c
      11'h2B: dout  = 8'b00000000; //   43 :   0 - 0x0
      11'h2C: dout  = 8'b00000000; //   44 :   0 - 0x0
      11'h2D: dout  = 8'b00000001; //   45 :   1 - 0x1
      11'h2E: dout  = 8'b00000011; //   46 :   3 - 0x3
      11'h2F: dout  = 8'b00011111; //   47 :  31 - 0x1f
      11'h30: dout  = 8'b00001000; //   48 :   8 - 0x8 -- Sprite 0x6
      11'h31: dout  = 8'b00100100; //   49 :  36 - 0x24
      11'h32: dout  = 8'b11100011; //   50 : 227 - 0xe3
      11'h33: dout  = 8'b11110000; //   51 : 240 - 0xf0
      11'h34: dout  = 8'b11111000; //   52 : 248 - 0xf8
      11'h35: dout  = 8'b01110000; //   53 : 112 - 0x70
      11'h36: dout  = 8'b01110000; //   54 : 112 - 0x70
      11'h37: dout  = 8'b00111000; //   55 :  56 - 0x38
      11'h38: dout  = 8'b00011111; //   56 :  31 - 0x1f -- Sprite 0x7
      11'h39: dout  = 8'b00011111; //   57 :  31 - 0x1f
      11'h3A: dout  = 8'b00011111; //   58 :  31 - 0x1f
      11'h3B: dout  = 8'b00011111; //   59 :  31 - 0x1f
      11'h3C: dout  = 8'b00000000; //   60 :   0 - 0x0
      11'h3D: dout  = 8'b00000000; //   61 :   0 - 0x0
      11'h3E: dout  = 8'b00000000; //   62 :   0 - 0x0
      11'h3F: dout  = 8'b00000000; //   63 :   0 - 0x0
      11'h40: dout  = 8'b00000000; //   64 :   0 - 0x0 -- Sprite 0x8
      11'h41: dout  = 8'b00000000; //   65 :   0 - 0x0
      11'h42: dout  = 8'b00000000; //   66 :   0 - 0x0
      11'h43: dout  = 8'b00000000; //   67 :   0 - 0x0
      11'h44: dout  = 8'b00000000; //   68 :   0 - 0x0
      11'h45: dout  = 8'b00000000; //   69 :   0 - 0x0
      11'h46: dout  = 8'b00001111; //   70 :  15 - 0xf
      11'h47: dout  = 8'b00011111; //   71 :  31 - 0x1f
      11'h48: dout  = 8'b00000000; //   72 :   0 - 0x0 -- Sprite 0x9
      11'h49: dout  = 8'b00000000; //   73 :   0 - 0x0
      11'h4A: dout  = 8'b00000000; //   74 :   0 - 0x0
      11'h4B: dout  = 8'b00010000; //   75 :  16 - 0x10
      11'h4C: dout  = 8'b00110000; //   76 :  48 - 0x30
      11'h4D: dout  = 8'b00000000; //   77 :   0 - 0x0
      11'h4E: dout  = 8'b11111000; //   78 : 248 - 0xf8
      11'h4F: dout  = 8'b11111110; //   79 : 254 - 0xfe
      11'h50: dout  = 8'b00011111; //   80 :  31 - 0x1f -- Sprite 0xa
      11'h51: dout  = 8'b00111111; //   81 :  63 - 0x3f
      11'h52: dout  = 8'b00111111; //   82 :  63 - 0x3f
      11'h53: dout  = 8'b00011111; //   83 :  31 - 0x1f
      11'h54: dout  = 8'b00000111; //   84 :   7 - 0x7
      11'h55: dout  = 8'b00001000; //   85 :   8 - 0x8
      11'h56: dout  = 8'b00010111; //   86 :  23 - 0x17
      11'h57: dout  = 8'b00010111; //   87 :  23 - 0x17
      11'h58: dout  = 8'b11111111; //   88 : 255 - 0xff -- Sprite 0xb
      11'h59: dout  = 8'b11111111; //   89 : 255 - 0xff
      11'h5A: dout  = 8'b11111110; //   90 : 254 - 0xfe
      11'h5B: dout  = 8'b11111110; //   91 : 254 - 0xfe
      11'h5C: dout  = 8'b11111100; //   92 : 252 - 0xfc
      11'h5D: dout  = 8'b11100000; //   93 : 224 - 0xe0
      11'h5E: dout  = 8'b01000000; //   94 :  64 - 0x40
      11'h5F: dout  = 8'b10100000; //   95 : 160 - 0xa0
      11'h60: dout  = 8'b00110111; //   96 :  55 - 0x37 -- Sprite 0xc
      11'h61: dout  = 8'b00100111; //   97 :  39 - 0x27
      11'h62: dout  = 8'b00100011; //   98 :  35 - 0x23
      11'h63: dout  = 8'b00000011; //   99 :   3 - 0x3
      11'h64: dout  = 8'b00000001; //  100 :   1 - 0x1
      11'h65: dout  = 8'b00000000; //  101 :   0 - 0x0
      11'h66: dout  = 8'b00000000; //  102 :   0 - 0x0
      11'h67: dout  = 8'b00000000; //  103 :   0 - 0x0
      11'h68: dout  = 8'b11001100; //  104 : 204 - 0xcc -- Sprite 0xd
      11'h69: dout  = 8'b11111111; //  105 : 255 - 0xff
      11'h6A: dout  = 8'b11111111; //  106 : 255 - 0xff
      11'h6B: dout  = 8'b11111111; //  107 : 255 - 0xff
      11'h6C: dout  = 8'b11111111; //  108 : 255 - 0xff
      11'h6D: dout  = 8'b01110000; //  109 : 112 - 0x70
      11'h6E: dout  = 8'b00000000; //  110 :   0 - 0x0
      11'h6F: dout  = 8'b00001000; //  111 :   8 - 0x8
      11'h70: dout  = 8'b11110000; //  112 : 240 - 0xf0 -- Sprite 0xe
      11'h71: dout  = 8'b11110000; //  113 : 240 - 0xf0
      11'h72: dout  = 8'b11110000; //  114 : 240 - 0xf0
      11'h73: dout  = 8'b11110000; //  115 : 240 - 0xf0
      11'h74: dout  = 8'b11110000; //  116 : 240 - 0xf0
      11'h75: dout  = 8'b11000000; //  117 : 192 - 0xc0
      11'h76: dout  = 8'b10000000; //  118 : 128 - 0x80
      11'h77: dout  = 8'b00000000; //  119 :   0 - 0x0
      11'h78: dout  = 8'b00010000; //  120 :  16 - 0x10 -- Sprite 0xf
      11'h79: dout  = 8'b01100000; //  121 :  96 - 0x60
      11'h7A: dout  = 8'b10000000; //  122 : 128 - 0x80
      11'h7B: dout  = 8'b00000000; //  123 :   0 - 0x0
      11'h7C: dout  = 8'b01111000; //  124 : 120 - 0x78
      11'h7D: dout  = 8'b01111000; //  125 : 120 - 0x78
      11'h7E: dout  = 8'b01111110; //  126 : 126 - 0x7e
      11'h7F: dout  = 8'b01111110; //  127 : 126 - 0x7e
      11'h80: dout  = 8'b00000000; //  128 :   0 - 0x0 -- Sprite 0x10
      11'h81: dout  = 8'b00000000; //  129 :   0 - 0x0
      11'h82: dout  = 8'b00000000; //  130 :   0 - 0x0
      11'h83: dout  = 8'b00000000; //  131 :   0 - 0x0
      11'h84: dout  = 8'b00000000; //  132 :   0 - 0x0
      11'h85: dout  = 8'b00011111; //  133 :  31 - 0x1f
      11'h86: dout  = 8'b00111111; //  134 :  63 - 0x3f
      11'h87: dout  = 8'b00111111; //  135 :  63 - 0x3f
      11'h88: dout  = 8'b00000000; //  136 :   0 - 0x0 -- Sprite 0x11
      11'h89: dout  = 8'b00000000; //  137 :   0 - 0x0
      11'h8A: dout  = 8'b00100000; //  138 :  32 - 0x20
      11'h8B: dout  = 8'b01100000; //  139 :  96 - 0x60
      11'h8C: dout  = 8'b00000000; //  140 :   0 - 0x0
      11'h8D: dout  = 8'b11110000; //  141 : 240 - 0xf0
      11'h8E: dout  = 8'b11111100; //  142 : 252 - 0xfc
      11'h8F: dout  = 8'b11111110; //  143 : 254 - 0xfe
      11'h90: dout  = 8'b01111111; //  144 : 127 - 0x7f -- Sprite 0x12
      11'h91: dout  = 8'b01111111; //  145 : 127 - 0x7f
      11'h92: dout  = 8'b00111111; //  146 :  63 - 0x3f
      11'h93: dout  = 8'b00011111; //  147 :  31 - 0x1f
      11'h94: dout  = 8'b00000000; //  148 :   0 - 0x0
      11'h95: dout  = 8'b00010110; //  149 :  22 - 0x16
      11'h96: dout  = 8'b00101111; //  150 :  47 - 0x2f
      11'h97: dout  = 8'b00101111; //  151 :  47 - 0x2f
      11'h98: dout  = 8'b11111110; //  152 : 254 - 0xfe -- Sprite 0x13
      11'h99: dout  = 8'b11111100; //  153 : 252 - 0xfc
      11'h9A: dout  = 8'b11111100; //  154 : 252 - 0xfc
      11'h9B: dout  = 8'b11111000; //  155 : 248 - 0xf8
      11'h9C: dout  = 8'b11000000; //  156 : 192 - 0xc0
      11'h9D: dout  = 8'b01100000; //  157 :  96 - 0x60
      11'h9E: dout  = 8'b00100000; //  158 :  32 - 0x20
      11'h9F: dout  = 8'b00110000; //  159 :  48 - 0x30
      11'hA0: dout  = 8'b00101111; //  160 :  47 - 0x2f -- Sprite 0x14
      11'hA1: dout  = 8'b00101111; //  161 :  47 - 0x2f
      11'hA2: dout  = 8'b00101111; //  162 :  47 - 0x2f
      11'hA3: dout  = 8'b00001111; //  163 :  15 - 0xf
      11'hA4: dout  = 8'b00000111; //  164 :   7 - 0x7
      11'hA5: dout  = 8'b00000011; //  165 :   3 - 0x3
      11'hA6: dout  = 8'b00000000; //  166 :   0 - 0x0
      11'hA7: dout  = 8'b00000000; //  167 :   0 - 0x0
      11'hA8: dout  = 8'b00010000; //  168 :  16 - 0x10 -- Sprite 0x15
      11'hA9: dout  = 8'b11110000; //  169 : 240 - 0xf0
      11'hAA: dout  = 8'b11110000; //  170 : 240 - 0xf0
      11'hAB: dout  = 8'b11110000; //  171 : 240 - 0xf0
      11'hAC: dout  = 8'b11110000; //  172 : 240 - 0xf0
      11'hAD: dout  = 8'b11100000; //  173 : 224 - 0xe0
      11'hAE: dout  = 8'b11000000; //  174 : 192 - 0xc0
      11'hAF: dout  = 8'b11100000; //  175 : 224 - 0xe0
      11'hB0: dout  = 8'b00000001; //  176 :   1 - 0x1 -- Sprite 0x16
      11'hB1: dout  = 8'b00000011; //  177 :   3 - 0x3
      11'hB2: dout  = 8'b00000001; //  178 :   1 - 0x1
      11'hB3: dout  = 8'b00000100; //  179 :   4 - 0x4
      11'hB4: dout  = 8'b00000111; //  180 :   7 - 0x7
      11'hB5: dout  = 8'b00001111; //  181 :  15 - 0xf
      11'hB6: dout  = 8'b00001111; //  182 :  15 - 0xf
      11'hB7: dout  = 8'b00000011; //  183 :   3 - 0x3
      11'hB8: dout  = 8'b11111000; //  184 : 248 - 0xf8 -- Sprite 0x17
      11'hB9: dout  = 8'b11110000; //  185 : 240 - 0xf0
      11'hBA: dout  = 8'b11100000; //  186 : 224 - 0xe0
      11'hBB: dout  = 8'b01110000; //  187 : 112 - 0x70
      11'hBC: dout  = 8'b10110000; //  188 : 176 - 0xb0
      11'hBD: dout  = 8'b10000000; //  189 : 128 - 0x80
      11'hBE: dout  = 8'b11100000; //  190 : 224 - 0xe0
      11'hBF: dout  = 8'b11100000; //  191 : 224 - 0xe0
      11'hC0: dout  = 8'b00000000; //  192 :   0 - 0x0 -- Sprite 0x18
      11'hC1: dout  = 8'b00110000; //  193 :  48 - 0x30
      11'hC2: dout  = 8'b01110000; //  194 : 112 - 0x70
      11'hC3: dout  = 8'b01111111; //  195 : 127 - 0x7f
      11'hC4: dout  = 8'b11111111; //  196 : 255 - 0xff
      11'hC5: dout  = 8'b11111111; //  197 : 255 - 0xff
      11'hC6: dout  = 8'b11110111; //  198 : 247 - 0xf7
      11'hC7: dout  = 8'b11110011; //  199 : 243 - 0xf3
      11'hC8: dout  = 8'b00000000; //  200 :   0 - 0x0 -- Sprite 0x19
      11'hC9: dout  = 8'b00011000; //  201 :  24 - 0x18
      11'hCA: dout  = 8'b00010000; //  202 :  16 - 0x10
      11'hCB: dout  = 8'b00000000; //  203 :   0 - 0x0
      11'hCC: dout  = 8'b11111000; //  204 : 248 - 0xf8
      11'hCD: dout  = 8'b11111000; //  205 : 248 - 0xf8
      11'hCE: dout  = 8'b11111110; //  206 : 254 - 0xfe
      11'hCF: dout  = 8'b11111111; //  207 : 255 - 0xff
      11'hD0: dout  = 8'b11100111; //  208 : 231 - 0xe7 -- Sprite 0x1a
      11'hD1: dout  = 8'b00001111; //  209 :  15 - 0xf
      11'hD2: dout  = 8'b00001111; //  210 :  15 - 0xf
      11'hD3: dout  = 8'b00011111; //  211 :  31 - 0x1f
      11'hD4: dout  = 8'b00011111; //  212 :  31 - 0x1f
      11'hD5: dout  = 8'b00011111; //  213 :  31 - 0x1f
      11'hD6: dout  = 8'b00001111; //  214 :  15 - 0xf
      11'hD7: dout  = 8'b00000111; //  215 :   7 - 0x7
      11'hD8: dout  = 8'b11111111; //  216 : 255 - 0xff -- Sprite 0x1b
      11'hD9: dout  = 8'b11111110; //  217 : 254 - 0xfe
      11'hDA: dout  = 8'b11111100; //  218 : 252 - 0xfc
      11'hDB: dout  = 8'b11000110; //  219 : 198 - 0xc6
      11'hDC: dout  = 8'b10001110; //  220 : 142 - 0x8e
      11'hDD: dout  = 8'b11101110; //  221 : 238 - 0xee
      11'hDE: dout  = 8'b11111111; //  222 : 255 - 0xff
      11'hDF: dout  = 8'b11111111; //  223 : 255 - 0xff
      11'hE0: dout  = 8'b00000011; //  224 :   3 - 0x3 -- Sprite 0x1c
      11'hE1: dout  = 8'b00000000; //  225 :   0 - 0x0
      11'hE2: dout  = 8'b00000000; //  226 :   0 - 0x0
      11'hE3: dout  = 8'b00001110; //  227 :  14 - 0xe
      11'hE4: dout  = 8'b00000111; //  228 :   7 - 0x7
      11'hE5: dout  = 8'b00111111; //  229 :  63 - 0x3f
      11'hE6: dout  = 8'b00111111; //  230 :  63 - 0x3f
      11'hE7: dout  = 8'b00111111; //  231 :  63 - 0x3f
      11'hE8: dout  = 8'b11111111; //  232 : 255 - 0xff -- Sprite 0x1d
      11'hE9: dout  = 8'b01111111; //  233 : 127 - 0x7f
      11'hEA: dout  = 8'b00111111; //  234 :  63 - 0x3f
      11'hEB: dout  = 8'b00001110; //  235 :  14 - 0xe
      11'hEC: dout  = 8'b11000000; //  236 : 192 - 0xc0
      11'hED: dout  = 8'b11000000; //  237 : 192 - 0xc0
      11'hEE: dout  = 8'b11100000; //  238 : 224 - 0xe0
      11'hEF: dout  = 8'b11100000; //  239 : 224 - 0xe0
      11'hF0: dout  = 8'b00000000; //  240 :   0 - 0x0 -- Sprite 0x1e
      11'hF1: dout  = 8'b10000000; //  241 : 128 - 0x80
      11'hF2: dout  = 8'b11001000; //  242 : 200 - 0xc8
      11'hF3: dout  = 8'b11111110; //  243 : 254 - 0xfe
      11'hF4: dout  = 8'b01111111; //  244 : 127 - 0x7f
      11'hF5: dout  = 8'b00111111; //  245 :  63 - 0x3f
      11'hF6: dout  = 8'b00011110; //  246 :  30 - 0x1e
      11'hF7: dout  = 8'b00001110; //  247 :  14 - 0xe
      11'hF8: dout  = 8'b11100000; //  248 : 224 - 0xe0 -- Sprite 0x1f
      11'hF9: dout  = 8'b00000000; //  249 :   0 - 0x0
      11'hFA: dout  = 8'b00000000; //  250 :   0 - 0x0
      11'hFB: dout  = 8'b00000000; //  251 :   0 - 0x0
      11'hFC: dout  = 8'b00000000; //  252 :   0 - 0x0
      11'hFD: dout  = 8'b00000000; //  253 :   0 - 0x0
      11'hFE: dout  = 8'b00000000; //  254 :   0 - 0x0
      11'hFF: dout  = 8'b00000000; //  255 :   0 - 0x0
      11'h100: dout  = 8'b00000000; //  256 :   0 - 0x0 -- Sprite 0x20
      11'h101: dout  = 8'b00000000; //  257 :   0 - 0x0
      11'h102: dout  = 8'b00000000; //  258 :   0 - 0x0
      11'h103: dout  = 8'b00000000; //  259 :   0 - 0x0
      11'h104: dout  = 8'b00000000; //  260 :   0 - 0x0
      11'h105: dout  = 8'b00000000; //  261 :   0 - 0x0
      11'h106: dout  = 8'b00011111; //  262 :  31 - 0x1f
      11'h107: dout  = 8'b00111111; //  263 :  63 - 0x3f
      11'h108: dout  = 8'b00001110; //  264 :  14 - 0xe -- Sprite 0x21
      11'h109: dout  = 8'b00011111; //  265 :  31 - 0x1f
      11'h10A: dout  = 8'b00011111; //  266 :  31 - 0x1f
      11'h10B: dout  = 8'b00011111; //  267 :  31 - 0x1f
      11'h10C: dout  = 8'b00011111; //  268 :  31 - 0x1f
      11'h10D: dout  = 8'b00000011; //  269 :   3 - 0x3
      11'h10E: dout  = 8'b11111111; //  270 : 255 - 0xff
      11'h10F: dout  = 8'b11111111; //  271 : 255 - 0xff
      11'h110: dout  = 8'b00111111; //  272 :  63 - 0x3f -- Sprite 0x22
      11'h111: dout  = 8'b00111111; //  273 :  63 - 0x3f
      11'h112: dout  = 8'b01111111; //  274 : 127 - 0x7f
      11'h113: dout  = 8'b01111111; //  275 : 127 - 0x7f
      11'h114: dout  = 8'b00011111; //  276 :  31 - 0x1f
      11'h115: dout  = 8'b00000000; //  277 :   0 - 0x0
      11'h116: dout  = 8'b01111110; //  278 : 126 - 0x7e
      11'h117: dout  = 8'b11111111; //  279 : 255 - 0xff
      11'h118: dout  = 8'b11111111; //  280 : 255 - 0xff -- Sprite 0x23
      11'h119: dout  = 8'b11111111; //  281 : 255 - 0xff
      11'h11A: dout  = 8'b11111110; //  282 : 254 - 0xfe
      11'h11B: dout  = 8'b11111110; //  283 : 254 - 0xfe
      11'h11C: dout  = 8'b11111110; //  284 : 254 - 0xfe
      11'h11D: dout  = 8'b11011110; //  285 : 222 - 0xde
      11'h11E: dout  = 8'b01011100; //  286 :  92 - 0x5c
      11'h11F: dout  = 8'b01101100; //  287 : 108 - 0x6c
      11'h120: dout  = 8'b11111111; //  288 : 255 - 0xff -- Sprite 0x24
      11'h121: dout  = 8'b11111111; //  289 : 255 - 0xff
      11'h122: dout  = 8'b11111110; //  290 : 254 - 0xfe
      11'h123: dout  = 8'b11111100; //  291 : 252 - 0xfc
      11'h124: dout  = 8'b11111000; //  292 : 248 - 0xf8
      11'h125: dout  = 8'b10110000; //  293 : 176 - 0xb0
      11'h126: dout  = 8'b01100000; //  294 :  96 - 0x60
      11'h127: dout  = 8'b00000000; //  295 :   0 - 0x0
      11'h128: dout  = 8'b00101000; //  296 :  40 - 0x28 -- Sprite 0x25
      11'h129: dout  = 8'b00110000; //  297 :  48 - 0x30
      11'h12A: dout  = 8'b00011000; //  298 :  24 - 0x18
      11'h12B: dout  = 8'b01000000; //  299 :  64 - 0x40
      11'h12C: dout  = 8'b00000000; //  300 :   0 - 0x0
      11'h12D: dout  = 8'b00000001; //  301 :   1 - 0x1
      11'h12E: dout  = 8'b00000011; //  302 :   3 - 0x3
      11'h12F: dout  = 8'b00001111; //  303 :  15 - 0xf
      11'h130: dout  = 8'b00010000; //  304 :  16 - 0x10 -- Sprite 0x26
      11'h131: dout  = 8'b11101100; //  305 : 236 - 0xec
      11'h132: dout  = 8'b11100011; //  306 : 227 - 0xe3
      11'h133: dout  = 8'b11100000; //  307 : 224 - 0xe0
      11'h134: dout  = 8'b11100000; //  308 : 224 - 0xe0
      11'h135: dout  = 8'b11100000; //  309 : 224 - 0xe0
      11'h136: dout  = 8'b11000000; //  310 : 192 - 0xc0
      11'h137: dout  = 8'b10000000; //  311 : 128 - 0x80
      11'h138: dout  = 8'b00001111; //  312 :  15 - 0xf -- Sprite 0x27
      11'h139: dout  = 8'b00001111; //  313 :  15 - 0xf
      11'h13A: dout  = 8'b00001111; //  314 :  15 - 0xf
      11'h13B: dout  = 8'b00001111; //  315 :  15 - 0xf
      11'h13C: dout  = 8'b00000000; //  316 :   0 - 0x0
      11'h13D: dout  = 8'b00000000; //  317 :   0 - 0x0
      11'h13E: dout  = 8'b00000000; //  318 :   0 - 0x0
      11'h13F: dout  = 8'b00000000; //  319 :   0 - 0x0
      11'h140: dout  = 8'b00011111; //  320 :  31 - 0x1f -- Sprite 0x28
      11'h141: dout  = 8'b00111111; //  321 :  63 - 0x3f
      11'h142: dout  = 8'b00111111; //  322 :  63 - 0x3f
      11'h143: dout  = 8'b00011111; //  323 :  31 - 0x1f
      11'h144: dout  = 8'b00000111; //  324 :   7 - 0x7
      11'h145: dout  = 8'b00001001; //  325 :   9 - 0x9
      11'h146: dout  = 8'b00010011; //  326 :  19 - 0x13
      11'h147: dout  = 8'b00010111; //  327 :  23 - 0x17
      11'h148: dout  = 8'b11111111; //  328 : 255 - 0xff -- Sprite 0x29
      11'h149: dout  = 8'b11111111; //  329 : 255 - 0xff
      11'h14A: dout  = 8'b11111110; //  330 : 254 - 0xfe
      11'h14B: dout  = 8'b11111111; //  331 : 255 - 0xff
      11'h14C: dout  = 8'b11111110; //  332 : 254 - 0xfe
      11'h14D: dout  = 8'b11111100; //  333 : 252 - 0xfc
      11'h14E: dout  = 8'b11111000; //  334 : 248 - 0xf8
      11'h14F: dout  = 8'b11100000; //  335 : 224 - 0xe0
      11'h150: dout  = 8'b00010111; //  336 :  23 - 0x17 -- Sprite 0x2a
      11'h151: dout  = 8'b00010111; //  337 :  23 - 0x17
      11'h152: dout  = 8'b00000011; //  338 :   3 - 0x3
      11'h153: dout  = 8'b00000000; //  339 :   0 - 0x0
      11'h154: dout  = 8'b00000000; //  340 :   0 - 0x0
      11'h155: dout  = 8'b00000000; //  341 :   0 - 0x0
      11'h156: dout  = 8'b00000000; //  342 :   0 - 0x0
      11'h157: dout  = 8'b00000000; //  343 :   0 - 0x0
      11'h158: dout  = 8'b11010000; //  344 : 208 - 0xd0 -- Sprite 0x2b
      11'h159: dout  = 8'b10010000; //  345 : 144 - 0x90
      11'h15A: dout  = 8'b00011000; //  346 :  24 - 0x18
      11'h15B: dout  = 8'b00001000; //  347 :   8 - 0x8
      11'h15C: dout  = 8'b01000000; //  348 :  64 - 0x40
      11'h15D: dout  = 8'b00000000; //  349 :   0 - 0x0
      11'h15E: dout  = 8'b00000000; //  350 :   0 - 0x0
      11'h15F: dout  = 8'b00000000; //  351 :   0 - 0x0
      11'h160: dout  = 8'b00110000; //  352 :  48 - 0x30 -- Sprite 0x2c
      11'h161: dout  = 8'b11110000; //  353 : 240 - 0xf0
      11'h162: dout  = 8'b11110000; //  354 : 240 - 0xf0
      11'h163: dout  = 8'b11110001; //  355 : 241 - 0xf1
      11'h164: dout  = 8'b11110110; //  356 : 246 - 0xf6
      11'h165: dout  = 8'b11000110; //  357 : 198 - 0xc6
      11'h166: dout  = 8'b10000100; //  358 : 132 - 0x84
      11'h167: dout  = 8'b00000000; //  359 :   0 - 0x0
      11'h168: dout  = 8'b00000000; //  360 :   0 - 0x0 -- Sprite 0x2d
      11'h169: dout  = 8'b00000000; //  361 :   0 - 0x0
      11'h16A: dout  = 8'b00000000; //  362 :   0 - 0x0
      11'h16B: dout  = 8'b00000000; //  363 :   0 - 0x0
      11'h16C: dout  = 8'b00000000; //  364 :   0 - 0x0
      11'h16D: dout  = 8'b00000000; //  365 :   0 - 0x0
      11'h16E: dout  = 8'b00000000; //  366 :   0 - 0x0
      11'h16F: dout  = 8'b00000000; //  367 :   0 - 0x0
      11'h170: dout  = 8'b00011111; //  368 :  31 - 0x1f -- Sprite 0x2e
      11'h171: dout  = 8'b00011111; //  369 :  31 - 0x1f
      11'h172: dout  = 8'b00111111; //  370 :  63 - 0x3f
      11'h173: dout  = 8'b00111110; //  371 :  62 - 0x3e
      11'h174: dout  = 8'b01111100; //  372 : 124 - 0x7c
      11'h175: dout  = 8'b01111000; //  373 : 120 - 0x78
      11'h176: dout  = 8'b11110000; //  374 : 240 - 0xf0
      11'h177: dout  = 8'b11100000; //  375 : 224 - 0xe0
      11'h178: dout  = 8'b10110000; //  376 : 176 - 0xb0 -- Sprite 0x2f
      11'h179: dout  = 8'b10010000; //  377 : 144 - 0x90
      11'h17A: dout  = 8'b00011000; //  378 :  24 - 0x18
      11'h17B: dout  = 8'b00001000; //  379 :   8 - 0x8
      11'h17C: dout  = 8'b01000000; //  380 :  64 - 0x40
      11'h17D: dout  = 8'b00000000; //  381 :   0 - 0x0
      11'h17E: dout  = 8'b00000000; //  382 :   0 - 0x0
      11'h17F: dout  = 8'b00000000; //  383 :   0 - 0x0
      11'h180: dout  = 8'b11000000; //  384 : 192 - 0xc0 -- Sprite 0x30
      11'h181: dout  = 8'b11100000; //  385 : 224 - 0xe0
      11'h182: dout  = 8'b11111100; //  386 : 252 - 0xfc
      11'h183: dout  = 8'b11111110; //  387 : 254 - 0xfe
      11'h184: dout  = 8'b11111111; //  388 : 255 - 0xff
      11'h185: dout  = 8'b01111111; //  389 : 127 - 0x7f
      11'h186: dout  = 8'b00000011; //  390 :   3 - 0x3
      11'h187: dout  = 8'b00000000; //  391 :   0 - 0x0
      11'h188: dout  = 8'b00000000; //  392 :   0 - 0x0 -- Sprite 0x31
      11'h189: dout  = 8'b00000000; //  393 :   0 - 0x0
      11'h18A: dout  = 8'b00010000; //  394 :  16 - 0x10
      11'h18B: dout  = 8'b00111000; //  395 :  56 - 0x38
      11'h18C: dout  = 8'b00111110; //  396 :  62 - 0x3e
      11'h18D: dout  = 8'b00111100; //  397 :  60 - 0x3c
      11'h18E: dout  = 8'b00111000; //  398 :  56 - 0x38
      11'h18F: dout  = 8'b00011000; //  399 :  24 - 0x18
      11'h190: dout  = 8'b00000000; //  400 :   0 - 0x0 -- Sprite 0x32
      11'h191: dout  = 8'b00000000; //  401 :   0 - 0x0
      11'h192: dout  = 8'b00000000; //  402 :   0 - 0x0
      11'h193: dout  = 8'b00000111; //  403 :   7 - 0x7
      11'h194: dout  = 8'b00001111; //  404 :  15 - 0xf
      11'h195: dout  = 8'b00001111; //  405 :  15 - 0xf
      11'h196: dout  = 8'b00001111; //  406 :  15 - 0xf
      11'h197: dout  = 8'b00000011; //  407 :   3 - 0x3
      11'h198: dout  = 8'b00000000; //  408 :   0 - 0x0 -- Sprite 0x33
      11'h199: dout  = 8'b00000000; //  409 :   0 - 0x0
      11'h19A: dout  = 8'b00000000; //  410 :   0 - 0x0
      11'h19B: dout  = 8'b11110000; //  411 : 240 - 0xf0
      11'h19C: dout  = 8'b11111100; //  412 : 252 - 0xfc
      11'h19D: dout  = 8'b11111110; //  413 : 254 - 0xfe
      11'h19E: dout  = 8'b11111100; //  414 : 252 - 0xfc
      11'h19F: dout  = 8'b11111000; //  415 : 248 - 0xf8
      11'h1A0: dout  = 8'b00000111; //  416 :   7 - 0x7 -- Sprite 0x34
      11'h1A1: dout  = 8'b00001111; //  417 :  15 - 0xf
      11'h1A2: dout  = 8'b00011011; //  418 :  27 - 0x1b
      11'h1A3: dout  = 8'b00011000; //  419 :  24 - 0x18
      11'h1A4: dout  = 8'b00010000; //  420 :  16 - 0x10
      11'h1A5: dout  = 8'b00110000; //  421 :  48 - 0x30
      11'h1A6: dout  = 8'b00100001; //  422 :  33 - 0x21
      11'h1A7: dout  = 8'b00000001; //  423 :   1 - 0x1
      11'h1A8: dout  = 8'b10101000; //  424 : 168 - 0xa8 -- Sprite 0x35
      11'h1A9: dout  = 8'b11111100; //  425 : 252 - 0xfc
      11'h1AA: dout  = 8'b11111000; //  426 : 248 - 0xf8
      11'h1AB: dout  = 8'b00000000; //  427 :   0 - 0x0
      11'h1AC: dout  = 8'b00000000; //  428 :   0 - 0x0
      11'h1AD: dout  = 8'b00000000; //  429 :   0 - 0x0
      11'h1AE: dout  = 8'b11000000; //  430 : 192 - 0xc0
      11'h1AF: dout  = 8'b11100000; //  431 : 224 - 0xe0
      11'h1B0: dout  = 8'b00000000; //  432 :   0 - 0x0 -- Sprite 0x36
      11'h1B1: dout  = 8'b00000000; //  433 :   0 - 0x0
      11'h1B2: dout  = 8'b00001111; //  434 :  15 - 0xf
      11'h1B3: dout  = 8'b00011111; //  435 :  31 - 0x1f
      11'h1B4: dout  = 8'b00011111; //  436 :  31 - 0x1f
      11'h1B5: dout  = 8'b00011111; //  437 :  31 - 0x1f
      11'h1B6: dout  = 8'b00000111; //  438 :   7 - 0x7
      11'h1B7: dout  = 8'b00111100; //  439 :  60 - 0x3c
      11'h1B8: dout  = 8'b00000000; //  440 :   0 - 0x0 -- Sprite 0x37
      11'h1B9: dout  = 8'b00000000; //  441 :   0 - 0x0
      11'h1BA: dout  = 8'b11100000; //  442 : 224 - 0xe0
      11'h1BB: dout  = 8'b11111000; //  443 : 248 - 0xf8
      11'h1BC: dout  = 8'b11111100; //  444 : 252 - 0xfc
      11'h1BD: dout  = 8'b11111000; //  445 : 248 - 0xf8
      11'h1BE: dout  = 8'b11110000; //  446 : 240 - 0xf0
      11'h1BF: dout  = 8'b11000000; //  447 : 192 - 0xc0
      11'h1C0: dout  = 8'b11111100; //  448 : 252 - 0xfc -- Sprite 0x38
      11'h1C1: dout  = 8'b11101101; //  449 : 237 - 0xed
      11'h1C2: dout  = 8'b11000000; //  450 : 192 - 0xc0
      11'h1C3: dout  = 8'b00000000; //  451 :   0 - 0x0
      11'h1C4: dout  = 8'b00000000; //  452 :   0 - 0x0
      11'h1C5: dout  = 8'b01100000; //  453 :  96 - 0x60
      11'h1C6: dout  = 8'b01110000; //  454 : 112 - 0x70
      11'h1C7: dout  = 8'b00111000; //  455 :  56 - 0x38
      11'h1C8: dout  = 8'b01111110; //  456 : 126 - 0x7e -- Sprite 0x39
      11'h1C9: dout  = 8'b00011110; //  457 :  30 - 0x1e
      11'h1CA: dout  = 8'b00000100; //  458 :   4 - 0x4
      11'h1CB: dout  = 8'b00001100; //  459 :  12 - 0xc
      11'h1CC: dout  = 8'b00001100; //  460 :  12 - 0xc
      11'h1CD: dout  = 8'b00001100; //  461 :  12 - 0xc
      11'h1CE: dout  = 8'b00000000; //  462 :   0 - 0x0
      11'h1CF: dout  = 8'b00000000; //  463 :   0 - 0x0
      11'h1D0: dout  = 8'b00000000; //  464 :   0 - 0x0 -- Sprite 0x3a
      11'h1D1: dout  = 8'b00000000; //  465 :   0 - 0x0
      11'h1D2: dout  = 8'b00001111; //  466 :  15 - 0xf
      11'h1D3: dout  = 8'b00011111; //  467 :  31 - 0x1f
      11'h1D4: dout  = 8'b00011111; //  468 :  31 - 0x1f
      11'h1D5: dout  = 8'b00011111; //  469 :  31 - 0x1f
      11'h1D6: dout  = 8'b00000111; //  470 :   7 - 0x7
      11'h1D7: dout  = 8'b00001101; //  471 :  13 - 0xd
      11'h1D8: dout  = 8'b00011110; //  472 :  30 - 0x1e -- Sprite 0x3b
      11'h1D9: dout  = 8'b00011100; //  473 :  28 - 0x1c
      11'h1DA: dout  = 8'b00011110; //  474 :  30 - 0x1e
      11'h1DB: dout  = 8'b00001111; //  475 :  15 - 0xf
      11'h1DC: dout  = 8'b00000111; //  476 :   7 - 0x7
      11'h1DD: dout  = 8'b00000000; //  477 :   0 - 0x0
      11'h1DE: dout  = 8'b00000111; //  478 :   7 - 0x7
      11'h1DF: dout  = 8'b00000111; //  479 :   7 - 0x7
      11'h1E0: dout  = 8'b01100000; //  480 :  96 - 0x60 -- Sprite 0x3c
      11'h1E1: dout  = 8'b10010000; //  481 : 144 - 0x90
      11'h1E2: dout  = 8'b00000000; //  482 :   0 - 0x0
      11'h1E3: dout  = 8'b10000000; //  483 : 128 - 0x80
      11'h1E4: dout  = 8'b00000000; //  484 :   0 - 0x0
      11'h1E5: dout  = 8'b11100000; //  485 : 224 - 0xe0
      11'h1E6: dout  = 8'b11110000; //  486 : 240 - 0xf0
      11'h1E7: dout  = 8'b10000000; //  487 : 128 - 0x80
      11'h1E8: dout  = 8'b00000000; //  488 :   0 - 0x0 -- Sprite 0x3d
      11'h1E9: dout  = 8'b00010000; //  489 :  16 - 0x10
      11'h1EA: dout  = 8'b00111111; //  490 :  63 - 0x3f
      11'h1EB: dout  = 8'b01111111; //  491 : 127 - 0x7f
      11'h1EC: dout  = 8'b01111111; //  492 : 127 - 0x7f
      11'h1ED: dout  = 8'b00111111; //  493 :  63 - 0x3f
      11'h1EE: dout  = 8'b00000011; //  494 :   3 - 0x3
      11'h1EF: dout  = 8'b00001111; //  495 :  15 - 0xf
      11'h1F0: dout  = 8'b00000000; //  496 :   0 - 0x0 -- Sprite 0x3e
      11'h1F1: dout  = 8'b00000000; //  497 :   0 - 0x0
      11'h1F2: dout  = 8'b11100000; //  498 : 224 - 0xe0
      11'h1F3: dout  = 8'b11111000; //  499 : 248 - 0xf8
      11'h1F4: dout  = 8'b11111100; //  500 : 252 - 0xfc
      11'h1F5: dout  = 8'b11111000; //  501 : 248 - 0xf8
      11'h1F6: dout  = 8'b10110000; //  502 : 176 - 0xb0
      11'h1F7: dout  = 8'b00111000; //  503 :  56 - 0x38
      11'h1F8: dout  = 8'b00011111; //  504 :  31 - 0x1f -- Sprite 0x3f
      11'h1F9: dout  = 8'b00000111; //  505 :   7 - 0x7
      11'h1FA: dout  = 8'b00000000; //  506 :   0 - 0x0
      11'h1FB: dout  = 8'b00001110; //  507 :  14 - 0xe
      11'h1FC: dout  = 8'b00001111; //  508 :  15 - 0xf
      11'h1FD: dout  = 8'b01010011; //  509 :  83 - 0x53
      11'h1FE: dout  = 8'b01111100; //  510 : 124 - 0x7c
      11'h1FF: dout  = 8'b00111100; //  511 :  60 - 0x3c
      11'h200: dout  = 8'b11111000; //  512 : 248 - 0xf8 -- Sprite 0x40
      11'h201: dout  = 8'b11111000; //  513 : 248 - 0xf8
      11'h202: dout  = 8'b11110000; //  514 : 240 - 0xf0
      11'h203: dout  = 8'b00000000; //  515 :   0 - 0x0
      11'h204: dout  = 8'b00000000; //  516 :   0 - 0x0
      11'h205: dout  = 8'b10000000; //  517 : 128 - 0x80
      11'h206: dout  = 8'b00000000; //  518 :   0 - 0x0
      11'h207: dout  = 8'b00000000; //  519 :   0 - 0x0
      11'h208: dout  = 8'b00000111; //  520 :   7 - 0x7 -- Sprite 0x41
      11'h209: dout  = 8'b00000111; //  521 :   7 - 0x7
      11'h20A: dout  = 8'b00000011; //  522 :   3 - 0x3
      11'h20B: dout  = 8'b11110111; //  523 : 247 - 0xf7
      11'h20C: dout  = 8'b11111111; //  524 : 255 - 0xff
      11'h20D: dout  = 8'b11111111; //  525 : 255 - 0xff
      11'h20E: dout  = 8'b11111110; //  526 : 254 - 0xfe
      11'h20F: dout  = 8'b11111100; //  527 : 252 - 0xfc
      11'h210: dout  = 8'b00111110; //  528 :  62 - 0x3e -- Sprite 0x42
      11'h211: dout  = 8'b01111111; //  529 : 127 - 0x7f
      11'h212: dout  = 8'b11111111; //  530 : 255 - 0xff
      11'h213: dout  = 8'b11100010; //  531 : 226 - 0xe2
      11'h214: dout  = 8'b01010000; //  532 :  80 - 0x50
      11'h215: dout  = 8'b00111000; //  533 :  56 - 0x38
      11'h216: dout  = 8'b01110000; //  534 : 112 - 0x70
      11'h217: dout  = 8'b01000000; //  535 :  64 - 0x40
      11'h218: dout  = 8'b11101000; //  536 : 232 - 0xe8 -- Sprite 0x43
      11'h219: dout  = 8'b01110001; //  537 : 113 - 0x71
      11'h21A: dout  = 8'b00000001; //  538 :   1 - 0x1
      11'h21B: dout  = 8'b01001011; //  539 :  75 - 0x4b
      11'h21C: dout  = 8'b00000011; //  540 :   3 - 0x3
      11'h21D: dout  = 8'b00000011; //  541 :   3 - 0x3
      11'h21E: dout  = 8'b00000000; //  542 :   0 - 0x0
      11'h21F: dout  = 8'b00000000; //  543 :   0 - 0x0
      11'h220: dout  = 8'b00000101; //  544 :   5 - 0x5 -- Sprite 0x44
      11'h221: dout  = 8'b00000011; //  545 :   3 - 0x3
      11'h222: dout  = 8'b00000001; //  546 :   1 - 0x1
      11'h223: dout  = 8'b00110000; //  547 :  48 - 0x30
      11'h224: dout  = 8'b00110000; //  548 :  48 - 0x30
      11'h225: dout  = 8'b00110000; //  549 :  48 - 0x30
      11'h226: dout  = 8'b00100110; //  550 :  38 - 0x26
      11'h227: dout  = 8'b00000100; //  551 :   4 - 0x4
      11'h228: dout  = 8'b11111110; //  552 : 254 - 0xfe -- Sprite 0x45
      11'h229: dout  = 8'b11111100; //  553 : 252 - 0xfc
      11'h22A: dout  = 8'b11100000; //  554 : 224 - 0xe0
      11'h22B: dout  = 8'b00000000; //  555 :   0 - 0x0
      11'h22C: dout  = 8'b00000000; //  556 :   0 - 0x0
      11'h22D: dout  = 8'b00000000; //  557 :   0 - 0x0
      11'h22E: dout  = 8'b00000000; //  558 :   0 - 0x0
      11'h22F: dout  = 8'b00000000; //  559 :   0 - 0x0
      11'h230: dout  = 8'b00000101; //  560 :   5 - 0x5 -- Sprite 0x46
      11'h231: dout  = 8'b00000011; //  561 :   3 - 0x3
      11'h232: dout  = 8'b00000001; //  562 :   1 - 0x1
      11'h233: dout  = 8'b00010000; //  563 :  16 - 0x10
      11'h234: dout  = 8'b00110000; //  564 :  48 - 0x30
      11'h235: dout  = 8'b00001100; //  565 :  12 - 0xc
      11'h236: dout  = 8'b00011100; //  566 :  28 - 0x1c
      11'h237: dout  = 8'b00011000; //  567 :  24 - 0x18
      11'h238: dout  = 8'b11000000; //  568 : 192 - 0xc0 -- Sprite 0x47
      11'h239: dout  = 8'b11100000; //  569 : 224 - 0xe0
      11'h23A: dout  = 8'b11110000; //  570 : 240 - 0xf0
      11'h23B: dout  = 8'b01111000; //  571 : 120 - 0x78
      11'h23C: dout  = 8'b00011000; //  572 :  24 - 0x18
      11'h23D: dout  = 8'b00001000; //  573 :   8 - 0x8
      11'h23E: dout  = 8'b00000000; //  574 :   0 - 0x0
      11'h23F: dout  = 8'b00000000; //  575 :   0 - 0x0
      11'h240: dout  = 8'b00000111; //  576 :   7 - 0x7 -- Sprite 0x48
      11'h241: dout  = 8'b00001111; //  577 :  15 - 0xf
      11'h242: dout  = 8'b00111110; //  578 :  62 - 0x3e
      11'h243: dout  = 8'b01111100; //  579 : 124 - 0x7c
      11'h244: dout  = 8'b00110000; //  580 :  48 - 0x30
      11'h245: dout  = 8'b00001100; //  581 :  12 - 0xc
      11'h246: dout  = 8'b00011100; //  582 :  28 - 0x1c
      11'h247: dout  = 8'b00011000; //  583 :  24 - 0x18
      11'h248: dout  = 8'b01100000; //  584 :  96 - 0x60 -- Sprite 0x49
      11'h249: dout  = 8'b01100000; //  585 :  96 - 0x60
      11'h24A: dout  = 8'b01100000; //  586 :  96 - 0x60
      11'h24B: dout  = 8'b10000000; //  587 : 128 - 0x80
      11'h24C: dout  = 8'b00000000; //  588 :   0 - 0x0
      11'h24D: dout  = 8'b00000000; //  589 :   0 - 0x0
      11'h24E: dout  = 8'b00000000; //  590 :   0 - 0x0
      11'h24F: dout  = 8'b00000000; //  591 :   0 - 0x0
      11'h250: dout  = 8'b01110011; //  592 : 115 - 0x73 -- Sprite 0x4a
      11'h251: dout  = 8'b11110011; //  593 : 243 - 0xf3
      11'h252: dout  = 8'b11110000; //  594 : 240 - 0xf0
      11'h253: dout  = 8'b11110100; //  595 : 244 - 0xf4
      11'h254: dout  = 8'b11110000; //  596 : 240 - 0xf0
      11'h255: dout  = 8'b11110000; //  597 : 240 - 0xf0
      11'h256: dout  = 8'b01110000; //  598 : 112 - 0x70
      11'h257: dout  = 8'b01100000; //  599 :  96 - 0x60
      11'h258: dout  = 8'b00000000; //  600 :   0 - 0x0 -- Sprite 0x4b
      11'h259: dout  = 8'b00000000; //  601 :   0 - 0x0
      11'h25A: dout  = 8'b00000000; //  602 :   0 - 0x0
      11'h25B: dout  = 8'b00000000; //  603 :   0 - 0x0
      11'h25C: dout  = 8'b00111100; //  604 :  60 - 0x3c
      11'h25D: dout  = 8'b00111100; //  605 :  60 - 0x3c
      11'h25E: dout  = 8'b11111100; //  606 : 252 - 0xfc
      11'h25F: dout  = 8'b11111100; //  607 : 252 - 0xfc
      11'h260: dout  = 8'b01111111; //  608 : 127 - 0x7f -- Sprite 0x4c
      11'h261: dout  = 8'b01111111; //  609 : 127 - 0x7f
      11'h262: dout  = 8'b00011111; //  610 :  31 - 0x1f
      11'h263: dout  = 8'b00000111; //  611 :   7 - 0x7
      11'h264: dout  = 8'b00001011; //  612 :  11 - 0xb
      11'h265: dout  = 8'b00011011; //  613 :  27 - 0x1b
      11'h266: dout  = 8'b00111011; //  614 :  59 - 0x3b
      11'h267: dout  = 8'b01111011; //  615 : 123 - 0x7b
      11'h268: dout  = 8'b11111100; //  616 : 252 - 0xfc -- Sprite 0x4d
      11'h269: dout  = 8'b11111100; //  617 : 252 - 0xfc
      11'h26A: dout  = 8'b11111000; //  618 : 248 - 0xf8
      11'h26B: dout  = 8'b11100000; //  619 : 224 - 0xe0
      11'h26C: dout  = 8'b11010000; //  620 : 208 - 0xd0
      11'h26D: dout  = 8'b11011000; //  621 : 216 - 0xd8
      11'h26E: dout  = 8'b11011100; //  622 : 220 - 0xdc
      11'h26F: dout  = 8'b11011110; //  623 : 222 - 0xde
      11'h270: dout  = 8'b11000100; //  624 : 196 - 0xc4 -- Sprite 0x4e
      11'h271: dout  = 8'b11100000; //  625 : 224 - 0xe0
      11'h272: dout  = 8'b11100000; //  626 : 224 - 0xe0
      11'h273: dout  = 8'b01000000; //  627 :  64 - 0x40
      11'h274: dout  = 8'b00000000; //  628 :   0 - 0x0
      11'h275: dout  = 8'b00111100; //  629 :  60 - 0x3c
      11'h276: dout  = 8'b00111100; //  630 :  60 - 0x3c
      11'h277: dout  = 8'b01111100; //  631 : 124 - 0x7c
      11'h278: dout  = 8'b00011101; //  632 :  29 - 0x1d -- Sprite 0x4f
      11'h279: dout  = 8'b00111100; //  633 :  60 - 0x3c
      11'h27A: dout  = 8'b00111010; //  634 :  58 - 0x3a
      11'h27B: dout  = 8'b00111000; //  635 :  56 - 0x38
      11'h27C: dout  = 8'b00110000; //  636 :  48 - 0x30
      11'h27D: dout  = 8'b00000000; //  637 :   0 - 0x0
      11'h27E: dout  = 8'b00011100; //  638 :  28 - 0x1c
      11'h27F: dout  = 8'b00111100; //  639 :  60 - 0x3c
      11'h280: dout  = 8'b00100010; //  640 :  34 - 0x22 -- Sprite 0x50
      11'h281: dout  = 8'b01010101; //  641 :  85 - 0x55
      11'h282: dout  = 8'b01010101; //  642 :  85 - 0x55
      11'h283: dout  = 8'b01010101; //  643 :  85 - 0x55
      11'h284: dout  = 8'b01010101; //  644 :  85 - 0x55
      11'h285: dout  = 8'b01010101; //  645 :  85 - 0x55
      11'h286: dout  = 8'b01110111; //  646 : 119 - 0x77
      11'h287: dout  = 8'b00100010; //  647 :  34 - 0x22
      11'h288: dout  = 8'b00000000; //  648 :   0 - 0x0 -- Sprite 0x51
      11'h289: dout  = 8'b00000000; //  649 :   0 - 0x0
      11'h28A: dout  = 8'b00000000; //  650 :   0 - 0x0
      11'h28B: dout  = 8'b00000000; //  651 :   0 - 0x0
      11'h28C: dout  = 8'b00000000; //  652 :   0 - 0x0
      11'h28D: dout  = 8'b00000000; //  653 :   0 - 0x0
      11'h28E: dout  = 8'b00000000; //  654 :   0 - 0x0
      11'h28F: dout  = 8'b00000000; //  655 :   0 - 0x0
      11'h290: dout  = 8'b00000000; //  656 :   0 - 0x0 -- Sprite 0x52
      11'h291: dout  = 8'b00000000; //  657 :   0 - 0x0
      11'h292: dout  = 8'b11001111; //  658 : 207 - 0xcf
      11'h293: dout  = 8'b00000111; //  659 :   7 - 0x7
      11'h294: dout  = 8'b01111111; //  660 : 127 - 0x7f
      11'h295: dout  = 8'b00000000; //  661 :   0 - 0x0
      11'h296: dout  = 8'b00000000; //  662 :   0 - 0x0
      11'h297: dout  = 8'b00000000; //  663 :   0 - 0x0
      11'h298: dout  = 8'b00000000; //  664 :   0 - 0x0 -- Sprite 0x53
      11'h299: dout  = 8'b00000000; //  665 :   0 - 0x0
      11'h29A: dout  = 8'b00111100; //  666 :  60 - 0x3c
      11'h29B: dout  = 8'b11111100; //  667 : 252 - 0xfc
      11'h29C: dout  = 8'b11111110; //  668 : 254 - 0xfe
      11'h29D: dout  = 8'b11100000; //  669 : 224 - 0xe0
      11'h29E: dout  = 8'b00000000; //  670 :   0 - 0x0
      11'h29F: dout  = 8'b00000000; //  671 :   0 - 0x0
      11'h2A0: dout  = 8'b01000000; //  672 :  64 - 0x40 -- Sprite 0x54
      11'h2A1: dout  = 8'b11100000; //  673 : 224 - 0xe0
      11'h2A2: dout  = 8'b01000000; //  674 :  64 - 0x40
      11'h2A3: dout  = 8'b00111111; //  675 :  63 - 0x3f
      11'h2A4: dout  = 8'b00111110; //  676 :  62 - 0x3e
      11'h2A5: dout  = 8'b00111110; //  677 :  62 - 0x3e
      11'h2A6: dout  = 8'b00110000; //  678 :  48 - 0x30
      11'h2A7: dout  = 8'b00111000; //  679 :  56 - 0x38
      11'h2A8: dout  = 8'b00000000; //  680 :   0 - 0x0 -- Sprite 0x55
      11'h2A9: dout  = 8'b00000000; //  681 :   0 - 0x0
      11'h2AA: dout  = 8'b00000000; //  682 :   0 - 0x0
      11'h2AB: dout  = 8'b11111000; //  683 : 248 - 0xf8
      11'h2AC: dout  = 8'b11111000; //  684 : 248 - 0xf8
      11'h2AD: dout  = 8'b11111000; //  685 : 248 - 0xf8
      11'h2AE: dout  = 8'b00011000; //  686 :  24 - 0x18
      11'h2AF: dout  = 8'b00111000; //  687 :  56 - 0x38
      11'h2B0: dout  = 8'b00111100; //  688 :  60 - 0x3c -- Sprite 0x56
      11'h2B1: dout  = 8'b00111001; //  689 :  57 - 0x39
      11'h2B2: dout  = 8'b00111011; //  690 :  59 - 0x3b
      11'h2B3: dout  = 8'b00111111; //  691 :  63 - 0x3f
      11'h2B4: dout  = 8'b00000000; //  692 :   0 - 0x0
      11'h2B5: dout  = 8'b00000000; //  693 :   0 - 0x0
      11'h2B6: dout  = 8'b00000000; //  694 :   0 - 0x0
      11'h2B7: dout  = 8'b00000000; //  695 :   0 - 0x0
      11'h2B8: dout  = 8'b01111000; //  696 : 120 - 0x78 -- Sprite 0x57
      11'h2B9: dout  = 8'b00111000; //  697 :  56 - 0x38
      11'h2BA: dout  = 8'b10111000; //  698 : 184 - 0xb8
      11'h2BB: dout  = 8'b11111000; //  699 : 248 - 0xf8
      11'h2BC: dout  = 8'b00000000; //  700 :   0 - 0x0
      11'h2BD: dout  = 8'b00000000; //  701 :   0 - 0x0
      11'h2BE: dout  = 8'b00000000; //  702 :   0 - 0x0
      11'h2BF: dout  = 8'b00000000; //  703 :   0 - 0x0
      11'h2C0: dout  = 8'b00111111; //  704 :  63 - 0x3f -- Sprite 0x58
      11'h2C1: dout  = 8'b00111111; //  705 :  63 - 0x3f
      11'h2C2: dout  = 8'b00001111; //  706 :  15 - 0xf
      11'h2C3: dout  = 8'b01110111; //  707 : 119 - 0x77
      11'h2C4: dout  = 8'b01110111; //  708 : 119 - 0x77
      11'h2C5: dout  = 8'b11110111; //  709 : 247 - 0xf7
      11'h2C6: dout  = 8'b11110111; //  710 : 247 - 0xf7
      11'h2C7: dout  = 8'b11110111; //  711 : 247 - 0xf7
      11'h2C8: dout  = 8'b11111111; //  712 : 255 - 0xff -- Sprite 0x59
      11'h2C9: dout  = 8'b11111110; //  713 : 254 - 0xfe
      11'h2CA: dout  = 8'b11111110; //  714 : 254 - 0xfe
      11'h2CB: dout  = 8'b11111110; //  715 : 254 - 0xfe
      11'h2CC: dout  = 8'b11111010; //  716 : 250 - 0xfa
      11'h2CD: dout  = 8'b11111010; //  717 : 250 - 0xfa
      11'h2CE: dout  = 8'b11110011; //  718 : 243 - 0xf3
      11'h2CF: dout  = 8'b11100111; //  719 : 231 - 0xe7
      11'h2D0: dout  = 8'b11110000; //  720 : 240 - 0xf0 -- Sprite 0x5a
      11'h2D1: dout  = 8'b11111000; //  721 : 248 - 0xf8
      11'h2D2: dout  = 8'b11111100; //  722 : 252 - 0xfc
      11'h2D3: dout  = 8'b01111100; //  723 : 124 - 0x7c
      11'h2D4: dout  = 8'b01111000; //  724 : 120 - 0x78
      11'h2D5: dout  = 8'b00111000; //  725 :  56 - 0x38
      11'h2D6: dout  = 8'b00111100; //  726 :  60 - 0x3c
      11'h2D7: dout  = 8'b11111100; //  727 : 252 - 0xfc
      11'h2D8: dout  = 8'b11111111; //  728 : 255 - 0xff -- Sprite 0x5b
      11'h2D9: dout  = 8'b00000000; //  729 :   0 - 0x0
      11'h2DA: dout  = 8'b11000011; //  730 : 195 - 0xc3
      11'h2DB: dout  = 8'b10000001; //  731 : 129 - 0x81
      11'h2DC: dout  = 8'b10000001; //  732 : 129 - 0x81
      11'h2DD: dout  = 8'b11000011; //  733 : 195 - 0xc3
      11'h2DE: dout  = 8'b11111111; //  734 : 255 - 0xff
      11'h2DF: dout  = 8'b00000000; //  735 :   0 - 0x0
      11'h2E0: dout  = 8'b00000000; //  736 :   0 - 0x0 -- Sprite 0x5c
      11'h2E1: dout  = 8'b00000000; //  737 :   0 - 0x0
      11'h2E2: dout  = 8'b00000000; //  738 :   0 - 0x0
      11'h2E3: dout  = 8'b00000000; //  739 :   0 - 0x0
      11'h2E4: dout  = 8'b00000000; //  740 :   0 - 0x0
      11'h2E5: dout  = 8'b00000000; //  741 :   0 - 0x0
      11'h2E6: dout  = 8'b00000000; //  742 :   0 - 0x0
      11'h2E7: dout  = 8'b00000000; //  743 :   0 - 0x0
      11'h2E8: dout  = 8'b00000000; //  744 :   0 - 0x0 -- Sprite 0x5d
      11'h2E9: dout  = 8'b00001011; //  745 :  11 - 0xb
      11'h2EA: dout  = 8'b00011111; //  746 :  31 - 0x1f
      11'h2EB: dout  = 8'b00011111; //  747 :  31 - 0x1f
      11'h2EC: dout  = 8'b00011110; //  748 :  30 - 0x1e
      11'h2ED: dout  = 8'b00111110; //  749 :  62 - 0x3e
      11'h2EE: dout  = 8'b00001100; //  750 :  12 - 0xc
      11'h2EF: dout  = 8'b00000100; //  751 :   4 - 0x4
      11'h2F0: dout  = 8'b00000000; //  752 :   0 - 0x0 -- Sprite 0x5e
      11'h2F1: dout  = 8'b00000000; //  753 :   0 - 0x0
      11'h2F2: dout  = 8'b00000000; //  754 :   0 - 0x0
      11'h2F3: dout  = 8'b00000000; //  755 :   0 - 0x0
      11'h2F4: dout  = 8'b00000000; //  756 :   0 - 0x0
      11'h2F5: dout  = 8'b00000000; //  757 :   0 - 0x0
      11'h2F6: dout  = 8'b00000000; //  758 :   0 - 0x0
      11'h2F7: dout  = 8'b00000000; //  759 :   0 - 0x0
      11'h2F8: dout  = 8'b00000011; //  760 :   3 - 0x3 -- Sprite 0x5f
      11'h2F9: dout  = 8'b00001111; //  761 :  15 - 0xf
      11'h2FA: dout  = 8'b00001111; //  762 :  15 - 0xf
      11'h2FB: dout  = 8'b00001111; //  763 :  15 - 0xf
      11'h2FC: dout  = 8'b00001111; //  764 :  15 - 0xf
      11'h2FD: dout  = 8'b00000000; //  765 :   0 - 0x0
      11'h2FE: dout  = 8'b00000000; //  766 :   0 - 0x0
      11'h2FF: dout  = 8'b00000000; //  767 :   0 - 0x0
      11'h300: dout  = 8'b00000000; //  768 :   0 - 0x0 -- Sprite 0x60
      11'h301: dout  = 8'b00011000; //  769 :  24 - 0x18
      11'h302: dout  = 8'b00111100; //  770 :  60 - 0x3c
      11'h303: dout  = 8'b01111110; //  771 : 126 - 0x7e
      11'h304: dout  = 8'b01110110; //  772 : 118 - 0x76
      11'h305: dout  = 8'b11111011; //  773 : 251 - 0xfb
      11'h306: dout  = 8'b11111011; //  774 : 251 - 0xfb
      11'h307: dout  = 8'b11111011; //  775 : 251 - 0xfb
      11'h308: dout  = 8'b00000000; //  776 :   0 - 0x0 -- Sprite 0x61
      11'h309: dout  = 8'b00010000; //  777 :  16 - 0x10
      11'h30A: dout  = 8'b00010000; //  778 :  16 - 0x10
      11'h30B: dout  = 8'b00100000; //  779 :  32 - 0x20
      11'h30C: dout  = 8'b00100000; //  780 :  32 - 0x20
      11'h30D: dout  = 8'b00100000; //  781 :  32 - 0x20
      11'h30E: dout  = 8'b00100000; //  782 :  32 - 0x20
      11'h30F: dout  = 8'b00100000; //  783 :  32 - 0x20
      11'h310: dout  = 8'b00000000; //  784 :   0 - 0x0 -- Sprite 0x62
      11'h311: dout  = 8'b00001000; //  785 :   8 - 0x8
      11'h312: dout  = 8'b00001000; //  786 :   8 - 0x8
      11'h313: dout  = 8'b00001000; //  787 :   8 - 0x8
      11'h314: dout  = 8'b00001000; //  788 :   8 - 0x8
      11'h315: dout  = 8'b00001000; //  789 :   8 - 0x8
      11'h316: dout  = 8'b00001000; //  790 :   8 - 0x8
      11'h317: dout  = 8'b00001000; //  791 :   8 - 0x8
      11'h318: dout  = 8'b00000000; //  792 :   0 - 0x0 -- Sprite 0x63
      11'h319: dout  = 8'b00010000; //  793 :  16 - 0x10
      11'h31A: dout  = 8'b00010000; //  794 :  16 - 0x10
      11'h31B: dout  = 8'b00111000; //  795 :  56 - 0x38
      11'h31C: dout  = 8'b00111000; //  796 :  56 - 0x38
      11'h31D: dout  = 8'b00111000; //  797 :  56 - 0x38
      11'h31E: dout  = 8'b00111000; //  798 :  56 - 0x38
      11'h31F: dout  = 8'b00111000; //  799 :  56 - 0x38
      11'h320: dout  = 8'b00000000; //  800 :   0 - 0x0 -- Sprite 0x64
      11'h321: dout  = 8'b00011000; //  801 :  24 - 0x18
      11'h322: dout  = 8'b00111100; //  802 :  60 - 0x3c
      11'h323: dout  = 8'b00001110; //  803 :  14 - 0xe
      11'h324: dout  = 8'b00001110; //  804 :  14 - 0xe
      11'h325: dout  = 8'b00000100; //  805 :   4 - 0x4
      11'h326: dout  = 8'b00000000; //  806 :   0 - 0x0
      11'h327: dout  = 8'b00000000; //  807 :   0 - 0x0
      11'h328: dout  = 8'b00000000; //  808 :   0 - 0x0 -- Sprite 0x65
      11'h329: dout  = 8'b00000000; //  809 :   0 - 0x0
      11'h32A: dout  = 8'b00000100; //  810 :   4 - 0x4
      11'h32B: dout  = 8'b00000110; //  811 :   6 - 0x6
      11'h32C: dout  = 8'b00011110; //  812 :  30 - 0x1e
      11'h32D: dout  = 8'b00111100; //  813 :  60 - 0x3c
      11'h32E: dout  = 8'b00011000; //  814 :  24 - 0x18
      11'h32F: dout  = 8'b00000000; //  815 :   0 - 0x0
      11'h330: dout  = 8'b00000000; //  816 :   0 - 0x0 -- Sprite 0x66
      11'h331: dout  = 8'b00000000; //  817 :   0 - 0x0
      11'h332: dout  = 8'b00000001; //  818 :   1 - 0x1
      11'h333: dout  = 8'b00001010; //  819 :  10 - 0xa
      11'h334: dout  = 8'b00010111; //  820 :  23 - 0x17
      11'h335: dout  = 8'b00001111; //  821 :  15 - 0xf
      11'h336: dout  = 8'b00101111; //  822 :  47 - 0x2f
      11'h337: dout  = 8'b00011111; //  823 :  31 - 0x1f
      11'h338: dout  = 8'b00000000; //  824 :   0 - 0x0 -- Sprite 0x67
      11'h339: dout  = 8'b00000000; //  825 :   0 - 0x0
      11'h33A: dout  = 8'b00000000; //  826 :   0 - 0x0
      11'h33B: dout  = 8'b00000000; //  827 :   0 - 0x0
      11'h33C: dout  = 8'b00000101; //  828 :   5 - 0x5
      11'h33D: dout  = 8'b00000111; //  829 :   7 - 0x7
      11'h33E: dout  = 8'b00001111; //  830 :  15 - 0xf
      11'h33F: dout  = 8'b00000111; //  831 :   7 - 0x7
      11'h340: dout  = 8'b00000000; //  832 :   0 - 0x0 -- Sprite 0x68
      11'h341: dout  = 8'b00000000; //  833 :   0 - 0x0
      11'h342: dout  = 8'b00000000; //  834 :   0 - 0x0
      11'h343: dout  = 8'b00000000; //  835 :   0 - 0x0
      11'h344: dout  = 8'b00000000; //  836 :   0 - 0x0
      11'h345: dout  = 8'b00000000; //  837 :   0 - 0x0
      11'h346: dout  = 8'b00000001; //  838 :   1 - 0x1
      11'h347: dout  = 8'b00000011; //  839 :   3 - 0x3
      11'h348: dout  = 8'b00000000; //  840 :   0 - 0x0 -- Sprite 0x69
      11'h349: dout  = 8'b01100000; //  841 :  96 - 0x60
      11'h34A: dout  = 8'b11110000; //  842 : 240 - 0xf0
      11'h34B: dout  = 8'b11111000; //  843 : 248 - 0xf8
      11'h34C: dout  = 8'b01111100; //  844 : 124 - 0x7c
      11'h34D: dout  = 8'b00111110; //  845 :  62 - 0x3e
      11'h34E: dout  = 8'b01111110; //  846 : 126 - 0x7e
      11'h34F: dout  = 8'b01111111; //  847 : 127 - 0x7f
      11'h350: dout  = 8'b00111111; //  848 :  63 - 0x3f -- Sprite 0x6a
      11'h351: dout  = 8'b01011111; //  849 :  95 - 0x5f
      11'h352: dout  = 8'b01111111; //  850 : 127 - 0x7f
      11'h353: dout  = 8'b00111110; //  851 :  62 - 0x3e
      11'h354: dout  = 8'b00001110; //  852 :  14 - 0xe
      11'h355: dout  = 8'b00001010; //  853 :  10 - 0xa
      11'h356: dout  = 8'b01010001; //  854 :  81 - 0x51
      11'h357: dout  = 8'b00100000; //  855 :  32 - 0x20
      11'h358: dout  = 8'b00000000; //  856 :   0 - 0x0 -- Sprite 0x6b
      11'h359: dout  = 8'b00000000; //  857 :   0 - 0x0
      11'h35A: dout  = 8'b00000000; //  858 :   0 - 0x0
      11'h35B: dout  = 8'b00000000; //  859 :   0 - 0x0
      11'h35C: dout  = 8'b00000000; //  860 :   0 - 0x0
      11'h35D: dout  = 8'b00000000; //  861 :   0 - 0x0
      11'h35E: dout  = 8'b00001110; //  862 :  14 - 0xe
      11'h35F: dout  = 8'b00011111; //  863 :  31 - 0x1f
      11'h360: dout  = 8'b00111111; //  864 :  63 - 0x3f -- Sprite 0x6c
      11'h361: dout  = 8'b01111111; //  865 : 127 - 0x7f
      11'h362: dout  = 8'b01111111; //  866 : 127 - 0x7f
      11'h363: dout  = 8'b11111110; //  867 : 254 - 0xfe
      11'h364: dout  = 8'b11101100; //  868 : 236 - 0xec
      11'h365: dout  = 8'b11001010; //  869 : 202 - 0xca
      11'h366: dout  = 8'b01010001; //  870 :  81 - 0x51
      11'h367: dout  = 8'b00100000; //  871 :  32 - 0x20
      11'h368: dout  = 8'b00000000; //  872 :   0 - 0x0 -- Sprite 0x6d
      11'h369: dout  = 8'b01000000; //  873 :  64 - 0x40
      11'h36A: dout  = 8'b01100011; //  874 :  99 - 0x63
      11'h36B: dout  = 8'b01110111; //  875 : 119 - 0x77
      11'h36C: dout  = 8'b01111100; //  876 : 124 - 0x7c
      11'h36D: dout  = 8'b00111000; //  877 :  56 - 0x38
      11'h36E: dout  = 8'b11111000; //  878 : 248 - 0xf8
      11'h36F: dout  = 8'b11100100; //  879 : 228 - 0xe4
      11'h370: dout  = 8'b00000000; //  880 :   0 - 0x0 -- Sprite 0x6e
      11'h371: dout  = 8'b00000000; //  881 :   0 - 0x0
      11'h372: dout  = 8'b00000011; //  882 :   3 - 0x3
      11'h373: dout  = 8'b00000111; //  883 :   7 - 0x7
      11'h374: dout  = 8'b00001100; //  884 :  12 - 0xc
      11'h375: dout  = 8'b00011000; //  885 :  24 - 0x18
      11'h376: dout  = 8'b11111000; //  886 : 248 - 0xf8
      11'h377: dout  = 8'b11100100; //  887 : 228 - 0xe4
      11'h378: dout  = 8'b00000011; //  888 :   3 - 0x3 -- Sprite 0x6f
      11'h379: dout  = 8'b01000100; //  889 :  68 - 0x44
      11'h37A: dout  = 8'b00101000; //  890 :  40 - 0x28
      11'h37B: dout  = 8'b00010000; //  891 :  16 - 0x10
      11'h37C: dout  = 8'b00001000; //  892 :   8 - 0x8
      11'h37D: dout  = 8'b00000100; //  893 :   4 - 0x4
      11'h37E: dout  = 8'b00000011; //  894 :   3 - 0x3
      11'h37F: dout  = 8'b00000100; //  895 :   4 - 0x4
      11'h380: dout  = 8'b00000011; //  896 :   3 - 0x3 -- Sprite 0x70
      11'h381: dout  = 8'b00000111; //  897 :   7 - 0x7
      11'h382: dout  = 8'b00001111; //  898 :  15 - 0xf
      11'h383: dout  = 8'b00011111; //  899 :  31 - 0x1f
      11'h384: dout  = 8'b00100111; //  900 :  39 - 0x27
      11'h385: dout  = 8'b01111011; //  901 : 123 - 0x7b
      11'h386: dout  = 8'b01111000; //  902 : 120 - 0x78
      11'h387: dout  = 8'b11111011; //  903 : 251 - 0xfb
      11'h388: dout  = 8'b11000000; //  904 : 192 - 0xc0 -- Sprite 0x71
      11'h389: dout  = 8'b11100000; //  905 : 224 - 0xe0
      11'h38A: dout  = 8'b11110000; //  906 : 240 - 0xf0
      11'h38B: dout  = 8'b11111000; //  907 : 248 - 0xf8
      11'h38C: dout  = 8'b11100100; //  908 : 228 - 0xe4
      11'h38D: dout  = 8'b11011110; //  909 : 222 - 0xde
      11'h38E: dout  = 8'b00011110; //  910 :  30 - 0x1e
      11'h38F: dout  = 8'b11011111; //  911 : 223 - 0xdf
      11'h390: dout  = 8'b11111111; //  912 : 255 - 0xff -- Sprite 0x72
      11'h391: dout  = 8'b11111111; //  913 : 255 - 0xff
      11'h392: dout  = 8'b01111111; //  914 : 127 - 0x7f
      11'h393: dout  = 8'b00001111; //  915 :  15 - 0xf
      11'h394: dout  = 8'b00001111; //  916 :  15 - 0xf
      11'h395: dout  = 8'b00000111; //  917 :   7 - 0x7
      11'h396: dout  = 8'b00000011; //  918 :   3 - 0x3
      11'h397: dout  = 8'b00000000; //  919 :   0 - 0x0
      11'h398: dout  = 8'b11111111; //  920 : 255 - 0xff -- Sprite 0x73
      11'h399: dout  = 8'b11111111; //  921 : 255 - 0xff
      11'h39A: dout  = 8'b11111110; //  922 : 254 - 0xfe
      11'h39B: dout  = 8'b11110000; //  923 : 240 - 0xf0
      11'h39C: dout  = 8'b11110000; //  924 : 240 - 0xf0
      11'h39D: dout  = 8'b11000000; //  925 : 192 - 0xc0
      11'h39E: dout  = 8'b10000000; //  926 : 128 - 0x80
      11'h39F: dout  = 8'b00000000; //  927 :   0 - 0x0
      11'h3A0: dout  = 8'b00000000; //  928 :   0 - 0x0 -- Sprite 0x74
      11'h3A1: dout  = 8'b00000000; //  929 :   0 - 0x0
      11'h3A2: dout  = 8'b00011000; //  930 :  24 - 0x18
      11'h3A3: dout  = 8'b00100100; //  931 :  36 - 0x24
      11'h3A4: dout  = 8'b00100100; //  932 :  36 - 0x24
      11'h3A5: dout  = 8'b00011000; //  933 :  24 - 0x18
      11'h3A6: dout  = 8'b00000000; //  934 :   0 - 0x0
      11'h3A7: dout  = 8'b00000000; //  935 :   0 - 0x0
      11'h3A8: dout  = 8'b00111100; //  936 :  60 - 0x3c -- Sprite 0x75
      11'h3A9: dout  = 8'b01111110; //  937 : 126 - 0x7e
      11'h3AA: dout  = 8'b11111111; //  938 : 255 - 0xff
      11'h3AB: dout  = 8'b11111111; //  939 : 255 - 0xff
      11'h3AC: dout  = 8'b11111111; //  940 : 255 - 0xff
      11'h3AD: dout  = 8'b11111111; //  941 : 255 - 0xff
      11'h3AE: dout  = 8'b01111110; //  942 : 126 - 0x7e
      11'h3AF: dout  = 8'b00111100; //  943 :  60 - 0x3c
      11'h3B0: dout  = 8'b00000011; //  944 :   3 - 0x3 -- Sprite 0x76
      11'h3B1: dout  = 8'b00000111; //  945 :   7 - 0x7
      11'h3B2: dout  = 8'b00001111; //  946 :  15 - 0xf
      11'h3B3: dout  = 8'b00011111; //  947 :  31 - 0x1f
      11'h3B4: dout  = 8'b00111111; //  948 :  63 - 0x3f
      11'h3B5: dout  = 8'b01100011; //  949 :  99 - 0x63
      11'h3B6: dout  = 8'b01000001; //  950 :  65 - 0x41
      11'h3B7: dout  = 8'b11000001; //  951 : 193 - 0xc1
      11'h3B8: dout  = 8'b11000000; //  952 : 192 - 0xc0 -- Sprite 0x77
      11'h3B9: dout  = 8'b10000000; //  953 : 128 - 0x80
      11'h3BA: dout  = 8'b00000000; //  954 :   0 - 0x0
      11'h3BB: dout  = 8'b00000000; //  955 :   0 - 0x0
      11'h3BC: dout  = 8'b10001100; //  956 : 140 - 0x8c
      11'h3BD: dout  = 8'b11111110; //  957 : 254 - 0xfe
      11'h3BE: dout  = 8'b11111110; //  958 : 254 - 0xfe
      11'h3BF: dout  = 8'b11110011; //  959 : 243 - 0xf3
      11'h3C0: dout  = 8'b11000001; //  960 : 193 - 0xc1 -- Sprite 0x78
      11'h3C1: dout  = 8'b11100011; //  961 : 227 - 0xe3
      11'h3C2: dout  = 8'b11111111; //  962 : 255 - 0xff
      11'h3C3: dout  = 8'b01000111; //  963 :  71 - 0x47
      11'h3C4: dout  = 8'b00001111; //  964 :  15 - 0xf
      11'h3C5: dout  = 8'b00001111; //  965 :  15 - 0xf
      11'h3C6: dout  = 8'b00001111; //  966 :  15 - 0xf
      11'h3C7: dout  = 8'b00000111; //  967 :   7 - 0x7
      11'h3C8: dout  = 8'b11110001; //  968 : 241 - 0xf1 -- Sprite 0x79
      11'h3C9: dout  = 8'b11111001; //  969 : 249 - 0xf9
      11'h3CA: dout  = 8'b11111111; //  970 : 255 - 0xff
      11'h3CB: dout  = 8'b11100010; //  971 : 226 - 0xe2
      11'h3CC: dout  = 8'b11110000; //  972 : 240 - 0xf0
      11'h3CD: dout  = 8'b11110000; //  973 : 240 - 0xf0
      11'h3CE: dout  = 8'b11110000; //  974 : 240 - 0xf0
      11'h3CF: dout  = 8'b11100000; //  975 : 224 - 0xe0
      11'h3D0: dout  = 8'b00010110; //  976 :  22 - 0x16 -- Sprite 0x7a
      11'h3D1: dout  = 8'b00011111; //  977 :  31 - 0x1f
      11'h3D2: dout  = 8'b00000000; //  978 :   0 - 0x0
      11'h3D3: dout  = 8'b00000000; //  979 :   0 - 0x0
      11'h3D4: dout  = 8'b00000101; //  980 :   5 - 0x5
      11'h3D5: dout  = 8'b00001101; //  981 :  13 - 0xd
      11'h3D6: dout  = 8'b00111111; //  982 :  63 - 0x3f
      11'h3D7: dout  = 8'b00011111; //  983 :  31 - 0x1f
      11'h3D8: dout  = 8'b10000000; //  984 : 128 - 0x80 -- Sprite 0x7b
      11'h3D9: dout  = 8'b10000000; //  985 : 128 - 0x80
      11'h3DA: dout  = 8'b00000000; //  986 :   0 - 0x0
      11'h3DB: dout  = 8'b00000000; //  987 :   0 - 0x0
      11'h3DC: dout  = 8'b00000000; //  988 :   0 - 0x0
      11'h3DD: dout  = 8'b10100000; //  989 : 160 - 0xa0
      11'h3DE: dout  = 8'b10100000; //  990 : 160 - 0xa0
      11'h3DF: dout  = 8'b11100000; //  991 : 224 - 0xe0
      11'h3E0: dout  = 8'b00000000; //  992 :   0 - 0x0 -- Sprite 0x7c
      11'h3E1: dout  = 8'b00000100; //  993 :   4 - 0x4
      11'h3E2: dout  = 8'b01001110; //  994 :  78 - 0x4e
      11'h3E3: dout  = 8'b10001100; //  995 : 140 - 0x8c
      11'h3E4: dout  = 8'b00001100; //  996 :  12 - 0xc
      11'h3E5: dout  = 8'b01111111; //  997 : 127 - 0x7f
      11'h3E6: dout  = 8'b11111111; //  998 : 255 - 0xff
      11'h3E7: dout  = 8'b11111111; //  999 : 255 - 0xff
      11'h3E8: dout  = 8'b00000000; // 1000 :   0 - 0x0 -- Sprite 0x7d
      11'h3E9: dout  = 8'b00000000; // 1001 :   0 - 0x0
      11'h3EA: dout  = 8'b00000000; // 1002 :   0 - 0x0
      11'h3EB: dout  = 8'b00000000; // 1003 :   0 - 0x0
      11'h3EC: dout  = 8'b00000000; // 1004 :   0 - 0x0
      11'h3ED: dout  = 8'b00000000; // 1005 :   0 - 0x0
      11'h3EE: dout  = 8'b00000001; // 1006 :   1 - 0x1
      11'h3EF: dout  = 8'b00000001; // 1007 :   1 - 0x1
      11'h3F0: dout  = 8'b11111111; // 1008 : 255 - 0xff -- Sprite 0x7e
      11'h3F1: dout  = 8'b01111111; // 1009 : 127 - 0x7f
      11'h3F2: dout  = 8'b00111111; // 1010 :  63 - 0x3f
      11'h3F3: dout  = 8'b00011111; // 1011 :  31 - 0x1f
      11'h3F4: dout  = 8'b00001111; // 1012 :  15 - 0xf
      11'h3F5: dout  = 8'b00000111; // 1013 :   7 - 0x7
      11'h3F6: dout  = 8'b00000011; // 1014 :   3 - 0x3
      11'h3F7: dout  = 8'b00000001; // 1015 :   1 - 0x1
      11'h3F8: dout  = 8'b11111111; // 1016 : 255 - 0xff -- Sprite 0x7f
      11'h3F9: dout  = 8'b10000011; // 1017 : 131 - 0x83
      11'h3FA: dout  = 8'b00101001; // 1018 :  41 - 0x29
      11'h3FB: dout  = 8'b01101101; // 1019 : 109 - 0x6d
      11'h3FC: dout  = 8'b01000101; // 1020 :  69 - 0x45
      11'h3FD: dout  = 8'b00010001; // 1021 :  17 - 0x11
      11'h3FE: dout  = 8'b00000001; // 1022 :   1 - 0x1
      11'h3FF: dout  = 8'b11000111; // 1023 : 199 - 0xc7
      11'h400: dout  = 8'b00001000; // 1024 :   8 - 0x8 -- Sprite 0x80
      11'h401: dout  = 8'b00001000; // 1025 :   8 - 0x8
      11'h402: dout  = 8'b00000010; // 1026 :   2 - 0x2
      11'h403: dout  = 8'b00011111; // 1027 :  31 - 0x1f
      11'h404: dout  = 8'b00100010; // 1028 :  34 - 0x22
      11'h405: dout  = 8'b00000010; // 1029 :   2 - 0x2
      11'h406: dout  = 8'b00000010; // 1030 :   2 - 0x2
      11'h407: dout  = 8'b00000000; // 1031 :   0 - 0x0
      11'h408: dout  = 8'b00001000; // 1032 :   8 - 0x8 -- Sprite 0x81
      11'h409: dout  = 8'b00001000; // 1033 :   8 - 0x8
      11'h40A: dout  = 8'b00001000; // 1034 :   8 - 0x8
      11'h40B: dout  = 8'b00001000; // 1035 :   8 - 0x8
      11'h40C: dout  = 8'b00001000; // 1036 :   8 - 0x8
      11'h40D: dout  = 8'b00001000; // 1037 :   8 - 0x8
      11'h40E: dout  = 8'b00001000; // 1038 :   8 - 0x8
      11'h40F: dout  = 8'b00001000; // 1039 :   8 - 0x8
      11'h410: dout  = 8'b00010000; // 1040 :  16 - 0x10 -- Sprite 0x82
      11'h411: dout  = 8'b00011110; // 1041 :  30 - 0x1e
      11'h412: dout  = 8'b00010000; // 1042 :  16 - 0x10
      11'h413: dout  = 8'b01010000; // 1043 :  80 - 0x50
      11'h414: dout  = 8'b00010000; // 1044 :  16 - 0x10
      11'h415: dout  = 8'b00001000; // 1045 :   8 - 0x8
      11'h416: dout  = 8'b00000000; // 1046 :   0 - 0x0
      11'h417: dout  = 8'b00000000; // 1047 :   0 - 0x0
      11'h418: dout  = 8'b00000000; // 1048 :   0 - 0x0 -- Sprite 0x83
      11'h419: dout  = 8'b00000000; // 1049 :   0 - 0x0
      11'h41A: dout  = 8'b00000000; // 1050 :   0 - 0x0
      11'h41B: dout  = 8'b11111110; // 1051 : 254 - 0xfe
      11'h41C: dout  = 8'b00000000; // 1052 :   0 - 0x0
      11'h41D: dout  = 8'b00000000; // 1053 :   0 - 0x0
      11'h41E: dout  = 8'b00000000; // 1054 :   0 - 0x0
      11'h41F: dout  = 8'b00000000; // 1055 :   0 - 0x0
      11'h420: dout  = 8'b00011100; // 1056 :  28 - 0x1c -- Sprite 0x84
      11'h421: dout  = 8'b00101010; // 1057 :  42 - 0x2a
      11'h422: dout  = 8'b01110111; // 1058 : 119 - 0x77
      11'h423: dout  = 8'b11101110; // 1059 : 238 - 0xee
      11'h424: dout  = 8'b11011101; // 1060 : 221 - 0xdd
      11'h425: dout  = 8'b10101010; // 1061 : 170 - 0xaa
      11'h426: dout  = 8'b01110100; // 1062 : 116 - 0x74
      11'h427: dout  = 8'b00101000; // 1063 :  40 - 0x28
      11'h428: dout  = 8'b11111111; // 1064 : 255 - 0xff -- Sprite 0x85
      11'h429: dout  = 8'b11111110; // 1065 : 254 - 0xfe
      11'h42A: dout  = 8'b11111110; // 1066 : 254 - 0xfe
      11'h42B: dout  = 8'b00000000; // 1067 :   0 - 0x0
      11'h42C: dout  = 8'b11101111; // 1068 : 239 - 0xef
      11'h42D: dout  = 8'b11101111; // 1069 : 239 - 0xef
      11'h42E: dout  = 8'b11101111; // 1070 : 239 - 0xef
      11'h42F: dout  = 8'b00000000; // 1071 :   0 - 0x0
      11'h430: dout  = 8'b11111110; // 1072 : 254 - 0xfe -- Sprite 0x86
      11'h431: dout  = 8'b11111110; // 1073 : 254 - 0xfe
      11'h432: dout  = 8'b11111110; // 1074 : 254 - 0xfe
      11'h433: dout  = 8'b00000000; // 1075 :   0 - 0x0
      11'h434: dout  = 8'b11101111; // 1076 : 239 - 0xef
      11'h435: dout  = 8'b11101111; // 1077 : 239 - 0xef
      11'h436: dout  = 8'b11101111; // 1078 : 239 - 0xef
      11'h437: dout  = 8'b00000000; // 1079 :   0 - 0x0
      11'h438: dout  = 8'b00000000; // 1080 :   0 - 0x0 -- Sprite 0x87
      11'h439: dout  = 8'b01111111; // 1081 : 127 - 0x7f
      11'h43A: dout  = 8'b01011111; // 1082 :  95 - 0x5f
      11'h43B: dout  = 8'b01111111; // 1083 : 127 - 0x7f
      11'h43C: dout  = 8'b01111111; // 1084 : 127 - 0x7f
      11'h43D: dout  = 8'b01111111; // 1085 : 127 - 0x7f
      11'h43E: dout  = 8'b01111111; // 1086 : 127 - 0x7f
      11'h43F: dout  = 8'b01111111; // 1087 : 127 - 0x7f
      11'h440: dout  = 8'b10111000; // 1088 : 184 - 0xb8 -- Sprite 0x88
      11'h441: dout  = 8'b10011110; // 1089 : 158 - 0x9e
      11'h442: dout  = 8'b10000000; // 1090 : 128 - 0x80
      11'h443: dout  = 8'b11000000; // 1091 : 192 - 0xc0
      11'h444: dout  = 8'b11100000; // 1092 : 224 - 0xe0
      11'h445: dout  = 8'b11110000; // 1093 : 240 - 0xf0
      11'h446: dout  = 8'b11111000; // 1094 : 248 - 0xf8
      11'h447: dout  = 8'b01111100; // 1095 : 124 - 0x7c
      11'h448: dout  = 8'b00000000; // 1096 :   0 - 0x0 -- Sprite 0x89
      11'h449: dout  = 8'b00100011; // 1097 :  35 - 0x23
      11'h44A: dout  = 8'b01010111; // 1098 :  87 - 0x57
      11'h44B: dout  = 8'b01001111; // 1099 :  79 - 0x4f
      11'h44C: dout  = 8'b01010111; // 1100 :  87 - 0x57
      11'h44D: dout  = 8'b00100111; // 1101 :  39 - 0x27
      11'h44E: dout  = 8'b11000011; // 1102 : 195 - 0xc3
      11'h44F: dout  = 8'b00100001; // 1103 :  33 - 0x21
      11'h450: dout  = 8'b00000000; // 1104 :   0 - 0x0 -- Sprite 0x8a
      11'h451: dout  = 8'b00110000; // 1105 :  48 - 0x30
      11'h452: dout  = 8'b01110000; // 1106 : 112 - 0x70
      11'h453: dout  = 8'b01110000; // 1107 : 112 - 0x70
      11'h454: dout  = 8'b11110000; // 1108 : 240 - 0xf0
      11'h455: dout  = 8'b11100000; // 1109 : 224 - 0xe0
      11'h456: dout  = 8'b11000000; // 1110 : 192 - 0xc0
      11'h457: dout  = 8'b00000000; // 1111 :   0 - 0x0
      11'h458: dout  = 8'b00010011; // 1112 :  19 - 0x13 -- Sprite 0x8b
      11'h459: dout  = 8'b00001111; // 1113 :  15 - 0xf
      11'h45A: dout  = 8'b00011110; // 1114 :  30 - 0x1e
      11'h45B: dout  = 8'b11110000; // 1115 : 240 - 0xf0
      11'h45C: dout  = 8'b11111100; // 1116 : 252 - 0xfc
      11'h45D: dout  = 8'b11111000; // 1117 : 248 - 0xf8
      11'h45E: dout  = 8'b11110000; // 1118 : 240 - 0xf0
      11'h45F: dout  = 8'b11100000; // 1119 : 224 - 0xe0
      11'h460: dout  = 8'b10111110; // 1120 : 190 - 0xbe -- Sprite 0x8c
      11'h461: dout  = 8'b10010000; // 1121 : 144 - 0x90
      11'h462: dout  = 8'b10000000; // 1122 : 128 - 0x80
      11'h463: dout  = 8'b11000000; // 1123 : 192 - 0xc0
      11'h464: dout  = 8'b11000000; // 1124 : 192 - 0xc0
      11'h465: dout  = 8'b10000000; // 1125 : 128 - 0x80
      11'h466: dout  = 8'b00000000; // 1126 :   0 - 0x0
      11'h467: dout  = 8'b00000000; // 1127 :   0 - 0x0
      11'h468: dout  = 8'b00000001; // 1128 :   1 - 0x1 -- Sprite 0x8d
      11'h469: dout  = 8'b00000001; // 1129 :   1 - 0x1
      11'h46A: dout  = 8'b00000011; // 1130 :   3 - 0x3
      11'h46B: dout  = 8'b00000011; // 1131 :   3 - 0x3
      11'h46C: dout  = 8'b00000111; // 1132 :   7 - 0x7
      11'h46D: dout  = 8'b01111111; // 1133 : 127 - 0x7f
      11'h46E: dout  = 8'b01111101; // 1134 : 125 - 0x7d
      11'h46F: dout  = 8'b00111101; // 1135 :  61 - 0x3d
      11'h470: dout  = 8'b00000110; // 1136 :   6 - 0x6 -- Sprite 0x8e
      11'h471: dout  = 8'b00000100; // 1137 :   4 - 0x4
      11'h472: dout  = 8'b00110000; // 1138 :  48 - 0x30
      11'h473: dout  = 8'b00100011; // 1139 :  35 - 0x23
      11'h474: dout  = 8'b00000110; // 1140 :   6 - 0x6
      11'h475: dout  = 8'b01100100; // 1141 : 100 - 0x64
      11'h476: dout  = 8'b01100000; // 1142 :  96 - 0x60
      11'h477: dout  = 8'b00000000; // 1143 :   0 - 0x0
      11'h478: dout  = 8'b00000000; // 1144 :   0 - 0x0 -- Sprite 0x8f
      11'h479: dout  = 8'b01100000; // 1145 :  96 - 0x60
      11'h47A: dout  = 8'b01100000; // 1146 :  96 - 0x60
      11'h47B: dout  = 8'b00000000; // 1147 :   0 - 0x0
      11'h47C: dout  = 8'b00100000; // 1148 :  32 - 0x20
      11'h47D: dout  = 8'b00110000; // 1149 :  48 - 0x30
      11'h47E: dout  = 8'b00000100; // 1150 :   4 - 0x4
      11'h47F: dout  = 8'b00000110; // 1151 :   6 - 0x6
      11'h480: dout  = 8'b00000000; // 1152 :   0 - 0x0 -- Sprite 0x90
      11'h481: dout  = 8'b00000001; // 1153 :   1 - 0x1
      11'h482: dout  = 8'b00000001; // 1154 :   1 - 0x1
      11'h483: dout  = 8'b00000000; // 1155 :   0 - 0x0
      11'h484: dout  = 8'b00000000; // 1156 :   0 - 0x0
      11'h485: dout  = 8'b00000000; // 1157 :   0 - 0x0
      11'h486: dout  = 8'b00000000; // 1158 :   0 - 0x0
      11'h487: dout  = 8'b00000000; // 1159 :   0 - 0x0
      11'h488: dout  = 8'b11111110; // 1160 : 254 - 0xfe -- Sprite 0x91
      11'h489: dout  = 8'b11111111; // 1161 : 255 - 0xff
      11'h48A: dout  = 8'b11111111; // 1162 : 255 - 0xff
      11'h48B: dout  = 8'b01000000; // 1163 :  64 - 0x40
      11'h48C: dout  = 8'b00000001; // 1164 :   1 - 0x1
      11'h48D: dout  = 8'b00000011; // 1165 :   3 - 0x3
      11'h48E: dout  = 8'b00000011; // 1166 :   3 - 0x3
      11'h48F: dout  = 8'b00000011; // 1167 :   3 - 0x3
      11'h490: dout  = 8'b00000001; // 1168 :   1 - 0x1 -- Sprite 0x92
      11'h491: dout  = 8'b00000001; // 1169 :   1 - 0x1
      11'h492: dout  = 8'b00000000; // 1170 :   0 - 0x0
      11'h493: dout  = 8'b00000000; // 1171 :   0 - 0x0
      11'h494: dout  = 8'b00000000; // 1172 :   0 - 0x0
      11'h495: dout  = 8'b00000000; // 1173 :   0 - 0x0
      11'h496: dout  = 8'b00000000; // 1174 :   0 - 0x0
      11'h497: dout  = 8'b00000000; // 1175 :   0 - 0x0
      11'h498: dout  = 8'b11100000; // 1176 : 224 - 0xe0 -- Sprite 0x93
      11'h499: dout  = 8'b11111110; // 1177 : 254 - 0xfe
      11'h49A: dout  = 8'b11111111; // 1178 : 255 - 0xff
      11'h49B: dout  = 8'b01111111; // 1179 : 127 - 0x7f
      11'h49C: dout  = 8'b00000011; // 1180 :   3 - 0x3
      11'h49D: dout  = 8'b00000010; // 1181 :   2 - 0x2
      11'h49E: dout  = 8'b00000000; // 1182 :   0 - 0x0
      11'h49F: dout  = 8'b00000000; // 1183 :   0 - 0x0
      11'h4A0: dout  = 8'b00000001; // 1184 :   1 - 0x1 -- Sprite 0x94
      11'h4A1: dout  = 8'b00001101; // 1185 :  13 - 0xd
      11'h4A2: dout  = 8'b00001000; // 1186 :   8 - 0x8
      11'h4A3: dout  = 8'b00000000; // 1187 :   0 - 0x0
      11'h4A4: dout  = 8'b00110110; // 1188 :  54 - 0x36
      11'h4A5: dout  = 8'b00101100; // 1189 :  44 - 0x2c
      11'h4A6: dout  = 8'b00001000; // 1190 :   8 - 0x8
      11'h4A7: dout  = 8'b01100000; // 1191 :  96 - 0x60
      11'h4A8: dout  = 8'b01100000; // 1192 :  96 - 0x60 -- Sprite 0x95
      11'h4A9: dout  = 8'b00000000; // 1193 :   0 - 0x0
      11'h4AA: dout  = 8'b00100000; // 1194 :  32 - 0x20
      11'h4AB: dout  = 8'b00110000; // 1195 :  48 - 0x30
      11'h4AC: dout  = 8'b00000000; // 1196 :   0 - 0x0
      11'h4AD: dout  = 8'b00001000; // 1197 :   8 - 0x8
      11'h4AE: dout  = 8'b00001101; // 1198 :  13 - 0xd
      11'h4AF: dout  = 8'b00000001; // 1199 :   1 - 0x1
      11'h4B0: dout  = 8'b00000001; // 1200 :   1 - 0x1 -- Sprite 0x96
      11'h4B1: dout  = 8'b00000001; // 1201 :   1 - 0x1
      11'h4B2: dout  = 8'b00000011; // 1202 :   3 - 0x3
      11'h4B3: dout  = 8'b01000011; // 1203 :  67 - 0x43
      11'h4B4: dout  = 8'b01100111; // 1204 : 103 - 0x67
      11'h4B5: dout  = 8'b01110111; // 1205 : 119 - 0x77
      11'h4B6: dout  = 8'b01111011; // 1206 : 123 - 0x7b
      11'h4B7: dout  = 8'b01111000; // 1207 : 120 - 0x78
      11'h4B8: dout  = 8'b00000000; // 1208 :   0 - 0x0 -- Sprite 0x97
      11'h4B9: dout  = 8'b00000000; // 1209 :   0 - 0x0
      11'h4BA: dout  = 8'b10000000; // 1210 : 128 - 0x80
      11'h4BB: dout  = 8'b10000100; // 1211 : 132 - 0x84
      11'h4BC: dout  = 8'b11001100; // 1212 : 204 - 0xcc
      11'h4BD: dout  = 8'b11011100; // 1213 : 220 - 0xdc
      11'h4BE: dout  = 8'b10111100; // 1214 : 188 - 0xbc
      11'h4BF: dout  = 8'b00111100; // 1215 :  60 - 0x3c
      11'h4C0: dout  = 8'b00110011; // 1216 :  51 - 0x33 -- Sprite 0x98
      11'h4C1: dout  = 8'b00000111; // 1217 :   7 - 0x7
      11'h4C2: dout  = 8'b00000111; // 1218 :   7 - 0x7
      11'h4C3: dout  = 8'b11100011; // 1219 : 227 - 0xe3
      11'h4C4: dout  = 8'b00111000; // 1220 :  56 - 0x38
      11'h4C5: dout  = 8'b00111111; // 1221 :  63 - 0x3f
      11'h4C6: dout  = 8'b00011100; // 1222 :  28 - 0x1c
      11'h4C7: dout  = 8'b00001100; // 1223 :  12 - 0xc
      11'h4C8: dout  = 8'b10011000; // 1224 : 152 - 0x98 -- Sprite 0x99
      11'h4C9: dout  = 8'b11000111; // 1225 : 199 - 0xc7
      11'h4CA: dout  = 8'b11001000; // 1226 : 200 - 0xc8
      11'h4CB: dout  = 8'b10010010; // 1227 : 146 - 0x92
      11'h4CC: dout  = 8'b00110000; // 1228 :  48 - 0x30
      11'h4CD: dout  = 8'b11111000; // 1229 : 248 - 0xf8
      11'h4CE: dout  = 8'b01110000; // 1230 : 112 - 0x70
      11'h4CF: dout  = 8'b01100000; // 1231 :  96 - 0x60
      11'h4D0: dout  = 8'b00000000; // 1232 :   0 - 0x0 -- Sprite 0x9a
      11'h4D1: dout  = 8'b00000001; // 1233 :   1 - 0x1
      11'h4D2: dout  = 8'b00000001; // 1234 :   1 - 0x1
      11'h4D3: dout  = 8'b00000011; // 1235 :   3 - 0x3
      11'h4D4: dout  = 8'b01000011; // 1236 :  67 - 0x43
      11'h4D5: dout  = 8'b01100111; // 1237 : 103 - 0x67
      11'h4D6: dout  = 8'b01110111; // 1238 : 119 - 0x77
      11'h4D7: dout  = 8'b01111011; // 1239 : 123 - 0x7b
      11'h4D8: dout  = 8'b00000000; // 1240 :   0 - 0x0 -- Sprite 0x9b
      11'h4D9: dout  = 8'b00000000; // 1241 :   0 - 0x0
      11'h4DA: dout  = 8'b00000000; // 1242 :   0 - 0x0
      11'h4DB: dout  = 8'b10000000; // 1243 : 128 - 0x80
      11'h4DC: dout  = 8'b10000100; // 1244 : 132 - 0x84
      11'h4DD: dout  = 8'b11001100; // 1245 : 204 - 0xcc
      11'h4DE: dout  = 8'b11011100; // 1246 : 220 - 0xdc
      11'h4DF: dout  = 8'b10111100; // 1247 : 188 - 0xbc
      11'h4E0: dout  = 8'b01111000; // 1248 : 120 - 0x78 -- Sprite 0x9c
      11'h4E1: dout  = 8'b00110011; // 1249 :  51 - 0x33
      11'h4E2: dout  = 8'b00000111; // 1250 :   7 - 0x7
      11'h4E3: dout  = 8'b00000111; // 1251 :   7 - 0x7
      11'h4E4: dout  = 8'b11100011; // 1252 : 227 - 0xe3
      11'h4E5: dout  = 8'b00111000; // 1253 :  56 - 0x38
      11'h4E6: dout  = 8'b01111111; // 1254 : 127 - 0x7f
      11'h4E7: dout  = 8'b11110000; // 1255 : 240 - 0xf0
      11'h4E8: dout  = 8'b00111100; // 1256 :  60 - 0x3c -- Sprite 0x9d
      11'h4E9: dout  = 8'b10011000; // 1257 : 152 - 0x98
      11'h4EA: dout  = 8'b11000111; // 1258 : 199 - 0xc7
      11'h4EB: dout  = 8'b11001000; // 1259 : 200 - 0xc8
      11'h4EC: dout  = 8'b10010010; // 1260 : 146 - 0x92
      11'h4ED: dout  = 8'b00110000; // 1261 :  48 - 0x30
      11'h4EE: dout  = 8'b11111000; // 1262 : 248 - 0xf8
      11'h4EF: dout  = 8'b00111100; // 1263 :  60 - 0x3c
      11'h4F0: dout  = 8'b00000000; // 1264 :   0 - 0x0 -- Sprite 0x9e
      11'h4F1: dout  = 8'b00010000; // 1265 :  16 - 0x10
      11'h4F2: dout  = 8'b01111111; // 1266 : 127 - 0x7f
      11'h4F3: dout  = 8'b01111111; // 1267 : 127 - 0x7f
      11'h4F4: dout  = 8'b01111111; // 1268 : 127 - 0x7f
      11'h4F5: dout  = 8'b00011111; // 1269 :  31 - 0x1f
      11'h4F6: dout  = 8'b00001111; // 1270 :  15 - 0xf
      11'h4F7: dout  = 8'b00001111; // 1271 :  15 - 0xf
      11'h4F8: dout  = 8'b00000011; // 1272 :   3 - 0x3 -- Sprite 0x9f
      11'h4F9: dout  = 8'b00110011; // 1273 :  51 - 0x33
      11'h4FA: dout  = 8'b00111001; // 1274 :  57 - 0x39
      11'h4FB: dout  = 8'b00111010; // 1275 :  58 - 0x3a
      11'h4FC: dout  = 8'b00111000; // 1276 :  56 - 0x38
      11'h4FD: dout  = 8'b00011000; // 1277 :  24 - 0x18
      11'h4FE: dout  = 8'b00000000; // 1278 :   0 - 0x0
      11'h4FF: dout  = 8'b00000000; // 1279 :   0 - 0x0
      11'h500: dout  = 8'b00010000; // 1280 :  16 - 0x10 -- Sprite 0xa0
      11'h501: dout  = 8'b00111000; // 1281 :  56 - 0x38
      11'h502: dout  = 8'b00111100; // 1282 :  60 - 0x3c
      11'h503: dout  = 8'b01110100; // 1283 : 116 - 0x74
      11'h504: dout  = 8'b01110110; // 1284 : 118 - 0x76
      11'h505: dout  = 8'b01110110; // 1285 : 118 - 0x76
      11'h506: dout  = 8'b01111110; // 1286 : 126 - 0x7e
      11'h507: dout  = 8'b01111101; // 1287 : 125 - 0x7d
      11'h508: dout  = 8'b00000000; // 1288 :   0 - 0x0 -- Sprite 0xa1
      11'h509: dout  = 8'b00000000; // 1289 :   0 - 0x0
      11'h50A: dout  = 8'b00010001; // 1290 :  17 - 0x11
      11'h50B: dout  = 8'b00001010; // 1291 :  10 - 0xa
      11'h50C: dout  = 8'b00110100; // 1292 :  52 - 0x34
      11'h50D: dout  = 8'b00101010; // 1293 :  42 - 0x2a
      11'h50E: dout  = 8'b01010001; // 1294 :  81 - 0x51
      11'h50F: dout  = 8'b00100000; // 1295 :  32 - 0x20
      11'h510: dout  = 8'b01111111; // 1296 : 127 - 0x7f -- Sprite 0xa2
      11'h511: dout  = 8'b01100111; // 1297 : 103 - 0x67
      11'h512: dout  = 8'b01100011; // 1298 :  99 - 0x63
      11'h513: dout  = 8'b01110000; // 1299 : 112 - 0x70
      11'h514: dout  = 8'b00111000; // 1300 :  56 - 0x38
      11'h515: dout  = 8'b00111110; // 1301 :  62 - 0x3e
      11'h516: dout  = 8'b01111100; // 1302 : 124 - 0x7c
      11'h517: dout  = 8'b10111000; // 1303 : 184 - 0xb8
      11'h518: dout  = 8'b01010001; // 1304 :  81 - 0x51 -- Sprite 0xa3
      11'h519: dout  = 8'b00001010; // 1305 :  10 - 0xa
      11'h51A: dout  = 8'b00000100; // 1306 :   4 - 0x4
      11'h51B: dout  = 8'b11101010; // 1307 : 234 - 0xea
      11'h51C: dout  = 8'b01111001; // 1308 : 121 - 0x79
      11'h51D: dout  = 8'b01111111; // 1309 : 127 - 0x7f
      11'h51E: dout  = 8'b01110000; // 1310 : 112 - 0x70
      11'h51F: dout  = 8'b00111001; // 1311 :  57 - 0x39
      11'h520: dout  = 8'b01011000; // 1312 :  88 - 0x58 -- Sprite 0xa4
      11'h521: dout  = 8'b00111000; // 1313 :  56 - 0x38
      11'h522: dout  = 8'b00010000; // 1314 :  16 - 0x10
      11'h523: dout  = 8'b00110000; // 1315 :  48 - 0x30
      11'h524: dout  = 8'b11110000; // 1316 : 240 - 0xf0
      11'h525: dout  = 8'b11110000; // 1317 : 240 - 0xf0
      11'h526: dout  = 8'b11100000; // 1318 : 224 - 0xe0
      11'h527: dout  = 8'b11000000; // 1319 : 192 - 0xc0
      11'h528: dout  = 8'b00000000; // 1320 :   0 - 0x0 -- Sprite 0xa5
      11'h529: dout  = 8'b00001000; // 1321 :   8 - 0x8
      11'h52A: dout  = 8'b00011100; // 1322 :  28 - 0x1c
      11'h52B: dout  = 8'b00111100; // 1323 :  60 - 0x3c
      11'h52C: dout  = 8'b01111010; // 1324 : 122 - 0x7a
      11'h52D: dout  = 8'b01111010; // 1325 : 122 - 0x7a
      11'h52E: dout  = 8'b01111010; // 1326 : 122 - 0x7a
      11'h52F: dout  = 8'b01111110; // 1327 : 126 - 0x7e
      11'h530: dout  = 8'b00000000; // 1328 :   0 - 0x0 -- Sprite 0xa6
      11'h531: dout  = 8'b00000000; // 1329 :   0 - 0x0
      11'h532: dout  = 8'b00000000; // 1330 :   0 - 0x0
      11'h533: dout  = 8'b00010001; // 1331 :  17 - 0x11
      11'h534: dout  = 8'b00001010; // 1332 :  10 - 0xa
      11'h535: dout  = 8'b00110100; // 1333 :  52 - 0x34
      11'h536: dout  = 8'b00101010; // 1334 :  42 - 0x2a
      11'h537: dout  = 8'b01010001; // 1335 :  81 - 0x51
      11'h538: dout  = 8'b01111111; // 1336 : 127 - 0x7f -- Sprite 0xa7
      11'h539: dout  = 8'b01111101; // 1337 : 125 - 0x7d
      11'h53A: dout  = 8'b00111111; // 1338 :  63 - 0x3f
      11'h53B: dout  = 8'b00110111; // 1339 :  55 - 0x37
      11'h53C: dout  = 8'b00110011; // 1340 :  51 - 0x33
      11'h53D: dout  = 8'b00111011; // 1341 :  59 - 0x3b
      11'h53E: dout  = 8'b00111010; // 1342 :  58 - 0x3a
      11'h53F: dout  = 8'b01111000; // 1343 : 120 - 0x78
      11'h540: dout  = 8'b00100000; // 1344 :  32 - 0x20 -- Sprite 0xa8
      11'h541: dout  = 8'b01010001; // 1345 :  81 - 0x51
      11'h542: dout  = 8'b00001010; // 1346 :  10 - 0xa
      11'h543: dout  = 8'b00000100; // 1347 :   4 - 0x4
      11'h544: dout  = 8'b11101010; // 1348 : 234 - 0xea
      11'h545: dout  = 8'b00111001; // 1349 :  57 - 0x39
      11'h546: dout  = 8'b01111111; // 1350 : 127 - 0x7f
      11'h547: dout  = 8'b11110000; // 1351 : 240 - 0xf0
      11'h548: dout  = 8'b10111100; // 1352 : 188 - 0xbc -- Sprite 0xa9
      11'h549: dout  = 8'b01011000; // 1353 :  88 - 0x58
      11'h54A: dout  = 8'b00111000; // 1354 :  56 - 0x38
      11'h54B: dout  = 8'b00010000; // 1355 :  16 - 0x10
      11'h54C: dout  = 8'b00110000; // 1356 :  48 - 0x30
      11'h54D: dout  = 8'b11111000; // 1357 : 248 - 0xf8
      11'h54E: dout  = 8'b11111100; // 1358 : 252 - 0xfc
      11'h54F: dout  = 8'b00111110; // 1359 :  62 - 0x3e
      11'h550: dout  = 8'b00000000; // 1360 :   0 - 0x0 -- Sprite 0xaa
      11'h551: dout  = 8'b00000000; // 1361 :   0 - 0x0
      11'h552: dout  = 8'b00000000; // 1362 :   0 - 0x0
      11'h553: dout  = 8'b00000110; // 1363 :   6 - 0x6
      11'h554: dout  = 8'b00001110; // 1364 :  14 - 0xe
      11'h555: dout  = 8'b00001100; // 1365 :  12 - 0xc
      11'h556: dout  = 8'b00000000; // 1366 :   0 - 0x0
      11'h557: dout  = 8'b00000000; // 1367 :   0 - 0x0
      11'h558: dout  = 8'b00000000; // 1368 :   0 - 0x0 -- Sprite 0xab
      11'h559: dout  = 8'b00000000; // 1369 :   0 - 0x0
      11'h55A: dout  = 8'b00000000; // 1370 :   0 - 0x0
      11'h55B: dout  = 8'b00000000; // 1371 :   0 - 0x0
      11'h55C: dout  = 8'b00000000; // 1372 :   0 - 0x0
      11'h55D: dout  = 8'b00000000; // 1373 :   0 - 0x0
      11'h55E: dout  = 8'b00001111; // 1374 :  15 - 0xf
      11'h55F: dout  = 8'b00011000; // 1375 :  24 - 0x18
      11'h560: dout  = 8'b00000000; // 1376 :   0 - 0x0 -- Sprite 0xac
      11'h561: dout  = 8'b00000000; // 1377 :   0 - 0x0
      11'h562: dout  = 8'b00000000; // 1378 :   0 - 0x0
      11'h563: dout  = 8'b00000000; // 1379 :   0 - 0x0
      11'h564: dout  = 8'b11111000; // 1380 : 248 - 0xf8
      11'h565: dout  = 8'b00111110; // 1381 :  62 - 0x3e
      11'h566: dout  = 8'b00111011; // 1382 :  59 - 0x3b
      11'h567: dout  = 8'b00011000; // 1383 :  24 - 0x18
      11'h568: dout  = 8'b00010000; // 1384 :  16 - 0x10 -- Sprite 0xad
      11'h569: dout  = 8'b00010100; // 1385 :  20 - 0x14
      11'h56A: dout  = 8'b00010000; // 1386 :  16 - 0x10
      11'h56B: dout  = 8'b00010000; // 1387 :  16 - 0x10
      11'h56C: dout  = 8'b00111000; // 1388 :  56 - 0x38
      11'h56D: dout  = 8'b01111000; // 1389 : 120 - 0x78
      11'h56E: dout  = 8'b11111000; // 1390 : 248 - 0xf8
      11'h56F: dout  = 8'b00110000; // 1391 :  48 - 0x30
      11'h570: dout  = 8'b00000000; // 1392 :   0 - 0x0 -- Sprite 0xae
      11'h571: dout  = 8'b00000000; // 1393 :   0 - 0x0
      11'h572: dout  = 8'b00000000; // 1394 :   0 - 0x0
      11'h573: dout  = 8'b00000000; // 1395 :   0 - 0x0
      11'h574: dout  = 8'b00000110; // 1396 :   6 - 0x6
      11'h575: dout  = 8'b00001110; // 1397 :  14 - 0xe
      11'h576: dout  = 8'b00001100; // 1398 :  12 - 0xc
      11'h577: dout  = 8'b00000000; // 1399 :   0 - 0x0
      11'h578: dout  = 8'b00000000; // 1400 :   0 - 0x0 -- Sprite 0xaf
      11'h579: dout  = 8'b00000000; // 1401 :   0 - 0x0
      11'h57A: dout  = 8'b00000000; // 1402 :   0 - 0x0
      11'h57B: dout  = 8'b00000000; // 1403 :   0 - 0x0
      11'h57C: dout  = 8'b00000000; // 1404 :   0 - 0x0
      11'h57D: dout  = 8'b00000000; // 1405 :   0 - 0x0
      11'h57E: dout  = 8'b00000000; // 1406 :   0 - 0x0
      11'h57F: dout  = 8'b00001111; // 1407 :  15 - 0xf
      11'h580: dout  = 8'b00000000; // 1408 :   0 - 0x0 -- Sprite 0xb0
      11'h581: dout  = 8'b00000000; // 1409 :   0 - 0x0
      11'h582: dout  = 8'b00000000; // 1410 :   0 - 0x0
      11'h583: dout  = 8'b00000000; // 1411 :   0 - 0x0
      11'h584: dout  = 8'b00000000; // 1412 :   0 - 0x0
      11'h585: dout  = 8'b11111000; // 1413 : 248 - 0xf8
      11'h586: dout  = 8'b01111110; // 1414 : 126 - 0x7e
      11'h587: dout  = 8'b11110011; // 1415 : 243 - 0xf3
      11'h588: dout  = 8'b00011000; // 1416 :  24 - 0x18 -- Sprite 0xb1
      11'h589: dout  = 8'b00010000; // 1417 :  16 - 0x10
      11'h58A: dout  = 8'b00010100; // 1418 :  20 - 0x14
      11'h58B: dout  = 8'b00010000; // 1419 :  16 - 0x10
      11'h58C: dout  = 8'b00010000; // 1420 :  16 - 0x10
      11'h58D: dout  = 8'b00111000; // 1421 :  56 - 0x38
      11'h58E: dout  = 8'b01111100; // 1422 : 124 - 0x7c
      11'h58F: dout  = 8'b11011110; // 1423 : 222 - 0xde
      11'h590: dout  = 8'b00000000; // 1424 :   0 - 0x0 -- Sprite 0xb2
      11'h591: dout  = 8'b00001101; // 1425 :  13 - 0xd
      11'h592: dout  = 8'b00011110; // 1426 :  30 - 0x1e
      11'h593: dout  = 8'b00011110; // 1427 :  30 - 0x1e
      11'h594: dout  = 8'b00011110; // 1428 :  30 - 0x1e
      11'h595: dout  = 8'b00011111; // 1429 :  31 - 0x1f
      11'h596: dout  = 8'b00001111; // 1430 :  15 - 0xf
      11'h597: dout  = 8'b00000111; // 1431 :   7 - 0x7
      11'h598: dout  = 8'b01111000; // 1432 : 120 - 0x78 -- Sprite 0xb3
      11'h599: dout  = 8'b11110000; // 1433 : 240 - 0xf0
      11'h59A: dout  = 8'b00000000; // 1434 :   0 - 0x0
      11'h59B: dout  = 8'b00011010; // 1435 :  26 - 0x1a
      11'h59C: dout  = 8'b00111111; // 1436 :  63 - 0x3f
      11'h59D: dout  = 8'b00110101; // 1437 :  53 - 0x35
      11'h59E: dout  = 8'b00110101; // 1438 :  53 - 0x35
      11'h59F: dout  = 8'b00111111; // 1439 :  63 - 0x3f
      11'h5A0: dout  = 8'b00000000; // 1440 :   0 - 0x0 -- Sprite 0xb4
      11'h5A1: dout  = 8'b00000000; // 1441 :   0 - 0x0
      11'h5A2: dout  = 8'b10000000; // 1442 : 128 - 0x80
      11'h5A3: dout  = 8'b11100000; // 1443 : 224 - 0xe0
      11'h5A4: dout  = 8'b11100000; // 1444 : 224 - 0xe0
      11'h5A5: dout  = 8'b01110000; // 1445 : 112 - 0x70
      11'h5A6: dout  = 8'b01110011; // 1446 : 115 - 0x73
      11'h5A7: dout  = 8'b00100001; // 1447 :  33 - 0x21
      11'h5A8: dout  = 8'b00011010; // 1448 :  26 - 0x1a -- Sprite 0xb5
      11'h5A9: dout  = 8'b00000111; // 1449 :   7 - 0x7
      11'h5AA: dout  = 8'b00001100; // 1450 :  12 - 0xc
      11'h5AB: dout  = 8'b00011000; // 1451 :  24 - 0x18
      11'h5AC: dout  = 8'b01111000; // 1452 : 120 - 0x78
      11'h5AD: dout  = 8'b11111110; // 1453 : 254 - 0xfe
      11'h5AE: dout  = 8'b11111100; // 1454 : 252 - 0xfc
      11'h5AF: dout  = 8'b11110000; // 1455 : 240 - 0xf0
      11'h5B0: dout  = 8'b00000000; // 1456 :   0 - 0x0 -- Sprite 0xb6
      11'h5B1: dout  = 8'b00000001; // 1457 :   1 - 0x1
      11'h5B2: dout  = 8'b00000010; // 1458 :   2 - 0x2
      11'h5B3: dout  = 8'b00000000; // 1459 :   0 - 0x0
      11'h5B4: dout  = 8'b00111000; // 1460 :  56 - 0x38
      11'h5B5: dout  = 8'b01111100; // 1461 : 124 - 0x7c
      11'h5B6: dout  = 8'b01111110; // 1462 : 126 - 0x7e
      11'h5B7: dout  = 8'b00111111; // 1463 :  63 - 0x3f
      11'h5B8: dout  = 8'b00111111; // 1464 :  63 - 0x3f -- Sprite 0xb7
      11'h5B9: dout  = 8'b01000000; // 1465 :  64 - 0x40
      11'h5BA: dout  = 8'b01100000; // 1466 :  96 - 0x60
      11'h5BB: dout  = 8'b01100000; // 1467 :  96 - 0x60
      11'h5BC: dout  = 8'b00100000; // 1468 :  32 - 0x20
      11'h5BD: dout  = 8'b00110000; // 1469 :  48 - 0x30
      11'h5BE: dout  = 8'b00010011; // 1470 :  19 - 0x13
      11'h5BF: dout  = 8'b00000001; // 1471 :   1 - 0x1
      11'h5C0: dout  = 8'b11000000; // 1472 : 192 - 0xc0 -- Sprite 0xb8
      11'h5C1: dout  = 8'b11100000; // 1473 : 224 - 0xe0
      11'h5C2: dout  = 8'b00110000; // 1474 :  48 - 0x30
      11'h5C3: dout  = 8'b11010000; // 1475 : 208 - 0xd0
      11'h5C4: dout  = 8'b11010000; // 1476 : 208 - 0xd0
      11'h5C5: dout  = 8'b11010000; // 1477 : 208 - 0xd0
      11'h5C6: dout  = 8'b11010000; // 1478 : 208 - 0xd0
      11'h5C7: dout  = 8'b00000000; // 1479 :   0 - 0x0
      11'h5C8: dout  = 8'b00000111; // 1480 :   7 - 0x7 -- Sprite 0xb9
      11'h5C9: dout  = 8'b00001111; // 1481 :  15 - 0xf
      11'h5CA: dout  = 8'b00000010; // 1482 :   2 - 0x2
      11'h5CB: dout  = 8'b00011101; // 1483 :  29 - 0x1d
      11'h5CC: dout  = 8'b00011111; // 1484 :  31 - 0x1f
      11'h5CD: dout  = 8'b00011010; // 1485 :  26 - 0x1a
      11'h5CE: dout  = 8'b00011010; // 1486 :  26 - 0x1a
      11'h5CF: dout  = 8'b00000010; // 1487 :   2 - 0x2
      11'h5D0: dout  = 8'b00111000; // 1488 :  56 - 0x38 -- Sprite 0xba
      11'h5D1: dout  = 8'b01111100; // 1489 : 124 - 0x7c
      11'h5D2: dout  = 8'b11111100; // 1490 : 252 - 0xfc
      11'h5D3: dout  = 8'b11111100; // 1491 : 252 - 0xfc
      11'h5D4: dout  = 8'b11111100; // 1492 : 252 - 0xfc
      11'h5D5: dout  = 8'b11111110; // 1493 : 254 - 0xfe
      11'h5D6: dout  = 8'b10111110; // 1494 : 190 - 0xbe
      11'h5D7: dout  = 8'b10111110; // 1495 : 190 - 0xbe
      11'h5D8: dout  = 8'b00011100; // 1496 :  28 - 0x1c -- Sprite 0xbb
      11'h5D9: dout  = 8'b00111110; // 1497 :  62 - 0x3e
      11'h5DA: dout  = 8'b00111111; // 1498 :  63 - 0x3f
      11'h5DB: dout  = 8'b00111111; // 1499 :  63 - 0x3f
      11'h5DC: dout  = 8'b00111111; // 1500 :  63 - 0x3f
      11'h5DD: dout  = 8'b01111111; // 1501 : 127 - 0x7f
      11'h5DE: dout  = 8'b01111101; // 1502 : 125 - 0x7d
      11'h5DF: dout  = 8'b01111101; // 1503 : 125 - 0x7d
      11'h5E0: dout  = 8'b01111101; // 1504 : 125 - 0x7d -- Sprite 0xbc
      11'h5E1: dout  = 8'b01111111; // 1505 : 127 - 0x7f
      11'h5E2: dout  = 8'b01011111; // 1506 :  95 - 0x5f
      11'h5E3: dout  = 8'b00111011; // 1507 :  59 - 0x3b
      11'h5E4: dout  = 8'b00111100; // 1508 :  60 - 0x3c
      11'h5E5: dout  = 8'b00111111; // 1509 :  63 - 0x3f
      11'h5E6: dout  = 8'b00011110; // 1510 :  30 - 0x1e
      11'h5E7: dout  = 8'b00000000; // 1511 :   0 - 0x0
      11'h5E8: dout  = 8'b00011100; // 1512 :  28 - 0x1c -- Sprite 0xbd
      11'h5E9: dout  = 8'b00111110; // 1513 :  62 - 0x3e
      11'h5EA: dout  = 8'b00111111; // 1514 :  63 - 0x3f
      11'h5EB: dout  = 8'b00011111; // 1515 :  31 - 0x1f
      11'h5EC: dout  = 8'b00111111; // 1516 :  63 - 0x3f
      11'h5ED: dout  = 8'b01111111; // 1517 : 127 - 0x7f
      11'h5EE: dout  = 8'b01111101; // 1518 : 125 - 0x7d
      11'h5EF: dout  = 8'b01111101; // 1519 : 125 - 0x7d
      11'h5F0: dout  = 8'b00000000; // 1520 :   0 - 0x0 -- Sprite 0xbe
      11'h5F1: dout  = 8'b00000000; // 1521 :   0 - 0x0
      11'h5F2: dout  = 8'b00000000; // 1522 :   0 - 0x0
      11'h5F3: dout  = 8'b01100000; // 1523 :  96 - 0x60
      11'h5F4: dout  = 8'b01100010; // 1524 :  98 - 0x62
      11'h5F5: dout  = 8'b01100101; // 1525 : 101 - 0x65
      11'h5F6: dout  = 8'b00111111; // 1526 :  63 - 0x3f
      11'h5F7: dout  = 8'b00011111; // 1527 :  31 - 0x1f
      11'h5F8: dout  = 8'b01110000; // 1528 : 112 - 0x70 -- Sprite 0xbf
      11'h5F9: dout  = 8'b00111100; // 1529 :  60 - 0x3c
      11'h5FA: dout  = 8'b00111100; // 1530 :  60 - 0x3c
      11'h5FB: dout  = 8'b00011000; // 1531 :  24 - 0x18
      11'h5FC: dout  = 8'b00000000; // 1532 :   0 - 0x0
      11'h5FD: dout  = 8'b00000000; // 1533 :   0 - 0x0
      11'h5FE: dout  = 8'b00000010; // 1534 :   2 - 0x2
      11'h5FF: dout  = 8'b00000111; // 1535 :   7 - 0x7
      11'h600: dout  = 8'b11001111; // 1536 : 207 - 0xcf -- Sprite 0xc0
      11'h601: dout  = 8'b01111010; // 1537 : 122 - 0x7a
      11'h602: dout  = 8'b01011010; // 1538 :  90 - 0x5a
      11'h603: dout  = 8'b00010000; // 1539 :  16 - 0x10
      11'h604: dout  = 8'b00000000; // 1540 :   0 - 0x0
      11'h605: dout  = 8'b00000000; // 1541 :   0 - 0x0
      11'h606: dout  = 8'b11000000; // 1542 : 192 - 0xc0
      11'h607: dout  = 8'b10000000; // 1543 : 128 - 0x80
      11'h608: dout  = 8'b10000101; // 1544 : 133 - 0x85 -- Sprite 0xc1
      11'h609: dout  = 8'b10000100; // 1545 : 132 - 0x84
      11'h60A: dout  = 8'b10000110; // 1546 : 134 - 0x86
      11'h60B: dout  = 8'b11000110; // 1547 : 198 - 0xc6
      11'h60C: dout  = 8'b11100111; // 1548 : 231 - 0xe7
      11'h60D: dout  = 8'b01110011; // 1549 : 115 - 0x73
      11'h60E: dout  = 8'b01110011; // 1550 : 115 - 0x73
      11'h60F: dout  = 8'b11100001; // 1551 : 225 - 0xe1
      11'h610: dout  = 8'b10000000; // 1552 : 128 - 0x80 -- Sprite 0xc2
      11'h611: dout  = 8'b01001110; // 1553 :  78 - 0x4e
      11'h612: dout  = 8'b01110111; // 1554 : 119 - 0x77
      11'h613: dout  = 8'b11110011; // 1555 : 243 - 0xf3
      11'h614: dout  = 8'b11111011; // 1556 : 251 - 0xfb
      11'h615: dout  = 8'b11111001; // 1557 : 249 - 0xf9
      11'h616: dout  = 8'b11111010; // 1558 : 250 - 0xfa
      11'h617: dout  = 8'b01111000; // 1559 : 120 - 0x78
      11'h618: dout  = 8'b00010001; // 1560 :  17 - 0x11 -- Sprite 0xc3
      11'h619: dout  = 8'b00111001; // 1561 :  57 - 0x39
      11'h61A: dout  = 8'b01111101; // 1562 : 125 - 0x7d
      11'h61B: dout  = 8'b00111001; // 1563 :  57 - 0x39
      11'h61C: dout  = 8'b00000000; // 1564 :   0 - 0x0
      11'h61D: dout  = 8'b00000000; // 1565 :   0 - 0x0
      11'h61E: dout  = 8'b11100000; // 1566 : 224 - 0xe0
      11'h61F: dout  = 8'b11100111; // 1567 : 231 - 0xe7
      11'h620: dout  = 8'b00000000; // 1568 :   0 - 0x0 -- Sprite 0xc4
      11'h621: dout  = 8'b00000000; // 1569 :   0 - 0x0
      11'h622: dout  = 8'b00000111; // 1570 :   7 - 0x7
      11'h623: dout  = 8'b00000111; // 1571 :   7 - 0x7
      11'h624: dout  = 8'b00010110; // 1572 :  22 - 0x16
      11'h625: dout  = 8'b00010000; // 1573 :  16 - 0x10
      11'h626: dout  = 8'b00000000; // 1574 :   0 - 0x0
      11'h627: dout  = 8'b00111000; // 1575 :  56 - 0x38
      11'h628: dout  = 8'b11001111; // 1576 : 207 - 0xcf -- Sprite 0xc5
      11'h629: dout  = 8'b00011111; // 1577 :  31 - 0x1f
      11'h62A: dout  = 8'b00010111; // 1578 :  23 - 0x17
      11'h62B: dout  = 8'b00010000; // 1579 :  16 - 0x10
      11'h62C: dout  = 8'b00110011; // 1580 :  51 - 0x33
      11'h62D: dout  = 8'b00110000; // 1581 :  48 - 0x30
      11'h62E: dout  = 8'b00110000; // 1582 :  48 - 0x30
      11'h62F: dout  = 8'b00100000; // 1583 :  32 - 0x20
      11'h630: dout  = 8'b00111000; // 1584 :  56 - 0x38 -- Sprite 0xc6
      11'h631: dout  = 8'b00110000; // 1585 :  48 - 0x30
      11'h632: dout  = 8'b01000000; // 1586 :  64 - 0x40
      11'h633: dout  = 8'b11000111; // 1587 : 199 - 0xc7
      11'h634: dout  = 8'b00000111; // 1588 :   7 - 0x7
      11'h635: dout  = 8'b01100110; // 1589 : 102 - 0x66
      11'h636: dout  = 8'b11100000; // 1590 : 224 - 0xe0
      11'h637: dout  = 8'b01101100; // 1591 : 108 - 0x6c
      11'h638: dout  = 8'b01100000; // 1592 :  96 - 0x60 -- Sprite 0xc7
      11'h639: dout  = 8'b11000000; // 1593 : 192 - 0xc0
      11'h63A: dout  = 8'b10000000; // 1594 : 128 - 0x80
      11'h63B: dout  = 8'b00000100; // 1595 :   4 - 0x4
      11'h63C: dout  = 8'b10011110; // 1596 : 158 - 0x9e
      11'h63D: dout  = 8'b11111111; // 1597 : 255 - 0xff
      11'h63E: dout  = 8'b11110000; // 1598 : 240 - 0xf0
      11'h63F: dout  = 8'b11111000; // 1599 : 248 - 0xf8
      11'h640: dout  = 8'b00100100; // 1600 :  36 - 0x24 -- Sprite 0xc8
      11'h641: dout  = 8'b00000001; // 1601 :   1 - 0x1
      11'h642: dout  = 8'b00000111; // 1602 :   7 - 0x7
      11'h643: dout  = 8'b11111110; // 1603 : 254 - 0xfe
      11'h644: dout  = 8'b11111111; // 1604 : 255 - 0xff
      11'h645: dout  = 8'b01111111; // 1605 : 127 - 0x7f
      11'h646: dout  = 8'b00111111; // 1606 :  63 - 0x3f
      11'h647: dout  = 8'b01111111; // 1607 : 127 - 0x7f
      11'h648: dout  = 8'b11001111; // 1608 : 207 - 0xcf -- Sprite 0xc9
      11'h649: dout  = 8'b01111010; // 1609 : 122 - 0x7a
      11'h64A: dout  = 8'b00001010; // 1610 :  10 - 0xa
      11'h64B: dout  = 8'b11111110; // 1611 : 254 - 0xfe
      11'h64C: dout  = 8'b11111100; // 1612 : 252 - 0xfc
      11'h64D: dout  = 8'b00000000; // 1613 :   0 - 0x0
      11'h64E: dout  = 8'b00000000; // 1614 :   0 - 0x0
      11'h64F: dout  = 8'b00000000; // 1615 :   0 - 0x0
      11'h650: dout  = 8'b10000101; // 1616 : 133 - 0x85 -- Sprite 0xca
      11'h651: dout  = 8'b10000110; // 1617 : 134 - 0x86
      11'h652: dout  = 8'b10000011; // 1618 : 131 - 0x83
      11'h653: dout  = 8'b11000011; // 1619 : 195 - 0xc3
      11'h654: dout  = 8'b11100001; // 1620 : 225 - 0xe1
      11'h655: dout  = 8'b01110000; // 1621 : 112 - 0x70
      11'h656: dout  = 8'b01110000; // 1622 : 112 - 0x70
      11'h657: dout  = 8'b11100000; // 1623 : 224 - 0xe0
      11'h658: dout  = 8'b01100000; // 1624 :  96 - 0x60 -- Sprite 0xcb
      11'h659: dout  = 8'b11000000; // 1625 : 192 - 0xc0
      11'h65A: dout  = 8'b10000000; // 1626 : 128 - 0x80
      11'h65B: dout  = 8'b00000000; // 1627 :   0 - 0x0
      11'h65C: dout  = 8'b10011000; // 1628 : 152 - 0x98
      11'h65D: dout  = 8'b11111100; // 1629 : 252 - 0xfc
      11'h65E: dout  = 8'b11111110; // 1630 : 254 - 0xfe
      11'h65F: dout  = 8'b11111111; // 1631 : 255 - 0xff
      11'h660: dout  = 8'b00100100; // 1632 :  36 - 0x24 -- Sprite 0xcc
      11'h661: dout  = 8'b00000000; // 1633 :   0 - 0x0
      11'h662: dout  = 8'b00000111; // 1634 :   7 - 0x7
      11'h663: dout  = 8'b11111110; // 1635 : 254 - 0xfe
      11'h664: dout  = 8'b11111111; // 1636 : 255 - 0xff
      11'h665: dout  = 8'b01111111; // 1637 : 127 - 0x7f
      11'h666: dout  = 8'b11111111; // 1638 : 255 - 0xff
      11'h667: dout  = 8'b00000011; // 1639 :   3 - 0x3
      11'h668: dout  = 8'b00000011; // 1640 :   3 - 0x3 -- Sprite 0xcd
      11'h669: dout  = 8'b00001111; // 1641 :  15 - 0xf
      11'h66A: dout  = 8'b00100011; // 1642 :  35 - 0x23
      11'h66B: dout  = 8'b01100010; // 1643 :  98 - 0x62
      11'h66C: dout  = 8'b01100100; // 1644 : 100 - 0x64
      11'h66D: dout  = 8'b00111100; // 1645 :  60 - 0x3c
      11'h66E: dout  = 8'b00011100; // 1646 :  28 - 0x1c
      11'h66F: dout  = 8'b00011110; // 1647 :  30 - 0x1e
      11'h670: dout  = 8'b00011111; // 1648 :  31 - 0x1f -- Sprite 0xce
      11'h671: dout  = 8'b00111101; // 1649 :  61 - 0x3d
      11'h672: dout  = 8'b01101101; // 1650 : 109 - 0x6d
      11'h673: dout  = 8'b01001111; // 1651 :  79 - 0x4f
      11'h674: dout  = 8'b11101110; // 1652 : 238 - 0xee
      11'h675: dout  = 8'b11110011; // 1653 : 243 - 0xf3
      11'h676: dout  = 8'b00100000; // 1654 :  32 - 0x20
      11'h677: dout  = 8'b00000011; // 1655 :   3 - 0x3
      11'h678: dout  = 8'b00000111; // 1656 :   7 - 0x7 -- Sprite 0xcf
      11'h679: dout  = 8'b00000111; // 1657 :   7 - 0x7
      11'h67A: dout  = 8'b00011111; // 1658 :  31 - 0x1f
      11'h67B: dout  = 8'b00111111; // 1659 :  63 - 0x3f
      11'h67C: dout  = 8'b00001111; // 1660 :  15 - 0xf
      11'h67D: dout  = 8'b01000111; // 1661 :  71 - 0x47
      11'h67E: dout  = 8'b00000011; // 1662 :   3 - 0x3
      11'h67F: dout  = 8'b00000000; // 1663 :   0 - 0x0
      11'h680: dout  = 8'b00000000; // 1664 :   0 - 0x0 -- Sprite 0xd0
      11'h681: dout  = 8'b00000000; // 1665 :   0 - 0x0
      11'h682: dout  = 8'b00000011; // 1666 :   3 - 0x3
      11'h683: dout  = 8'b00000111; // 1667 :   7 - 0x7
      11'h684: dout  = 8'b00001111; // 1668 :  15 - 0xf
      11'h685: dout  = 8'b00001111; // 1669 :  15 - 0xf
      11'h686: dout  = 8'b00011111; // 1670 :  31 - 0x1f
      11'h687: dout  = 8'b00011111; // 1671 :  31 - 0x1f
      11'h688: dout  = 8'b00000000; // 1672 :   0 - 0x0 -- Sprite 0xd1
      11'h689: dout  = 8'b00100011; // 1673 :  35 - 0x23
      11'h68A: dout  = 8'b01010111; // 1674 :  87 - 0x57
      11'h68B: dout  = 8'b01001111; // 1675 :  79 - 0x4f
      11'h68C: dout  = 8'b01010111; // 1676 :  87 - 0x57
      11'h68D: dout  = 8'b00101111; // 1677 :  47 - 0x2f
      11'h68E: dout  = 8'b11011111; // 1678 : 223 - 0xdf
      11'h68F: dout  = 8'b00100001; // 1679 :  33 - 0x21
      11'h690: dout  = 8'b00000000; // 1680 :   0 - 0x0 -- Sprite 0xd2
      11'h691: dout  = 8'b00000000; // 1681 :   0 - 0x0
      11'h692: dout  = 8'b00000000; // 1682 :   0 - 0x0
      11'h693: dout  = 8'b00000000; // 1683 :   0 - 0x0
      11'h694: dout  = 8'b10000000; // 1684 : 128 - 0x80
      11'h695: dout  = 8'b10000000; // 1685 : 128 - 0x80
      11'h696: dout  = 8'b00000000; // 1686 :   0 - 0x0
      11'h697: dout  = 8'b00000000; // 1687 :   0 - 0x0
      11'h698: dout  = 8'b00100011; // 1688 :  35 - 0x23 -- Sprite 0xd3
      11'h699: dout  = 8'b00001111; // 1689 :  15 - 0xf
      11'h69A: dout  = 8'b00011110; // 1690 :  30 - 0x1e
      11'h69B: dout  = 8'b11110000; // 1691 : 240 - 0xf0
      11'h69C: dout  = 8'b00011100; // 1692 :  28 - 0x1c
      11'h69D: dout  = 8'b00111111; // 1693 :  63 - 0x3f
      11'h69E: dout  = 8'b00011111; // 1694 :  31 - 0x1f
      11'h69F: dout  = 8'b00011110; // 1695 :  30 - 0x1e
      11'h6A0: dout  = 8'b00000000; // 1696 :   0 - 0x0 -- Sprite 0xd4
      11'h6A1: dout  = 8'b10000000; // 1697 : 128 - 0x80
      11'h6A2: dout  = 8'b00011000; // 1698 :  24 - 0x18
      11'h6A3: dout  = 8'b00110000; // 1699 :  48 - 0x30
      11'h6A4: dout  = 8'b00110100; // 1700 :  52 - 0x34
      11'h6A5: dout  = 8'b11111110; // 1701 : 254 - 0xfe
      11'h6A6: dout  = 8'b11111110; // 1702 : 254 - 0xfe
      11'h6A7: dout  = 8'b11111110; // 1703 : 254 - 0xfe
      11'h6A8: dout  = 8'b00000000; // 1704 :   0 - 0x0 -- Sprite 0xd5
      11'h6A9: dout  = 8'b00000000; // 1705 :   0 - 0x0
      11'h6AA: dout  = 8'b00000001; // 1706 :   1 - 0x1
      11'h6AB: dout  = 8'b00000100; // 1707 :   4 - 0x4
      11'h6AC: dout  = 8'b00000110; // 1708 :   6 - 0x6
      11'h6AD: dout  = 8'b00000110; // 1709 :   6 - 0x6
      11'h6AE: dout  = 8'b00000111; // 1710 :   7 - 0x7
      11'h6AF: dout  = 8'b00000111; // 1711 :   7 - 0x7
      11'h6B0: dout  = 8'b00001111; // 1712 :  15 - 0xf -- Sprite 0xd6
      11'h6B1: dout  = 8'b00111111; // 1713 :  63 - 0x3f
      11'h6B2: dout  = 8'b01111111; // 1714 : 127 - 0x7f
      11'h6B3: dout  = 8'b11111000; // 1715 : 248 - 0xf8
      11'h6B4: dout  = 8'b11111000; // 1716 : 248 - 0xf8
      11'h6B5: dout  = 8'b01111111; // 1717 : 127 - 0x7f
      11'h6B6: dout  = 8'b00111111; // 1718 :  63 - 0x3f
      11'h6B7: dout  = 8'b00001111; // 1719 :  15 - 0xf
      11'h6B8: dout  = 8'b00011111; // 1720 :  31 - 0x1f -- Sprite 0xd7
      11'h6B9: dout  = 8'b00011111; // 1721 :  31 - 0x1f
      11'h6BA: dout  = 8'b00011111; // 1722 :  31 - 0x1f
      11'h6BB: dout  = 8'b00001011; // 1723 :  11 - 0xb
      11'h6BC: dout  = 8'b00000001; // 1724 :   1 - 0x1
      11'h6BD: dout  = 8'b00000001; // 1725 :   1 - 0x1
      11'h6BE: dout  = 8'b00000000; // 1726 :   0 - 0x0
      11'h6BF: dout  = 8'b00000000; // 1727 :   0 - 0x0
      11'h6C0: dout  = 8'b00000011; // 1728 :   3 - 0x3 -- Sprite 0xd8
      11'h6C1: dout  = 8'b00011111; // 1729 :  31 - 0x1f
      11'h6C2: dout  = 8'b00111111; // 1730 :  63 - 0x3f
      11'h6C3: dout  = 8'b00111111; // 1731 :  63 - 0x3f
      11'h6C4: dout  = 8'b01111000; // 1732 : 120 - 0x78
      11'h6C5: dout  = 8'b00000000; // 1733 :   0 - 0x0
      11'h6C6: dout  = 8'b00000011; // 1734 :   3 - 0x3
      11'h6C7: dout  = 8'b11111111; // 1735 : 255 - 0xff
      11'h6C8: dout  = 8'b00000000; // 1736 :   0 - 0x0 -- Sprite 0xd9
      11'h6C9: dout  = 8'b00000000; // 1737 :   0 - 0x0
      11'h6CA: dout  = 8'b00000000; // 1738 :   0 - 0x0
      11'h6CB: dout  = 8'b00000000; // 1739 :   0 - 0x0
      11'h6CC: dout  = 8'b00000000; // 1740 :   0 - 0x0
      11'h6CD: dout  = 8'b00000000; // 1741 :   0 - 0x0
      11'h6CE: dout  = 8'b00000000; // 1742 :   0 - 0x0
      11'h6CF: dout  = 8'b00000000; // 1743 :   0 - 0x0
      11'h6D0: dout  = 8'b00100011; // 1744 :  35 - 0x23 -- Sprite 0xda
      11'h6D1: dout  = 8'b00100111; // 1745 :  39 - 0x27
      11'h6D2: dout  = 8'b00011111; // 1746 :  31 - 0x1f
      11'h6D3: dout  = 8'b00000111; // 1747 :   7 - 0x7
      11'h6D4: dout  = 8'b00001111; // 1748 :  15 - 0xf
      11'h6D5: dout  = 8'b00011111; // 1749 :  31 - 0x1f
      11'h6D6: dout  = 8'b01111111; // 1750 : 127 - 0x7f
      11'h6D7: dout  = 8'b00111111; // 1751 :  63 - 0x3f
      11'h6D8: dout  = 8'b11100000; // 1752 : 224 - 0xe0 -- Sprite 0xdb
      11'h6D9: dout  = 8'b10000000; // 1753 : 128 - 0x80
      11'h6DA: dout  = 8'b10000000; // 1754 : 128 - 0x80
      11'h6DB: dout  = 8'b01000000; // 1755 :  64 - 0x40
      11'h6DC: dout  = 8'b11100000; // 1756 : 224 - 0xe0
      11'h6DD: dout  = 8'b11100000; // 1757 : 224 - 0xe0
      11'h6DE: dout  = 8'b11100000; // 1758 : 224 - 0xe0
      11'h6DF: dout  = 8'b11000000; // 1759 : 192 - 0xc0
      11'h6E0: dout  = 8'b00000011; // 1760 :   3 - 0x3 -- Sprite 0xdc
      11'h6E1: dout  = 8'b00000111; // 1761 :   7 - 0x7
      11'h6E2: dout  = 8'b00001111; // 1762 :  15 - 0xf
      11'h6E3: dout  = 8'b00011111; // 1763 :  31 - 0x1f
      11'h6E4: dout  = 8'b00111111; // 1764 :  63 - 0x3f
      11'h6E5: dout  = 8'b01111111; // 1765 : 127 - 0x7f
      11'h6E6: dout  = 8'b11111111; // 1766 : 255 - 0xff
      11'h6E7: dout  = 8'b00011111; // 1767 :  31 - 0x1f
      11'h6E8: dout  = 8'b00011111; // 1768 :  31 - 0x1f -- Sprite 0xdd
      11'h6E9: dout  = 8'b00010000; // 1769 :  16 - 0x10
      11'h6EA: dout  = 8'b00001100; // 1770 :  12 - 0xc
      11'h6EB: dout  = 8'b00010010; // 1771 :  18 - 0x12
      11'h6EC: dout  = 8'b00010010; // 1772 :  18 - 0x12
      11'h6ED: dout  = 8'b00101100; // 1773 :  44 - 0x2c
      11'h6EE: dout  = 8'b00111111; // 1774 :  63 - 0x3f
      11'h6EF: dout  = 8'b00111111; // 1775 :  63 - 0x3f
      11'h6F0: dout  = 8'b00110111; // 1776 :  55 - 0x37 -- Sprite 0xde
      11'h6F1: dout  = 8'b00110110; // 1777 :  54 - 0x36
      11'h6F2: dout  = 8'b00110110; // 1778 :  54 - 0x36
      11'h6F3: dout  = 8'b00110110; // 1779 :  54 - 0x36
      11'h6F4: dout  = 8'b00010110; // 1780 :  22 - 0x16
      11'h6F5: dout  = 8'b00010110; // 1781 :  22 - 0x16
      11'h6F6: dout  = 8'b00010010; // 1782 :  18 - 0x12
      11'h6F7: dout  = 8'b00000010; // 1783 :   2 - 0x2
      11'h6F8: dout  = 8'b00010000; // 1784 :  16 - 0x10 -- Sprite 0xdf
      11'h6F9: dout  = 8'b01111110; // 1785 : 126 - 0x7e
      11'h6FA: dout  = 8'b11111111; // 1786 : 255 - 0xff
      11'h6FB: dout  = 8'b11111111; // 1787 : 255 - 0xff
      11'h6FC: dout  = 8'b11110110; // 1788 : 246 - 0xf6
      11'h6FD: dout  = 8'b01110110; // 1789 : 118 - 0x76
      11'h6FE: dout  = 8'b00111010; // 1790 :  58 - 0x3a
      11'h6FF: dout  = 8'b00011010; // 1791 :  26 - 0x1a
      11'h700: dout  = 8'b00000000; // 1792 :   0 - 0x0 -- Sprite 0xe0
      11'h701: dout  = 8'b00000000; // 1793 :   0 - 0x0
      11'h702: dout  = 8'b00111000; // 1794 :  56 - 0x38
      11'h703: dout  = 8'b00000100; // 1795 :   4 - 0x4
      11'h704: dout  = 8'b00000000; // 1796 :   0 - 0x0
      11'h705: dout  = 8'b00000000; // 1797 :   0 - 0x0
      11'h706: dout  = 8'b00000000; // 1798 :   0 - 0x0
      11'h707: dout  = 8'b00000000; // 1799 :   0 - 0x0
      11'h708: dout  = 8'b00000000; // 1800 :   0 - 0x0 -- Sprite 0xe1
      11'h709: dout  = 8'b00000000; // 1801 :   0 - 0x0
      11'h70A: dout  = 8'b00000000; // 1802 :   0 - 0x0
      11'h70B: dout  = 8'b00111000; // 1803 :  56 - 0x38
      11'h70C: dout  = 8'b01000000; // 1804 :  64 - 0x40
      11'h70D: dout  = 8'b00000000; // 1805 :   0 - 0x0
      11'h70E: dout  = 8'b00000000; // 1806 :   0 - 0x0
      11'h70F: dout  = 8'b00000000; // 1807 :   0 - 0x0
      11'h710: dout  = 8'b11111100; // 1808 : 252 - 0xfc -- Sprite 0xe2
      11'h711: dout  = 8'b10100000; // 1809 : 160 - 0xa0
      11'h712: dout  = 8'b10000000; // 1810 : 128 - 0x80
      11'h713: dout  = 8'b10000000; // 1811 : 128 - 0x80
      11'h714: dout  = 8'b00000000; // 1812 :   0 - 0x0
      11'h715: dout  = 8'b00000000; // 1813 :   0 - 0x0
      11'h716: dout  = 8'b00000000; // 1814 :   0 - 0x0
      11'h717: dout  = 8'b00000000; // 1815 :   0 - 0x0
      11'h718: dout  = 8'b00000111; // 1816 :   7 - 0x7 -- Sprite 0xe3
      11'h719: dout  = 8'b00100111; // 1817 :  39 - 0x27
      11'h71A: dout  = 8'b01010111; // 1818 :  87 - 0x57
      11'h71B: dout  = 8'b01001111; // 1819 :  79 - 0x4f
      11'h71C: dout  = 8'b01010111; // 1820 :  87 - 0x57
      11'h71D: dout  = 8'b00100111; // 1821 :  39 - 0x27
      11'h71E: dout  = 8'b11000001; // 1822 : 193 - 0xc1
      11'h71F: dout  = 8'b00100001; // 1823 :  33 - 0x21
      11'h720: dout  = 8'b00011101; // 1824 :  29 - 0x1d -- Sprite 0xe4
      11'h721: dout  = 8'b00001111; // 1825 :  15 - 0xf
      11'h722: dout  = 8'b00001111; // 1826 :  15 - 0xf
      11'h723: dout  = 8'b00011111; // 1827 :  31 - 0x1f
      11'h724: dout  = 8'b00011111; // 1828 :  31 - 0x1f
      11'h725: dout  = 8'b00011110; // 1829 :  30 - 0x1e
      11'h726: dout  = 8'b00111000; // 1830 :  56 - 0x38
      11'h727: dout  = 8'b00110000; // 1831 :  48 - 0x30
      11'h728: dout  = 8'b00000000; // 1832 :   0 - 0x0 -- Sprite 0xe5
      11'h729: dout  = 8'b00000000; // 1833 :   0 - 0x0
      11'h72A: dout  = 8'b00111000; // 1834 :  56 - 0x38
      11'h72B: dout  = 8'b00010000; // 1835 :  16 - 0x10
      11'h72C: dout  = 8'b01001100; // 1836 :  76 - 0x4c
      11'h72D: dout  = 8'b00011000; // 1837 :  24 - 0x18
      11'h72E: dout  = 8'b10000110; // 1838 : 134 - 0x86
      11'h72F: dout  = 8'b00100100; // 1839 :  36 - 0x24
      11'h730: dout  = 8'b00000000; // 1840 :   0 - 0x0 -- Sprite 0xe6
      11'h731: dout  = 8'b01000010; // 1841 :  66 - 0x42
      11'h732: dout  = 8'b00001010; // 1842 :  10 - 0xa
      11'h733: dout  = 8'b01000000; // 1843 :  64 - 0x40
      11'h734: dout  = 8'b00010000; // 1844 :  16 - 0x10
      11'h735: dout  = 8'b00000010; // 1845 :   2 - 0x2
      11'h736: dout  = 8'b00001000; // 1846 :   8 - 0x8
      11'h737: dout  = 8'b00000010; // 1847 :   2 - 0x2
      11'h738: dout  = 8'b00000000; // 1848 :   0 - 0x0 -- Sprite 0xe7
      11'h739: dout  = 8'b00000000; // 1849 :   0 - 0x0
      11'h73A: dout  = 8'b10000000; // 1850 : 128 - 0x80
      11'h73B: dout  = 8'b01000000; // 1851 :  64 - 0x40
      11'h73C: dout  = 8'b00001000; // 1852 :   8 - 0x8
      11'h73D: dout  = 8'b00001100; // 1853 :  12 - 0xc
      11'h73E: dout  = 8'b00001010; // 1854 :  10 - 0xa
      11'h73F: dout  = 8'b10000100; // 1855 : 132 - 0x84
      11'h740: dout  = 8'b00000000; // 1856 :   0 - 0x0 -- Sprite 0xe8
      11'h741: dout  = 8'b00000000; // 1857 :   0 - 0x0
      11'h742: dout  = 8'b11001111; // 1858 : 207 - 0xcf
      11'h743: dout  = 8'b00100000; // 1859 :  32 - 0x20
      11'h744: dout  = 8'b00100000; // 1860 :  32 - 0x20
      11'h745: dout  = 8'b00100000; // 1861 :  32 - 0x20
      11'h746: dout  = 8'b00100110; // 1862 :  38 - 0x26
      11'h747: dout  = 8'b00101110; // 1863 :  46 - 0x2e
      11'h748: dout  = 8'b11100000; // 1864 : 224 - 0xe0 -- Sprite 0xe9
      11'h749: dout  = 8'b11100000; // 1865 : 224 - 0xe0
      11'h74A: dout  = 8'b11000000; // 1866 : 192 - 0xc0
      11'h74B: dout  = 8'b00000000; // 1867 :   0 - 0x0
      11'h74C: dout  = 8'b00000000; // 1868 :   0 - 0x0
      11'h74D: dout  = 8'b00000000; // 1869 :   0 - 0x0
      11'h74E: dout  = 8'b00000000; // 1870 :   0 - 0x0
      11'h74F: dout  = 8'b00000000; // 1871 :   0 - 0x0
      11'h750: dout  = 8'b00101111; // 1872 :  47 - 0x2f -- Sprite 0xea
      11'h751: dout  = 8'b00100011; // 1873 :  35 - 0x23
      11'h752: dout  = 8'b00100001; // 1874 :  33 - 0x21
      11'h753: dout  = 8'b00100000; // 1875 :  32 - 0x20
      11'h754: dout  = 8'b00100000; // 1876 :  32 - 0x20
      11'h755: dout  = 8'b00000000; // 1877 :   0 - 0x0
      11'h756: dout  = 8'b00000000; // 1878 :   0 - 0x0
      11'h757: dout  = 8'b00000000; // 1879 :   0 - 0x0
      11'h758: dout  = 8'b11000001; // 1880 : 193 - 0xc1 -- Sprite 0xeb
      11'h759: dout  = 8'b10110001; // 1881 : 177 - 0xb1
      11'h75A: dout  = 8'b01011001; // 1882 :  89 - 0x59
      11'h75B: dout  = 8'b01101101; // 1883 : 109 - 0x6d
      11'h75C: dout  = 8'b00110101; // 1884 :  53 - 0x35
      11'h75D: dout  = 8'b00111011; // 1885 :  59 - 0x3b
      11'h75E: dout  = 8'b00011111; // 1886 :  31 - 0x1f
      11'h75F: dout  = 8'b00000011; // 1887 :   3 - 0x3
      11'h760: dout  = 8'b00000000; // 1888 :   0 - 0x0 -- Sprite 0xec
      11'h761: dout  = 8'b00000010; // 1889 :   2 - 0x2
      11'h762: dout  = 8'b00000000; // 1890 :   0 - 0x0
      11'h763: dout  = 8'b00001000; // 1891 :   8 - 0x8
      11'h764: dout  = 8'b00000010; // 1892 :   2 - 0x2
      11'h765: dout  = 8'b00000000; // 1893 :   0 - 0x0
      11'h766: dout  = 8'b00101000; // 1894 :  40 - 0x28
      11'h767: dout  = 8'b00000000; // 1895 :   0 - 0x0
      11'h768: dout  = 8'b00000100; // 1896 :   4 - 0x4 -- Sprite 0xed
      11'h769: dout  = 8'b00010000; // 1897 :  16 - 0x10
      11'h76A: dout  = 8'b00000010; // 1898 :   2 - 0x2
      11'h76B: dout  = 8'b00010000; // 1899 :  16 - 0x10
      11'h76C: dout  = 8'b00000100; // 1900 :   4 - 0x4
      11'h76D: dout  = 8'b00000000; // 1901 :   0 - 0x0
      11'h76E: dout  = 8'b00001010; // 1902 :  10 - 0xa
      11'h76F: dout  = 8'b00000000; // 1903 :   0 - 0x0
      11'h770: dout  = 8'b11000001; // 1904 : 193 - 0xc1 -- Sprite 0xee
      11'h771: dout  = 8'b10110001; // 1905 : 177 - 0xb1
      11'h772: dout  = 8'b01011001; // 1906 :  89 - 0x59
      11'h773: dout  = 8'b01101101; // 1907 : 109 - 0x6d
      11'h774: dout  = 8'b00110101; // 1908 :  53 - 0x35
      11'h775: dout  = 8'b00111011; // 1909 :  59 - 0x3b
      11'h776: dout  = 8'b00011111; // 1910 :  31 - 0x1f
      11'h777: dout  = 8'b00000011; // 1911 :   3 - 0x3
      11'h778: dout  = 8'b00000000; // 1912 :   0 - 0x0 -- Sprite 0xef
      11'h779: dout  = 8'b00001111; // 1913 :  15 - 0xf
      11'h77A: dout  = 8'b00011111; // 1914 :  31 - 0x1f
      11'h77B: dout  = 8'b11111111; // 1915 : 255 - 0xff
      11'h77C: dout  = 8'b11111100; // 1916 : 252 - 0xfc
      11'h77D: dout  = 8'b01100011; // 1917 :  99 - 0x63
      11'h77E: dout  = 8'b00011111; // 1918 :  31 - 0x1f
      11'h77F: dout  = 8'b00000011; // 1919 :   3 - 0x3
      11'h780: dout  = 8'b00000000; // 1920 :   0 - 0x0 -- Sprite 0xf0
      11'h781: dout  = 8'b00000000; // 1921 :   0 - 0x0
      11'h782: dout  = 8'b11111110; // 1922 : 254 - 0xfe
      11'h783: dout  = 8'b11000110; // 1923 : 198 - 0xc6
      11'h784: dout  = 8'b11000110; // 1924 : 198 - 0xc6
      11'h785: dout  = 8'b11111110; // 1925 : 254 - 0xfe
      11'h786: dout  = 8'b00000000; // 1926 :   0 - 0x0
      11'h787: dout  = 8'b00000000; // 1927 :   0 - 0x0
      11'h788: dout  = 8'b00000000; // 1928 :   0 - 0x0 -- Sprite 0xf1
      11'h789: dout  = 8'b00000000; // 1929 :   0 - 0x0
      11'h78A: dout  = 8'b00000110; // 1930 :   6 - 0x6
      11'h78B: dout  = 8'b00000110; // 1931 :   6 - 0x6
      11'h78C: dout  = 8'b00001100; // 1932 :  12 - 0xc
      11'h78D: dout  = 8'b00011000; // 1933 :  24 - 0x18
      11'h78E: dout  = 8'b01110000; // 1934 : 112 - 0x70
      11'h78F: dout  = 8'b01100000; // 1935 :  96 - 0x60
      11'h790: dout  = 8'b00000000; // 1936 :   0 - 0x0 -- Sprite 0xf2
      11'h791: dout  = 8'b00000000; // 1937 :   0 - 0x0
      11'h792: dout  = 8'b00000110; // 1938 :   6 - 0x6
      11'h793: dout  = 8'b00000110; // 1939 :   6 - 0x6
      11'h794: dout  = 8'b00000100; // 1940 :   4 - 0x4
      11'h795: dout  = 8'b00000100; // 1941 :   4 - 0x4
      11'h796: dout  = 8'b00001000; // 1942 :   8 - 0x8
      11'h797: dout  = 8'b00001000; // 1943 :   8 - 0x8
      11'h798: dout  = 8'b00001000; // 1944 :   8 - 0x8 -- Sprite 0xf3
      11'h799: dout  = 8'b00010000; // 1945 :  16 - 0x10
      11'h79A: dout  = 8'b00110000; // 1946 :  48 - 0x30
      11'h79B: dout  = 8'b00110000; // 1947 :  48 - 0x30
      11'h79C: dout  = 8'b00110000; // 1948 :  48 - 0x30
      11'h79D: dout  = 8'b00110000; // 1949 :  48 - 0x30
      11'h79E: dout  = 8'b00010000; // 1950 :  16 - 0x10
      11'h79F: dout  = 8'b00001000; // 1951 :   8 - 0x8
      11'h7A0: dout  = 8'b00000000; // 1952 :   0 - 0x0 -- Sprite 0xf4
      11'h7A1: dout  = 8'b00000000; // 1953 :   0 - 0x0
      11'h7A2: dout  = 8'b00000001; // 1954 :   1 - 0x1
      11'h7A3: dout  = 8'b00000011; // 1955 :   3 - 0x3
      11'h7A4: dout  = 8'b00000001; // 1956 :   1 - 0x1
      11'h7A5: dout  = 8'b00000000; // 1957 :   0 - 0x0
      11'h7A6: dout  = 8'b00000000; // 1958 :   0 - 0x0
      11'h7A7: dout  = 8'b00000000; // 1959 :   0 - 0x0
      11'h7A8: dout  = 8'b00000011; // 1960 :   3 - 0x3 -- Sprite 0xf5
      11'h7A9: dout  = 8'b00001110; // 1961 :  14 - 0xe
      11'h7AA: dout  = 8'b11111000; // 1962 : 248 - 0xf8
      11'h7AB: dout  = 8'b00000000; // 1963 :   0 - 0x0
      11'h7AC: dout  = 8'b00000000; // 1964 :   0 - 0x0
      11'h7AD: dout  = 8'b00000000; // 1965 :   0 - 0x0
      11'h7AE: dout  = 8'b00000000; // 1966 :   0 - 0x0
      11'h7AF: dout  = 8'b00000000; // 1967 :   0 - 0x0
      11'h7B0: dout  = 8'b00100010; // 1968 :  34 - 0x22 -- Sprite 0xf6
      11'h7B1: dout  = 8'b01100101; // 1969 : 101 - 0x65
      11'h7B2: dout  = 8'b00100101; // 1970 :  37 - 0x25
      11'h7B3: dout  = 8'b00100101; // 1971 :  37 - 0x25
      11'h7B4: dout  = 8'b00100101; // 1972 :  37 - 0x25
      11'h7B5: dout  = 8'b00100101; // 1973 :  37 - 0x25
      11'h7B6: dout  = 8'b01110111; // 1974 : 119 - 0x77
      11'h7B7: dout  = 8'b01110010; // 1975 : 114 - 0x72
      11'h7B8: dout  = 8'b01100010; // 1976 :  98 - 0x62 -- Sprite 0xf7
      11'h7B9: dout  = 8'b10010101; // 1977 : 149 - 0x95
      11'h7BA: dout  = 8'b00010101; // 1978 :  21 - 0x15
      11'h7BB: dout  = 8'b00100101; // 1979 :  37 - 0x25
      11'h7BC: dout  = 8'b01000101; // 1980 :  69 - 0x45
      11'h7BD: dout  = 8'b10000101; // 1981 : 133 - 0x85
      11'h7BE: dout  = 8'b11110111; // 1982 : 247 - 0xf7
      11'h7BF: dout  = 8'b11110010; // 1983 : 242 - 0xf2
      11'h7C0: dout  = 8'b10100010; // 1984 : 162 - 0xa2 -- Sprite 0xf8
      11'h7C1: dout  = 8'b10100101; // 1985 : 165 - 0xa5
      11'h7C2: dout  = 8'b10100101; // 1986 : 165 - 0xa5
      11'h7C3: dout  = 8'b10100101; // 1987 : 165 - 0xa5
      11'h7C4: dout  = 8'b11110101; // 1988 : 245 - 0xf5
      11'h7C5: dout  = 8'b11110101; // 1989 : 245 - 0xf5
      11'h7C6: dout  = 8'b00100111; // 1990 :  39 - 0x27
      11'h7C7: dout  = 8'b00100010; // 1991 :  34 - 0x22
      11'h7C8: dout  = 8'b11110010; // 1992 : 242 - 0xf2 -- Sprite 0xf9
      11'h7C9: dout  = 8'b10000101; // 1993 : 133 - 0x85
      11'h7CA: dout  = 8'b10000101; // 1994 : 133 - 0x85
      11'h7CB: dout  = 8'b11100101; // 1995 : 229 - 0xe5
      11'h7CC: dout  = 8'b00010101; // 1996 :  21 - 0x15
      11'h7CD: dout  = 8'b00010101; // 1997 :  21 - 0x15
      11'h7CE: dout  = 8'b11110111; // 1998 : 247 - 0xf7
      11'h7CF: dout  = 8'b11100010; // 1999 : 226 - 0xe2
      11'h7D0: dout  = 8'b01100010; // 2000 :  98 - 0x62 -- Sprite 0xfa
      11'h7D1: dout  = 8'b10010101; // 2001 : 149 - 0x95
      11'h7D2: dout  = 8'b01010101; // 2002 :  85 - 0x55
      11'h7D3: dout  = 8'b01100101; // 2003 : 101 - 0x65
      11'h7D4: dout  = 8'b10110101; // 2004 : 181 - 0xb5
      11'h7D5: dout  = 8'b10010101; // 2005 : 149 - 0x95
      11'h7D6: dout  = 8'b10010111; // 2006 : 151 - 0x97
      11'h7D7: dout  = 8'b01100010; // 2007 :  98 - 0x62
      11'h7D8: dout  = 8'b00100000; // 2008 :  32 - 0x20 -- Sprite 0xfb
      11'h7D9: dout  = 8'b01010000; // 2009 :  80 - 0x50
      11'h7DA: dout  = 8'b01010000; // 2010 :  80 - 0x50
      11'h7DB: dout  = 8'b01010000; // 2011 :  80 - 0x50
      11'h7DC: dout  = 8'b01010000; // 2012 :  80 - 0x50
      11'h7DD: dout  = 8'b01010000; // 2013 :  80 - 0x50
      11'h7DE: dout  = 8'b01110000; // 2014 : 112 - 0x70
      11'h7DF: dout  = 8'b00100000; // 2015 :  32 - 0x20
      11'h7E0: dout  = 8'b00000000; // 2016 :   0 - 0x0 -- Sprite 0xfc
      11'h7E1: dout  = 8'b00000000; // 2017 :   0 - 0x0
      11'h7E2: dout  = 8'b00000000; // 2018 :   0 - 0x0
      11'h7E3: dout  = 8'b00000000; // 2019 :   0 - 0x0
      11'h7E4: dout  = 8'b00000000; // 2020 :   0 - 0x0
      11'h7E5: dout  = 8'b00000000; // 2021 :   0 - 0x0
      11'h7E6: dout  = 8'b00000000; // 2022 :   0 - 0x0
      11'h7E7: dout  = 8'b00000000; // 2023 :   0 - 0x0
      11'h7E8: dout  = 8'b01100110; // 2024 : 102 - 0x66 -- Sprite 0xfd
      11'h7E9: dout  = 8'b11100110; // 2025 : 230 - 0xe6
      11'h7EA: dout  = 8'b01100110; // 2026 : 102 - 0x66
      11'h7EB: dout  = 8'b01100110; // 2027 : 102 - 0x66
      11'h7EC: dout  = 8'b01100110; // 2028 : 102 - 0x66
      11'h7ED: dout  = 8'b01100111; // 2029 : 103 - 0x67
      11'h7EE: dout  = 8'b11110011; // 2030 : 243 - 0xf3
      11'h7EF: dout  = 8'b00000000; // 2031 :   0 - 0x0
      11'h7F0: dout  = 8'b01011110; // 2032 :  94 - 0x5e -- Sprite 0xfe
      11'h7F1: dout  = 8'b01011001; // 2033 :  89 - 0x59
      11'h7F2: dout  = 8'b01011001; // 2034 :  89 - 0x59
      11'h7F3: dout  = 8'b01011001; // 2035 :  89 - 0x59
      11'h7F4: dout  = 8'b01011110; // 2036 :  94 - 0x5e
      11'h7F5: dout  = 8'b11011000; // 2037 : 216 - 0xd8
      11'h7F6: dout  = 8'b10011000; // 2038 : 152 - 0x98
      11'h7F7: dout  = 8'b00000000; // 2039 :   0 - 0x0
      11'h7F8: dout  = 8'b00000000; // 2040 :   0 - 0x0 -- Sprite 0xff
      11'h7F9: dout  = 8'b00000000; // 2041 :   0 - 0x0
      11'h7FA: dout  = 8'b00000000; // 2042 :   0 - 0x0
      11'h7FB: dout  = 8'b00000000; // 2043 :   0 - 0x0
      11'h7FC: dout  = 8'b00000000; // 2044 :   0 - 0x0
      11'h7FD: dout  = 8'b00000100; // 2045 :   4 - 0x4
      11'h7FE: dout  = 8'b00001000; // 2046 :   8 - 0x8
      11'h7FF: dout  = 8'b00000000; // 2047 :   0 - 0x0
    endcase
  end

endmodule
