---   Background Pattern table COLOR PLANE 0
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
--- Autcmatically generated VHDL ROM from a NES memory file----


---  Original memory dump file name: pacman_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_PACMAN_BG_PLN0 is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(11-1 downto 0);  --2048 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_PACMAN_BG_PLN0;

architecture BEHAVIORAL of ROM_PTABLE_PACMAN_BG_PLN0 is
  signal addr_int  : natural range 0 to 2**11-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Background pattern Table COLOR PLANE 0
    "00000000", --    0 -  0x0  :    0 - 0x0 -- Background 0x0
    "00000000", --    1 -  0x1  :    0 - 0x0
    "00000000", --    2 -  0x2  :    0 - 0x0
    "00000000", --    3 -  0x3  :    0 - 0x0
    "00000000", --    4 -  0x4  :    0 - 0x0
    "00000000", --    5 -  0x5  :    0 - 0x0
    "00000000", --    6 -  0x6  :    0 - 0x0
    "00000000", --    7 -  0x7  :    0 - 0x0
    "00000000", --    8 -  0x8  :    0 - 0x0 -- Background 0x1
    "00111000", --    9 -  0x9  :   56 - 0x38
    "01111100", --   10 -  0xa  :  124 - 0x7c
    "11111110", --   11 -  0xb  :  254 - 0xfe
    "11111110", --   12 -  0xc  :  254 - 0xfe
    "11111110", --   13 -  0xd  :  254 - 0xfe
    "01111100", --   14 -  0xe  :  124 - 0x7c
    "00111000", --   15 -  0xf  :   56 - 0x38
    "00000000", --   16 - 0x10  :    0 - 0x0 -- Background 0x2
    "00000000", --   17 - 0x11  :    0 - 0x0
    "00000000", --   18 - 0x12  :    0 - 0x0
    "00000000", --   19 - 0x13  :    0 - 0x0
    "00000000", --   20 - 0x14  :    0 - 0x0
    "00000000", --   21 - 0x15  :    0 - 0x0
    "00000000", --   22 - 0x16  :    0 - 0x0
    "00000000", --   23 - 0x17  :    0 - 0x0
    "00000000", --   24 - 0x18  :    0 - 0x0 -- Background 0x3
    "00000000", --   25 - 0x19  :    0 - 0x0
    "00000000", --   26 - 0x1a  :    0 - 0x0
    "00011000", --   27 - 0x1b  :   24 - 0x18
    "00011000", --   28 - 0x1c  :   24 - 0x18
    "00000000", --   29 - 0x1d  :    0 - 0x0
    "00000000", --   30 - 0x1e  :    0 - 0x0
    "00000000", --   31 - 0x1f  :    0 - 0x0
    "00000000", --   32 - 0x20  :    0 - 0x0 -- Background 0x4
    "00000000", --   33 - 0x21  :    0 - 0x0
    "00000000", --   34 - 0x22  :    0 - 0x0
    "00000000", --   35 - 0x23  :    0 - 0x0
    "00000000", --   36 - 0x24  :    0 - 0x0
    "00000000", --   37 - 0x25  :    0 - 0x0
    "00000000", --   38 - 0x26  :    0 - 0x0
    "00000000", --   39 - 0x27  :    0 - 0x0
    "00000000", --   40 - 0x28  :    0 - 0x0 -- Background 0x5
    "00000000", --   41 - 0x29  :    0 - 0x0
    "00000000", --   42 - 0x2a  :    0 - 0x0
    "00000000", --   43 - 0x2b  :    0 - 0x0
    "00000000", --   44 - 0x2c  :    0 - 0x0
    "00000000", --   45 - 0x2d  :    0 - 0x0
    "00000000", --   46 - 0x2e  :    0 - 0x0
    "00000000", --   47 - 0x2f  :    0 - 0x0
    "00000000", --   48 - 0x30  :    0 - 0x0 -- Background 0x6
    "00000000", --   49 - 0x31  :    0 - 0x0
    "00000000", --   50 - 0x32  :    0 - 0x0
    "00000000", --   51 - 0x33  :    0 - 0x0
    "00000000", --   52 - 0x34  :    0 - 0x0
    "00000000", --   53 - 0x35  :    0 - 0x0
    "00000000", --   54 - 0x36  :    0 - 0x0
    "00000000", --   55 - 0x37  :    0 - 0x0
    "00000000", --   56 - 0x38  :    0 - 0x0 -- Background 0x7
    "00000000", --   57 - 0x39  :    0 - 0x0
    "00000000", --   58 - 0x3a  :    0 - 0x0
    "00000000", --   59 - 0x3b  :    0 - 0x0
    "00000000", --   60 - 0x3c  :    0 - 0x0
    "00000000", --   61 - 0x3d  :    0 - 0x0
    "00000000", --   62 - 0x3e  :    0 - 0x0
    "00000000", --   63 - 0x3f  :    0 - 0x0
    "00000000", --   64 - 0x40  :    0 - 0x0 -- Background 0x8
    "00000000", --   65 - 0x41  :    0 - 0x0
    "00000000", --   66 - 0x42  :    0 - 0x0
    "00000000", --   67 - 0x43  :    0 - 0x0
    "00000000", --   68 - 0x44  :    0 - 0x0
    "00000000", --   69 - 0x45  :    0 - 0x0
    "00000000", --   70 - 0x46  :    0 - 0x0
    "00000000", --   71 - 0x47  :    0 - 0x0
    "00000000", --   72 - 0x48  :    0 - 0x0 -- Background 0x9
    "00000000", --   73 - 0x49  :    0 - 0x0
    "00000000", --   74 - 0x4a  :    0 - 0x0
    "00011000", --   75 - 0x4b  :   24 - 0x18
    "00011000", --   76 - 0x4c  :   24 - 0x18
    "00000000", --   77 - 0x4d  :    0 - 0x0
    "00000000", --   78 - 0x4e  :    0 - 0x0
    "00000000", --   79 - 0x4f  :    0 - 0x0
    "00000000", --   80 - 0x50  :    0 - 0x0 -- Background 0xa
    "00000000", --   81 - 0x51  :    0 - 0x0
    "00000000", --   82 - 0x52  :    0 - 0x0
    "00000000", --   83 - 0x53  :    0 - 0x0
    "00000000", --   84 - 0x54  :    0 - 0x0
    "00000000", --   85 - 0x55  :    0 - 0x0
    "00000000", --   86 - 0x56  :    0 - 0x0
    "00000000", --   87 - 0x57  :    0 - 0x0
    "00000000", --   88 - 0x58  :    0 - 0x0 -- Background 0xb
    "00000000", --   89 - 0x59  :    0 - 0x0
    "00000000", --   90 - 0x5a  :    0 - 0x0
    "00000000", --   91 - 0x5b  :    0 - 0x0
    "00000000", --   92 - 0x5c  :    0 - 0x0
    "00000000", --   93 - 0x5d  :    0 - 0x0
    "00000000", --   94 - 0x5e  :    0 - 0x0
    "00000000", --   95 - 0x5f  :    0 - 0x0
    "00000000", --   96 - 0x60  :    0 - 0x0 -- Background 0xc
    "00000000", --   97 - 0x61  :    0 - 0x0
    "00000000", --   98 - 0x62  :    0 - 0x0
    "00000000", --   99 - 0x63  :    0 - 0x0
    "00000000", --  100 - 0x64  :    0 - 0x0
    "00000000", --  101 - 0x65  :    0 - 0x0
    "00000000", --  102 - 0x66  :    0 - 0x0
    "00000000", --  103 - 0x67  :    0 - 0x0
    "00000000", --  104 - 0x68  :    0 - 0x0 -- Background 0xd
    "00000000", --  105 - 0x69  :    0 - 0x0
    "00000000", --  106 - 0x6a  :    0 - 0x0
    "00000000", --  107 - 0x6b  :    0 - 0x0
    "00000000", --  108 - 0x6c  :    0 - 0x0
    "00000000", --  109 - 0x6d  :    0 - 0x0
    "00000000", --  110 - 0x6e  :    0 - 0x0
    "00000000", --  111 - 0x6f  :    0 - 0x0
    "00000000", --  112 - 0x70  :    0 - 0x0 -- Background 0xe
    "00000000", --  113 - 0x71  :    0 - 0x0
    "00000000", --  114 - 0x72  :    0 - 0x0
    "00000000", --  115 - 0x73  :    0 - 0x0
    "00000000", --  116 - 0x74  :    0 - 0x0
    "00000000", --  117 - 0x75  :    0 - 0x0
    "00000000", --  118 - 0x76  :    0 - 0x0
    "00000000", --  119 - 0x77  :    0 - 0x0
    "00000000", --  120 - 0x78  :    0 - 0x0 -- Background 0xf
    "00000000", --  121 - 0x79  :    0 - 0x0
    "00000000", --  122 - 0x7a  :    0 - 0x0
    "00000000", --  123 - 0x7b  :    0 - 0x0
    "00000000", --  124 - 0x7c  :    0 - 0x0
    "00000000", --  125 - 0x7d  :    0 - 0x0
    "00000000", --  126 - 0x7e  :    0 - 0x0
    "00000000", --  127 - 0x7f  :    0 - 0x0
    "00000000", --  128 - 0x80  :    0 - 0x0 -- Background 0x10
    "00000000", --  129 - 0x81  :    0 - 0x0
    "11111111", --  130 - 0x82  :  255 - 0xff
    "00000000", --  131 - 0x83  :    0 - 0x0
    "00000000", --  132 - 0x84  :    0 - 0x0
    "11111111", --  133 - 0x85  :  255 - 0xff
    "00000000", --  134 - 0x86  :    0 - 0x0
    "00000000", --  135 - 0x87  :    0 - 0x0
    "00100100", --  136 - 0x88  :   36 - 0x24 -- Background 0x11
    "00100100", --  137 - 0x89  :   36 - 0x24
    "00100100", --  138 - 0x8a  :   36 - 0x24
    "00100100", --  139 - 0x8b  :   36 - 0x24
    "00100100", --  140 - 0x8c  :   36 - 0x24
    "00100100", --  141 - 0x8d  :   36 - 0x24
    "00100100", --  142 - 0x8e  :   36 - 0x24
    "00100100", --  143 - 0x8f  :   36 - 0x24
    "00100100", --  144 - 0x90  :   36 - 0x24 -- Background 0x12
    "00100100", --  145 - 0x91  :   36 - 0x24
    "11000011", --  146 - 0x92  :  195 - 0xc3
    "00000000", --  147 - 0x93  :    0 - 0x0
    "00000000", --  148 - 0x94  :    0 - 0x0
    "11111111", --  149 - 0x95  :  255 - 0xff
    "00000000", --  150 - 0x96  :    0 - 0x0
    "00000000", --  151 - 0x97  :    0 - 0x0
    "00000000", --  152 - 0x98  :    0 - 0x0 -- Background 0x13
    "00000000", --  153 - 0x99  :    0 - 0x0
    "11111111", --  154 - 0x9a  :  255 - 0xff
    "00000000", --  155 - 0x9b  :    0 - 0x0
    "00000000", --  156 - 0x9c  :    0 - 0x0
    "11000011", --  157 - 0x9d  :  195 - 0xc3
    "00100100", --  158 - 0x9e  :   36 - 0x24
    "00100100", --  159 - 0x9f  :   36 - 0x24
    "00100100", --  160 - 0xa0  :   36 - 0x24 -- Background 0x14
    "00100100", --  161 - 0xa1  :   36 - 0x24
    "11000100", --  162 - 0xa2  :  196 - 0xc4
    "00000100", --  163 - 0xa3  :    4 - 0x4
    "00000100", --  164 - 0xa4  :    4 - 0x4
    "11000100", --  165 - 0xa5  :  196 - 0xc4
    "00100100", --  166 - 0xa6  :   36 - 0x24
    "00100100", --  167 - 0xa7  :   36 - 0x24
    "00100100", --  168 - 0xa8  :   36 - 0x24 -- Background 0x15
    "00100100", --  169 - 0xa9  :   36 - 0x24
    "00100011", --  170 - 0xaa  :   35 - 0x23
    "00100000", --  171 - 0xab  :   32 - 0x20
    "00100000", --  172 - 0xac  :   32 - 0x20
    "00100011", --  173 - 0xad  :   35 - 0x23
    "00100100", --  174 - 0xae  :   36 - 0x24
    "00100100", --  175 - 0xaf  :   36 - 0x24
    "00000000", --  176 - 0xb0  :    0 - 0x0 -- Background 0x16
    "00000000", --  177 - 0xb1  :    0 - 0x0
    "00001111", --  178 - 0xb2  :   15 - 0xf
    "00010000", --  179 - 0xb3  :   16 - 0x10
    "11110000", --  180 - 0xb4  :  240 - 0xf0
    "00001111", --  181 - 0xb5  :   15 - 0xf
    "00000000", --  182 - 0xb6  :    0 - 0x0
    "00000000", --  183 - 0xb7  :    0 - 0x0
    "00000000", --  184 - 0xb8  :    0 - 0x0 -- Background 0x17
    "00000000", --  185 - 0xb9  :    0 - 0x0
    "11110000", --  186 - 0xba  :  240 - 0xf0
    "00001000", --  187 - 0xbb  :    8 - 0x8
    "00001111", --  188 - 0xbc  :   15 - 0xf
    "11110000", --  189 - 0xbd  :  240 - 0xf0
    "00000000", --  190 - 0xbe  :    0 - 0x0
    "00000000", --  191 - 0xbf  :    0 - 0x0
    "00000000", --  192 - 0xc0  :    0 - 0x0 -- Background 0x18
    "00000000", --  193 - 0xc1  :    0 - 0x0
    "11110000", --  194 - 0xc2  :  240 - 0xf0
    "00001000", --  195 - 0xc3  :    8 - 0x8
    "00001000", --  196 - 0xc4  :    8 - 0x8
    "11110000", --  197 - 0xc5  :  240 - 0xf0
    "00000000", --  198 - 0xc6  :    0 - 0x0
    "00000000", --  199 - 0xc7  :    0 - 0x0
    "00000000", --  200 - 0xc8  :    0 - 0x0 -- Background 0x19
    "00000000", --  201 - 0xc9  :    0 - 0x0
    "00001111", --  202 - 0xca  :   15 - 0xf
    "00010000", --  203 - 0xcb  :   16 - 0x10
    "00010000", --  204 - 0xcc  :   16 - 0x10
    "00001111", --  205 - 0xcd  :   15 - 0xf
    "00000000", --  206 - 0xce  :    0 - 0x0
    "00000000", --  207 - 0xcf  :    0 - 0x0
    "00100100", --  208 - 0xd0  :   36 - 0x24 -- Background 0x1a
    "00100100", --  209 - 0xd1  :   36 - 0x24
    "00100100", --  210 - 0xd2  :   36 - 0x24
    "00100100", --  211 - 0xd3  :   36 - 0x24
    "00011000", --  212 - 0xd4  :   24 - 0x18
    "00000000", --  213 - 0xd5  :    0 - 0x0
    "00000000", --  214 - 0xd6  :    0 - 0x0
    "00000000", --  215 - 0xd7  :    0 - 0x0
    "00000000", --  216 - 0xd8  :    0 - 0x0 -- Background 0x1b
    "00000000", --  217 - 0xd9  :    0 - 0x0
    "00000000", --  218 - 0xda  :    0 - 0x0
    "00011000", --  219 - 0xdb  :   24 - 0x18
    "00100100", --  220 - 0xdc  :   36 - 0x24
    "00100100", --  221 - 0xdd  :   36 - 0x24
    "00100100", --  222 - 0xde  :   36 - 0x24
    "00100100", --  223 - 0xdf  :   36 - 0x24
    "00100100", --  224 - 0xe0  :   36 - 0x24 -- Background 0x1c
    "00100100", --  225 - 0xe1  :   36 - 0x24
    "11000100", --  226 - 0xe2  :  196 - 0xc4
    "00000100", --  227 - 0xe3  :    4 - 0x4
    "00001000", --  228 - 0xe4  :    8 - 0x8
    "11110000", --  229 - 0xe5  :  240 - 0xf0
    "00000000", --  230 - 0xe6  :    0 - 0x0
    "00000000", --  231 - 0xe7  :    0 - 0x0
    "00000000", --  232 - 0xe8  :    0 - 0x0 -- Background 0x1d
    "00000000", --  233 - 0xe9  :    0 - 0x0
    "11110000", --  234 - 0xea  :  240 - 0xf0
    "00001000", --  235 - 0xeb  :    8 - 0x8
    "00000100", --  236 - 0xec  :    4 - 0x4
    "11000100", --  237 - 0xed  :  196 - 0xc4
    "00100100", --  238 - 0xee  :   36 - 0x24
    "00100100", --  239 - 0xef  :   36 - 0x24
    "00100100", --  240 - 0xf0  :   36 - 0x24 -- Background 0x1e
    "00100100", --  241 - 0xf1  :   36 - 0x24
    "00100011", --  242 - 0xf2  :   35 - 0x23
    "00100000", --  243 - 0xf3  :   32 - 0x20
    "00010000", --  244 - 0xf4  :   16 - 0x10
    "00001111", --  245 - 0xf5  :   15 - 0xf
    "00000000", --  246 - 0xf6  :    0 - 0x0
    "00000000", --  247 - 0xf7  :    0 - 0x0
    "00000000", --  248 - 0xf8  :    0 - 0x0 -- Background 0x1f
    "00000000", --  249 - 0xf9  :    0 - 0x0
    "00001111", --  250 - 0xfa  :   15 - 0xf
    "00010000", --  251 - 0xfb  :   16 - 0x10
    "00100000", --  252 - 0xfc  :   32 - 0x20
    "00100011", --  253 - 0xfd  :   35 - 0x23
    "00100100", --  254 - 0xfe  :   36 - 0x24
    "00100100", --  255 - 0xff  :   36 - 0x24
    "00000000", --  256 - 0x100  :    0 - 0x0 -- Background 0x20
    "00000000", --  257 - 0x101  :    0 - 0x0
    "00000000", --  258 - 0x102  :    0 - 0x0
    "00000000", --  259 - 0x103  :    0 - 0x0
    "00000000", --  260 - 0x104  :    0 - 0x0
    "00000000", --  261 - 0x105  :    0 - 0x0
    "00000000", --  262 - 0x106  :    0 - 0x0
    "00000000", --  263 - 0x107  :    0 - 0x0
    "00000000", --  264 - 0x108  :    0 - 0x0 -- Background 0x21
    "00000000", --  265 - 0x109  :    0 - 0x0
    "11110000", --  266 - 0x10a  :  240 - 0xf0
    "00001000", --  267 - 0x10b  :    8 - 0x8
    "00001000", --  268 - 0x10c  :    8 - 0x8
    "11110000", --  269 - 0x10d  :  240 - 0xf0
    "00000000", --  270 - 0x10e  :    0 - 0x0
    "00000000", --  271 - 0x10f  :    0 - 0x0
    "00000000", --  272 - 0x110  :    0 - 0x0 -- Background 0x22
    "00000000", --  273 - 0x111  :    0 - 0x0
    "00001111", --  274 - 0x112  :   15 - 0xf
    "00010000", --  275 - 0x113  :   16 - 0x10
    "00010000", --  276 - 0x114  :   16 - 0x10
    "00001111", --  277 - 0x115  :   15 - 0xf
    "00000000", --  278 - 0x116  :    0 - 0x0
    "00000000", --  279 - 0x117  :    0 - 0x0
    "11111111", --  280 - 0x118  :  255 - 0xff -- Background 0x23
    "11111111", --  281 - 0x119  :  255 - 0xff
    "11100001", --  282 - 0x11a  :  225 - 0xe1
    "11100001", --  283 - 0x11b  :  225 - 0xe1
    "11100001", --  284 - 0x11c  :  225 - 0xe1
    "11100001", --  285 - 0x11d  :  225 - 0xe1
    "11100001", --  286 - 0x11e  :  225 - 0xe1
    "11100001", --  287 - 0x11f  :  225 - 0xe1
    "10000111", --  288 - 0x120  :  135 - 0x87 -- Background 0x24
    "11000111", --  289 - 0x121  :  199 - 0xc7
    "11000000", --  290 - 0x122  :  192 - 0xc0
    "11000111", --  291 - 0x123  :  199 - 0xc7
    "11001111", --  292 - 0x124  :  207 - 0xcf
    "11001110", --  293 - 0x125  :  206 - 0xce
    "11001111", --  294 - 0x126  :  207 - 0xcf
    "11000111", --  295 - 0x127  :  199 - 0xc7
    "11111000", --  296 - 0x128  :  248 - 0xf8 -- Background 0x25
    "11111100", --  297 - 0x129  :  252 - 0xfc
    "00011100", --  298 - 0x12a  :   28 - 0x1c
    "11111100", --  299 - 0x12b  :  252 - 0xfc
    "11111100", --  300 - 0x12c  :  252 - 0xfc
    "00011100", --  301 - 0x12d  :   28 - 0x1c
    "11111100", --  302 - 0x12e  :  252 - 0xfc
    "11111100", --  303 - 0x12f  :  252 - 0xfc
    "11111111", --  304 - 0x130  :  255 - 0xff -- Background 0x26
    "11111111", --  305 - 0x131  :  255 - 0xff
    "11100111", --  306 - 0x132  :  231 - 0xe7
    "11100111", --  307 - 0x133  :  231 - 0xe7
    "11100111", --  308 - 0x134  :  231 - 0xe7
    "11100111", --  309 - 0x135  :  231 - 0xe7
    "11100111", --  310 - 0x136  :  231 - 0xe7
    "11100111", --  311 - 0x137  :  231 - 0xe7
    "11110000", --  312 - 0x138  :  240 - 0xf0 -- Background 0x27
    "11111001", --  313 - 0x139  :  249 - 0xf9
    "00111001", --  314 - 0x13a  :   57 - 0x39
    "00111001", --  315 - 0x13b  :   57 - 0x39
    "00111001", --  316 - 0x13c  :   57 - 0x39
    "00111001", --  317 - 0x13d  :   57 - 0x39
    "00111001", --  318 - 0x13e  :   57 - 0x39
    "00111000", --  319 - 0x13f  :   56 - 0x38
    "11111111", --  320 - 0x140  :  255 - 0xff -- Background 0x28
    "11111111", --  321 - 0x141  :  255 - 0xff
    "11000000", --  322 - 0x142  :  192 - 0xc0
    "11000000", --  323 - 0x143  :  192 - 0xc0
    "11000000", --  324 - 0x144  :  192 - 0xc0
    "11000000", --  325 - 0x145  :  192 - 0xc0
    "11111111", --  326 - 0x146  :  255 - 0xff
    "11111111", --  327 - 0x147  :  255 - 0xff
    "00011111", --  328 - 0x148  :   31 - 0x1f -- Background 0x29
    "00111111", --  329 - 0x149  :   63 - 0x3f
    "00110000", --  330 - 0x14a  :   48 - 0x30
    "00110000", --  331 - 0x14b  :   48 - 0x30
    "00110000", --  332 - 0x14c  :   48 - 0x30
    "00110000", --  333 - 0x14d  :   48 - 0x30
    "00111111", --  334 - 0x14e  :   63 - 0x3f
    "00011111", --  335 - 0x14f  :   31 - 0x1f
    "11100011", --  336 - 0x150  :  227 - 0xe3 -- Background 0x2a
    "11110011", --  337 - 0x151  :  243 - 0xf3
    "01110000", --  338 - 0x152  :  112 - 0x70
    "01110000", --  339 - 0x153  :  112 - 0x70
    "01110000", --  340 - 0x154  :  112 - 0x70
    "01110000", --  341 - 0x155  :  112 - 0x70
    "11110000", --  342 - 0x156  :  240 - 0xf0
    "11100000", --  343 - 0x157  :  224 - 0xe0
    "11111110", --  344 - 0x158  :  254 - 0xfe -- Background 0x2b
    "11111110", --  345 - 0x159  :  254 - 0xfe
    "01110000", --  346 - 0x15a  :  112 - 0x70
    "01110000", --  347 - 0x15b  :  112 - 0x70
    "01110000", --  348 - 0x15c  :  112 - 0x70
    "01110000", --  349 - 0x15d  :  112 - 0x70
    "01110000", --  350 - 0x15e  :  112 - 0x70
    "01110000", --  351 - 0x15f  :  112 - 0x70
    "00000000", --  352 - 0x160  :    0 - 0x0 -- Background 0x2c
    "00000000", --  353 - 0x161  :    0 - 0x0
    "00000000", --  354 - 0x162  :    0 - 0x0
    "00000000", --  355 - 0x163  :    0 - 0x0
    "11111111", --  356 - 0x164  :  255 - 0xff
    "00000000", --  357 - 0x165  :    0 - 0x0
    "00000000", --  358 - 0x166  :    0 - 0x0
    "00000000", --  359 - 0x167  :    0 - 0x0
    "00000000", --  360 - 0x168  :    0 - 0x0 -- Background 0x2d
    "00000000", --  361 - 0x169  :    0 - 0x0
    "00000000", --  362 - 0x16a  :    0 - 0x0
    "00000000", --  363 - 0x16b  :    0 - 0x0
    "00000000", --  364 - 0x16c  :    0 - 0x0
    "00000000", --  365 - 0x16d  :    0 - 0x0
    "00000000", --  366 - 0x16e  :    0 - 0x0
    "00000000", --  367 - 0x16f  :    0 - 0x0
    "00000000", --  368 - 0x170  :    0 - 0x0 -- Background 0x2e
    "00000000", --  369 - 0x171  :    0 - 0x0
    "00000000", --  370 - 0x172  :    0 - 0x0
    "00011000", --  371 - 0x173  :   24 - 0x18
    "00011000", --  372 - 0x174  :   24 - 0x18
    "00000000", --  373 - 0x175  :    0 - 0x0
    "00000000", --  374 - 0x176  :    0 - 0x0
    "00000000", --  375 - 0x177  :    0 - 0x0
    "00000000", --  376 - 0x178  :    0 - 0x0 -- Background 0x2f
    "00000000", --  377 - 0x179  :    0 - 0x0
    "00000000", --  378 - 0x17a  :    0 - 0x0
    "00000000", --  379 - 0x17b  :    0 - 0x0
    "00000000", --  380 - 0x17c  :    0 - 0x0
    "00000000", --  381 - 0x17d  :    0 - 0x0
    "00000000", --  382 - 0x17e  :    0 - 0x0
    "00000000", --  383 - 0x17f  :    0 - 0x0
    "00011100", --  384 - 0x180  :   28 - 0x1c -- Background 0x30
    "00100110", --  385 - 0x181  :   38 - 0x26
    "01100011", --  386 - 0x182  :   99 - 0x63
    "01100011", --  387 - 0x183  :   99 - 0x63
    "01100011", --  388 - 0x184  :   99 - 0x63
    "00110010", --  389 - 0x185  :   50 - 0x32
    "00011100", --  390 - 0x186  :   28 - 0x1c
    "00000000", --  391 - 0x187  :    0 - 0x0
    "00001100", --  392 - 0x188  :   12 - 0xc -- Background 0x31
    "00011100", --  393 - 0x189  :   28 - 0x1c
    "00001100", --  394 - 0x18a  :   12 - 0xc
    "00001100", --  395 - 0x18b  :   12 - 0xc
    "00001100", --  396 - 0x18c  :   12 - 0xc
    "00001100", --  397 - 0x18d  :   12 - 0xc
    "00111111", --  398 - 0x18e  :   63 - 0x3f
    "00000000", --  399 - 0x18f  :    0 - 0x0
    "00111110", --  400 - 0x190  :   62 - 0x3e -- Background 0x32
    "01100011", --  401 - 0x191  :   99 - 0x63
    "00000111", --  402 - 0x192  :    7 - 0x7
    "00011110", --  403 - 0x193  :   30 - 0x1e
    "00111100", --  404 - 0x194  :   60 - 0x3c
    "01110000", --  405 - 0x195  :  112 - 0x70
    "01111111", --  406 - 0x196  :  127 - 0x7f
    "00000000", --  407 - 0x197  :    0 - 0x0
    "00111111", --  408 - 0x198  :   63 - 0x3f -- Background 0x33
    "00000110", --  409 - 0x199  :    6 - 0x6
    "00001100", --  410 - 0x19a  :   12 - 0xc
    "00011110", --  411 - 0x19b  :   30 - 0x1e
    "00000011", --  412 - 0x19c  :    3 - 0x3
    "01100011", --  413 - 0x19d  :   99 - 0x63
    "00111110", --  414 - 0x19e  :   62 - 0x3e
    "00000000", --  415 - 0x19f  :    0 - 0x0
    "00001110", --  416 - 0x1a0  :   14 - 0xe -- Background 0x34
    "00011110", --  417 - 0x1a1  :   30 - 0x1e
    "00110110", --  418 - 0x1a2  :   54 - 0x36
    "01100110", --  419 - 0x1a3  :  102 - 0x66
    "01111111", --  420 - 0x1a4  :  127 - 0x7f
    "00000110", --  421 - 0x1a5  :    6 - 0x6
    "00000110", --  422 - 0x1a6  :    6 - 0x6
    "00000000", --  423 - 0x1a7  :    0 - 0x0
    "01111110", --  424 - 0x1a8  :  126 - 0x7e -- Background 0x35
    "01100000", --  425 - 0x1a9  :   96 - 0x60
    "01111110", --  426 - 0x1aa  :  126 - 0x7e
    "00000011", --  427 - 0x1ab  :    3 - 0x3
    "00000011", --  428 - 0x1ac  :    3 - 0x3
    "01100011", --  429 - 0x1ad  :   99 - 0x63
    "00111110", --  430 - 0x1ae  :   62 - 0x3e
    "00000000", --  431 - 0x1af  :    0 - 0x0
    "00011110", --  432 - 0x1b0  :   30 - 0x1e -- Background 0x36
    "00110000", --  433 - 0x1b1  :   48 - 0x30
    "01100000", --  434 - 0x1b2  :   96 - 0x60
    "01111110", --  435 - 0x1b3  :  126 - 0x7e
    "01100011", --  436 - 0x1b4  :   99 - 0x63
    "01100011", --  437 - 0x1b5  :   99 - 0x63
    "00111110", --  438 - 0x1b6  :   62 - 0x3e
    "00000000", --  439 - 0x1b7  :    0 - 0x0
    "01111111", --  440 - 0x1b8  :  127 - 0x7f -- Background 0x37
    "01100011", --  441 - 0x1b9  :   99 - 0x63
    "00000110", --  442 - 0x1ba  :    6 - 0x6
    "00001100", --  443 - 0x1bb  :   12 - 0xc
    "00011000", --  444 - 0x1bc  :   24 - 0x18
    "00011000", --  445 - 0x1bd  :   24 - 0x18
    "00011000", --  446 - 0x1be  :   24 - 0x18
    "00000000", --  447 - 0x1bf  :    0 - 0x0
    "00111100", --  448 - 0x1c0  :   60 - 0x3c -- Background 0x38
    "01100010", --  449 - 0x1c1  :   98 - 0x62
    "01110010", --  450 - 0x1c2  :  114 - 0x72
    "00111100", --  451 - 0x1c3  :   60 - 0x3c
    "01001111", --  452 - 0x1c4  :   79 - 0x4f
    "01000011", --  453 - 0x1c5  :   67 - 0x43
    "00111110", --  454 - 0x1c6  :   62 - 0x3e
    "00000000", --  455 - 0x1c7  :    0 - 0x0
    "00111110", --  456 - 0x1c8  :   62 - 0x3e -- Background 0x39
    "01100011", --  457 - 0x1c9  :   99 - 0x63
    "01100011", --  458 - 0x1ca  :   99 - 0x63
    "00111111", --  459 - 0x1cb  :   63 - 0x3f
    "00000011", --  460 - 0x1cc  :    3 - 0x3
    "00000110", --  461 - 0x1cd  :    6 - 0x6
    "00111100", --  462 - 0x1ce  :   60 - 0x3c
    "00000000", --  463 - 0x1cf  :    0 - 0x0
    "00000000", --  464 - 0x1d0  :    0 - 0x0 -- Background 0x3a
    "00000000", --  465 - 0x1d1  :    0 - 0x0
    "00000000", --  466 - 0x1d2  :    0 - 0x0
    "01111110", --  467 - 0x1d3  :  126 - 0x7e
    "00000000", --  468 - 0x1d4  :    0 - 0x0
    "00000000", --  469 - 0x1d5  :    0 - 0x0
    "00000000", --  470 - 0x1d6  :    0 - 0x0
    "00000000", --  471 - 0x1d7  :    0 - 0x0
    "00000000", --  472 - 0x1d8  :    0 - 0x0 -- Background 0x3b
    "00000010", --  473 - 0x1d9  :    2 - 0x2
    "00000100", --  474 - 0x1da  :    4 - 0x4
    "00001000", --  475 - 0x1db  :    8 - 0x8
    "00010000", --  476 - 0x1dc  :   16 - 0x10
    "00100000", --  477 - 0x1dd  :   32 - 0x20
    "00000000", --  478 - 0x1de  :    0 - 0x0
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "00000000", --  480 - 0x1e0  :    0 - 0x0 -- Background 0x3c
    "00000111", --  481 - 0x1e1  :    7 - 0x7
    "00011111", --  482 - 0x1e2  :   31 - 0x1f
    "00111111", --  483 - 0x1e3  :   63 - 0x3f
    "00111111", --  484 - 0x1e4  :   63 - 0x3f
    "00001111", --  485 - 0x1e5  :   15 - 0xf
    "00000011", --  486 - 0x1e6  :    3 - 0x3
    "00000000", --  487 - 0x1e7  :    0 - 0x0
    "00000000", --  488 - 0x1e8  :    0 - 0x0 -- Background 0x3d
    "11000000", --  489 - 0x1e9  :  192 - 0xc0
    "11110000", --  490 - 0x1ea  :  240 - 0xf0
    "11111000", --  491 - 0x1eb  :  248 - 0xf8
    "11111000", --  492 - 0x1ec  :  248 - 0xf8
    "11111100", --  493 - 0x1ed  :  252 - 0xfc
    "11111100", --  494 - 0x1ee  :  252 - 0xfc
    "11111100", --  495 - 0x1ef  :  252 - 0xfc
    "00000000", --  496 - 0x1f0  :    0 - 0x0 -- Background 0x3e
    "00000011", --  497 - 0x1f1  :    3 - 0x3
    "00001111", --  498 - 0x1f2  :   15 - 0xf
    "00111111", --  499 - 0x1f3  :   63 - 0x3f
    "00111111", --  500 - 0x1f4  :   63 - 0x3f
    "00011111", --  501 - 0x1f5  :   31 - 0x1f
    "00000111", --  502 - 0x1f6  :    7 - 0x7
    "00000000", --  503 - 0x1f7  :    0 - 0x0
    "11111100", --  504 - 0x1f8  :  252 - 0xfc -- Background 0x3f
    "11111100", --  505 - 0x1f9  :  252 - 0xfc
    "11111100", --  506 - 0x1fa  :  252 - 0xfc
    "11111000", --  507 - 0x1fb  :  248 - 0xf8
    "11111000", --  508 - 0x1fc  :  248 - 0xf8
    "11110000", --  509 - 0x1fd  :  240 - 0xf0
    "11000000", --  510 - 0x1fe  :  192 - 0xc0
    "00000000", --  511 - 0x1ff  :    0 - 0x0
    "00000000", --  512 - 0x200  :    0 - 0x0 -- Background 0x40
    "00000000", --  513 - 0x201  :    0 - 0x0
    "00000000", --  514 - 0x202  :    0 - 0x0
    "00000000", --  515 - 0x203  :    0 - 0x0
    "00000000", --  516 - 0x204  :    0 - 0x0
    "00000000", --  517 - 0x205  :    0 - 0x0
    "00000000", --  518 - 0x206  :    0 - 0x0
    "00000000", --  519 - 0x207  :    0 - 0x0
    "00011100", --  520 - 0x208  :   28 - 0x1c -- Background 0x41
    "00110110", --  521 - 0x209  :   54 - 0x36
    "01100011", --  522 - 0x20a  :   99 - 0x63
    "01100011", --  523 - 0x20b  :   99 - 0x63
    "01111111", --  524 - 0x20c  :  127 - 0x7f
    "01100011", --  525 - 0x20d  :   99 - 0x63
    "01100011", --  526 - 0x20e  :   99 - 0x63
    "00000000", --  527 - 0x20f  :    0 - 0x0
    "01111110", --  528 - 0x210  :  126 - 0x7e -- Background 0x42
    "01100011", --  529 - 0x211  :   99 - 0x63
    "01100011", --  530 - 0x212  :   99 - 0x63
    "01111110", --  531 - 0x213  :  126 - 0x7e
    "01100011", --  532 - 0x214  :   99 - 0x63
    "01100011", --  533 - 0x215  :   99 - 0x63
    "01111110", --  534 - 0x216  :  126 - 0x7e
    "00000000", --  535 - 0x217  :    0 - 0x0
    "00011110", --  536 - 0x218  :   30 - 0x1e -- Background 0x43
    "00110011", --  537 - 0x219  :   51 - 0x33
    "01100000", --  538 - 0x21a  :   96 - 0x60
    "01100000", --  539 - 0x21b  :   96 - 0x60
    "01100000", --  540 - 0x21c  :   96 - 0x60
    "00110011", --  541 - 0x21d  :   51 - 0x33
    "00011110", --  542 - 0x21e  :   30 - 0x1e
    "00000000", --  543 - 0x21f  :    0 - 0x0
    "01111100", --  544 - 0x220  :  124 - 0x7c -- Background 0x44
    "01100110", --  545 - 0x221  :  102 - 0x66
    "01100011", --  546 - 0x222  :   99 - 0x63
    "01100011", --  547 - 0x223  :   99 - 0x63
    "01100011", --  548 - 0x224  :   99 - 0x63
    "01100110", --  549 - 0x225  :  102 - 0x66
    "01111100", --  550 - 0x226  :  124 - 0x7c
    "00000000", --  551 - 0x227  :    0 - 0x0
    "01111111", --  552 - 0x228  :  127 - 0x7f -- Background 0x45
    "01100000", --  553 - 0x229  :   96 - 0x60
    "01100000", --  554 - 0x22a  :   96 - 0x60
    "01111110", --  555 - 0x22b  :  126 - 0x7e
    "01100000", --  556 - 0x22c  :   96 - 0x60
    "01100000", --  557 - 0x22d  :   96 - 0x60
    "01111111", --  558 - 0x22e  :  127 - 0x7f
    "00000000", --  559 - 0x22f  :    0 - 0x0
    "01111111", --  560 - 0x230  :  127 - 0x7f -- Background 0x46
    "01100000", --  561 - 0x231  :   96 - 0x60
    "01100000", --  562 - 0x232  :   96 - 0x60
    "01111110", --  563 - 0x233  :  126 - 0x7e
    "01100000", --  564 - 0x234  :   96 - 0x60
    "01100000", --  565 - 0x235  :   96 - 0x60
    "01100000", --  566 - 0x236  :   96 - 0x60
    "00000000", --  567 - 0x237  :    0 - 0x0
    "00011111", --  568 - 0x238  :   31 - 0x1f -- Background 0x47
    "00110000", --  569 - 0x239  :   48 - 0x30
    "01100000", --  570 - 0x23a  :   96 - 0x60
    "01100111", --  571 - 0x23b  :  103 - 0x67
    "01100011", --  572 - 0x23c  :   99 - 0x63
    "00110011", --  573 - 0x23d  :   51 - 0x33
    "00011111", --  574 - 0x23e  :   31 - 0x1f
    "00000000", --  575 - 0x23f  :    0 - 0x0
    "01100011", --  576 - 0x240  :   99 - 0x63 -- Background 0x48
    "01100011", --  577 - 0x241  :   99 - 0x63
    "01100011", --  578 - 0x242  :   99 - 0x63
    "01111111", --  579 - 0x243  :  127 - 0x7f
    "01100011", --  580 - 0x244  :   99 - 0x63
    "01100011", --  581 - 0x245  :   99 - 0x63
    "01100011", --  582 - 0x246  :   99 - 0x63
    "00000000", --  583 - 0x247  :    0 - 0x0
    "00111111", --  584 - 0x248  :   63 - 0x3f -- Background 0x49
    "00001100", --  585 - 0x249  :   12 - 0xc
    "00001100", --  586 - 0x24a  :   12 - 0xc
    "00001100", --  587 - 0x24b  :   12 - 0xc
    "00001100", --  588 - 0x24c  :   12 - 0xc
    "00001100", --  589 - 0x24d  :   12 - 0xc
    "00111111", --  590 - 0x24e  :   63 - 0x3f
    "00000000", --  591 - 0x24f  :    0 - 0x0
    "00000011", --  592 - 0x250  :    3 - 0x3 -- Background 0x4a
    "00000011", --  593 - 0x251  :    3 - 0x3
    "00000011", --  594 - 0x252  :    3 - 0x3
    "00000011", --  595 - 0x253  :    3 - 0x3
    "00000011", --  596 - 0x254  :    3 - 0x3
    "01100011", --  597 - 0x255  :   99 - 0x63
    "00111110", --  598 - 0x256  :   62 - 0x3e
    "00000000", --  599 - 0x257  :    0 - 0x0
    "01100011", --  600 - 0x258  :   99 - 0x63 -- Background 0x4b
    "01100110", --  601 - 0x259  :  102 - 0x66
    "01101100", --  602 - 0x25a  :  108 - 0x6c
    "01111000", --  603 - 0x25b  :  120 - 0x78
    "01111100", --  604 - 0x25c  :  124 - 0x7c
    "01100110", --  605 - 0x25d  :  102 - 0x66
    "01100011", --  606 - 0x25e  :   99 - 0x63
    "00000000", --  607 - 0x25f  :    0 - 0x0
    "01100000", --  608 - 0x260  :   96 - 0x60 -- Background 0x4c
    "01100000", --  609 - 0x261  :   96 - 0x60
    "01100000", --  610 - 0x262  :   96 - 0x60
    "01100000", --  611 - 0x263  :   96 - 0x60
    "01100000", --  612 - 0x264  :   96 - 0x60
    "01100000", --  613 - 0x265  :   96 - 0x60
    "01111111", --  614 - 0x266  :  127 - 0x7f
    "00000000", --  615 - 0x267  :    0 - 0x0
    "01100011", --  616 - 0x268  :   99 - 0x63 -- Background 0x4d
    "01110111", --  617 - 0x269  :  119 - 0x77
    "01111111", --  618 - 0x26a  :  127 - 0x7f
    "01111111", --  619 - 0x26b  :  127 - 0x7f
    "01101011", --  620 - 0x26c  :  107 - 0x6b
    "01100011", --  621 - 0x26d  :   99 - 0x63
    "01100011", --  622 - 0x26e  :   99 - 0x63
    "00000000", --  623 - 0x26f  :    0 - 0x0
    "01100011", --  624 - 0x270  :   99 - 0x63 -- Background 0x4e
    "01110011", --  625 - 0x271  :  115 - 0x73
    "01111011", --  626 - 0x272  :  123 - 0x7b
    "01111111", --  627 - 0x273  :  127 - 0x7f
    "01101111", --  628 - 0x274  :  111 - 0x6f
    "01100111", --  629 - 0x275  :  103 - 0x67
    "01100011", --  630 - 0x276  :   99 - 0x63
    "00000000", --  631 - 0x277  :    0 - 0x0
    "00111110", --  632 - 0x278  :   62 - 0x3e -- Background 0x4f
    "01100011", --  633 - 0x279  :   99 - 0x63
    "01100011", --  634 - 0x27a  :   99 - 0x63
    "01100011", --  635 - 0x27b  :   99 - 0x63
    "01100011", --  636 - 0x27c  :   99 - 0x63
    "01100011", --  637 - 0x27d  :   99 - 0x63
    "00111110", --  638 - 0x27e  :   62 - 0x3e
    "00000000", --  639 - 0x27f  :    0 - 0x0
    "01111110", --  640 - 0x280  :  126 - 0x7e -- Background 0x50
    "01100011", --  641 - 0x281  :   99 - 0x63
    "01100011", --  642 - 0x282  :   99 - 0x63
    "01100011", --  643 - 0x283  :   99 - 0x63
    "01111110", --  644 - 0x284  :  126 - 0x7e
    "01100000", --  645 - 0x285  :   96 - 0x60
    "01100000", --  646 - 0x286  :   96 - 0x60
    "00000000", --  647 - 0x287  :    0 - 0x0
    "00111110", --  648 - 0x288  :   62 - 0x3e -- Background 0x51
    "01100011", --  649 - 0x289  :   99 - 0x63
    "01100011", --  650 - 0x28a  :   99 - 0x63
    "01100011", --  651 - 0x28b  :   99 - 0x63
    "01101111", --  652 - 0x28c  :  111 - 0x6f
    "01100110", --  653 - 0x28d  :  102 - 0x66
    "00111101", --  654 - 0x28e  :   61 - 0x3d
    "00000000", --  655 - 0x28f  :    0 - 0x0
    "01111110", --  656 - 0x290  :  126 - 0x7e -- Background 0x52
    "01100011", --  657 - 0x291  :   99 - 0x63
    "01100011", --  658 - 0x292  :   99 - 0x63
    "01100111", --  659 - 0x293  :  103 - 0x67
    "01111100", --  660 - 0x294  :  124 - 0x7c
    "01101110", --  661 - 0x295  :  110 - 0x6e
    "01100111", --  662 - 0x296  :  103 - 0x67
    "00000000", --  663 - 0x297  :    0 - 0x0
    "00111100", --  664 - 0x298  :   60 - 0x3c -- Background 0x53
    "01100110", --  665 - 0x299  :  102 - 0x66
    "01100000", --  666 - 0x29a  :   96 - 0x60
    "00111110", --  667 - 0x29b  :   62 - 0x3e
    "00000011", --  668 - 0x29c  :    3 - 0x3
    "01100011", --  669 - 0x29d  :   99 - 0x63
    "00111110", --  670 - 0x29e  :   62 - 0x3e
    "00000000", --  671 - 0x29f  :    0 - 0x0
    "00111111", --  672 - 0x2a0  :   63 - 0x3f -- Background 0x54
    "00001100", --  673 - 0x2a1  :   12 - 0xc
    "00001100", --  674 - 0x2a2  :   12 - 0xc
    "00001100", --  675 - 0x2a3  :   12 - 0xc
    "00001100", --  676 - 0x2a4  :   12 - 0xc
    "00001100", --  677 - 0x2a5  :   12 - 0xc
    "00001100", --  678 - 0x2a6  :   12 - 0xc
    "00000000", --  679 - 0x2a7  :    0 - 0x0
    "01100011", --  680 - 0x2a8  :   99 - 0x63 -- Background 0x55
    "01100011", --  681 - 0x2a9  :   99 - 0x63
    "01100011", --  682 - 0x2aa  :   99 - 0x63
    "01100011", --  683 - 0x2ab  :   99 - 0x63
    "01100011", --  684 - 0x2ac  :   99 - 0x63
    "01100011", --  685 - 0x2ad  :   99 - 0x63
    "00111110", --  686 - 0x2ae  :   62 - 0x3e
    "00000000", --  687 - 0x2af  :    0 - 0x0
    "01100011", --  688 - 0x2b0  :   99 - 0x63 -- Background 0x56
    "01100011", --  689 - 0x2b1  :   99 - 0x63
    "01100011", --  690 - 0x2b2  :   99 - 0x63
    "01110111", --  691 - 0x2b3  :  119 - 0x77
    "00111110", --  692 - 0x2b4  :   62 - 0x3e
    "00011100", --  693 - 0x2b5  :   28 - 0x1c
    "00001000", --  694 - 0x2b6  :    8 - 0x8
    "00000000", --  695 - 0x2b7  :    0 - 0x0
    "01100011", --  696 - 0x2b8  :   99 - 0x63 -- Background 0x57
    "01100011", --  697 - 0x2b9  :   99 - 0x63
    "01101011", --  698 - 0x2ba  :  107 - 0x6b
    "01111111", --  699 - 0x2bb  :  127 - 0x7f
    "01111111", --  700 - 0x2bc  :  127 - 0x7f
    "01110111", --  701 - 0x2bd  :  119 - 0x77
    "01100011", --  702 - 0x2be  :   99 - 0x63
    "00000000", --  703 - 0x2bf  :    0 - 0x0
    "01100011", --  704 - 0x2c0  :   99 - 0x63 -- Background 0x58
    "01110111", --  705 - 0x2c1  :  119 - 0x77
    "00111110", --  706 - 0x2c2  :   62 - 0x3e
    "00011100", --  707 - 0x2c3  :   28 - 0x1c
    "00111110", --  708 - 0x2c4  :   62 - 0x3e
    "01110111", --  709 - 0x2c5  :  119 - 0x77
    "01100011", --  710 - 0x2c6  :   99 - 0x63
    "00000000", --  711 - 0x2c7  :    0 - 0x0
    "00110011", --  712 - 0x2c8  :   51 - 0x33 -- Background 0x59
    "00110011", --  713 - 0x2c9  :   51 - 0x33
    "00110011", --  714 - 0x2ca  :   51 - 0x33
    "00011110", --  715 - 0x2cb  :   30 - 0x1e
    "00001100", --  716 - 0x2cc  :   12 - 0xc
    "00001100", --  717 - 0x2cd  :   12 - 0xc
    "00001100", --  718 - 0x2ce  :   12 - 0xc
    "00000000", --  719 - 0x2cf  :    0 - 0x0
    "01111111", --  720 - 0x2d0  :  127 - 0x7f -- Background 0x5a
    "00000111", --  721 - 0x2d1  :    7 - 0x7
    "00001110", --  722 - 0x2d2  :   14 - 0xe
    "00011100", --  723 - 0x2d3  :   28 - 0x1c
    "00111000", --  724 - 0x2d4  :   56 - 0x38
    "01110000", --  725 - 0x2d5  :  112 - 0x70
    "01111111", --  726 - 0x2d6  :  127 - 0x7f
    "00000000", --  727 - 0x2d7  :    0 - 0x0
    "00000000", --  728 - 0x2d8  :    0 - 0x0 -- Background 0x5b
    "00000000", --  729 - 0x2d9  :    0 - 0x0
    "00000000", --  730 - 0x2da  :    0 - 0x0
    "00000000", --  731 - 0x2db  :    0 - 0x0
    "00000000", --  732 - 0x2dc  :    0 - 0x0
    "00110000", --  733 - 0x2dd  :   48 - 0x30
    "00110000", --  734 - 0x2de  :   48 - 0x30
    "00000000", --  735 - 0x2df  :    0 - 0x0
    "11000000", --  736 - 0x2e0  :  192 - 0xc0 -- Background 0x5c
    "11110000", --  737 - 0x2e1  :  240 - 0xf0
    "11111100", --  738 - 0x2e2  :  252 - 0xfc
    "11111111", --  739 - 0x2e3  :  255 - 0xff
    "11111100", --  740 - 0x2e4  :  252 - 0xfc
    "11110000", --  741 - 0x2e5  :  240 - 0xf0
    "11000000", --  742 - 0x2e6  :  192 - 0xc0
    "00000000", --  743 - 0x2e7  :    0 - 0x0
    "00111100", --  744 - 0x2e8  :   60 - 0x3c -- Background 0x5d
    "01000010", --  745 - 0x2e9  :   66 - 0x42
    "10011001", --  746 - 0x2ea  :  153 - 0x99
    "10100001", --  747 - 0x2eb  :  161 - 0xa1
    "10100001", --  748 - 0x2ec  :  161 - 0xa1
    "10011001", --  749 - 0x2ed  :  153 - 0x99
    "01000010", --  750 - 0x2ee  :   66 - 0x42
    "00111100", --  751 - 0x2ef  :   60 - 0x3c
    "00000000", --  752 - 0x2f0  :    0 - 0x0 -- Background 0x5e
    "00000000", --  753 - 0x2f1  :    0 - 0x0
    "00010000", --  754 - 0x2f2  :   16 - 0x10
    "00010000", --  755 - 0x2f3  :   16 - 0x10
    "00010000", --  756 - 0x2f4  :   16 - 0x10
    "00010000", --  757 - 0x2f5  :   16 - 0x10
    "00000000", --  758 - 0x2f6  :    0 - 0x0
    "00000000", --  759 - 0x2f7  :    0 - 0x0
    "00110110", --  760 - 0x2f8  :   54 - 0x36 -- Background 0x5f
    "00110110", --  761 - 0x2f9  :   54 - 0x36
    "00010010", --  762 - 0x2fa  :   18 - 0x12
    "00000000", --  763 - 0x2fb  :    0 - 0x0
    "00000000", --  764 - 0x2fc  :    0 - 0x0
    "00000000", --  765 - 0x2fd  :    0 - 0x0
    "00000000", --  766 - 0x2fe  :    0 - 0x0
    "00000000", --  767 - 0x2ff  :    0 - 0x0
    "00000000", --  768 - 0x300  :    0 - 0x0 -- Background 0x60
    "00000000", --  769 - 0x301  :    0 - 0x0
    "00000000", --  770 - 0x302  :    0 - 0x0
    "00000000", --  771 - 0x303  :    0 - 0x0
    "00000000", --  772 - 0x304  :    0 - 0x0
    "00000001", --  773 - 0x305  :    1 - 0x1
    "00011110", --  774 - 0x306  :   30 - 0x1e
    "00111011", --  775 - 0x307  :   59 - 0x3b
    "00000000", --  776 - 0x308  :    0 - 0x0 -- Background 0x61
    "00000000", --  777 - 0x309  :    0 - 0x0
    "00001100", --  778 - 0x30a  :   12 - 0xc
    "00111100", --  779 - 0x30b  :   60 - 0x3c
    "11010000", --  780 - 0x30c  :  208 - 0xd0
    "00010000", --  781 - 0x30d  :   16 - 0x10
    "00100000", --  782 - 0x30e  :   32 - 0x20
    "01000000", --  783 - 0x30f  :   64 - 0x40
    "00111110", --  784 - 0x310  :   62 - 0x3e -- Background 0x62
    "00101101", --  785 - 0x311  :   45 - 0x2d
    "00110101", --  786 - 0x312  :   53 - 0x35
    "00011101", --  787 - 0x313  :   29 - 0x1d
    "00000001", --  788 - 0x314  :    1 - 0x1
    "00000000", --  789 - 0x315  :    0 - 0x0
    "00000000", --  790 - 0x316  :    0 - 0x0
    "00000000", --  791 - 0x317  :    0 - 0x0
    "10110000", --  792 - 0x318  :  176 - 0xb0 -- Background 0x63
    "10111000", --  793 - 0x319  :  184 - 0xb8
    "11111000", --  794 - 0x31a  :  248 - 0xf8
    "01111000", --  795 - 0x31b  :  120 - 0x78
    "10011000", --  796 - 0x31c  :  152 - 0x98
    "11110000", --  797 - 0x31d  :  240 - 0xf0
    "00000000", --  798 - 0x31e  :    0 - 0x0
    "00000000", --  799 - 0x31f  :    0 - 0x0
    "00000000", --  800 - 0x320  :    0 - 0x0 -- Background 0x64
    "00000000", --  801 - 0x321  :    0 - 0x0
    "00000111", --  802 - 0x322  :    7 - 0x7
    "00000011", --  803 - 0x323  :    3 - 0x3
    "00001101", --  804 - 0x324  :   13 - 0xd
    "00011110", --  805 - 0x325  :   30 - 0x1e
    "00010111", --  806 - 0x326  :   23 - 0x17
    "00011101", --  807 - 0x327  :   29 - 0x1d
    "00000000", --  808 - 0x328  :    0 - 0x0 -- Background 0x65
    "10000000", --  809 - 0x329  :  128 - 0x80
    "01110000", --  810 - 0x32a  :  112 - 0x70
    "11100000", --  811 - 0x32b  :  224 - 0xe0
    "11011000", --  812 - 0x32c  :  216 - 0xd8
    "10111100", --  813 - 0x32d  :  188 - 0xbc
    "01110100", --  814 - 0x32e  :  116 - 0x74
    "11011100", --  815 - 0x32f  :  220 - 0xdc
    "00011111", --  816 - 0x330  :   31 - 0x1f -- Background 0x66
    "00001011", --  817 - 0x331  :   11 - 0xb
    "00001111", --  818 - 0x332  :   15 - 0xf
    "00000101", --  819 - 0x333  :    5 - 0x5
    "00000011", --  820 - 0x334  :    3 - 0x3
    "00000001", --  821 - 0x335  :    1 - 0x1
    "00000000", --  822 - 0x336  :    0 - 0x0
    "00000000", --  823 - 0x337  :    0 - 0x0
    "11111100", --  824 - 0x338  :  252 - 0xfc -- Background 0x67
    "01101000", --  825 - 0x339  :  104 - 0x68
    "11111000", --  826 - 0x33a  :  248 - 0xf8
    "10110000", --  827 - 0x33b  :  176 - 0xb0
    "11100000", --  828 - 0x33c  :  224 - 0xe0
    "10000000", --  829 - 0x33d  :  128 - 0x80
    "00000000", --  830 - 0x33e  :    0 - 0x0
    "00000000", --  831 - 0x33f  :    0 - 0x0
    "00000000", --  832 - 0x340  :    0 - 0x0 -- Background 0x68
    "00000000", --  833 - 0x341  :    0 - 0x0
    "00000000", --  834 - 0x342  :    0 - 0x0
    "00000000", --  835 - 0x343  :    0 - 0x0
    "00000000", --  836 - 0x344  :    0 - 0x0
    "00000000", --  837 - 0x345  :    0 - 0x0
    "00000000", --  838 - 0x346  :    0 - 0x0
    "00000000", --  839 - 0x347  :    0 - 0x0
    "00000000", --  840 - 0x348  :    0 - 0x0 -- Background 0x69
    "00000000", --  841 - 0x349  :    0 - 0x0
    "00000000", --  842 - 0x34a  :    0 - 0x0
    "00000000", --  843 - 0x34b  :    0 - 0x0
    "00000000", --  844 - 0x34c  :    0 - 0x0
    "00000000", --  845 - 0x34d  :    0 - 0x0
    "00000000", --  846 - 0x34e  :    0 - 0x0
    "00000000", --  847 - 0x34f  :    0 - 0x0
    "00000000", --  848 - 0x350  :    0 - 0x0 -- Background 0x6a
    "00000000", --  849 - 0x351  :    0 - 0x0
    "00000000", --  850 - 0x352  :    0 - 0x0
    "00000000", --  851 - 0x353  :    0 - 0x0
    "00000000", --  852 - 0x354  :    0 - 0x0
    "00000000", --  853 - 0x355  :    0 - 0x0
    "00000000", --  854 - 0x356  :    0 - 0x0
    "00000000", --  855 - 0x357  :    0 - 0x0
    "00000000", --  856 - 0x358  :    0 - 0x0 -- Background 0x6b
    "00000000", --  857 - 0x359  :    0 - 0x0
    "00000000", --  858 - 0x35a  :    0 - 0x0
    "00000000", --  859 - 0x35b  :    0 - 0x0
    "00000000", --  860 - 0x35c  :    0 - 0x0
    "00000000", --  861 - 0x35d  :    0 - 0x0
    "00000000", --  862 - 0x35e  :    0 - 0x0
    "00000000", --  863 - 0x35f  :    0 - 0x0
    "00000000", --  864 - 0x360  :    0 - 0x0 -- Background 0x6c
    "00000000", --  865 - 0x361  :    0 - 0x0
    "00000001", --  866 - 0x362  :    1 - 0x1
    "00011101", --  867 - 0x363  :   29 - 0x1d
    "00111110", --  868 - 0x364  :   62 - 0x3e
    "00111111", --  869 - 0x365  :   63 - 0x3f
    "00111111", --  870 - 0x366  :   63 - 0x3f
    "00111111", --  871 - 0x367  :   63 - 0x3f
    "00000000", --  872 - 0x368  :    0 - 0x0 -- Background 0x6d
    "10000000", --  873 - 0x369  :  128 - 0x80
    "00000000", --  874 - 0x36a  :    0 - 0x0
    "01110000", --  875 - 0x36b  :  112 - 0x70
    "11111000", --  876 - 0x36c  :  248 - 0xf8
    "11111100", --  877 - 0x36d  :  252 - 0xfc
    "11111100", --  878 - 0x36e  :  252 - 0xfc
    "11111100", --  879 - 0x36f  :  252 - 0xfc
    "00111111", --  880 - 0x370  :   63 - 0x3f -- Background 0x6e
    "00111111", --  881 - 0x371  :   63 - 0x3f
    "00011111", --  882 - 0x372  :   31 - 0x1f
    "00011111", --  883 - 0x373  :   31 - 0x1f
    "00001111", --  884 - 0x374  :   15 - 0xf
    "00000110", --  885 - 0x375  :    6 - 0x6
    "00000000", --  886 - 0x376  :    0 - 0x0
    "00000000", --  887 - 0x377  :    0 - 0x0
    "11101100", --  888 - 0x378  :  236 - 0xec -- Background 0x6f
    "11101100", --  889 - 0x379  :  236 - 0xec
    "11011000", --  890 - 0x37a  :  216 - 0xd8
    "11111000", --  891 - 0x37b  :  248 - 0xf8
    "11110000", --  892 - 0x37c  :  240 - 0xf0
    "11100000", --  893 - 0x37d  :  224 - 0xe0
    "00000000", --  894 - 0x37e  :    0 - 0x0
    "00000000", --  895 - 0x37f  :    0 - 0x0
    "00000000", --  896 - 0x380  :    0 - 0x0 -- Background 0x70
    "00000100", --  897 - 0x381  :    4 - 0x4
    "00000011", --  898 - 0x382  :    3 - 0x3
    "00000000", --  899 - 0x383  :    0 - 0x0
    "00000001", --  900 - 0x384  :    1 - 0x1
    "00000111", --  901 - 0x385  :    7 - 0x7
    "00001111", --  902 - 0x386  :   15 - 0xf
    "00001100", --  903 - 0x387  :   12 - 0xc
    "00000000", --  904 - 0x388  :    0 - 0x0 -- Background 0x71
    "00000000", --  905 - 0x389  :    0 - 0x0
    "11100000", --  906 - 0x38a  :  224 - 0xe0
    "10000000", --  907 - 0x38b  :  128 - 0x80
    "01000000", --  908 - 0x38c  :   64 - 0x40
    "11110000", --  909 - 0x38d  :  240 - 0xf0
    "10011000", --  910 - 0x38e  :  152 - 0x98
    "11111000", --  911 - 0x38f  :  248 - 0xf8
    "00011111", --  912 - 0x390  :   31 - 0x1f -- Background 0x72
    "00010011", --  913 - 0x391  :   19 - 0x13
    "00011111", --  914 - 0x392  :   31 - 0x1f
    "00001111", --  915 - 0x393  :   15 - 0xf
    "00001001", --  916 - 0x394  :    9 - 0x9
    "00000111", --  917 - 0x395  :    7 - 0x7
    "00000001", --  918 - 0x396  :    1 - 0x1
    "00000000", --  919 - 0x397  :    0 - 0x0
    "11100100", --  920 - 0x398  :  228 - 0xe4 -- Background 0x73
    "00111100", --  921 - 0x399  :   60 - 0x3c
    "11100100", --  922 - 0x39a  :  228 - 0xe4
    "00111000", --  923 - 0x39b  :   56 - 0x38
    "11111000", --  924 - 0x39c  :  248 - 0xf8
    "11110000", --  925 - 0x39d  :  240 - 0xf0
    "11000000", --  926 - 0x39e  :  192 - 0xc0
    "00000000", --  927 - 0x39f  :    0 - 0x0
    "00000000", --  928 - 0x3a0  :    0 - 0x0 -- Background 0x74
    "00000000", --  929 - 0x3a1  :    0 - 0x0
    "00000000", --  930 - 0x3a2  :    0 - 0x0
    "00000000", --  931 - 0x3a3  :    0 - 0x0
    "00000000", --  932 - 0x3a4  :    0 - 0x0
    "00000000", --  933 - 0x3a5  :    0 - 0x0
    "00000000", --  934 - 0x3a6  :    0 - 0x0
    "00000000", --  935 - 0x3a7  :    0 - 0x0
    "00000000", --  936 - 0x3a8  :    0 - 0x0 -- Background 0x75
    "00000000", --  937 - 0x3a9  :    0 - 0x0
    "00000000", --  938 - 0x3aa  :    0 - 0x0
    "00000000", --  939 - 0x3ab  :    0 - 0x0
    "00000000", --  940 - 0x3ac  :    0 - 0x0
    "00000000", --  941 - 0x3ad  :    0 - 0x0
    "00000000", --  942 - 0x3ae  :    0 - 0x0
    "00000000", --  943 - 0x3af  :    0 - 0x0
    "00000000", --  944 - 0x3b0  :    0 - 0x0 -- Background 0x76
    "00000000", --  945 - 0x3b1  :    0 - 0x0
    "00000000", --  946 - 0x3b2  :    0 - 0x0
    "00000000", --  947 - 0x3b3  :    0 - 0x0
    "00000000", --  948 - 0x3b4  :    0 - 0x0
    "00000000", --  949 - 0x3b5  :    0 - 0x0
    "00000000", --  950 - 0x3b6  :    0 - 0x0
    "00000000", --  951 - 0x3b7  :    0 - 0x0
    "00000000", --  952 - 0x3b8  :    0 - 0x0 -- Background 0x77
    "00000000", --  953 - 0x3b9  :    0 - 0x0
    "00000000", --  954 - 0x3ba  :    0 - 0x0
    "00000000", --  955 - 0x3bb  :    0 - 0x0
    "00000000", --  956 - 0x3bc  :    0 - 0x0
    "00000000", --  957 - 0x3bd  :    0 - 0x0
    "00000000", --  958 - 0x3be  :    0 - 0x0
    "00000000", --  959 - 0x3bf  :    0 - 0x0
    "00000000", --  960 - 0x3c0  :    0 - 0x0 -- Background 0x78
    "00000000", --  961 - 0x3c1  :    0 - 0x0
    "00000000", --  962 - 0x3c2  :    0 - 0x0
    "00000000", --  963 - 0x3c3  :    0 - 0x0
    "00000000", --  964 - 0x3c4  :    0 - 0x0
    "00000000", --  965 - 0x3c5  :    0 - 0x0
    "00000000", --  966 - 0x3c6  :    0 - 0x0
    "00000000", --  967 - 0x3c7  :    0 - 0x0
    "00000000", --  968 - 0x3c8  :    0 - 0x0 -- Background 0x79
    "00000000", --  969 - 0x3c9  :    0 - 0x0
    "00000000", --  970 - 0x3ca  :    0 - 0x0
    "00000000", --  971 - 0x3cb  :    0 - 0x0
    "00000000", --  972 - 0x3cc  :    0 - 0x0
    "00000000", --  973 - 0x3cd  :    0 - 0x0
    "00000000", --  974 - 0x3ce  :    0 - 0x0
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "00000000", --  976 - 0x3d0  :    0 - 0x0 -- Background 0x7a
    "00000000", --  977 - 0x3d1  :    0 - 0x0
    "00000000", --  978 - 0x3d2  :    0 - 0x0
    "00000000", --  979 - 0x3d3  :    0 - 0x0
    "00000000", --  980 - 0x3d4  :    0 - 0x0
    "00000000", --  981 - 0x3d5  :    0 - 0x0
    "00000000", --  982 - 0x3d6  :    0 - 0x0
    "00000000", --  983 - 0x3d7  :    0 - 0x0
    "00000000", --  984 - 0x3d8  :    0 - 0x0 -- Background 0x7b
    "00000000", --  985 - 0x3d9  :    0 - 0x0
    "00000000", --  986 - 0x3da  :    0 - 0x0
    "00000000", --  987 - 0x3db  :    0 - 0x0
    "00000000", --  988 - 0x3dc  :    0 - 0x0
    "00000000", --  989 - 0x3dd  :    0 - 0x0
    "00000000", --  990 - 0x3de  :    0 - 0x0
    "00000000", --  991 - 0x3df  :    0 - 0x0
    "00000000", --  992 - 0x3e0  :    0 - 0x0 -- Background 0x7c
    "00000001", --  993 - 0x3e1  :    1 - 0x1
    "00000110", --  994 - 0x3e2  :    6 - 0x6
    "00000111", --  995 - 0x3e3  :    7 - 0x7
    "00000111", --  996 - 0x3e4  :    7 - 0x7
    "00000111", --  997 - 0x3e5  :    7 - 0x7
    "00000001", --  998 - 0x3e6  :    1 - 0x1
    "00000011", --  999 - 0x3e7  :    3 - 0x3
    "00000000", -- 1000 - 0x3e8  :    0 - 0x0 -- Background 0x7d
    "11000000", -- 1001 - 0x3e9  :  192 - 0xc0
    "00110000", -- 1002 - 0x3ea  :   48 - 0x30
    "11110000", -- 1003 - 0x3eb  :  240 - 0xf0
    "11110000", -- 1004 - 0x3ec  :  240 - 0xf0
    "11110000", -- 1005 - 0x3ed  :  240 - 0xf0
    "01000000", -- 1006 - 0x3ee  :   64 - 0x40
    "01000000", -- 1007 - 0x3ef  :   64 - 0x40
    "00000001", -- 1008 - 0x3f0  :    1 - 0x1 -- Background 0x7e
    "00000000", -- 1009 - 0x3f1  :    0 - 0x0
    "00000001", -- 1010 - 0x3f2  :    1 - 0x1
    "00000011", -- 1011 - 0x3f3  :    3 - 0x3
    "00000001", -- 1012 - 0x3f4  :    1 - 0x1
    "00000000", -- 1013 - 0x3f5  :    0 - 0x0
    "00000000", -- 1014 - 0x3f6  :    0 - 0x0
    "00000000", -- 1015 - 0x3f7  :    0 - 0x0
    "01000000", -- 1016 - 0x3f8  :   64 - 0x40 -- Background 0x7f
    "01000000", -- 1017 - 0x3f9  :   64 - 0x40
    "01000000", -- 1018 - 0x3fa  :   64 - 0x40
    "01000000", -- 1019 - 0x3fb  :   64 - 0x40
    "01000000", -- 1020 - 0x3fc  :   64 - 0x40
    "10000000", -- 1021 - 0x3fd  :  128 - 0x80
    "00000000", -- 1022 - 0x3fe  :    0 - 0x0
    "00000000", -- 1023 - 0x3ff  :    0 - 0x0
    "11111111", -- 1024 - 0x400  :  255 - 0xff -- Background 0x80
    "11111111", -- 1025 - 0x401  :  255 - 0xff
    "11111111", -- 1026 - 0x402  :  255 - 0xff
    "11111111", -- 1027 - 0x403  :  255 - 0xff
    "11000000", -- 1028 - 0x404  :  192 - 0xc0
    "11000000", -- 1029 - 0x405  :  192 - 0xc0
    "11000000", -- 1030 - 0x406  :  192 - 0xc0
    "11000111", -- 1031 - 0x407  :  199 - 0xc7
    "11111111", -- 1032 - 0x408  :  255 - 0xff -- Background 0x81
    "11111111", -- 1033 - 0x409  :  255 - 0xff
    "11111111", -- 1034 - 0x40a  :  255 - 0xff
    "11111111", -- 1035 - 0x40b  :  255 - 0xff
    "00000000", -- 1036 - 0x40c  :    0 - 0x0
    "00000000", -- 1037 - 0x40d  :    0 - 0x0
    "00000000", -- 1038 - 0x40e  :    0 - 0x0
    "11111111", -- 1039 - 0x40f  :  255 - 0xff
    "11111111", -- 1040 - 0x410  :  255 - 0xff -- Background 0x82
    "11111111", -- 1041 - 0x411  :  255 - 0xff
    "11111111", -- 1042 - 0x412  :  255 - 0xff
    "11111111", -- 1043 - 0x413  :  255 - 0xff
    "01111111", -- 1044 - 0x414  :  127 - 0x7f
    "00111111", -- 1045 - 0x415  :   63 - 0x3f
    "00011111", -- 1046 - 0x416  :   31 - 0x1f
    "11001111", -- 1047 - 0x417  :  207 - 0xcf
    "11111111", -- 1048 - 0x418  :  255 - 0xff -- Background 0x83
    "11111111", -- 1049 - 0x419  :  255 - 0xff
    "11111111", -- 1050 - 0x41a  :  255 - 0xff
    "11110111", -- 1051 - 0x41b  :  247 - 0xf7
    "11110111", -- 1052 - 0x41c  :  247 - 0xf7
    "11100010", -- 1053 - 0x41d  :  226 - 0xe2
    "11100000", -- 1054 - 0x41e  :  224 - 0xe0
    "11000110", -- 1055 - 0x41f  :  198 - 0xc6
    "11111111", -- 1056 - 0x420  :  255 - 0xff -- Background 0x84
    "11111111", -- 1057 - 0x421  :  255 - 0xff
    "11111111", -- 1058 - 0x422  :  255 - 0xff
    "11111111", -- 1059 - 0x423  :  255 - 0xff
    "10111111", -- 1060 - 0x424  :  191 - 0xbf
    "10111111", -- 1061 - 0x425  :  191 - 0xbf
    "00011111", -- 1062 - 0x426  :   31 - 0x1f
    "00011111", -- 1063 - 0x427  :   31 - 0x1f
    "11111111", -- 1064 - 0x428  :  255 - 0xff -- Background 0x85
    "11111111", -- 1065 - 0x429  :  255 - 0xff
    "11111111", -- 1066 - 0x42a  :  255 - 0xff
    "11111111", -- 1067 - 0x42b  :  255 - 0xff
    "11111110", -- 1068 - 0x42c  :  254 - 0xfe
    "11111000", -- 1069 - 0x42d  :  248 - 0xf8
    "11100000", -- 1070 - 0x42e  :  224 - 0xe0
    "11000000", -- 1071 - 0x42f  :  192 - 0xc0
    "11111111", -- 1072 - 0x430  :  255 - 0xff -- Background 0x86
    "11111111", -- 1073 - 0x431  :  255 - 0xff
    "11111111", -- 1074 - 0x432  :  255 - 0xff
    "11111111", -- 1075 - 0x433  :  255 - 0xff
    "00000111", -- 1076 - 0x434  :    7 - 0x7
    "00000000", -- 1077 - 0x435  :    0 - 0x0
    "00111111", -- 1078 - 0x436  :   63 - 0x3f
    "11111111", -- 1079 - 0x437  :  255 - 0xff
    "11111111", -- 1080 - 0x438  :  255 - 0xff -- Background 0x87
    "11111111", -- 1081 - 0x439  :  255 - 0xff
    "11111111", -- 1082 - 0x43a  :  255 - 0xff
    "11111111", -- 1083 - 0x43b  :  255 - 0xff
    "11111111", -- 1084 - 0x43c  :  255 - 0xff
    "11111111", -- 1085 - 0x43d  :  255 - 0xff
    "00111111", -- 1086 - 0x43e  :   63 - 0x3f
    "11001111", -- 1087 - 0x43f  :  207 - 0xcf
    "11111111", -- 1088 - 0x440  :  255 - 0xff -- Background 0x88
    "11111111", -- 1089 - 0x441  :  255 - 0xff
    "11111111", -- 1090 - 0x442  :  255 - 0xff
    "11111111", -- 1091 - 0x443  :  255 - 0xff
    "11111111", -- 1092 - 0x444  :  255 - 0xff
    "11111111", -- 1093 - 0x445  :  255 - 0xff
    "11111111", -- 1094 - 0x446  :  255 - 0xff
    "11111111", -- 1095 - 0x447  :  255 - 0xff
    "11111111", -- 1096 - 0x448  :  255 - 0xff -- Background 0x89
    "11111111", -- 1097 - 0x449  :  255 - 0xff
    "11111111", -- 1098 - 0x44a  :  255 - 0xff
    "01110111", -- 1099 - 0x44b  :  119 - 0x77
    "00010011", -- 1100 - 0x44c  :   19 - 0x13
    "00000001", -- 1101 - 0x44d  :    1 - 0x1
    "00010000", -- 1102 - 0x44e  :   16 - 0x10
    "00011000", -- 1103 - 0x44f  :   24 - 0x18
    "11111111", -- 1104 - 0x450  :  255 - 0xff -- Background 0x8a
    "11111111", -- 1105 - 0x451  :  255 - 0xff
    "11111111", -- 1106 - 0x452  :  255 - 0xff
    "11111111", -- 1107 - 0x453  :  255 - 0xff
    "11111111", -- 1108 - 0x454  :  255 - 0xff
    "11111111", -- 1109 - 0x455  :  255 - 0xff
    "11111111", -- 1110 - 0x456  :  255 - 0xff
    "01111111", -- 1111 - 0x457  :  127 - 0x7f
    "11111111", -- 1112 - 0x458  :  255 - 0xff -- Background 0x8b
    "11111111", -- 1113 - 0x459  :  255 - 0xff
    "11111111", -- 1114 - 0x45a  :  255 - 0xff
    "11110111", -- 1115 - 0x45b  :  247 - 0xf7
    "11100101", -- 1116 - 0x45c  :  229 - 0xe5
    "11000001", -- 1117 - 0x45d  :  193 - 0xc1
    "10000100", -- 1118 - 0x45e  :  132 - 0x84
    "00001100", -- 1119 - 0x45f  :   12 - 0xc
    "11111111", -- 1120 - 0x460  :  255 - 0xff -- Background 0x8c
    "11111111", -- 1121 - 0x461  :  255 - 0xff
    "11111111", -- 1122 - 0x462  :  255 - 0xff
    "11111111", -- 1123 - 0x463  :  255 - 0xff
    "11111111", -- 1124 - 0x464  :  255 - 0xff
    "01111111", -- 1125 - 0x465  :  127 - 0x7f
    "01111110", -- 1126 - 0x466  :  126 - 0x7e
    "01111110", -- 1127 - 0x467  :  126 - 0x7e
    "11111111", -- 1128 - 0x468  :  255 - 0xff -- Background 0x8d
    "11111111", -- 1129 - 0x469  :  255 - 0xff
    "10111111", -- 1130 - 0x46a  :  191 - 0xbf
    "10110111", -- 1131 - 0x46b  :  183 - 0xb7
    "00010111", -- 1132 - 0x46c  :   23 - 0x17
    "00000011", -- 1133 - 0x46d  :    3 - 0x3
    "00100011", -- 1134 - 0x46e  :   35 - 0x23
    "00100001", -- 1135 - 0x46f  :   33 - 0x21
    "11111111", -- 1136 - 0x470  :  255 - 0xff -- Background 0x8e
    "11111111", -- 1137 - 0x471  :  255 - 0xff
    "11111011", -- 1138 - 0x472  :  251 - 0xfb
    "11111001", -- 1139 - 0x473  :  249 - 0xf9
    "11111000", -- 1140 - 0x474  :  248 - 0xf8
    "11111000", -- 1141 - 0x475  :  248 - 0xf8
    "11111000", -- 1142 - 0x476  :  248 - 0xf8
    "11111000", -- 1143 - 0x477  :  248 - 0xf8
    "11111111", -- 1144 - 0x478  :  255 - 0xff -- Background 0x8f
    "11111111", -- 1145 - 0x479  :  255 - 0xff
    "01111000", -- 1146 - 0x47a  :  120 - 0x78
    "00111000", -- 1147 - 0x47b  :   56 - 0x38
    "00011000", -- 1148 - 0x47c  :   24 - 0x18
    "00001000", -- 1149 - 0x47d  :    8 - 0x8
    "10000000", -- 1150 - 0x47e  :  128 - 0x80
    "11000000", -- 1151 - 0x47f  :  192 - 0xc0
    "11111111", -- 1152 - 0x480  :  255 - 0xff -- Background 0x90
    "11111111", -- 1153 - 0x481  :  255 - 0xff
    "00000001", -- 1154 - 0x482  :    1 - 0x1
    "00000001", -- 1155 - 0x483  :    1 - 0x1
    "00000001", -- 1156 - 0x484  :    1 - 0x1
    "00000000", -- 1157 - 0x485  :    0 - 0x0
    "11111111", -- 1158 - 0x486  :  255 - 0xff
    "11111111", -- 1159 - 0x487  :  255 - 0xff
    "11111111", -- 1160 - 0x488  :  255 - 0xff -- Background 0x91
    "11111111", -- 1161 - 0x489  :  255 - 0xff
    "11111111", -- 1162 - 0x48a  :  255 - 0xff
    "11111111", -- 1163 - 0x48b  :  255 - 0xff
    "11111111", -- 1164 - 0x48c  :  255 - 0xff
    "11111111", -- 1165 - 0x48d  :  255 - 0xff
    "01111111", -- 1166 - 0x48e  :  127 - 0x7f
    "00111111", -- 1167 - 0x48f  :   63 - 0x3f
    "11000111", -- 1168 - 0x490  :  199 - 0xc7 -- Background 0x92
    "11000111", -- 1169 - 0x491  :  199 - 0xc7
    "11000111", -- 1170 - 0x492  :  199 - 0xc7
    "11000111", -- 1171 - 0x493  :  199 - 0xc7
    "11000111", -- 1172 - 0x494  :  199 - 0xc7
    "11000111", -- 1173 - 0x495  :  199 - 0xc7
    "11000111", -- 1174 - 0x496  :  199 - 0xc7
    "11000111", -- 1175 - 0x497  :  199 - 0xc7
    "11111111", -- 1176 - 0x498  :  255 - 0xff -- Background 0x93
    "11111111", -- 1177 - 0x499  :  255 - 0xff
    "11111111", -- 1178 - 0x49a  :  255 - 0xff
    "11111111", -- 1179 - 0x49b  :  255 - 0xff
    "11111001", -- 1180 - 0x49c  :  249 - 0xf9
    "11111001", -- 1181 - 0x49d  :  249 - 0xf9
    "11111111", -- 1182 - 0x49e  :  255 - 0xff
    "11111111", -- 1183 - 0x49f  :  255 - 0xff
    "11110111", -- 1184 - 0x4a0  :  247 - 0xf7 -- Background 0x94
    "11111011", -- 1185 - 0x4a1  :  251 - 0xfb
    "11111011", -- 1186 - 0x4a2  :  251 - 0xfb
    "11111101", -- 1187 - 0x4a3  :  253 - 0xfd
    "11111100", -- 1188 - 0x4a4  :  252 - 0xfc
    "11111100", -- 1189 - 0x4a5  :  252 - 0xfc
    "01111100", -- 1190 - 0x4a6  :  124 - 0x7c
    "01111100", -- 1191 - 0x4a7  :  124 - 0x7c
    "11000111", -- 1192 - 0x4a8  :  199 - 0xc7 -- Background 0x95
    "10001111", -- 1193 - 0x4a9  :  143 - 0x8f
    "10001111", -- 1194 - 0x4aa  :  143 - 0x8f
    "00011111", -- 1195 - 0x4ab  :   31 - 0x1f
    "00011111", -- 1196 - 0x4ac  :   31 - 0x1f
    "00111111", -- 1197 - 0x4ad  :   63 - 0x3f
    "00111111", -- 1198 - 0x4ae  :   63 - 0x3f
    "01111111", -- 1199 - 0x4af  :  127 - 0x7f
    "00001111", -- 1200 - 0x4b0  :   15 - 0xf -- Background 0x96
    "00001111", -- 1201 - 0x4b1  :   15 - 0xf
    "10000111", -- 1202 - 0x4b2  :  135 - 0x87
    "10000111", -- 1203 - 0x4b3  :  135 - 0x87
    "11000010", -- 1204 - 0x4b4  :  194 - 0xc2
    "11000010", -- 1205 - 0x4b5  :  194 - 0xc2
    "11100000", -- 1206 - 0x4b6  :  224 - 0xe0
    "11100000", -- 1207 - 0x4b7  :  224 - 0xe0
    "10000011", -- 1208 - 0x4b8  :  131 - 0x83 -- Background 0x97
    "10001111", -- 1209 - 0x4b9  :  143 - 0x8f
    "00001111", -- 1210 - 0x4ba  :   15 - 0xf
    "00011111", -- 1211 - 0x4bb  :   31 - 0x1f
    "00011111", -- 1212 - 0x4bc  :   31 - 0x1f
    "00111111", -- 1213 - 0x4bd  :   63 - 0x3f
    "00111111", -- 1214 - 0x4be  :   63 - 0x3f
    "00111111", -- 1215 - 0x4bf  :   63 - 0x3f
    "11111111", -- 1216 - 0x4c0  :  255 - 0xff -- Background 0x98
    "11111111", -- 1217 - 0x4c1  :  255 - 0xff
    "11111111", -- 1218 - 0x4c2  :  255 - 0xff
    "11111110", -- 1219 - 0x4c3  :  254 - 0xfe
    "11111001", -- 1220 - 0x4c4  :  249 - 0xf9
    "11100111", -- 1221 - 0x4c5  :  231 - 0xe7
    "11111100", -- 1222 - 0x4c6  :  252 - 0xfc
    "11110000", -- 1223 - 0x4c7  :  240 - 0xf0
    "11110111", -- 1224 - 0x4c8  :  247 - 0xf7 -- Background 0x99
    "11111011", -- 1225 - 0x4c9  :  251 - 0xfb
    "11111011", -- 1226 - 0x4ca  :  251 - 0xfb
    "01110011", -- 1227 - 0x4cb  :  115 - 0x73
    "11000001", -- 1228 - 0x4cc  :  193 - 0xc1
    "00000011", -- 1229 - 0x4cd  :    3 - 0x3
    "00001111", -- 1230 - 0x4ce  :   15 - 0xf
    "00111111", -- 1231 - 0x4cf  :   63 - 0x3f
    "11111111", -- 1232 - 0x4d0  :  255 - 0xff -- Background 0x9a
    "11111111", -- 1233 - 0x4d1  :  255 - 0xff
    "11111111", -- 1234 - 0x4d2  :  255 - 0xff
    "10000000", -- 1235 - 0x4d3  :  128 - 0x80
    "10000000", -- 1236 - 0x4d4  :  128 - 0x80
    "10000000", -- 1237 - 0x4d5  :  128 - 0x80
    "10001111", -- 1238 - 0x4d6  :  143 - 0x8f
    "10001111", -- 1239 - 0x4d7  :  143 - 0x8f
    "11111111", -- 1240 - 0x4d8  :  255 - 0xff -- Background 0x9b
    "11111111", -- 1241 - 0x4d9  :  255 - 0xff
    "11111111", -- 1242 - 0x4da  :  255 - 0xff
    "00001111", -- 1243 - 0x4db  :   15 - 0xf
    "00001111", -- 1244 - 0x4dc  :   15 - 0xf
    "00000111", -- 1245 - 0x4dd  :    7 - 0x7
    "11110111", -- 1246 - 0x4de  :  247 - 0xf7
    "11110001", -- 1247 - 0x4df  :  241 - 0xf1
    "00011100", -- 1248 - 0x4e0  :   28 - 0x1c -- Background 0x9c
    "00011110", -- 1249 - 0x4e1  :   30 - 0x1e
    "00011111", -- 1250 - 0x4e2  :   31 - 0x1f
    "00011111", -- 1251 - 0x4e3  :   31 - 0x1f
    "00011111", -- 1252 - 0x4e4  :   31 - 0x1f
    "00011111", -- 1253 - 0x4e5  :   31 - 0x1f
    "00011111", -- 1254 - 0x4e6  :   31 - 0x1f
    "00011111", -- 1255 - 0x4e7  :   31 - 0x1f
    "00111110", -- 1256 - 0x4e8  :   62 - 0x3e -- Background 0x9d
    "00011100", -- 1257 - 0x4e9  :   28 - 0x1c
    "00001000", -- 1258 - 0x4ea  :    8 - 0x8
    "10000000", -- 1259 - 0x4eb  :  128 - 0x80
    "11000001", -- 1260 - 0x4ec  :  193 - 0xc1
    "11100011", -- 1261 - 0x4ed  :  227 - 0xe3
    "11110111", -- 1262 - 0x4ee  :  247 - 0xf7
    "11111111", -- 1263 - 0x4ef  :  255 - 0xff
    "00011100", -- 1264 - 0x4f0  :   28 - 0x1c -- Background 0x9e
    "00111100", -- 1265 - 0x4f1  :   60 - 0x3c
    "01111100", -- 1266 - 0x4f2  :  124 - 0x7c
    "11111100", -- 1267 - 0x4f3  :  252 - 0xfc
    "11111100", -- 1268 - 0x4f4  :  252 - 0xfc
    "11111100", -- 1269 - 0x4f5  :  252 - 0xfc
    "11111100", -- 1270 - 0x4f6  :  252 - 0xfc
    "11111100", -- 1271 - 0x4f7  :  252 - 0xfc
    "01111100", -- 1272 - 0x4f8  :  124 - 0x7c -- Background 0x9f
    "01111100", -- 1273 - 0x4f9  :  124 - 0x7c
    "01111000", -- 1274 - 0x4fa  :  120 - 0x78
    "01111000", -- 1275 - 0x4fb  :  120 - 0x78
    "01110001", -- 1276 - 0x4fc  :  113 - 0x71
    "01110001", -- 1277 - 0x4fd  :  113 - 0x71
    "01100011", -- 1278 - 0x4fe  :   99 - 0x63
    "01100011", -- 1279 - 0x4ff  :   99 - 0x63
    "01110001", -- 1280 - 0x500  :  113 - 0x71 -- Background 0xa0
    "01110000", -- 1281 - 0x501  :  112 - 0x70
    "11111000", -- 1282 - 0x502  :  248 - 0xf8
    "11111000", -- 1283 - 0x503  :  248 - 0xf8
    "11111100", -- 1284 - 0x504  :  252 - 0xfc
    "11111100", -- 1285 - 0x505  :  252 - 0xfc
    "11111110", -- 1286 - 0x506  :  254 - 0xfe
    "11111110", -- 1287 - 0x507  :  254 - 0xfe
    "11111000", -- 1288 - 0x508  :  248 - 0xf8 -- Background 0xa1
    "11111000", -- 1289 - 0x509  :  248 - 0xf8
    "11111000", -- 1290 - 0x50a  :  248 - 0xf8
    "01111000", -- 1291 - 0x50b  :  120 - 0x78
    "01111000", -- 1292 - 0x50c  :  120 - 0x78
    "00111000", -- 1293 - 0x50d  :   56 - 0x38
    "00111000", -- 1294 - 0x50e  :   56 - 0x38
    "00011000", -- 1295 - 0x50f  :   24 - 0x18
    "11100000", -- 1296 - 0x510  :  224 - 0xe0 -- Background 0xa2
    "11110000", -- 1297 - 0x511  :  240 - 0xf0
    "11111000", -- 1298 - 0x512  :  248 - 0xf8
    "11111000", -- 1299 - 0x513  :  248 - 0xf8
    "11111100", -- 1300 - 0x514  :  252 - 0xfc
    "11111100", -- 1301 - 0x515  :  252 - 0xfc
    "11111110", -- 1302 - 0x516  :  254 - 0xfe
    "11111111", -- 1303 - 0x517  :  255 - 0xff
    "11111111", -- 1304 - 0x518  :  255 - 0xff -- Background 0xa3
    "11111111", -- 1305 - 0x519  :  255 - 0xff
    "11111111", -- 1306 - 0x51a  :  255 - 0xff
    "11111111", -- 1307 - 0x51b  :  255 - 0xff
    "11111111", -- 1308 - 0x51c  :  255 - 0xff
    "11111111", -- 1309 - 0x51d  :  255 - 0xff
    "11111111", -- 1310 - 0x51e  :  255 - 0xff
    "11111111", -- 1311 - 0x51f  :  255 - 0xff
    "00011111", -- 1312 - 0x520  :   31 - 0x1f -- Background 0xa4
    "00011111", -- 1313 - 0x521  :   31 - 0x1f
    "00011111", -- 1314 - 0x522  :   31 - 0x1f
    "00011111", -- 1315 - 0x523  :   31 - 0x1f
    "00011111", -- 1316 - 0x524  :   31 - 0x1f
    "00011111", -- 1317 - 0x525  :   31 - 0x1f
    "00011111", -- 1318 - 0x526  :   31 - 0x1f
    "00011111", -- 1319 - 0x527  :   31 - 0x1f
    "11111000", -- 1320 - 0x528  :  248 - 0xf8 -- Background 0xa5
    "11111111", -- 1321 - 0x529  :  255 - 0xff
    "11111111", -- 1322 - 0x52a  :  255 - 0xff
    "11111000", -- 1323 - 0x52b  :  248 - 0xf8
    "11111000", -- 1324 - 0x52c  :  248 - 0xf8
    "11111000", -- 1325 - 0x52d  :  248 - 0xf8
    "11111000", -- 1326 - 0x52e  :  248 - 0xf8
    "11111000", -- 1327 - 0x52f  :  248 - 0xf8
    "11111100", -- 1328 - 0x530  :  252 - 0xfc -- Background 0xa6
    "11111000", -- 1329 - 0x531  :  248 - 0xf8
    "11110000", -- 1330 - 0x532  :  240 - 0xf0
    "00000001", -- 1331 - 0x533  :    1 - 0x1
    "00000001", -- 1332 - 0x534  :    1 - 0x1
    "00000011", -- 1333 - 0x535  :    3 - 0x3
    "11000011", -- 1334 - 0x536  :  195 - 0xc3
    "10000111", -- 1335 - 0x537  :  135 - 0x87
    "01111111", -- 1336 - 0x538  :  127 - 0x7f -- Background 0xa7
    "11111001", -- 1337 - 0x539  :  249 - 0xf9
    "11111001", -- 1338 - 0x53a  :  249 - 0xf9
    "11111111", -- 1339 - 0x53b  :  255 - 0xff
    "11111110", -- 1340 - 0x53c  :  254 - 0xfe
    "11111100", -- 1341 - 0x53d  :  252 - 0xfc
    "11111111", -- 1342 - 0x53e  :  255 - 0xff
    "11111111", -- 1343 - 0x53f  :  255 - 0xff
    "11110000", -- 1344 - 0x540  :  240 - 0xf0 -- Background 0xa8
    "11110000", -- 1345 - 0x541  :  240 - 0xf0
    "11111000", -- 1346 - 0x542  :  248 - 0xf8
    "01111000", -- 1347 - 0x543  :  120 - 0x78
    "11111100", -- 1348 - 0x544  :  252 - 0xfc
    "11110100", -- 1349 - 0x545  :  244 - 0xf4
    "11110110", -- 1350 - 0x546  :  246 - 0xf6
    "11111010", -- 1351 - 0x547  :  250 - 0xfa
    "00111111", -- 1352 - 0x548  :   63 - 0x3f -- Background 0xa9
    "00111111", -- 1353 - 0x549  :   63 - 0x3f
    "00111111", -- 1354 - 0x54a  :   63 - 0x3f
    "00111111", -- 1355 - 0x54b  :   63 - 0x3f
    "00111111", -- 1356 - 0x54c  :   63 - 0x3f
    "00011111", -- 1357 - 0x54d  :   31 - 0x1f
    "00001111", -- 1358 - 0x54e  :   15 - 0xf
    "00000111", -- 1359 - 0x54f  :    7 - 0x7
    "11100000", -- 1360 - 0x550  :  224 - 0xe0 -- Background 0xaa
    "11111000", -- 1361 - 0x551  :  248 - 0xf8
    "11111111", -- 1362 - 0x552  :  255 - 0xff
    "11110011", -- 1363 - 0x553  :  243 - 0xf3
    "11111100", -- 1364 - 0x554  :  252 - 0xfc
    "11111111", -- 1365 - 0x555  :  255 - 0xff
    "11111111", -- 1366 - 0x556  :  255 - 0xff
    "11111111", -- 1367 - 0x557  :  255 - 0xff
    "11111111", -- 1368 - 0x558  :  255 - 0xff -- Background 0xab
    "11111111", -- 1369 - 0x559  :  255 - 0xff
    "00111111", -- 1370 - 0x55a  :   63 - 0x3f
    "11001111", -- 1371 - 0x55b  :  207 - 0xcf
    "11110011", -- 1372 - 0x55c  :  243 - 0xf3
    "00111101", -- 1373 - 0x55d  :   61 - 0x3d
    "11011000", -- 1374 - 0x55e  :  216 - 0xd8
    "10110000", -- 1375 - 0x55f  :  176 - 0xb0
    "10001111", -- 1376 - 0x560  :  143 - 0x8f -- Background 0xac
    "11101111", -- 1377 - 0x561  :  239 - 0xef
    "11100000", -- 1378 - 0x562  :  224 - 0xe0
    "11111000", -- 1379 - 0x563  :  248 - 0xf8
    "11111000", -- 1380 - 0x564  :  248 - 0xf8
    "11111111", -- 1381 - 0x565  :  255 - 0xff
    "11111111", -- 1382 - 0x566  :  255 - 0xff
    "11111111", -- 1383 - 0x567  :  255 - 0xff
    "11110001", -- 1384 - 0x568  :  241 - 0xf1 -- Background 0xad
    "11110001", -- 1385 - 0x569  :  241 - 0xf1
    "00000001", -- 1386 - 0x56a  :    1 - 0x1
    "00000001", -- 1387 - 0x56b  :    1 - 0x1
    "00000001", -- 1388 - 0x56c  :    1 - 0x1
    "11111111", -- 1389 - 0x56d  :  255 - 0xff
    "11111111", -- 1390 - 0x56e  :  255 - 0xff
    "11111111", -- 1391 - 0x56f  :  255 - 0xff
    "00011111", -- 1392 - 0x570  :   31 - 0x1f -- Background 0xae
    "00011111", -- 1393 - 0x571  :   31 - 0x1f
    "00011111", -- 1394 - 0x572  :   31 - 0x1f
    "00011111", -- 1395 - 0x573  :   31 - 0x1f
    "00011111", -- 1396 - 0x574  :   31 - 0x1f
    "00011111", -- 1397 - 0x575  :   31 - 0x1f
    "00011111", -- 1398 - 0x576  :   31 - 0x1f
    "00011111", -- 1399 - 0x577  :   31 - 0x1f
    "11111100", -- 1400 - 0x578  :  252 - 0xfc -- Background 0xaf
    "11111100", -- 1401 - 0x579  :  252 - 0xfc
    "11111100", -- 1402 - 0x57a  :  252 - 0xfc
    "11111100", -- 1403 - 0x57b  :  252 - 0xfc
    "11110100", -- 1404 - 0x57c  :  244 - 0xf4
    "11110100", -- 1405 - 0x57d  :  244 - 0xf4
    "11110100", -- 1406 - 0x57e  :  244 - 0xf4
    "11110100", -- 1407 - 0x57f  :  244 - 0xf4
    "00001100", -- 1408 - 0x580  :   12 - 0xc -- Background 0xb0
    "00011100", -- 1409 - 0x581  :   28 - 0x1c
    "00001100", -- 1410 - 0x582  :   12 - 0xc
    "00001100", -- 1411 - 0x583  :   12 - 0xc
    "00001100", -- 1412 - 0x584  :   12 - 0xc
    "00001100", -- 1413 - 0x585  :   12 - 0xc
    "00111111", -- 1414 - 0x586  :   63 - 0x3f
    "00000000", -- 1415 - 0x587  :    0 - 0x0
    "00111110", -- 1416 - 0x588  :   62 - 0x3e -- Background 0xb1
    "01100011", -- 1417 - 0x589  :   99 - 0x63
    "00000111", -- 1418 - 0x58a  :    7 - 0x7
    "00011110", -- 1419 - 0x58b  :   30 - 0x1e
    "00111100", -- 1420 - 0x58c  :   60 - 0x3c
    "01110000", -- 1421 - 0x58d  :  112 - 0x70
    "01111111", -- 1422 - 0x58e  :  127 - 0x7f
    "00000000", -- 1423 - 0x58f  :    0 - 0x0
    "01111110", -- 1424 - 0x590  :  126 - 0x7e -- Background 0xb2
    "01100011", -- 1425 - 0x591  :   99 - 0x63
    "01100011", -- 1426 - 0x592  :   99 - 0x63
    "01100011", -- 1427 - 0x593  :   99 - 0x63
    "01111110", -- 1428 - 0x594  :  126 - 0x7e
    "01100000", -- 1429 - 0x595  :   96 - 0x60
    "01100000", -- 1430 - 0x596  :   96 - 0x60
    "00000000", -- 1431 - 0x597  :    0 - 0x0
    "01100011", -- 1432 - 0x598  :   99 - 0x63 -- Background 0xb3
    "01100011", -- 1433 - 0x599  :   99 - 0x63
    "01100011", -- 1434 - 0x59a  :   99 - 0x63
    "01100011", -- 1435 - 0x59b  :   99 - 0x63
    "01100011", -- 1436 - 0x59c  :   99 - 0x63
    "01100011", -- 1437 - 0x59d  :   99 - 0x63
    "00111110", -- 1438 - 0x59e  :   62 - 0x3e
    "00000000", -- 1439 - 0x59f  :    0 - 0x0
    "01100011", -- 1440 - 0x5a0  :   99 - 0x63 -- Background 0xb4
    "01100011", -- 1441 - 0x5a1  :   99 - 0x63
    "01100011", -- 1442 - 0x5a2  :   99 - 0x63
    "01111111", -- 1443 - 0x5a3  :  127 - 0x7f
    "01100011", -- 1444 - 0x5a4  :   99 - 0x63
    "01100011", -- 1445 - 0x5a5  :   99 - 0x63
    "01100011", -- 1446 - 0x5a6  :   99 - 0x63
    "00000000", -- 1447 - 0x5a7  :    0 - 0x0
    "00111111", -- 1448 - 0x5a8  :   63 - 0x3f -- Background 0xb5
    "00001100", -- 1449 - 0x5a9  :   12 - 0xc
    "00001100", -- 1450 - 0x5aa  :   12 - 0xc
    "00001100", -- 1451 - 0x5ab  :   12 - 0xc
    "00001100", -- 1452 - 0x5ac  :   12 - 0xc
    "00001100", -- 1453 - 0x5ad  :   12 - 0xc
    "00111111", -- 1454 - 0x5ae  :   63 - 0x3f
    "00000000", -- 1455 - 0x5af  :    0 - 0x0
    "00000000", -- 1456 - 0x5b0  :    0 - 0x0 -- Background 0xb6
    "00000000", -- 1457 - 0x5b1  :    0 - 0x0
    "00000000", -- 1458 - 0x5b2  :    0 - 0x0
    "01111110", -- 1459 - 0x5b3  :  126 - 0x7e
    "00000000", -- 1460 - 0x5b4  :    0 - 0x0
    "00000000", -- 1461 - 0x5b5  :    0 - 0x0
    "00000000", -- 1462 - 0x5b6  :    0 - 0x0
    "00000000", -- 1463 - 0x5b7  :    0 - 0x0
    "00111100", -- 1464 - 0x5b8  :   60 - 0x3c -- Background 0xb7
    "01100110", -- 1465 - 0x5b9  :  102 - 0x66
    "01100000", -- 1466 - 0x5ba  :   96 - 0x60
    "00111110", -- 1467 - 0x5bb  :   62 - 0x3e
    "00000011", -- 1468 - 0x5bc  :    3 - 0x3
    "01100011", -- 1469 - 0x5bd  :   99 - 0x63
    "00111110", -- 1470 - 0x5be  :   62 - 0x3e
    "00000000", -- 1471 - 0x5bf  :    0 - 0x0
    "00011110", -- 1472 - 0x5c0  :   30 - 0x1e -- Background 0xb8
    "00110011", -- 1473 - 0x5c1  :   51 - 0x33
    "01100000", -- 1474 - 0x5c2  :   96 - 0x60
    "01100000", -- 1475 - 0x5c3  :   96 - 0x60
    "01100000", -- 1476 - 0x5c4  :   96 - 0x60
    "00110011", -- 1477 - 0x5c5  :   51 - 0x33
    "00011110", -- 1478 - 0x5c6  :   30 - 0x1e
    "00000000", -- 1479 - 0x5c7  :    0 - 0x0
    "00111110", -- 1480 - 0x5c8  :   62 - 0x3e -- Background 0xb9
    "01100011", -- 1481 - 0x5c9  :   99 - 0x63
    "01100011", -- 1482 - 0x5ca  :   99 - 0x63
    "01100011", -- 1483 - 0x5cb  :   99 - 0x63
    "01100011", -- 1484 - 0x5cc  :   99 - 0x63
    "01100011", -- 1485 - 0x5cd  :   99 - 0x63
    "00111110", -- 1486 - 0x5ce  :   62 - 0x3e
    "00000000", -- 1487 - 0x5cf  :    0 - 0x0
    "01111110", -- 1488 - 0x5d0  :  126 - 0x7e -- Background 0xba
    "01100011", -- 1489 - 0x5d1  :   99 - 0x63
    "01100011", -- 1490 - 0x5d2  :   99 - 0x63
    "01100111", -- 1491 - 0x5d3  :  103 - 0x67
    "01111100", -- 1492 - 0x5d4  :  124 - 0x7c
    "01101110", -- 1493 - 0x5d5  :  110 - 0x6e
    "01100111", -- 1494 - 0x5d6  :  103 - 0x67
    "00000000", -- 1495 - 0x5d7  :    0 - 0x0
    "01111111", -- 1496 - 0x5d8  :  127 - 0x7f -- Background 0xbb
    "01100000", -- 1497 - 0x5d9  :   96 - 0x60
    "01100000", -- 1498 - 0x5da  :   96 - 0x60
    "01111110", -- 1499 - 0x5db  :  126 - 0x7e
    "01100000", -- 1500 - 0x5dc  :   96 - 0x60
    "01100000", -- 1501 - 0x5dd  :   96 - 0x60
    "01111111", -- 1502 - 0x5de  :  127 - 0x7f
    "00000000", -- 1503 - 0x5df  :    0 - 0x0
    "00000000", -- 1504 - 0x5e0  :    0 - 0x0 -- Background 0xbc
    "00100010", -- 1505 - 0x5e1  :   34 - 0x22
    "01100101", -- 1506 - 0x5e2  :  101 - 0x65
    "00100101", -- 1507 - 0x5e3  :   37 - 0x25
    "00100101", -- 1508 - 0x5e4  :   37 - 0x25
    "01110010", -- 1509 - 0x5e5  :  114 - 0x72
    "00000000", -- 1510 - 0x5e6  :    0 - 0x0
    "00000000", -- 1511 - 0x5e7  :    0 - 0x0
    "00000000", -- 1512 - 0x5e8  :    0 - 0x0 -- Background 0xbd
    "01110010", -- 1513 - 0x5e9  :  114 - 0x72
    "01000101", -- 1514 - 0x5ea  :   69 - 0x45
    "01100101", -- 1515 - 0x5eb  :  101 - 0x65
    "00010101", -- 1516 - 0x5ec  :   21 - 0x15
    "01100010", -- 1517 - 0x5ed  :   98 - 0x62
    "00000000", -- 1518 - 0x5ee  :    0 - 0x0
    "00000000", -- 1519 - 0x5ef  :    0 - 0x0
    "00000000", -- 1520 - 0x5f0  :    0 - 0x0 -- Background 0xbe
    "01100111", -- 1521 - 0x5f1  :  103 - 0x67
    "01010010", -- 1522 - 0x5f2  :   82 - 0x52
    "01100010", -- 1523 - 0x5f3  :   98 - 0x62
    "01000010", -- 1524 - 0x5f4  :   66 - 0x42
    "01000010", -- 1525 - 0x5f5  :   66 - 0x42
    "00000000", -- 1526 - 0x5f6  :    0 - 0x0
    "00000000", -- 1527 - 0x5f7  :    0 - 0x0
    "00000000", -- 1528 - 0x5f8  :    0 - 0x0 -- Background 0xbf
    "01100000", -- 1529 - 0x5f9  :   96 - 0x60
    "10000000", -- 1530 - 0x5fa  :  128 - 0x80
    "01000000", -- 1531 - 0x5fb  :   64 - 0x40
    "00100000", -- 1532 - 0x5fc  :   32 - 0x20
    "11000110", -- 1533 - 0x5fd  :  198 - 0xc6
    "00000000", -- 1534 - 0x5fe  :    0 - 0x0
    "00000000", -- 1535 - 0x5ff  :    0 - 0x0
    "01100011", -- 1536 - 0x600  :   99 - 0x63 -- Background 0xc0
    "01100110", -- 1537 - 0x601  :  102 - 0x66
    "01101100", -- 1538 - 0x602  :  108 - 0x6c
    "01111000", -- 1539 - 0x603  :  120 - 0x78
    "01111100", -- 1540 - 0x604  :  124 - 0x7c
    "01100110", -- 1541 - 0x605  :  102 - 0x66
    "01100011", -- 1542 - 0x606  :   99 - 0x63
    "00000000", -- 1543 - 0x607  :    0 - 0x0
    "00111111", -- 1544 - 0x608  :   63 - 0x3f -- Background 0xc1
    "00001100", -- 1545 - 0x609  :   12 - 0xc
    "00001100", -- 1546 - 0x60a  :   12 - 0xc
    "00001100", -- 1547 - 0x60b  :   12 - 0xc
    "00001100", -- 1548 - 0x60c  :   12 - 0xc
    "00001100", -- 1549 - 0x60d  :   12 - 0xc
    "00111111", -- 1550 - 0x60e  :   63 - 0x3f
    "00000000", -- 1551 - 0x60f  :    0 - 0x0
    "01100011", -- 1552 - 0x610  :   99 - 0x63 -- Background 0xc2
    "01110111", -- 1553 - 0x611  :  119 - 0x77
    "01111111", -- 1554 - 0x612  :  127 - 0x7f
    "01111111", -- 1555 - 0x613  :  127 - 0x7f
    "01101011", -- 1556 - 0x614  :  107 - 0x6b
    "01100011", -- 1557 - 0x615  :   99 - 0x63
    "01100011", -- 1558 - 0x616  :   99 - 0x63
    "00000000", -- 1559 - 0x617  :    0 - 0x0
    "00011100", -- 1560 - 0x618  :   28 - 0x1c -- Background 0xc3
    "00110110", -- 1561 - 0x619  :   54 - 0x36
    "01100011", -- 1562 - 0x61a  :   99 - 0x63
    "01100011", -- 1563 - 0x61b  :   99 - 0x63
    "01111111", -- 1564 - 0x61c  :  127 - 0x7f
    "01100011", -- 1565 - 0x61d  :   99 - 0x63
    "01100011", -- 1566 - 0x61e  :   99 - 0x63
    "00000000", -- 1567 - 0x61f  :    0 - 0x0
    "00011111", -- 1568 - 0x620  :   31 - 0x1f -- Background 0xc4
    "00110000", -- 1569 - 0x621  :   48 - 0x30
    "01100000", -- 1570 - 0x622  :   96 - 0x60
    "01100111", -- 1571 - 0x623  :  103 - 0x67
    "01100011", -- 1572 - 0x624  :   99 - 0x63
    "00110011", -- 1573 - 0x625  :   51 - 0x33
    "00011111", -- 1574 - 0x626  :   31 - 0x1f
    "00000000", -- 1575 - 0x627  :    0 - 0x0
    "01100011", -- 1576 - 0x628  :   99 - 0x63 -- Background 0xc5
    "01100011", -- 1577 - 0x629  :   99 - 0x63
    "01100011", -- 1578 - 0x62a  :   99 - 0x63
    "01100011", -- 1579 - 0x62b  :   99 - 0x63
    "01100011", -- 1580 - 0x62c  :   99 - 0x63
    "01100011", -- 1581 - 0x62d  :   99 - 0x63
    "00111110", -- 1582 - 0x62e  :   62 - 0x3e
    "00000000", -- 1583 - 0x62f  :    0 - 0x0
    "01111110", -- 1584 - 0x630  :  126 - 0x7e -- Background 0xc6
    "01100011", -- 1585 - 0x631  :   99 - 0x63
    "01100011", -- 1586 - 0x632  :   99 - 0x63
    "01100111", -- 1587 - 0x633  :  103 - 0x67
    "01111100", -- 1588 - 0x634  :  124 - 0x7c
    "01101110", -- 1589 - 0x635  :  110 - 0x6e
    "01100111", -- 1590 - 0x636  :  103 - 0x67
    "00000000", -- 1591 - 0x637  :    0 - 0x0
    "01111111", -- 1592 - 0x638  :  127 - 0x7f -- Background 0xc7
    "01100000", -- 1593 - 0x639  :   96 - 0x60
    "01100000", -- 1594 - 0x63a  :   96 - 0x60
    "01111110", -- 1595 - 0x63b  :  126 - 0x7e
    "01100000", -- 1596 - 0x63c  :   96 - 0x60
    "01100000", -- 1597 - 0x63d  :   96 - 0x60
    "01111111", -- 1598 - 0x63e  :  127 - 0x7f
    "00000000", -- 1599 - 0x63f  :    0 - 0x0
    "00110110", -- 1600 - 0x640  :   54 - 0x36 -- Background 0xc8
    "00110110", -- 1601 - 0x641  :   54 - 0x36
    "00010010", -- 1602 - 0x642  :   18 - 0x12
    "00000000", -- 1603 - 0x643  :    0 - 0x0
    "00000000", -- 1604 - 0x644  :    0 - 0x0
    "00000000", -- 1605 - 0x645  :    0 - 0x0
    "00000000", -- 1606 - 0x646  :    0 - 0x0
    "00000000", -- 1607 - 0x647  :    0 - 0x0
    "00111110", -- 1608 - 0x648  :   62 - 0x3e -- Background 0xc9
    "01100011", -- 1609 - 0x649  :   99 - 0x63
    "01100011", -- 1610 - 0x64a  :   99 - 0x63
    "01100011", -- 1611 - 0x64b  :   99 - 0x63
    "01100011", -- 1612 - 0x64c  :   99 - 0x63
    "01100011", -- 1613 - 0x64d  :   99 - 0x63
    "00111110", -- 1614 - 0x64e  :   62 - 0x3e
    "00000000", -- 1615 - 0x64f  :    0 - 0x0
    "00111100", -- 1616 - 0x650  :   60 - 0x3c -- Background 0xca
    "01100110", -- 1617 - 0x651  :  102 - 0x66
    "01100000", -- 1618 - 0x652  :   96 - 0x60
    "00111110", -- 1619 - 0x653  :   62 - 0x3e
    "00000011", -- 1620 - 0x654  :    3 - 0x3
    "01100011", -- 1621 - 0x655  :   99 - 0x63
    "00111110", -- 1622 - 0x656  :   62 - 0x3e
    "00000000", -- 1623 - 0x657  :    0 - 0x0
    "00000000", -- 1624 - 0x658  :    0 - 0x0 -- Background 0xcb
    "00000000", -- 1625 - 0x659  :    0 - 0x0
    "00000000", -- 1626 - 0x65a  :    0 - 0x0
    "00000000", -- 1627 - 0x65b  :    0 - 0x0
    "00000000", -- 1628 - 0x65c  :    0 - 0x0
    "00000000", -- 1629 - 0x65d  :    0 - 0x0
    "00000000", -- 1630 - 0x65e  :    0 - 0x0
    "00000000", -- 1631 - 0x65f  :    0 - 0x0
    "00000000", -- 1632 - 0x660  :    0 - 0x0 -- Background 0xcc
    "00000000", -- 1633 - 0x661  :    0 - 0x0
    "00000000", -- 1634 - 0x662  :    0 - 0x0
    "00000000", -- 1635 - 0x663  :    0 - 0x0
    "00000000", -- 1636 - 0x664  :    0 - 0x0
    "00000000", -- 1637 - 0x665  :    0 - 0x0
    "00000000", -- 1638 - 0x666  :    0 - 0x0
    "00000000", -- 1639 - 0x667  :    0 - 0x0
    "00000000", -- 1640 - 0x668  :    0 - 0x0 -- Background 0xcd
    "00000000", -- 1641 - 0x669  :    0 - 0x0
    "00000000", -- 1642 - 0x66a  :    0 - 0x0
    "00000000", -- 1643 - 0x66b  :    0 - 0x0
    "00000000", -- 1644 - 0x66c  :    0 - 0x0
    "00000000", -- 1645 - 0x66d  :    0 - 0x0
    "00000000", -- 1646 - 0x66e  :    0 - 0x0
    "00000000", -- 1647 - 0x66f  :    0 - 0x0
    "00000000", -- 1648 - 0x670  :    0 - 0x0 -- Background 0xce
    "00000000", -- 1649 - 0x671  :    0 - 0x0
    "00000000", -- 1650 - 0x672  :    0 - 0x0
    "00000000", -- 1651 - 0x673  :    0 - 0x0
    "00000000", -- 1652 - 0x674  :    0 - 0x0
    "00000000", -- 1653 - 0x675  :    0 - 0x0
    "00000000", -- 1654 - 0x676  :    0 - 0x0
    "00000000", -- 1655 - 0x677  :    0 - 0x0
    "00000000", -- 1656 - 0x678  :    0 - 0x0 -- Background 0xcf
    "00000000", -- 1657 - 0x679  :    0 - 0x0
    "00000000", -- 1658 - 0x67a  :    0 - 0x0
    "00000000", -- 1659 - 0x67b  :    0 - 0x0
    "00000000", -- 1660 - 0x67c  :    0 - 0x0
    "00000000", -- 1661 - 0x67d  :    0 - 0x0
    "00000000", -- 1662 - 0x67e  :    0 - 0x0
    "00000000", -- 1663 - 0x67f  :    0 - 0x0
    "01000111", -- 1664 - 0x680  :   71 - 0x47 -- Background 0xd0
    "01000111", -- 1665 - 0x681  :   71 - 0x47
    "00001111", -- 1666 - 0x682  :   15 - 0xf
    "00001111", -- 1667 - 0x683  :   15 - 0xf
    "00011111", -- 1668 - 0x684  :   31 - 0x1f
    "00011111", -- 1669 - 0x685  :   31 - 0x1f
    "00111111", -- 1670 - 0x686  :   63 - 0x3f
    "00111111", -- 1671 - 0x687  :   63 - 0x3f
    "11111111", -- 1672 - 0x688  :  255 - 0xff -- Background 0xd1
    "11001111", -- 1673 - 0x689  :  207 - 0xcf
    "11001111", -- 1674 - 0x68a  :  207 - 0xcf
    "11111011", -- 1675 - 0x68b  :  251 - 0xfb
    "11110111", -- 1676 - 0x68c  :  247 - 0xf7
    "11100111", -- 1677 - 0x68d  :  231 - 0xe7
    "11111111", -- 1678 - 0x68e  :  255 - 0xff
    "11111111", -- 1679 - 0x68f  :  255 - 0xff
    "00011000", -- 1680 - 0x690  :   24 - 0x18 -- Background 0xd2
    "00001000", -- 1681 - 0x691  :    8 - 0x8
    "10001000", -- 1682 - 0x692  :  136 - 0x88
    "10000000", -- 1683 - 0x693  :  128 - 0x80
    "01000000", -- 1684 - 0x694  :   64 - 0x40
    "01000000", -- 1685 - 0x695  :   64 - 0x40
    "10100000", -- 1686 - 0x696  :  160 - 0xa0
    "10100000", -- 1687 - 0x697  :  160 - 0xa0
    "11111111", -- 1688 - 0x698  :  255 - 0xff -- Background 0xd3
    "11111111", -- 1689 - 0x699  :  255 - 0xff
    "11111111", -- 1690 - 0x69a  :  255 - 0xff
    "11111111", -- 1691 - 0x69b  :  255 - 0xff
    "11111101", -- 1692 - 0x69c  :  253 - 0xfd
    "11111101", -- 1693 - 0x69d  :  253 - 0xfd
    "11111101", -- 1694 - 0x69e  :  253 - 0xfd
    "11111101", -- 1695 - 0x69f  :  253 - 0xfd
    "11000111", -- 1696 - 0x6a0  :  199 - 0xc7 -- Background 0xd4
    "11110111", -- 1697 - 0x6a1  :  247 - 0xf7
    "11110000", -- 1698 - 0x6a2  :  240 - 0xf0
    "11111000", -- 1699 - 0x6a3  :  248 - 0xf8
    "11111000", -- 1700 - 0x6a4  :  248 - 0xf8
    "11111111", -- 1701 - 0x6a5  :  255 - 0xff
    "11111111", -- 1702 - 0x6a6  :  255 - 0xff
    "11111111", -- 1703 - 0x6a7  :  255 - 0xff
    "11111000", -- 1704 - 0x6a8  :  248 - 0xf8 -- Background 0xd5
    "11111000", -- 1705 - 0x6a9  :  248 - 0xf8
    "00000000", -- 1706 - 0x6aa  :    0 - 0x0
    "00000000", -- 1707 - 0x6ab  :    0 - 0x0
    "00000000", -- 1708 - 0x6ac  :    0 - 0x0
    "11111111", -- 1709 - 0x6ad  :  255 - 0xff
    "11111111", -- 1710 - 0x6ae  :  255 - 0xff
    "11111111", -- 1711 - 0x6af  :  255 - 0xff
    "10001111", -- 1712 - 0x6b0  :  143 - 0x8f -- Background 0xd6
    "11101111", -- 1713 - 0x6b1  :  239 - 0xef
    "11000000", -- 1714 - 0x6b2  :  192 - 0xc0
    "11110000", -- 1715 - 0x6b3  :  240 - 0xf0
    "11100000", -- 1716 - 0x6b4  :  224 - 0xe0
    "11111111", -- 1717 - 0x6b5  :  255 - 0xff
    "11111111", -- 1718 - 0x6b6  :  255 - 0xff
    "11111111", -- 1719 - 0x6b7  :  255 - 0xff
    "11111111", -- 1720 - 0x6b8  :  255 - 0xff -- Background 0xd7
    "11111111", -- 1721 - 0x6b9  :  255 - 0xff
    "00000000", -- 1722 - 0x6ba  :    0 - 0x0
    "00000000", -- 1723 - 0x6bb  :    0 - 0x0
    "00000000", -- 1724 - 0x6bc  :    0 - 0x0
    "11111111", -- 1725 - 0x6bd  :  255 - 0xff
    "11111111", -- 1726 - 0x6be  :  255 - 0xff
    "11111111", -- 1727 - 0x6bf  :  255 - 0xff
    "11000011", -- 1728 - 0x6c0  :  195 - 0xc3 -- Background 0xd8
    "11111111", -- 1729 - 0x6c1  :  255 - 0xff
    "00000000", -- 1730 - 0x6c2  :    0 - 0x0
    "00000000", -- 1731 - 0x6c3  :    0 - 0x0
    "00000000", -- 1732 - 0x6c4  :    0 - 0x0
    "11111111", -- 1733 - 0x6c5  :  255 - 0xff
    "11111111", -- 1734 - 0x6c6  :  255 - 0xff
    "11111111", -- 1735 - 0x6c7  :  255 - 0xff
    "00000011", -- 1736 - 0x6c8  :    3 - 0x3 -- Background 0xd9
    "10000001", -- 1737 - 0x6c9  :  129 - 0x81
    "00000000", -- 1738 - 0x6ca  :    0 - 0x0
    "00000000", -- 1739 - 0x6cb  :    0 - 0x0
    "00000011", -- 1740 - 0x6cc  :    3 - 0x3
    "11111111", -- 1741 - 0x6cd  :  255 - 0xff
    "11111111", -- 1742 - 0x6ce  :  255 - 0xff
    "11111111", -- 1743 - 0x6cf  :  255 - 0xff
    "11111111", -- 1744 - 0x6d0  :  255 - 0xff -- Background 0xda
    "11111111", -- 1745 - 0x6d1  :  255 - 0xff
    "01111110", -- 1746 - 0x6d2  :  126 - 0x7e
    "00000000", -- 1747 - 0x6d3  :    0 - 0x0
    "00000000", -- 1748 - 0x6d4  :    0 - 0x0
    "11100000", -- 1749 - 0x6d5  :  224 - 0xe0
    "11111111", -- 1750 - 0x6d6  :  255 - 0xff
    "11111111", -- 1751 - 0x6d7  :  255 - 0xff
    "01100001", -- 1752 - 0x6d8  :   97 - 0x61 -- Background 0xdb
    "11000011", -- 1753 - 0x6d9  :  195 - 0xc3
    "00000111", -- 1754 - 0x6da  :    7 - 0x7
    "00001111", -- 1755 - 0x6db  :   15 - 0xf
    "00011111", -- 1756 - 0x6dc  :   31 - 0x1f
    "01111111", -- 1757 - 0x6dd  :  127 - 0x7f
    "11111111", -- 1758 - 0x6de  :  255 - 0xff
    "11111111", -- 1759 - 0x6df  :  255 - 0xff
    "00011111", -- 1760 - 0x6e0  :   31 - 0x1f -- Background 0xdc
    "11011111", -- 1761 - 0x6e1  :  223 - 0xdf
    "11000000", -- 1762 - 0x6e2  :  192 - 0xc0
    "11110000", -- 1763 - 0x6e3  :  240 - 0xf0
    "11110000", -- 1764 - 0x6e4  :  240 - 0xf0
    "11111111", -- 1765 - 0x6e5  :  255 - 0xff
    "11111111", -- 1766 - 0x6e6  :  255 - 0xff
    "11111111", -- 1767 - 0x6e7  :  255 - 0xff
    "10000100", -- 1768 - 0x6e8  :  132 - 0x84 -- Background 0xdd
    "11111100", -- 1769 - 0x6e9  :  252 - 0xfc
    "00000000", -- 1770 - 0x6ea  :    0 - 0x0
    "00000000", -- 1771 - 0x6eb  :    0 - 0x0
    "00000000", -- 1772 - 0x6ec  :    0 - 0x0
    "11111111", -- 1773 - 0x6ed  :  255 - 0xff
    "11111111", -- 1774 - 0x6ee  :  255 - 0xff
    "11111111", -- 1775 - 0x6ef  :  255 - 0xff
    "01111111", -- 1776 - 0x6f0  :  127 - 0x7f -- Background 0xde
    "01111111", -- 1777 - 0x6f1  :  127 - 0x7f
    "00000000", -- 1778 - 0x6f2  :    0 - 0x0
    "00000000", -- 1779 - 0x6f3  :    0 - 0x0
    "00000000", -- 1780 - 0x6f4  :    0 - 0x0
    "11111111", -- 1781 - 0x6f5  :  255 - 0xff
    "11111111", -- 1782 - 0x6f6  :  255 - 0xff
    "11111111", -- 1783 - 0x6f7  :  255 - 0xff
    "11111100", -- 1784 - 0x6f8  :  252 - 0xfc -- Background 0xdf
    "11111111", -- 1785 - 0x6f9  :  255 - 0xff
    "00000000", -- 1786 - 0x6fa  :    0 - 0x0
    "00000000", -- 1787 - 0x6fb  :    0 - 0x0
    "00000000", -- 1788 - 0x6fc  :    0 - 0x0
    "11111111", -- 1789 - 0x6fd  :  255 - 0xff
    "11111111", -- 1790 - 0x6fe  :  255 - 0xff
    "11111111", -- 1791 - 0x6ff  :  255 - 0xff
    "00110000", -- 1792 - 0x700  :   48 - 0x30 -- Background 0xe0
    "11110000", -- 1793 - 0x701  :  240 - 0xf0
    "00000000", -- 1794 - 0x702  :    0 - 0x0
    "00000000", -- 1795 - 0x703  :    0 - 0x0
    "00000000", -- 1796 - 0x704  :    0 - 0x0
    "11111111", -- 1797 - 0x705  :  255 - 0xff
    "11111111", -- 1798 - 0x706  :  255 - 0xff
    "11111111", -- 1799 - 0x707  :  255 - 0xff
    "11111111", -- 1800 - 0x708  :  255 - 0xff -- Background 0xe1
    "11111111", -- 1801 - 0x709  :  255 - 0xff
    "00000000", -- 1802 - 0x70a  :    0 - 0x0
    "00000000", -- 1803 - 0x70b  :    0 - 0x0
    "00000000", -- 1804 - 0x70c  :    0 - 0x0
    "11111111", -- 1805 - 0x70d  :  255 - 0xff
    "11111111", -- 1806 - 0x70e  :  255 - 0xff
    "11111111", -- 1807 - 0x70f  :  255 - 0xff
    "11100001", -- 1808 - 0x710  :  225 - 0xe1 -- Background 0xe2
    "11111111", -- 1809 - 0x711  :  255 - 0xff
    "00000000", -- 1810 - 0x712  :    0 - 0x0
    "00000000", -- 1811 - 0x713  :    0 - 0x0
    "00000000", -- 1812 - 0x714  :    0 - 0x0
    "11111111", -- 1813 - 0x715  :  255 - 0xff
    "11111111", -- 1814 - 0x716  :  255 - 0xff
    "11111111", -- 1815 - 0x717  :  255 - 0xff
    "00011111", -- 1816 - 0x718  :   31 - 0x1f -- Background 0xe3
    "00011111", -- 1817 - 0x719  :   31 - 0x1f
    "00011111", -- 1818 - 0x71a  :   31 - 0x1f
    "00011111", -- 1819 - 0x71b  :   31 - 0x1f
    "00011111", -- 1820 - 0x71c  :   31 - 0x1f
    "11111111", -- 1821 - 0x71d  :  255 - 0xff
    "11111111", -- 1822 - 0x71e  :  255 - 0xff
    "11111111", -- 1823 - 0x71f  :  255 - 0xff
    "00000000", -- 1824 - 0x720  :    0 - 0x0 -- Background 0xe4
    "00011111", -- 1825 - 0x721  :   31 - 0x1f
    "00111111", -- 1826 - 0x722  :   63 - 0x3f
    "01111000", -- 1827 - 0x723  :  120 - 0x78
    "01110111", -- 1828 - 0x724  :  119 - 0x77
    "01101111", -- 1829 - 0x725  :  111 - 0x6f
    "01101111", -- 1830 - 0x726  :  111 - 0x6f
    "01101111", -- 1831 - 0x727  :  111 - 0x6f
    "00000000", -- 1832 - 0x728  :    0 - 0x0 -- Background 0xe5
    "11111000", -- 1833 - 0x729  :  248 - 0xf8
    "11111100", -- 1834 - 0x72a  :  252 - 0xfc
    "00011110", -- 1835 - 0x72b  :   30 - 0x1e
    "11101110", -- 1836 - 0x72c  :  238 - 0xee
    "11110110", -- 1837 - 0x72d  :  246 - 0xf6
    "11110110", -- 1838 - 0x72e  :  246 - 0xf6
    "11110110", -- 1839 - 0x72f  :  246 - 0xf6
    "11110110", -- 1840 - 0x730  :  246 - 0xf6 -- Background 0xe6
    "11110110", -- 1841 - 0x731  :  246 - 0xf6
    "11110110", -- 1842 - 0x732  :  246 - 0xf6
    "11101110", -- 1843 - 0x733  :  238 - 0xee
    "00011110", -- 1844 - 0x734  :   30 - 0x1e
    "11111100", -- 1845 - 0x735  :  252 - 0xfc
    "11111000", -- 1846 - 0x736  :  248 - 0xf8
    "00000000", -- 1847 - 0x737  :    0 - 0x0
    "01101111", -- 1848 - 0x738  :  111 - 0x6f -- Background 0xe7
    "01101111", -- 1849 - 0x739  :  111 - 0x6f
    "01101111", -- 1850 - 0x73a  :  111 - 0x6f
    "01110111", -- 1851 - 0x73b  :  119 - 0x77
    "01111000", -- 1852 - 0x73c  :  120 - 0x78
    "00111111", -- 1853 - 0x73d  :   63 - 0x3f
    "00011111", -- 1854 - 0x73e  :   31 - 0x1f
    "00000000", -- 1855 - 0x73f  :    0 - 0x0
    "00000000", -- 1856 - 0x740  :    0 - 0x0 -- Background 0xe8
    "11111111", -- 1857 - 0x741  :  255 - 0xff
    "11111111", -- 1858 - 0x742  :  255 - 0xff
    "00000000", -- 1859 - 0x743  :    0 - 0x0
    "11111111", -- 1860 - 0x744  :  255 - 0xff
    "11111111", -- 1861 - 0x745  :  255 - 0xff
    "11111111", -- 1862 - 0x746  :  255 - 0xff
    "11111111", -- 1863 - 0x747  :  255 - 0xff
    "11110110", -- 1864 - 0x748  :  246 - 0xf6 -- Background 0xe9
    "11110110", -- 1865 - 0x749  :  246 - 0xf6
    "11110110", -- 1866 - 0x74a  :  246 - 0xf6
    "11110110", -- 1867 - 0x74b  :  246 - 0xf6
    "11110110", -- 1868 - 0x74c  :  246 - 0xf6
    "11110110", -- 1869 - 0x74d  :  246 - 0xf6
    "11110110", -- 1870 - 0x74e  :  246 - 0xf6
    "11110110", -- 1871 - 0x74f  :  246 - 0xf6
    "11111111", -- 1872 - 0x750  :  255 - 0xff -- Background 0xea
    "11111111", -- 1873 - 0x751  :  255 - 0xff
    "11111111", -- 1874 - 0x752  :  255 - 0xff
    "11111111", -- 1875 - 0x753  :  255 - 0xff
    "00000000", -- 1876 - 0x754  :    0 - 0x0
    "11111111", -- 1877 - 0x755  :  255 - 0xff
    "11111111", -- 1878 - 0x756  :  255 - 0xff
    "00000000", -- 1879 - 0x757  :    0 - 0x0
    "01101111", -- 1880 - 0x758  :  111 - 0x6f -- Background 0xeb
    "01101111", -- 1881 - 0x759  :  111 - 0x6f
    "01101111", -- 1882 - 0x75a  :  111 - 0x6f
    "01101111", -- 1883 - 0x75b  :  111 - 0x6f
    "01101111", -- 1884 - 0x75c  :  111 - 0x6f
    "01101111", -- 1885 - 0x75d  :  111 - 0x6f
    "01101111", -- 1886 - 0x75e  :  111 - 0x6f
    "01101111", -- 1887 - 0x75f  :  111 - 0x6f
    "00000000", -- 1888 - 0x760  :    0 - 0x0 -- Background 0xec
    "00000000", -- 1889 - 0x761  :    0 - 0x0
    "00000000", -- 1890 - 0x762  :    0 - 0x0
    "00000000", -- 1891 - 0x763  :    0 - 0x0
    "00000000", -- 1892 - 0x764  :    0 - 0x0
    "00000000", -- 1893 - 0x765  :    0 - 0x0
    "00000000", -- 1894 - 0x766  :    0 - 0x0
    "00000000", -- 1895 - 0x767  :    0 - 0x0
    "00000000", -- 1896 - 0x768  :    0 - 0x0 -- Background 0xed
    "00000000", -- 1897 - 0x769  :    0 - 0x0
    "00000000", -- 1898 - 0x76a  :    0 - 0x0
    "00000000", -- 1899 - 0x76b  :    0 - 0x0
    "00000000", -- 1900 - 0x76c  :    0 - 0x0
    "00000000", -- 1901 - 0x76d  :    0 - 0x0
    "00000000", -- 1902 - 0x76e  :    0 - 0x0
    "00000000", -- 1903 - 0x76f  :    0 - 0x0
    "00000000", -- 1904 - 0x770  :    0 - 0x0 -- Background 0xee
    "00000000", -- 1905 - 0x771  :    0 - 0x0
    "00000000", -- 1906 - 0x772  :    0 - 0x0
    "00000000", -- 1907 - 0x773  :    0 - 0x0
    "00000000", -- 1908 - 0x774  :    0 - 0x0
    "00000000", -- 1909 - 0x775  :    0 - 0x0
    "00000000", -- 1910 - 0x776  :    0 - 0x0
    "00000000", -- 1911 - 0x777  :    0 - 0x0
    "00000000", -- 1912 - 0x778  :    0 - 0x0 -- Background 0xef
    "00000000", -- 1913 - 0x779  :    0 - 0x0
    "00000000", -- 1914 - 0x77a  :    0 - 0x0
    "00000000", -- 1915 - 0x77b  :    0 - 0x0
    "00000000", -- 1916 - 0x77c  :    0 - 0x0
    "00000000", -- 1917 - 0x77d  :    0 - 0x0
    "00000000", -- 1918 - 0x77e  :    0 - 0x0
    "00000000", -- 1919 - 0x77f  :    0 - 0x0
    "11111111", -- 1920 - 0x780  :  255 - 0xff -- Background 0xf0
    "11111111", -- 1921 - 0x781  :  255 - 0xff
    "11111111", -- 1922 - 0x782  :  255 - 0xff
    "11111111", -- 1923 - 0x783  :  255 - 0xff
    "11111111", -- 1924 - 0x784  :  255 - 0xff
    "11111111", -- 1925 - 0x785  :  255 - 0xff
    "11111111", -- 1926 - 0x786  :  255 - 0xff
    "11111111", -- 1927 - 0x787  :  255 - 0xff
    "11111111", -- 1928 - 0x788  :  255 - 0xff -- Background 0xf1
    "11111111", -- 1929 - 0x789  :  255 - 0xff
    "11111111", -- 1930 - 0x78a  :  255 - 0xff
    "11111111", -- 1931 - 0x78b  :  255 - 0xff
    "11111111", -- 1932 - 0x78c  :  255 - 0xff
    "11111111", -- 1933 - 0x78d  :  255 - 0xff
    "11111111", -- 1934 - 0x78e  :  255 - 0xff
    "11111111", -- 1935 - 0x78f  :  255 - 0xff
    "11111111", -- 1936 - 0x790  :  255 - 0xff -- Background 0xf2
    "11111111", -- 1937 - 0x791  :  255 - 0xff
    "11111111", -- 1938 - 0x792  :  255 - 0xff
    "11111111", -- 1939 - 0x793  :  255 - 0xff
    "11111111", -- 1940 - 0x794  :  255 - 0xff
    "11111111", -- 1941 - 0x795  :  255 - 0xff
    "11111111", -- 1942 - 0x796  :  255 - 0xff
    "11111111", -- 1943 - 0x797  :  255 - 0xff
    "11111111", -- 1944 - 0x798  :  255 - 0xff -- Background 0xf3
    "11111111", -- 1945 - 0x799  :  255 - 0xff
    "11111111", -- 1946 - 0x79a  :  255 - 0xff
    "11111111", -- 1947 - 0x79b  :  255 - 0xff
    "11111111", -- 1948 - 0x79c  :  255 - 0xff
    "11111111", -- 1949 - 0x79d  :  255 - 0xff
    "11111111", -- 1950 - 0x79e  :  255 - 0xff
    "11111111", -- 1951 - 0x79f  :  255 - 0xff
    "11111111", -- 1952 - 0x7a0  :  255 - 0xff -- Background 0xf4
    "11111111", -- 1953 - 0x7a1  :  255 - 0xff
    "11111111", -- 1954 - 0x7a2  :  255 - 0xff
    "11111111", -- 1955 - 0x7a3  :  255 - 0xff
    "11111111", -- 1956 - 0x7a4  :  255 - 0xff
    "11111111", -- 1957 - 0x7a5  :  255 - 0xff
    "11111111", -- 1958 - 0x7a6  :  255 - 0xff
    "11111111", -- 1959 - 0x7a7  :  255 - 0xff
    "11111111", -- 1960 - 0x7a8  :  255 - 0xff -- Background 0xf5
    "11111111", -- 1961 - 0x7a9  :  255 - 0xff
    "11111111", -- 1962 - 0x7aa  :  255 - 0xff
    "11111111", -- 1963 - 0x7ab  :  255 - 0xff
    "11111111", -- 1964 - 0x7ac  :  255 - 0xff
    "11111111", -- 1965 - 0x7ad  :  255 - 0xff
    "11111111", -- 1966 - 0x7ae  :  255 - 0xff
    "11111111", -- 1967 - 0x7af  :  255 - 0xff
    "11111111", -- 1968 - 0x7b0  :  255 - 0xff -- Background 0xf6
    "11111111", -- 1969 - 0x7b1  :  255 - 0xff
    "11111111", -- 1970 - 0x7b2  :  255 - 0xff
    "11111111", -- 1971 - 0x7b3  :  255 - 0xff
    "11111111", -- 1972 - 0x7b4  :  255 - 0xff
    "11111111", -- 1973 - 0x7b5  :  255 - 0xff
    "11111111", -- 1974 - 0x7b6  :  255 - 0xff
    "11111111", -- 1975 - 0x7b7  :  255 - 0xff
    "11111111", -- 1976 - 0x7b8  :  255 - 0xff -- Background 0xf7
    "11111111", -- 1977 - 0x7b9  :  255 - 0xff
    "11111111", -- 1978 - 0x7ba  :  255 - 0xff
    "11111111", -- 1979 - 0x7bb  :  255 - 0xff
    "11111111", -- 1980 - 0x7bc  :  255 - 0xff
    "11111111", -- 1981 - 0x7bd  :  255 - 0xff
    "11111111", -- 1982 - 0x7be  :  255 - 0xff
    "11111111", -- 1983 - 0x7bf  :  255 - 0xff
    "11111111", -- 1984 - 0x7c0  :  255 - 0xff -- Background 0xf8
    "11111111", -- 1985 - 0x7c1  :  255 - 0xff
    "11111111", -- 1986 - 0x7c2  :  255 - 0xff
    "11111111", -- 1987 - 0x7c3  :  255 - 0xff
    "11111111", -- 1988 - 0x7c4  :  255 - 0xff
    "11111111", -- 1989 - 0x7c5  :  255 - 0xff
    "11111111", -- 1990 - 0x7c6  :  255 - 0xff
    "11111111", -- 1991 - 0x7c7  :  255 - 0xff
    "11111111", -- 1992 - 0x7c8  :  255 - 0xff -- Background 0xf9
    "11111111", -- 1993 - 0x7c9  :  255 - 0xff
    "11111111", -- 1994 - 0x7ca  :  255 - 0xff
    "11111111", -- 1995 - 0x7cb  :  255 - 0xff
    "11111111", -- 1996 - 0x7cc  :  255 - 0xff
    "11111111", -- 1997 - 0x7cd  :  255 - 0xff
    "11111111", -- 1998 - 0x7ce  :  255 - 0xff
    "11111111", -- 1999 - 0x7cf  :  255 - 0xff
    "11111111", -- 2000 - 0x7d0  :  255 - 0xff -- Background 0xfa
    "11111111", -- 2001 - 0x7d1  :  255 - 0xff
    "11111111", -- 2002 - 0x7d2  :  255 - 0xff
    "11111111", -- 2003 - 0x7d3  :  255 - 0xff
    "11111111", -- 2004 - 0x7d4  :  255 - 0xff
    "11111111", -- 2005 - 0x7d5  :  255 - 0xff
    "11111111", -- 2006 - 0x7d6  :  255 - 0xff
    "11111111", -- 2007 - 0x7d7  :  255 - 0xff
    "11111111", -- 2008 - 0x7d8  :  255 - 0xff -- Background 0xfb
    "11111111", -- 2009 - 0x7d9  :  255 - 0xff
    "11111111", -- 2010 - 0x7da  :  255 - 0xff
    "11111111", -- 2011 - 0x7db  :  255 - 0xff
    "11111111", -- 2012 - 0x7dc  :  255 - 0xff
    "11111111", -- 2013 - 0x7dd  :  255 - 0xff
    "11111111", -- 2014 - 0x7de  :  255 - 0xff
    "11111111", -- 2015 - 0x7df  :  255 - 0xff
    "11111111", -- 2016 - 0x7e0  :  255 - 0xff -- Background 0xfc
    "11111111", -- 2017 - 0x7e1  :  255 - 0xff
    "11111111", -- 2018 - 0x7e2  :  255 - 0xff
    "11111111", -- 2019 - 0x7e3  :  255 - 0xff
    "11111111", -- 2020 - 0x7e4  :  255 - 0xff
    "11111111", -- 2021 - 0x7e5  :  255 - 0xff
    "11111111", -- 2022 - 0x7e6  :  255 - 0xff
    "11111111", -- 2023 - 0x7e7  :  255 - 0xff
    "11111111", -- 2024 - 0x7e8  :  255 - 0xff -- Background 0xfd
    "11111111", -- 2025 - 0x7e9  :  255 - 0xff
    "11111111", -- 2026 - 0x7ea  :  255 - 0xff
    "11111111", -- 2027 - 0x7eb  :  255 - 0xff
    "11111111", -- 2028 - 0x7ec  :  255 - 0xff
    "11111111", -- 2029 - 0x7ed  :  255 - 0xff
    "11111111", -- 2030 - 0x7ee  :  255 - 0xff
    "11111111", -- 2031 - 0x7ef  :  255 - 0xff
    "11111111", -- 2032 - 0x7f0  :  255 - 0xff -- Background 0xfe
    "11111111", -- 2033 - 0x7f1  :  255 - 0xff
    "11111111", -- 2034 - 0x7f2  :  255 - 0xff
    "11111111", -- 2035 - 0x7f3  :  255 - 0xff
    "11111111", -- 2036 - 0x7f4  :  255 - 0xff
    "11111111", -- 2037 - 0x7f5  :  255 - 0xff
    "11111111", -- 2038 - 0x7f6  :  255 - 0xff
    "11111111", -- 2039 - 0x7f7  :  255 - 0xff
    "11111111", -- 2040 - 0x7f8  :  255 - 0xff -- Background 0xff
    "11111111", -- 2041 - 0x7f9  :  255 - 0xff
    "11111111", -- 2042 - 0x7fa  :  255 - 0xff
    "11111111", -- 2043 - 0x7fb  :  255 - 0xff
    "11111111", -- 2044 - 0x7fc  :  255 - 0xff
    "11111111", -- 2045 - 0x7fd  :  255 - 0xff
    "11111111", -- 2046 - 0x7fe  :  255 - 0xff
    "11111111"  -- 2047 - 0x7ff  :  255 - 0xff
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
