------- ROM creada automaticamente por ppm2rom -----------
------- Felipe Machado -----------------------------------
------- Departamento de Tecnologia Electronica -----------
------- Universidad Rey Juan Carlos ----------------------
------- http://gtebim.es ---------------------------------
----------------------------------------------------------
--------Datos de la imagen -------------------------------
--- Fichero original    : laberinto_40x30.pbm 
--- Filas    : 30 
--- Columnas : 40 
--- Color    :  Blanco y negro. 2 niveles (1 bit)



------ Puertos -------------------------------------------
-- Entradas ----------------------------------------------
--    clk  :  senal de reloj
--    addr :  direccion de la memoria
-- Salidas  ----------------------------------------------
--    dout :  dato de 40 bits de la direccion addr (un ciclo despues)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM1b_1f_laberinto_40x30 is
  port (
    clk  : in  std_logic;   -- reloj
    addr : in  std_logic_vector(5-1 downto 0);
    dout : out std_logic_vector(40-1 downto 0) 
  );
end ROM1b_1f_laberinto_40x30;


architecture BEHAVIORAL of ROM1b_1f_laberinto_40x30 is
  signal addr_int  : natural range 0 to 2**5-1;
  type memostruct is array (natural range<>) of std_logic_vector(40-1 downto 0);
  constant filaimg : memostruct := (
       "0000000010000000001000000000000100000000",
       "0111111111111111111111110001111111111110",
       "0100000010000000010000011011000000100010",
       "0101111011111111111000010001011111111010",
       "0100000010000000001101111111110010101010",
       "0101111111111011111111001001010110101010",
       "0100100000010001001001101101010000111010",
       "1111111111111111101111000101011111100011",
       "0100000100000100100001111101010001111110",
       "0101110101111110101100001001000001001010",
       "0100000100010000101111111111111111101010",
       "0111111111010111111000001100000010101010",
       "0100100100010010001011111111111010101110",
       "0100100111111110101011111111111010101000",
       "1101111110000000101000000000000010101010",
       "0101000011101111101111111111111110101111",
       "0100011110100000101000000000000010100010",
       "0111110010111110001111111011111110111110",
       "0101010010000011111000001010000010001000",
       "0101011111111010001011101110111011111100",
       "0101000001000010101000000100000010000110",
       "0101111101111110101111111111111111110010",
       "1100001001001000101000011011000010010111",
       "0111111111101011101011010001011010010100",
       "0100000100001000101011010101011010010100",
       "0101001111111110101011010001011010010100",
       "0101111000000010001011011111011010010110",
       "0101000000111111111000010001000010010010",
       "0111111111100000011111111111111111111110",
       "0000000010000000001000000000000100000000"
        );

begin

  addr_int <= TO_INTEGER(unsigned(addr));

  P_ROM: process (clk)
  begin
    if clk'event and clk='1' then
      dout <= filaimg(addr_int);
    end if;
  end process;

end BEHAVIORAL;

