//-   Sprites Pattern table COLOR PLANE 0
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
//- Autcmatically generated verilog ROM from a NES memory file----


//-  Original memory dump file name: pacman_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_PTABLE_PACMAN_SPR_PLN0
  (
     input     clk,   // clock
     input      [11-1:0] addr,  //2048 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Sprite pattern Table COLOR PLANE 0
      11'h0: dout <= 8'b00000000; //    0 :   0 - 0x0 -- Sprite 0x0
      11'h1: dout <= 8'b00000011; //    1 :   3 - 0x3
      11'h2: dout <= 8'b00001111; //    2 :  15 - 0xf
      11'h3: dout <= 8'b00011111; //    3 :  31 - 0x1f
      11'h4: dout <= 8'b00111111; //    4 :  63 - 0x3f
      11'h5: dout <= 8'b00111111; //    5 :  63 - 0x3f
      11'h6: dout <= 8'b01111111; //    6 : 127 - 0x7f
      11'h7: dout <= 8'b01111111; //    7 : 127 - 0x7f
      11'h8: dout <= 8'b00000000; //    8 :   0 - 0x0 -- Sprite 0x1
      11'h9: dout <= 8'b11000000; //    9 : 192 - 0xc0
      11'hA: dout <= 8'b11110000; //   10 : 240 - 0xf0
      11'hB: dout <= 8'b11111000; //   11 : 248 - 0xf8
      11'hC: dout <= 8'b11111000; //   12 : 248 - 0xf8
      11'hD: dout <= 8'b11111100; //   13 : 252 - 0xfc
      11'hE: dout <= 8'b11111100; //   14 : 252 - 0xfc
      11'hF: dout <= 8'b11111100; //   15 : 252 - 0xfc
      11'h10: dout <= 8'b00000000; //   16 :   0 - 0x0 -- Sprite 0x2
      11'h11: dout <= 8'b00000111; //   17 :   7 - 0x7
      11'h12: dout <= 8'b00011111; //   18 :  31 - 0x1f
      11'h13: dout <= 8'b00111111; //   19 :  63 - 0x3f
      11'h14: dout <= 8'b00111111; //   20 :  63 - 0x3f
      11'h15: dout <= 8'b00001111; //   21 :  15 - 0xf
      11'h16: dout <= 8'b00000011; //   22 :   3 - 0x3
      11'h17: dout <= 8'b00000000; //   23 :   0 - 0x0
      11'h18: dout <= 8'b00000000; //   24 :   0 - 0x0 -- Sprite 0x3
      11'h19: dout <= 8'b00000000; //   25 :   0 - 0x0
      11'h1A: dout <= 8'b00000111; //   26 :   7 - 0x7
      11'h1B: dout <= 8'b00011111; //   27 :  31 - 0x1f
      11'h1C: dout <= 8'b00111111; //   28 :  63 - 0x3f
      11'h1D: dout <= 8'b00111111; //   29 :  63 - 0x3f
      11'h1E: dout <= 8'b01111111; //   30 : 127 - 0x7f
      11'h1F: dout <= 8'b01111111; //   31 : 127 - 0x7f
      11'h20: dout <= 8'b01111110; //   32 : 126 - 0x7e -- Sprite 0x4
      11'h21: dout <= 8'b01111110; //   33 : 126 - 0x7e
      11'h22: dout <= 8'b01111100; //   34 : 124 - 0x7c
      11'h23: dout <= 8'b00111100; //   35 :  60 - 0x3c
      11'h24: dout <= 8'b00111000; //   36 :  56 - 0x38
      11'h25: dout <= 8'b00011000; //   37 :  24 - 0x18
      11'h26: dout <= 8'b00000000; //   38 :   0 - 0x0
      11'h27: dout <= 8'b00000000; //   39 :   0 - 0x0
      11'h28: dout <= 8'b00000000; //   40 :   0 - 0x0 -- Sprite 0x5
      11'h29: dout <= 8'b11000000; //   41 : 192 - 0xc0
      11'h2A: dout <= 8'b11110000; //   42 : 240 - 0xf0
      11'h2B: dout <= 8'b11111000; //   43 : 248 - 0xf8
      11'h2C: dout <= 8'b11111000; //   44 : 248 - 0xf8
      11'h2D: dout <= 8'b11111100; //   45 : 252 - 0xfc
      11'h2E: dout <= 8'b01111100; //   46 : 124 - 0x7c
      11'h2F: dout <= 8'b00111100; //   47 :  60 - 0x3c
      11'h30: dout <= 8'b00000000; //   48 :   0 - 0x0 -- Sprite 0x6
      11'h31: dout <= 8'b00000111; //   49 :   7 - 0x7
      11'h32: dout <= 8'b00000111; //   50 :   7 - 0x7
      11'h33: dout <= 8'b00000011; //   51 :   3 - 0x3
      11'h34: dout <= 8'b00000001; //   52 :   1 - 0x1
      11'h35: dout <= 8'b00000000; //   53 :   0 - 0x0
      11'h36: dout <= 8'b00000000; //   54 :   0 - 0x0
      11'h37: dout <= 8'b00000000; //   55 :   0 - 0x0
      11'h38: dout <= 8'b00000000; //   56 :   0 - 0x0 -- Sprite 0x7
      11'h39: dout <= 8'b00000000; //   57 :   0 - 0x0
      11'h3A: dout <= 8'b00000111; //   58 :   7 - 0x7
      11'h3B: dout <= 8'b00011111; //   59 :  31 - 0x1f
      11'h3C: dout <= 8'b00111111; //   60 :  63 - 0x3f
      11'h3D: dout <= 8'b00111111; //   61 :  63 - 0x3f
      11'h3E: dout <= 8'b01111110; //   62 : 126 - 0x7e
      11'h3F: dout <= 8'b01111100; //   63 : 124 - 0x7c
      11'h40: dout <= 8'b01111000; //   64 : 120 - 0x78 -- Sprite 0x8
      11'h41: dout <= 8'b01110000; //   65 : 112 - 0x70
      11'h42: dout <= 8'b01100000; //   66 :  96 - 0x60
      11'h43: dout <= 8'b00000000; //   67 :   0 - 0x0
      11'h44: dout <= 8'b00000000; //   68 :   0 - 0x0
      11'h45: dout <= 8'b00000000; //   69 :   0 - 0x0
      11'h46: dout <= 8'b00000000; //   70 :   0 - 0x0
      11'h47: dout <= 8'b00000000; //   71 :   0 - 0x0
      11'h48: dout <= 8'b00000000; //   72 :   0 - 0x0 -- Sprite 0x9
      11'h49: dout <= 8'b00000000; //   73 :   0 - 0x0
      11'h4A: dout <= 8'b00000000; //   74 :   0 - 0x0
      11'h4B: dout <= 8'b00000000; //   75 :   0 - 0x0
      11'h4C: dout <= 8'b00000000; //   76 :   0 - 0x0
      11'h4D: dout <= 8'b01000000; //   77 :  64 - 0x40
      11'h4E: dout <= 8'b11110000; //   78 : 240 - 0xf0
      11'h4F: dout <= 8'b11111000; //   79 : 248 - 0xf8
      11'h50: dout <= 8'b11111110; //   80 : 254 - 0xfe -- Sprite 0xa
      11'h51: dout <= 8'b01111111; //   81 : 127 - 0x7f
      11'h52: dout <= 8'b01111111; //   82 : 127 - 0x7f
      11'h53: dout <= 8'b00111111; //   83 :  63 - 0x3f
      11'h54: dout <= 8'b00001110; //   84 :  14 - 0xe
      11'h55: dout <= 8'b00000000; //   85 :   0 - 0x0
      11'h56: dout <= 8'b00000000; //   86 :   0 - 0x0
      11'h57: dout <= 8'b00000000; //   87 :   0 - 0x0
      11'h58: dout <= 8'b00000000; //   88 :   0 - 0x0 -- Sprite 0xb
      11'h59: dout <= 8'b00000000; //   89 :   0 - 0x0
      11'h5A: dout <= 8'b00000000; //   90 :   0 - 0x0
      11'h5B: dout <= 8'b00000000; //   91 :   0 - 0x0
      11'h5C: dout <= 8'b00000000; //   92 :   0 - 0x0
      11'h5D: dout <= 8'b00000000; //   93 :   0 - 0x0
      11'h5E: dout <= 8'b00000000; //   94 :   0 - 0x0
      11'h5F: dout <= 8'b11100000; //   95 : 224 - 0xe0
      11'h60: dout <= 8'b11111100; //   96 : 252 - 0xfc -- Sprite 0xc
      11'h61: dout <= 8'b11111111; //   97 : 255 - 0xff
      11'h62: dout <= 8'b01111111; //   98 : 127 - 0x7f
      11'h63: dout <= 8'b00111111; //   99 :  63 - 0x3f
      11'h64: dout <= 8'b00001110; //  100 :  14 - 0xe
      11'h65: dout <= 8'b00000000; //  101 :   0 - 0x0
      11'h66: dout <= 8'b00000000; //  102 :   0 - 0x0
      11'h67: dout <= 8'b00000000; //  103 :   0 - 0x0
      11'h68: dout <= 8'b11110000; //  104 : 240 - 0xf0 -- Sprite 0xd
      11'h69: dout <= 8'b11111111; //  105 : 255 - 0xff
      11'h6A: dout <= 8'b11111111; //  106 : 255 - 0xff
      11'h6B: dout <= 8'b01111111; //  107 : 127 - 0x7f
      11'h6C: dout <= 8'b00011110; //  108 :  30 - 0x1e
      11'h6D: dout <= 8'b00000000; //  109 :   0 - 0x0
      11'h6E: dout <= 8'b00000000; //  110 :   0 - 0x0
      11'h6F: dout <= 8'b00000000; //  111 :   0 - 0x0
      11'h70: dout <= 8'b00000000; //  112 :   0 - 0x0 -- Sprite 0xe
      11'h71: dout <= 8'b00001111; //  113 :  15 - 0xf
      11'h72: dout <= 8'b11111111; //  114 : 255 - 0xff
      11'h73: dout <= 8'b11111111; //  115 : 255 - 0xff
      11'h74: dout <= 8'b01111111; //  116 : 127 - 0x7f
      11'h75: dout <= 8'b00011110; //  117 :  30 - 0x1e
      11'h76: dout <= 8'b00000000; //  118 :   0 - 0x0
      11'h77: dout <= 8'b00000000; //  119 :   0 - 0x0
      11'h78: dout <= 8'b00000000; //  120 :   0 - 0x0 -- Sprite 0xf
      11'h79: dout <= 8'b00000011; //  121 :   3 - 0x3
      11'h7A: dout <= 8'b00001111; //  122 :  15 - 0xf
      11'h7B: dout <= 8'b01111111; //  123 : 127 - 0x7f
      11'h7C: dout <= 8'b11111111; //  124 : 255 - 0xff
      11'h7D: dout <= 8'b01111110; //  125 : 126 - 0x7e
      11'h7E: dout <= 8'b00011100; //  126 :  28 - 0x1c
      11'h7F: dout <= 8'b00000000; //  127 :   0 - 0x0
      11'h80: dout <= 8'b00000000; //  128 :   0 - 0x0 -- Sprite 0x10
      11'h81: dout <= 8'b00000001; //  129 :   1 - 0x1
      11'h82: dout <= 8'b00000011; //  130 :   3 - 0x3
      11'h83: dout <= 8'b00001111; //  131 :  15 - 0xf
      11'h84: dout <= 8'b00011111; //  132 :  31 - 0x1f
      11'h85: dout <= 8'b01111111; //  133 : 127 - 0x7f
      11'h86: dout <= 8'b01111110; //  134 : 126 - 0x7e
      11'h87: dout <= 8'b00111100; //  135 :  60 - 0x3c
      11'h88: dout <= 8'b00000000; //  136 :   0 - 0x0 -- Sprite 0x11
      11'h89: dout <= 8'b00000001; //  137 :   1 - 0x1
      11'h8A: dout <= 8'b00000011; //  138 :   3 - 0x3
      11'h8B: dout <= 8'b00000111; //  139 :   7 - 0x7
      11'h8C: dout <= 8'b00000111; //  140 :   7 - 0x7
      11'h8D: dout <= 8'b00001111; //  141 :  15 - 0xf
      11'h8E: dout <= 8'b00011111; //  142 :  31 - 0x1f
      11'h8F: dout <= 8'b00001110; //  143 :  14 - 0xe
      11'h90: dout <= 8'b00000000; //  144 :   0 - 0x0 -- Sprite 0x12
      11'h91: dout <= 8'b00000000; //  145 :   0 - 0x0
      11'h92: dout <= 8'b00000001; //  146 :   1 - 0x1
      11'h93: dout <= 8'b00000011; //  147 :   3 - 0x3
      11'h94: dout <= 8'b00000011; //  148 :   3 - 0x3
      11'h95: dout <= 8'b00000011; //  149 :   3 - 0x3
      11'h96: dout <= 8'b00000111; //  150 :   7 - 0x7
      11'h97: dout <= 8'b00000010; //  151 :   2 - 0x2
      11'h98: dout <= 8'b00000000; //  152 :   0 - 0x0 -- Sprite 0x13
      11'h99: dout <= 8'b00000000; //  153 :   0 - 0x0
      11'h9A: dout <= 8'b00000001; //  154 :   1 - 0x1
      11'h9B: dout <= 8'b00000001; //  155 :   1 - 0x1
      11'h9C: dout <= 8'b00000001; //  156 :   1 - 0x1
      11'h9D: dout <= 8'b00000001; //  157 :   1 - 0x1
      11'h9E: dout <= 8'b00000001; //  158 :   1 - 0x1
      11'h9F: dout <= 8'b00000001; //  159 :   1 - 0x1
      11'hA0: dout <= 8'b00000000; //  160 :   0 - 0x0 -- Sprite 0x14
      11'hA1: dout <= 8'b00000000; //  161 :   0 - 0x0
      11'hA2: dout <= 8'b00000000; //  162 :   0 - 0x0
      11'hA3: dout <= 8'b00000000; //  163 :   0 - 0x0
      11'hA4: dout <= 8'b00000000; //  164 :   0 - 0x0
      11'hA5: dout <= 8'b00000000; //  165 :   0 - 0x0
      11'hA6: dout <= 8'b00000100; //  166 :   4 - 0x4
      11'hA7: dout <= 8'b00000010; //  167 :   2 - 0x2
      11'hA8: dout <= 8'b00000000; //  168 :   0 - 0x0 -- Sprite 0x15
      11'hA9: dout <= 8'b00000000; //  169 :   0 - 0x0
      11'hAA: dout <= 8'b00000000; //  170 :   0 - 0x0
      11'hAB: dout <= 8'b00000000; //  171 :   0 - 0x0
      11'hAC: dout <= 8'b00000000; //  172 :   0 - 0x0
      11'hAD: dout <= 8'b00000000; //  173 :   0 - 0x0
      11'hAE: dout <= 8'b00100000; //  174 :  32 - 0x20
      11'hAF: dout <= 8'b01001000; //  175 :  72 - 0x48
      11'hB0: dout <= 8'b00010000; //  176 :  16 - 0x10 -- Sprite 0x16
      11'hB1: dout <= 8'b00001000; //  177 :   8 - 0x8
      11'hB2: dout <= 8'b00000000; //  178 :   0 - 0x0
      11'hB3: dout <= 8'b00110000; //  179 :  48 - 0x30
      11'hB4: dout <= 8'b00000000; //  180 :   0 - 0x0
      11'hB5: dout <= 8'b00001000; //  181 :   8 - 0x8
      11'hB6: dout <= 8'b00010010; //  182 :  18 - 0x12
      11'hB7: dout <= 8'b00000100; //  183 :   4 - 0x4
      11'hB8: dout <= 8'b00010000; //  184 :  16 - 0x10 -- Sprite 0x17
      11'hB9: dout <= 8'b00000000; //  185 :   0 - 0x0
      11'hBA: dout <= 8'b00001100; //  186 :  12 - 0xc
      11'hBB: dout <= 8'b00000000; //  187 :   0 - 0x0
      11'hBC: dout <= 8'b00010000; //  188 :  16 - 0x10
      11'hBD: dout <= 8'b00001000; //  189 :   8 - 0x8
      11'hBE: dout <= 8'b01000000; //  190 :  64 - 0x40
      11'hBF: dout <= 8'b00100000; //  191 :  32 - 0x20
      11'hC0: dout <= 8'b00000000; //  192 :   0 - 0x0 -- Sprite 0x18
      11'hC1: dout <= 8'b00000000; //  193 :   0 - 0x0
      11'hC2: dout <= 8'b00000011; //  194 :   3 - 0x3
      11'hC3: dout <= 8'b00000011; //  195 :   3 - 0x3
      11'hC4: dout <= 8'b00000001; //  196 :   1 - 0x1
      11'hC5: dout <= 8'b00100001; //  197 :  33 - 0x21
      11'hC6: dout <= 8'b00100001; //  198 :  33 - 0x21
      11'hC7: dout <= 8'b01110011; //  199 : 115 - 0x73
      11'hC8: dout <= 8'b01111111; //  200 : 127 - 0x7f -- Sprite 0x19
      11'hC9: dout <= 8'b01111111; //  201 : 127 - 0x7f
      11'hCA: dout <= 8'b01111111; //  202 : 127 - 0x7f
      11'hCB: dout <= 8'b01111111; //  203 : 127 - 0x7f
      11'hCC: dout <= 8'b01101110; //  204 : 110 - 0x6e
      11'hCD: dout <= 8'b01000110; //  205 :  70 - 0x46
      11'hCE: dout <= 8'b00000000; //  206 :   0 - 0x0
      11'hCF: dout <= 8'b00000000; //  207 :   0 - 0x0
      11'hD0: dout <= 8'b01111111; //  208 : 127 - 0x7f -- Sprite 0x1a
      11'hD1: dout <= 8'b01111111; //  209 : 127 - 0x7f
      11'hD2: dout <= 8'b01111111; //  210 : 127 - 0x7f
      11'hD3: dout <= 8'b01111111; //  211 : 127 - 0x7f
      11'hD4: dout <= 8'b01111011; //  212 : 123 - 0x7b
      11'hD5: dout <= 8'b00110001; //  213 :  49 - 0x31
      11'hD6: dout <= 8'b00000000; //  214 :   0 - 0x0
      11'hD7: dout <= 8'b00000000; //  215 :   0 - 0x0
      11'hD8: dout <= 8'b00000000; //  216 :   0 - 0x0 -- Sprite 0x1b
      11'hD9: dout <= 8'b00000011; //  217 :   3 - 0x3
      11'hDA: dout <= 8'b00001111; //  218 :  15 - 0xf
      11'hDB: dout <= 8'b00011111; //  219 :  31 - 0x1f
      11'hDC: dout <= 8'b00100111; //  220 :  39 - 0x27
      11'hDD: dout <= 8'b00000011; //  221 :   3 - 0x3
      11'hDE: dout <= 8'b00000011; //  222 :   3 - 0x3
      11'hDF: dout <= 8'b01000011; //  223 :  67 - 0x43
      11'hE0: dout <= 8'b00000000; //  224 :   0 - 0x0 -- Sprite 0x1c
      11'hE1: dout <= 8'b11000000; //  225 : 192 - 0xc0
      11'hE2: dout <= 8'b11110000; //  226 : 240 - 0xf0
      11'hE3: dout <= 8'b11111000; //  227 : 248 - 0xf8
      11'hE4: dout <= 8'b10011100; //  228 : 156 - 0x9c
      11'hE5: dout <= 8'b00001100; //  229 :  12 - 0xc
      11'hE6: dout <= 8'b00001100; //  230 :  12 - 0xc
      11'hE7: dout <= 8'b00001110; //  231 :  14 - 0xe
      11'hE8: dout <= 8'b01100111; //  232 : 103 - 0x67 -- Sprite 0x1d
      11'hE9: dout <= 8'b01111111; //  233 : 127 - 0x7f
      11'hEA: dout <= 8'b01111111; //  234 : 127 - 0x7f
      11'hEB: dout <= 8'b01111111; //  235 : 127 - 0x7f
      11'hEC: dout <= 8'b01101110; //  236 : 110 - 0x6e
      11'hED: dout <= 8'b01000110; //  237 :  70 - 0x46
      11'hEE: dout <= 8'b00000000; //  238 :   0 - 0x0
      11'hEF: dout <= 8'b00000000; //  239 :   0 - 0x0
      11'hF0: dout <= 8'b01100111; //  240 : 103 - 0x67 -- Sprite 0x1e
      11'hF1: dout <= 8'b01111111; //  241 : 127 - 0x7f
      11'hF2: dout <= 8'b01111111; //  242 : 127 - 0x7f
      11'hF3: dout <= 8'b01111111; //  243 : 127 - 0x7f
      11'hF4: dout <= 8'b01111011; //  244 : 123 - 0x7b
      11'hF5: dout <= 8'b00110001; //  245 :  49 - 0x31
      11'hF6: dout <= 8'b00000000; //  246 :   0 - 0x0
      11'hF7: dout <= 8'b00000000; //  247 :   0 - 0x0
      11'hF8: dout <= 8'b10011110; //  248 : 158 - 0x9e -- Sprite 0x1f
      11'hF9: dout <= 8'b11111110; //  249 : 254 - 0xfe
      11'hFA: dout <= 8'b11111110; //  250 : 254 - 0xfe
      11'hFB: dout <= 8'b11111110; //  251 : 254 - 0xfe
      11'hFC: dout <= 8'b01110110; //  252 : 118 - 0x76
      11'hFD: dout <= 8'b01100010; //  253 :  98 - 0x62
      11'hFE: dout <= 8'b00000000; //  254 :   0 - 0x0
      11'hFF: dout <= 8'b00000000; //  255 :   0 - 0x0
      11'h100: dout <= 8'b10011110; //  256 : 158 - 0x9e -- Sprite 0x20
      11'h101: dout <= 8'b11111110; //  257 : 254 - 0xfe
      11'h102: dout <= 8'b11111110; //  258 : 254 - 0xfe
      11'h103: dout <= 8'b11111110; //  259 : 254 - 0xfe
      11'h104: dout <= 8'b11011110; //  260 : 222 - 0xde
      11'h105: dout <= 8'b10001100; //  261 : 140 - 0x8c
      11'h106: dout <= 8'b00000000; //  262 :   0 - 0x0
      11'h107: dout <= 8'b00000000; //  263 :   0 - 0x0
      11'h108: dout <= 8'b00000000; //  264 :   0 - 0x0 -- Sprite 0x21
      11'h109: dout <= 8'b00000011; //  265 :   3 - 0x3
      11'h10A: dout <= 8'b00001111; //  266 :  15 - 0xf
      11'h10B: dout <= 8'b00011111; //  267 :  31 - 0x1f
      11'h10C: dout <= 8'b00111111; //  268 :  63 - 0x3f
      11'h10D: dout <= 8'b00110011; //  269 :  51 - 0x33
      11'h10E: dout <= 8'b00100001; //  270 :  33 - 0x21
      11'h10F: dout <= 8'b01100001; //  271 :  97 - 0x61
      11'h110: dout <= 8'b01100001; //  272 :  97 - 0x61 -- Sprite 0x22
      11'h111: dout <= 8'b01110011; //  273 : 115 - 0x73
      11'h112: dout <= 8'b01111111; //  274 : 127 - 0x7f
      11'h113: dout <= 8'b01111111; //  275 : 127 - 0x7f
      11'h114: dout <= 8'b01101110; //  276 : 110 - 0x6e
      11'h115: dout <= 8'b01000110; //  277 :  70 - 0x46
      11'h116: dout <= 8'b00000000; //  278 :   0 - 0x0
      11'h117: dout <= 8'b00000000; //  279 :   0 - 0x0
      11'h118: dout <= 8'b01100001; //  280 :  97 - 0x61 -- Sprite 0x23
      11'h119: dout <= 8'b01110011; //  281 : 115 - 0x73
      11'h11A: dout <= 8'b01111111; //  282 : 127 - 0x7f
      11'h11B: dout <= 8'b01111111; //  283 : 127 - 0x7f
      11'h11C: dout <= 8'b01110111; //  284 : 119 - 0x77
      11'h11D: dout <= 8'b00100011; //  285 :  35 - 0x23
      11'h11E: dout <= 8'b00000000; //  286 :   0 - 0x0
      11'h11F: dout <= 8'b00000000; //  287 :   0 - 0x0
      11'h120: dout <= 8'b00000000; //  288 :   0 - 0x0 -- Sprite 0x24
      11'h121: dout <= 8'b00000011; //  289 :   3 - 0x3
      11'h122: dout <= 8'b00001111; //  290 :  15 - 0xf
      11'h123: dout <= 8'b00011111; //  291 :  31 - 0x1f
      11'h124: dout <= 8'b00111111; //  292 :  63 - 0x3f
      11'h125: dout <= 8'b00111111; //  293 :  63 - 0x3f
      11'h126: dout <= 8'b00111111; //  294 :  63 - 0x3f
      11'h127: dout <= 8'b01111111; //  295 : 127 - 0x7f
      11'h128: dout <= 8'b01111111; //  296 : 127 - 0x7f -- Sprite 0x25
      11'h129: dout <= 8'b01111111; //  297 : 127 - 0x7f
      11'h12A: dout <= 8'b01111111; //  298 : 127 - 0x7f
      11'h12B: dout <= 8'b01111111; //  299 : 127 - 0x7f
      11'h12C: dout <= 8'b01101110; //  300 : 110 - 0x6e
      11'h12D: dout <= 8'b01000110; //  301 :  70 - 0x46
      11'h12E: dout <= 8'b00000000; //  302 :   0 - 0x0
      11'h12F: dout <= 8'b00000000; //  303 :   0 - 0x0
      11'h130: dout <= 8'b01111111; //  304 : 127 - 0x7f -- Sprite 0x26
      11'h131: dout <= 8'b01111111; //  305 : 127 - 0x7f
      11'h132: dout <= 8'b01111111; //  306 : 127 - 0x7f
      11'h133: dout <= 8'b01111111; //  307 : 127 - 0x7f
      11'h134: dout <= 8'b01111011; //  308 : 123 - 0x7b
      11'h135: dout <= 8'b00110001; //  309 :  49 - 0x31
      11'h136: dout <= 8'b00000000; //  310 :   0 - 0x0
      11'h137: dout <= 8'b00000000; //  311 :   0 - 0x0
      11'h138: dout <= 8'b00000000; //  312 :   0 - 0x0 -- Sprite 0x27
      11'h139: dout <= 8'b00000000; //  313 :   0 - 0x0
      11'h13A: dout <= 8'b00000000; //  314 :   0 - 0x0
      11'h13B: dout <= 8'b00000000; //  315 :   0 - 0x0
      11'h13C: dout <= 8'b00000000; //  316 :   0 - 0x0
      11'h13D: dout <= 8'b00000000; //  317 :   0 - 0x0
      11'h13E: dout <= 8'b00000000; //  318 :   0 - 0x0
      11'h13F: dout <= 8'b00000000; //  319 :   0 - 0x0
      11'h140: dout <= 8'b00000000; //  320 :   0 - 0x0 -- Sprite 0x28
      11'h141: dout <= 8'b00000000; //  321 :   0 - 0x0
      11'h142: dout <= 8'b00000000; //  322 :   0 - 0x0
      11'h143: dout <= 8'b00000000; //  323 :   0 - 0x0
      11'h144: dout <= 8'b00000000; //  324 :   0 - 0x0
      11'h145: dout <= 8'b00000000; //  325 :   0 - 0x0
      11'h146: dout <= 8'b00000000; //  326 :   0 - 0x0
      11'h147: dout <= 8'b00000000; //  327 :   0 - 0x0
      11'h148: dout <= 8'b00000000; //  328 :   0 - 0x0 -- Sprite 0x29
      11'h149: dout <= 8'b00000000; //  329 :   0 - 0x0
      11'h14A: dout <= 8'b00000000; //  330 :   0 - 0x0
      11'h14B: dout <= 8'b00000000; //  331 :   0 - 0x0
      11'h14C: dout <= 8'b00000000; //  332 :   0 - 0x0
      11'h14D: dout <= 8'b00000000; //  333 :   0 - 0x0
      11'h14E: dout <= 8'b00000000; //  334 :   0 - 0x0
      11'h14F: dout <= 8'b00000000; //  335 :   0 - 0x0
      11'h150: dout <= 8'b00000000; //  336 :   0 - 0x0 -- Sprite 0x2a
      11'h151: dout <= 8'b00000000; //  337 :   0 - 0x0
      11'h152: dout <= 8'b00000000; //  338 :   0 - 0x0
      11'h153: dout <= 8'b00000000; //  339 :   0 - 0x0
      11'h154: dout <= 8'b00000000; //  340 :   0 - 0x0
      11'h155: dout <= 8'b00000000; //  341 :   0 - 0x0
      11'h156: dout <= 8'b00000000; //  342 :   0 - 0x0
      11'h157: dout <= 8'b00000000; //  343 :   0 - 0x0
      11'h158: dout <= 8'b00000000; //  344 :   0 - 0x0 -- Sprite 0x2b
      11'h159: dout <= 8'b00000000; //  345 :   0 - 0x0
      11'h15A: dout <= 8'b00000000; //  346 :   0 - 0x0
      11'h15B: dout <= 8'b00000000; //  347 :   0 - 0x0
      11'h15C: dout <= 8'b00000000; //  348 :   0 - 0x0
      11'h15D: dout <= 8'b00000000; //  349 :   0 - 0x0
      11'h15E: dout <= 8'b00000000; //  350 :   0 - 0x0
      11'h15F: dout <= 8'b00000000; //  351 :   0 - 0x0
      11'h160: dout <= 8'b00000000; //  352 :   0 - 0x0 -- Sprite 0x2c
      11'h161: dout <= 8'b00000000; //  353 :   0 - 0x0
      11'h162: dout <= 8'b00000000; //  354 :   0 - 0x0
      11'h163: dout <= 8'b00000000; //  355 :   0 - 0x0
      11'h164: dout <= 8'b00000000; //  356 :   0 - 0x0
      11'h165: dout <= 8'b00000000; //  357 :   0 - 0x0
      11'h166: dout <= 8'b00000000; //  358 :   0 - 0x0
      11'h167: dout <= 8'b00000000; //  359 :   0 - 0x0
      11'h168: dout <= 8'b00000000; //  360 :   0 - 0x0 -- Sprite 0x2d
      11'h169: dout <= 8'b00000000; //  361 :   0 - 0x0
      11'h16A: dout <= 8'b00000000; //  362 :   0 - 0x0
      11'h16B: dout <= 8'b00000000; //  363 :   0 - 0x0
      11'h16C: dout <= 8'b00000000; //  364 :   0 - 0x0
      11'h16D: dout <= 8'b00000000; //  365 :   0 - 0x0
      11'h16E: dout <= 8'b00000000; //  366 :   0 - 0x0
      11'h16F: dout <= 8'b00000000; //  367 :   0 - 0x0
      11'h170: dout <= 8'b00000000; //  368 :   0 - 0x0 -- Sprite 0x2e
      11'h171: dout <= 8'b00000000; //  369 :   0 - 0x0
      11'h172: dout <= 8'b00000000; //  370 :   0 - 0x0
      11'h173: dout <= 8'b00000000; //  371 :   0 - 0x0
      11'h174: dout <= 8'b00000000; //  372 :   0 - 0x0
      11'h175: dout <= 8'b00000000; //  373 :   0 - 0x0
      11'h176: dout <= 8'b00000000; //  374 :   0 - 0x0
      11'h177: dout <= 8'b00000000; //  375 :   0 - 0x0
      11'h178: dout <= 8'b00000000; //  376 :   0 - 0x0 -- Sprite 0x2f
      11'h179: dout <= 8'b00000000; //  377 :   0 - 0x0
      11'h17A: dout <= 8'b00000000; //  378 :   0 - 0x0
      11'h17B: dout <= 8'b00000000; //  379 :   0 - 0x0
      11'h17C: dout <= 8'b00000000; //  380 :   0 - 0x0
      11'h17D: dout <= 8'b00000000; //  381 :   0 - 0x0
      11'h17E: dout <= 8'b00000000; //  382 :   0 - 0x0
      11'h17F: dout <= 8'b00000000; //  383 :   0 - 0x0
      11'h180: dout <= 8'b00000000; //  384 :   0 - 0x0 -- Sprite 0x30
      11'h181: dout <= 8'b00000000; //  385 :   0 - 0x0
      11'h182: dout <= 8'b00000000; //  386 :   0 - 0x0
      11'h183: dout <= 8'b00000000; //  387 :   0 - 0x0
      11'h184: dout <= 8'b00000000; //  388 :   0 - 0x0
      11'h185: dout <= 8'b00000000; //  389 :   0 - 0x0
      11'h186: dout <= 8'b00000000; //  390 :   0 - 0x0
      11'h187: dout <= 8'b00000000; //  391 :   0 - 0x0
      11'h188: dout <= 8'b00000000; //  392 :   0 - 0x0 -- Sprite 0x31
      11'h189: dout <= 8'b00000000; //  393 :   0 - 0x0
      11'h18A: dout <= 8'b00000000; //  394 :   0 - 0x0
      11'h18B: dout <= 8'b00000000; //  395 :   0 - 0x0
      11'h18C: dout <= 8'b00000000; //  396 :   0 - 0x0
      11'h18D: dout <= 8'b00000000; //  397 :   0 - 0x0
      11'h18E: dout <= 8'b00000000; //  398 :   0 - 0x0
      11'h18F: dout <= 8'b00000000; //  399 :   0 - 0x0
      11'h190: dout <= 8'b00000000; //  400 :   0 - 0x0 -- Sprite 0x32
      11'h191: dout <= 8'b00000000; //  401 :   0 - 0x0
      11'h192: dout <= 8'b00000000; //  402 :   0 - 0x0
      11'h193: dout <= 8'b00000000; //  403 :   0 - 0x0
      11'h194: dout <= 8'b00000000; //  404 :   0 - 0x0
      11'h195: dout <= 8'b00000000; //  405 :   0 - 0x0
      11'h196: dout <= 8'b00000000; //  406 :   0 - 0x0
      11'h197: dout <= 8'b00000000; //  407 :   0 - 0x0
      11'h198: dout <= 8'b00000000; //  408 :   0 - 0x0 -- Sprite 0x33
      11'h199: dout <= 8'b00000000; //  409 :   0 - 0x0
      11'h19A: dout <= 8'b00000000; //  410 :   0 - 0x0
      11'h19B: dout <= 8'b00000000; //  411 :   0 - 0x0
      11'h19C: dout <= 8'b00000000; //  412 :   0 - 0x0
      11'h19D: dout <= 8'b00000000; //  413 :   0 - 0x0
      11'h19E: dout <= 8'b00000000; //  414 :   0 - 0x0
      11'h19F: dout <= 8'b00000000; //  415 :   0 - 0x0
      11'h1A0: dout <= 8'b00000000; //  416 :   0 - 0x0 -- Sprite 0x34
      11'h1A1: dout <= 8'b00000000; //  417 :   0 - 0x0
      11'h1A2: dout <= 8'b00000000; //  418 :   0 - 0x0
      11'h1A3: dout <= 8'b00000000; //  419 :   0 - 0x0
      11'h1A4: dout <= 8'b00000000; //  420 :   0 - 0x0
      11'h1A5: dout <= 8'b00000000; //  421 :   0 - 0x0
      11'h1A6: dout <= 8'b00000000; //  422 :   0 - 0x0
      11'h1A7: dout <= 8'b00000000; //  423 :   0 - 0x0
      11'h1A8: dout <= 8'b00000000; //  424 :   0 - 0x0 -- Sprite 0x35
      11'h1A9: dout <= 8'b00000000; //  425 :   0 - 0x0
      11'h1AA: dout <= 8'b00000000; //  426 :   0 - 0x0
      11'h1AB: dout <= 8'b00000000; //  427 :   0 - 0x0
      11'h1AC: dout <= 8'b00000000; //  428 :   0 - 0x0
      11'h1AD: dout <= 8'b00000000; //  429 :   0 - 0x0
      11'h1AE: dout <= 8'b00000000; //  430 :   0 - 0x0
      11'h1AF: dout <= 8'b00000000; //  431 :   0 - 0x0
      11'h1B0: dout <= 8'b00000000; //  432 :   0 - 0x0 -- Sprite 0x36
      11'h1B1: dout <= 8'b00000000; //  433 :   0 - 0x0
      11'h1B2: dout <= 8'b00000000; //  434 :   0 - 0x0
      11'h1B3: dout <= 8'b00000000; //  435 :   0 - 0x0
      11'h1B4: dout <= 8'b00000000; //  436 :   0 - 0x0
      11'h1B5: dout <= 8'b00000000; //  437 :   0 - 0x0
      11'h1B6: dout <= 8'b00000000; //  438 :   0 - 0x0
      11'h1B7: dout <= 8'b00000000; //  439 :   0 - 0x0
      11'h1B8: dout <= 8'b00000000; //  440 :   0 - 0x0 -- Sprite 0x37
      11'h1B9: dout <= 8'b00000000; //  441 :   0 - 0x0
      11'h1BA: dout <= 8'b00000000; //  442 :   0 - 0x0
      11'h1BB: dout <= 8'b00000000; //  443 :   0 - 0x0
      11'h1BC: dout <= 8'b00000000; //  444 :   0 - 0x0
      11'h1BD: dout <= 8'b00000000; //  445 :   0 - 0x0
      11'h1BE: dout <= 8'b00000000; //  446 :   0 - 0x0
      11'h1BF: dout <= 8'b00000000; //  447 :   0 - 0x0
      11'h1C0: dout <= 8'b00000000; //  448 :   0 - 0x0 -- Sprite 0x38
      11'h1C1: dout <= 8'b00000000; //  449 :   0 - 0x0
      11'h1C2: dout <= 8'b00000000; //  450 :   0 - 0x0
      11'h1C3: dout <= 8'b00000000; //  451 :   0 - 0x0
      11'h1C4: dout <= 8'b00000000; //  452 :   0 - 0x0
      11'h1C5: dout <= 8'b00000000; //  453 :   0 - 0x0
      11'h1C6: dout <= 8'b00000000; //  454 :   0 - 0x0
      11'h1C7: dout <= 8'b00000000; //  455 :   0 - 0x0
      11'h1C8: dout <= 8'b00000000; //  456 :   0 - 0x0 -- Sprite 0x39
      11'h1C9: dout <= 8'b00000000; //  457 :   0 - 0x0
      11'h1CA: dout <= 8'b00000000; //  458 :   0 - 0x0
      11'h1CB: dout <= 8'b00000000; //  459 :   0 - 0x0
      11'h1CC: dout <= 8'b00000000; //  460 :   0 - 0x0
      11'h1CD: dout <= 8'b00000000; //  461 :   0 - 0x0
      11'h1CE: dout <= 8'b00000000; //  462 :   0 - 0x0
      11'h1CF: dout <= 8'b00000000; //  463 :   0 - 0x0
      11'h1D0: dout <= 8'b00000000; //  464 :   0 - 0x0 -- Sprite 0x3a
      11'h1D1: dout <= 8'b00000000; //  465 :   0 - 0x0
      11'h1D2: dout <= 8'b00000000; //  466 :   0 - 0x0
      11'h1D3: dout <= 8'b00000000; //  467 :   0 - 0x0
      11'h1D4: dout <= 8'b00000000; //  468 :   0 - 0x0
      11'h1D5: dout <= 8'b00000000; //  469 :   0 - 0x0
      11'h1D6: dout <= 8'b00000000; //  470 :   0 - 0x0
      11'h1D7: dout <= 8'b00000000; //  471 :   0 - 0x0
      11'h1D8: dout <= 8'b00000000; //  472 :   0 - 0x0 -- Sprite 0x3b
      11'h1D9: dout <= 8'b00000000; //  473 :   0 - 0x0
      11'h1DA: dout <= 8'b00000000; //  474 :   0 - 0x0
      11'h1DB: dout <= 8'b00000000; //  475 :   0 - 0x0
      11'h1DC: dout <= 8'b00000000; //  476 :   0 - 0x0
      11'h1DD: dout <= 8'b00000000; //  477 :   0 - 0x0
      11'h1DE: dout <= 8'b00000000; //  478 :   0 - 0x0
      11'h1DF: dout <= 8'b00000000; //  479 :   0 - 0x0
      11'h1E0: dout <= 8'b00000000; //  480 :   0 - 0x0 -- Sprite 0x3c
      11'h1E1: dout <= 8'b00000000; //  481 :   0 - 0x0
      11'h1E2: dout <= 8'b00000000; //  482 :   0 - 0x0
      11'h1E3: dout <= 8'b00000000; //  483 :   0 - 0x0
      11'h1E4: dout <= 8'b00000000; //  484 :   0 - 0x0
      11'h1E5: dout <= 8'b00000000; //  485 :   0 - 0x0
      11'h1E6: dout <= 8'b00000000; //  486 :   0 - 0x0
      11'h1E7: dout <= 8'b00000000; //  487 :   0 - 0x0
      11'h1E8: dout <= 8'b00000000; //  488 :   0 - 0x0 -- Sprite 0x3d
      11'h1E9: dout <= 8'b00000000; //  489 :   0 - 0x0
      11'h1EA: dout <= 8'b00000000; //  490 :   0 - 0x0
      11'h1EB: dout <= 8'b00000000; //  491 :   0 - 0x0
      11'h1EC: dout <= 8'b00000000; //  492 :   0 - 0x0
      11'h1ED: dout <= 8'b00000000; //  493 :   0 - 0x0
      11'h1EE: dout <= 8'b00000000; //  494 :   0 - 0x0
      11'h1EF: dout <= 8'b00000000; //  495 :   0 - 0x0
      11'h1F0: dout <= 8'b00000000; //  496 :   0 - 0x0 -- Sprite 0x3e
      11'h1F1: dout <= 8'b00000000; //  497 :   0 - 0x0
      11'h1F2: dout <= 8'b00000000; //  498 :   0 - 0x0
      11'h1F3: dout <= 8'b00000000; //  499 :   0 - 0x0
      11'h1F4: dout <= 8'b00000000; //  500 :   0 - 0x0
      11'h1F5: dout <= 8'b00000000; //  501 :   0 - 0x0
      11'h1F6: dout <= 8'b00000000; //  502 :   0 - 0x0
      11'h1F7: dout <= 8'b00000000; //  503 :   0 - 0x0
      11'h1F8: dout <= 8'b00000000; //  504 :   0 - 0x0 -- Sprite 0x3f
      11'h1F9: dout <= 8'b00000000; //  505 :   0 - 0x0
      11'h1FA: dout <= 8'b00000000; //  506 :   0 - 0x0
      11'h1FB: dout <= 8'b00000000; //  507 :   0 - 0x0
      11'h1FC: dout <= 8'b00000000; //  508 :   0 - 0x0
      11'h1FD: dout <= 8'b00000000; //  509 :   0 - 0x0
      11'h1FE: dout <= 8'b00000000; //  510 :   0 - 0x0
      11'h1FF: dout <= 8'b00000000; //  511 :   0 - 0x0
      11'h200: dout <= 8'b00000000; //  512 :   0 - 0x0 -- Sprite 0x40
      11'h201: dout <= 8'b00000000; //  513 :   0 - 0x0
      11'h202: dout <= 8'b00000000; //  514 :   0 - 0x0
      11'h203: dout <= 8'b00000000; //  515 :   0 - 0x0
      11'h204: dout <= 8'b00000000; //  516 :   0 - 0x0
      11'h205: dout <= 8'b00000000; //  517 :   0 - 0x0
      11'h206: dout <= 8'b00000000; //  518 :   0 - 0x0
      11'h207: dout <= 8'b00000000; //  519 :   0 - 0x0
      11'h208: dout <= 8'b00000000; //  520 :   0 - 0x0 -- Sprite 0x41
      11'h209: dout <= 8'b00000000; //  521 :   0 - 0x0
      11'h20A: dout <= 8'b00000000; //  522 :   0 - 0x0
      11'h20B: dout <= 8'b00000000; //  523 :   0 - 0x0
      11'h20C: dout <= 8'b00000000; //  524 :   0 - 0x0
      11'h20D: dout <= 8'b00000000; //  525 :   0 - 0x0
      11'h20E: dout <= 8'b00000000; //  526 :   0 - 0x0
      11'h20F: dout <= 8'b00000000; //  527 :   0 - 0x0
      11'h210: dout <= 8'b00000000; //  528 :   0 - 0x0 -- Sprite 0x42
      11'h211: dout <= 8'b00000000; //  529 :   0 - 0x0
      11'h212: dout <= 8'b00000000; //  530 :   0 - 0x0
      11'h213: dout <= 8'b00000000; //  531 :   0 - 0x0
      11'h214: dout <= 8'b00000000; //  532 :   0 - 0x0
      11'h215: dout <= 8'b00000000; //  533 :   0 - 0x0
      11'h216: dout <= 8'b00000000; //  534 :   0 - 0x0
      11'h217: dout <= 8'b00000000; //  535 :   0 - 0x0
      11'h218: dout <= 8'b00000000; //  536 :   0 - 0x0 -- Sprite 0x43
      11'h219: dout <= 8'b00000000; //  537 :   0 - 0x0
      11'h21A: dout <= 8'b00000000; //  538 :   0 - 0x0
      11'h21B: dout <= 8'b00000000; //  539 :   0 - 0x0
      11'h21C: dout <= 8'b00000000; //  540 :   0 - 0x0
      11'h21D: dout <= 8'b00000000; //  541 :   0 - 0x0
      11'h21E: dout <= 8'b00000000; //  542 :   0 - 0x0
      11'h21F: dout <= 8'b00000000; //  543 :   0 - 0x0
      11'h220: dout <= 8'b00000000; //  544 :   0 - 0x0 -- Sprite 0x44
      11'h221: dout <= 8'b00000000; //  545 :   0 - 0x0
      11'h222: dout <= 8'b00000000; //  546 :   0 - 0x0
      11'h223: dout <= 8'b00000000; //  547 :   0 - 0x0
      11'h224: dout <= 8'b00000000; //  548 :   0 - 0x0
      11'h225: dout <= 8'b00000000; //  549 :   0 - 0x0
      11'h226: dout <= 8'b00000000; //  550 :   0 - 0x0
      11'h227: dout <= 8'b00000000; //  551 :   0 - 0x0
      11'h228: dout <= 8'b00000000; //  552 :   0 - 0x0 -- Sprite 0x45
      11'h229: dout <= 8'b00000000; //  553 :   0 - 0x0
      11'h22A: dout <= 8'b00000000; //  554 :   0 - 0x0
      11'h22B: dout <= 8'b00000000; //  555 :   0 - 0x0
      11'h22C: dout <= 8'b00000000; //  556 :   0 - 0x0
      11'h22D: dout <= 8'b00000000; //  557 :   0 - 0x0
      11'h22E: dout <= 8'b00000000; //  558 :   0 - 0x0
      11'h22F: dout <= 8'b00000000; //  559 :   0 - 0x0
      11'h230: dout <= 8'b00000000; //  560 :   0 - 0x0 -- Sprite 0x46
      11'h231: dout <= 8'b00000000; //  561 :   0 - 0x0
      11'h232: dout <= 8'b00000000; //  562 :   0 - 0x0
      11'h233: dout <= 8'b00000000; //  563 :   0 - 0x0
      11'h234: dout <= 8'b00000000; //  564 :   0 - 0x0
      11'h235: dout <= 8'b00000000; //  565 :   0 - 0x0
      11'h236: dout <= 8'b00000000; //  566 :   0 - 0x0
      11'h237: dout <= 8'b00000000; //  567 :   0 - 0x0
      11'h238: dout <= 8'b00000000; //  568 :   0 - 0x0 -- Sprite 0x47
      11'h239: dout <= 8'b00000000; //  569 :   0 - 0x0
      11'h23A: dout <= 8'b00000000; //  570 :   0 - 0x0
      11'h23B: dout <= 8'b00000000; //  571 :   0 - 0x0
      11'h23C: dout <= 8'b00000000; //  572 :   0 - 0x0
      11'h23D: dout <= 8'b00000000; //  573 :   0 - 0x0
      11'h23E: dout <= 8'b00000000; //  574 :   0 - 0x0
      11'h23F: dout <= 8'b00000000; //  575 :   0 - 0x0
      11'h240: dout <= 8'b00000000; //  576 :   0 - 0x0 -- Sprite 0x48
      11'h241: dout <= 8'b00000000; //  577 :   0 - 0x0
      11'h242: dout <= 8'b00000000; //  578 :   0 - 0x0
      11'h243: dout <= 8'b00000000; //  579 :   0 - 0x0
      11'h244: dout <= 8'b00000000; //  580 :   0 - 0x0
      11'h245: dout <= 8'b00000000; //  581 :   0 - 0x0
      11'h246: dout <= 8'b00000000; //  582 :   0 - 0x0
      11'h247: dout <= 8'b00000000; //  583 :   0 - 0x0
      11'h248: dout <= 8'b00000000; //  584 :   0 - 0x0 -- Sprite 0x49
      11'h249: dout <= 8'b00000000; //  585 :   0 - 0x0
      11'h24A: dout <= 8'b00000000; //  586 :   0 - 0x0
      11'h24B: dout <= 8'b00000000; //  587 :   0 - 0x0
      11'h24C: dout <= 8'b00000000; //  588 :   0 - 0x0
      11'h24D: dout <= 8'b00000000; //  589 :   0 - 0x0
      11'h24E: dout <= 8'b00000000; //  590 :   0 - 0x0
      11'h24F: dout <= 8'b00000000; //  591 :   0 - 0x0
      11'h250: dout <= 8'b00000000; //  592 :   0 - 0x0 -- Sprite 0x4a
      11'h251: dout <= 8'b00000000; //  593 :   0 - 0x0
      11'h252: dout <= 8'b00000000; //  594 :   0 - 0x0
      11'h253: dout <= 8'b00000000; //  595 :   0 - 0x0
      11'h254: dout <= 8'b00000000; //  596 :   0 - 0x0
      11'h255: dout <= 8'b00000000; //  597 :   0 - 0x0
      11'h256: dout <= 8'b00000000; //  598 :   0 - 0x0
      11'h257: dout <= 8'b00000000; //  599 :   0 - 0x0
      11'h258: dout <= 8'b00000000; //  600 :   0 - 0x0 -- Sprite 0x4b
      11'h259: dout <= 8'b00000000; //  601 :   0 - 0x0
      11'h25A: dout <= 8'b00000000; //  602 :   0 - 0x0
      11'h25B: dout <= 8'b00000000; //  603 :   0 - 0x0
      11'h25C: dout <= 8'b00000000; //  604 :   0 - 0x0
      11'h25D: dout <= 8'b00000000; //  605 :   0 - 0x0
      11'h25E: dout <= 8'b00000000; //  606 :   0 - 0x0
      11'h25F: dout <= 8'b00000000; //  607 :   0 - 0x0
      11'h260: dout <= 8'b00000000; //  608 :   0 - 0x0 -- Sprite 0x4c
      11'h261: dout <= 8'b00000000; //  609 :   0 - 0x0
      11'h262: dout <= 8'b00000000; //  610 :   0 - 0x0
      11'h263: dout <= 8'b00000000; //  611 :   0 - 0x0
      11'h264: dout <= 8'b00000000; //  612 :   0 - 0x0
      11'h265: dout <= 8'b00000000; //  613 :   0 - 0x0
      11'h266: dout <= 8'b00000000; //  614 :   0 - 0x0
      11'h267: dout <= 8'b00000000; //  615 :   0 - 0x0
      11'h268: dout <= 8'b00000000; //  616 :   0 - 0x0 -- Sprite 0x4d
      11'h269: dout <= 8'b00000000; //  617 :   0 - 0x0
      11'h26A: dout <= 8'b00000000; //  618 :   0 - 0x0
      11'h26B: dout <= 8'b00000001; //  619 :   1 - 0x1
      11'h26C: dout <= 8'b00000011; //  620 :   3 - 0x3
      11'h26D: dout <= 8'b00000111; //  621 :   7 - 0x7
      11'h26E: dout <= 8'b00001111; //  622 :  15 - 0xf
      11'h26F: dout <= 8'b00011111; //  623 :  31 - 0x1f
      11'h270: dout <= 8'b00000000; //  624 :   0 - 0x0 -- Sprite 0x4e
      11'h271: dout <= 8'b00001111; //  625 :  15 - 0xf
      11'h272: dout <= 8'b01111111; //  626 : 127 - 0x7f
      11'h273: dout <= 8'b11111111; //  627 : 255 - 0xff
      11'h274: dout <= 8'b11111111; //  628 : 255 - 0xff
      11'h275: dout <= 8'b11111111; //  629 : 255 - 0xff
      11'h276: dout <= 8'b11111111; //  630 : 255 - 0xff
      11'h277: dout <= 8'b11111111; //  631 : 255 - 0xff
      11'h278: dout <= 8'b00011111; //  632 :  31 - 0x1f -- Sprite 0x4f
      11'h279: dout <= 8'b00111111; //  633 :  63 - 0x3f
      11'h27A: dout <= 8'b00111111; //  634 :  63 - 0x3f
      11'h27B: dout <= 8'b00111111; //  635 :  63 - 0x3f
      11'h27C: dout <= 8'b01111111; //  636 : 127 - 0x7f
      11'h27D: dout <= 8'b01111111; //  637 : 127 - 0x7f
      11'h27E: dout <= 8'b01111111; //  638 : 127 - 0x7f
      11'h27F: dout <= 8'b01111111; //  639 : 127 - 0x7f
      11'h280: dout <= 8'b11111111; //  640 : 255 - 0xff -- Sprite 0x50
      11'h281: dout <= 8'b11111111; //  641 : 255 - 0xff
      11'h282: dout <= 8'b11111111; //  642 : 255 - 0xff
      11'h283: dout <= 8'b11111111; //  643 : 255 - 0xff
      11'h284: dout <= 8'b11111111; //  644 : 255 - 0xff
      11'h285: dout <= 8'b11111111; //  645 : 255 - 0xff
      11'h286: dout <= 8'b11111111; //  646 : 255 - 0xff
      11'h287: dout <= 8'b11111111; //  647 : 255 - 0xff
      11'h288: dout <= 8'b11111111; //  648 : 255 - 0xff -- Sprite 0x51
      11'h289: dout <= 8'b11111111; //  649 : 255 - 0xff
      11'h28A: dout <= 8'b11111111; //  650 : 255 - 0xff
      11'h28B: dout <= 8'b11111111; //  651 : 255 - 0xff
      11'h28C: dout <= 8'b11111111; //  652 : 255 - 0xff
      11'h28D: dout <= 8'b11111111; //  653 : 255 - 0xff
      11'h28E: dout <= 8'b11111111; //  654 : 255 - 0xff
      11'h28F: dout <= 8'b11111110; //  655 : 254 - 0xfe
      11'h290: dout <= 8'b00000000; //  656 :   0 - 0x0 -- Sprite 0x52
      11'h291: dout <= 8'b00000000; //  657 :   0 - 0x0
      11'h292: dout <= 8'b00000000; //  658 :   0 - 0x0
      11'h293: dout <= 8'b10000000; //  659 : 128 - 0x80
      11'h294: dout <= 8'b11000000; //  660 : 192 - 0xc0
      11'h295: dout <= 8'b11100000; //  661 : 224 - 0xe0
      11'h296: dout <= 8'b11110000; //  662 : 240 - 0xf0
      11'h297: dout <= 8'b11110000; //  663 : 240 - 0xf0
      11'h298: dout <= 8'b11111111; //  664 : 255 - 0xff -- Sprite 0x53
      11'h299: dout <= 8'b11111111; //  665 : 255 - 0xff
      11'h29A: dout <= 8'b11111110; //  666 : 254 - 0xfe
      11'h29B: dout <= 8'b11111100; //  667 : 252 - 0xfc
      11'h29C: dout <= 8'b11110000; //  668 : 240 - 0xf0
      11'h29D: dout <= 8'b11100000; //  669 : 224 - 0xe0
      11'h29E: dout <= 8'b10000000; //  670 : 128 - 0x80
      11'h29F: dout <= 8'b00000000; //  671 :   0 - 0x0
      11'h2A0: dout <= 8'b11000000; //  672 : 192 - 0xc0 -- Sprite 0x54
      11'h2A1: dout <= 8'b10000000; //  673 : 128 - 0x80
      11'h2A2: dout <= 8'b00000000; //  674 :   0 - 0x0
      11'h2A3: dout <= 8'b00000000; //  675 :   0 - 0x0
      11'h2A4: dout <= 8'b00000000; //  676 :   0 - 0x0
      11'h2A5: dout <= 8'b00000000; //  677 :   0 - 0x0
      11'h2A6: dout <= 8'b00000000; //  678 :   0 - 0x0
      11'h2A7: dout <= 8'b00000000; //  679 :   0 - 0x0
      11'h2A8: dout <= 8'b00000000; //  680 :   0 - 0x0 -- Sprite 0x55
      11'h2A9: dout <= 8'b11110000; //  681 : 240 - 0xf0
      11'h2AA: dout <= 8'b11111110; //  682 : 254 - 0xfe
      11'h2AB: dout <= 8'b11111110; //  683 : 254 - 0xfe
      11'h2AC: dout <= 8'b11111110; //  684 : 254 - 0xfe
      11'h2AD: dout <= 8'b11111100; //  685 : 252 - 0xfc
      11'h2AE: dout <= 8'b11111000; //  686 : 248 - 0xf8
      11'h2AF: dout <= 8'b11111000; //  687 : 248 - 0xf8
      11'h2B0: dout <= 8'b11110000; //  688 : 240 - 0xf0 -- Sprite 0x56
      11'h2B1: dout <= 8'b11100000; //  689 : 224 - 0xe0
      11'h2B2: dout <= 8'b11100000; //  690 : 224 - 0xe0
      11'h2B3: dout <= 8'b11000000; //  691 : 192 - 0xc0
      11'h2B4: dout <= 8'b10000000; //  692 : 128 - 0x80
      11'h2B5: dout <= 8'b10000000; //  693 : 128 - 0x80
      11'h2B6: dout <= 8'b00000000; //  694 :   0 - 0x0
      11'h2B7: dout <= 8'b00000000; //  695 :   0 - 0x0
      11'h2B8: dout <= 8'b00000000; //  696 :   0 - 0x0 -- Sprite 0x57
      11'h2B9: dout <= 8'b00000000; //  697 :   0 - 0x0
      11'h2BA: dout <= 8'b00000000; //  698 :   0 - 0x0
      11'h2BB: dout <= 8'b00000000; //  699 :   0 - 0x0
      11'h2BC: dout <= 8'b00000000; //  700 :   0 - 0x0
      11'h2BD: dout <= 8'b00000000; //  701 :   0 - 0x0
      11'h2BE: dout <= 8'b00000000; //  702 :   0 - 0x0
      11'h2BF: dout <= 8'b00000100; //  703 :   4 - 0x4
      11'h2C0: dout <= 8'b00000110; //  704 :   6 - 0x6 -- Sprite 0x58
      11'h2C1: dout <= 8'b00000110; //  705 :   6 - 0x6
      11'h2C2: dout <= 8'b00000111; //  706 :   7 - 0x7
      11'h2C3: dout <= 8'b00000111; //  707 :   7 - 0x7
      11'h2C4: dout <= 8'b00000111; //  708 :   7 - 0x7
      11'h2C5: dout <= 8'b00000111; //  709 :   7 - 0x7
      11'h2C6: dout <= 8'b00000000; //  710 :   0 - 0x0
      11'h2C7: dout <= 8'b00000000; //  711 :   0 - 0x0
      11'h2C8: dout <= 8'b00000000; //  712 :   0 - 0x0 -- Sprite 0x59
      11'h2C9: dout <= 8'b00000000; //  713 :   0 - 0x0
      11'h2CA: dout <= 8'b00000000; //  714 :   0 - 0x0
      11'h2CB: dout <= 8'b00000000; //  715 :   0 - 0x0
      11'h2CC: dout <= 8'b00000000; //  716 :   0 - 0x0
      11'h2CD: dout <= 8'b00000000; //  717 :   0 - 0x0
      11'h2CE: dout <= 8'b00000000; //  718 :   0 - 0x0
      11'h2CF: dout <= 8'b00010000; //  719 :  16 - 0x10
      11'h2D0: dout <= 8'b00011100; //  720 :  28 - 0x1c -- Sprite 0x5a
      11'h2D1: dout <= 8'b00011110; //  721 :  30 - 0x1e
      11'h2D2: dout <= 8'b00011111; //  722 :  31 - 0x1f
      11'h2D3: dout <= 8'b00011111; //  723 :  31 - 0x1f
      11'h2D4: dout <= 8'b00011111; //  724 :  31 - 0x1f
      11'h2D5: dout <= 8'b00011111; //  725 :  31 - 0x1f
      11'h2D6: dout <= 8'b00000000; //  726 :   0 - 0x0
      11'h2D7: dout <= 8'b00000000; //  727 :   0 - 0x0
      11'h2D8: dout <= 8'b00000000; //  728 :   0 - 0x0 -- Sprite 0x5b
      11'h2D9: dout <= 8'b00000000; //  729 :   0 - 0x0
      11'h2DA: dout <= 8'b00000000; //  730 :   0 - 0x0
      11'h2DB: dout <= 8'b00000000; //  731 :   0 - 0x0
      11'h2DC: dout <= 8'b00000000; //  732 :   0 - 0x0
      11'h2DD: dout <= 8'b00000000; //  733 :   0 - 0x0
      11'h2DE: dout <= 8'b00000000; //  734 :   0 - 0x0
      11'h2DF: dout <= 8'b11000000; //  735 : 192 - 0xc0
      11'h2E0: dout <= 8'b11110000; //  736 : 240 - 0xf0 -- Sprite 0x5c
      11'h2E1: dout <= 8'b11111100; //  737 : 252 - 0xfc
      11'h2E2: dout <= 8'b11111111; //  738 : 255 - 0xff
      11'h2E3: dout <= 8'b11111111; //  739 : 255 - 0xff
      11'h2E4: dout <= 8'b11111111; //  740 : 255 - 0xff
      11'h2E5: dout <= 8'b11111111; //  741 : 255 - 0xff
      11'h2E6: dout <= 8'b00000000; //  742 :   0 - 0x0
      11'h2E7: dout <= 8'b00000000; //  743 :   0 - 0x0
      11'h2E8: dout <= 8'b00000000; //  744 :   0 - 0x0 -- Sprite 0x5d
      11'h2E9: dout <= 8'b00000000; //  745 :   0 - 0x0
      11'h2EA: dout <= 8'b00000001; //  746 :   1 - 0x1
      11'h2EB: dout <= 8'b00000011; //  747 :   3 - 0x3
      11'h2EC: dout <= 8'b00001111; //  748 :  15 - 0xf
      11'h2ED: dout <= 8'b00001111; //  749 :  15 - 0xf
      11'h2EE: dout <= 8'b00000000; //  750 :   0 - 0x0
      11'h2EF: dout <= 8'b00000000; //  751 :   0 - 0x0
      11'h2F0: dout <= 8'b11111100; //  752 : 252 - 0xfc -- Sprite 0x5e
      11'h2F1: dout <= 8'b11111100; //  753 : 252 - 0xfc
      11'h2F2: dout <= 8'b11111100; //  754 : 252 - 0xfc
      11'h2F3: dout <= 8'b11111100; //  755 : 252 - 0xfc
      11'h2F4: dout <= 8'b11111000; //  756 : 248 - 0xf8
      11'h2F5: dout <= 8'b11111100; //  757 : 252 - 0xfc
      11'h2F6: dout <= 8'b00111100; //  758 :  60 - 0x3c
      11'h2F7: dout <= 8'b00000000; //  759 :   0 - 0x0
      11'h2F8: dout <= 8'b00000100; //  760 :   4 - 0x4 -- Sprite 0x5f
      11'h2F9: dout <= 8'b00001100; //  761 :  12 - 0xc
      11'h2FA: dout <= 8'b00011100; //  762 :  28 - 0x1c
      11'h2FB: dout <= 8'b00001100; //  763 :  12 - 0xc
      11'h2FC: dout <= 8'b00011000; //  764 :  24 - 0x18
      11'h2FD: dout <= 8'b00111100; //  765 :  60 - 0x3c
      11'h2FE: dout <= 8'b00111100; //  766 :  60 - 0x3c
      11'h2FF: dout <= 8'b00000000; //  767 :   0 - 0x0
      11'h300: dout <= 8'b00000000; //  768 :   0 - 0x0 -- Sprite 0x60
      11'h301: dout <= 8'b00000011; //  769 :   3 - 0x3
      11'h302: dout <= 8'b00001111; //  770 :  15 - 0xf
      11'h303: dout <= 8'b00010011; //  771 :  19 - 0x13
      11'h304: dout <= 8'b00100001; //  772 :  33 - 0x21
      11'h305: dout <= 8'b00100001; //  773 :  33 - 0x21
      11'h306: dout <= 8'b00100001; //  774 :  33 - 0x21
      11'h307: dout <= 8'b01110011; //  775 : 115 - 0x73
      11'h308: dout <= 8'b00000000; //  776 :   0 - 0x0 -- Sprite 0x61
      11'h309: dout <= 8'b11000000; //  777 : 192 - 0xc0
      11'h30A: dout <= 8'b11110000; //  778 : 240 - 0xf0
      11'h30B: dout <= 8'b11001000; //  779 : 200 - 0xc8
      11'h30C: dout <= 8'b10000100; //  780 : 132 - 0x84
      11'h30D: dout <= 8'b10000100; //  781 : 132 - 0x84
      11'h30E: dout <= 8'b10000100; //  782 : 132 - 0x84
      11'h30F: dout <= 8'b11001110; //  783 : 206 - 0xce
      11'h310: dout <= 8'b10010100; //  784 : 148 - 0x94 -- Sprite 0x62
      11'h311: dout <= 8'b11101010; //  785 : 234 - 0xea
      11'h312: dout <= 8'b11011110; //  786 : 222 - 0xde
      11'h313: dout <= 8'b11101110; //  787 : 238 - 0xee
      11'h314: dout <= 8'b11011110; //  788 : 222 - 0xde
      11'h315: dout <= 8'b01100110; //  789 : 102 - 0x66
      11'h316: dout <= 8'b01000010; //  790 :  66 - 0x42
      11'h317: dout <= 8'b00000000; //  791 :   0 - 0x0
      11'h318: dout <= 8'b10010100; //  792 : 148 - 0x94 -- Sprite 0x63
      11'h319: dout <= 8'b11101010; //  793 : 234 - 0xea
      11'h31A: dout <= 8'b11011110; //  794 : 222 - 0xde
      11'h31B: dout <= 8'b11101110; //  795 : 238 - 0xee
      11'h31C: dout <= 8'b11011110; //  796 : 222 - 0xde
      11'h31D: dout <= 8'b11001110; //  797 : 206 - 0xce
      11'h31E: dout <= 8'b10001100; //  798 : 140 - 0x8c
      11'h31F: dout <= 8'b00000000; //  799 :   0 - 0x0
      11'h320: dout <= 8'b00000000; //  800 :   0 - 0x0 -- Sprite 0x64
      11'h321: dout <= 8'b00000000; //  801 :   0 - 0x0
      11'h322: dout <= 8'b00000000; //  802 :   0 - 0x0
      11'h323: dout <= 8'b00000000; //  803 :   0 - 0x0
      11'h324: dout <= 8'b00000000; //  804 :   0 - 0x0
      11'h325: dout <= 8'b00000000; //  805 :   0 - 0x0
      11'h326: dout <= 8'b00000000; //  806 :   0 - 0x0
      11'h327: dout <= 8'b00000001; //  807 :   1 - 0x1
      11'h328: dout <= 8'b00000000; //  808 :   0 - 0x0 -- Sprite 0x65
      11'h329: dout <= 8'b00000000; //  809 :   0 - 0x0
      11'h32A: dout <= 8'b00000000; //  810 :   0 - 0x0
      11'h32B: dout <= 8'b00000000; //  811 :   0 - 0x0
      11'h32C: dout <= 8'b00000000; //  812 :   0 - 0x0
      11'h32D: dout <= 8'b00110110; //  813 :  54 - 0x36
      11'h32E: dout <= 8'b00110110; //  814 :  54 - 0x36
      11'h32F: dout <= 8'b10010000; //  815 : 144 - 0x90
      11'h330: dout <= 8'b00000001; //  816 :   1 - 0x1 -- Sprite 0x66
      11'h331: dout <= 8'b00000011; //  817 :   3 - 0x3
      11'h332: dout <= 8'b00000111; //  818 :   7 - 0x7
      11'h333: dout <= 8'b00000111; //  819 :   7 - 0x7
      11'h334: dout <= 8'b00011111; //  820 :  31 - 0x1f
      11'h335: dout <= 8'b00011111; //  821 :  31 - 0x1f
      11'h336: dout <= 8'b00011100; //  822 :  28 - 0x1c
      11'h337: dout <= 8'b00000000; //  823 :   0 - 0x0
      11'h338: dout <= 8'b11111000; //  824 : 248 - 0xf8 -- Sprite 0x67
      11'h339: dout <= 8'b11111000; //  825 : 248 - 0xf8
      11'h33A: dout <= 8'b11111000; //  826 : 248 - 0xf8
      11'h33B: dout <= 8'b11111000; //  827 : 248 - 0xf8
      11'h33C: dout <= 8'b11111110; //  828 : 254 - 0xfe
      11'h33D: dout <= 8'b11111110; //  829 : 254 - 0xfe
      11'h33E: dout <= 8'b00001110; //  830 :  14 - 0xe
      11'h33F: dout <= 8'b00000000; //  831 :   0 - 0x0
      11'h340: dout <= 8'b00000111; //  832 :   7 - 0x7 -- Sprite 0x68
      11'h341: dout <= 8'b00001111; //  833 :  15 - 0xf
      11'h342: dout <= 8'b00011111; //  834 :  31 - 0x1f
      11'h343: dout <= 8'b00011111; //  835 :  31 - 0x1f
      11'h344: dout <= 8'b00111111; //  836 :  63 - 0x3f
      11'h345: dout <= 8'b00111111; //  837 :  63 - 0x3f
      11'h346: dout <= 8'b00111000; //  838 :  56 - 0x38
      11'h347: dout <= 8'b00000000; //  839 :   0 - 0x0
      11'h348: dout <= 8'b11111000; //  840 : 248 - 0xf8 -- Sprite 0x69
      11'h349: dout <= 8'b11110000; //  841 : 240 - 0xf0
      11'h34A: dout <= 8'b11110000; //  842 : 240 - 0xf0
      11'h34B: dout <= 8'b11100000; //  843 : 224 - 0xe0
      11'h34C: dout <= 8'b11111000; //  844 : 248 - 0xf8
      11'h34D: dout <= 8'b11111000; //  845 : 248 - 0xf8
      11'h34E: dout <= 8'b00111000; //  846 :  56 - 0x38
      11'h34F: dout <= 8'b00000000; //  847 :   0 - 0x0
      11'h350: dout <= 8'b00000000; //  848 :   0 - 0x0 -- Sprite 0x6a
      11'h351: dout <= 8'b00011111; //  849 :  31 - 0x1f
      11'h352: dout <= 8'b01111111; //  850 : 127 - 0x7f
      11'h353: dout <= 8'b00111111; //  851 :  63 - 0x3f
      11'h354: dout <= 8'b00001111; //  852 :  15 - 0xf
      11'h355: dout <= 8'b00000111; //  853 :   7 - 0x7
      11'h356: dout <= 8'b00000000; //  854 :   0 - 0x0
      11'h357: dout <= 8'b00000000; //  855 :   0 - 0x0
      11'h358: dout <= 8'b00000000; //  856 :   0 - 0x0 -- Sprite 0x6b
      11'h359: dout <= 8'b00000000; //  857 :   0 - 0x0
      11'h35A: dout <= 8'b11000000; //  858 : 192 - 0xc0
      11'h35B: dout <= 8'b11110000; //  859 : 240 - 0xf0
      11'h35C: dout <= 8'b11111000; //  860 : 248 - 0xf8
      11'h35D: dout <= 8'b11111000; //  861 : 248 - 0xf8
      11'h35E: dout <= 8'b11100000; //  862 : 224 - 0xe0
      11'h35F: dout <= 8'b00000000; //  863 :   0 - 0x0
      11'h360: dout <= 8'b00000000; //  864 :   0 - 0x0 -- Sprite 0x6c
      11'h361: dout <= 8'b00000000; //  865 :   0 - 0x0
      11'h362: dout <= 8'b00000000; //  866 :   0 - 0x0
      11'h363: dout <= 8'b00000000; //  867 :   0 - 0x0
      11'h364: dout <= 8'b00000000; //  868 :   0 - 0x0
      11'h365: dout <= 8'b00000000; //  869 :   0 - 0x0
      11'h366: dout <= 8'b00000000; //  870 :   0 - 0x0
      11'h367: dout <= 8'b00000000; //  871 :   0 - 0x0
      11'h368: dout <= 8'b00000000; //  872 :   0 - 0x0 -- Sprite 0x6d
      11'h369: dout <= 8'b00000000; //  873 :   0 - 0x0
      11'h36A: dout <= 8'b00000000; //  874 :   0 - 0x0
      11'h36B: dout <= 8'b00000000; //  875 :   0 - 0x0
      11'h36C: dout <= 8'b00000000; //  876 :   0 - 0x0
      11'h36D: dout <= 8'b00000000; //  877 :   0 - 0x0
      11'h36E: dout <= 8'b00000000; //  878 :   0 - 0x0
      11'h36F: dout <= 8'b00000000; //  879 :   0 - 0x0
      11'h370: dout <= 8'b00000000; //  880 :   0 - 0x0 -- Sprite 0x6e
      11'h371: dout <= 8'b00000000; //  881 :   0 - 0x0
      11'h372: dout <= 8'b00000000; //  882 :   0 - 0x0
      11'h373: dout <= 8'b00000000; //  883 :   0 - 0x0
      11'h374: dout <= 8'b00000000; //  884 :   0 - 0x0
      11'h375: dout <= 8'b00000000; //  885 :   0 - 0x0
      11'h376: dout <= 8'b00000000; //  886 :   0 - 0x0
      11'h377: dout <= 8'b00000000; //  887 :   0 - 0x0
      11'h378: dout <= 8'b00000000; //  888 :   0 - 0x0 -- Sprite 0x6f
      11'h379: dout <= 8'b00000000; //  889 :   0 - 0x0
      11'h37A: dout <= 8'b00000000; //  890 :   0 - 0x0
      11'h37B: dout <= 8'b00000000; //  891 :   0 - 0x0
      11'h37C: dout <= 8'b00000000; //  892 :   0 - 0x0
      11'h37D: dout <= 8'b00000000; //  893 :   0 - 0x0
      11'h37E: dout <= 8'b00000000; //  894 :   0 - 0x0
      11'h37F: dout <= 8'b00000000; //  895 :   0 - 0x0
      11'h380: dout <= 8'b11111111; //  896 : 255 - 0xff -- Sprite 0x70
      11'h381: dout <= 8'b11111111; //  897 : 255 - 0xff
      11'h382: dout <= 8'b11111111; //  898 : 255 - 0xff
      11'h383: dout <= 8'b11111111; //  899 : 255 - 0xff
      11'h384: dout <= 8'b11111111; //  900 : 255 - 0xff
      11'h385: dout <= 8'b11111111; //  901 : 255 - 0xff
      11'h386: dout <= 8'b11111111; //  902 : 255 - 0xff
      11'h387: dout <= 8'b11111111; //  903 : 255 - 0xff
      11'h388: dout <= 8'b11111111; //  904 : 255 - 0xff -- Sprite 0x71
      11'h389: dout <= 8'b11111111; //  905 : 255 - 0xff
      11'h38A: dout <= 8'b11111111; //  906 : 255 - 0xff
      11'h38B: dout <= 8'b11111111; //  907 : 255 - 0xff
      11'h38C: dout <= 8'b11111111; //  908 : 255 - 0xff
      11'h38D: dout <= 8'b11111111; //  909 : 255 - 0xff
      11'h38E: dout <= 8'b11111111; //  910 : 255 - 0xff
      11'h38F: dout <= 8'b11111111; //  911 : 255 - 0xff
      11'h390: dout <= 8'b11111111; //  912 : 255 - 0xff -- Sprite 0x72
      11'h391: dout <= 8'b11111111; //  913 : 255 - 0xff
      11'h392: dout <= 8'b11111111; //  914 : 255 - 0xff
      11'h393: dout <= 8'b11111111; //  915 : 255 - 0xff
      11'h394: dout <= 8'b11111111; //  916 : 255 - 0xff
      11'h395: dout <= 8'b11111111; //  917 : 255 - 0xff
      11'h396: dout <= 8'b11111111; //  918 : 255 - 0xff
      11'h397: dout <= 8'b11111111; //  919 : 255 - 0xff
      11'h398: dout <= 8'b11111111; //  920 : 255 - 0xff -- Sprite 0x73
      11'h399: dout <= 8'b11111111; //  921 : 255 - 0xff
      11'h39A: dout <= 8'b11111111; //  922 : 255 - 0xff
      11'h39B: dout <= 8'b11111111; //  923 : 255 - 0xff
      11'h39C: dout <= 8'b11111111; //  924 : 255 - 0xff
      11'h39D: dout <= 8'b11111111; //  925 : 255 - 0xff
      11'h39E: dout <= 8'b11111111; //  926 : 255 - 0xff
      11'h39F: dout <= 8'b11111111; //  927 : 255 - 0xff
      11'h3A0: dout <= 8'b11111111; //  928 : 255 - 0xff -- Sprite 0x74
      11'h3A1: dout <= 8'b11111111; //  929 : 255 - 0xff
      11'h3A2: dout <= 8'b11111111; //  930 : 255 - 0xff
      11'h3A3: dout <= 8'b11111111; //  931 : 255 - 0xff
      11'h3A4: dout <= 8'b11111111; //  932 : 255 - 0xff
      11'h3A5: dout <= 8'b11111111; //  933 : 255 - 0xff
      11'h3A6: dout <= 8'b11111111; //  934 : 255 - 0xff
      11'h3A7: dout <= 8'b11111111; //  935 : 255 - 0xff
      11'h3A8: dout <= 8'b11111111; //  936 : 255 - 0xff -- Sprite 0x75
      11'h3A9: dout <= 8'b11111111; //  937 : 255 - 0xff
      11'h3AA: dout <= 8'b11111111; //  938 : 255 - 0xff
      11'h3AB: dout <= 8'b11111111; //  939 : 255 - 0xff
      11'h3AC: dout <= 8'b11111111; //  940 : 255 - 0xff
      11'h3AD: dout <= 8'b11111111; //  941 : 255 - 0xff
      11'h3AE: dout <= 8'b11111111; //  942 : 255 - 0xff
      11'h3AF: dout <= 8'b11111111; //  943 : 255 - 0xff
      11'h3B0: dout <= 8'b11111111; //  944 : 255 - 0xff -- Sprite 0x76
      11'h3B1: dout <= 8'b11111111; //  945 : 255 - 0xff
      11'h3B2: dout <= 8'b11111111; //  946 : 255 - 0xff
      11'h3B3: dout <= 8'b11111111; //  947 : 255 - 0xff
      11'h3B4: dout <= 8'b11111111; //  948 : 255 - 0xff
      11'h3B5: dout <= 8'b11111111; //  949 : 255 - 0xff
      11'h3B6: dout <= 8'b11111111; //  950 : 255 - 0xff
      11'h3B7: dout <= 8'b11111111; //  951 : 255 - 0xff
      11'h3B8: dout <= 8'b11111111; //  952 : 255 - 0xff -- Sprite 0x77
      11'h3B9: dout <= 8'b11111111; //  953 : 255 - 0xff
      11'h3BA: dout <= 8'b11111111; //  954 : 255 - 0xff
      11'h3BB: dout <= 8'b11111111; //  955 : 255 - 0xff
      11'h3BC: dout <= 8'b11111111; //  956 : 255 - 0xff
      11'h3BD: dout <= 8'b11111111; //  957 : 255 - 0xff
      11'h3BE: dout <= 8'b11111111; //  958 : 255 - 0xff
      11'h3BF: dout <= 8'b11111111; //  959 : 255 - 0xff
      11'h3C0: dout <= 8'b11111111; //  960 : 255 - 0xff -- Sprite 0x78
      11'h3C1: dout <= 8'b11111111; //  961 : 255 - 0xff
      11'h3C2: dout <= 8'b11111111; //  962 : 255 - 0xff
      11'h3C3: dout <= 8'b11111111; //  963 : 255 - 0xff
      11'h3C4: dout <= 8'b11111111; //  964 : 255 - 0xff
      11'h3C5: dout <= 8'b11111111; //  965 : 255 - 0xff
      11'h3C6: dout <= 8'b11111111; //  966 : 255 - 0xff
      11'h3C7: dout <= 8'b11111111; //  967 : 255 - 0xff
      11'h3C8: dout <= 8'b11111111; //  968 : 255 - 0xff -- Sprite 0x79
      11'h3C9: dout <= 8'b11111111; //  969 : 255 - 0xff
      11'h3CA: dout <= 8'b11111111; //  970 : 255 - 0xff
      11'h3CB: dout <= 8'b11111111; //  971 : 255 - 0xff
      11'h3CC: dout <= 8'b11111111; //  972 : 255 - 0xff
      11'h3CD: dout <= 8'b11111111; //  973 : 255 - 0xff
      11'h3CE: dout <= 8'b11111111; //  974 : 255 - 0xff
      11'h3CF: dout <= 8'b11111111; //  975 : 255 - 0xff
      11'h3D0: dout <= 8'b11111111; //  976 : 255 - 0xff -- Sprite 0x7a
      11'h3D1: dout <= 8'b11111111; //  977 : 255 - 0xff
      11'h3D2: dout <= 8'b11111111; //  978 : 255 - 0xff
      11'h3D3: dout <= 8'b11111111; //  979 : 255 - 0xff
      11'h3D4: dout <= 8'b11111111; //  980 : 255 - 0xff
      11'h3D5: dout <= 8'b11111111; //  981 : 255 - 0xff
      11'h3D6: dout <= 8'b11111111; //  982 : 255 - 0xff
      11'h3D7: dout <= 8'b11111111; //  983 : 255 - 0xff
      11'h3D8: dout <= 8'b11111111; //  984 : 255 - 0xff -- Sprite 0x7b
      11'h3D9: dout <= 8'b11111111; //  985 : 255 - 0xff
      11'h3DA: dout <= 8'b11111111; //  986 : 255 - 0xff
      11'h3DB: dout <= 8'b11111111; //  987 : 255 - 0xff
      11'h3DC: dout <= 8'b11111111; //  988 : 255 - 0xff
      11'h3DD: dout <= 8'b11111111; //  989 : 255 - 0xff
      11'h3DE: dout <= 8'b11111111; //  990 : 255 - 0xff
      11'h3DF: dout <= 8'b11111111; //  991 : 255 - 0xff
      11'h3E0: dout <= 8'b11111111; //  992 : 255 - 0xff -- Sprite 0x7c
      11'h3E1: dout <= 8'b11111111; //  993 : 255 - 0xff
      11'h3E2: dout <= 8'b11111111; //  994 : 255 - 0xff
      11'h3E3: dout <= 8'b11111111; //  995 : 255 - 0xff
      11'h3E4: dout <= 8'b11111111; //  996 : 255 - 0xff
      11'h3E5: dout <= 8'b11111111; //  997 : 255 - 0xff
      11'h3E6: dout <= 8'b11111111; //  998 : 255 - 0xff
      11'h3E7: dout <= 8'b11111111; //  999 : 255 - 0xff
      11'h3E8: dout <= 8'b11111111; // 1000 : 255 - 0xff -- Sprite 0x7d
      11'h3E9: dout <= 8'b11111111; // 1001 : 255 - 0xff
      11'h3EA: dout <= 8'b11111111; // 1002 : 255 - 0xff
      11'h3EB: dout <= 8'b11111111; // 1003 : 255 - 0xff
      11'h3EC: dout <= 8'b11111111; // 1004 : 255 - 0xff
      11'h3ED: dout <= 8'b11111111; // 1005 : 255 - 0xff
      11'h3EE: dout <= 8'b11111111; // 1006 : 255 - 0xff
      11'h3EF: dout <= 8'b11111111; // 1007 : 255 - 0xff
      11'h3F0: dout <= 8'b11111111; // 1008 : 255 - 0xff -- Sprite 0x7e
      11'h3F1: dout <= 8'b11111111; // 1009 : 255 - 0xff
      11'h3F2: dout <= 8'b11111111; // 1010 : 255 - 0xff
      11'h3F3: dout <= 8'b11111111; // 1011 : 255 - 0xff
      11'h3F4: dout <= 8'b11111111; // 1012 : 255 - 0xff
      11'h3F5: dout <= 8'b11111111; // 1013 : 255 - 0xff
      11'h3F6: dout <= 8'b11111111; // 1014 : 255 - 0xff
      11'h3F7: dout <= 8'b11111111; // 1015 : 255 - 0xff
      11'h3F8: dout <= 8'b11111111; // 1016 : 255 - 0xff -- Sprite 0x7f
      11'h3F9: dout <= 8'b11111111; // 1017 : 255 - 0xff
      11'h3FA: dout <= 8'b11111111; // 1018 : 255 - 0xff
      11'h3FB: dout <= 8'b11111111; // 1019 : 255 - 0xff
      11'h3FC: dout <= 8'b11111111; // 1020 : 255 - 0xff
      11'h3FD: dout <= 8'b11111111; // 1021 : 255 - 0xff
      11'h3FE: dout <= 8'b11111111; // 1022 : 255 - 0xff
      11'h3FF: dout <= 8'b11111111; // 1023 : 255 - 0xff
      11'h400: dout <= 8'b11111111; // 1024 : 255 - 0xff -- Sprite 0x80
      11'h401: dout <= 8'b11111111; // 1025 : 255 - 0xff
      11'h402: dout <= 8'b11111111; // 1026 : 255 - 0xff
      11'h403: dout <= 8'b11111111; // 1027 : 255 - 0xff
      11'h404: dout <= 8'b11111111; // 1028 : 255 - 0xff
      11'h405: dout <= 8'b11111111; // 1029 : 255 - 0xff
      11'h406: dout <= 8'b11111111; // 1030 : 255 - 0xff
      11'h407: dout <= 8'b11111111; // 1031 : 255 - 0xff
      11'h408: dout <= 8'b11111111; // 1032 : 255 - 0xff -- Sprite 0x81
      11'h409: dout <= 8'b11111111; // 1033 : 255 - 0xff
      11'h40A: dout <= 8'b11111111; // 1034 : 255 - 0xff
      11'h40B: dout <= 8'b11111111; // 1035 : 255 - 0xff
      11'h40C: dout <= 8'b11111111; // 1036 : 255 - 0xff
      11'h40D: dout <= 8'b11111111; // 1037 : 255 - 0xff
      11'h40E: dout <= 8'b11111111; // 1038 : 255 - 0xff
      11'h40F: dout <= 8'b11111111; // 1039 : 255 - 0xff
      11'h410: dout <= 8'b11111111; // 1040 : 255 - 0xff -- Sprite 0x82
      11'h411: dout <= 8'b11111111; // 1041 : 255 - 0xff
      11'h412: dout <= 8'b11111111; // 1042 : 255 - 0xff
      11'h413: dout <= 8'b11111111; // 1043 : 255 - 0xff
      11'h414: dout <= 8'b11111111; // 1044 : 255 - 0xff
      11'h415: dout <= 8'b11111111; // 1045 : 255 - 0xff
      11'h416: dout <= 8'b11111111; // 1046 : 255 - 0xff
      11'h417: dout <= 8'b11111111; // 1047 : 255 - 0xff
      11'h418: dout <= 8'b11111111; // 1048 : 255 - 0xff -- Sprite 0x83
      11'h419: dout <= 8'b11111111; // 1049 : 255 - 0xff
      11'h41A: dout <= 8'b11111111; // 1050 : 255 - 0xff
      11'h41B: dout <= 8'b11111111; // 1051 : 255 - 0xff
      11'h41C: dout <= 8'b11111111; // 1052 : 255 - 0xff
      11'h41D: dout <= 8'b11111111; // 1053 : 255 - 0xff
      11'h41E: dout <= 8'b11111111; // 1054 : 255 - 0xff
      11'h41F: dout <= 8'b11111111; // 1055 : 255 - 0xff
      11'h420: dout <= 8'b11111111; // 1056 : 255 - 0xff -- Sprite 0x84
      11'h421: dout <= 8'b11111111; // 1057 : 255 - 0xff
      11'h422: dout <= 8'b11111111; // 1058 : 255 - 0xff
      11'h423: dout <= 8'b11111111; // 1059 : 255 - 0xff
      11'h424: dout <= 8'b11111111; // 1060 : 255 - 0xff
      11'h425: dout <= 8'b11111111; // 1061 : 255 - 0xff
      11'h426: dout <= 8'b11111111; // 1062 : 255 - 0xff
      11'h427: dout <= 8'b11111111; // 1063 : 255 - 0xff
      11'h428: dout <= 8'b11111111; // 1064 : 255 - 0xff -- Sprite 0x85
      11'h429: dout <= 8'b11111111; // 1065 : 255 - 0xff
      11'h42A: dout <= 8'b11111111; // 1066 : 255 - 0xff
      11'h42B: dout <= 8'b11111111; // 1067 : 255 - 0xff
      11'h42C: dout <= 8'b11111111; // 1068 : 255 - 0xff
      11'h42D: dout <= 8'b11111111; // 1069 : 255 - 0xff
      11'h42E: dout <= 8'b11111111; // 1070 : 255 - 0xff
      11'h42F: dout <= 8'b11111111; // 1071 : 255 - 0xff
      11'h430: dout <= 8'b11111111; // 1072 : 255 - 0xff -- Sprite 0x86
      11'h431: dout <= 8'b11111111; // 1073 : 255 - 0xff
      11'h432: dout <= 8'b11111111; // 1074 : 255 - 0xff
      11'h433: dout <= 8'b11111111; // 1075 : 255 - 0xff
      11'h434: dout <= 8'b11111111; // 1076 : 255 - 0xff
      11'h435: dout <= 8'b11111111; // 1077 : 255 - 0xff
      11'h436: dout <= 8'b11111111; // 1078 : 255 - 0xff
      11'h437: dout <= 8'b11111111; // 1079 : 255 - 0xff
      11'h438: dout <= 8'b11111111; // 1080 : 255 - 0xff -- Sprite 0x87
      11'h439: dout <= 8'b11111111; // 1081 : 255 - 0xff
      11'h43A: dout <= 8'b11111111; // 1082 : 255 - 0xff
      11'h43B: dout <= 8'b11111111; // 1083 : 255 - 0xff
      11'h43C: dout <= 8'b11111111; // 1084 : 255 - 0xff
      11'h43D: dout <= 8'b11111111; // 1085 : 255 - 0xff
      11'h43E: dout <= 8'b11111111; // 1086 : 255 - 0xff
      11'h43F: dout <= 8'b11111111; // 1087 : 255 - 0xff
      11'h440: dout <= 8'b11111111; // 1088 : 255 - 0xff -- Sprite 0x88
      11'h441: dout <= 8'b11111111; // 1089 : 255 - 0xff
      11'h442: dout <= 8'b11111111; // 1090 : 255 - 0xff
      11'h443: dout <= 8'b11111111; // 1091 : 255 - 0xff
      11'h444: dout <= 8'b11111111; // 1092 : 255 - 0xff
      11'h445: dout <= 8'b11111111; // 1093 : 255 - 0xff
      11'h446: dout <= 8'b11111111; // 1094 : 255 - 0xff
      11'h447: dout <= 8'b11111111; // 1095 : 255 - 0xff
      11'h448: dout <= 8'b11111111; // 1096 : 255 - 0xff -- Sprite 0x89
      11'h449: dout <= 8'b11111111; // 1097 : 255 - 0xff
      11'h44A: dout <= 8'b11111111; // 1098 : 255 - 0xff
      11'h44B: dout <= 8'b11111111; // 1099 : 255 - 0xff
      11'h44C: dout <= 8'b11111111; // 1100 : 255 - 0xff
      11'h44D: dout <= 8'b11111111; // 1101 : 255 - 0xff
      11'h44E: dout <= 8'b11111111; // 1102 : 255 - 0xff
      11'h44F: dout <= 8'b11111111; // 1103 : 255 - 0xff
      11'h450: dout <= 8'b11111111; // 1104 : 255 - 0xff -- Sprite 0x8a
      11'h451: dout <= 8'b11111111; // 1105 : 255 - 0xff
      11'h452: dout <= 8'b11111111; // 1106 : 255 - 0xff
      11'h453: dout <= 8'b11111111; // 1107 : 255 - 0xff
      11'h454: dout <= 8'b11111111; // 1108 : 255 - 0xff
      11'h455: dout <= 8'b11111111; // 1109 : 255 - 0xff
      11'h456: dout <= 8'b11111111; // 1110 : 255 - 0xff
      11'h457: dout <= 8'b11111111; // 1111 : 255 - 0xff
      11'h458: dout <= 8'b11111111; // 1112 : 255 - 0xff -- Sprite 0x8b
      11'h459: dout <= 8'b11111111; // 1113 : 255 - 0xff
      11'h45A: dout <= 8'b11111111; // 1114 : 255 - 0xff
      11'h45B: dout <= 8'b11111111; // 1115 : 255 - 0xff
      11'h45C: dout <= 8'b11111111; // 1116 : 255 - 0xff
      11'h45D: dout <= 8'b11111111; // 1117 : 255 - 0xff
      11'h45E: dout <= 8'b11111111; // 1118 : 255 - 0xff
      11'h45F: dout <= 8'b11111111; // 1119 : 255 - 0xff
      11'h460: dout <= 8'b11111111; // 1120 : 255 - 0xff -- Sprite 0x8c
      11'h461: dout <= 8'b11111111; // 1121 : 255 - 0xff
      11'h462: dout <= 8'b11111111; // 1122 : 255 - 0xff
      11'h463: dout <= 8'b11111111; // 1123 : 255 - 0xff
      11'h464: dout <= 8'b11111111; // 1124 : 255 - 0xff
      11'h465: dout <= 8'b11111111; // 1125 : 255 - 0xff
      11'h466: dout <= 8'b11111111; // 1126 : 255 - 0xff
      11'h467: dout <= 8'b11111111; // 1127 : 255 - 0xff
      11'h468: dout <= 8'b11111111; // 1128 : 255 - 0xff -- Sprite 0x8d
      11'h469: dout <= 8'b11111111; // 1129 : 255 - 0xff
      11'h46A: dout <= 8'b11111111; // 1130 : 255 - 0xff
      11'h46B: dout <= 8'b11111111; // 1131 : 255 - 0xff
      11'h46C: dout <= 8'b11111111; // 1132 : 255 - 0xff
      11'h46D: dout <= 8'b11111111; // 1133 : 255 - 0xff
      11'h46E: dout <= 8'b11111111; // 1134 : 255 - 0xff
      11'h46F: dout <= 8'b11111111; // 1135 : 255 - 0xff
      11'h470: dout <= 8'b11111111; // 1136 : 255 - 0xff -- Sprite 0x8e
      11'h471: dout <= 8'b11111111; // 1137 : 255 - 0xff
      11'h472: dout <= 8'b11111111; // 1138 : 255 - 0xff
      11'h473: dout <= 8'b11111111; // 1139 : 255 - 0xff
      11'h474: dout <= 8'b11111111; // 1140 : 255 - 0xff
      11'h475: dout <= 8'b11111111; // 1141 : 255 - 0xff
      11'h476: dout <= 8'b11111111; // 1142 : 255 - 0xff
      11'h477: dout <= 8'b11111111; // 1143 : 255 - 0xff
      11'h478: dout <= 8'b11111111; // 1144 : 255 - 0xff -- Sprite 0x8f
      11'h479: dout <= 8'b11111111; // 1145 : 255 - 0xff
      11'h47A: dout <= 8'b11111111; // 1146 : 255 - 0xff
      11'h47B: dout <= 8'b11111111; // 1147 : 255 - 0xff
      11'h47C: dout <= 8'b11111111; // 1148 : 255 - 0xff
      11'h47D: dout <= 8'b11111111; // 1149 : 255 - 0xff
      11'h47E: dout <= 8'b11111111; // 1150 : 255 - 0xff
      11'h47F: dout <= 8'b11111111; // 1151 : 255 - 0xff
      11'h480: dout <= 8'b00000000; // 1152 :   0 - 0x0 -- Sprite 0x90
      11'h481: dout <= 8'b00000000; // 1153 :   0 - 0x0
      11'h482: dout <= 8'b00000000; // 1154 :   0 - 0x0
      11'h483: dout <= 8'b00000000; // 1155 :   0 - 0x0
      11'h484: dout <= 8'b00000000; // 1156 :   0 - 0x0
      11'h485: dout <= 8'b00000001; // 1157 :   1 - 0x1
      11'h486: dout <= 8'b00011110; // 1158 :  30 - 0x1e
      11'h487: dout <= 8'b00111011; // 1159 :  59 - 0x3b
      11'h488: dout <= 8'b00000000; // 1160 :   0 - 0x0 -- Sprite 0x91
      11'h489: dout <= 8'b00000000; // 1161 :   0 - 0x0
      11'h48A: dout <= 8'b00001100; // 1162 :  12 - 0xc
      11'h48B: dout <= 8'b00111100; // 1163 :  60 - 0x3c
      11'h48C: dout <= 8'b11010000; // 1164 : 208 - 0xd0
      11'h48D: dout <= 8'b00010000; // 1165 :  16 - 0x10
      11'h48E: dout <= 8'b00100000; // 1166 :  32 - 0x20
      11'h48F: dout <= 8'b01000000; // 1167 :  64 - 0x40
      11'h490: dout <= 8'b00111110; // 1168 :  62 - 0x3e -- Sprite 0x92
      11'h491: dout <= 8'b00101101; // 1169 :  45 - 0x2d
      11'h492: dout <= 8'b00110101; // 1170 :  53 - 0x35
      11'h493: dout <= 8'b00011101; // 1171 :  29 - 0x1d
      11'h494: dout <= 8'b00000001; // 1172 :   1 - 0x1
      11'h495: dout <= 8'b00000000; // 1173 :   0 - 0x0
      11'h496: dout <= 8'b00000000; // 1174 :   0 - 0x0
      11'h497: dout <= 8'b00000000; // 1175 :   0 - 0x0
      11'h498: dout <= 8'b10110000; // 1176 : 176 - 0xb0 -- Sprite 0x93
      11'h499: dout <= 8'b10111000; // 1177 : 184 - 0xb8
      11'h49A: dout <= 8'b11111000; // 1178 : 248 - 0xf8
      11'h49B: dout <= 8'b01111000; // 1179 : 120 - 0x78
      11'h49C: dout <= 8'b10011000; // 1180 : 152 - 0x98
      11'h49D: dout <= 8'b11110000; // 1181 : 240 - 0xf0
      11'h49E: dout <= 8'b00000000; // 1182 :   0 - 0x0
      11'h49F: dout <= 8'b00000000; // 1183 :   0 - 0x0
      11'h4A0: dout <= 8'b00000000; // 1184 :   0 - 0x0 -- Sprite 0x94
      11'h4A1: dout <= 8'b00000000; // 1185 :   0 - 0x0
      11'h4A2: dout <= 8'b00000111; // 1186 :   7 - 0x7
      11'h4A3: dout <= 8'b00000011; // 1187 :   3 - 0x3
      11'h4A4: dout <= 8'b00001101; // 1188 :  13 - 0xd
      11'h4A5: dout <= 8'b00011110; // 1189 :  30 - 0x1e
      11'h4A6: dout <= 8'b00010111; // 1190 :  23 - 0x17
      11'h4A7: dout <= 8'b00011101; // 1191 :  29 - 0x1d
      11'h4A8: dout <= 8'b00000000; // 1192 :   0 - 0x0 -- Sprite 0x95
      11'h4A9: dout <= 8'b10000000; // 1193 : 128 - 0x80
      11'h4AA: dout <= 8'b01110000; // 1194 : 112 - 0x70
      11'h4AB: dout <= 8'b11100000; // 1195 : 224 - 0xe0
      11'h4AC: dout <= 8'b11011000; // 1196 : 216 - 0xd8
      11'h4AD: dout <= 8'b10111100; // 1197 : 188 - 0xbc
      11'h4AE: dout <= 8'b01110100; // 1198 : 116 - 0x74
      11'h4AF: dout <= 8'b11011100; // 1199 : 220 - 0xdc
      11'h4B0: dout <= 8'b00011111; // 1200 :  31 - 0x1f -- Sprite 0x96
      11'h4B1: dout <= 8'b00001011; // 1201 :  11 - 0xb
      11'h4B2: dout <= 8'b00001111; // 1202 :  15 - 0xf
      11'h4B3: dout <= 8'b00000101; // 1203 :   5 - 0x5
      11'h4B4: dout <= 8'b00000011; // 1204 :   3 - 0x3
      11'h4B5: dout <= 8'b00000001; // 1205 :   1 - 0x1
      11'h4B6: dout <= 8'b00000000; // 1206 :   0 - 0x0
      11'h4B7: dout <= 8'b00000000; // 1207 :   0 - 0x0
      11'h4B8: dout <= 8'b11111100; // 1208 : 252 - 0xfc -- Sprite 0x97
      11'h4B9: dout <= 8'b01101000; // 1209 : 104 - 0x68
      11'h4BA: dout <= 8'b11111000; // 1210 : 248 - 0xf8
      11'h4BB: dout <= 8'b10110000; // 1211 : 176 - 0xb0
      11'h4BC: dout <= 8'b11100000; // 1212 : 224 - 0xe0
      11'h4BD: dout <= 8'b10000000; // 1213 : 128 - 0x80
      11'h4BE: dout <= 8'b00000000; // 1214 :   0 - 0x0
      11'h4BF: dout <= 8'b00000000; // 1215 :   0 - 0x0
      11'h4C0: dout <= 8'b00000000; // 1216 :   0 - 0x0 -- Sprite 0x98
      11'h4C1: dout <= 8'b00000000; // 1217 :   0 - 0x0
      11'h4C2: dout <= 8'b00000000; // 1218 :   0 - 0x0
      11'h4C3: dout <= 8'b00000001; // 1219 :   1 - 0x1
      11'h4C4: dout <= 8'b00000001; // 1220 :   1 - 0x1
      11'h4C5: dout <= 8'b00001011; // 1221 :  11 - 0xb
      11'h4C6: dout <= 8'b00011100; // 1222 :  28 - 0x1c
      11'h4C7: dout <= 8'b00111111; // 1223 :  63 - 0x3f
      11'h4C8: dout <= 8'b00000000; // 1224 :   0 - 0x0 -- Sprite 0x99
      11'h4C9: dout <= 8'b00000000; // 1225 :   0 - 0x0
      11'h4CA: dout <= 8'b00110000; // 1226 :  48 - 0x30
      11'h4CB: dout <= 8'b01111000; // 1227 : 120 - 0x78
      11'h4CC: dout <= 8'b10000000; // 1228 : 128 - 0x80
      11'h4CD: dout <= 8'b11110000; // 1229 : 240 - 0xf0
      11'h4CE: dout <= 8'b11111000; // 1230 : 248 - 0xf8
      11'h4CF: dout <= 8'b11111100; // 1231 : 252 - 0xfc
      11'h4D0: dout <= 8'b00111111; // 1232 :  63 - 0x3f -- Sprite 0x9a
      11'h4D1: dout <= 8'b00111111; // 1233 :  63 - 0x3f
      11'h4D2: dout <= 8'b00111111; // 1234 :  63 - 0x3f
      11'h4D3: dout <= 8'b00011111; // 1235 :  31 - 0x1f
      11'h4D4: dout <= 8'b00011111; // 1236 :  31 - 0x1f
      11'h4D5: dout <= 8'b00000111; // 1237 :   7 - 0x7
      11'h4D6: dout <= 8'b00000000; // 1238 :   0 - 0x0
      11'h4D7: dout <= 8'b00000000; // 1239 :   0 - 0x0
      11'h4D8: dout <= 8'b11111100; // 1240 : 252 - 0xfc -- Sprite 0x9b
      11'h4D9: dout <= 8'b11101100; // 1241 : 236 - 0xec
      11'h4DA: dout <= 8'b11101100; // 1242 : 236 - 0xec
      11'h4DB: dout <= 8'b11011000; // 1243 : 216 - 0xd8
      11'h4DC: dout <= 8'b11111000; // 1244 : 248 - 0xf8
      11'h4DD: dout <= 8'b11100000; // 1245 : 224 - 0xe0
      11'h4DE: dout <= 8'b00000000; // 1246 :   0 - 0x0
      11'h4DF: dout <= 8'b00000000; // 1247 :   0 - 0x0
      11'h4E0: dout <= 8'b00000000; // 1248 :   0 - 0x0 -- Sprite 0x9c
      11'h4E1: dout <= 8'b00000000; // 1249 :   0 - 0x0
      11'h4E2: dout <= 8'b00000001; // 1250 :   1 - 0x1
      11'h4E3: dout <= 8'b00011101; // 1251 :  29 - 0x1d
      11'h4E4: dout <= 8'b00111110; // 1252 :  62 - 0x3e
      11'h4E5: dout <= 8'b00111111; // 1253 :  63 - 0x3f
      11'h4E6: dout <= 8'b00111111; // 1254 :  63 - 0x3f
      11'h4E7: dout <= 8'b00111111; // 1255 :  63 - 0x3f
      11'h4E8: dout <= 8'b00000000; // 1256 :   0 - 0x0 -- Sprite 0x9d
      11'h4E9: dout <= 8'b10000000; // 1257 : 128 - 0x80
      11'h4EA: dout <= 8'b00000000; // 1258 :   0 - 0x0
      11'h4EB: dout <= 8'b01110000; // 1259 : 112 - 0x70
      11'h4EC: dout <= 8'b11111000; // 1260 : 248 - 0xf8
      11'h4ED: dout <= 8'b11111100; // 1261 : 252 - 0xfc
      11'h4EE: dout <= 8'b11111100; // 1262 : 252 - 0xfc
      11'h4EF: dout <= 8'b11111100; // 1263 : 252 - 0xfc
      11'h4F0: dout <= 8'b00111111; // 1264 :  63 - 0x3f -- Sprite 0x9e
      11'h4F1: dout <= 8'b00111111; // 1265 :  63 - 0x3f
      11'h4F2: dout <= 8'b00011111; // 1266 :  31 - 0x1f
      11'h4F3: dout <= 8'b00011111; // 1267 :  31 - 0x1f
      11'h4F4: dout <= 8'b00001111; // 1268 :  15 - 0xf
      11'h4F5: dout <= 8'b00000110; // 1269 :   6 - 0x6
      11'h4F6: dout <= 8'b00000000; // 1270 :   0 - 0x0
      11'h4F7: dout <= 8'b00000000; // 1271 :   0 - 0x0
      11'h4F8: dout <= 8'b11101100; // 1272 : 236 - 0xec -- Sprite 0x9f
      11'h4F9: dout <= 8'b11101100; // 1273 : 236 - 0xec
      11'h4FA: dout <= 8'b11011000; // 1274 : 216 - 0xd8
      11'h4FB: dout <= 8'b11111000; // 1275 : 248 - 0xf8
      11'h4FC: dout <= 8'b11110000; // 1276 : 240 - 0xf0
      11'h4FD: dout <= 8'b11100000; // 1277 : 224 - 0xe0
      11'h4FE: dout <= 8'b00000000; // 1278 :   0 - 0x0
      11'h4FF: dout <= 8'b00000000; // 1279 :   0 - 0x0
      11'h500: dout <= 8'b00000000; // 1280 :   0 - 0x0 -- Sprite 0xa0
      11'h501: dout <= 8'b00000100; // 1281 :   4 - 0x4
      11'h502: dout <= 8'b00000011; // 1282 :   3 - 0x3
      11'h503: dout <= 8'b00000000; // 1283 :   0 - 0x0
      11'h504: dout <= 8'b00000001; // 1284 :   1 - 0x1
      11'h505: dout <= 8'b00000111; // 1285 :   7 - 0x7
      11'h506: dout <= 8'b00001111; // 1286 :  15 - 0xf
      11'h507: dout <= 8'b00001100; // 1287 :  12 - 0xc
      11'h508: dout <= 8'b00000000; // 1288 :   0 - 0x0 -- Sprite 0xa1
      11'h509: dout <= 8'b00000000; // 1289 :   0 - 0x0
      11'h50A: dout <= 8'b11100000; // 1290 : 224 - 0xe0
      11'h50B: dout <= 8'b10000000; // 1291 : 128 - 0x80
      11'h50C: dout <= 8'b01000000; // 1292 :  64 - 0x40
      11'h50D: dout <= 8'b11110000; // 1293 : 240 - 0xf0
      11'h50E: dout <= 8'b10011000; // 1294 : 152 - 0x98
      11'h50F: dout <= 8'b11111000; // 1295 : 248 - 0xf8
      11'h510: dout <= 8'b00011111; // 1296 :  31 - 0x1f -- Sprite 0xa2
      11'h511: dout <= 8'b00010011; // 1297 :  19 - 0x13
      11'h512: dout <= 8'b00011111; // 1298 :  31 - 0x1f
      11'h513: dout <= 8'b00001111; // 1299 :  15 - 0xf
      11'h514: dout <= 8'b00001001; // 1300 :   9 - 0x9
      11'h515: dout <= 8'b00000111; // 1301 :   7 - 0x7
      11'h516: dout <= 8'b00000001; // 1302 :   1 - 0x1
      11'h517: dout <= 8'b00000000; // 1303 :   0 - 0x0
      11'h518: dout <= 8'b11100100; // 1304 : 228 - 0xe4 -- Sprite 0xa3
      11'h519: dout <= 8'b00111100; // 1305 :  60 - 0x3c
      11'h51A: dout <= 8'b11100100; // 1306 : 228 - 0xe4
      11'h51B: dout <= 8'b00111000; // 1307 :  56 - 0x38
      11'h51C: dout <= 8'b11111000; // 1308 : 248 - 0xf8
      11'h51D: dout <= 8'b11110000; // 1309 : 240 - 0xf0
      11'h51E: dout <= 8'b11000000; // 1310 : 192 - 0xc0
      11'h51F: dout <= 8'b00000000; // 1311 :   0 - 0x0
      11'h520: dout <= 8'b00000000; // 1312 :   0 - 0x0 -- Sprite 0xa4
      11'h521: dout <= 8'b00000000; // 1313 :   0 - 0x0
      11'h522: dout <= 8'b00000000; // 1314 :   0 - 0x0
      11'h523: dout <= 8'b00000000; // 1315 :   0 - 0x0
      11'h524: dout <= 8'b00010001; // 1316 :  17 - 0x11
      11'h525: dout <= 8'b00010011; // 1317 :  19 - 0x13
      11'h526: dout <= 8'b00011111; // 1318 :  31 - 0x1f
      11'h527: dout <= 8'b00011111; // 1319 :  31 - 0x1f
      11'h528: dout <= 8'b00000000; // 1320 :   0 - 0x0 -- Sprite 0xa5
      11'h529: dout <= 8'b00000000; // 1321 :   0 - 0x0
      11'h52A: dout <= 8'b00000000; // 1322 :   0 - 0x0
      11'h52B: dout <= 8'b10000000; // 1323 : 128 - 0x80
      11'h52C: dout <= 8'b11000100; // 1324 : 196 - 0xc4
      11'h52D: dout <= 8'b11100100; // 1325 : 228 - 0xe4
      11'h52E: dout <= 8'b11111100; // 1326 : 252 - 0xfc
      11'h52F: dout <= 8'b11111100; // 1327 : 252 - 0xfc
      11'h530: dout <= 8'b00011111; // 1328 :  31 - 0x1f -- Sprite 0xa6
      11'h531: dout <= 8'b00001110; // 1329 :  14 - 0xe
      11'h532: dout <= 8'b00000110; // 1330 :   6 - 0x6
      11'h533: dout <= 8'b00000010; // 1331 :   2 - 0x2
      11'h534: dout <= 8'b00000000; // 1332 :   0 - 0x0
      11'h535: dout <= 8'b00000000; // 1333 :   0 - 0x0
      11'h536: dout <= 8'b00000000; // 1334 :   0 - 0x0
      11'h537: dout <= 8'b00000000; // 1335 :   0 - 0x0
      11'h538: dout <= 8'b11111100; // 1336 : 252 - 0xfc -- Sprite 0xa7
      11'h539: dout <= 8'b10111000; // 1337 : 184 - 0xb8
      11'h53A: dout <= 8'b10110000; // 1338 : 176 - 0xb0
      11'h53B: dout <= 8'b10100000; // 1339 : 160 - 0xa0
      11'h53C: dout <= 8'b10000000; // 1340 : 128 - 0x80
      11'h53D: dout <= 8'b00000000; // 1341 :   0 - 0x0
      11'h53E: dout <= 8'b00000000; // 1342 :   0 - 0x0
      11'h53F: dout <= 8'b00000000; // 1343 :   0 - 0x0
      11'h540: dout <= 8'b00000000; // 1344 :   0 - 0x0 -- Sprite 0xa8
      11'h541: dout <= 8'b00000000; // 1345 :   0 - 0x0
      11'h542: dout <= 8'b00000000; // 1346 :   0 - 0x0
      11'h543: dout <= 8'b00000001; // 1347 :   1 - 0x1
      11'h544: dout <= 8'b00000011; // 1348 :   3 - 0x3
      11'h545: dout <= 8'b00000110; // 1349 :   6 - 0x6
      11'h546: dout <= 8'b00000110; // 1350 :   6 - 0x6
      11'h547: dout <= 8'b00001111; // 1351 :  15 - 0xf
      11'h548: dout <= 8'b00000000; // 1352 :   0 - 0x0 -- Sprite 0xa9
      11'h549: dout <= 8'b00011000; // 1353 :  24 - 0x18
      11'h54A: dout <= 8'b11110100; // 1354 : 244 - 0xf4
      11'h54B: dout <= 8'b11111000; // 1355 : 248 - 0xf8
      11'h54C: dout <= 8'b00111000; // 1356 :  56 - 0x38
      11'h54D: dout <= 8'b01111100; // 1357 : 124 - 0x7c
      11'h54E: dout <= 8'b11111100; // 1358 : 252 - 0xfc
      11'h54F: dout <= 8'b11111100; // 1359 : 252 - 0xfc
      11'h550: dout <= 8'b00001111; // 1360 :  15 - 0xf -- Sprite 0xaa
      11'h551: dout <= 8'b00011111; // 1361 :  31 - 0x1f
      11'h552: dout <= 8'b00110000; // 1362 :  48 - 0x30
      11'h553: dout <= 8'b00111000; // 1363 :  56 - 0x38
      11'h554: dout <= 8'b00011101; // 1364 :  29 - 0x1d
      11'h555: dout <= 8'b00000011; // 1365 :   3 - 0x3
      11'h556: dout <= 8'b00000011; // 1366 :   3 - 0x3
      11'h557: dout <= 8'b00000000; // 1367 :   0 - 0x0
      11'h558: dout <= 8'b11111100; // 1368 : 252 - 0xfc -- Sprite 0xab
      11'h559: dout <= 8'b11111100; // 1369 : 252 - 0xfc
      11'h55A: dout <= 8'b01111100; // 1370 : 124 - 0x7c
      11'h55B: dout <= 8'b10001110; // 1371 : 142 - 0x8e
      11'h55C: dout <= 8'b10000110; // 1372 : 134 - 0x86
      11'h55D: dout <= 8'b10011100; // 1373 : 156 - 0x9c
      11'h55E: dout <= 8'b01111000; // 1374 : 120 - 0x78
      11'h55F: dout <= 8'b00000000; // 1375 :   0 - 0x0
      11'h560: dout <= 8'b00000000; // 1376 :   0 - 0x0 -- Sprite 0xac
      11'h561: dout <= 8'b00000001; // 1377 :   1 - 0x1
      11'h562: dout <= 8'b00000110; // 1378 :   6 - 0x6
      11'h563: dout <= 8'b00000111; // 1379 :   7 - 0x7
      11'h564: dout <= 8'b00000111; // 1380 :   7 - 0x7
      11'h565: dout <= 8'b00000111; // 1381 :   7 - 0x7
      11'h566: dout <= 8'b00000001; // 1382 :   1 - 0x1
      11'h567: dout <= 8'b00000011; // 1383 :   3 - 0x3
      11'h568: dout <= 8'b00000000; // 1384 :   0 - 0x0 -- Sprite 0xad
      11'h569: dout <= 8'b11000000; // 1385 : 192 - 0xc0
      11'h56A: dout <= 8'b00110000; // 1386 :  48 - 0x30
      11'h56B: dout <= 8'b11110000; // 1387 : 240 - 0xf0
      11'h56C: dout <= 8'b11110000; // 1388 : 240 - 0xf0
      11'h56D: dout <= 8'b11110000; // 1389 : 240 - 0xf0
      11'h56E: dout <= 8'b01000000; // 1390 :  64 - 0x40
      11'h56F: dout <= 8'b01000000; // 1391 :  64 - 0x40
      11'h570: dout <= 8'b00000001; // 1392 :   1 - 0x1 -- Sprite 0xae
      11'h571: dout <= 8'b00000000; // 1393 :   0 - 0x0
      11'h572: dout <= 8'b00000001; // 1394 :   1 - 0x1
      11'h573: dout <= 8'b00000011; // 1395 :   3 - 0x3
      11'h574: dout <= 8'b00000001; // 1396 :   1 - 0x1
      11'h575: dout <= 8'b00000000; // 1397 :   0 - 0x0
      11'h576: dout <= 8'b00000000; // 1398 :   0 - 0x0
      11'h577: dout <= 8'b00000000; // 1399 :   0 - 0x0
      11'h578: dout <= 8'b01000000; // 1400 :  64 - 0x40 -- Sprite 0xaf
      11'h579: dout <= 8'b01000000; // 1401 :  64 - 0x40
      11'h57A: dout <= 8'b01000000; // 1402 :  64 - 0x40
      11'h57B: dout <= 8'b01000000; // 1403 :  64 - 0x40
      11'h57C: dout <= 8'b01000000; // 1404 :  64 - 0x40
      11'h57D: dout <= 8'b10000000; // 1405 : 128 - 0x80
      11'h57E: dout <= 8'b00000000; // 1406 :   0 - 0x0
      11'h57F: dout <= 8'b00000000; // 1407 :   0 - 0x0
      11'h580: dout <= 8'b01111110; // 1408 : 126 - 0x7e -- Sprite 0xb0
      11'h581: dout <= 8'b01100011; // 1409 :  99 - 0x63
      11'h582: dout <= 8'b01100011; // 1410 :  99 - 0x63
      11'h583: dout <= 8'b01100011; // 1411 :  99 - 0x63
      11'h584: dout <= 8'b01111110; // 1412 : 126 - 0x7e
      11'h585: dout <= 8'b01100000; // 1413 :  96 - 0x60
      11'h586: dout <= 8'b01100000; // 1414 :  96 - 0x60
      11'h587: dout <= 8'b00000000; // 1415 :   0 - 0x0
      11'h588: dout <= 8'b01100000; // 1416 :  96 - 0x60 -- Sprite 0xb1
      11'h589: dout <= 8'b01100000; // 1417 :  96 - 0x60
      11'h58A: dout <= 8'b01100000; // 1418 :  96 - 0x60
      11'h58B: dout <= 8'b01100000; // 1419 :  96 - 0x60
      11'h58C: dout <= 8'b01100000; // 1420 :  96 - 0x60
      11'h58D: dout <= 8'b01100000; // 1421 :  96 - 0x60
      11'h58E: dout <= 8'b01111111; // 1422 : 127 - 0x7f
      11'h58F: dout <= 8'b00000000; // 1423 :   0 - 0x0
      11'h590: dout <= 8'b00011100; // 1424 :  28 - 0x1c -- Sprite 0xb2
      11'h591: dout <= 8'b00110110; // 1425 :  54 - 0x36
      11'h592: dout <= 8'b01100011; // 1426 :  99 - 0x63
      11'h593: dout <= 8'b01100011; // 1427 :  99 - 0x63
      11'h594: dout <= 8'b01111111; // 1428 : 127 - 0x7f
      11'h595: dout <= 8'b01100011; // 1429 :  99 - 0x63
      11'h596: dout <= 8'b01100011; // 1430 :  99 - 0x63
      11'h597: dout <= 8'b00000000; // 1431 :   0 - 0x0
      11'h598: dout <= 8'b00110011; // 1432 :  51 - 0x33 -- Sprite 0xb3
      11'h599: dout <= 8'b00110011; // 1433 :  51 - 0x33
      11'h59A: dout <= 8'b00110011; // 1434 :  51 - 0x33
      11'h59B: dout <= 8'b00011110; // 1435 :  30 - 0x1e
      11'h59C: dout <= 8'b00001100; // 1436 :  12 - 0xc
      11'h59D: dout <= 8'b00001100; // 1437 :  12 - 0xc
      11'h59E: dout <= 8'b00001100; // 1438 :  12 - 0xc
      11'h59F: dout <= 8'b00000000; // 1439 :   0 - 0x0
      11'h5A0: dout <= 8'b01111111; // 1440 : 127 - 0x7f -- Sprite 0xb4
      11'h5A1: dout <= 8'b01100000; // 1441 :  96 - 0x60
      11'h5A2: dout <= 8'b01100000; // 1442 :  96 - 0x60
      11'h5A3: dout <= 8'b01111110; // 1443 : 126 - 0x7e
      11'h5A4: dout <= 8'b01100000; // 1444 :  96 - 0x60
      11'h5A5: dout <= 8'b01100000; // 1445 :  96 - 0x60
      11'h5A6: dout <= 8'b01111111; // 1446 : 127 - 0x7f
      11'h5A7: dout <= 8'b00000000; // 1447 :   0 - 0x0
      11'h5A8: dout <= 8'b01111110; // 1448 : 126 - 0x7e -- Sprite 0xb5
      11'h5A9: dout <= 8'b01100011; // 1449 :  99 - 0x63
      11'h5AA: dout <= 8'b01100011; // 1450 :  99 - 0x63
      11'h5AB: dout <= 8'b01100111; // 1451 : 103 - 0x67
      11'h5AC: dout <= 8'b01111100; // 1452 : 124 - 0x7c
      11'h5AD: dout <= 8'b01101110; // 1453 : 110 - 0x6e
      11'h5AE: dout <= 8'b01100111; // 1454 : 103 - 0x67
      11'h5AF: dout <= 8'b00000000; // 1455 :   0 - 0x0
      11'h5B0: dout <= 8'b00111110; // 1456 :  62 - 0x3e -- Sprite 0xb6
      11'h5B1: dout <= 8'b01100011; // 1457 :  99 - 0x63
      11'h5B2: dout <= 8'b01100011; // 1458 :  99 - 0x63
      11'h5B3: dout <= 8'b01100011; // 1459 :  99 - 0x63
      11'h5B4: dout <= 8'b01100011; // 1460 :  99 - 0x63
      11'h5B5: dout <= 8'b01100011; // 1461 :  99 - 0x63
      11'h5B6: dout <= 8'b00111110; // 1462 :  62 - 0x3e
      11'h5B7: dout <= 8'b00000000; // 1463 :   0 - 0x0
      11'h5B8: dout <= 8'b01100011; // 1464 :  99 - 0x63 -- Sprite 0xb7
      11'h5B9: dout <= 8'b01110011; // 1465 : 115 - 0x73
      11'h5BA: dout <= 8'b01111011; // 1466 : 123 - 0x7b
      11'h5BB: dout <= 8'b01111111; // 1467 : 127 - 0x7f
      11'h5BC: dout <= 8'b01101111; // 1468 : 111 - 0x6f
      11'h5BD: dout <= 8'b01100111; // 1469 : 103 - 0x67
      11'h5BE: dout <= 8'b01100011; // 1470 :  99 - 0x63
      11'h5BF: dout <= 8'b00000000; // 1471 :   0 - 0x0
      11'h5C0: dout <= 8'b00111111; // 1472 :  63 - 0x3f -- Sprite 0xb8
      11'h5C1: dout <= 8'b00001100; // 1473 :  12 - 0xc
      11'h5C2: dout <= 8'b00001100; // 1474 :  12 - 0xc
      11'h5C3: dout <= 8'b00001100; // 1475 :  12 - 0xc
      11'h5C4: dout <= 8'b00001100; // 1476 :  12 - 0xc
      11'h5C5: dout <= 8'b00001100; // 1477 :  12 - 0xc
      11'h5C6: dout <= 8'b00001100; // 1478 :  12 - 0xc
      11'h5C7: dout <= 8'b00000000; // 1479 :   0 - 0x0
      11'h5C8: dout <= 8'b01100011; // 1480 :  99 - 0x63 -- Sprite 0xb9
      11'h5C9: dout <= 8'b01100011; // 1481 :  99 - 0x63
      11'h5CA: dout <= 8'b01101011; // 1482 : 107 - 0x6b
      11'h5CB: dout <= 8'b01111111; // 1483 : 127 - 0x7f
      11'h5CC: dout <= 8'b01111111; // 1484 : 127 - 0x7f
      11'h5CD: dout <= 8'b01110111; // 1485 : 119 - 0x77
      11'h5CE: dout <= 8'b01100011; // 1486 :  99 - 0x63
      11'h5CF: dout <= 8'b00000000; // 1487 :   0 - 0x0
      11'h5D0: dout <= 8'b01111100; // 1488 : 124 - 0x7c -- Sprite 0xba
      11'h5D1: dout <= 8'b01100110; // 1489 : 102 - 0x66
      11'h5D2: dout <= 8'b01100011; // 1490 :  99 - 0x63
      11'h5D3: dout <= 8'b01100011; // 1491 :  99 - 0x63
      11'h5D4: dout <= 8'b01100011; // 1492 :  99 - 0x63
      11'h5D5: dout <= 8'b01100110; // 1493 : 102 - 0x66
      11'h5D6: dout <= 8'b01111100; // 1494 : 124 - 0x7c
      11'h5D7: dout <= 8'b00000000; // 1495 :   0 - 0x0
      11'h5D8: dout <= 8'b00011100; // 1496 :  28 - 0x1c -- Sprite 0xbb
      11'h5D9: dout <= 8'b00011100; // 1497 :  28 - 0x1c
      11'h5DA: dout <= 8'b00011100; // 1498 :  28 - 0x1c
      11'h5DB: dout <= 8'b00011000; // 1499 :  24 - 0x18
      11'h5DC: dout <= 8'b00011000; // 1500 :  24 - 0x18
      11'h5DD: dout <= 8'b00000000; // 1501 :   0 - 0x0
      11'h5DE: dout <= 8'b00011000; // 1502 :  24 - 0x18
      11'h5DF: dout <= 8'b00000000; // 1503 :   0 - 0x0
      11'h5E0: dout <= 8'b00011111; // 1504 :  31 - 0x1f -- Sprite 0xbc
      11'h5E1: dout <= 8'b00110000; // 1505 :  48 - 0x30
      11'h5E2: dout <= 8'b01100000; // 1506 :  96 - 0x60
      11'h5E3: dout <= 8'b01100111; // 1507 : 103 - 0x67
      11'h5E4: dout <= 8'b01100011; // 1508 :  99 - 0x63
      11'h5E5: dout <= 8'b00110011; // 1509 :  51 - 0x33
      11'h5E6: dout <= 8'b00011111; // 1510 :  31 - 0x1f
      11'h5E7: dout <= 8'b00000000; // 1511 :   0 - 0x0
      11'h5E8: dout <= 8'b01100011; // 1512 :  99 - 0x63 -- Sprite 0xbd
      11'h5E9: dout <= 8'b01110111; // 1513 : 119 - 0x77
      11'h5EA: dout <= 8'b01111111; // 1514 : 127 - 0x7f
      11'h5EB: dout <= 8'b01111111; // 1515 : 127 - 0x7f
      11'h5EC: dout <= 8'b01101011; // 1516 : 107 - 0x6b
      11'h5ED: dout <= 8'b01100011; // 1517 :  99 - 0x63
      11'h5EE: dout <= 8'b01100011; // 1518 :  99 - 0x63
      11'h5EF: dout <= 8'b00000000; // 1519 :   0 - 0x0
      11'h5F0: dout <= 8'b01100011; // 1520 :  99 - 0x63 -- Sprite 0xbe
      11'h5F1: dout <= 8'b01100011; // 1521 :  99 - 0x63
      11'h5F2: dout <= 8'b01100011; // 1522 :  99 - 0x63
      11'h5F3: dout <= 8'b01110111; // 1523 : 119 - 0x77
      11'h5F4: dout <= 8'b00111110; // 1524 :  62 - 0x3e
      11'h5F5: dout <= 8'b00011100; // 1525 :  28 - 0x1c
      11'h5F6: dout <= 8'b00001000; // 1526 :   8 - 0x8
      11'h5F7: dout <= 8'b00000000; // 1527 :   0 - 0x0
      11'h5F8: dout <= 8'b00000000; // 1528 :   0 - 0x0 -- Sprite 0xbf
      11'h5F9: dout <= 8'b00000000; // 1529 :   0 - 0x0
      11'h5FA: dout <= 8'b00000000; // 1530 :   0 - 0x0
      11'h5FB: dout <= 8'b00000000; // 1531 :   0 - 0x0
      11'h5FC: dout <= 8'b00000000; // 1532 :   0 - 0x0
      11'h5FD: dout <= 8'b00000000; // 1533 :   0 - 0x0
      11'h5FE: dout <= 8'b00000000; // 1534 :   0 - 0x0
      11'h5FF: dout <= 8'b00000000; // 1535 :   0 - 0x0
      11'h600: dout <= 8'b00011111; // 1536 :  31 - 0x1f -- Sprite 0xc0
      11'h601: dout <= 8'b00110000; // 1537 :  48 - 0x30
      11'h602: dout <= 8'b01100000; // 1538 :  96 - 0x60
      11'h603: dout <= 8'b01100111; // 1539 : 103 - 0x67
      11'h604: dout <= 8'b01100011; // 1540 :  99 - 0x63
      11'h605: dout <= 8'b00110011; // 1541 :  51 - 0x33
      11'h606: dout <= 8'b00011111; // 1542 :  31 - 0x1f
      11'h607: dout <= 8'b00000000; // 1543 :   0 - 0x0
      11'h608: dout <= 8'b00011100; // 1544 :  28 - 0x1c -- Sprite 0xc1
      11'h609: dout <= 8'b00110110; // 1545 :  54 - 0x36
      11'h60A: dout <= 8'b01100011; // 1546 :  99 - 0x63
      11'h60B: dout <= 8'b01100011; // 1547 :  99 - 0x63
      11'h60C: dout <= 8'b01111111; // 1548 : 127 - 0x7f
      11'h60D: dout <= 8'b01100011; // 1549 :  99 - 0x63
      11'h60E: dout <= 8'b01100011; // 1550 :  99 - 0x63
      11'h60F: dout <= 8'b00000000; // 1551 :   0 - 0x0
      11'h610: dout <= 8'b01100011; // 1552 :  99 - 0x63 -- Sprite 0xc2
      11'h611: dout <= 8'b01110111; // 1553 : 119 - 0x77
      11'h612: dout <= 8'b01111111; // 1554 : 127 - 0x7f
      11'h613: dout <= 8'b01111111; // 1555 : 127 - 0x7f
      11'h614: dout <= 8'b01101011; // 1556 : 107 - 0x6b
      11'h615: dout <= 8'b01100011; // 1557 :  99 - 0x63
      11'h616: dout <= 8'b01100011; // 1558 :  99 - 0x63
      11'h617: dout <= 8'b00000000; // 1559 :   0 - 0x0
      11'h618: dout <= 8'b01111111; // 1560 : 127 - 0x7f -- Sprite 0xc3
      11'h619: dout <= 8'b01100000; // 1561 :  96 - 0x60
      11'h61A: dout <= 8'b01100000; // 1562 :  96 - 0x60
      11'h61B: dout <= 8'b01111110; // 1563 : 126 - 0x7e
      11'h61C: dout <= 8'b01100000; // 1564 :  96 - 0x60
      11'h61D: dout <= 8'b01100000; // 1565 :  96 - 0x60
      11'h61E: dout <= 8'b01111111; // 1566 : 127 - 0x7f
      11'h61F: dout <= 8'b00000000; // 1567 :   0 - 0x0
      11'h620: dout <= 8'b00111110; // 1568 :  62 - 0x3e -- Sprite 0xc4
      11'h621: dout <= 8'b01100011; // 1569 :  99 - 0x63
      11'h622: dout <= 8'b01100011; // 1570 :  99 - 0x63
      11'h623: dout <= 8'b01100011; // 1571 :  99 - 0x63
      11'h624: dout <= 8'b01100011; // 1572 :  99 - 0x63
      11'h625: dout <= 8'b01100011; // 1573 :  99 - 0x63
      11'h626: dout <= 8'b00111110; // 1574 :  62 - 0x3e
      11'h627: dout <= 8'b00000000; // 1575 :   0 - 0x0
      11'h628: dout <= 8'b01100011; // 1576 :  99 - 0x63 -- Sprite 0xc5
      11'h629: dout <= 8'b01100011; // 1577 :  99 - 0x63
      11'h62A: dout <= 8'b01100011; // 1578 :  99 - 0x63
      11'h62B: dout <= 8'b01110111; // 1579 : 119 - 0x77
      11'h62C: dout <= 8'b00111110; // 1580 :  62 - 0x3e
      11'h62D: dout <= 8'b00011100; // 1581 :  28 - 0x1c
      11'h62E: dout <= 8'b00001000; // 1582 :   8 - 0x8
      11'h62F: dout <= 8'b00000000; // 1583 :   0 - 0x0
      11'h630: dout <= 8'b01111110; // 1584 : 126 - 0x7e -- Sprite 0xc6
      11'h631: dout <= 8'b01100011; // 1585 :  99 - 0x63
      11'h632: dout <= 8'b01100011; // 1586 :  99 - 0x63
      11'h633: dout <= 8'b01100111; // 1587 : 103 - 0x67
      11'h634: dout <= 8'b01111100; // 1588 : 124 - 0x7c
      11'h635: dout <= 8'b01101110; // 1589 : 110 - 0x6e
      11'h636: dout <= 8'b01100111; // 1590 : 103 - 0x67
      11'h637: dout <= 8'b00000000; // 1591 :   0 - 0x0
      11'h638: dout <= 8'b00110011; // 1592 :  51 - 0x33 -- Sprite 0xc7
      11'h639: dout <= 8'b00110011; // 1593 :  51 - 0x33
      11'h63A: dout <= 8'b00110011; // 1594 :  51 - 0x33
      11'h63B: dout <= 8'b00011110; // 1595 :  30 - 0x1e
      11'h63C: dout <= 8'b00001100; // 1596 :  12 - 0xc
      11'h63D: dout <= 8'b00001100; // 1597 :  12 - 0xc
      11'h63E: dout <= 8'b00001100; // 1598 :  12 - 0xc
      11'h63F: dout <= 8'b00000000; // 1599 :   0 - 0x0
      11'h640: dout <= 8'b00000000; // 1600 :   0 - 0x0 -- Sprite 0xc8
      11'h641: dout <= 8'b00000000; // 1601 :   0 - 0x0
      11'h642: dout <= 8'b00000000; // 1602 :   0 - 0x0
      11'h643: dout <= 8'b00000000; // 1603 :   0 - 0x0
      11'h644: dout <= 8'b00000000; // 1604 :   0 - 0x0
      11'h645: dout <= 8'b00000000; // 1605 :   0 - 0x0
      11'h646: dout <= 8'b00000000; // 1606 :   0 - 0x0
      11'h647: dout <= 8'b00000000; // 1607 :   0 - 0x0
      11'h648: dout <= 8'b00000000; // 1608 :   0 - 0x0 -- Sprite 0xc9
      11'h649: dout <= 8'b00000000; // 1609 :   0 - 0x0
      11'h64A: dout <= 8'b00000000; // 1610 :   0 - 0x0
      11'h64B: dout <= 8'b00000000; // 1611 :   0 - 0x0
      11'h64C: dout <= 8'b00000000; // 1612 :   0 - 0x0
      11'h64D: dout <= 8'b00000000; // 1613 :   0 - 0x0
      11'h64E: dout <= 8'b00000000; // 1614 :   0 - 0x0
      11'h64F: dout <= 8'b00000000; // 1615 :   0 - 0x0
      11'h650: dout <= 8'b00000000; // 1616 :   0 - 0x0 -- Sprite 0xca
      11'h651: dout <= 8'b00000000; // 1617 :   0 - 0x0
      11'h652: dout <= 8'b00000000; // 1618 :   0 - 0x0
      11'h653: dout <= 8'b00000000; // 1619 :   0 - 0x0
      11'h654: dout <= 8'b00000000; // 1620 :   0 - 0x0
      11'h655: dout <= 8'b00000000; // 1621 :   0 - 0x0
      11'h656: dout <= 8'b00000000; // 1622 :   0 - 0x0
      11'h657: dout <= 8'b00000000; // 1623 :   0 - 0x0
      11'h658: dout <= 8'b00000000; // 1624 :   0 - 0x0 -- Sprite 0xcb
      11'h659: dout <= 8'b00000000; // 1625 :   0 - 0x0
      11'h65A: dout <= 8'b00000000; // 1626 :   0 - 0x0
      11'h65B: dout <= 8'b00000000; // 1627 :   0 - 0x0
      11'h65C: dout <= 8'b00000000; // 1628 :   0 - 0x0
      11'h65D: dout <= 8'b00000000; // 1629 :   0 - 0x0
      11'h65E: dout <= 8'b00000000; // 1630 :   0 - 0x0
      11'h65F: dout <= 8'b00000000; // 1631 :   0 - 0x0
      11'h660: dout <= 8'b00000000; // 1632 :   0 - 0x0 -- Sprite 0xcc
      11'h661: dout <= 8'b00000000; // 1633 :   0 - 0x0
      11'h662: dout <= 8'b00000000; // 1634 :   0 - 0x0
      11'h663: dout <= 8'b00000000; // 1635 :   0 - 0x0
      11'h664: dout <= 8'b00000000; // 1636 :   0 - 0x0
      11'h665: dout <= 8'b00000000; // 1637 :   0 - 0x0
      11'h666: dout <= 8'b00000000; // 1638 :   0 - 0x0
      11'h667: dout <= 8'b00000000; // 1639 :   0 - 0x0
      11'h668: dout <= 8'b00000000; // 1640 :   0 - 0x0 -- Sprite 0xcd
      11'h669: dout <= 8'b00000000; // 1641 :   0 - 0x0
      11'h66A: dout <= 8'b00000000; // 1642 :   0 - 0x0
      11'h66B: dout <= 8'b00000000; // 1643 :   0 - 0x0
      11'h66C: dout <= 8'b00000000; // 1644 :   0 - 0x0
      11'h66D: dout <= 8'b00000000; // 1645 :   0 - 0x0
      11'h66E: dout <= 8'b00000000; // 1646 :   0 - 0x0
      11'h66F: dout <= 8'b00000000; // 1647 :   0 - 0x0
      11'h670: dout <= 8'b00000000; // 1648 :   0 - 0x0 -- Sprite 0xce
      11'h671: dout <= 8'b00000000; // 1649 :   0 - 0x0
      11'h672: dout <= 8'b00000000; // 1650 :   0 - 0x0
      11'h673: dout <= 8'b00000000; // 1651 :   0 - 0x0
      11'h674: dout <= 8'b00000000; // 1652 :   0 - 0x0
      11'h675: dout <= 8'b00000000; // 1653 :   0 - 0x0
      11'h676: dout <= 8'b00000000; // 1654 :   0 - 0x0
      11'h677: dout <= 8'b00000000; // 1655 :   0 - 0x0
      11'h678: dout <= 8'b00000000; // 1656 :   0 - 0x0 -- Sprite 0xcf
      11'h679: dout <= 8'b00000000; // 1657 :   0 - 0x0
      11'h67A: dout <= 8'b00000000; // 1658 :   0 - 0x0
      11'h67B: dout <= 8'b00000000; // 1659 :   0 - 0x0
      11'h67C: dout <= 8'b00000000; // 1660 :   0 - 0x0
      11'h67D: dout <= 8'b00000000; // 1661 :   0 - 0x0
      11'h67E: dout <= 8'b00000000; // 1662 :   0 - 0x0
      11'h67F: dout <= 8'b00000000; // 1663 :   0 - 0x0
      11'h680: dout <= 8'b11111111; // 1664 : 255 - 0xff -- Sprite 0xd0
      11'h681: dout <= 8'b11111111; // 1665 : 255 - 0xff
      11'h682: dout <= 8'b11111111; // 1666 : 255 - 0xff
      11'h683: dout <= 8'b11111111; // 1667 : 255 - 0xff
      11'h684: dout <= 8'b11111111; // 1668 : 255 - 0xff
      11'h685: dout <= 8'b11111111; // 1669 : 255 - 0xff
      11'h686: dout <= 8'b11111111; // 1670 : 255 - 0xff
      11'h687: dout <= 8'b11111111; // 1671 : 255 - 0xff
      11'h688: dout <= 8'b11111111; // 1672 : 255 - 0xff -- Sprite 0xd1
      11'h689: dout <= 8'b11111111; // 1673 : 255 - 0xff
      11'h68A: dout <= 8'b11111111; // 1674 : 255 - 0xff
      11'h68B: dout <= 8'b11111111; // 1675 : 255 - 0xff
      11'h68C: dout <= 8'b11111111; // 1676 : 255 - 0xff
      11'h68D: dout <= 8'b11111111; // 1677 : 255 - 0xff
      11'h68E: dout <= 8'b11111111; // 1678 : 255 - 0xff
      11'h68F: dout <= 8'b11111111; // 1679 : 255 - 0xff
      11'h690: dout <= 8'b11111111; // 1680 : 255 - 0xff -- Sprite 0xd2
      11'h691: dout <= 8'b11111111; // 1681 : 255 - 0xff
      11'h692: dout <= 8'b11111111; // 1682 : 255 - 0xff
      11'h693: dout <= 8'b11111111; // 1683 : 255 - 0xff
      11'h694: dout <= 8'b11111111; // 1684 : 255 - 0xff
      11'h695: dout <= 8'b11111111; // 1685 : 255 - 0xff
      11'h696: dout <= 8'b11111111; // 1686 : 255 - 0xff
      11'h697: dout <= 8'b11111111; // 1687 : 255 - 0xff
      11'h698: dout <= 8'b11111111; // 1688 : 255 - 0xff -- Sprite 0xd3
      11'h699: dout <= 8'b11111111; // 1689 : 255 - 0xff
      11'h69A: dout <= 8'b11111111; // 1690 : 255 - 0xff
      11'h69B: dout <= 8'b11111111; // 1691 : 255 - 0xff
      11'h69C: dout <= 8'b11111111; // 1692 : 255 - 0xff
      11'h69D: dout <= 8'b11111111; // 1693 : 255 - 0xff
      11'h69E: dout <= 8'b11111111; // 1694 : 255 - 0xff
      11'h69F: dout <= 8'b11111111; // 1695 : 255 - 0xff
      11'h6A0: dout <= 8'b11111111; // 1696 : 255 - 0xff -- Sprite 0xd4
      11'h6A1: dout <= 8'b11111111; // 1697 : 255 - 0xff
      11'h6A2: dout <= 8'b11111111; // 1698 : 255 - 0xff
      11'h6A3: dout <= 8'b11111111; // 1699 : 255 - 0xff
      11'h6A4: dout <= 8'b11111111; // 1700 : 255 - 0xff
      11'h6A5: dout <= 8'b11111111; // 1701 : 255 - 0xff
      11'h6A6: dout <= 8'b11111111; // 1702 : 255 - 0xff
      11'h6A7: dout <= 8'b11111111; // 1703 : 255 - 0xff
      11'h6A8: dout <= 8'b11111111; // 1704 : 255 - 0xff -- Sprite 0xd5
      11'h6A9: dout <= 8'b11111111; // 1705 : 255 - 0xff
      11'h6AA: dout <= 8'b11111111; // 1706 : 255 - 0xff
      11'h6AB: dout <= 8'b11111111; // 1707 : 255 - 0xff
      11'h6AC: dout <= 8'b11111111; // 1708 : 255 - 0xff
      11'h6AD: dout <= 8'b11111111; // 1709 : 255 - 0xff
      11'h6AE: dout <= 8'b11111111; // 1710 : 255 - 0xff
      11'h6AF: dout <= 8'b11111111; // 1711 : 255 - 0xff
      11'h6B0: dout <= 8'b11111111; // 1712 : 255 - 0xff -- Sprite 0xd6
      11'h6B1: dout <= 8'b11111111; // 1713 : 255 - 0xff
      11'h6B2: dout <= 8'b11111111; // 1714 : 255 - 0xff
      11'h6B3: dout <= 8'b11111111; // 1715 : 255 - 0xff
      11'h6B4: dout <= 8'b11111111; // 1716 : 255 - 0xff
      11'h6B5: dout <= 8'b11111111; // 1717 : 255 - 0xff
      11'h6B6: dout <= 8'b11111111; // 1718 : 255 - 0xff
      11'h6B7: dout <= 8'b11111111; // 1719 : 255 - 0xff
      11'h6B8: dout <= 8'b11111111; // 1720 : 255 - 0xff -- Sprite 0xd7
      11'h6B9: dout <= 8'b11111111; // 1721 : 255 - 0xff
      11'h6BA: dout <= 8'b11111111; // 1722 : 255 - 0xff
      11'h6BB: dout <= 8'b11111111; // 1723 : 255 - 0xff
      11'h6BC: dout <= 8'b11111111; // 1724 : 255 - 0xff
      11'h6BD: dout <= 8'b11111111; // 1725 : 255 - 0xff
      11'h6BE: dout <= 8'b11111111; // 1726 : 255 - 0xff
      11'h6BF: dout <= 8'b11111111; // 1727 : 255 - 0xff
      11'h6C0: dout <= 8'b11111111; // 1728 : 255 - 0xff -- Sprite 0xd8
      11'h6C1: dout <= 8'b11111111; // 1729 : 255 - 0xff
      11'h6C2: dout <= 8'b11111111; // 1730 : 255 - 0xff
      11'h6C3: dout <= 8'b11111111; // 1731 : 255 - 0xff
      11'h6C4: dout <= 8'b11111111; // 1732 : 255 - 0xff
      11'h6C5: dout <= 8'b11111111; // 1733 : 255 - 0xff
      11'h6C6: dout <= 8'b11111111; // 1734 : 255 - 0xff
      11'h6C7: dout <= 8'b11111111; // 1735 : 255 - 0xff
      11'h6C8: dout <= 8'b11111111; // 1736 : 255 - 0xff -- Sprite 0xd9
      11'h6C9: dout <= 8'b11111111; // 1737 : 255 - 0xff
      11'h6CA: dout <= 8'b11111111; // 1738 : 255 - 0xff
      11'h6CB: dout <= 8'b11111111; // 1739 : 255 - 0xff
      11'h6CC: dout <= 8'b11111111; // 1740 : 255 - 0xff
      11'h6CD: dout <= 8'b11111111; // 1741 : 255 - 0xff
      11'h6CE: dout <= 8'b11111111; // 1742 : 255 - 0xff
      11'h6CF: dout <= 8'b11111111; // 1743 : 255 - 0xff
      11'h6D0: dout <= 8'b11111111; // 1744 : 255 - 0xff -- Sprite 0xda
      11'h6D1: dout <= 8'b11111111; // 1745 : 255 - 0xff
      11'h6D2: dout <= 8'b11111111; // 1746 : 255 - 0xff
      11'h6D3: dout <= 8'b11111111; // 1747 : 255 - 0xff
      11'h6D4: dout <= 8'b11111111; // 1748 : 255 - 0xff
      11'h6D5: dout <= 8'b11111111; // 1749 : 255 - 0xff
      11'h6D6: dout <= 8'b11111111; // 1750 : 255 - 0xff
      11'h6D7: dout <= 8'b11111111; // 1751 : 255 - 0xff
      11'h6D8: dout <= 8'b11111111; // 1752 : 255 - 0xff -- Sprite 0xdb
      11'h6D9: dout <= 8'b11111111; // 1753 : 255 - 0xff
      11'h6DA: dout <= 8'b11111111; // 1754 : 255 - 0xff
      11'h6DB: dout <= 8'b11111111; // 1755 : 255 - 0xff
      11'h6DC: dout <= 8'b11111111; // 1756 : 255 - 0xff
      11'h6DD: dout <= 8'b11111111; // 1757 : 255 - 0xff
      11'h6DE: dout <= 8'b11111111; // 1758 : 255 - 0xff
      11'h6DF: dout <= 8'b11111111; // 1759 : 255 - 0xff
      11'h6E0: dout <= 8'b11111111; // 1760 : 255 - 0xff -- Sprite 0xdc
      11'h6E1: dout <= 8'b11111111; // 1761 : 255 - 0xff
      11'h6E2: dout <= 8'b11111111; // 1762 : 255 - 0xff
      11'h6E3: dout <= 8'b11111111; // 1763 : 255 - 0xff
      11'h6E4: dout <= 8'b11111111; // 1764 : 255 - 0xff
      11'h6E5: dout <= 8'b11111111; // 1765 : 255 - 0xff
      11'h6E6: dout <= 8'b11111111; // 1766 : 255 - 0xff
      11'h6E7: dout <= 8'b11111111; // 1767 : 255 - 0xff
      11'h6E8: dout <= 8'b11111111; // 1768 : 255 - 0xff -- Sprite 0xdd
      11'h6E9: dout <= 8'b11111111; // 1769 : 255 - 0xff
      11'h6EA: dout <= 8'b11111111; // 1770 : 255 - 0xff
      11'h6EB: dout <= 8'b11111111; // 1771 : 255 - 0xff
      11'h6EC: dout <= 8'b11111111; // 1772 : 255 - 0xff
      11'h6ED: dout <= 8'b11111111; // 1773 : 255 - 0xff
      11'h6EE: dout <= 8'b11111111; // 1774 : 255 - 0xff
      11'h6EF: dout <= 8'b11111111; // 1775 : 255 - 0xff
      11'h6F0: dout <= 8'b11111111; // 1776 : 255 - 0xff -- Sprite 0xde
      11'h6F1: dout <= 8'b11111111; // 1777 : 255 - 0xff
      11'h6F2: dout <= 8'b11111111; // 1778 : 255 - 0xff
      11'h6F3: dout <= 8'b11111111; // 1779 : 255 - 0xff
      11'h6F4: dout <= 8'b11111111; // 1780 : 255 - 0xff
      11'h6F5: dout <= 8'b11111111; // 1781 : 255 - 0xff
      11'h6F6: dout <= 8'b11111111; // 1782 : 255 - 0xff
      11'h6F7: dout <= 8'b11111111; // 1783 : 255 - 0xff
      11'h6F8: dout <= 8'b11111111; // 1784 : 255 - 0xff -- Sprite 0xdf
      11'h6F9: dout <= 8'b11111111; // 1785 : 255 - 0xff
      11'h6FA: dout <= 8'b11111111; // 1786 : 255 - 0xff
      11'h6FB: dout <= 8'b11111111; // 1787 : 255 - 0xff
      11'h6FC: dout <= 8'b11111111; // 1788 : 255 - 0xff
      11'h6FD: dout <= 8'b11111111; // 1789 : 255 - 0xff
      11'h6FE: dout <= 8'b11111111; // 1790 : 255 - 0xff
      11'h6FF: dout <= 8'b11111111; // 1791 : 255 - 0xff
      11'h700: dout <= 8'b11111111; // 1792 : 255 - 0xff -- Sprite 0xe0
      11'h701: dout <= 8'b11111111; // 1793 : 255 - 0xff
      11'h702: dout <= 8'b11111111; // 1794 : 255 - 0xff
      11'h703: dout <= 8'b11111111; // 1795 : 255 - 0xff
      11'h704: dout <= 8'b11111111; // 1796 : 255 - 0xff
      11'h705: dout <= 8'b11111111; // 1797 : 255 - 0xff
      11'h706: dout <= 8'b11111111; // 1798 : 255 - 0xff
      11'h707: dout <= 8'b11111111; // 1799 : 255 - 0xff
      11'h708: dout <= 8'b11111111; // 1800 : 255 - 0xff -- Sprite 0xe1
      11'h709: dout <= 8'b11111111; // 1801 : 255 - 0xff
      11'h70A: dout <= 8'b11111111; // 1802 : 255 - 0xff
      11'h70B: dout <= 8'b11111111; // 1803 : 255 - 0xff
      11'h70C: dout <= 8'b11111111; // 1804 : 255 - 0xff
      11'h70D: dout <= 8'b11111111; // 1805 : 255 - 0xff
      11'h70E: dout <= 8'b11111111; // 1806 : 255 - 0xff
      11'h70F: dout <= 8'b11111111; // 1807 : 255 - 0xff
      11'h710: dout <= 8'b11111111; // 1808 : 255 - 0xff -- Sprite 0xe2
      11'h711: dout <= 8'b11111111; // 1809 : 255 - 0xff
      11'h712: dout <= 8'b11111111; // 1810 : 255 - 0xff
      11'h713: dout <= 8'b11111111; // 1811 : 255 - 0xff
      11'h714: dout <= 8'b11111111; // 1812 : 255 - 0xff
      11'h715: dout <= 8'b11111111; // 1813 : 255 - 0xff
      11'h716: dout <= 8'b11111111; // 1814 : 255 - 0xff
      11'h717: dout <= 8'b11111111; // 1815 : 255 - 0xff
      11'h718: dout <= 8'b11111111; // 1816 : 255 - 0xff -- Sprite 0xe3
      11'h719: dout <= 8'b11111111; // 1817 : 255 - 0xff
      11'h71A: dout <= 8'b11111111; // 1818 : 255 - 0xff
      11'h71B: dout <= 8'b11111111; // 1819 : 255 - 0xff
      11'h71C: dout <= 8'b11111111; // 1820 : 255 - 0xff
      11'h71D: dout <= 8'b11111111; // 1821 : 255 - 0xff
      11'h71E: dout <= 8'b11111111; // 1822 : 255 - 0xff
      11'h71F: dout <= 8'b11111111; // 1823 : 255 - 0xff
      11'h720: dout <= 8'b11111111; // 1824 : 255 - 0xff -- Sprite 0xe4
      11'h721: dout <= 8'b11111111; // 1825 : 255 - 0xff
      11'h722: dout <= 8'b11111111; // 1826 : 255 - 0xff
      11'h723: dout <= 8'b11111111; // 1827 : 255 - 0xff
      11'h724: dout <= 8'b11111111; // 1828 : 255 - 0xff
      11'h725: dout <= 8'b11111111; // 1829 : 255 - 0xff
      11'h726: dout <= 8'b11111111; // 1830 : 255 - 0xff
      11'h727: dout <= 8'b11111111; // 1831 : 255 - 0xff
      11'h728: dout <= 8'b11111111; // 1832 : 255 - 0xff -- Sprite 0xe5
      11'h729: dout <= 8'b11111111; // 1833 : 255 - 0xff
      11'h72A: dout <= 8'b11111111; // 1834 : 255 - 0xff
      11'h72B: dout <= 8'b11111111; // 1835 : 255 - 0xff
      11'h72C: dout <= 8'b11111111; // 1836 : 255 - 0xff
      11'h72D: dout <= 8'b11111111; // 1837 : 255 - 0xff
      11'h72E: dout <= 8'b11111111; // 1838 : 255 - 0xff
      11'h72F: dout <= 8'b11111111; // 1839 : 255 - 0xff
      11'h730: dout <= 8'b11111111; // 1840 : 255 - 0xff -- Sprite 0xe6
      11'h731: dout <= 8'b11111111; // 1841 : 255 - 0xff
      11'h732: dout <= 8'b11111111; // 1842 : 255 - 0xff
      11'h733: dout <= 8'b11111111; // 1843 : 255 - 0xff
      11'h734: dout <= 8'b11111111; // 1844 : 255 - 0xff
      11'h735: dout <= 8'b11111111; // 1845 : 255 - 0xff
      11'h736: dout <= 8'b11111111; // 1846 : 255 - 0xff
      11'h737: dout <= 8'b11111111; // 1847 : 255 - 0xff
      11'h738: dout <= 8'b11111111; // 1848 : 255 - 0xff -- Sprite 0xe7
      11'h739: dout <= 8'b11111111; // 1849 : 255 - 0xff
      11'h73A: dout <= 8'b11111111; // 1850 : 255 - 0xff
      11'h73B: dout <= 8'b11111111; // 1851 : 255 - 0xff
      11'h73C: dout <= 8'b11111111; // 1852 : 255 - 0xff
      11'h73D: dout <= 8'b11111111; // 1853 : 255 - 0xff
      11'h73E: dout <= 8'b11111111; // 1854 : 255 - 0xff
      11'h73F: dout <= 8'b11111111; // 1855 : 255 - 0xff
      11'h740: dout <= 8'b11111111; // 1856 : 255 - 0xff -- Sprite 0xe8
      11'h741: dout <= 8'b11111111; // 1857 : 255 - 0xff
      11'h742: dout <= 8'b11111111; // 1858 : 255 - 0xff
      11'h743: dout <= 8'b11111111; // 1859 : 255 - 0xff
      11'h744: dout <= 8'b11111111; // 1860 : 255 - 0xff
      11'h745: dout <= 8'b11111111; // 1861 : 255 - 0xff
      11'h746: dout <= 8'b11111111; // 1862 : 255 - 0xff
      11'h747: dout <= 8'b11111111; // 1863 : 255 - 0xff
      11'h748: dout <= 8'b11111111; // 1864 : 255 - 0xff -- Sprite 0xe9
      11'h749: dout <= 8'b11111111; // 1865 : 255 - 0xff
      11'h74A: dout <= 8'b11111111; // 1866 : 255 - 0xff
      11'h74B: dout <= 8'b11111111; // 1867 : 255 - 0xff
      11'h74C: dout <= 8'b11111111; // 1868 : 255 - 0xff
      11'h74D: dout <= 8'b11111111; // 1869 : 255 - 0xff
      11'h74E: dout <= 8'b11111111; // 1870 : 255 - 0xff
      11'h74F: dout <= 8'b11111111; // 1871 : 255 - 0xff
      11'h750: dout <= 8'b11111111; // 1872 : 255 - 0xff -- Sprite 0xea
      11'h751: dout <= 8'b11111111; // 1873 : 255 - 0xff
      11'h752: dout <= 8'b11111111; // 1874 : 255 - 0xff
      11'h753: dout <= 8'b11111111; // 1875 : 255 - 0xff
      11'h754: dout <= 8'b11111111; // 1876 : 255 - 0xff
      11'h755: dout <= 8'b11111111; // 1877 : 255 - 0xff
      11'h756: dout <= 8'b11111111; // 1878 : 255 - 0xff
      11'h757: dout <= 8'b11111111; // 1879 : 255 - 0xff
      11'h758: dout <= 8'b11111111; // 1880 : 255 - 0xff -- Sprite 0xeb
      11'h759: dout <= 8'b11111111; // 1881 : 255 - 0xff
      11'h75A: dout <= 8'b11111111; // 1882 : 255 - 0xff
      11'h75B: dout <= 8'b11111111; // 1883 : 255 - 0xff
      11'h75C: dout <= 8'b11111111; // 1884 : 255 - 0xff
      11'h75D: dout <= 8'b11111111; // 1885 : 255 - 0xff
      11'h75E: dout <= 8'b11111111; // 1886 : 255 - 0xff
      11'h75F: dout <= 8'b11111111; // 1887 : 255 - 0xff
      11'h760: dout <= 8'b11111111; // 1888 : 255 - 0xff -- Sprite 0xec
      11'h761: dout <= 8'b11111111; // 1889 : 255 - 0xff
      11'h762: dout <= 8'b11111111; // 1890 : 255 - 0xff
      11'h763: dout <= 8'b11111111; // 1891 : 255 - 0xff
      11'h764: dout <= 8'b11111111; // 1892 : 255 - 0xff
      11'h765: dout <= 8'b11111111; // 1893 : 255 - 0xff
      11'h766: dout <= 8'b11111111; // 1894 : 255 - 0xff
      11'h767: dout <= 8'b11111111; // 1895 : 255 - 0xff
      11'h768: dout <= 8'b11111111; // 1896 : 255 - 0xff -- Sprite 0xed
      11'h769: dout <= 8'b11111111; // 1897 : 255 - 0xff
      11'h76A: dout <= 8'b11111111; // 1898 : 255 - 0xff
      11'h76B: dout <= 8'b11111111; // 1899 : 255 - 0xff
      11'h76C: dout <= 8'b11111111; // 1900 : 255 - 0xff
      11'h76D: dout <= 8'b11111111; // 1901 : 255 - 0xff
      11'h76E: dout <= 8'b11111111; // 1902 : 255 - 0xff
      11'h76F: dout <= 8'b11111111; // 1903 : 255 - 0xff
      11'h770: dout <= 8'b11111111; // 1904 : 255 - 0xff -- Sprite 0xee
      11'h771: dout <= 8'b11111111; // 1905 : 255 - 0xff
      11'h772: dout <= 8'b11111111; // 1906 : 255 - 0xff
      11'h773: dout <= 8'b11111111; // 1907 : 255 - 0xff
      11'h774: dout <= 8'b11111111; // 1908 : 255 - 0xff
      11'h775: dout <= 8'b11111111; // 1909 : 255 - 0xff
      11'h776: dout <= 8'b11111111; // 1910 : 255 - 0xff
      11'h777: dout <= 8'b11111111; // 1911 : 255 - 0xff
      11'h778: dout <= 8'b11111111; // 1912 : 255 - 0xff -- Sprite 0xef
      11'h779: dout <= 8'b11111111; // 1913 : 255 - 0xff
      11'h77A: dout <= 8'b11111111; // 1914 : 255 - 0xff
      11'h77B: dout <= 8'b11111111; // 1915 : 255 - 0xff
      11'h77C: dout <= 8'b11111111; // 1916 : 255 - 0xff
      11'h77D: dout <= 8'b11111111; // 1917 : 255 - 0xff
      11'h77E: dout <= 8'b11111111; // 1918 : 255 - 0xff
      11'h77F: dout <= 8'b11111111; // 1919 : 255 - 0xff
      11'h780: dout <= 8'b11111111; // 1920 : 255 - 0xff -- Sprite 0xf0
      11'h781: dout <= 8'b11111111; // 1921 : 255 - 0xff
      11'h782: dout <= 8'b11111111; // 1922 : 255 - 0xff
      11'h783: dout <= 8'b11111111; // 1923 : 255 - 0xff
      11'h784: dout <= 8'b11111111; // 1924 : 255 - 0xff
      11'h785: dout <= 8'b11111111; // 1925 : 255 - 0xff
      11'h786: dout <= 8'b11111111; // 1926 : 255 - 0xff
      11'h787: dout <= 8'b11111111; // 1927 : 255 - 0xff
      11'h788: dout <= 8'b11111111; // 1928 : 255 - 0xff -- Sprite 0xf1
      11'h789: dout <= 8'b11111111; // 1929 : 255 - 0xff
      11'h78A: dout <= 8'b11111111; // 1930 : 255 - 0xff
      11'h78B: dout <= 8'b11111111; // 1931 : 255 - 0xff
      11'h78C: dout <= 8'b11111111; // 1932 : 255 - 0xff
      11'h78D: dout <= 8'b11111111; // 1933 : 255 - 0xff
      11'h78E: dout <= 8'b11111111; // 1934 : 255 - 0xff
      11'h78F: dout <= 8'b11111111; // 1935 : 255 - 0xff
      11'h790: dout <= 8'b11111111; // 1936 : 255 - 0xff -- Sprite 0xf2
      11'h791: dout <= 8'b11111111; // 1937 : 255 - 0xff
      11'h792: dout <= 8'b11111111; // 1938 : 255 - 0xff
      11'h793: dout <= 8'b11111111; // 1939 : 255 - 0xff
      11'h794: dout <= 8'b11111111; // 1940 : 255 - 0xff
      11'h795: dout <= 8'b11111111; // 1941 : 255 - 0xff
      11'h796: dout <= 8'b11111111; // 1942 : 255 - 0xff
      11'h797: dout <= 8'b11111111; // 1943 : 255 - 0xff
      11'h798: dout <= 8'b11111111; // 1944 : 255 - 0xff -- Sprite 0xf3
      11'h799: dout <= 8'b11111111; // 1945 : 255 - 0xff
      11'h79A: dout <= 8'b11111111; // 1946 : 255 - 0xff
      11'h79B: dout <= 8'b11111111; // 1947 : 255 - 0xff
      11'h79C: dout <= 8'b11111111; // 1948 : 255 - 0xff
      11'h79D: dout <= 8'b11111111; // 1949 : 255 - 0xff
      11'h79E: dout <= 8'b11111111; // 1950 : 255 - 0xff
      11'h79F: dout <= 8'b11111111; // 1951 : 255 - 0xff
      11'h7A0: dout <= 8'b11111111; // 1952 : 255 - 0xff -- Sprite 0xf4
      11'h7A1: dout <= 8'b11111111; // 1953 : 255 - 0xff
      11'h7A2: dout <= 8'b11111111; // 1954 : 255 - 0xff
      11'h7A3: dout <= 8'b11111111; // 1955 : 255 - 0xff
      11'h7A4: dout <= 8'b11111111; // 1956 : 255 - 0xff
      11'h7A5: dout <= 8'b11111111; // 1957 : 255 - 0xff
      11'h7A6: dout <= 8'b11111111; // 1958 : 255 - 0xff
      11'h7A7: dout <= 8'b11111111; // 1959 : 255 - 0xff
      11'h7A8: dout <= 8'b11111111; // 1960 : 255 - 0xff -- Sprite 0xf5
      11'h7A9: dout <= 8'b11111111; // 1961 : 255 - 0xff
      11'h7AA: dout <= 8'b11111111; // 1962 : 255 - 0xff
      11'h7AB: dout <= 8'b11111111; // 1963 : 255 - 0xff
      11'h7AC: dout <= 8'b11111111; // 1964 : 255 - 0xff
      11'h7AD: dout <= 8'b11111111; // 1965 : 255 - 0xff
      11'h7AE: dout <= 8'b11111111; // 1966 : 255 - 0xff
      11'h7AF: dout <= 8'b11111111; // 1967 : 255 - 0xff
      11'h7B0: dout <= 8'b11111111; // 1968 : 255 - 0xff -- Sprite 0xf6
      11'h7B1: dout <= 8'b11111111; // 1969 : 255 - 0xff
      11'h7B2: dout <= 8'b11111111; // 1970 : 255 - 0xff
      11'h7B3: dout <= 8'b11111111; // 1971 : 255 - 0xff
      11'h7B4: dout <= 8'b11111111; // 1972 : 255 - 0xff
      11'h7B5: dout <= 8'b11111111; // 1973 : 255 - 0xff
      11'h7B6: dout <= 8'b11111111; // 1974 : 255 - 0xff
      11'h7B7: dout <= 8'b11111111; // 1975 : 255 - 0xff
      11'h7B8: dout <= 8'b11111111; // 1976 : 255 - 0xff -- Sprite 0xf7
      11'h7B9: dout <= 8'b11111111; // 1977 : 255 - 0xff
      11'h7BA: dout <= 8'b11111111; // 1978 : 255 - 0xff
      11'h7BB: dout <= 8'b11111111; // 1979 : 255 - 0xff
      11'h7BC: dout <= 8'b11111111; // 1980 : 255 - 0xff
      11'h7BD: dout <= 8'b11111111; // 1981 : 255 - 0xff
      11'h7BE: dout <= 8'b11111111; // 1982 : 255 - 0xff
      11'h7BF: dout <= 8'b11111111; // 1983 : 255 - 0xff
      11'h7C0: dout <= 8'b11111111; // 1984 : 255 - 0xff -- Sprite 0xf8
      11'h7C1: dout <= 8'b11111111; // 1985 : 255 - 0xff
      11'h7C2: dout <= 8'b11111111; // 1986 : 255 - 0xff
      11'h7C3: dout <= 8'b11111111; // 1987 : 255 - 0xff
      11'h7C4: dout <= 8'b11111111; // 1988 : 255 - 0xff
      11'h7C5: dout <= 8'b11111111; // 1989 : 255 - 0xff
      11'h7C6: dout <= 8'b11111111; // 1990 : 255 - 0xff
      11'h7C7: dout <= 8'b11111111; // 1991 : 255 - 0xff
      11'h7C8: dout <= 8'b11111111; // 1992 : 255 - 0xff -- Sprite 0xf9
      11'h7C9: dout <= 8'b11111111; // 1993 : 255 - 0xff
      11'h7CA: dout <= 8'b11111111; // 1994 : 255 - 0xff
      11'h7CB: dout <= 8'b11111111; // 1995 : 255 - 0xff
      11'h7CC: dout <= 8'b11111111; // 1996 : 255 - 0xff
      11'h7CD: dout <= 8'b11111111; // 1997 : 255 - 0xff
      11'h7CE: dout <= 8'b11111111; // 1998 : 255 - 0xff
      11'h7CF: dout <= 8'b11111111; // 1999 : 255 - 0xff
      11'h7D0: dout <= 8'b11111111; // 2000 : 255 - 0xff -- Sprite 0xfa
      11'h7D1: dout <= 8'b11111111; // 2001 : 255 - 0xff
      11'h7D2: dout <= 8'b11111111; // 2002 : 255 - 0xff
      11'h7D3: dout <= 8'b11111111; // 2003 : 255 - 0xff
      11'h7D4: dout <= 8'b11111111; // 2004 : 255 - 0xff
      11'h7D5: dout <= 8'b11111111; // 2005 : 255 - 0xff
      11'h7D6: dout <= 8'b11111111; // 2006 : 255 - 0xff
      11'h7D7: dout <= 8'b11111111; // 2007 : 255 - 0xff
      11'h7D8: dout <= 8'b11111111; // 2008 : 255 - 0xff -- Sprite 0xfb
      11'h7D9: dout <= 8'b11111111; // 2009 : 255 - 0xff
      11'h7DA: dout <= 8'b11111111; // 2010 : 255 - 0xff
      11'h7DB: dout <= 8'b11111111; // 2011 : 255 - 0xff
      11'h7DC: dout <= 8'b11111111; // 2012 : 255 - 0xff
      11'h7DD: dout <= 8'b11111111; // 2013 : 255 - 0xff
      11'h7DE: dout <= 8'b11111111; // 2014 : 255 - 0xff
      11'h7DF: dout <= 8'b11111111; // 2015 : 255 - 0xff
      11'h7E0: dout <= 8'b11111111; // 2016 : 255 - 0xff -- Sprite 0xfc
      11'h7E1: dout <= 8'b11111111; // 2017 : 255 - 0xff
      11'h7E2: dout <= 8'b11111111; // 2018 : 255 - 0xff
      11'h7E3: dout <= 8'b11111111; // 2019 : 255 - 0xff
      11'h7E4: dout <= 8'b11111111; // 2020 : 255 - 0xff
      11'h7E5: dout <= 8'b11111111; // 2021 : 255 - 0xff
      11'h7E6: dout <= 8'b11111111; // 2022 : 255 - 0xff
      11'h7E7: dout <= 8'b11111111; // 2023 : 255 - 0xff
      11'h7E8: dout <= 8'b11111111; // 2024 : 255 - 0xff -- Sprite 0xfd
      11'h7E9: dout <= 8'b11111111; // 2025 : 255 - 0xff
      11'h7EA: dout <= 8'b11111111; // 2026 : 255 - 0xff
      11'h7EB: dout <= 8'b11111111; // 2027 : 255 - 0xff
      11'h7EC: dout <= 8'b11111111; // 2028 : 255 - 0xff
      11'h7ED: dout <= 8'b11111111; // 2029 : 255 - 0xff
      11'h7EE: dout <= 8'b11111111; // 2030 : 255 - 0xff
      11'h7EF: dout <= 8'b11111111; // 2031 : 255 - 0xff
      11'h7F0: dout <= 8'b11111111; // 2032 : 255 - 0xff -- Sprite 0xfe
      11'h7F1: dout <= 8'b11111111; // 2033 : 255 - 0xff
      11'h7F2: dout <= 8'b11111111; // 2034 : 255 - 0xff
      11'h7F3: dout <= 8'b11111111; // 2035 : 255 - 0xff
      11'h7F4: dout <= 8'b11111111; // 2036 : 255 - 0xff
      11'h7F5: dout <= 8'b11111111; // 2037 : 255 - 0xff
      11'h7F6: dout <= 8'b11111111; // 2038 : 255 - 0xff
      11'h7F7: dout <= 8'b11111111; // 2039 : 255 - 0xff
      11'h7F8: dout <= 8'b11111111; // 2040 : 255 - 0xff -- Sprite 0xff
      11'h7F9: dout <= 8'b11111111; // 2041 : 255 - 0xff
      11'h7FA: dout <= 8'b11111111; // 2042 : 255 - 0xff
      11'h7FB: dout <= 8'b11111111; // 2043 : 255 - 0xff
      11'h7FC: dout <= 8'b11111111; // 2044 : 255 - 0xff
      11'h7FD: dout <= 8'b11111111; // 2045 : 255 - 0xff
      11'h7FE: dout <= 8'b11111111; // 2046 : 255 - 0xff
      11'h7FF: dout <= 8'b11111111; // 2047 : 255 - 0xff
    endcase
  end

endmodule
