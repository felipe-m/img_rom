------- ROM creada automaticamente por ppm2rom -----------
------- Felipe Machado -----------------------------------
------- Departamento de Tecnologia Electronica -----------
------- Universidad Rey Juan Carlos ----------------------
------- http://gtebim.es ---------------------------------
----------------------------------------------------------
--------Datos de la imagen -------------------------------
--- Fichero original    : hor_ver_128.pgm 
--- Filas    : 128 
--- Columnas : 128 
--- Color    :  8 bits



------ Puertos -------------------------------------------
-- Entradas ----------------------------------------------
--    clk  :  senal de reloj
--    addr :  direccion de la memoria
-- Salidas  ----------------------------------------------
--    dout :  dato de 8 bits de la direccion addr (un ciclo despues)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM8b_hor_ver_128 is
  port (
    clk  : in  std_logic;   -- reloj
    addr : in  std_logic_vector(14-1 downto 0);
    dout : out std_logic_vector(8-1 downto 0) 
  );
end ROM8b_hor_ver_128;


architecture BEHAVIORAL of ROM8b_hor_ver_128 is
  signal addr_int  : natural range 0 to 2**14-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant filaimg : memostruct := (
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010011",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "01010011",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "01010010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "00000110",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11010011",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "00000010",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "01000111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "10001101",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "00000001",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "01110111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "11111111",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000",
       "00000000"
        );

begin

  addr_int <= TO_INTEGER(unsigned(addr));

  P_ROM: process (clk)
  begin
    if clk'event and clk='1' then
      dout <= filaimg(addr_int);
    end if;
  end process;

end BEHAVIORAL;

