//- Autcmatically generated verilog ROM from a NES memory file----
//-   PATTERN TABLE WITH ONLY ONE COLOR PLANE
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables


//-  Original memory dump file name: nova_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_PTABLE_NOVA_color1
  (
     input     clk,   // clock
     input      [12-1:0] addr,  //4096 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                              //  address:   value 
                              //    dec  : dec - hex
          // Sprite pattern Table
      12'h0: dout <= 8'b00000000; //    0 :   0 - 0x0 -- Sprite 0x0
      12'h1: dout <= 8'b01111111; //    1 : 127 - 0x7f
      12'h2: dout <= 8'b01111111; //    2 : 127 - 0x7f
      12'h3: dout <= 8'b01111111; //    3 : 127 - 0x7f
      12'h4: dout <= 8'b01111111; //    4 : 127 - 0x7f
      12'h5: dout <= 8'b01111111; //    5 : 127 - 0x7f
      12'h6: dout <= 8'b01101010; //    6 : 106 - 0x6a
      12'h7: dout <= 8'b00000000; //    7 :   0 - 0x0
      12'h8: dout <= 8'b00000000; //    8 :   0 - 0x0 -- Sprite 0x1
      12'h9: dout <= 8'b01111011; //    9 : 123 - 0x7b
      12'hA: dout <= 8'b01110011; //   10 : 115 - 0x73
      12'hB: dout <= 8'b01111011; //   11 : 123 - 0x7b
      12'hC: dout <= 8'b01110011; //   12 : 115 - 0x73
      12'hD: dout <= 8'b01111011; //   13 : 123 - 0x7b
      12'hE: dout <= 8'b01010011; //   14 :  83 - 0x53
      12'hF: dout <= 8'b00000000; //   15 :   0 - 0x0
      12'h10: dout <= 8'b00000000; //   16 :   0 - 0x0 -- Sprite 0x2
      12'h11: dout <= 8'b11011110; //   17 : 222 - 0xde
      12'h12: dout <= 8'b10011110; //   18 : 158 - 0x9e
      12'h13: dout <= 8'b11011100; //   19 : 220 - 0xdc
      12'h14: dout <= 8'b10011110; //   20 : 158 - 0x9e
      12'h15: dout <= 8'b11011100; //   21 : 220 - 0xdc
      12'h16: dout <= 8'b10011010; //   22 : 154 - 0x9a
      12'h17: dout <= 8'b00000000; //   23 :   0 - 0x0
      12'h18: dout <= 8'b00000000; //   24 :   0 - 0x0 -- Sprite 0x3
      12'h19: dout <= 8'b11111110; //   25 : 254 - 0xfe
      12'h1A: dout <= 8'b11111100; //   26 : 252 - 0xfc
      12'h1B: dout <= 8'b11111110; //   27 : 254 - 0xfe
      12'h1C: dout <= 8'b11111100; //   28 : 252 - 0xfc
      12'h1D: dout <= 8'b11111110; //   29 : 254 - 0xfe
      12'h1E: dout <= 8'b01010100; //   30 :  84 - 0x54
      12'h1F: dout <= 8'b00000000; //   31 :   0 - 0x0
      12'h20: dout <= 8'b00000000; //   32 :   0 - 0x0 -- Sprite 0x4
      12'h21: dout <= 8'b01111111; //   33 : 127 - 0x7f
      12'h22: dout <= 8'b01011111; //   34 :  95 - 0x5f
      12'h23: dout <= 8'b01111001; //   35 : 121 - 0x79
      12'h24: dout <= 8'b01111001; //   36 : 121 - 0x79
      12'h25: dout <= 8'b01001001; //   37 :  73 - 0x49
      12'h26: dout <= 8'b01001111; //   38 :  79 - 0x4f
      12'h27: dout <= 8'b01001110; //   39 :  78 - 0x4e
      12'h28: dout <= 8'b01111000; //   40 : 120 - 0x78 -- Sprite 0x5
      12'h29: dout <= 8'b01110000; //   41 : 112 - 0x70
      12'h2A: dout <= 8'b01100000; //   42 :  96 - 0x60
      12'h2B: dout <= 8'b01100000; //   43 :  96 - 0x60
      12'h2C: dout <= 8'b01110001; //   44 : 113 - 0x71
      12'h2D: dout <= 8'b01011111; //   45 :  95 - 0x5f
      12'h2E: dout <= 8'b01111111; //   46 : 127 - 0x7f
      12'h2F: dout <= 8'b00000000; //   47 :   0 - 0x0
      12'h30: dout <= 8'b00000000; //   48 :   0 - 0x0 -- Sprite 0x6
      12'h31: dout <= 8'b11111110; //   49 : 254 - 0xfe
      12'h32: dout <= 8'b11111010; //   50 : 250 - 0xfa
      12'h33: dout <= 8'b10011110; //   51 : 158 - 0x9e
      12'h34: dout <= 8'b10011110; //   52 : 158 - 0x9e
      12'h35: dout <= 8'b10010010; //   53 : 146 - 0x92
      12'h36: dout <= 8'b11110010; //   54 : 242 - 0xf2
      12'h37: dout <= 8'b01110010; //   55 : 114 - 0x72
      12'h38: dout <= 8'b00011110; //   56 :  30 - 0x1e -- Sprite 0x7
      12'h39: dout <= 8'b00001110; //   57 :  14 - 0xe
      12'h3A: dout <= 8'b00000110; //   58 :   6 - 0x6
      12'h3B: dout <= 8'b00000110; //   59 :   6 - 0x6
      12'h3C: dout <= 8'b10001110; //   60 : 142 - 0x8e
      12'h3D: dout <= 8'b11111010; //   61 : 250 - 0xfa
      12'h3E: dout <= 8'b11111110; //   62 : 254 - 0xfe
      12'h3F: dout <= 8'b00000000; //   63 :   0 - 0x0
      12'h40: dout <= 8'b00000000; //   64 :   0 - 0x0 -- Sprite 0x8
      12'h41: dout <= 8'b01111111; //   65 : 127 - 0x7f
      12'h42: dout <= 8'b01011111; //   66 :  95 - 0x5f
      12'h43: dout <= 8'b01111111; //   67 : 127 - 0x7f
      12'h44: dout <= 8'b01111111; //   68 : 127 - 0x7f
      12'h45: dout <= 8'b01111111; //   69 : 127 - 0x7f
      12'h46: dout <= 8'b01111111; //   70 : 127 - 0x7f
      12'h47: dout <= 8'b01111111; //   71 : 127 - 0x7f
      12'h48: dout <= 8'b01111111; //   72 : 127 - 0x7f -- Sprite 0x9
      12'h49: dout <= 8'b01111111; //   73 : 127 - 0x7f
      12'h4A: dout <= 8'b01111111; //   74 : 127 - 0x7f
      12'h4B: dout <= 8'b01111111; //   75 : 127 - 0x7f
      12'h4C: dout <= 8'b01111111; //   76 : 127 - 0x7f
      12'h4D: dout <= 8'b01011111; //   77 :  95 - 0x5f
      12'h4E: dout <= 8'b01111111; //   78 : 127 - 0x7f
      12'h4F: dout <= 8'b00000000; //   79 :   0 - 0x0
      12'h50: dout <= 8'b00000000; //   80 :   0 - 0x0 -- Sprite 0xa
      12'h51: dout <= 8'b11111110; //   81 : 254 - 0xfe
      12'h52: dout <= 8'b11111010; //   82 : 250 - 0xfa
      12'h53: dout <= 8'b11111110; //   83 : 254 - 0xfe
      12'h54: dout <= 8'b11111110; //   84 : 254 - 0xfe
      12'h55: dout <= 8'b11111110; //   85 : 254 - 0xfe
      12'h56: dout <= 8'b11111110; //   86 : 254 - 0xfe
      12'h57: dout <= 8'b11111110; //   87 : 254 - 0xfe
      12'h58: dout <= 8'b11111110; //   88 : 254 - 0xfe -- Sprite 0xb
      12'h59: dout <= 8'b11111110; //   89 : 254 - 0xfe
      12'h5A: dout <= 8'b11111110; //   90 : 254 - 0xfe
      12'h5B: dout <= 8'b11111110; //   91 : 254 - 0xfe
      12'h5C: dout <= 8'b11111110; //   92 : 254 - 0xfe
      12'h5D: dout <= 8'b11111010; //   93 : 250 - 0xfa
      12'h5E: dout <= 8'b11111110; //   94 : 254 - 0xfe
      12'h5F: dout <= 8'b00000000; //   95 :   0 - 0x0
      12'h60: dout <= 8'b00000000; //   96 :   0 - 0x0 -- Sprite 0xc
      12'h61: dout <= 8'b00111111; //   97 :  63 - 0x3f
      12'h62: dout <= 8'b01011111; //   98 :  95 - 0x5f
      12'h63: dout <= 8'b01101111; //   99 : 111 - 0x6f
      12'h64: dout <= 8'b01110000; //  100 : 112 - 0x70
      12'h65: dout <= 8'b01110111; //  101 : 119 - 0x77
      12'h66: dout <= 8'b01110111; //  102 : 119 - 0x77
      12'h67: dout <= 8'b01110111; //  103 : 119 - 0x77
      12'h68: dout <= 8'b01110111; //  104 : 119 - 0x77 -- Sprite 0xd
      12'h69: dout <= 8'b01110111; //  105 : 119 - 0x77
      12'h6A: dout <= 8'b01110111; //  106 : 119 - 0x77
      12'h6B: dout <= 8'b01110000; //  107 : 112 - 0x70
      12'h6C: dout <= 8'b01101111; //  108 : 111 - 0x6f
      12'h6D: dout <= 8'b01011111; //  109 :  95 - 0x5f
      12'h6E: dout <= 8'b00010101; //  110 :  21 - 0x15
      12'h6F: dout <= 8'b00000000; //  111 :   0 - 0x0
      12'h70: dout <= 8'b00000000; //  112 :   0 - 0x0 -- Sprite 0xe
      12'h71: dout <= 8'b11111100; //  113 : 252 - 0xfc
      12'h72: dout <= 8'b11111000; //  114 : 248 - 0xf8
      12'h73: dout <= 8'b11110110; //  115 : 246 - 0xf6
      12'h74: dout <= 8'b00001100; //  116 :  12 - 0xc
      12'h75: dout <= 8'b11101110; //  117 : 238 - 0xee
      12'h76: dout <= 8'b11101100; //  118 : 236 - 0xec
      12'h77: dout <= 8'b11101110; //  119 : 238 - 0xee
      12'h78: dout <= 8'b11101100; //  120 : 236 - 0xec -- Sprite 0xf
      12'h79: dout <= 8'b11101110; //  121 : 238 - 0xee
      12'h7A: dout <= 8'b11101100; //  122 : 236 - 0xec
      12'h7B: dout <= 8'b00001110; //  123 :  14 - 0xe
      12'h7C: dout <= 8'b11110100; //  124 : 244 - 0xf4
      12'h7D: dout <= 8'b11111010; //  125 : 250 - 0xfa
      12'h7E: dout <= 8'b01010100; //  126 :  84 - 0x54
      12'h7F: dout <= 8'b00000000; //  127 :   0 - 0x0
      12'h80: dout <= 8'b01100000; //  128 :  96 - 0x60 -- Sprite 0x10
      12'h81: dout <= 8'b01100000; //  129 :  96 - 0x60
      12'h82: dout <= 8'b01100000; //  130 :  96 - 0x60
      12'h83: dout <= 8'b01101111; //  131 : 111 - 0x6f
      12'h84: dout <= 8'b01101010; //  132 : 106 - 0x6a
      12'h85: dout <= 8'b01100000; //  133 :  96 - 0x60
      12'h86: dout <= 8'b01100000; //  134 :  96 - 0x60
      12'h87: dout <= 8'b01100000; //  135 :  96 - 0x60
      12'h88: dout <= 8'b00000110; //  136 :   6 - 0x6 -- Sprite 0x11
      12'h89: dout <= 8'b00000100; //  137 :   4 - 0x4
      12'h8A: dout <= 8'b00000110; //  138 :   6 - 0x6
      12'h8B: dout <= 8'b11110100; //  139 : 244 - 0xf4
      12'h8C: dout <= 8'b10100110; //  140 : 166 - 0xa6
      12'h8D: dout <= 8'b00000100; //  141 :   4 - 0x4
      12'h8E: dout <= 8'b00000110; //  142 :   6 - 0x6
      12'h8F: dout <= 8'b00000100; //  143 :   4 - 0x4
      12'h90: dout <= 8'b00000000; //  144 :   0 - 0x0 -- Sprite 0x12
      12'h91: dout <= 8'b00001000; //  145 :   8 - 0x8
      12'h92: dout <= 8'b00001000; //  146 :   8 - 0x8
      12'h93: dout <= 8'b00011100; //  147 :  28 - 0x1c
      12'h94: dout <= 8'b00011100; //  148 :  28 - 0x1c
      12'h95: dout <= 8'b00111100; //  149 :  60 - 0x3c
      12'h96: dout <= 8'b00111100; //  150 :  60 - 0x3c
      12'h97: dout <= 8'b00111100; //  151 :  60 - 0x3c
      12'h98: dout <= 8'b00111100; //  152 :  60 - 0x3c -- Sprite 0x13
      12'h99: dout <= 8'b01111110; //  153 : 126 - 0x7e
      12'h9A: dout <= 8'b01111110; //  154 : 126 - 0x7e
      12'h9B: dout <= 8'b01111110; //  155 : 126 - 0x7e
      12'h9C: dout <= 8'b01111110; //  156 : 126 - 0x7e
      12'h9D: dout <= 8'b01111110; //  157 : 126 - 0x7e
      12'h9E: dout <= 8'b01111110; //  158 : 126 - 0x7e
      12'h9F: dout <= 8'b00000000; //  159 :   0 - 0x0
      12'hA0: dout <= 8'b00000000; //  160 :   0 - 0x0 -- Sprite 0x14
      12'hA1: dout <= 8'b00000000; //  161 :   0 - 0x0
      12'hA2: dout <= 8'b00000101; //  162 :   5 - 0x5
      12'hA3: dout <= 8'b00000011; //  163 :   3 - 0x3
      12'hA4: dout <= 8'b00000000; //  164 :   0 - 0x0
      12'hA5: dout <= 8'b00000000; //  165 :   0 - 0x0
      12'hA6: dout <= 8'b00000010; //  166 :   2 - 0x2
      12'hA7: dout <= 8'b00001111; //  167 :  15 - 0xf
      12'hA8: dout <= 8'b00011100; //  168 :  28 - 0x1c -- Sprite 0x15
      12'hA9: dout <= 8'b00111010; //  169 :  58 - 0x3a
      12'hAA: dout <= 8'b00111100; //  170 :  60 - 0x3c
      12'hAB: dout <= 8'b00111111; //  171 :  63 - 0x3f
      12'hAC: dout <= 8'b00111000; //  172 :  56 - 0x38
      12'hAD: dout <= 8'b00011110; //  173 :  30 - 0x1e
      12'hAE: dout <= 8'b00001111; //  174 :  15 - 0xf
      12'hAF: dout <= 8'b00000000; //  175 :   0 - 0x0
      12'hB0: dout <= 8'b00000000; //  176 :   0 - 0x0 -- Sprite 0x16
      12'hB1: dout <= 8'b00000000; //  177 :   0 - 0x0
      12'hB2: dout <= 8'b01000000; //  178 :  64 - 0x40
      12'hB3: dout <= 8'b11000000; //  179 : 192 - 0xc0
      12'hB4: dout <= 8'b00000000; //  180 :   0 - 0x0
      12'hB5: dout <= 8'b10000000; //  181 : 128 - 0x80
      12'hB6: dout <= 8'b11000000; //  182 : 192 - 0xc0
      12'hB7: dout <= 8'b01110000; //  183 : 112 - 0x70
      12'hB8: dout <= 8'b00011000; //  184 :  24 - 0x18 -- Sprite 0x17
      12'hB9: dout <= 8'b11111100; //  185 : 252 - 0xfc
      12'hBA: dout <= 8'b00111100; //  186 :  60 - 0x3c
      12'hBB: dout <= 8'b01011100; //  187 :  92 - 0x5c
      12'hBC: dout <= 8'b00111100; //  188 :  60 - 0x3c
      12'hBD: dout <= 8'b11111000; //  189 : 248 - 0xf8
      12'hBE: dout <= 8'b11110000; //  190 : 240 - 0xf0
      12'hBF: dout <= 8'b00000000; //  191 :   0 - 0x0
      12'hC0: dout <= 8'b00000000; //  192 :   0 - 0x0 -- Sprite 0x18
      12'hC1: dout <= 8'b00111111; //  193 :  63 - 0x3f
      12'hC2: dout <= 8'b00111111; //  194 :  63 - 0x3f
      12'hC3: dout <= 8'b01111111; //  195 : 127 - 0x7f
      12'hC4: dout <= 8'b01111111; //  196 : 127 - 0x7f
      12'hC5: dout <= 8'b00000000; //  197 :   0 - 0x0
      12'hC6: dout <= 8'b00000000; //  198 :   0 - 0x0
      12'hC7: dout <= 8'b00000000; //  199 :   0 - 0x0
      12'hC8: dout <= 8'b00000000; //  200 :   0 - 0x0 -- Sprite 0x19
      12'hC9: dout <= 8'b11111100; //  201 : 252 - 0xfc
      12'hCA: dout <= 8'b11111100; //  202 : 252 - 0xfc
      12'hCB: dout <= 8'b11111110; //  203 : 254 - 0xfe
      12'hCC: dout <= 8'b11111110; //  204 : 254 - 0xfe
      12'hCD: dout <= 8'b00000000; //  205 :   0 - 0x0
      12'hCE: dout <= 8'b00000000; //  206 :   0 - 0x0
      12'hCF: dout <= 8'b00000000; //  207 :   0 - 0x0
      12'hD0: dout <= 8'b00000000; //  208 :   0 - 0x0 -- Sprite 0x1a
      12'hD1: dout <= 8'b00000000; //  209 :   0 - 0x0
      12'hD2: dout <= 8'b00000000; //  210 :   0 - 0x0
      12'hD3: dout <= 8'b00111111; //  211 :  63 - 0x3f
      12'hD4: dout <= 8'b00111111; //  212 :  63 - 0x3f
      12'hD5: dout <= 8'b01111111; //  213 : 127 - 0x7f
      12'hD6: dout <= 8'b01111111; //  214 : 127 - 0x7f
      12'hD7: dout <= 8'b00000000; //  215 :   0 - 0x0
      12'hD8: dout <= 8'b00000000; //  216 :   0 - 0x0 -- Sprite 0x1b
      12'hD9: dout <= 8'b00000000; //  217 :   0 - 0x0
      12'hDA: dout <= 8'b00000000; //  218 :   0 - 0x0
      12'hDB: dout <= 8'b11111100; //  219 : 252 - 0xfc
      12'hDC: dout <= 8'b11111100; //  220 : 252 - 0xfc
      12'hDD: dout <= 8'b11111110; //  221 : 254 - 0xfe
      12'hDE: dout <= 8'b11111110; //  222 : 254 - 0xfe
      12'hDF: dout <= 8'b00000000; //  223 :   0 - 0x0
      12'hE0: dout <= 8'b00000000; //  224 :   0 - 0x0 -- Sprite 0x1c
      12'hE1: dout <= 8'b01111111; //  225 : 127 - 0x7f
      12'hE2: dout <= 8'b01111111; //  226 : 127 - 0x7f
      12'hE3: dout <= 8'b01111111; //  227 : 127 - 0x7f
      12'hE4: dout <= 8'b01100100; //  228 : 100 - 0x64
      12'hE5: dout <= 8'b01011011; //  229 :  91 - 0x5b
      12'hE6: dout <= 8'b01011001; //  230 :  89 - 0x59
      12'hE7: dout <= 8'b01111111; //  231 : 127 - 0x7f
      12'hE8: dout <= 8'b01111111; //  232 : 127 - 0x7f -- Sprite 0x1d
      12'hE9: dout <= 8'b00000000; //  233 :   0 - 0x0
      12'hEA: dout <= 8'b00000001; //  234 :   1 - 0x1
      12'hEB: dout <= 8'b00000001; //  235 :   1 - 0x1
      12'hEC: dout <= 8'b00000001; //  236 :   1 - 0x1
      12'hED: dout <= 8'b00000001; //  237 :   1 - 0x1
      12'hEE: dout <= 8'b00000001; //  238 :   1 - 0x1
      12'hEF: dout <= 8'b00000000; //  239 :   0 - 0x0
      12'hF0: dout <= 8'b00000000; //  240 :   0 - 0x0 -- Sprite 0x1e
      12'hF1: dout <= 8'b11111110; //  241 : 254 - 0xfe
      12'hF2: dout <= 8'b11111110; //  242 : 254 - 0xfe
      12'hF3: dout <= 8'b11111110; //  243 : 254 - 0xfe
      12'hF4: dout <= 8'b10111110; //  244 : 190 - 0xbe
      12'hF5: dout <= 8'b00001010; //  245 :  10 - 0xa
      12'hF6: dout <= 8'b11100010; //  246 : 226 - 0xe2
      12'hF7: dout <= 8'b11111110; //  247 : 254 - 0xfe
      12'hF8: dout <= 8'b11111110; //  248 : 254 - 0xfe -- Sprite 0x1f
      12'hF9: dout <= 8'b00000000; //  249 :   0 - 0x0
      12'hFA: dout <= 8'b10000000; //  250 : 128 - 0x80
      12'hFB: dout <= 8'b10000000; //  251 : 128 - 0x80
      12'hFC: dout <= 8'b10000000; //  252 : 128 - 0x80
      12'hFD: dout <= 8'b10000000; //  253 : 128 - 0x80
      12'hFE: dout <= 8'b10000000; //  254 : 128 - 0x80
      12'hFF: dout <= 8'b00000000; //  255 :   0 - 0x0
      12'h100: dout <= 8'b00000000; //  256 :   0 - 0x0 -- Sprite 0x20
      12'h101: dout <= 8'b00000000; //  257 :   0 - 0x0
      12'h102: dout <= 8'b00000000; //  258 :   0 - 0x0
      12'h103: dout <= 8'b00000000; //  259 :   0 - 0x0
      12'h104: dout <= 8'b00000000; //  260 :   0 - 0x0
      12'h105: dout <= 8'b00000000; //  261 :   0 - 0x0
      12'h106: dout <= 8'b00000000; //  262 :   0 - 0x0
      12'h107: dout <= 8'b00000000; //  263 :   0 - 0x0
      12'h108: dout <= 8'b00000000; //  264 :   0 - 0x0 -- Sprite 0x21
      12'h109: dout <= 8'b00000000; //  265 :   0 - 0x0
      12'h10A: dout <= 8'b00000000; //  266 :   0 - 0x0
      12'h10B: dout <= 8'b00000000; //  267 :   0 - 0x0
      12'h10C: dout <= 8'b00000000; //  268 :   0 - 0x0
      12'h10D: dout <= 8'b00000000; //  269 :   0 - 0x0
      12'h10E: dout <= 8'b00000000; //  270 :   0 - 0x0
      12'h10F: dout <= 8'b00000000; //  271 :   0 - 0x0
      12'h110: dout <= 8'b00000000; //  272 :   0 - 0x0 -- Sprite 0x22
      12'h111: dout <= 8'b00000000; //  273 :   0 - 0x0
      12'h112: dout <= 8'b00011000; //  274 :  24 - 0x18
      12'h113: dout <= 8'b00010000; //  275 :  16 - 0x10
      12'h114: dout <= 8'b00011010; //  276 :  26 - 0x1a
      12'h115: dout <= 8'b00010001; //  277 :  17 - 0x11
      12'h116: dout <= 8'b00011010; //  278 :  26 - 0x1a
      12'h117: dout <= 8'b00000000; //  279 :   0 - 0x0
      12'h118: dout <= 8'b00000000; //  280 :   0 - 0x0 -- Sprite 0x23
      12'h119: dout <= 8'b00000000; //  281 :   0 - 0x0
      12'h11A: dout <= 8'b00000000; //  282 :   0 - 0x0
      12'h11B: dout <= 8'b00101000; //  283 :  40 - 0x28
      12'h11C: dout <= 8'b10001100; //  284 : 140 - 0x8c
      12'h11D: dout <= 8'b00101000; //  285 :  40 - 0x28
      12'h11E: dout <= 8'b10101100; //  286 : 172 - 0xac
      12'h11F: dout <= 8'b00000000; //  287 :   0 - 0x0
      12'h120: dout <= 8'b00000000; //  288 :   0 - 0x0 -- Sprite 0x24
      12'h121: dout <= 8'b00000000; //  289 :   0 - 0x0
      12'h122: dout <= 8'b00000000; //  290 :   0 - 0x0
      12'h123: dout <= 8'b00000000; //  291 :   0 - 0x0
      12'h124: dout <= 8'b00000000; //  292 :   0 - 0x0
      12'h125: dout <= 8'b00000000; //  293 :   0 - 0x0
      12'h126: dout <= 8'b00000000; //  294 :   0 - 0x0
      12'h127: dout <= 8'b00000000; //  295 :   0 - 0x0
      12'h128: dout <= 8'b00011100; //  296 :  28 - 0x1c -- Sprite 0x25
      12'h129: dout <= 8'b00111001; //  297 :  57 - 0x39
      12'h12A: dout <= 8'b00111111; //  298 :  63 - 0x3f
      12'h12B: dout <= 8'b00111110; //  299 :  62 - 0x3e
      12'h12C: dout <= 8'b00111111; //  300 :  63 - 0x3f
      12'h12D: dout <= 8'b00011110; //  301 :  30 - 0x1e
      12'h12E: dout <= 8'b00001111; //  302 :  15 - 0xf
      12'h12F: dout <= 8'b00000000; //  303 :   0 - 0x0
      12'h130: dout <= 8'b00000000; //  304 :   0 - 0x0 -- Sprite 0x26
      12'h131: dout <= 8'b00000000; //  305 :   0 - 0x0
      12'h132: dout <= 8'b01000000; //  306 :  64 - 0x40
      12'h133: dout <= 8'b11000000; //  307 : 192 - 0xc0
      12'h134: dout <= 8'b00000000; //  308 :   0 - 0x0
      12'h135: dout <= 8'b10000000; //  309 : 128 - 0x80
      12'h136: dout <= 8'b11000000; //  310 : 192 - 0xc0
      12'h137: dout <= 8'b11110000; //  311 : 240 - 0xf0
      12'h138: dout <= 8'b00111000; //  312 :  56 - 0x38 -- Sprite 0x27
      12'h139: dout <= 8'b10011100; //  313 : 156 - 0x9c
      12'h13A: dout <= 8'b10011100; //  314 : 156 - 0x9c
      12'h13B: dout <= 8'b00111100; //  315 :  60 - 0x3c
      12'h13C: dout <= 8'b11111100; //  316 : 252 - 0xfc
      12'h13D: dout <= 8'b01111000; //  317 : 120 - 0x78
      12'h13E: dout <= 8'b11110000; //  318 : 240 - 0xf0
      12'h13F: dout <= 8'b00000000; //  319 :   0 - 0x0
      12'h140: dout <= 8'b00000000; //  320 :   0 - 0x0 -- Sprite 0x28
      12'h141: dout <= 8'b00111110; //  321 :  62 - 0x3e
      12'h142: dout <= 8'b01011101; //  322 :  93 - 0x5d
      12'h143: dout <= 8'b01101011; //  323 : 107 - 0x6b
      12'h144: dout <= 8'b01110101; //  324 : 117 - 0x75
      12'h145: dout <= 8'b01110001; //  325 : 113 - 0x71
      12'h146: dout <= 8'b01110101; //  326 : 117 - 0x75
      12'h147: dout <= 8'b01110100; //  327 : 116 - 0x74
      12'h148: dout <= 8'b01110000; //  328 : 112 - 0x70 -- Sprite 0x29
      12'h149: dout <= 8'b01110111; //  329 : 119 - 0x77
      12'h14A: dout <= 8'b01110111; //  330 : 119 - 0x77
      12'h14B: dout <= 8'b01110000; //  331 : 112 - 0x70
      12'h14C: dout <= 8'b01101111; //  332 : 111 - 0x6f
      12'h14D: dout <= 8'b01011111; //  333 :  95 - 0x5f
      12'h14E: dout <= 8'b00010101; //  334 :  21 - 0x15
      12'h14F: dout <= 8'b00000000; //  335 :   0 - 0x0
      12'h150: dout <= 8'b00000000; //  336 :   0 - 0x0 -- Sprite 0x2a
      12'h151: dout <= 8'b01111100; //  337 : 124 - 0x7c
      12'h152: dout <= 8'b10111000; //  338 : 184 - 0xb8
      12'h153: dout <= 8'b11010110; //  339 : 214 - 0xd6
      12'h154: dout <= 8'b10101100; //  340 : 172 - 0xac
      12'h155: dout <= 8'b10001110; //  341 : 142 - 0x8e
      12'h156: dout <= 8'b10101100; //  342 : 172 - 0xac
      12'h157: dout <= 8'b00101110; //  343 :  46 - 0x2e
      12'h158: dout <= 8'b00001100; //  344 :  12 - 0xc -- Sprite 0x2b
      12'h159: dout <= 8'b11101110; //  345 : 238 - 0xee
      12'h15A: dout <= 8'b11101100; //  346 : 236 - 0xec
      12'h15B: dout <= 8'b00001110; //  347 :  14 - 0xe
      12'h15C: dout <= 8'b11110100; //  348 : 244 - 0xf4
      12'h15D: dout <= 8'b11111010; //  349 : 250 - 0xfa
      12'h15E: dout <= 8'b01010100; //  350 :  84 - 0x54
      12'h15F: dout <= 8'b00000000; //  351 :   0 - 0x0
      12'h160: dout <= 8'b00000000; //  352 :   0 - 0x0 -- Sprite 0x2c
      12'h161: dout <= 8'b00000000; //  353 :   0 - 0x0
      12'h162: dout <= 8'b00000000; //  354 :   0 - 0x0
      12'h163: dout <= 8'b00000000; //  355 :   0 - 0x0
      12'h164: dout <= 8'b00000000; //  356 :   0 - 0x0
      12'h165: dout <= 8'b00000000; //  357 :   0 - 0x0
      12'h166: dout <= 8'b00000000; //  358 :   0 - 0x0
      12'h167: dout <= 8'b00000000; //  359 :   0 - 0x0
      12'h168: dout <= 8'b00011110; //  360 :  30 - 0x1e -- Sprite 0x2d
      12'h169: dout <= 8'b00111110; //  361 :  62 - 0x3e
      12'h16A: dout <= 8'b00111110; //  362 :  62 - 0x3e
      12'h16B: dout <= 8'b00111110; //  363 :  62 - 0x3e
      12'h16C: dout <= 8'b00111111; //  364 :  63 - 0x3f
      12'h16D: dout <= 8'b00011110; //  365 :  30 - 0x1e
      12'h16E: dout <= 8'b00001111; //  366 :  15 - 0xf
      12'h16F: dout <= 8'b00000000; //  367 :   0 - 0x0
      12'h170: dout <= 8'b00000000; //  368 :   0 - 0x0 -- Sprite 0x2e
      12'h171: dout <= 8'b00000000; //  369 :   0 - 0x0
      12'h172: dout <= 8'b00000000; //  370 :   0 - 0x0
      12'h173: dout <= 8'b00000000; //  371 :   0 - 0x0
      12'h174: dout <= 8'b00000000; //  372 :   0 - 0x0
      12'h175: dout <= 8'b00000000; //  373 :   0 - 0x0
      12'h176: dout <= 8'b00000000; //  374 :   0 - 0x0
      12'h177: dout <= 8'b00000000; //  375 :   0 - 0x0
      12'h178: dout <= 8'b01111000; //  376 : 120 - 0x78 -- Sprite 0x2f
      12'h179: dout <= 8'b01111100; //  377 : 124 - 0x7c
      12'h17A: dout <= 8'b01111100; //  378 : 124 - 0x7c
      12'h17B: dout <= 8'b01111100; //  379 : 124 - 0x7c
      12'h17C: dout <= 8'b11111100; //  380 : 252 - 0xfc
      12'h17D: dout <= 8'b01111000; //  381 : 120 - 0x78
      12'h17E: dout <= 8'b11110000; //  382 : 240 - 0xf0
      12'h17F: dout <= 8'b00000000; //  383 :   0 - 0x0
      12'h180: dout <= 8'b00000000; //  384 :   0 - 0x0 -- Sprite 0x30
      12'h181: dout <= 8'b00011000; //  385 :  24 - 0x18
      12'h182: dout <= 8'b00111100; //  386 :  60 - 0x3c
      12'h183: dout <= 8'b01011010; //  387 :  90 - 0x5a
      12'h184: dout <= 8'b00011000; //  388 :  24 - 0x18
      12'h185: dout <= 8'b00011000; //  389 :  24 - 0x18
      12'h186: dout <= 8'b00011000; //  390 :  24 - 0x18
      12'h187: dout <= 8'b00000000; //  391 :   0 - 0x0
      12'h188: dout <= 8'b00000000; //  392 :   0 - 0x0 -- Sprite 0x31
      12'h189: dout <= 8'b00011000; //  393 :  24 - 0x18
      12'h18A: dout <= 8'b00011000; //  394 :  24 - 0x18
      12'h18B: dout <= 8'b00011000; //  395 :  24 - 0x18
      12'h18C: dout <= 8'b01011010; //  396 :  90 - 0x5a
      12'h18D: dout <= 8'b00111100; //  397 :  60 - 0x3c
      12'h18E: dout <= 8'b00011000; //  398 :  24 - 0x18
      12'h18F: dout <= 8'b00000000; //  399 :   0 - 0x0
      12'h190: dout <= 8'b00000001; //  400 :   1 - 0x1 -- Sprite 0x32
      12'h191: dout <= 8'b00000001; //  401 :   1 - 0x1
      12'h192: dout <= 8'b00000000; //  402 :   0 - 0x0
      12'h193: dout <= 8'b00000001; //  403 :   1 - 0x1
      12'h194: dout <= 8'b00000001; //  404 :   1 - 0x1
      12'h195: dout <= 8'b00000001; //  405 :   1 - 0x1
      12'h196: dout <= 8'b00000000; //  406 :   0 - 0x0
      12'h197: dout <= 8'b00000001; //  407 :   1 - 0x1
      12'h198: dout <= 8'b10000000; //  408 : 128 - 0x80 -- Sprite 0x33
      12'h199: dout <= 8'b00000000; //  409 :   0 - 0x0
      12'h19A: dout <= 8'b10000000; //  410 : 128 - 0x80
      12'h19B: dout <= 8'b10000000; //  411 : 128 - 0x80
      12'h19C: dout <= 8'b10000000; //  412 : 128 - 0x80
      12'h19D: dout <= 8'b00000000; //  413 :   0 - 0x0
      12'h19E: dout <= 8'b10000000; //  414 : 128 - 0x80
      12'h19F: dout <= 8'b10000000; //  415 : 128 - 0x80
      12'h1A0: dout <= 8'b00000000; //  416 :   0 - 0x0 -- Sprite 0x34
      12'h1A1: dout <= 8'b00000000; //  417 :   0 - 0x0
      12'h1A2: dout <= 8'b00011000; //  418 :  24 - 0x18
      12'h1A3: dout <= 8'b00111100; //  419 :  60 - 0x3c
      12'h1A4: dout <= 8'b00111110; //  420 :  62 - 0x3e
      12'h1A5: dout <= 8'b01111111; //  421 : 127 - 0x7f
      12'h1A6: dout <= 8'b01111111; //  422 : 127 - 0x7f
      12'h1A7: dout <= 8'b01111111; //  423 : 127 - 0x7f
      12'h1A8: dout <= 8'b00111111; //  424 :  63 - 0x3f -- Sprite 0x35
      12'h1A9: dout <= 8'b00111111; //  425 :  63 - 0x3f
      12'h1AA: dout <= 8'b00011111; //  426 :  31 - 0x1f
      12'h1AB: dout <= 8'b00001111; //  427 :  15 - 0xf
      12'h1AC: dout <= 8'b00000111; //  428 :   7 - 0x7
      12'h1AD: dout <= 8'b00000011; //  429 :   3 - 0x3
      12'h1AE: dout <= 8'b00000001; //  430 :   1 - 0x1
      12'h1AF: dout <= 8'b00000000; //  431 :   0 - 0x0
      12'h1B0: dout <= 8'b00000000; //  432 :   0 - 0x0 -- Sprite 0x36
      12'h1B1: dout <= 8'b00000000; //  433 :   0 - 0x0
      12'h1B2: dout <= 8'b00011000; //  434 :  24 - 0x18
      12'h1B3: dout <= 8'b00111100; //  435 :  60 - 0x3c
      12'h1B4: dout <= 8'b01111100; //  436 : 124 - 0x7c
      12'h1B5: dout <= 8'b11111110; //  437 : 254 - 0xfe
      12'h1B6: dout <= 8'b11111110; //  438 : 254 - 0xfe
      12'h1B7: dout <= 8'b11111110; //  439 : 254 - 0xfe
      12'h1B8: dout <= 8'b11111100; //  440 : 252 - 0xfc -- Sprite 0x37
      12'h1B9: dout <= 8'b11111100; //  441 : 252 - 0xfc
      12'h1BA: dout <= 8'b11111000; //  442 : 248 - 0xf8
      12'h1BB: dout <= 8'b11110000; //  443 : 240 - 0xf0
      12'h1BC: dout <= 8'b11100000; //  444 : 224 - 0xe0
      12'h1BD: dout <= 8'b11000000; //  445 : 192 - 0xc0
      12'h1BE: dout <= 8'b10000000; //  446 : 128 - 0x80
      12'h1BF: dout <= 8'b00000000; //  447 :   0 - 0x0
      12'h1C0: dout <= 8'b00000000; //  448 :   0 - 0x0 -- Sprite 0x38
      12'h1C1: dout <= 8'b00000000; //  449 :   0 - 0x0
      12'h1C2: dout <= 8'b00000110; //  450 :   6 - 0x6
      12'h1C3: dout <= 8'b00000111; //  451 :   7 - 0x7
      12'h1C4: dout <= 8'b00000111; //  452 :   7 - 0x7
      12'h1C5: dout <= 8'b00000011; //  453 :   3 - 0x3
      12'h1C6: dout <= 8'b00000001; //  454 :   1 - 0x1
      12'h1C7: dout <= 8'b00000000; //  455 :   0 - 0x0
      12'h1C8: dout <= 8'b00000000; //  456 :   0 - 0x0 -- Sprite 0x39
      12'h1C9: dout <= 8'b00000000; //  457 :   0 - 0x0
      12'h1CA: dout <= 8'b00000000; //  458 :   0 - 0x0
      12'h1CB: dout <= 8'b00000000; //  459 :   0 - 0x0
      12'h1CC: dout <= 8'b00000000; //  460 :   0 - 0x0
      12'h1CD: dout <= 8'b00000000; //  461 :   0 - 0x0
      12'h1CE: dout <= 8'b00000000; //  462 :   0 - 0x0
      12'h1CF: dout <= 8'b00000000; //  463 :   0 - 0x0
      12'h1D0: dout <= 8'b00000000; //  464 :   0 - 0x0 -- Sprite 0x3a
      12'h1D1: dout <= 8'b00000000; //  465 :   0 - 0x0
      12'h1D2: dout <= 8'b01100000; //  466 :  96 - 0x60
      12'h1D3: dout <= 8'b11100000; //  467 : 224 - 0xe0
      12'h1D4: dout <= 8'b11100000; //  468 : 224 - 0xe0
      12'h1D5: dout <= 8'b11000000; //  469 : 192 - 0xc0
      12'h1D6: dout <= 8'b10000000; //  470 : 128 - 0x80
      12'h1D7: dout <= 8'b00000000; //  471 :   0 - 0x0
      12'h1D8: dout <= 8'b00000000; //  472 :   0 - 0x0 -- Sprite 0x3b
      12'h1D9: dout <= 8'b00101010; //  473 :  42 - 0x2a
      12'h1DA: dout <= 8'b01000000; //  474 :  64 - 0x40
      12'h1DB: dout <= 8'b00000010; //  475 :   2 - 0x2
      12'h1DC: dout <= 8'b01000000; //  476 :  64 - 0x40
      12'h1DD: dout <= 8'b00000010; //  477 :   2 - 0x2
      12'h1DE: dout <= 8'b01010100; //  478 :  84 - 0x54
      12'h1DF: dout <= 8'b00000000; //  479 :   0 - 0x0
      12'h1E0: dout <= 8'b00000000; //  480 :   0 - 0x0 -- Sprite 0x3c
      12'h1E1: dout <= 8'b00000000; //  481 :   0 - 0x0
      12'h1E2: dout <= 8'b00000000; //  482 :   0 - 0x0
      12'h1E3: dout <= 8'b00000000; //  483 :   0 - 0x0
      12'h1E4: dout <= 8'b00000000; //  484 :   0 - 0x0
      12'h1E5: dout <= 8'b00000000; //  485 :   0 - 0x0
      12'h1E6: dout <= 8'b00000000; //  486 :   0 - 0x0
      12'h1E7: dout <= 8'b00000000; //  487 :   0 - 0x0
      12'h1E8: dout <= 8'b11111111; //  488 : 255 - 0xff -- Sprite 0x3d
      12'h1E9: dout <= 8'b11111111; //  489 : 255 - 0xff
      12'h1EA: dout <= 8'b11111111; //  490 : 255 - 0xff
      12'h1EB: dout <= 8'b11111111; //  491 : 255 - 0xff
      12'h1EC: dout <= 8'b11111111; //  492 : 255 - 0xff
      12'h1ED: dout <= 8'b11111111; //  493 : 255 - 0xff
      12'h1EE: dout <= 8'b11111111; //  494 : 255 - 0xff
      12'h1EF: dout <= 8'b11111111; //  495 : 255 - 0xff
      12'h1F0: dout <= 8'b11111111; //  496 : 255 - 0xff -- Sprite 0x3e
      12'h1F1: dout <= 8'b11111111; //  497 : 255 - 0xff
      12'h1F2: dout <= 8'b11111111; //  498 : 255 - 0xff
      12'h1F3: dout <= 8'b11111111; //  499 : 255 - 0xff
      12'h1F4: dout <= 8'b11111111; //  500 : 255 - 0xff
      12'h1F5: dout <= 8'b11111111; //  501 : 255 - 0xff
      12'h1F6: dout <= 8'b11111111; //  502 : 255 - 0xff
      12'h1F7: dout <= 8'b11111111; //  503 : 255 - 0xff
      12'h1F8: dout <= 8'b00000000; //  504 :   0 - 0x0 -- Sprite 0x3f
      12'h1F9: dout <= 8'b00000000; //  505 :   0 - 0x0
      12'h1FA: dout <= 8'b00000000; //  506 :   0 - 0x0
      12'h1FB: dout <= 8'b00000000; //  507 :   0 - 0x0
      12'h1FC: dout <= 8'b00000000; //  508 :   0 - 0x0
      12'h1FD: dout <= 8'b00000000; //  509 :   0 - 0x0
      12'h1FE: dout <= 8'b00000000; //  510 :   0 - 0x0
      12'h1FF: dout <= 8'b00000000; //  511 :   0 - 0x0
      12'h200: dout <= 8'b00000000; //  512 :   0 - 0x0 -- Sprite 0x40
      12'h201: dout <= 8'b00000000; //  513 :   0 - 0x0
      12'h202: dout <= 8'b00000000; //  514 :   0 - 0x0
      12'h203: dout <= 8'b00000000; //  515 :   0 - 0x0
      12'h204: dout <= 8'b00000000; //  516 :   0 - 0x0
      12'h205: dout <= 8'b00000000; //  517 :   0 - 0x0
      12'h206: dout <= 8'b00000000; //  518 :   0 - 0x0
      12'h207: dout <= 8'b00000000; //  519 :   0 - 0x0
      12'h208: dout <= 8'b00000000; //  520 :   0 - 0x0 -- Sprite 0x41
      12'h209: dout <= 8'b00000000; //  521 :   0 - 0x0
      12'h20A: dout <= 8'b00000000; //  522 :   0 - 0x0
      12'h20B: dout <= 8'b00000000; //  523 :   0 - 0x0
      12'h20C: dout <= 8'b00000000; //  524 :   0 - 0x0
      12'h20D: dout <= 8'b00000000; //  525 :   0 - 0x0
      12'h20E: dout <= 8'b00000000; //  526 :   0 - 0x0
      12'h20F: dout <= 8'b00000000; //  527 :   0 - 0x0
      12'h210: dout <= 8'b00000000; //  528 :   0 - 0x0 -- Sprite 0x42
      12'h211: dout <= 8'b00000000; //  529 :   0 - 0x0
      12'h212: dout <= 8'b00000000; //  530 :   0 - 0x0
      12'h213: dout <= 8'b00000000; //  531 :   0 - 0x0
      12'h214: dout <= 8'b00000000; //  532 :   0 - 0x0
      12'h215: dout <= 8'b00000000; //  533 :   0 - 0x0
      12'h216: dout <= 8'b00000000; //  534 :   0 - 0x0
      12'h217: dout <= 8'b00000000; //  535 :   0 - 0x0
      12'h218: dout <= 8'b00000000; //  536 :   0 - 0x0 -- Sprite 0x43
      12'h219: dout <= 8'b00000000; //  537 :   0 - 0x0
      12'h21A: dout <= 8'b00000000; //  538 :   0 - 0x0
      12'h21B: dout <= 8'b00000000; //  539 :   0 - 0x0
      12'h21C: dout <= 8'b00000000; //  540 :   0 - 0x0
      12'h21D: dout <= 8'b00000000; //  541 :   0 - 0x0
      12'h21E: dout <= 8'b00000000; //  542 :   0 - 0x0
      12'h21F: dout <= 8'b00000000; //  543 :   0 - 0x0
      12'h220: dout <= 8'b00000000; //  544 :   0 - 0x0 -- Sprite 0x44
      12'h221: dout <= 8'b00000000; //  545 :   0 - 0x0
      12'h222: dout <= 8'b00000000; //  546 :   0 - 0x0
      12'h223: dout <= 8'b00000000; //  547 :   0 - 0x0
      12'h224: dout <= 8'b00000000; //  548 :   0 - 0x0
      12'h225: dout <= 8'b00000000; //  549 :   0 - 0x0
      12'h226: dout <= 8'b00000000; //  550 :   0 - 0x0
      12'h227: dout <= 8'b00000000; //  551 :   0 - 0x0
      12'h228: dout <= 8'b00000000; //  552 :   0 - 0x0 -- Sprite 0x45
      12'h229: dout <= 8'b00000000; //  553 :   0 - 0x0
      12'h22A: dout <= 8'b00000000; //  554 :   0 - 0x0
      12'h22B: dout <= 8'b00000000; //  555 :   0 - 0x0
      12'h22C: dout <= 8'b00000000; //  556 :   0 - 0x0
      12'h22D: dout <= 8'b00000000; //  557 :   0 - 0x0
      12'h22E: dout <= 8'b00000000; //  558 :   0 - 0x0
      12'h22F: dout <= 8'b00000000; //  559 :   0 - 0x0
      12'h230: dout <= 8'b00000000; //  560 :   0 - 0x0 -- Sprite 0x46
      12'h231: dout <= 8'b00000000; //  561 :   0 - 0x0
      12'h232: dout <= 8'b00000000; //  562 :   0 - 0x0
      12'h233: dout <= 8'b00000000; //  563 :   0 - 0x0
      12'h234: dout <= 8'b00000000; //  564 :   0 - 0x0
      12'h235: dout <= 8'b00000000; //  565 :   0 - 0x0
      12'h236: dout <= 8'b00000000; //  566 :   0 - 0x0
      12'h237: dout <= 8'b00000000; //  567 :   0 - 0x0
      12'h238: dout <= 8'b00000000; //  568 :   0 - 0x0 -- Sprite 0x47
      12'h239: dout <= 8'b00000000; //  569 :   0 - 0x0
      12'h23A: dout <= 8'b00000000; //  570 :   0 - 0x0
      12'h23B: dout <= 8'b00000000; //  571 :   0 - 0x0
      12'h23C: dout <= 8'b00000000; //  572 :   0 - 0x0
      12'h23D: dout <= 8'b00000000; //  573 :   0 - 0x0
      12'h23E: dout <= 8'b00000000; //  574 :   0 - 0x0
      12'h23F: dout <= 8'b00000000; //  575 :   0 - 0x0
      12'h240: dout <= 8'b00000000; //  576 :   0 - 0x0 -- Sprite 0x48
      12'h241: dout <= 8'b00000000; //  577 :   0 - 0x0
      12'h242: dout <= 8'b00000000; //  578 :   0 - 0x0
      12'h243: dout <= 8'b00000000; //  579 :   0 - 0x0
      12'h244: dout <= 8'b00000000; //  580 :   0 - 0x0
      12'h245: dout <= 8'b00000000; //  581 :   0 - 0x0
      12'h246: dout <= 8'b00000000; //  582 :   0 - 0x0
      12'h247: dout <= 8'b00000000; //  583 :   0 - 0x0
      12'h248: dout <= 8'b00000000; //  584 :   0 - 0x0 -- Sprite 0x49
      12'h249: dout <= 8'b00000000; //  585 :   0 - 0x0
      12'h24A: dout <= 8'b00000000; //  586 :   0 - 0x0
      12'h24B: dout <= 8'b00000000; //  587 :   0 - 0x0
      12'h24C: dout <= 8'b00000000; //  588 :   0 - 0x0
      12'h24D: dout <= 8'b00000000; //  589 :   0 - 0x0
      12'h24E: dout <= 8'b00000000; //  590 :   0 - 0x0
      12'h24F: dout <= 8'b00000000; //  591 :   0 - 0x0
      12'h250: dout <= 8'b00000000; //  592 :   0 - 0x0 -- Sprite 0x4a
      12'h251: dout <= 8'b00000000; //  593 :   0 - 0x0
      12'h252: dout <= 8'b00000000; //  594 :   0 - 0x0
      12'h253: dout <= 8'b00000000; //  595 :   0 - 0x0
      12'h254: dout <= 8'b00000000; //  596 :   0 - 0x0
      12'h255: dout <= 8'b00000000; //  597 :   0 - 0x0
      12'h256: dout <= 8'b00000000; //  598 :   0 - 0x0
      12'h257: dout <= 8'b00000000; //  599 :   0 - 0x0
      12'h258: dout <= 8'b00000000; //  600 :   0 - 0x0 -- Sprite 0x4b
      12'h259: dout <= 8'b00000000; //  601 :   0 - 0x0
      12'h25A: dout <= 8'b00000000; //  602 :   0 - 0x0
      12'h25B: dout <= 8'b00000000; //  603 :   0 - 0x0
      12'h25C: dout <= 8'b00000000; //  604 :   0 - 0x0
      12'h25D: dout <= 8'b00000000; //  605 :   0 - 0x0
      12'h25E: dout <= 8'b00000000; //  606 :   0 - 0x0
      12'h25F: dout <= 8'b00000000; //  607 :   0 - 0x0
      12'h260: dout <= 8'b00000000; //  608 :   0 - 0x0 -- Sprite 0x4c
      12'h261: dout <= 8'b00000000; //  609 :   0 - 0x0
      12'h262: dout <= 8'b00000000; //  610 :   0 - 0x0
      12'h263: dout <= 8'b00000000; //  611 :   0 - 0x0
      12'h264: dout <= 8'b00000000; //  612 :   0 - 0x0
      12'h265: dout <= 8'b00000000; //  613 :   0 - 0x0
      12'h266: dout <= 8'b00000000; //  614 :   0 - 0x0
      12'h267: dout <= 8'b00000000; //  615 :   0 - 0x0
      12'h268: dout <= 8'b00000000; //  616 :   0 - 0x0 -- Sprite 0x4d
      12'h269: dout <= 8'b00000000; //  617 :   0 - 0x0
      12'h26A: dout <= 8'b00000000; //  618 :   0 - 0x0
      12'h26B: dout <= 8'b00000000; //  619 :   0 - 0x0
      12'h26C: dout <= 8'b00000000; //  620 :   0 - 0x0
      12'h26D: dout <= 8'b00000000; //  621 :   0 - 0x0
      12'h26E: dout <= 8'b00000000; //  622 :   0 - 0x0
      12'h26F: dout <= 8'b00000000; //  623 :   0 - 0x0
      12'h270: dout <= 8'b00000000; //  624 :   0 - 0x0 -- Sprite 0x4e
      12'h271: dout <= 8'b00000000; //  625 :   0 - 0x0
      12'h272: dout <= 8'b00000000; //  626 :   0 - 0x0
      12'h273: dout <= 8'b00000000; //  627 :   0 - 0x0
      12'h274: dout <= 8'b00000000; //  628 :   0 - 0x0
      12'h275: dout <= 8'b00000000; //  629 :   0 - 0x0
      12'h276: dout <= 8'b00000000; //  630 :   0 - 0x0
      12'h277: dout <= 8'b00000000; //  631 :   0 - 0x0
      12'h278: dout <= 8'b00000000; //  632 :   0 - 0x0 -- Sprite 0x4f
      12'h279: dout <= 8'b00000000; //  633 :   0 - 0x0
      12'h27A: dout <= 8'b00000000; //  634 :   0 - 0x0
      12'h27B: dout <= 8'b00000000; //  635 :   0 - 0x0
      12'h27C: dout <= 8'b00000000; //  636 :   0 - 0x0
      12'h27D: dout <= 8'b00000000; //  637 :   0 - 0x0
      12'h27E: dout <= 8'b00000000; //  638 :   0 - 0x0
      12'h27F: dout <= 8'b00000000; //  639 :   0 - 0x0
      12'h280: dout <= 8'b00000000; //  640 :   0 - 0x0 -- Sprite 0x50
      12'h281: dout <= 8'b00111111; //  641 :  63 - 0x3f
      12'h282: dout <= 8'b01111111; //  642 : 127 - 0x7f
      12'h283: dout <= 8'b01111111; //  643 : 127 - 0x7f
      12'h284: dout <= 8'b01111111; //  644 : 127 - 0x7f
      12'h285: dout <= 8'b00111100; //  645 :  60 - 0x3c
      12'h286: dout <= 8'b00000000; //  646 :   0 - 0x0
      12'h287: dout <= 8'b01000000; //  647 :  64 - 0x40
      12'h288: dout <= 8'b00000000; //  648 :   0 - 0x0 -- Sprite 0x51
      12'h289: dout <= 8'b11111100; //  649 : 252 - 0xfc
      12'h28A: dout <= 8'b11111110; //  650 : 254 - 0xfe
      12'h28B: dout <= 8'b11111110; //  651 : 254 - 0xfe
      12'h28C: dout <= 8'b11111110; //  652 : 254 - 0xfe
      12'h28D: dout <= 8'b00111100; //  653 :  60 - 0x3c
      12'h28E: dout <= 8'b00000000; //  654 :   0 - 0x0
      12'h28F: dout <= 8'b00000010; //  655 :   2 - 0x2
      12'h290: dout <= 8'b00000000; //  656 :   0 - 0x0 -- Sprite 0x52
      12'h291: dout <= 8'b00000000; //  657 :   0 - 0x0
      12'h292: dout <= 8'b00000011; //  658 :   3 - 0x3
      12'h293: dout <= 8'b00000111; //  659 :   7 - 0x7
      12'h294: dout <= 8'b00001111; //  660 :  15 - 0xf
      12'h295: dout <= 8'b00011111; //  661 :  31 - 0x1f
      12'h296: dout <= 8'b00111111; //  662 :  63 - 0x3f
      12'h297: dout <= 8'b00110000; //  663 :  48 - 0x30
      12'h298: dout <= 8'b00000000; //  664 :   0 - 0x0 -- Sprite 0x53
      12'h299: dout <= 8'b00000000; //  665 :   0 - 0x0
      12'h29A: dout <= 8'b10100000; //  666 : 160 - 0xa0
      12'h29B: dout <= 8'b10110000; //  667 : 176 - 0xb0
      12'h29C: dout <= 8'b10110000; //  668 : 176 - 0xb0
      12'h29D: dout <= 8'b10111000; //  669 : 184 - 0xb8
      12'h29E: dout <= 8'b01111100; //  670 : 124 - 0x7c
      12'h29F: dout <= 8'b01111100; //  671 : 124 - 0x7c
      12'h2A0: dout <= 8'b00000000; //  672 :   0 - 0x0 -- Sprite 0x54
      12'h2A1: dout <= 8'b00100001; //  673 :  33 - 0x21
      12'h2A2: dout <= 8'b01110001; //  674 : 113 - 0x71
      12'h2A3: dout <= 8'b00111010; //  675 :  58 - 0x3a
      12'h2A4: dout <= 8'b01101101; //  676 : 109 - 0x6d
      12'h2A5: dout <= 8'b00111000; //  677 :  56 - 0x38
      12'h2A6: dout <= 8'b00011101; //  678 :  29 - 0x1d
      12'h2A7: dout <= 8'b00101111; //  679 :  47 - 0x2f
      12'h2A8: dout <= 8'b00000000; //  680 :   0 - 0x0 -- Sprite 0x55
      12'h2A9: dout <= 8'b00100001; //  681 :  33 - 0x21
      12'h2AA: dout <= 8'b01110001; //  682 : 113 - 0x71
      12'h2AB: dout <= 8'b00111010; //  683 :  58 - 0x3a
      12'h2AC: dout <= 8'b01101101; //  684 : 109 - 0x6d
      12'h2AD: dout <= 8'b10111000; //  685 : 184 - 0xb8
      12'h2AE: dout <= 8'b00011101; //  686 :  29 - 0x1d
      12'h2AF: dout <= 8'b10101111; //  687 : 175 - 0xaf
      12'h2B0: dout <= 8'b00000000; //  688 :   0 - 0x0 -- Sprite 0x56
      12'h2B1: dout <= 8'b00100000; //  689 :  32 - 0x20
      12'h2B2: dout <= 8'b01110000; //  690 : 112 - 0x70
      12'h2B3: dout <= 8'b00111010; //  691 :  58 - 0x3a
      12'h2B4: dout <= 8'b01101100; //  692 : 108 - 0x6c
      12'h2B5: dout <= 8'b10111000; //  693 : 184 - 0xb8
      12'h2B6: dout <= 8'b00011100; //  694 :  28 - 0x1c
      12'h2B7: dout <= 8'b10101110; //  695 : 174 - 0xae
      12'h2B8: dout <= 8'b00000000; //  696 :   0 - 0x0 -- Sprite 0x57
      12'h2B9: dout <= 8'b01111111; //  697 : 127 - 0x7f
      12'h2BA: dout <= 8'b01001100; //  698 :  76 - 0x4c
      12'h2BB: dout <= 8'b00110011; //  699 :  51 - 0x33
      12'h2BC: dout <= 8'b00000000; //  700 :   0 - 0x0
      12'h2BD: dout <= 8'b00000000; //  701 :   0 - 0x0
      12'h2BE: dout <= 8'b00000000; //  702 :   0 - 0x0
      12'h2BF: dout <= 8'b00000000; //  703 :   0 - 0x0
      12'h2C0: dout <= 8'b00000000; //  704 :   0 - 0x0 -- Sprite 0x58
      12'h2C1: dout <= 8'b11111111; //  705 : 255 - 0xff
      12'h2C2: dout <= 8'b11001100; //  706 : 204 - 0xcc
      12'h2C3: dout <= 8'b00110011; //  707 :  51 - 0x33
      12'h2C4: dout <= 8'b11001100; //  708 : 204 - 0xcc
      12'h2C5: dout <= 8'b00000000; //  709 :   0 - 0x0
      12'h2C6: dout <= 8'b00000000; //  710 :   0 - 0x0
      12'h2C7: dout <= 8'b00000000; //  711 :   0 - 0x0
      12'h2C8: dout <= 8'b00000000; //  712 :   0 - 0x0 -- Sprite 0x59
      12'h2C9: dout <= 8'b11111110; //  713 : 254 - 0xfe
      12'h2CA: dout <= 8'b11001100; //  714 : 204 - 0xcc
      12'h2CB: dout <= 8'b00110000; //  715 :  48 - 0x30
      12'h2CC: dout <= 8'b11000000; //  716 : 192 - 0xc0
      12'h2CD: dout <= 8'b00000000; //  717 :   0 - 0x0
      12'h2CE: dout <= 8'b00000000; //  718 :   0 - 0x0
      12'h2CF: dout <= 8'b00000000; //  719 :   0 - 0x0
      12'h2D0: dout <= 8'b00000000; //  720 :   0 - 0x0 -- Sprite 0x5a
      12'h2D1: dout <= 8'b00000000; //  721 :   0 - 0x0
      12'h2D2: dout <= 8'b00000000; //  722 :   0 - 0x0
      12'h2D3: dout <= 8'b00000000; //  723 :   0 - 0x0
      12'h2D4: dout <= 8'b00000000; //  724 :   0 - 0x0
      12'h2D5: dout <= 8'b00000000; //  725 :   0 - 0x0
      12'h2D6: dout <= 8'b00000000; //  726 :   0 - 0x0
      12'h2D7: dout <= 8'b00000000; //  727 :   0 - 0x0
      12'h2D8: dout <= 8'b00000000; //  728 :   0 - 0x0 -- Sprite 0x5b
      12'h2D9: dout <= 8'b00000000; //  729 :   0 - 0x0
      12'h2DA: dout <= 8'b00000000; //  730 :   0 - 0x0
      12'h2DB: dout <= 8'b00000000; //  731 :   0 - 0x0
      12'h2DC: dout <= 8'b00000001; //  732 :   1 - 0x1
      12'h2DD: dout <= 8'b00000001; //  733 :   1 - 0x1
      12'h2DE: dout <= 8'b00000011; //  734 :   3 - 0x3
      12'h2DF: dout <= 8'b00000011; //  735 :   3 - 0x3
      12'h2E0: dout <= 8'b00000000; //  736 :   0 - 0x0 -- Sprite 0x5c
      12'h2E1: dout <= 8'b00000000; //  737 :   0 - 0x0
      12'h2E2: dout <= 8'b00000001; //  738 :   1 - 0x1
      12'h2E3: dout <= 8'b01111110; //  739 : 126 - 0x7e
      12'h2E4: dout <= 8'b11111111; //  740 : 255 - 0xff
      12'h2E5: dout <= 8'b11111111; //  741 : 255 - 0xff
      12'h2E6: dout <= 8'b11111111; //  742 : 255 - 0xff
      12'h2E7: dout <= 8'b11111111; //  743 : 255 - 0xff
      12'h2E8: dout <= 8'b00000000; //  744 :   0 - 0x0 -- Sprite 0x5d
      12'h2E9: dout <= 8'b11111111; //  745 : 255 - 0xff
      12'h2EA: dout <= 8'b11111111; //  746 : 255 - 0xff
      12'h2EB: dout <= 8'b11111111; //  747 : 255 - 0xff
      12'h2EC: dout <= 8'b01111111; //  748 : 127 - 0x7f
      12'h2ED: dout <= 8'b11111111; //  749 : 255 - 0xff
      12'h2EE: dout <= 8'b11111111; //  750 : 255 - 0xff
      12'h2EF: dout <= 8'b11111111; //  751 : 255 - 0xff
      12'h2F0: dout <= 8'b00000000; //  752 :   0 - 0x0 -- Sprite 0x5e
      12'h2F1: dout <= 8'b00000000; //  753 :   0 - 0x0
      12'h2F2: dout <= 8'b10000000; //  754 : 128 - 0x80
      12'h2F3: dout <= 8'b01111110; //  755 : 126 - 0x7e
      12'h2F4: dout <= 8'b10111111; //  756 : 191 - 0xbf
      12'h2F5: dout <= 8'b11111111; //  757 : 255 - 0xff
      12'h2F6: dout <= 8'b11111111; //  758 : 255 - 0xff
      12'h2F7: dout <= 8'b11111111; //  759 : 255 - 0xff
      12'h2F8: dout <= 8'b00000000; //  760 :   0 - 0x0 -- Sprite 0x5f
      12'h2F9: dout <= 8'b00000000; //  761 :   0 - 0x0
      12'h2FA: dout <= 8'b00000000; //  762 :   0 - 0x0
      12'h2FB: dout <= 8'b00000000; //  763 :   0 - 0x0
      12'h2FC: dout <= 8'b10000000; //  764 : 128 - 0x80
      12'h2FD: dout <= 8'b10000000; //  765 : 128 - 0x80
      12'h2FE: dout <= 8'b11000000; //  766 : 192 - 0xc0
      12'h2FF: dout <= 8'b11000000; //  767 : 192 - 0xc0
      12'h300: dout <= 8'b01111111; //  768 : 127 - 0x7f -- Sprite 0x60
      12'h301: dout <= 8'b01111111; //  769 : 127 - 0x7f
      12'h302: dout <= 8'b01111101; //  770 : 125 - 0x7d
      12'h303: dout <= 8'b01111111; //  771 : 127 - 0x7f
      12'h304: dout <= 8'b00111111; //  772 :  63 - 0x3f
      12'h305: dout <= 8'b01111111; //  773 : 127 - 0x7f
      12'h306: dout <= 8'b01111111; //  774 : 127 - 0x7f
      12'h307: dout <= 8'b01110111; //  775 : 119 - 0x77
      12'h308: dout <= 8'b11111110; //  776 : 254 - 0xfe -- Sprite 0x61
      12'h309: dout <= 8'b11111110; //  777 : 254 - 0xfe
      12'h30A: dout <= 8'b11111100; //  778 : 252 - 0xfc
      12'h30B: dout <= 8'b11111110; //  779 : 254 - 0xfe
      12'h30C: dout <= 8'b10111110; //  780 : 190 - 0xbe
      12'h30D: dout <= 8'b11111110; //  781 : 254 - 0xfe
      12'h30E: dout <= 8'b11111110; //  782 : 254 - 0xfe
      12'h30F: dout <= 8'b11110110; //  783 : 246 - 0xf6
      12'h310: dout <= 8'b00000111; //  784 :   7 - 0x7 -- Sprite 0x62
      12'h311: dout <= 8'b00011111; //  785 :  31 - 0x1f
      12'h312: dout <= 8'b00111111; //  786 :  63 - 0x3f
      12'h313: dout <= 8'b00111111; //  787 :  63 - 0x3f
      12'h314: dout <= 8'b00111111; //  788 :  63 - 0x3f
      12'h315: dout <= 8'b00011111; //  789 :  31 - 0x1f
      12'h316: dout <= 8'b00001111; //  790 :  15 - 0xf
      12'h317: dout <= 8'b00000000; //  791 :   0 - 0x0
      12'h318: dout <= 8'b01111110; //  792 : 126 - 0x7e -- Sprite 0x63
      12'h319: dout <= 8'b01111100; //  793 : 124 - 0x7c
      12'h31A: dout <= 8'b00111110; //  794 :  62 - 0x3e
      12'h31B: dout <= 8'b10111100; //  795 : 188 - 0xbc
      12'h31C: dout <= 8'b10111110; //  796 : 190 - 0xbe
      12'h31D: dout <= 8'b10011100; //  797 : 156 - 0x9c
      12'h31E: dout <= 8'b11011000; //  798 : 216 - 0xd8
      12'h31F: dout <= 8'b00000000; //  799 :   0 - 0x0
      12'h320: dout <= 8'b01000110; //  800 :  70 - 0x46 -- Sprite 0x64
      12'h321: dout <= 8'b01101011; //  801 : 107 - 0x6b
      12'h322: dout <= 8'b01110001; //  802 : 113 - 0x71
      12'h323: dout <= 8'b00111010; //  803 :  58 - 0x3a
      12'h324: dout <= 8'b01101101; //  804 : 109 - 0x6d
      12'h325: dout <= 8'b00111000; //  805 :  56 - 0x38
      12'h326: dout <= 8'b00011101; //  806 :  29 - 0x1d
      12'h327: dout <= 8'b00101111; //  807 :  47 - 0x2f
      12'h328: dout <= 8'b01000110; //  808 :  70 - 0x46 -- Sprite 0x65
      12'h329: dout <= 8'b11101011; //  809 : 235 - 0xeb
      12'h32A: dout <= 8'b01110001; //  810 : 113 - 0x71
      12'h32B: dout <= 8'b00111010; //  811 :  58 - 0x3a
      12'h32C: dout <= 8'b01101101; //  812 : 109 - 0x6d
      12'h32D: dout <= 8'b10111000; //  813 : 184 - 0xb8
      12'h32E: dout <= 8'b00011101; //  814 :  29 - 0x1d
      12'h32F: dout <= 8'b10101111; //  815 : 175 - 0xaf
      12'h330: dout <= 8'b01000110; //  816 :  70 - 0x46 -- Sprite 0x66
      12'h331: dout <= 8'b11101010; //  817 : 234 - 0xea
      12'h332: dout <= 8'b01110000; //  818 : 112 - 0x70
      12'h333: dout <= 8'b00111010; //  819 :  58 - 0x3a
      12'h334: dout <= 8'b01101100; //  820 : 108 - 0x6c
      12'h335: dout <= 8'b10111000; //  821 : 184 - 0xb8
      12'h336: dout <= 8'b00011100; //  822 :  28 - 0x1c
      12'h337: dout <= 8'b10101110; //  823 : 174 - 0xae
      12'h338: dout <= 8'b00000000; //  824 :   0 - 0x0 -- Sprite 0x67
      12'h339: dout <= 8'b01111111; //  825 : 127 - 0x7f
      12'h33A: dout <= 8'b01111111; //  826 : 127 - 0x7f
      12'h33B: dout <= 8'b00110011; //  827 :  51 - 0x33
      12'h33C: dout <= 8'b00000000; //  828 :   0 - 0x0
      12'h33D: dout <= 8'b00000000; //  829 :   0 - 0x0
      12'h33E: dout <= 8'b00000000; //  830 :   0 - 0x0
      12'h33F: dout <= 8'b00000000; //  831 :   0 - 0x0
      12'h340: dout <= 8'b00000000; //  832 :   0 - 0x0 -- Sprite 0x68
      12'h341: dout <= 8'b11111111; //  833 : 255 - 0xff
      12'h342: dout <= 8'b11111111; //  834 : 255 - 0xff
      12'h343: dout <= 8'b11111111; //  835 : 255 - 0xff
      12'h344: dout <= 8'b11001100; //  836 : 204 - 0xcc
      12'h345: dout <= 8'b00000000; //  837 :   0 - 0x0
      12'h346: dout <= 8'b00000000; //  838 :   0 - 0x0
      12'h347: dout <= 8'b00000000; //  839 :   0 - 0x0
      12'h348: dout <= 8'b00000000; //  840 :   0 - 0x0 -- Sprite 0x69
      12'h349: dout <= 8'b11111110; //  841 : 254 - 0xfe
      12'h34A: dout <= 8'b11111110; //  842 : 254 - 0xfe
      12'h34B: dout <= 8'b11110000; //  843 : 240 - 0xf0
      12'h34C: dout <= 8'b11000000; //  844 : 192 - 0xc0
      12'h34D: dout <= 8'b00000000; //  845 :   0 - 0x0
      12'h34E: dout <= 8'b00000000; //  846 :   0 - 0x0
      12'h34F: dout <= 8'b00000000; //  847 :   0 - 0x0
      12'h350: dout <= 8'b00000000; //  848 :   0 - 0x0 -- Sprite 0x6a
      12'h351: dout <= 8'b00000000; //  849 :   0 - 0x0
      12'h352: dout <= 8'b00000000; //  850 :   0 - 0x0
      12'h353: dout <= 8'b00000000; //  851 :   0 - 0x0
      12'h354: dout <= 8'b00000000; //  852 :   0 - 0x0
      12'h355: dout <= 8'b00000000; //  853 :   0 - 0x0
      12'h356: dout <= 8'b00000000; //  854 :   0 - 0x0
      12'h357: dout <= 8'b00000000; //  855 :   0 - 0x0
      12'h358: dout <= 8'b00111101; //  856 :  61 - 0x3d -- Sprite 0x6b
      12'h359: dout <= 8'b01111111; //  857 : 127 - 0x7f
      12'h35A: dout <= 8'b01111111; //  858 : 127 - 0x7f
      12'h35B: dout <= 8'b01111111; //  859 : 127 - 0x7f
      12'h35C: dout <= 8'b00111111; //  860 :  63 - 0x3f
      12'h35D: dout <= 8'b00001111; //  861 :  15 - 0xf
      12'h35E: dout <= 8'b00000000; //  862 :   0 - 0x0
      12'h35F: dout <= 8'b00000000; //  863 :   0 - 0x0
      12'h360: dout <= 8'b11111111; //  864 : 255 - 0xff -- Sprite 0x6c
      12'h361: dout <= 8'b11111111; //  865 : 255 - 0xff
      12'h362: dout <= 8'b11111111; //  866 : 255 - 0xff
      12'h363: dout <= 8'b11111111; //  867 : 255 - 0xff
      12'h364: dout <= 8'b11111111; //  868 : 255 - 0xff
      12'h365: dout <= 8'b11111111; //  869 : 255 - 0xff
      12'h366: dout <= 8'b11111110; //  870 : 254 - 0xfe
      12'h367: dout <= 8'b00000000; //  871 :   0 - 0x0
      12'h368: dout <= 8'b00000000; //  872 :   0 - 0x0 -- Sprite 0x6d
      12'h369: dout <= 8'b00000000; //  873 :   0 - 0x0
      12'h36A: dout <= 8'b00000000; //  874 :   0 - 0x0
      12'h36B: dout <= 8'b00000000; //  875 :   0 - 0x0
      12'h36C: dout <= 8'b00000000; //  876 :   0 - 0x0
      12'h36D: dout <= 8'b00000000; //  877 :   0 - 0x0
      12'h36E: dout <= 8'b00000000; //  878 :   0 - 0x0
      12'h36F: dout <= 8'b00000000; //  879 :   0 - 0x0
      12'h370: dout <= 8'b00000000; //  880 :   0 - 0x0 -- Sprite 0x6e
      12'h371: dout <= 8'b00000000; //  881 :   0 - 0x0
      12'h372: dout <= 8'b00000000; //  882 :   0 - 0x0
      12'h373: dout <= 8'b00000000; //  883 :   0 - 0x0
      12'h374: dout <= 8'b00000000; //  884 :   0 - 0x0
      12'h375: dout <= 8'b00000000; //  885 :   0 - 0x0
      12'h376: dout <= 8'b00000000; //  886 :   0 - 0x0
      12'h377: dout <= 8'b00000000; //  887 :   0 - 0x0
      12'h378: dout <= 8'b10111000; //  888 : 184 - 0xb8 -- Sprite 0x6f
      12'h379: dout <= 8'b11111100; //  889 : 252 - 0xfc
      12'h37A: dout <= 8'b11111110; //  890 : 254 - 0xfe
      12'h37B: dout <= 8'b11111110; //  891 : 254 - 0xfe
      12'h37C: dout <= 8'b11111100; //  892 : 252 - 0xfc
      12'h37D: dout <= 8'b11110000; //  893 : 240 - 0xf0
      12'h37E: dout <= 8'b00000000; //  894 :   0 - 0x0
      12'h37F: dout <= 8'b00000000; //  895 :   0 - 0x0
      12'h380: dout <= 8'b00000000; //  896 :   0 - 0x0 -- Sprite 0x70
      12'h381: dout <= 8'b00111111; //  897 :  63 - 0x3f
      12'h382: dout <= 8'b01111111; //  898 : 127 - 0x7f
      12'h383: dout <= 8'b01111111; //  899 : 127 - 0x7f
      12'h384: dout <= 8'b00011100; //  900 :  28 - 0x1c
      12'h385: dout <= 8'b00000000; //  901 :   0 - 0x0
      12'h386: dout <= 8'b00000000; //  902 :   0 - 0x0
      12'h387: dout <= 8'b00000000; //  903 :   0 - 0x0
      12'h388: dout <= 8'b00000000; //  904 :   0 - 0x0 -- Sprite 0x71
      12'h389: dout <= 8'b11111111; //  905 : 255 - 0xff
      12'h38A: dout <= 8'b11111111; //  906 : 255 - 0xff
      12'h38B: dout <= 8'b11111111; //  907 : 255 - 0xff
      12'h38C: dout <= 8'b11111111; //  908 : 255 - 0xff
      12'h38D: dout <= 8'b00111100; //  909 :  60 - 0x3c
      12'h38E: dout <= 8'b00000000; //  910 :   0 - 0x0
      12'h38F: dout <= 8'b00000000; //  911 :   0 - 0x0
      12'h390: dout <= 8'b00000000; //  912 :   0 - 0x0 -- Sprite 0x72
      12'h391: dout <= 8'b11111100; //  913 : 252 - 0xfc
      12'h392: dout <= 8'b11111110; //  914 : 254 - 0xfe
      12'h393: dout <= 8'b11111110; //  915 : 254 - 0xfe
      12'h394: dout <= 8'b00111000; //  916 :  56 - 0x38
      12'h395: dout <= 8'b00000000; //  917 :   0 - 0x0
      12'h396: dout <= 8'b00000000; //  918 :   0 - 0x0
      12'h397: dout <= 8'b00000000; //  919 :   0 - 0x0
      12'h398: dout <= 8'b11111111; //  920 : 255 - 0xff -- Sprite 0x73
      12'h399: dout <= 8'b11111111; //  921 : 255 - 0xff
      12'h39A: dout <= 8'b11111101; //  922 : 253 - 0xfd
      12'h39B: dout <= 8'b11111111; //  923 : 255 - 0xff
      12'h39C: dout <= 8'b10111111; //  924 : 191 - 0xbf
      12'h39D: dout <= 8'b11111111; //  925 : 255 - 0xff
      12'h39E: dout <= 8'b11111111; //  926 : 255 - 0xff
      12'h39F: dout <= 8'b11110111; //  927 : 247 - 0xf7
      12'h3A0: dout <= 8'b01000110; //  928 :  70 - 0x46 -- Sprite 0x74
      12'h3A1: dout <= 8'b01101011; //  929 : 107 - 0x6b
      12'h3A2: dout <= 8'b01110001; //  930 : 113 - 0x71
      12'h3A3: dout <= 8'b00111010; //  931 :  58 - 0x3a
      12'h3A4: dout <= 8'b01101101; //  932 : 109 - 0x6d
      12'h3A5: dout <= 8'b00111000; //  933 :  56 - 0x38
      12'h3A6: dout <= 8'b00011101; //  934 :  29 - 0x1d
      12'h3A7: dout <= 8'b00000000; //  935 :   0 - 0x0
      12'h3A8: dout <= 8'b01000110; //  936 :  70 - 0x46 -- Sprite 0x75
      12'h3A9: dout <= 8'b11101011; //  937 : 235 - 0xeb
      12'h3AA: dout <= 8'b01110001; //  938 : 113 - 0x71
      12'h3AB: dout <= 8'b00111010; //  939 :  58 - 0x3a
      12'h3AC: dout <= 8'b01101101; //  940 : 109 - 0x6d
      12'h3AD: dout <= 8'b10111000; //  941 : 184 - 0xb8
      12'h3AE: dout <= 8'b00011101; //  942 :  29 - 0x1d
      12'h3AF: dout <= 8'b00000000; //  943 :   0 - 0x0
      12'h3B0: dout <= 8'b01000110; //  944 :  70 - 0x46 -- Sprite 0x76
      12'h3B1: dout <= 8'b11101010; //  945 : 234 - 0xea
      12'h3B2: dout <= 8'b01110000; //  946 : 112 - 0x70
      12'h3B3: dout <= 8'b00111010; //  947 :  58 - 0x3a
      12'h3B4: dout <= 8'b01101100; //  948 : 108 - 0x6c
      12'h3B5: dout <= 8'b10111000; //  949 : 184 - 0xb8
      12'h3B6: dout <= 8'b00011100; //  950 :  28 - 0x1c
      12'h3B7: dout <= 8'b00000000; //  951 :   0 - 0x0
      12'h3B8: dout <= 8'b10000001; //  952 : 129 - 0x81 -- Sprite 0x77
      12'h3B9: dout <= 8'b11111111; //  953 : 255 - 0xff
      12'h3BA: dout <= 8'b11111101; //  954 : 253 - 0xfd
      12'h3BB: dout <= 8'b11111111; //  955 : 255 - 0xff
      12'h3BC: dout <= 8'b10111111; //  956 : 191 - 0xbf
      12'h3BD: dout <= 8'b11111111; //  957 : 255 - 0xff
      12'h3BE: dout <= 8'b11111111; //  958 : 255 - 0xff
      12'h3BF: dout <= 8'b11110111; //  959 : 247 - 0xf7
      12'h3C0: dout <= 8'b00000000; //  960 :   0 - 0x0 -- Sprite 0x78
      12'h3C1: dout <= 8'b00000000; //  961 :   0 - 0x0
      12'h3C2: dout <= 8'b00000000; //  962 :   0 - 0x0
      12'h3C3: dout <= 8'b00000000; //  963 :   0 - 0x0
      12'h3C4: dout <= 8'b00000000; //  964 :   0 - 0x0
      12'h3C5: dout <= 8'b00000000; //  965 :   0 - 0x0
      12'h3C6: dout <= 8'b00000000; //  966 :   0 - 0x0
      12'h3C7: dout <= 8'b00000000; //  967 :   0 - 0x0
      12'h3C8: dout <= 8'b00000000; //  968 :   0 - 0x0 -- Sprite 0x79
      12'h3C9: dout <= 8'b00000000; //  969 :   0 - 0x0
      12'h3CA: dout <= 8'b00000000; //  970 :   0 - 0x0
      12'h3CB: dout <= 8'b00000000; //  971 :   0 - 0x0
      12'h3CC: dout <= 8'b00000000; //  972 :   0 - 0x0
      12'h3CD: dout <= 8'b00000000; //  973 :   0 - 0x0
      12'h3CE: dout <= 8'b00000000; //  974 :   0 - 0x0
      12'h3CF: dout <= 8'b00000000; //  975 :   0 - 0x0
      12'h3D0: dout <= 8'b00000000; //  976 :   0 - 0x0 -- Sprite 0x7a
      12'h3D1: dout <= 8'b00000000; //  977 :   0 - 0x0
      12'h3D2: dout <= 8'b00000000; //  978 :   0 - 0x0
      12'h3D3: dout <= 8'b00000000; //  979 :   0 - 0x0
      12'h3D4: dout <= 8'b00000000; //  980 :   0 - 0x0
      12'h3D5: dout <= 8'b00000000; //  981 :   0 - 0x0
      12'h3D6: dout <= 8'b00000000; //  982 :   0 - 0x0
      12'h3D7: dout <= 8'b00000000; //  983 :   0 - 0x0
      12'h3D8: dout <= 8'b00000000; //  984 :   0 - 0x0 -- Sprite 0x7b
      12'h3D9: dout <= 8'b00000000; //  985 :   0 - 0x0
      12'h3DA: dout <= 8'b00000000; //  986 :   0 - 0x0
      12'h3DB: dout <= 8'b00000000; //  987 :   0 - 0x0
      12'h3DC: dout <= 8'b00000000; //  988 :   0 - 0x0
      12'h3DD: dout <= 8'b00000000; //  989 :   0 - 0x0
      12'h3DE: dout <= 8'b00000000; //  990 :   0 - 0x0
      12'h3DF: dout <= 8'b00000000; //  991 :   0 - 0x0
      12'h3E0: dout <= 8'b00000000; //  992 :   0 - 0x0 -- Sprite 0x7c
      12'h3E1: dout <= 8'b00100010; //  993 :  34 - 0x22
      12'h3E2: dout <= 8'b01110111; //  994 : 119 - 0x77
      12'h3E3: dout <= 8'b11111111; //  995 : 255 - 0xff
      12'h3E4: dout <= 8'b11111011; //  996 : 251 - 0xfb
      12'h3E5: dout <= 8'b11110101; //  997 : 245 - 0xf5
      12'h3E6: dout <= 8'b11101111; //  998 : 239 - 0xef
      12'h3E7: dout <= 8'b11111111; //  999 : 255 - 0xff
      12'h3E8: dout <= 8'b00000000; // 1000 :   0 - 0x0 -- Sprite 0x7d
      12'h3E9: dout <= 8'b01110011; // 1001 : 115 - 0x73
      12'h3EA: dout <= 8'b11111111; // 1002 : 255 - 0xff
      12'h3EB: dout <= 8'b11111111; // 1003 : 255 - 0xff
      12'h3EC: dout <= 8'b11111011; // 1004 : 251 - 0xfb
      12'h3ED: dout <= 8'b11111101; // 1005 : 253 - 0xfd
      12'h3EE: dout <= 8'b11101111; // 1006 : 239 - 0xef
      12'h3EF: dout <= 8'b11111111; // 1007 : 255 - 0xff
      12'h3F0: dout <= 8'b11011111; // 1008 : 223 - 0xdf -- Sprite 0x7e
      12'h3F1: dout <= 8'b10101111; // 1009 : 175 - 0xaf
      12'h3F2: dout <= 8'b01111111; // 1010 : 127 - 0x7f
      12'h3F3: dout <= 8'b11111111; // 1011 : 255 - 0xff
      12'h3F4: dout <= 8'b11111011; // 1012 : 251 - 0xfb
      12'h3F5: dout <= 8'b11110101; // 1013 : 245 - 0xf5
      12'h3F6: dout <= 8'b11101111; // 1014 : 239 - 0xef
      12'h3F7: dout <= 8'b11111111; // 1015 : 255 - 0xff
      12'h3F8: dout <= 8'b00000000; // 1016 :   0 - 0x0 -- Sprite 0x7f
      12'h3F9: dout <= 8'b10101111; // 1017 : 175 - 0xaf
      12'h3FA: dout <= 8'b01111111; // 1018 : 127 - 0x7f
      12'h3FB: dout <= 8'b11111111; // 1019 : 255 - 0xff
      12'h3FC: dout <= 8'b11111011; // 1020 : 251 - 0xfb
      12'h3FD: dout <= 8'b11110101; // 1021 : 245 - 0xf5
      12'h3FE: dout <= 8'b11101111; // 1022 : 239 - 0xef
      12'h3FF: dout <= 8'b11111111; // 1023 : 255 - 0xff
      12'h400: dout <= 8'b00000000; // 1024 :   0 - 0x0 -- Sprite 0x80
      12'h401: dout <= 8'b01111111; // 1025 : 127 - 0x7f
      12'h402: dout <= 8'b00110000; // 1026 :  48 - 0x30
      12'h403: dout <= 8'b00110000; // 1027 :  48 - 0x30
      12'h404: dout <= 8'b00110000; // 1028 :  48 - 0x30
      12'h405: dout <= 8'b01111111; // 1029 : 127 - 0x7f
      12'h406: dout <= 8'b00110000; // 1030 :  48 - 0x30
      12'h407: dout <= 8'b00110000; // 1031 :  48 - 0x30
      12'h408: dout <= 8'b00000000; // 1032 :   0 - 0x0 -- Sprite 0x81
      12'h409: dout <= 8'b01111111; // 1033 : 127 - 0x7f
      12'h40A: dout <= 8'b00000000; // 1034 :   0 - 0x0
      12'h40B: dout <= 8'b01111111; // 1035 : 127 - 0x7f
      12'h40C: dout <= 8'b01111111; // 1036 : 127 - 0x7f
      12'h40D: dout <= 8'b00100000; // 1037 :  32 - 0x20
      12'h40E: dout <= 8'b01000000; // 1038 :  64 - 0x40
      12'h40F: dout <= 8'b00000000; // 1039 :   0 - 0x0
      12'h410: dout <= 8'b00000000; // 1040 :   0 - 0x0 -- Sprite 0x82
      12'h411: dout <= 8'b11111110; // 1041 : 254 - 0xfe
      12'h412: dout <= 8'b00001100; // 1042 :  12 - 0xc
      12'h413: dout <= 8'b00001100; // 1043 :  12 - 0xc
      12'h414: dout <= 8'b00001100; // 1044 :  12 - 0xc
      12'h415: dout <= 8'b11111110; // 1045 : 254 - 0xfe
      12'h416: dout <= 8'b00001100; // 1046 :  12 - 0xc
      12'h417: dout <= 8'b00001100; // 1047 :  12 - 0xc
      12'h418: dout <= 8'b00000000; // 1048 :   0 - 0x0 -- Sprite 0x83
      12'h419: dout <= 8'b11111111; // 1049 : 255 - 0xff
      12'h41A: dout <= 8'b00000000; // 1050 :   0 - 0x0
      12'h41B: dout <= 8'b11111111; // 1051 : 255 - 0xff
      12'h41C: dout <= 8'b11111111; // 1052 : 255 - 0xff
      12'h41D: dout <= 8'b00000000; // 1053 :   0 - 0x0
      12'h41E: dout <= 8'b00000000; // 1054 :   0 - 0x0
      12'h41F: dout <= 8'b00000000; // 1055 :   0 - 0x0
      12'h420: dout <= 8'b00000000; // 1056 :   0 - 0x0 -- Sprite 0x84
      12'h421: dout <= 8'b11111111; // 1057 : 255 - 0xff
      12'h422: dout <= 8'b11111111; // 1058 : 255 - 0xff
      12'h423: dout <= 8'b11111111; // 1059 : 255 - 0xff
      12'h424: dout <= 8'b11111111; // 1060 : 255 - 0xff
      12'h425: dout <= 8'b11101111; // 1061 : 239 - 0xef
      12'h426: dout <= 8'b10111011; // 1062 : 187 - 0xbb
      12'h427: dout <= 8'b00000000; // 1063 :   0 - 0x0
      12'h428: dout <= 8'b00000000; // 1064 :   0 - 0x0 -- Sprite 0x85
      12'h429: dout <= 8'b11111110; // 1065 : 254 - 0xfe
      12'h42A: dout <= 8'b00000000; // 1066 :   0 - 0x0
      12'h42B: dout <= 8'b11111110; // 1067 : 254 - 0xfe
      12'h42C: dout <= 8'b11111110; // 1068 : 254 - 0xfe
      12'h42D: dout <= 8'b00001100; // 1069 :  12 - 0xc
      12'h42E: dout <= 8'b00000010; // 1070 :   2 - 0x2
      12'h42F: dout <= 8'b00000000; // 1071 :   0 - 0x0
      12'h430: dout <= 8'b00000000; // 1072 :   0 - 0x0 -- Sprite 0x86
      12'h431: dout <= 8'b00000000; // 1073 :   0 - 0x0
      12'h432: dout <= 8'b00000000; // 1074 :   0 - 0x0
      12'h433: dout <= 8'b00000000; // 1075 :   0 - 0x0
      12'h434: dout <= 8'b00000000; // 1076 :   0 - 0x0
      12'h435: dout <= 8'b00000000; // 1077 :   0 - 0x0
      12'h436: dout <= 8'b00000000; // 1078 :   0 - 0x0
      12'h437: dout <= 8'b00000000; // 1079 :   0 - 0x0
      12'h438: dout <= 8'b00000000; // 1080 :   0 - 0x0 -- Sprite 0x87
      12'h439: dout <= 8'b00000000; // 1081 :   0 - 0x0
      12'h43A: dout <= 8'b00000000; // 1082 :   0 - 0x0
      12'h43B: dout <= 8'b00000000; // 1083 :   0 - 0x0
      12'h43C: dout <= 8'b00000000; // 1084 :   0 - 0x0
      12'h43D: dout <= 8'b00000000; // 1085 :   0 - 0x0
      12'h43E: dout <= 8'b00000000; // 1086 :   0 - 0x0
      12'h43F: dout <= 8'b00000000; // 1087 :   0 - 0x0
      12'h440: dout <= 8'b00000000; // 1088 :   0 - 0x0 -- Sprite 0x88
      12'h441: dout <= 8'b00000111; // 1089 :   7 - 0x7
      12'h442: dout <= 8'b00011111; // 1090 :  31 - 0x1f
      12'h443: dout <= 8'b00111100; // 1091 :  60 - 0x3c
      12'h444: dout <= 8'b00110001; // 1092 :  49 - 0x31
      12'h445: dout <= 8'b01110100; // 1093 : 116 - 0x74
      12'h446: dout <= 8'b01100101; // 1094 : 101 - 0x65
      12'h447: dout <= 8'b01101010; // 1095 : 106 - 0x6a
      12'h448: dout <= 8'b01100100; // 1096 : 100 - 0x64 -- Sprite 0x89
      12'h449: dout <= 8'b01101101; // 1097 : 109 - 0x6d
      12'h44A: dout <= 8'b01110010; // 1098 : 114 - 0x72
      12'h44B: dout <= 8'b00110000; // 1099 :  48 - 0x30
      12'h44C: dout <= 8'b00111100; // 1100 :  60 - 0x3c
      12'h44D: dout <= 8'b00011111; // 1101 :  31 - 0x1f
      12'h44E: dout <= 8'b00000111; // 1102 :   7 - 0x7
      12'h44F: dout <= 8'b00000000; // 1103 :   0 - 0x0
      12'h450: dout <= 8'b00000000; // 1104 :   0 - 0x0 -- Sprite 0x8a
      12'h451: dout <= 8'b11100000; // 1105 : 224 - 0xe0
      12'h452: dout <= 8'b11111000; // 1106 : 248 - 0xf8
      12'h453: dout <= 8'b00111100; // 1107 :  60 - 0x3c
      12'h454: dout <= 8'b01001100; // 1108 :  76 - 0x4c
      12'h455: dout <= 8'b01101110; // 1109 : 110 - 0x6e
      12'h456: dout <= 8'b00100110; // 1110 :  38 - 0x26
      12'h457: dout <= 8'b01000110; // 1111 :  70 - 0x46
      12'h458: dout <= 8'b10010110; // 1112 : 150 - 0x96 -- Sprite 0x8b
      12'h459: dout <= 8'b01100110; // 1113 : 102 - 0x66
      12'h45A: dout <= 8'b10101110; // 1114 : 174 - 0xae
      12'h45B: dout <= 8'b01001100; // 1115 :  76 - 0x4c
      12'h45C: dout <= 8'b00111100; // 1116 :  60 - 0x3c
      12'h45D: dout <= 8'b11111000; // 1117 : 248 - 0xf8
      12'h45E: dout <= 8'b11100000; // 1118 : 224 - 0xe0
      12'h45F: dout <= 8'b00000000; // 1119 :   0 - 0x0
      12'h460: dout <= 8'b00000000; // 1120 :   0 - 0x0 -- Sprite 0x8c
      12'h461: dout <= 8'b00000111; // 1121 :   7 - 0x7
      12'h462: dout <= 8'b00011111; // 1122 :  31 - 0x1f
      12'h463: dout <= 8'b00111111; // 1123 :  63 - 0x3f
      12'h464: dout <= 8'b00111111; // 1124 :  63 - 0x3f
      12'h465: dout <= 8'b01111111; // 1125 : 127 - 0x7f
      12'h466: dout <= 8'b01111111; // 1126 : 127 - 0x7f
      12'h467: dout <= 8'b01111111; // 1127 : 127 - 0x7f
      12'h468: dout <= 8'b01111111; // 1128 : 127 - 0x7f -- Sprite 0x8d
      12'h469: dout <= 8'b01111111; // 1129 : 127 - 0x7f
      12'h46A: dout <= 8'b01111111; // 1130 : 127 - 0x7f
      12'h46B: dout <= 8'b00111111; // 1131 :  63 - 0x3f
      12'h46C: dout <= 8'b00111111; // 1132 :  63 - 0x3f
      12'h46D: dout <= 8'b00011111; // 1133 :  31 - 0x1f
      12'h46E: dout <= 8'b00000111; // 1134 :   7 - 0x7
      12'h46F: dout <= 8'b00000000; // 1135 :   0 - 0x0
      12'h470: dout <= 8'b00000000; // 1136 :   0 - 0x0 -- Sprite 0x8e
      12'h471: dout <= 8'b11100000; // 1137 : 224 - 0xe0
      12'h472: dout <= 8'b11111000; // 1138 : 248 - 0xf8
      12'h473: dout <= 8'b11111100; // 1139 : 252 - 0xfc
      12'h474: dout <= 8'b11111100; // 1140 : 252 - 0xfc
      12'h475: dout <= 8'b11111110; // 1141 : 254 - 0xfe
      12'h476: dout <= 8'b11111110; // 1142 : 254 - 0xfe
      12'h477: dout <= 8'b11111110; // 1143 : 254 - 0xfe
      12'h478: dout <= 8'b11111110; // 1144 : 254 - 0xfe -- Sprite 0x8f
      12'h479: dout <= 8'b11111110; // 1145 : 254 - 0xfe
      12'h47A: dout <= 8'b11111110; // 1146 : 254 - 0xfe
      12'h47B: dout <= 8'b11111100; // 1147 : 252 - 0xfc
      12'h47C: dout <= 8'b11111100; // 1148 : 252 - 0xfc
      12'h47D: dout <= 8'b11111000; // 1149 : 248 - 0xf8
      12'h47E: dout <= 8'b11100000; // 1150 : 224 - 0xe0
      12'h47F: dout <= 8'b00000000; // 1151 :   0 - 0x0
      12'h480: dout <= 8'b00000000; // 1152 :   0 - 0x0 -- Sprite 0x90
      12'h481: dout <= 8'b00000000; // 1153 :   0 - 0x0
      12'h482: dout <= 8'b00000000; // 1154 :   0 - 0x0
      12'h483: dout <= 8'b00000000; // 1155 :   0 - 0x0
      12'h484: dout <= 8'b00010000; // 1156 :  16 - 0x10
      12'h485: dout <= 8'b00011100; // 1157 :  28 - 0x1c
      12'h486: dout <= 8'b00001110; // 1158 :  14 - 0xe
      12'h487: dout <= 8'b00000111; // 1159 :   7 - 0x7
      12'h488: dout <= 8'b00000011; // 1160 :   3 - 0x3 -- Sprite 0x91
      12'h489: dout <= 8'b00000001; // 1161 :   1 - 0x1
      12'h48A: dout <= 8'b00110000; // 1162 :  48 - 0x30
      12'h48B: dout <= 8'b00001111; // 1163 :  15 - 0xf
      12'h48C: dout <= 8'b00000011; // 1164 :   3 - 0x3
      12'h48D: dout <= 8'b00000000; // 1165 :   0 - 0x0
      12'h48E: dout <= 8'b01111111; // 1166 : 127 - 0x7f
      12'h48F: dout <= 8'b00000000; // 1167 :   0 - 0x0
      12'h490: dout <= 8'b00000000; // 1168 :   0 - 0x0 -- Sprite 0x92
      12'h491: dout <= 8'b01000010; // 1169 :  66 - 0x42
      12'h492: dout <= 8'b01000010; // 1170 :  66 - 0x42
      12'h493: dout <= 8'b01100110; // 1171 : 102 - 0x66
      12'h494: dout <= 8'b01100110; // 1172 : 102 - 0x66
      12'h495: dout <= 8'b01100110; // 1173 : 102 - 0x66
      12'h496: dout <= 8'b11111110; // 1174 : 254 - 0xfe
      12'h497: dout <= 8'b11111111; // 1175 : 255 - 0xff
      12'h498: dout <= 8'b01111110; // 1176 : 126 - 0x7e -- Sprite 0x93
      12'h499: dout <= 8'b01111110; // 1177 : 126 - 0x7e
      12'h49A: dout <= 8'b01111110; // 1178 : 126 - 0x7e
      12'h49B: dout <= 8'b01111110; // 1179 : 126 - 0x7e
      12'h49C: dout <= 8'b01111110; // 1180 : 126 - 0x7e
      12'h49D: dout <= 8'b01111110; // 1181 : 126 - 0x7e
      12'h49E: dout <= 8'b01111110; // 1182 : 126 - 0x7e
      12'h49F: dout <= 8'b01111110; // 1183 : 126 - 0x7e
      12'h4A0: dout <= 8'b00000000; // 1184 :   0 - 0x0 -- Sprite 0x94
      12'h4A1: dout <= 8'b00000000; // 1185 :   0 - 0x0
      12'h4A2: dout <= 8'b00000000; // 1186 :   0 - 0x0
      12'h4A3: dout <= 8'b00000000; // 1187 :   0 - 0x0
      12'h4A4: dout <= 8'b00001000; // 1188 :   8 - 0x8
      12'h4A5: dout <= 8'b00111000; // 1189 :  56 - 0x38
      12'h4A6: dout <= 8'b01110000; // 1190 : 112 - 0x70
      12'h4A7: dout <= 8'b11100000; // 1191 : 224 - 0xe0
      12'h4A8: dout <= 8'b11000000; // 1192 : 192 - 0xc0 -- Sprite 0x95
      12'h4A9: dout <= 8'b10000000; // 1193 : 128 - 0x80
      12'h4AA: dout <= 8'b00001100; // 1194 :  12 - 0xc
      12'h4AB: dout <= 8'b11110000; // 1195 : 240 - 0xf0
      12'h4AC: dout <= 8'b11000000; // 1196 : 192 - 0xc0
      12'h4AD: dout <= 8'b00000000; // 1197 :   0 - 0x0
      12'h4AE: dout <= 8'b11111110; // 1198 : 254 - 0xfe
      12'h4AF: dout <= 8'b00000000; // 1199 :   0 - 0x0
      12'h4B0: dout <= 8'b00000000; // 1200 :   0 - 0x0 -- Sprite 0x96
      12'h4B1: dout <= 8'b00111111; // 1201 :  63 - 0x3f
      12'h4B2: dout <= 8'b01111111; // 1202 : 127 - 0x7f
      12'h4B3: dout <= 8'b01111111; // 1203 : 127 - 0x7f
      12'h4B4: dout <= 8'b01111111; // 1204 : 127 - 0x7f
      12'h4B5: dout <= 8'b01111111; // 1205 : 127 - 0x7f
      12'h4B6: dout <= 8'b01111111; // 1206 : 127 - 0x7f
      12'h4B7: dout <= 8'b01111111; // 1207 : 127 - 0x7f
      12'h4B8: dout <= 8'b01111111; // 1208 : 127 - 0x7f -- Sprite 0x97
      12'h4B9: dout <= 8'b01111111; // 1209 : 127 - 0x7f
      12'h4BA: dout <= 8'b00111111; // 1210 :  63 - 0x3f
      12'h4BB: dout <= 8'b01111111; // 1211 : 127 - 0x7f
      12'h4BC: dout <= 8'b01111111; // 1212 : 127 - 0x7f
      12'h4BD: dout <= 8'b01111111; // 1213 : 127 - 0x7f
      12'h4BE: dout <= 8'b01111111; // 1214 : 127 - 0x7f
      12'h4BF: dout <= 8'b01111111; // 1215 : 127 - 0x7f
      12'h4C0: dout <= 8'b00000000; // 1216 :   0 - 0x0 -- Sprite 0x98
      12'h4C1: dout <= 8'b11011111; // 1217 : 223 - 0xdf
      12'h4C2: dout <= 8'b11111111; // 1218 : 255 - 0xff
      12'h4C3: dout <= 8'b11111111; // 1219 : 255 - 0xff
      12'h4C4: dout <= 8'b11111111; // 1220 : 255 - 0xff
      12'h4C5: dout <= 8'b11111111; // 1221 : 255 - 0xff
      12'h4C6: dout <= 8'b11111111; // 1222 : 255 - 0xff
      12'h4C7: dout <= 8'b11111111; // 1223 : 255 - 0xff
      12'h4C8: dout <= 8'b11111111; // 1224 : 255 - 0xff -- Sprite 0x99
      12'h4C9: dout <= 8'b11111111; // 1225 : 255 - 0xff
      12'h4CA: dout <= 8'b10111111; // 1226 : 191 - 0xbf
      12'h4CB: dout <= 8'b11111111; // 1227 : 255 - 0xff
      12'h4CC: dout <= 8'b11111111; // 1228 : 255 - 0xff
      12'h4CD: dout <= 8'b11111111; // 1229 : 255 - 0xff
      12'h4CE: dout <= 8'b11111111; // 1230 : 255 - 0xff
      12'h4CF: dout <= 8'b11111111; // 1231 : 255 - 0xff
      12'h4D0: dout <= 8'b00000000; // 1232 :   0 - 0x0 -- Sprite 0x9a
      12'h4D1: dout <= 8'b10111100; // 1233 : 188 - 0xbc
      12'h4D2: dout <= 8'b11111110; // 1234 : 254 - 0xfe
      12'h4D3: dout <= 8'b11111110; // 1235 : 254 - 0xfe
      12'h4D4: dout <= 8'b11111110; // 1236 : 254 - 0xfe
      12'h4D5: dout <= 8'b11111110; // 1237 : 254 - 0xfe
      12'h4D6: dout <= 8'b11111110; // 1238 : 254 - 0xfe
      12'h4D7: dout <= 8'b11111110; // 1239 : 254 - 0xfe
      12'h4D8: dout <= 8'b11111110; // 1240 : 254 - 0xfe -- Sprite 0x9b
      12'h4D9: dout <= 8'b11111110; // 1241 : 254 - 0xfe
      12'h4DA: dout <= 8'b10111110; // 1242 : 190 - 0xbe
      12'h4DB: dout <= 8'b11111110; // 1243 : 254 - 0xfe
      12'h4DC: dout <= 8'b11111110; // 1244 : 254 - 0xfe
      12'h4DD: dout <= 8'b11111110; // 1245 : 254 - 0xfe
      12'h4DE: dout <= 8'b11111110; // 1246 : 254 - 0xfe
      12'h4DF: dout <= 8'b11111110; // 1247 : 254 - 0xfe
      12'h4E0: dout <= 8'b00000000; // 1248 :   0 - 0x0 -- Sprite 0x9c
      12'h4E1: dout <= 8'b00111111; // 1249 :  63 - 0x3f
      12'h4E2: dout <= 8'b01011111; // 1250 :  95 - 0x5f
      12'h4E3: dout <= 8'b01101111; // 1251 : 111 - 0x6f
      12'h4E4: dout <= 8'b01110111; // 1252 : 119 - 0x77
      12'h4E5: dout <= 8'b01111011; // 1253 : 123 - 0x7b
      12'h4E6: dout <= 8'b00010101; // 1254 :  21 - 0x15
      12'h4E7: dout <= 8'b00000000; // 1255 :   0 - 0x0
      12'h4E8: dout <= 8'b00000000; // 1256 :   0 - 0x0 -- Sprite 0x9d
      12'h4E9: dout <= 8'b10111110; // 1257 : 190 - 0xbe
      12'h4EA: dout <= 8'b11011110; // 1258 : 222 - 0xde
      12'h4EB: dout <= 8'b11101110; // 1259 : 238 - 0xee
      12'h4EC: dout <= 8'b11110110; // 1260 : 246 - 0xf6
      12'h4ED: dout <= 8'b11111010; // 1261 : 250 - 0xfa
      12'h4EE: dout <= 8'b01010100; // 1262 :  84 - 0x54
      12'h4EF: dout <= 8'b00000000; // 1263 :   0 - 0x0
      12'h4F0: dout <= 8'b00000000; // 1264 :   0 - 0x0 -- Sprite 0x9e
      12'h4F1: dout <= 8'b10111111; // 1265 : 191 - 0xbf
      12'h4F2: dout <= 8'b11011111; // 1266 : 223 - 0xdf
      12'h4F3: dout <= 8'b11101111; // 1267 : 239 - 0xef
      12'h4F4: dout <= 8'b11110111; // 1268 : 247 - 0xf7
      12'h4F5: dout <= 8'b11111011; // 1269 : 251 - 0xfb
      12'h4F6: dout <= 8'b01010101; // 1270 :  85 - 0x55
      12'h4F7: dout <= 8'b00000000; // 1271 :   0 - 0x0
      12'h4F8: dout <= 8'b00000000; // 1272 :   0 - 0x0 -- Sprite 0x9f
      12'h4F9: dout <= 8'b00000000; // 1273 :   0 - 0x0
      12'h4FA: dout <= 8'b00000000; // 1274 :   0 - 0x0
      12'h4FB: dout <= 8'b00000000; // 1275 :   0 - 0x0
      12'h4FC: dout <= 8'b00000000; // 1276 :   0 - 0x0
      12'h4FD: dout <= 8'b00000000; // 1277 :   0 - 0x0
      12'h4FE: dout <= 8'b00000000; // 1278 :   0 - 0x0
      12'h4FF: dout <= 8'b00000000; // 1279 :   0 - 0x0
      12'h500: dout <= 8'b00000000; // 1280 :   0 - 0x0 -- Sprite 0xa0
      12'h501: dout <= 8'b01111111; // 1281 : 127 - 0x7f
      12'h502: dout <= 8'b00000000; // 1282 :   0 - 0x0
      12'h503: dout <= 8'b00000001; // 1283 :   1 - 0x1
      12'h504: dout <= 8'b00000001; // 1284 :   1 - 0x1
      12'h505: dout <= 8'b00000001; // 1285 :   1 - 0x1
      12'h506: dout <= 8'b00000001; // 1286 :   1 - 0x1
      12'h507: dout <= 8'b00000001; // 1287 :   1 - 0x1
      12'h508: dout <= 8'b00000001; // 1288 :   1 - 0x1 -- Sprite 0xa1
      12'h509: dout <= 8'b00000001; // 1289 :   1 - 0x1
      12'h50A: dout <= 8'b00000001; // 1290 :   1 - 0x1
      12'h50B: dout <= 8'b00000001; // 1291 :   1 - 0x1
      12'h50C: dout <= 8'b00000001; // 1292 :   1 - 0x1
      12'h50D: dout <= 8'b00000001; // 1293 :   1 - 0x1
      12'h50E: dout <= 8'b00000001; // 1294 :   1 - 0x1
      12'h50F: dout <= 8'b00000001; // 1295 :   1 - 0x1
      12'h510: dout <= 8'b00000000; // 1296 :   0 - 0x0 -- Sprite 0xa2
      12'h511: dout <= 8'b11111110; // 1297 : 254 - 0xfe
      12'h512: dout <= 8'b00000000; // 1298 :   0 - 0x0
      12'h513: dout <= 8'b10000000; // 1299 : 128 - 0x80
      12'h514: dout <= 8'b10000000; // 1300 : 128 - 0x80
      12'h515: dout <= 8'b10000000; // 1301 : 128 - 0x80
      12'h516: dout <= 8'b10000000; // 1302 : 128 - 0x80
      12'h517: dout <= 8'b10000000; // 1303 : 128 - 0x80
      12'h518: dout <= 8'b10000000; // 1304 : 128 - 0x80 -- Sprite 0xa3
      12'h519: dout <= 8'b10000000; // 1305 : 128 - 0x80
      12'h51A: dout <= 8'b10000000; // 1306 : 128 - 0x80
      12'h51B: dout <= 8'b10000000; // 1307 : 128 - 0x80
      12'h51C: dout <= 8'b10000000; // 1308 : 128 - 0x80
      12'h51D: dout <= 8'b10000000; // 1309 : 128 - 0x80
      12'h51E: dout <= 8'b10000000; // 1310 : 128 - 0x80
      12'h51F: dout <= 8'b10000000; // 1311 : 128 - 0x80
      12'h520: dout <= 8'b00000000; // 1312 :   0 - 0x0 -- Sprite 0xa4
      12'h521: dout <= 8'b00110000; // 1313 :  48 - 0x30
      12'h522: dout <= 8'b00111000; // 1314 :  56 - 0x38
      12'h523: dout <= 8'b01111000; // 1315 : 120 - 0x78
      12'h524: dout <= 8'b01111100; // 1316 : 124 - 0x7c
      12'h525: dout <= 8'b01111101; // 1317 : 125 - 0x7d
      12'h526: dout <= 8'b00011101; // 1318 :  29 - 0x1d
      12'h527: dout <= 8'b00001101; // 1319 :  13 - 0xd
      12'h528: dout <= 8'b00001101; // 1320 :  13 - 0xd -- Sprite 0xa5
      12'h529: dout <= 8'b00011101; // 1321 :  29 - 0x1d
      12'h52A: dout <= 8'b00111101; // 1322 :  61 - 0x3d
      12'h52B: dout <= 8'b00111111; // 1323 :  63 - 0x3f
      12'h52C: dout <= 8'b00111111; // 1324 :  63 - 0x3f
      12'h52D: dout <= 8'b00011111; // 1325 :  31 - 0x1f
      12'h52E: dout <= 8'b00000001; // 1326 :   1 - 0x1
      12'h52F: dout <= 8'b00000000; // 1327 :   0 - 0x0
      12'h530: dout <= 8'b00000000; // 1328 :   0 - 0x0 -- Sprite 0xa6
      12'h531: dout <= 8'b00000000; // 1329 :   0 - 0x0
      12'h532: dout <= 8'b11100000; // 1330 : 224 - 0xe0
      12'h533: dout <= 8'b11111000; // 1331 : 248 - 0xf8
      12'h534: dout <= 8'b11111000; // 1332 : 248 - 0xf8
      12'h535: dout <= 8'b11110000; // 1333 : 240 - 0xf0
      12'h536: dout <= 8'b11000000; // 1334 : 192 - 0xc0
      12'h537: dout <= 8'b11000000; // 1335 : 192 - 0xc0
      12'h538: dout <= 8'b11000000; // 1336 : 192 - 0xc0 -- Sprite 0xa7
      12'h539: dout <= 8'b11110000; // 1337 : 240 - 0xf0
      12'h53A: dout <= 8'b11110000; // 1338 : 240 - 0xf0
      12'h53B: dout <= 8'b11000000; // 1339 : 192 - 0xc0
      12'h53C: dout <= 8'b11000000; // 1340 : 192 - 0xc0
      12'h53D: dout <= 8'b11000000; // 1341 : 192 - 0xc0
      12'h53E: dout <= 8'b11000000; // 1342 : 192 - 0xc0
      12'h53F: dout <= 8'b00000000; // 1343 :   0 - 0x0
      12'h540: dout <= 8'b00000000; // 1344 :   0 - 0x0 -- Sprite 0xa8
      12'h541: dout <= 8'b01100000; // 1345 :  96 - 0x60
      12'h542: dout <= 8'b01100000; // 1346 :  96 - 0x60
      12'h543: dout <= 8'b01100000; // 1347 :  96 - 0x60
      12'h544: dout <= 8'b01100000; // 1348 :  96 - 0x60
      12'h545: dout <= 8'b01100000; // 1349 :  96 - 0x60
      12'h546: dout <= 8'b01100000; // 1350 :  96 - 0x60
      12'h547: dout <= 8'b01100000; // 1351 :  96 - 0x60
      12'h548: dout <= 8'b01100000; // 1352 :  96 - 0x60 -- Sprite 0xa9
      12'h549: dout <= 8'b01100000; // 1353 :  96 - 0x60
      12'h54A: dout <= 8'b01100000; // 1354 :  96 - 0x60
      12'h54B: dout <= 8'b01100000; // 1355 :  96 - 0x60
      12'h54C: dout <= 8'b01100000; // 1356 :  96 - 0x60
      12'h54D: dout <= 8'b01100000; // 1357 :  96 - 0x60
      12'h54E: dout <= 8'b01100000; // 1358 :  96 - 0x60
      12'h54F: dout <= 8'b00000000; // 1359 :   0 - 0x0
      12'h550: dout <= 8'b00000000; // 1360 :   0 - 0x0 -- Sprite 0xaa
      12'h551: dout <= 8'b00000000; // 1361 :   0 - 0x0
      12'h552: dout <= 8'b00000000; // 1362 :   0 - 0x0
      12'h553: dout <= 8'b00000000; // 1363 :   0 - 0x0
      12'h554: dout <= 8'b00000000; // 1364 :   0 - 0x0
      12'h555: dout <= 8'b00000000; // 1365 :   0 - 0x0
      12'h556: dout <= 8'b00000000; // 1366 :   0 - 0x0
      12'h557: dout <= 8'b00000000; // 1367 :   0 - 0x0
      12'h558: dout <= 8'b00000000; // 1368 :   0 - 0x0 -- Sprite 0xab
      12'h559: dout <= 8'b00000000; // 1369 :   0 - 0x0
      12'h55A: dout <= 8'b00000000; // 1370 :   0 - 0x0
      12'h55B: dout <= 8'b00000000; // 1371 :   0 - 0x0
      12'h55C: dout <= 8'b00000000; // 1372 :   0 - 0x0
      12'h55D: dout <= 8'b00000000; // 1373 :   0 - 0x0
      12'h55E: dout <= 8'b00000000; // 1374 :   0 - 0x0
      12'h55F: dout <= 8'b00000000; // 1375 :   0 - 0x0
      12'h560: dout <= 8'b00000000; // 1376 :   0 - 0x0 -- Sprite 0xac
      12'h561: dout <= 8'b00000110; // 1377 :   6 - 0x6
      12'h562: dout <= 8'b00000110; // 1378 :   6 - 0x6
      12'h563: dout <= 8'b00000110; // 1379 :   6 - 0x6
      12'h564: dout <= 8'b00000110; // 1380 :   6 - 0x6
      12'h565: dout <= 8'b00000110; // 1381 :   6 - 0x6
      12'h566: dout <= 8'b00000110; // 1382 :   6 - 0x6
      12'h567: dout <= 8'b00000110; // 1383 :   6 - 0x6
      12'h568: dout <= 8'b00000110; // 1384 :   6 - 0x6 -- Sprite 0xad
      12'h569: dout <= 8'b00000110; // 1385 :   6 - 0x6
      12'h56A: dout <= 8'b00000110; // 1386 :   6 - 0x6
      12'h56B: dout <= 8'b00000110; // 1387 :   6 - 0x6
      12'h56C: dout <= 8'b00000110; // 1388 :   6 - 0x6
      12'h56D: dout <= 8'b00000110; // 1389 :   6 - 0x6
      12'h56E: dout <= 8'b00000110; // 1390 :   6 - 0x6
      12'h56F: dout <= 8'b00000000; // 1391 :   0 - 0x0
      12'h570: dout <= 8'b00000000; // 1392 :   0 - 0x0 -- Sprite 0xae
      12'h571: dout <= 8'b00000001; // 1393 :   1 - 0x1
      12'h572: dout <= 8'b00000011; // 1394 :   3 - 0x3
      12'h573: dout <= 8'b00000010; // 1395 :   2 - 0x2
      12'h574: dout <= 8'b00000010; // 1396 :   2 - 0x2
      12'h575: dout <= 8'b00000000; // 1397 :   0 - 0x0
      12'h576: dout <= 8'b00000011; // 1398 :   3 - 0x3
      12'h577: dout <= 8'b00000010; // 1399 :   2 - 0x2
      12'h578: dout <= 8'b00000001; // 1400 :   1 - 0x1 -- Sprite 0xaf
      12'h579: dout <= 8'b00000011; // 1401 :   3 - 0x3
      12'h57A: dout <= 8'b00000101; // 1402 :   5 - 0x5
      12'h57B: dout <= 8'b00000100; // 1403 :   4 - 0x4
      12'h57C: dout <= 8'b00000101; // 1404 :   5 - 0x5
      12'h57D: dout <= 8'b00001101; // 1405 :  13 - 0xd
      12'h57E: dout <= 8'b00001100; // 1406 :  12 - 0xc
      12'h57F: dout <= 8'b00000001; // 1407 :   1 - 0x1
      12'h580: dout <= 8'b00000000; // 1408 :   0 - 0x0 -- Sprite 0xb0
      12'h581: dout <= 8'b00000000; // 1409 :   0 - 0x0
      12'h582: dout <= 8'b01000000; // 1410 :  64 - 0x40
      12'h583: dout <= 8'b11110000; // 1411 : 240 - 0xf0
      12'h584: dout <= 8'b11101000; // 1412 : 232 - 0xe8
      12'h585: dout <= 8'b10010000; // 1413 : 144 - 0x90
      12'h586: dout <= 8'b01010000; // 1414 :  80 - 0x50
      12'h587: dout <= 8'b11010000; // 1415 : 208 - 0xd0
      12'h588: dout <= 8'b11111000; // 1416 : 248 - 0xf8 -- Sprite 0xb1
      12'h589: dout <= 8'b11000000; // 1417 : 192 - 0xc0
      12'h58A: dout <= 8'b11100000; // 1418 : 224 - 0xe0
      12'h58B: dout <= 8'b01000000; // 1419 :  64 - 0x40
      12'h58C: dout <= 8'b10000000; // 1420 : 128 - 0x80
      12'h58D: dout <= 8'b11000000; // 1421 : 192 - 0xc0
      12'h58E: dout <= 8'b11100000; // 1422 : 224 - 0xe0
      12'h58F: dout <= 8'b01110000; // 1423 : 112 - 0x70
      12'h590: dout <= 8'b00000001; // 1424 :   1 - 0x1 -- Sprite 0xb2
      12'h591: dout <= 8'b00001101; // 1425 :  13 - 0xd
      12'h592: dout <= 8'b00001101; // 1426 :  13 - 0xd
      12'h593: dout <= 8'b00000011; // 1427 :   3 - 0x3
      12'h594: dout <= 8'b00000011; // 1428 :   3 - 0x3
      12'h595: dout <= 8'b00000111; // 1429 :   7 - 0x7
      12'h596: dout <= 8'b00000111; // 1430 :   7 - 0x7
      12'h597: dout <= 8'b00000000; // 1431 :   0 - 0x0
      12'h598: dout <= 8'b00111111; // 1432 :  63 - 0x3f -- Sprite 0xb3
      12'h599: dout <= 8'b00111111; // 1433 :  63 - 0x3f
      12'h59A: dout <= 8'b00111111; // 1434 :  63 - 0x3f
      12'h59B: dout <= 8'b00111111; // 1435 :  63 - 0x3f
      12'h59C: dout <= 8'b00111111; // 1436 :  63 - 0x3f
      12'h59D: dout <= 8'b00111111; // 1437 :  63 - 0x3f
      12'h59E: dout <= 8'b00110101; // 1438 :  53 - 0x35
      12'h59F: dout <= 8'b00000000; // 1439 :   0 - 0x0
      12'h5A0: dout <= 8'b10110000; // 1440 : 176 - 0xb0 -- Sprite 0xb4
      12'h5A1: dout <= 8'b11000000; // 1441 : 192 - 0xc0
      12'h5A2: dout <= 8'b11100000; // 1442 : 224 - 0xe0
      12'h5A3: dout <= 8'b11100000; // 1443 : 224 - 0xe0
      12'h5A4: dout <= 8'b11110000; // 1444 : 240 - 0xf0
      12'h5A5: dout <= 8'b11110000; // 1445 : 240 - 0xf0
      12'h5A6: dout <= 8'b11110000; // 1446 : 240 - 0xf0
      12'h5A7: dout <= 8'b00000000; // 1447 :   0 - 0x0
      12'h5A8: dout <= 8'b11111100; // 1448 : 252 - 0xfc -- Sprite 0xb5
      12'h5A9: dout <= 8'b11111000; // 1449 : 248 - 0xf8
      12'h5AA: dout <= 8'b11111100; // 1450 : 252 - 0xfc
      12'h5AB: dout <= 8'b11111000; // 1451 : 248 - 0xf8
      12'h5AC: dout <= 8'b11111100; // 1452 : 252 - 0xfc
      12'h5AD: dout <= 8'b11111000; // 1453 : 248 - 0xf8
      12'h5AE: dout <= 8'b01010100; // 1454 :  84 - 0x54
      12'h5AF: dout <= 8'b00000000; // 1455 :   0 - 0x0
      12'h5B0: dout <= 8'b00000000; // 1456 :   0 - 0x0 -- Sprite 0xb6
      12'h5B1: dout <= 8'b01111111; // 1457 : 127 - 0x7f
      12'h5B2: dout <= 8'b01111111; // 1458 : 127 - 0x7f
      12'h5B3: dout <= 8'b01111111; // 1459 : 127 - 0x7f
      12'h5B4: dout <= 8'b01111111; // 1460 : 127 - 0x7f
      12'h5B5: dout <= 8'b01111111; // 1461 : 127 - 0x7f
      12'h5B6: dout <= 8'b01101010; // 1462 : 106 - 0x6a
      12'h5B7: dout <= 8'b00000000; // 1463 :   0 - 0x0
      12'h5B8: dout <= 8'b00000000; // 1464 :   0 - 0x0 -- Sprite 0xb7
      12'h5B9: dout <= 8'b01111011; // 1465 : 123 - 0x7b
      12'h5BA: dout <= 8'b01110011; // 1466 : 115 - 0x73
      12'h5BB: dout <= 8'b01111011; // 1467 : 123 - 0x7b
      12'h5BC: dout <= 8'b01110011; // 1468 : 115 - 0x73
      12'h5BD: dout <= 8'b01111011; // 1469 : 123 - 0x7b
      12'h5BE: dout <= 8'b01010011; // 1470 :  83 - 0x53
      12'h5BF: dout <= 8'b00000000; // 1471 :   0 - 0x0
      12'h5C0: dout <= 8'b00000000; // 1472 :   0 - 0x0 -- Sprite 0xb8
      12'h5C1: dout <= 8'b11011110; // 1473 : 222 - 0xde
      12'h5C2: dout <= 8'b10011110; // 1474 : 158 - 0x9e
      12'h5C3: dout <= 8'b11011100; // 1475 : 220 - 0xdc
      12'h5C4: dout <= 8'b10011110; // 1476 : 158 - 0x9e
      12'h5C5: dout <= 8'b11011100; // 1477 : 220 - 0xdc
      12'h5C6: dout <= 8'b10011010; // 1478 : 154 - 0x9a
      12'h5C7: dout <= 8'b00000000; // 1479 :   0 - 0x0
      12'h5C8: dout <= 8'b00000000; // 1480 :   0 - 0x0 -- Sprite 0xb9
      12'h5C9: dout <= 8'b11111110; // 1481 : 254 - 0xfe
      12'h5CA: dout <= 8'b11111100; // 1482 : 252 - 0xfc
      12'h5CB: dout <= 8'b11111110; // 1483 : 254 - 0xfe
      12'h5CC: dout <= 8'b11111100; // 1484 : 252 - 0xfc
      12'h5CD: dout <= 8'b11111110; // 1485 : 254 - 0xfe
      12'h5CE: dout <= 8'b01010100; // 1486 :  84 - 0x54
      12'h5CF: dout <= 8'b00000000; // 1487 :   0 - 0x0
      12'h5D0: dout <= 8'b00000000; // 1488 :   0 - 0x0 -- Sprite 0xba
      12'h5D1: dout <= 8'b01111111; // 1489 : 127 - 0x7f
      12'h5D2: dout <= 8'b01111111; // 1490 : 127 - 0x7f
      12'h5D3: dout <= 8'b00000000; // 1491 :   0 - 0x0
      12'h5D4: dout <= 8'b01111111; // 1492 : 127 - 0x7f
      12'h5D5: dout <= 8'b01111111; // 1493 : 127 - 0x7f
      12'h5D6: dout <= 8'b01101010; // 1494 : 106 - 0x6a
      12'h5D7: dout <= 8'b00000000; // 1495 :   0 - 0x0
      12'h5D8: dout <= 8'b00000000; // 1496 :   0 - 0x0 -- Sprite 0xbb
      12'h5D9: dout <= 8'b00000000; // 1497 :   0 - 0x0
      12'h5DA: dout <= 8'b00000000; // 1498 :   0 - 0x0
      12'h5DB: dout <= 8'b00000000; // 1499 :   0 - 0x0
      12'h5DC: dout <= 8'b00000000; // 1500 :   0 - 0x0
      12'h5DD: dout <= 8'b00000000; // 1501 :   0 - 0x0
      12'h5DE: dout <= 8'b00000000; // 1502 :   0 - 0x0
      12'h5DF: dout <= 8'b00000000; // 1503 :   0 - 0x0
      12'h5E0: dout <= 8'b00000000; // 1504 :   0 - 0x0 -- Sprite 0xbc
      12'h5E1: dout <= 8'b11111110; // 1505 : 254 - 0xfe
      12'h5E2: dout <= 8'b11111110; // 1506 : 254 - 0xfe
      12'h5E3: dout <= 8'b00000000; // 1507 :   0 - 0x0
      12'h5E4: dout <= 8'b10011110; // 1508 : 158 - 0x9e
      12'h5E5: dout <= 8'b11011100; // 1509 : 220 - 0xdc
      12'h5E6: dout <= 8'b10011010; // 1510 : 154 - 0x9a
      12'h5E7: dout <= 8'b00000000; // 1511 :   0 - 0x0
      12'h5E8: dout <= 8'b00000000; // 1512 :   0 - 0x0 -- Sprite 0xbd
      12'h5E9: dout <= 8'b00000000; // 1513 :   0 - 0x0
      12'h5EA: dout <= 8'b00000000; // 1514 :   0 - 0x0
      12'h5EB: dout <= 8'b00000000; // 1515 :   0 - 0x0
      12'h5EC: dout <= 8'b00000000; // 1516 :   0 - 0x0
      12'h5ED: dout <= 8'b00000000; // 1517 :   0 - 0x0
      12'h5EE: dout <= 8'b00000000; // 1518 :   0 - 0x0
      12'h5EF: dout <= 8'b00000000; // 1519 :   0 - 0x0
      12'h5F0: dout <= 8'b00000000; // 1520 :   0 - 0x0 -- Sprite 0xbe
      12'h5F1: dout <= 8'b00000000; // 1521 :   0 - 0x0
      12'h5F2: dout <= 8'b00000000; // 1522 :   0 - 0x0
      12'h5F3: dout <= 8'b00000000; // 1523 :   0 - 0x0
      12'h5F4: dout <= 8'b00000000; // 1524 :   0 - 0x0
      12'h5F5: dout <= 8'b00000000; // 1525 :   0 - 0x0
      12'h5F6: dout <= 8'b00000000; // 1526 :   0 - 0x0
      12'h5F7: dout <= 8'b00000000; // 1527 :   0 - 0x0
      12'h5F8: dout <= 8'b00000000; // 1528 :   0 - 0x0 -- Sprite 0xbf
      12'h5F9: dout <= 8'b00000000; // 1529 :   0 - 0x0
      12'h5FA: dout <= 8'b00000000; // 1530 :   0 - 0x0
      12'h5FB: dout <= 8'b00000000; // 1531 :   0 - 0x0
      12'h5FC: dout <= 8'b00000000; // 1532 :   0 - 0x0
      12'h5FD: dout <= 8'b00000000; // 1533 :   0 - 0x0
      12'h5FE: dout <= 8'b00000000; // 1534 :   0 - 0x0
      12'h5FF: dout <= 8'b00000000; // 1535 :   0 - 0x0
      12'h600: dout <= 8'b00000000; // 1536 :   0 - 0x0 -- Sprite 0xc0
      12'h601: dout <= 8'b00000000; // 1537 :   0 - 0x0
      12'h602: dout <= 8'b00000000; // 1538 :   0 - 0x0
      12'h603: dout <= 8'b00000000; // 1539 :   0 - 0x0
      12'h604: dout <= 8'b00000000; // 1540 :   0 - 0x0
      12'h605: dout <= 8'b00000000; // 1541 :   0 - 0x0
      12'h606: dout <= 8'b00000000; // 1542 :   0 - 0x0
      12'h607: dout <= 8'b00000000; // 1543 :   0 - 0x0
      12'h608: dout <= 8'b00000000; // 1544 :   0 - 0x0 -- Sprite 0xc1
      12'h609: dout <= 8'b00000000; // 1545 :   0 - 0x0
      12'h60A: dout <= 8'b00000000; // 1546 :   0 - 0x0
      12'h60B: dout <= 8'b00000000; // 1547 :   0 - 0x0
      12'h60C: dout <= 8'b00000000; // 1548 :   0 - 0x0
      12'h60D: dout <= 8'b00000000; // 1549 :   0 - 0x0
      12'h60E: dout <= 8'b00000000; // 1550 :   0 - 0x0
      12'h60F: dout <= 8'b00000000; // 1551 :   0 - 0x0
      12'h610: dout <= 8'b00000000; // 1552 :   0 - 0x0 -- Sprite 0xc2
      12'h611: dout <= 8'b00000000; // 1553 :   0 - 0x0
      12'h612: dout <= 8'b00000000; // 1554 :   0 - 0x0
      12'h613: dout <= 8'b00000000; // 1555 :   0 - 0x0
      12'h614: dout <= 8'b00000000; // 1556 :   0 - 0x0
      12'h615: dout <= 8'b00000000; // 1557 :   0 - 0x0
      12'h616: dout <= 8'b00000000; // 1558 :   0 - 0x0
      12'h617: dout <= 8'b00000000; // 1559 :   0 - 0x0
      12'h618: dout <= 8'b00000000; // 1560 :   0 - 0x0 -- Sprite 0xc3
      12'h619: dout <= 8'b00000000; // 1561 :   0 - 0x0
      12'h61A: dout <= 8'b00000000; // 1562 :   0 - 0x0
      12'h61B: dout <= 8'b00000000; // 1563 :   0 - 0x0
      12'h61C: dout <= 8'b00000000; // 1564 :   0 - 0x0
      12'h61D: dout <= 8'b00000000; // 1565 :   0 - 0x0
      12'h61E: dout <= 8'b00000000; // 1566 :   0 - 0x0
      12'h61F: dout <= 8'b00000000; // 1567 :   0 - 0x0
      12'h620: dout <= 8'b00000000; // 1568 :   0 - 0x0 -- Sprite 0xc4
      12'h621: dout <= 8'b00000000; // 1569 :   0 - 0x0
      12'h622: dout <= 8'b00000000; // 1570 :   0 - 0x0
      12'h623: dout <= 8'b00000000; // 1571 :   0 - 0x0
      12'h624: dout <= 8'b00000000; // 1572 :   0 - 0x0
      12'h625: dout <= 8'b00000000; // 1573 :   0 - 0x0
      12'h626: dout <= 8'b00000000; // 1574 :   0 - 0x0
      12'h627: dout <= 8'b00000000; // 1575 :   0 - 0x0
      12'h628: dout <= 8'b00000000; // 1576 :   0 - 0x0 -- Sprite 0xc5
      12'h629: dout <= 8'b00000000; // 1577 :   0 - 0x0
      12'h62A: dout <= 8'b00000000; // 1578 :   0 - 0x0
      12'h62B: dout <= 8'b00000001; // 1579 :   1 - 0x1
      12'h62C: dout <= 8'b00000111; // 1580 :   7 - 0x7
      12'h62D: dout <= 8'b00001111; // 1581 :  15 - 0xf
      12'h62E: dout <= 8'b00001111; // 1582 :  15 - 0xf
      12'h62F: dout <= 8'b00011111; // 1583 :  31 - 0x1f
      12'h630: dout <= 8'b00000000; // 1584 :   0 - 0x0 -- Sprite 0xc6
      12'h631: dout <= 8'b00011111; // 1585 :  31 - 0x1f
      12'h632: dout <= 8'b01111111; // 1586 : 127 - 0x7f
      12'h633: dout <= 8'b11111111; // 1587 : 255 - 0xff
      12'h634: dout <= 8'b11111111; // 1588 : 255 - 0xff
      12'h635: dout <= 8'b11111111; // 1589 : 255 - 0xff
      12'h636: dout <= 8'b11111111; // 1590 : 255 - 0xff
      12'h637: dout <= 8'b11111111; // 1591 : 255 - 0xff
      12'h638: dout <= 8'b00011111; // 1592 :  31 - 0x1f -- Sprite 0xc7
      12'h639: dout <= 8'b00111111; // 1593 :  63 - 0x3f
      12'h63A: dout <= 8'b00111111; // 1594 :  63 - 0x3f
      12'h63B: dout <= 8'b01111111; // 1595 : 127 - 0x7f
      12'h63C: dout <= 8'b01111111; // 1596 : 127 - 0x7f
      12'h63D: dout <= 8'b01111111; // 1597 : 127 - 0x7f
      12'h63E: dout <= 8'b01111111; // 1598 : 127 - 0x7f
      12'h63F: dout <= 8'b01111111; // 1599 : 127 - 0x7f
      12'h640: dout <= 8'b00000000; // 1600 :   0 - 0x0 -- Sprite 0xc8
      12'h641: dout <= 8'b11111111; // 1601 : 255 - 0xff
      12'h642: dout <= 8'b11111111; // 1602 : 255 - 0xff
      12'h643: dout <= 8'b11111111; // 1603 : 255 - 0xff
      12'h644: dout <= 8'b11111111; // 1604 : 255 - 0xff
      12'h645: dout <= 8'b11111111; // 1605 : 255 - 0xff
      12'h646: dout <= 8'b11111111; // 1606 : 255 - 0xff
      12'h647: dout <= 8'b11111111; // 1607 : 255 - 0xff
      12'h648: dout <= 8'b11101000; // 1608 : 232 - 0xe8 -- Sprite 0xc9
      12'h649: dout <= 8'b11010100; // 1609 : 212 - 0xd4
      12'h64A: dout <= 8'b11101000; // 1610 : 232 - 0xe8
      12'h64B: dout <= 8'b11010100; // 1611 : 212 - 0xd4
      12'h64C: dout <= 8'b11101010; // 1612 : 234 - 0xea
      12'h64D: dout <= 8'b11010100; // 1613 : 212 - 0xd4
      12'h64E: dout <= 8'b11101010; // 1614 : 234 - 0xea
      12'h64F: dout <= 8'b11010100; // 1615 : 212 - 0xd4
      12'h650: dout <= 8'b00000000; // 1616 :   0 - 0x0 -- Sprite 0xca
      12'h651: dout <= 8'b00000000; // 1617 :   0 - 0x0
      12'h652: dout <= 8'b00000000; // 1618 :   0 - 0x0
      12'h653: dout <= 8'b00000000; // 1619 :   0 - 0x0
      12'h654: dout <= 8'b00000000; // 1620 :   0 - 0x0
      12'h655: dout <= 8'b00000000; // 1621 :   0 - 0x0
      12'h656: dout <= 8'b00000000; // 1622 :   0 - 0x0
      12'h657: dout <= 8'b00000000; // 1623 :   0 - 0x0
      12'h658: dout <= 8'b00000000; // 1624 :   0 - 0x0 -- Sprite 0xcb
      12'h659: dout <= 8'b00000000; // 1625 :   0 - 0x0
      12'h65A: dout <= 8'b00000000; // 1626 :   0 - 0x0
      12'h65B: dout <= 8'b00000000; // 1627 :   0 - 0x0
      12'h65C: dout <= 8'b00000000; // 1628 :   0 - 0x0
      12'h65D: dout <= 8'b00000000; // 1629 :   0 - 0x0
      12'h65E: dout <= 8'b00000000; // 1630 :   0 - 0x0
      12'h65F: dout <= 8'b00000000; // 1631 :   0 - 0x0
      12'h660: dout <= 8'b00000000; // 1632 :   0 - 0x0 -- Sprite 0xcc
      12'h661: dout <= 8'b00000000; // 1633 :   0 - 0x0
      12'h662: dout <= 8'b00000000; // 1634 :   0 - 0x0
      12'h663: dout <= 8'b00000000; // 1635 :   0 - 0x0
      12'h664: dout <= 8'b00000101; // 1636 :   5 - 0x5
      12'h665: dout <= 8'b00000010; // 1637 :   2 - 0x2
      12'h666: dout <= 8'b00000001; // 1638 :   1 - 0x1
      12'h667: dout <= 8'b00000000; // 1639 :   0 - 0x0
      12'h668: dout <= 8'b00000000; // 1640 :   0 - 0x0 -- Sprite 0xcd
      12'h669: dout <= 8'b00000000; // 1641 :   0 - 0x0
      12'h66A: dout <= 8'b00000000; // 1642 :   0 - 0x0
      12'h66B: dout <= 8'b10000000; // 1643 : 128 - 0x80
      12'h66C: dout <= 8'b01010000; // 1644 :  80 - 0x50
      12'h66D: dout <= 8'b10100000; // 1645 : 160 - 0xa0
      12'h66E: dout <= 8'b01000000; // 1646 :  64 - 0x40
      12'h66F: dout <= 8'b10000000; // 1647 : 128 - 0x80
      12'h670: dout <= 8'b00000000; // 1648 :   0 - 0x0 -- Sprite 0xce
      12'h671: dout <= 8'b00000000; // 1649 :   0 - 0x0
      12'h672: dout <= 8'b00000000; // 1650 :   0 - 0x0
      12'h673: dout <= 8'b00000000; // 1651 :   0 - 0x0
      12'h674: dout <= 8'b00110000; // 1652 :  48 - 0x30
      12'h675: dout <= 8'b01111111; // 1653 : 127 - 0x7f
      12'h676: dout <= 8'b00110000; // 1654 :  48 - 0x30
      12'h677: dout <= 8'b00110000; // 1655 :  48 - 0x30
      12'h678: dout <= 8'b00000000; // 1656 :   0 - 0x0 -- Sprite 0xcf
      12'h679: dout <= 8'b00000000; // 1657 :   0 - 0x0
      12'h67A: dout <= 8'b00000000; // 1658 :   0 - 0x0
      12'h67B: dout <= 8'b00000000; // 1659 :   0 - 0x0
      12'h67C: dout <= 8'b00001100; // 1660 :  12 - 0xc
      12'h67D: dout <= 8'b11111110; // 1661 : 254 - 0xfe
      12'h67E: dout <= 8'b00001100; // 1662 :  12 - 0xc
      12'h67F: dout <= 8'b00001100; // 1663 :  12 - 0xc
      12'h680: dout <= 8'b00000000; // 1664 :   0 - 0x0 -- Sprite 0xd0
      12'h681: dout <= 8'b00000000; // 1665 :   0 - 0x0
      12'h682: dout <= 8'b00000000; // 1666 :   0 - 0x0
      12'h683: dout <= 8'b00000000; // 1667 :   0 - 0x0
      12'h684: dout <= 8'b00000000; // 1668 :   0 - 0x0
      12'h685: dout <= 8'b00000000; // 1669 :   0 - 0x0
      12'h686: dout <= 8'b00000000; // 1670 :   0 - 0x0
      12'h687: dout <= 8'b00000000; // 1671 :   0 - 0x0
      12'h688: dout <= 8'b00000000; // 1672 :   0 - 0x0 -- Sprite 0xd1
      12'h689: dout <= 8'b00000000; // 1673 :   0 - 0x0
      12'h68A: dout <= 8'b00000000; // 1674 :   0 - 0x0
      12'h68B: dout <= 8'b00000000; // 1675 :   0 - 0x0
      12'h68C: dout <= 8'b00000000; // 1676 :   0 - 0x0
      12'h68D: dout <= 8'b00000000; // 1677 :   0 - 0x0
      12'h68E: dout <= 8'b00000000; // 1678 :   0 - 0x0
      12'h68F: dout <= 8'b00000000; // 1679 :   0 - 0x0
      12'h690: dout <= 8'b00000111; // 1680 :   7 - 0x7 -- Sprite 0xd2
      12'h691: dout <= 8'b00000111; // 1681 :   7 - 0x7
      12'h692: dout <= 8'b00000111; // 1682 :   7 - 0x7
      12'h693: dout <= 8'b00000111; // 1683 :   7 - 0x7
      12'h694: dout <= 8'b00000111; // 1684 :   7 - 0x7
      12'h695: dout <= 8'b00000111; // 1685 :   7 - 0x7
      12'h696: dout <= 8'b00000111; // 1686 :   7 - 0x7
      12'h697: dout <= 8'b00000111; // 1687 :   7 - 0x7
      12'h698: dout <= 8'b11100000; // 1688 : 224 - 0xe0 -- Sprite 0xd3
      12'h699: dout <= 8'b11100000; // 1689 : 224 - 0xe0
      12'h69A: dout <= 8'b11000000; // 1690 : 192 - 0xc0
      12'h69B: dout <= 8'b11100000; // 1691 : 224 - 0xe0
      12'h69C: dout <= 8'b10100000; // 1692 : 160 - 0xa0
      12'h69D: dout <= 8'b11100000; // 1693 : 224 - 0xe0
      12'h69E: dout <= 8'b11000000; // 1694 : 192 - 0xc0
      12'h69F: dout <= 8'b11100000; // 1695 : 224 - 0xe0
      12'h6A0: dout <= 8'b00000000; // 1696 :   0 - 0x0 -- Sprite 0xd4
      12'h6A1: dout <= 8'b00000000; // 1697 :   0 - 0x0
      12'h6A2: dout <= 8'b00000000; // 1698 :   0 - 0x0
      12'h6A3: dout <= 8'b00000000; // 1699 :   0 - 0x0
      12'h6A4: dout <= 8'b00000000; // 1700 :   0 - 0x0
      12'h6A5: dout <= 8'b00000000; // 1701 :   0 - 0x0
      12'h6A6: dout <= 8'b00000000; // 1702 :   0 - 0x0
      12'h6A7: dout <= 8'b00000000; // 1703 :   0 - 0x0
      12'h6A8: dout <= 8'b00000000; // 1704 :   0 - 0x0 -- Sprite 0xd5
      12'h6A9: dout <= 8'b11111000; // 1705 : 248 - 0xf8
      12'h6AA: dout <= 8'b11111110; // 1706 : 254 - 0xfe
      12'h6AB: dout <= 8'b11111111; // 1707 : 255 - 0xff
      12'h6AC: dout <= 8'b11111111; // 1708 : 255 - 0xff
      12'h6AD: dout <= 8'b11111111; // 1709 : 255 - 0xff
      12'h6AE: dout <= 8'b11111111; // 1710 : 255 - 0xff
      12'h6AF: dout <= 8'b11111111; // 1711 : 255 - 0xff
      12'h6B0: dout <= 8'b00000000; // 1712 :   0 - 0x0 -- Sprite 0xd6
      12'h6B1: dout <= 8'b00000000; // 1713 :   0 - 0x0
      12'h6B2: dout <= 8'b00000000; // 1714 :   0 - 0x0
      12'h6B3: dout <= 8'b10000000; // 1715 : 128 - 0x80
      12'h6B4: dout <= 8'b10100000; // 1716 : 160 - 0xa0
      12'h6B5: dout <= 8'b01010000; // 1717 :  80 - 0x50
      12'h6B6: dout <= 8'b10100000; // 1718 : 160 - 0xa0
      12'h6B7: dout <= 8'b11010000; // 1719 : 208 - 0xd0
      12'h6B8: dout <= 8'b01111111; // 1720 : 127 - 0x7f -- Sprite 0xd7
      12'h6B9: dout <= 8'b01111111; // 1721 : 127 - 0x7f
      12'h6BA: dout <= 8'b01111111; // 1722 : 127 - 0x7f
      12'h6BB: dout <= 8'b00111111; // 1723 :  63 - 0x3f
      12'h6BC: dout <= 8'b00111111; // 1724 :  63 - 0x3f
      12'h6BD: dout <= 8'b00001111; // 1725 :  15 - 0xf
      12'h6BE: dout <= 8'b00000111; // 1726 :   7 - 0x7
      12'h6BF: dout <= 8'b00000000; // 1727 :   0 - 0x0
      12'h6C0: dout <= 8'b11111111; // 1728 : 255 - 0xff -- Sprite 0xd8
      12'h6C1: dout <= 8'b11111111; // 1729 : 255 - 0xff
      12'h6C2: dout <= 8'b11111111; // 1730 : 255 - 0xff
      12'h6C3: dout <= 8'b11111111; // 1731 : 255 - 0xff
      12'h6C4: dout <= 8'b11111111; // 1732 : 255 - 0xff
      12'h6C5: dout <= 8'b11111111; // 1733 : 255 - 0xff
      12'h6C6: dout <= 8'b11111111; // 1734 : 255 - 0xff
      12'h6C7: dout <= 8'b00000000; // 1735 :   0 - 0x0
      12'h6C8: dout <= 8'b11101010; // 1736 : 234 - 0xea -- Sprite 0xd9
      12'h6C9: dout <= 8'b11010100; // 1737 : 212 - 0xd4
      12'h6CA: dout <= 8'b11101010; // 1738 : 234 - 0xea
      12'h6CB: dout <= 8'b11010100; // 1739 : 212 - 0xd4
      12'h6CC: dout <= 8'b10101000; // 1740 : 168 - 0xa8
      12'h6CD: dout <= 8'b01010000; // 1741 :  80 - 0x50
      12'h6CE: dout <= 8'b10100000; // 1742 : 160 - 0xa0
      12'h6CF: dout <= 8'b00000000; // 1743 :   0 - 0x0
      12'h6D0: dout <= 8'b00000000; // 1744 :   0 - 0x0 -- Sprite 0xda
      12'h6D1: dout <= 8'b00000000; // 1745 :   0 - 0x0
      12'h6D2: dout <= 8'b00001100; // 1746 :  12 - 0xc
      12'h6D3: dout <= 8'b00000000; // 1747 :   0 - 0x0
      12'h6D4: dout <= 8'b00000000; // 1748 :   0 - 0x0
      12'h6D5: dout <= 8'b00000000; // 1749 :   0 - 0x0
      12'h6D6: dout <= 8'b00000000; // 1750 :   0 - 0x0
      12'h6D7: dout <= 8'b00000000; // 1751 :   0 - 0x0
      12'h6D8: dout <= 8'b00000000; // 1752 :   0 - 0x0 -- Sprite 0xdb
      12'h6D9: dout <= 8'b10000000; // 1753 : 128 - 0x80
      12'h6DA: dout <= 8'b10000000; // 1754 : 128 - 0x80
      12'h6DB: dout <= 8'b10000000; // 1755 : 128 - 0x80
      12'h6DC: dout <= 8'b10011000; // 1756 : 152 - 0x98
      12'h6DD: dout <= 8'b10000000; // 1757 : 128 - 0x80
      12'h6DE: dout <= 8'b10000000; // 1758 : 128 - 0x80
      12'h6DF: dout <= 8'b10000000; // 1759 : 128 - 0x80
      12'h6E0: dout <= 8'b00000000; // 1760 :   0 - 0x0 -- Sprite 0xdc
      12'h6E1: dout <= 8'b00000000; // 1761 :   0 - 0x0
      12'h6E2: dout <= 8'b00000000; // 1762 :   0 - 0x0
      12'h6E3: dout <= 8'b00000000; // 1763 :   0 - 0x0
      12'h6E4: dout <= 8'b00000010; // 1764 :   2 - 0x2
      12'h6E5: dout <= 8'b00000011; // 1765 :   3 - 0x3
      12'h6E6: dout <= 8'b00000011; // 1766 :   3 - 0x3
      12'h6E7: dout <= 8'b00000001; // 1767 :   1 - 0x1
      12'h6E8: dout <= 8'b00000000; // 1768 :   0 - 0x0 -- Sprite 0xdd
      12'h6E9: dout <= 8'b00000000; // 1769 :   0 - 0x0
      12'h6EA: dout <= 8'b00000000; // 1770 :   0 - 0x0
      12'h6EB: dout <= 8'b00000000; // 1771 :   0 - 0x0
      12'h6EC: dout <= 8'b10100000; // 1772 : 160 - 0xa0
      12'h6ED: dout <= 8'b11100000; // 1773 : 224 - 0xe0
      12'h6EE: dout <= 8'b11100000; // 1774 : 224 - 0xe0
      12'h6EF: dout <= 8'b11000000; // 1775 : 192 - 0xc0
      12'h6F0: dout <= 8'b00110000; // 1776 :  48 - 0x30 -- Sprite 0xde
      12'h6F1: dout <= 8'b01111111; // 1777 : 127 - 0x7f
      12'h6F2: dout <= 8'b00110000; // 1778 :  48 - 0x30
      12'h6F3: dout <= 8'b00110000; // 1779 :  48 - 0x30
      12'h6F4: dout <= 8'b00110000; // 1780 :  48 - 0x30
      12'h6F5: dout <= 8'b00110000; // 1781 :  48 - 0x30
      12'h6F6: dout <= 8'b00110000; // 1782 :  48 - 0x30
      12'h6F7: dout <= 8'b00110000; // 1783 :  48 - 0x30
      12'h6F8: dout <= 8'b00001100; // 1784 :  12 - 0xc -- Sprite 0xdf
      12'h6F9: dout <= 8'b11111110; // 1785 : 254 - 0xfe
      12'h6FA: dout <= 8'b00001100; // 1786 :  12 - 0xc
      12'h6FB: dout <= 8'b00001100; // 1787 :  12 - 0xc
      12'h6FC: dout <= 8'b00001100; // 1788 :  12 - 0xc
      12'h6FD: dout <= 8'b00001100; // 1789 :  12 - 0xc
      12'h6FE: dout <= 8'b00001100; // 1790 :  12 - 0xc
      12'h6FF: dout <= 8'b00001100; // 1791 :  12 - 0xc
      12'h700: dout <= 8'b00000000; // 1792 :   0 - 0x0 -- Sprite 0xe0
      12'h701: dout <= 8'b00000000; // 1793 :   0 - 0x0
      12'h702: dout <= 8'b00000000; // 1794 :   0 - 0x0
      12'h703: dout <= 8'b00000000; // 1795 :   0 - 0x0
      12'h704: dout <= 8'b00000000; // 1796 :   0 - 0x0
      12'h705: dout <= 8'b00000000; // 1797 :   0 - 0x0
      12'h706: dout <= 8'b00000000; // 1798 :   0 - 0x0
      12'h707: dout <= 8'b00000000; // 1799 :   0 - 0x0
      12'h708: dout <= 8'b00000000; // 1800 :   0 - 0x0 -- Sprite 0xe1
      12'h709: dout <= 8'b00000000; // 1801 :   0 - 0x0
      12'h70A: dout <= 8'b00000000; // 1802 :   0 - 0x0
      12'h70B: dout <= 8'b00000000; // 1803 :   0 - 0x0
      12'h70C: dout <= 8'b00000000; // 1804 :   0 - 0x0
      12'h70D: dout <= 8'b00000000; // 1805 :   0 - 0x0
      12'h70E: dout <= 8'b00000000; // 1806 :   0 - 0x0
      12'h70F: dout <= 8'b00000000; // 1807 :   0 - 0x0
      12'h710: dout <= 8'b00000000; // 1808 :   0 - 0x0 -- Sprite 0xe2
      12'h711: dout <= 8'b00000000; // 1809 :   0 - 0x0
      12'h712: dout <= 8'b00000000; // 1810 :   0 - 0x0
      12'h713: dout <= 8'b00000000; // 1811 :   0 - 0x0
      12'h714: dout <= 8'b00000000; // 1812 :   0 - 0x0
      12'h715: dout <= 8'b00000000; // 1813 :   0 - 0x0
      12'h716: dout <= 8'b00000000; // 1814 :   0 - 0x0
      12'h717: dout <= 8'b00000000; // 1815 :   0 - 0x0
      12'h718: dout <= 8'b00000000; // 1816 :   0 - 0x0 -- Sprite 0xe3
      12'h719: dout <= 8'b00000000; // 1817 :   0 - 0x0
      12'h71A: dout <= 8'b00000000; // 1818 :   0 - 0x0
      12'h71B: dout <= 8'b00000000; // 1819 :   0 - 0x0
      12'h71C: dout <= 8'b00000000; // 1820 :   0 - 0x0
      12'h71D: dout <= 8'b00000000; // 1821 :   0 - 0x0
      12'h71E: dout <= 8'b00000000; // 1822 :   0 - 0x0
      12'h71F: dout <= 8'b00000000; // 1823 :   0 - 0x0
      12'h720: dout <= 8'b00000000; // 1824 :   0 - 0x0 -- Sprite 0xe4
      12'h721: dout <= 8'b00000000; // 1825 :   0 - 0x0
      12'h722: dout <= 8'b00000000; // 1826 :   0 - 0x0
      12'h723: dout <= 8'b00000000; // 1827 :   0 - 0x0
      12'h724: dout <= 8'b00000000; // 1828 :   0 - 0x0
      12'h725: dout <= 8'b00000000; // 1829 :   0 - 0x0
      12'h726: dout <= 8'b00000000; // 1830 :   0 - 0x0
      12'h727: dout <= 8'b00000000; // 1831 :   0 - 0x0
      12'h728: dout <= 8'b00000000; // 1832 :   0 - 0x0 -- Sprite 0xe5
      12'h729: dout <= 8'b00000000; // 1833 :   0 - 0x0
      12'h72A: dout <= 8'b00000000; // 1834 :   0 - 0x0
      12'h72B: dout <= 8'b00000000; // 1835 :   0 - 0x0
      12'h72C: dout <= 8'b00000000; // 1836 :   0 - 0x0
      12'h72D: dout <= 8'b00000000; // 1837 :   0 - 0x0
      12'h72E: dout <= 8'b00000000; // 1838 :   0 - 0x0
      12'h72F: dout <= 8'b00000000; // 1839 :   0 - 0x0
      12'h730: dout <= 8'b00000000; // 1840 :   0 - 0x0 -- Sprite 0xe6
      12'h731: dout <= 8'b00000000; // 1841 :   0 - 0x0
      12'h732: dout <= 8'b00000000; // 1842 :   0 - 0x0
      12'h733: dout <= 8'b00000000; // 1843 :   0 - 0x0
      12'h734: dout <= 8'b00000000; // 1844 :   0 - 0x0
      12'h735: dout <= 8'b00000000; // 1845 :   0 - 0x0
      12'h736: dout <= 8'b00000000; // 1846 :   0 - 0x0
      12'h737: dout <= 8'b00000000; // 1847 :   0 - 0x0
      12'h738: dout <= 8'b00000000; // 1848 :   0 - 0x0 -- Sprite 0xe7
      12'h739: dout <= 8'b00000000; // 1849 :   0 - 0x0
      12'h73A: dout <= 8'b00000000; // 1850 :   0 - 0x0
      12'h73B: dout <= 8'b00000000; // 1851 :   0 - 0x0
      12'h73C: dout <= 8'b00000000; // 1852 :   0 - 0x0
      12'h73D: dout <= 8'b00000000; // 1853 :   0 - 0x0
      12'h73E: dout <= 8'b00000000; // 1854 :   0 - 0x0
      12'h73F: dout <= 8'b00000000; // 1855 :   0 - 0x0
      12'h740: dout <= 8'b00000000; // 1856 :   0 - 0x0 -- Sprite 0xe8
      12'h741: dout <= 8'b00000000; // 1857 :   0 - 0x0
      12'h742: dout <= 8'b00000000; // 1858 :   0 - 0x0
      12'h743: dout <= 8'b00000000; // 1859 :   0 - 0x0
      12'h744: dout <= 8'b00000000; // 1860 :   0 - 0x0
      12'h745: dout <= 8'b00000000; // 1861 :   0 - 0x0
      12'h746: dout <= 8'b00000000; // 1862 :   0 - 0x0
      12'h747: dout <= 8'b00000000; // 1863 :   0 - 0x0
      12'h748: dout <= 8'b00000000; // 1864 :   0 - 0x0 -- Sprite 0xe9
      12'h749: dout <= 8'b00000000; // 1865 :   0 - 0x0
      12'h74A: dout <= 8'b00000000; // 1866 :   0 - 0x0
      12'h74B: dout <= 8'b00000000; // 1867 :   0 - 0x0
      12'h74C: dout <= 8'b00000000; // 1868 :   0 - 0x0
      12'h74D: dout <= 8'b00000000; // 1869 :   0 - 0x0
      12'h74E: dout <= 8'b00000000; // 1870 :   0 - 0x0
      12'h74F: dout <= 8'b00000000; // 1871 :   0 - 0x0
      12'h750: dout <= 8'b00000000; // 1872 :   0 - 0x0 -- Sprite 0xea
      12'h751: dout <= 8'b00000000; // 1873 :   0 - 0x0
      12'h752: dout <= 8'b00000000; // 1874 :   0 - 0x0
      12'h753: dout <= 8'b00000000; // 1875 :   0 - 0x0
      12'h754: dout <= 8'b00000000; // 1876 :   0 - 0x0
      12'h755: dout <= 8'b00000000; // 1877 :   0 - 0x0
      12'h756: dout <= 8'b00000000; // 1878 :   0 - 0x0
      12'h757: dout <= 8'b00000000; // 1879 :   0 - 0x0
      12'h758: dout <= 8'b00000000; // 1880 :   0 - 0x0 -- Sprite 0xeb
      12'h759: dout <= 8'b00000000; // 1881 :   0 - 0x0
      12'h75A: dout <= 8'b00000000; // 1882 :   0 - 0x0
      12'h75B: dout <= 8'b00000000; // 1883 :   0 - 0x0
      12'h75C: dout <= 8'b00000000; // 1884 :   0 - 0x0
      12'h75D: dout <= 8'b00000000; // 1885 :   0 - 0x0
      12'h75E: dout <= 8'b00000000; // 1886 :   0 - 0x0
      12'h75F: dout <= 8'b00000000; // 1887 :   0 - 0x0
      12'h760: dout <= 8'b00000000; // 1888 :   0 - 0x0 -- Sprite 0xec
      12'h761: dout <= 8'b00000000; // 1889 :   0 - 0x0
      12'h762: dout <= 8'b00000000; // 1890 :   0 - 0x0
      12'h763: dout <= 8'b00000000; // 1891 :   0 - 0x0
      12'h764: dout <= 8'b00000000; // 1892 :   0 - 0x0
      12'h765: dout <= 8'b00000000; // 1893 :   0 - 0x0
      12'h766: dout <= 8'b00000000; // 1894 :   0 - 0x0
      12'h767: dout <= 8'b00000000; // 1895 :   0 - 0x0
      12'h768: dout <= 8'b00000000; // 1896 :   0 - 0x0 -- Sprite 0xed
      12'h769: dout <= 8'b00000000; // 1897 :   0 - 0x0
      12'h76A: dout <= 8'b00000000; // 1898 :   0 - 0x0
      12'h76B: dout <= 8'b00000000; // 1899 :   0 - 0x0
      12'h76C: dout <= 8'b00000000; // 1900 :   0 - 0x0
      12'h76D: dout <= 8'b00000000; // 1901 :   0 - 0x0
      12'h76E: dout <= 8'b00000000; // 1902 :   0 - 0x0
      12'h76F: dout <= 8'b00000000; // 1903 :   0 - 0x0
      12'h770: dout <= 8'b00000000; // 1904 :   0 - 0x0 -- Sprite 0xee
      12'h771: dout <= 8'b00000000; // 1905 :   0 - 0x0
      12'h772: dout <= 8'b00000000; // 1906 :   0 - 0x0
      12'h773: dout <= 8'b00000000; // 1907 :   0 - 0x0
      12'h774: dout <= 8'b00000000; // 1908 :   0 - 0x0
      12'h775: dout <= 8'b00000000; // 1909 :   0 - 0x0
      12'h776: dout <= 8'b00000000; // 1910 :   0 - 0x0
      12'h777: dout <= 8'b00000000; // 1911 :   0 - 0x0
      12'h778: dout <= 8'b00000000; // 1912 :   0 - 0x0 -- Sprite 0xef
      12'h779: dout <= 8'b00000000; // 1913 :   0 - 0x0
      12'h77A: dout <= 8'b00000000; // 1914 :   0 - 0x0
      12'h77B: dout <= 8'b00000000; // 1915 :   0 - 0x0
      12'h77C: dout <= 8'b00000000; // 1916 :   0 - 0x0
      12'h77D: dout <= 8'b00000000; // 1917 :   0 - 0x0
      12'h77E: dout <= 8'b00000000; // 1918 :   0 - 0x0
      12'h77F: dout <= 8'b00000000; // 1919 :   0 - 0x0
      12'h780: dout <= 8'b00000000; // 1920 :   0 - 0x0 -- Sprite 0xf0
      12'h781: dout <= 8'b00000000; // 1921 :   0 - 0x0
      12'h782: dout <= 8'b00000000; // 1922 :   0 - 0x0
      12'h783: dout <= 8'b00000000; // 1923 :   0 - 0x0
      12'h784: dout <= 8'b00000000; // 1924 :   0 - 0x0
      12'h785: dout <= 8'b00000000; // 1925 :   0 - 0x0
      12'h786: dout <= 8'b00000000; // 1926 :   0 - 0x0
      12'h787: dout <= 8'b00000000; // 1927 :   0 - 0x0
      12'h788: dout <= 8'b00000000; // 1928 :   0 - 0x0 -- Sprite 0xf1
      12'h789: dout <= 8'b00000000; // 1929 :   0 - 0x0
      12'h78A: dout <= 8'b00000000; // 1930 :   0 - 0x0
      12'h78B: dout <= 8'b00000000; // 1931 :   0 - 0x0
      12'h78C: dout <= 8'b00000000; // 1932 :   0 - 0x0
      12'h78D: dout <= 8'b00000000; // 1933 :   0 - 0x0
      12'h78E: dout <= 8'b00000000; // 1934 :   0 - 0x0
      12'h78F: dout <= 8'b00000000; // 1935 :   0 - 0x0
      12'h790: dout <= 8'b00000000; // 1936 :   0 - 0x0 -- Sprite 0xf2
      12'h791: dout <= 8'b00000000; // 1937 :   0 - 0x0
      12'h792: dout <= 8'b00000000; // 1938 :   0 - 0x0
      12'h793: dout <= 8'b00000000; // 1939 :   0 - 0x0
      12'h794: dout <= 8'b00000000; // 1940 :   0 - 0x0
      12'h795: dout <= 8'b00000000; // 1941 :   0 - 0x0
      12'h796: dout <= 8'b00000000; // 1942 :   0 - 0x0
      12'h797: dout <= 8'b00000000; // 1943 :   0 - 0x0
      12'h798: dout <= 8'b00000000; // 1944 :   0 - 0x0 -- Sprite 0xf3
      12'h799: dout <= 8'b00000000; // 1945 :   0 - 0x0
      12'h79A: dout <= 8'b00000000; // 1946 :   0 - 0x0
      12'h79B: dout <= 8'b00000000; // 1947 :   0 - 0x0
      12'h79C: dout <= 8'b00000000; // 1948 :   0 - 0x0
      12'h79D: dout <= 8'b00000000; // 1949 :   0 - 0x0
      12'h79E: dout <= 8'b00000000; // 1950 :   0 - 0x0
      12'h79F: dout <= 8'b00000000; // 1951 :   0 - 0x0
      12'h7A0: dout <= 8'b00000000; // 1952 :   0 - 0x0 -- Sprite 0xf4
      12'h7A1: dout <= 8'b00000000; // 1953 :   0 - 0x0
      12'h7A2: dout <= 8'b00000000; // 1954 :   0 - 0x0
      12'h7A3: dout <= 8'b00000000; // 1955 :   0 - 0x0
      12'h7A4: dout <= 8'b00000000; // 1956 :   0 - 0x0
      12'h7A5: dout <= 8'b00000000; // 1957 :   0 - 0x0
      12'h7A6: dout <= 8'b00000000; // 1958 :   0 - 0x0
      12'h7A7: dout <= 8'b00000000; // 1959 :   0 - 0x0
      12'h7A8: dout <= 8'b00000000; // 1960 :   0 - 0x0 -- Sprite 0xf5
      12'h7A9: dout <= 8'b00000000; // 1961 :   0 - 0x0
      12'h7AA: dout <= 8'b00000000; // 1962 :   0 - 0x0
      12'h7AB: dout <= 8'b00000000; // 1963 :   0 - 0x0
      12'h7AC: dout <= 8'b00000000; // 1964 :   0 - 0x0
      12'h7AD: dout <= 8'b00000000; // 1965 :   0 - 0x0
      12'h7AE: dout <= 8'b00000000; // 1966 :   0 - 0x0
      12'h7AF: dout <= 8'b00000000; // 1967 :   0 - 0x0
      12'h7B0: dout <= 8'b00000000; // 1968 :   0 - 0x0 -- Sprite 0xf6
      12'h7B1: dout <= 8'b00000000; // 1969 :   0 - 0x0
      12'h7B2: dout <= 8'b00000000; // 1970 :   0 - 0x0
      12'h7B3: dout <= 8'b00000000; // 1971 :   0 - 0x0
      12'h7B4: dout <= 8'b00000000; // 1972 :   0 - 0x0
      12'h7B5: dout <= 8'b00000000; // 1973 :   0 - 0x0
      12'h7B6: dout <= 8'b00000000; // 1974 :   0 - 0x0
      12'h7B7: dout <= 8'b00000000; // 1975 :   0 - 0x0
      12'h7B8: dout <= 8'b00000000; // 1976 :   0 - 0x0 -- Sprite 0xf7
      12'h7B9: dout <= 8'b00000000; // 1977 :   0 - 0x0
      12'h7BA: dout <= 8'b00000000; // 1978 :   0 - 0x0
      12'h7BB: dout <= 8'b00000000; // 1979 :   0 - 0x0
      12'h7BC: dout <= 8'b00000000; // 1980 :   0 - 0x0
      12'h7BD: dout <= 8'b00000000; // 1981 :   0 - 0x0
      12'h7BE: dout <= 8'b00000000; // 1982 :   0 - 0x0
      12'h7BF: dout <= 8'b00000000; // 1983 :   0 - 0x0
      12'h7C0: dout <= 8'b00000000; // 1984 :   0 - 0x0 -- Sprite 0xf8
      12'h7C1: dout <= 8'b00000000; // 1985 :   0 - 0x0
      12'h7C2: dout <= 8'b00000000; // 1986 :   0 - 0x0
      12'h7C3: dout <= 8'b00000000; // 1987 :   0 - 0x0
      12'h7C4: dout <= 8'b00000000; // 1988 :   0 - 0x0
      12'h7C5: dout <= 8'b00000000; // 1989 :   0 - 0x0
      12'h7C6: dout <= 8'b00000000; // 1990 :   0 - 0x0
      12'h7C7: dout <= 8'b00000000; // 1991 :   0 - 0x0
      12'h7C8: dout <= 8'b00000000; // 1992 :   0 - 0x0 -- Sprite 0xf9
      12'h7C9: dout <= 8'b00000000; // 1993 :   0 - 0x0
      12'h7CA: dout <= 8'b00000000; // 1994 :   0 - 0x0
      12'h7CB: dout <= 8'b00000000; // 1995 :   0 - 0x0
      12'h7CC: dout <= 8'b00000000; // 1996 :   0 - 0x0
      12'h7CD: dout <= 8'b00000000; // 1997 :   0 - 0x0
      12'h7CE: dout <= 8'b00000000; // 1998 :   0 - 0x0
      12'h7CF: dout <= 8'b00000000; // 1999 :   0 - 0x0
      12'h7D0: dout <= 8'b00000000; // 2000 :   0 - 0x0 -- Sprite 0xfa
      12'h7D1: dout <= 8'b00000000; // 2001 :   0 - 0x0
      12'h7D2: dout <= 8'b00000000; // 2002 :   0 - 0x0
      12'h7D3: dout <= 8'b00000000; // 2003 :   0 - 0x0
      12'h7D4: dout <= 8'b00000000; // 2004 :   0 - 0x0
      12'h7D5: dout <= 8'b00000000; // 2005 :   0 - 0x0
      12'h7D6: dout <= 8'b00000000; // 2006 :   0 - 0x0
      12'h7D7: dout <= 8'b00000000; // 2007 :   0 - 0x0
      12'h7D8: dout <= 8'b00000000; // 2008 :   0 - 0x0 -- Sprite 0xfb
      12'h7D9: dout <= 8'b00000000; // 2009 :   0 - 0x0
      12'h7DA: dout <= 8'b00000000; // 2010 :   0 - 0x0
      12'h7DB: dout <= 8'b00000000; // 2011 :   0 - 0x0
      12'h7DC: dout <= 8'b00000000; // 2012 :   0 - 0x0
      12'h7DD: dout <= 8'b00000000; // 2013 :   0 - 0x0
      12'h7DE: dout <= 8'b00000000; // 2014 :   0 - 0x0
      12'h7DF: dout <= 8'b00000000; // 2015 :   0 - 0x0
      12'h7E0: dout <= 8'b00000000; // 2016 :   0 - 0x0 -- Sprite 0xfc
      12'h7E1: dout <= 8'b00000000; // 2017 :   0 - 0x0
      12'h7E2: dout <= 8'b00000000; // 2018 :   0 - 0x0
      12'h7E3: dout <= 8'b00000000; // 2019 :   0 - 0x0
      12'h7E4: dout <= 8'b00000000; // 2020 :   0 - 0x0
      12'h7E5: dout <= 8'b00000000; // 2021 :   0 - 0x0
      12'h7E6: dout <= 8'b00000000; // 2022 :   0 - 0x0
      12'h7E7: dout <= 8'b00000000; // 2023 :   0 - 0x0
      12'h7E8: dout <= 8'b00000000; // 2024 :   0 - 0x0 -- Sprite 0xfd
      12'h7E9: dout <= 8'b00000000; // 2025 :   0 - 0x0
      12'h7EA: dout <= 8'b00000000; // 2026 :   0 - 0x0
      12'h7EB: dout <= 8'b00000000; // 2027 :   0 - 0x0
      12'h7EC: dout <= 8'b00000000; // 2028 :   0 - 0x0
      12'h7ED: dout <= 8'b00000000; // 2029 :   0 - 0x0
      12'h7EE: dout <= 8'b00000000; // 2030 :   0 - 0x0
      12'h7EF: dout <= 8'b00000000; // 2031 :   0 - 0x0
      12'h7F0: dout <= 8'b00000000; // 2032 :   0 - 0x0 -- Sprite 0xfe
      12'h7F1: dout <= 8'b00000000; // 2033 :   0 - 0x0
      12'h7F2: dout <= 8'b00000000; // 2034 :   0 - 0x0
      12'h7F3: dout <= 8'b00000000; // 2035 :   0 - 0x0
      12'h7F4: dout <= 8'b00000000; // 2036 :   0 - 0x0
      12'h7F5: dout <= 8'b00000000; // 2037 :   0 - 0x0
      12'h7F6: dout <= 8'b00000000; // 2038 :   0 - 0x0
      12'h7F7: dout <= 8'b00000000; // 2039 :   0 - 0x0
      12'h7F8: dout <= 8'b00000000; // 2040 :   0 - 0x0 -- Sprite 0xff
      12'h7F9: dout <= 8'b00000000; // 2041 :   0 - 0x0
      12'h7FA: dout <= 8'b00000000; // 2042 :   0 - 0x0
      12'h7FB: dout <= 8'b00000000; // 2043 :   0 - 0x0
      12'h7FC: dout <= 8'b00000000; // 2044 :   0 - 0x0
      12'h7FD: dout <= 8'b00000000; // 2045 :   0 - 0x0
      12'h7FE: dout <= 8'b00000000; // 2046 :   0 - 0x0
      12'h7FF: dout <= 8'b00000000; // 2047 :   0 - 0x0
          // Background pattern Table
      12'h800: dout <= 8'b00000000; // 2048 :   0 - 0x0 -- Background 0x0
      12'h801: dout <= 8'b00000000; // 2049 :   0 - 0x0
      12'h802: dout <= 8'b00000011; // 2050 :   3 - 0x3
      12'h803: dout <= 8'b00000001; // 2051 :   1 - 0x1
      12'h804: dout <= 8'b00000001; // 2052 :   1 - 0x1
      12'h805: dout <= 8'b00000000; // 2053 :   0 - 0x0
      12'h806: dout <= 8'b00000011; // 2054 :   3 - 0x3
      12'h807: dout <= 8'b00000001; // 2055 :   1 - 0x1
      12'h808: dout <= 8'b00000000; // 2056 :   0 - 0x0 -- Background 0x1
      12'h809: dout <= 8'b00000000; // 2057 :   0 - 0x0
      12'h80A: dout <= 8'b00111000; // 2058 :  56 - 0x38
      12'h80B: dout <= 8'b10110100; // 2059 : 180 - 0xb4
      12'h80C: dout <= 8'b10101000; // 2060 : 168 - 0xa8
      12'h80D: dout <= 8'b11010100; // 2061 : 212 - 0xd4
      12'h80E: dout <= 8'b01110100; // 2062 : 116 - 0x74
      12'h80F: dout <= 8'b01111110; // 2063 : 126 - 0x7e
      12'h810: dout <= 8'b00111000; // 2064 :  56 - 0x38 -- Background 0x2
      12'h811: dout <= 8'b01111000; // 2065 : 120 - 0x78
      12'h812: dout <= 8'b01111100; // 2066 : 124 - 0x7c
      12'h813: dout <= 8'b01111110; // 2067 : 126 - 0x7e
      12'h814: dout <= 8'b01111110; // 2068 : 126 - 0x7e
      12'h815: dout <= 8'b01111110; // 2069 : 126 - 0x7e
      12'h816: dout <= 8'b00111110; // 2070 :  62 - 0x3e
      12'h817: dout <= 8'b00011110; // 2071 :  30 - 0x1e
      12'h818: dout <= 8'b11110110; // 2072 : 246 - 0xf6 -- Background 0x3
      12'h819: dout <= 8'b11110000; // 2073 : 240 - 0xf0
      12'h81A: dout <= 8'b00111000; // 2074 :  56 - 0x38
      12'h81B: dout <= 8'b11010000; // 2075 : 208 - 0xd0
      12'h81C: dout <= 8'b11100000; // 2076 : 224 - 0xe0
      12'h81D: dout <= 8'b01110000; // 2077 : 112 - 0x70
      12'h81E: dout <= 8'b10111000; // 2078 : 184 - 0xb8
      12'h81F: dout <= 8'b01000000; // 2079 :  64 - 0x40
      12'h820: dout <= 8'b00011100; // 2080 :  28 - 0x1c -- Background 0x4
      12'h821: dout <= 8'b00011100; // 2081 :  28 - 0x1c
      12'h822: dout <= 8'b00011110; // 2082 :  30 - 0x1e
      12'h823: dout <= 8'b00011111; // 2083 :  31 - 0x1f
      12'h824: dout <= 8'b00001100; // 2084 :  12 - 0xc
      12'h825: dout <= 8'b00000000; // 2085 :   0 - 0x0
      12'h826: dout <= 8'b00000000; // 2086 :   0 - 0x0
      12'h827: dout <= 8'b00000000; // 2087 :   0 - 0x0
      12'h828: dout <= 8'b10101000; // 2088 : 168 - 0xa8 -- Background 0x5
      12'h829: dout <= 8'b01010000; // 2089 :  80 - 0x50
      12'h82A: dout <= 8'b10101000; // 2090 : 168 - 0xa8
      12'h82B: dout <= 8'b00000000; // 2091 :   0 - 0x0
      12'h82C: dout <= 8'b01100000; // 2092 :  96 - 0x60
      12'h82D: dout <= 8'b01100000; // 2093 :  96 - 0x60
      12'h82E: dout <= 8'b01110000; // 2094 : 112 - 0x70
      12'h82F: dout <= 8'b00000000; // 2095 :   0 - 0x0
      12'h830: dout <= 8'b00011100; // 2096 :  28 - 0x1c -- Background 0x6
      12'h831: dout <= 8'b00011100; // 2097 :  28 - 0x1c
      12'h832: dout <= 8'b00011110; // 2098 :  30 - 0x1e
      12'h833: dout <= 8'b00011111; // 2099 :  31 - 0x1f
      12'h834: dout <= 8'b00001100; // 2100 :  12 - 0xc
      12'h835: dout <= 8'b00000000; // 2101 :   0 - 0x0
      12'h836: dout <= 8'b00000001; // 2102 :   1 - 0x1
      12'h837: dout <= 8'b00000000; // 2103 :   0 - 0x0
      12'h838: dout <= 8'b10101000; // 2104 : 168 - 0xa8 -- Background 0x7
      12'h839: dout <= 8'b01010000; // 2105 :  80 - 0x50
      12'h83A: dout <= 8'b10101000; // 2106 : 168 - 0xa8
      12'h83B: dout <= 8'b00000000; // 2107 :   0 - 0x0
      12'h83C: dout <= 8'b01011000; // 2108 :  88 - 0x58
      12'h83D: dout <= 8'b11011000; // 2109 : 216 - 0xd8
      12'h83E: dout <= 8'b10001100; // 2110 : 140 - 0x8c
      12'h83F: dout <= 8'b00000000; // 2111 :   0 - 0x0
      12'h840: dout <= 8'b00011100; // 2112 :  28 - 0x1c -- Background 0x8
      12'h841: dout <= 8'b00011100; // 2113 :  28 - 0x1c
      12'h842: dout <= 8'b00011110; // 2114 :  30 - 0x1e
      12'h843: dout <= 8'b00011111; // 2115 :  31 - 0x1f
      12'h844: dout <= 8'b00001100; // 2116 :  12 - 0xc
      12'h845: dout <= 8'b00000000; // 2117 :   0 - 0x0
      12'h846: dout <= 8'b00000000; // 2118 :   0 - 0x0
      12'h847: dout <= 8'b00000000; // 2119 :   0 - 0x0
      12'h848: dout <= 8'b10101000; // 2120 : 168 - 0xa8 -- Background 0x9
      12'h849: dout <= 8'b01010100; // 2121 :  84 - 0x54
      12'h84A: dout <= 8'b10101000; // 2122 : 168 - 0xa8
      12'h84B: dout <= 8'b00000000; // 2123 :   0 - 0x0
      12'h84C: dout <= 8'b01101110; // 2124 : 110 - 0x6e
      12'h84D: dout <= 8'b11000000; // 2125 : 192 - 0xc0
      12'h84E: dout <= 8'b10000000; // 2126 : 128 - 0x80
      12'h84F: dout <= 8'b00000000; // 2127 :   0 - 0x0
      12'h850: dout <= 8'b00011100; // 2128 :  28 - 0x1c -- Background 0xa
      12'h851: dout <= 8'b00011100; // 2129 :  28 - 0x1c
      12'h852: dout <= 8'b00011110; // 2130 :  30 - 0x1e
      12'h853: dout <= 8'b00011111; // 2131 :  31 - 0x1f
      12'h854: dout <= 8'b00001100; // 2132 :  12 - 0xc
      12'h855: dout <= 8'b00000001; // 2133 :   1 - 0x1
      12'h856: dout <= 8'b00000000; // 2134 :   0 - 0x0
      12'h857: dout <= 8'b00000000; // 2135 :   0 - 0x0
      12'h858: dout <= 8'b10101000; // 2136 : 168 - 0xa8 -- Background 0xb
      12'h859: dout <= 8'b01010100; // 2137 :  84 - 0x54
      12'h85A: dout <= 8'b10101000; // 2138 : 168 - 0xa8
      12'h85B: dout <= 8'b00000000; // 2139 :   0 - 0x0
      12'h85C: dout <= 8'b11011000; // 2140 : 216 - 0xd8
      12'h85D: dout <= 8'b11011100; // 2141 : 220 - 0xdc
      12'h85E: dout <= 8'b00001100; // 2142 :  12 - 0xc
      12'h85F: dout <= 8'b00000000; // 2143 :   0 - 0x0
      12'h860: dout <= 8'b11110110; // 2144 : 246 - 0xf6 -- Background 0xc
      12'h861: dout <= 8'b11110000; // 2145 : 240 - 0xf0
      12'h862: dout <= 8'b00000000; // 2146 :   0 - 0x0
      12'h863: dout <= 8'b11111100; // 2147 : 252 - 0xfc
      12'h864: dout <= 8'b11111000; // 2148 : 248 - 0xf8
      12'h865: dout <= 8'b00000000; // 2149 :   0 - 0x0
      12'h866: dout <= 8'b10101000; // 2150 : 168 - 0xa8
      12'h867: dout <= 8'b01010100; // 2151 :  84 - 0x54
      12'h868: dout <= 8'b00111000; // 2152 :  56 - 0x38 -- Background 0xd
      12'h869: dout <= 8'b01111000; // 2153 : 120 - 0x78
      12'h86A: dout <= 8'b01111100; // 2154 : 124 - 0x7c
      12'h86B: dout <= 8'b01111101; // 2155 : 125 - 0x7d
      12'h86C: dout <= 8'b01111101; // 2156 : 125 - 0x7d
      12'h86D: dout <= 8'b01111011; // 2157 : 123 - 0x7b
      12'h86E: dout <= 8'b00111011; // 2158 :  59 - 0x3b
      12'h86F: dout <= 8'b00011011; // 2159 :  27 - 0x1b
      12'h870: dout <= 8'b11110110; // 2160 : 246 - 0xf6 -- Background 0xe
      12'h871: dout <= 8'b11110000; // 2161 : 240 - 0xf0
      12'h872: dout <= 8'b01111000; // 2162 : 120 - 0x78
      12'h873: dout <= 8'b01110000; // 2163 : 112 - 0x70
      12'h874: dout <= 8'b10100000; // 2164 : 160 - 0xa0
      12'h875: dout <= 8'b10010000; // 2165 : 144 - 0x90
      12'h876: dout <= 8'b00101000; // 2166 :  40 - 0x28
      12'h877: dout <= 8'b01010100; // 2167 :  84 - 0x54
      12'h878: dout <= 8'b00000000; // 2168 :   0 - 0x0 -- Background 0xf
      12'h879: dout <= 8'b00000000; // 2169 :   0 - 0x0
      12'h87A: dout <= 8'b00000011; // 2170 :   3 - 0x3
      12'h87B: dout <= 8'b00000001; // 2171 :   1 - 0x1
      12'h87C: dout <= 8'b00000001; // 2172 :   1 - 0x1
      12'h87D: dout <= 8'b00000000; // 2173 :   0 - 0x0
      12'h87E: dout <= 8'b00000011; // 2174 :   3 - 0x3
      12'h87F: dout <= 8'b00000001; // 2175 :   1 - 0x1
      12'h880: dout <= 8'b00000000; // 2176 :   0 - 0x0 -- Background 0x10
      12'h881: dout <= 8'b00000011; // 2177 :   3 - 0x3
      12'h882: dout <= 8'b00001111; // 2178 :  15 - 0xf
      12'h883: dout <= 8'b00001111; // 2179 :  15 - 0xf
      12'h884: dout <= 8'b00001111; // 2180 :  15 - 0xf
      12'h885: dout <= 8'b00011111; // 2181 :  31 - 0x1f
      12'h886: dout <= 8'b00011111; // 2182 :  31 - 0x1f
      12'h887: dout <= 8'b00011110; // 2183 :  30 - 0x1e
      12'h888: dout <= 8'b00110110; // 2184 :  54 - 0x36 -- Background 0x11
      12'h889: dout <= 8'b10110000; // 2185 : 176 - 0xb0
      12'h88A: dout <= 8'b10111000; // 2186 : 184 - 0xb8
      12'h88B: dout <= 8'b10010000; // 2187 : 144 - 0x90
      12'h88C: dout <= 8'b10100000; // 2188 : 160 - 0xa0
      12'h88D: dout <= 8'b01110000; // 2189 : 112 - 0x70
      12'h88E: dout <= 8'b00111000; // 2190 :  56 - 0x38
      12'h88F: dout <= 8'b01000000; // 2191 :  64 - 0x40
      12'h890: dout <= 8'b00011100; // 2192 :  28 - 0x1c -- Background 0x12
      12'h891: dout <= 8'b00011100; // 2193 :  28 - 0x1c
      12'h892: dout <= 8'b00011110; // 2194 :  30 - 0x1e
      12'h893: dout <= 8'b00011111; // 2195 :  31 - 0x1f
      12'h894: dout <= 8'b00001100; // 2196 :  12 - 0xc
      12'h895: dout <= 8'b00000000; // 2197 :   0 - 0x0
      12'h896: dout <= 8'b00000000; // 2198 :   0 - 0x0
      12'h897: dout <= 8'b00000000; // 2199 :   0 - 0x0
      12'h898: dout <= 8'b00000000; // 2200 :   0 - 0x0 -- Background 0x13
      12'h899: dout <= 8'b00000000; // 2201 :   0 - 0x0
      12'h89A: dout <= 8'b00000000; // 2202 :   0 - 0x0
      12'h89B: dout <= 8'b00000011; // 2203 :   3 - 0x3
      12'h89C: dout <= 8'b00000111; // 2204 :   7 - 0x7
      12'h89D: dout <= 8'b00001111; // 2205 :  15 - 0xf
      12'h89E: dout <= 8'b00001111; // 2206 :  15 - 0xf
      12'h89F: dout <= 8'b00011111; // 2207 :  31 - 0x1f
      12'h8A0: dout <= 8'b11110110; // 2208 : 246 - 0xf6 -- Background 0x14
      12'h8A1: dout <= 8'b00000000; // 2209 :   0 - 0x0
      12'h8A2: dout <= 8'b11111000; // 2210 : 248 - 0xf8
      12'h8A3: dout <= 8'b11111110; // 2211 : 254 - 0xfe
      12'h8A4: dout <= 8'b11111110; // 2212 : 254 - 0xfe
      12'h8A5: dout <= 8'b11111110; // 2213 : 254 - 0xfe
      12'h8A6: dout <= 8'b11111000; // 2214 : 248 - 0xf8
      12'h8A7: dout <= 8'b00000000; // 2215 :   0 - 0x0
      12'h8A8: dout <= 8'b00000011; // 2216 :   3 - 0x3 -- Background 0x15
      12'h8A9: dout <= 8'b00000011; // 2217 :   3 - 0x3
      12'h8AA: dout <= 8'b00000000; // 2218 :   0 - 0x0
      12'h8AB: dout <= 8'b00000011; // 2219 :   3 - 0x3
      12'h8AC: dout <= 8'b00000011; // 2220 :   3 - 0x3
      12'h8AD: dout <= 8'b00000000; // 2221 :   0 - 0x0
      12'h8AE: dout <= 8'b00001111; // 2222 :  15 - 0xf
      12'h8AF: dout <= 8'b00111111; // 2223 :  63 - 0x3f
      12'h8B0: dout <= 8'b11011000; // 2224 : 216 - 0xd8 -- Background 0x16
      12'h8B1: dout <= 8'b11000000; // 2225 : 192 - 0xc0
      12'h8B2: dout <= 8'b11100000; // 2226 : 224 - 0xe0
      12'h8B3: dout <= 8'b01000000; // 2227 :  64 - 0x40
      12'h8B4: dout <= 8'b10000000; // 2228 : 128 - 0x80
      12'h8B5: dout <= 8'b00000000; // 2229 :   0 - 0x0
      12'h8B6: dout <= 8'b11100000; // 2230 : 224 - 0xe0
      12'h8B7: dout <= 8'b11111100; // 2231 : 252 - 0xfc
      12'h8B8: dout <= 8'b01111111; // 2232 : 127 - 0x7f -- Background 0x17
      12'h8B9: dout <= 8'b01111111; // 2233 : 127 - 0x7f
      12'h8BA: dout <= 8'b01111111; // 2234 : 127 - 0x7f
      12'h8BB: dout <= 8'b01111100; // 2235 : 124 - 0x7c
      12'h8BC: dout <= 8'b00110000; // 2236 :  48 - 0x30
      12'h8BD: dout <= 8'b00000001; // 2237 :   1 - 0x1
      12'h8BE: dout <= 8'b00000001; // 2238 :   1 - 0x1
      12'h8BF: dout <= 8'b00000000; // 2239 :   0 - 0x0
      12'h8C0: dout <= 8'b11111100; // 2240 : 252 - 0xfc -- Background 0x18
      12'h8C1: dout <= 8'b11111110; // 2241 : 254 - 0xfe
      12'h8C2: dout <= 8'b11111100; // 2242 : 252 - 0xfc
      12'h8C3: dout <= 8'b00000000; // 2243 :   0 - 0x0
      12'h8C4: dout <= 8'b00000000; // 2244 :   0 - 0x0
      12'h8C5: dout <= 8'b10000000; // 2245 : 128 - 0x80
      12'h8C6: dout <= 8'b11000000; // 2246 : 192 - 0xc0
      12'h8C7: dout <= 8'b00000000; // 2247 :   0 - 0x0
      12'h8C8: dout <= 8'b00000111; // 2248 :   7 - 0x7 -- Background 0x19
      12'h8C9: dout <= 8'b00000111; // 2249 :   7 - 0x7
      12'h8CA: dout <= 8'b00000001; // 2250 :   1 - 0x1
      12'h8CB: dout <= 8'b00000110; // 2251 :   6 - 0x6
      12'h8CC: dout <= 8'b00000111; // 2252 :   7 - 0x7
      12'h8CD: dout <= 8'b00000110; // 2253 :   6 - 0x6
      12'h8CE: dout <= 8'b00000000; // 2254 :   0 - 0x0
      12'h8CF: dout <= 8'b00001111; // 2255 :  15 - 0xf
      12'h8D0: dout <= 8'b10110000; // 2256 : 176 - 0xb0 -- Background 0x1a
      12'h8D1: dout <= 8'b10000000; // 2257 : 128 - 0x80
      12'h8D2: dout <= 8'b11000000; // 2258 : 192 - 0xc0
      12'h8D3: dout <= 8'b10000000; // 2259 : 128 - 0x80
      12'h8D4: dout <= 8'b00000000; // 2260 :   0 - 0x0
      12'h8D5: dout <= 8'b00000000; // 2261 :   0 - 0x0
      12'h8D6: dout <= 8'b00000000; // 2262 :   0 - 0x0
      12'h8D7: dout <= 8'b11100000; // 2263 : 224 - 0xe0
      12'h8D8: dout <= 8'b00111111; // 2264 :  63 - 0x3f -- Background 0x1b
      12'h8D9: dout <= 8'b00111111; // 2265 :  63 - 0x3f
      12'h8DA: dout <= 8'b01111111; // 2266 : 127 - 0x7f
      12'h8DB: dout <= 8'b01111111; // 2267 : 127 - 0x7f
      12'h8DC: dout <= 8'b00111111; // 2268 :  63 - 0x3f
      12'h8DD: dout <= 8'b00000000; // 2269 :   0 - 0x0
      12'h8DE: dout <= 8'b00000011; // 2270 :   3 - 0x3
      12'h8DF: dout <= 8'b00000000; // 2271 :   0 - 0x0
      12'h8E0: dout <= 8'b11111111; // 2272 : 255 - 0xff -- Background 0x1c
      12'h8E1: dout <= 8'b11111111; // 2273 : 255 - 0xff
      12'h8E2: dout <= 8'b11111111; // 2274 : 255 - 0xff
      12'h8E3: dout <= 8'b11111111; // 2275 : 255 - 0xff
      12'h8E4: dout <= 8'b11111111; // 2276 : 255 - 0xff
      12'h8E5: dout <= 8'b00000000; // 2277 :   0 - 0x0
      12'h8E6: dout <= 8'b10000000; // 2278 : 128 - 0x80
      12'h8E7: dout <= 8'b00000000; // 2279 :   0 - 0x0
      12'h8E8: dout <= 8'b00000000; // 2280 :   0 - 0x0 -- Background 0x1d
      12'h8E9: dout <= 8'b11000000; // 2281 : 192 - 0xc0
      12'h8EA: dout <= 8'b11000000; // 2282 : 192 - 0xc0
      12'h8EB: dout <= 8'b11000000; // 2283 : 192 - 0xc0
      12'h8EC: dout <= 8'b10000000; // 2284 : 128 - 0x80
      12'h8ED: dout <= 8'b00000000; // 2285 :   0 - 0x0
      12'h8EE: dout <= 8'b00000000; // 2286 :   0 - 0x0
      12'h8EF: dout <= 8'b00000000; // 2287 :   0 - 0x0
      12'h8F0: dout <= 8'b11100000; // 2288 : 224 - 0xe0 -- Background 0x1e
      12'h8F1: dout <= 8'b10011100; // 2289 : 156 - 0x9c
      12'h8F2: dout <= 8'b00111000; // 2290 :  56 - 0x38
      12'h8F3: dout <= 8'b11100000; // 2291 : 224 - 0xe0
      12'h8F4: dout <= 8'b11001000; // 2292 : 200 - 0xc8
      12'h8F5: dout <= 8'b00010100; // 2293 :  20 - 0x14
      12'h8F6: dout <= 8'b10101000; // 2294 : 168 - 0xa8
      12'h8F7: dout <= 8'b01010100; // 2295 :  84 - 0x54
      12'h8F8: dout <= 8'b00000000; // 2296 :   0 - 0x0 -- Background 0x1f
      12'h8F9: dout <= 8'b00000000; // 2297 :   0 - 0x0
      12'h8FA: dout <= 8'b00111000; // 2298 :  56 - 0x38
      12'h8FB: dout <= 8'b10110100; // 2299 : 180 - 0xb4
      12'h8FC: dout <= 8'b10101000; // 2300 : 168 - 0xa8
      12'h8FD: dout <= 8'b11010100; // 2301 : 212 - 0xd4
      12'h8FE: dout <= 8'b01110100; // 2302 : 116 - 0x74
      12'h8FF: dout <= 8'b00011110; // 2303 :  30 - 0x1e
      12'h900: dout <= 8'b00000000; // 2304 :   0 - 0x0 -- Background 0x20
      12'h901: dout <= 8'b00000000; // 2305 :   0 - 0x0
      12'h902: dout <= 8'b00001100; // 2306 :  12 - 0xc
      12'h903: dout <= 8'b00000111; // 2307 :   7 - 0x7
      12'h904: dout <= 8'b00001111; // 2308 :  15 - 0xf
      12'h905: dout <= 8'b00000111; // 2309 :   7 - 0x7
      12'h906: dout <= 8'b00001111; // 2310 :  15 - 0xf
      12'h907: dout <= 8'b00001111; // 2311 :  15 - 0xf
      12'h908: dout <= 8'b00000000; // 2312 :   0 - 0x0 -- Background 0x21
      12'h909: dout <= 8'b00000000; // 2313 :   0 - 0x0
      12'h90A: dout <= 8'b00110000; // 2314 :  48 - 0x30
      12'h90B: dout <= 8'b11100000; // 2315 : 224 - 0xe0
      12'h90C: dout <= 8'b11110000; // 2316 : 240 - 0xf0
      12'h90D: dout <= 8'b11100000; // 2317 : 224 - 0xe0
      12'h90E: dout <= 8'b11110000; // 2318 : 240 - 0xf0
      12'h90F: dout <= 8'b11110000; // 2319 : 240 - 0xf0
      12'h910: dout <= 8'b00000111; // 2320 :   7 - 0x7 -- Background 0x22
      12'h911: dout <= 8'b00000011; // 2321 :   3 - 0x3
      12'h912: dout <= 8'b00011000; // 2322 :  24 - 0x18
      12'h913: dout <= 8'b00010101; // 2323 :  21 - 0x15
      12'h914: dout <= 8'b00000010; // 2324 :   2 - 0x2
      12'h915: dout <= 8'b00000101; // 2325 :   5 - 0x5
      12'h916: dout <= 8'b00000010; // 2326 :   2 - 0x2
      12'h917: dout <= 8'b00000100; // 2327 :   4 - 0x4
      12'h918: dout <= 8'b11100000; // 2328 : 224 - 0xe0 -- Background 0x23
      12'h919: dout <= 8'b11000000; // 2329 : 192 - 0xc0
      12'h91A: dout <= 8'b00111100; // 2330 :  60 - 0x3c
      12'h91B: dout <= 8'b01111100; // 2331 : 124 - 0x7c
      12'h91C: dout <= 8'b01111100; // 2332 : 124 - 0x7c
      12'h91D: dout <= 8'b01111100; // 2333 : 124 - 0x7c
      12'h91E: dout <= 8'b11101100; // 2334 : 236 - 0xec
      12'h91F: dout <= 8'b11100000; // 2335 : 224 - 0xe0
      12'h920: dout <= 8'b00000010; // 2336 :   2 - 0x2 -- Background 0x24
      12'h921: dout <= 8'b00000101; // 2337 :   5 - 0x5
      12'h922: dout <= 8'b00001011; // 2338 :  11 - 0xb
      12'h923: dout <= 8'b00001011; // 2339 :  11 - 0xb
      12'h924: dout <= 8'b00001101; // 2340 :  13 - 0xd
      12'h925: dout <= 8'b00011000; // 2341 :  24 - 0x18
      12'h926: dout <= 8'b00111000; // 2342 :  56 - 0x38
      12'h927: dout <= 8'b00000000; // 2343 :   0 - 0x0
      12'h928: dout <= 8'b11100000; // 2344 : 224 - 0xe0 -- Background 0x25
      12'h929: dout <= 8'b11100000; // 2345 : 224 - 0xe0
      12'h92A: dout <= 8'b11100000; // 2346 : 224 - 0xe0
      12'h92B: dout <= 8'b11010000; // 2347 : 208 - 0xd0
      12'h92C: dout <= 8'b10111000; // 2348 : 184 - 0xb8
      12'h92D: dout <= 8'b00111000; // 2349 :  56 - 0x38
      12'h92E: dout <= 8'b00000000; // 2350 :   0 - 0x0
      12'h92F: dout <= 8'b00000000; // 2351 :   0 - 0x0
      12'h930: dout <= 8'b00000000; // 2352 :   0 - 0x0 -- Background 0x26
      12'h931: dout <= 8'b00000000; // 2353 :   0 - 0x0
      12'h932: dout <= 8'b00000000; // 2354 :   0 - 0x0
      12'h933: dout <= 8'b00000000; // 2355 :   0 - 0x0
      12'h934: dout <= 8'b00000000; // 2356 :   0 - 0x0
      12'h935: dout <= 8'b00000000; // 2357 :   0 - 0x0
      12'h936: dout <= 8'b00000000; // 2358 :   0 - 0x0
      12'h937: dout <= 8'b00000000; // 2359 :   0 - 0x0
      12'h938: dout <= 8'b00000000; // 2360 :   0 - 0x0 -- Background 0x27
      12'h939: dout <= 8'b00000000; // 2361 :   0 - 0x0
      12'h93A: dout <= 8'b00000000; // 2362 :   0 - 0x0
      12'h93B: dout <= 8'b00000000; // 2363 :   0 - 0x0
      12'h93C: dout <= 8'b00000000; // 2364 :   0 - 0x0
      12'h93D: dout <= 8'b00000000; // 2365 :   0 - 0x0
      12'h93E: dout <= 8'b00000000; // 2366 :   0 - 0x0
      12'h93F: dout <= 8'b00000000; // 2367 :   0 - 0x0
      12'h940: dout <= 8'b00000000; // 2368 :   0 - 0x0 -- Background 0x28
      12'h941: dout <= 8'b00000000; // 2369 :   0 - 0x0
      12'h942: dout <= 8'b00000000; // 2370 :   0 - 0x0
      12'h943: dout <= 8'b00000000; // 2371 :   0 - 0x0
      12'h944: dout <= 8'b00000000; // 2372 :   0 - 0x0
      12'h945: dout <= 8'b00000000; // 2373 :   0 - 0x0
      12'h946: dout <= 8'b00000000; // 2374 :   0 - 0x0
      12'h947: dout <= 8'b00000000; // 2375 :   0 - 0x0
      12'h948: dout <= 8'b00011111; // 2376 :  31 - 0x1f -- Background 0x29
      12'h949: dout <= 8'b00011111; // 2377 :  31 - 0x1f
      12'h94A: dout <= 8'b00011111; // 2378 :  31 - 0x1f
      12'h94B: dout <= 8'b00011111; // 2379 :  31 - 0x1f
      12'h94C: dout <= 8'b00001100; // 2380 :  12 - 0xc
      12'h94D: dout <= 8'b00000000; // 2381 :   0 - 0x0
      12'h94E: dout <= 8'b00000001; // 2382 :   1 - 0x1
      12'h94F: dout <= 8'b00000000; // 2383 :   0 - 0x0
      12'h950: dout <= 8'b00011111; // 2384 :  31 - 0x1f -- Background 0x2a
      12'h951: dout <= 8'b00011111; // 2385 :  31 - 0x1f
      12'h952: dout <= 8'b00011111; // 2386 :  31 - 0x1f
      12'h953: dout <= 8'b00011111; // 2387 :  31 - 0x1f
      12'h954: dout <= 8'b00001100; // 2388 :  12 - 0xc
      12'h955: dout <= 8'b00000000; // 2389 :   0 - 0x0
      12'h956: dout <= 8'b00000000; // 2390 :   0 - 0x0
      12'h957: dout <= 8'b00000000; // 2391 :   0 - 0x0
      12'h958: dout <= 8'b00000000; // 2392 :   0 - 0x0 -- Background 0x2b
      12'h959: dout <= 8'b00000000; // 2393 :   0 - 0x0
      12'h95A: dout <= 8'b00000000; // 2394 :   0 - 0x0
      12'h95B: dout <= 8'b00000000; // 2395 :   0 - 0x0
      12'h95C: dout <= 8'b00000000; // 2396 :   0 - 0x0
      12'h95D: dout <= 8'b00000000; // 2397 :   0 - 0x0
      12'h95E: dout <= 8'b00000000; // 2398 :   0 - 0x0
      12'h95F: dout <= 8'b00000000; // 2399 :   0 - 0x0
      12'h960: dout <= 8'b00000000; // 2400 :   0 - 0x0 -- Background 0x2c
      12'h961: dout <= 8'b00000000; // 2401 :   0 - 0x0
      12'h962: dout <= 8'b00000000; // 2402 :   0 - 0x0
      12'h963: dout <= 8'b00000000; // 2403 :   0 - 0x0
      12'h964: dout <= 8'b00000000; // 2404 :   0 - 0x0
      12'h965: dout <= 8'b00000000; // 2405 :   0 - 0x0
      12'h966: dout <= 8'b00000000; // 2406 :   0 - 0x0
      12'h967: dout <= 8'b00000000; // 2407 :   0 - 0x0
      12'h968: dout <= 8'b00000000; // 2408 :   0 - 0x0 -- Background 0x2d
      12'h969: dout <= 8'b01111110; // 2409 : 126 - 0x7e
      12'h96A: dout <= 8'b01000010; // 2410 :  66 - 0x42
      12'h96B: dout <= 8'b01000010; // 2411 :  66 - 0x42
      12'h96C: dout <= 8'b01000010; // 2412 :  66 - 0x42
      12'h96D: dout <= 8'b01000010; // 2413 :  66 - 0x42
      12'h96E: dout <= 8'b01111110; // 2414 : 126 - 0x7e
      12'h96F: dout <= 8'b00000000; // 2415 :   0 - 0x0
      12'h970: dout <= 8'b00000000; // 2416 :   0 - 0x0 -- Background 0x2e
      12'h971: dout <= 8'b00000000; // 2417 :   0 - 0x0
      12'h972: dout <= 8'b00000000; // 2418 :   0 - 0x0
      12'h973: dout <= 8'b00000000; // 2419 :   0 - 0x0
      12'h974: dout <= 8'b00000000; // 2420 :   0 - 0x0
      12'h975: dout <= 8'b00000000; // 2421 :   0 - 0x0
      12'h976: dout <= 8'b00000000; // 2422 :   0 - 0x0
      12'h977: dout <= 8'b00000000; // 2423 :   0 - 0x0
      12'h978: dout <= 8'b01100110; // 2424 : 102 - 0x66 -- Background 0x2f
      12'h979: dout <= 8'b01100000; // 2425 :  96 - 0x60
      12'h97A: dout <= 8'b01101000; // 2426 : 104 - 0x68
      12'h97B: dout <= 8'b11100000; // 2427 : 224 - 0xe0
      12'h97C: dout <= 8'b11000000; // 2428 : 192 - 0xc0
      12'h97D: dout <= 8'b00010000; // 2429 :  16 - 0x10
      12'h97E: dout <= 8'b00101000; // 2430 :  40 - 0x28
      12'h97F: dout <= 8'b01010000; // 2431 :  80 - 0x50
      12'h980: dout <= 8'b11110110; // 2432 : 246 - 0xf6 -- Background 0x30
      12'h981: dout <= 8'b11110000; // 2433 : 240 - 0xf0
      12'h982: dout <= 8'b00111000; // 2434 :  56 - 0x38
      12'h983: dout <= 8'b11010000; // 2435 : 208 - 0xd0
      12'h984: dout <= 8'b11000000; // 2436 : 192 - 0xc0
      12'h985: dout <= 8'b11111000; // 2437 : 248 - 0xf8
      12'h986: dout <= 8'b01111000; // 2438 : 120 - 0x78
      12'h987: dout <= 8'b00000000; // 2439 :   0 - 0x0
      12'h988: dout <= 8'b11110110; // 2440 : 246 - 0xf6 -- Background 0x31
      12'h989: dout <= 8'b11110000; // 2441 : 240 - 0xf0
      12'h98A: dout <= 8'b00111000; // 2442 :  56 - 0x38
      12'h98B: dout <= 8'b11010000; // 2443 : 208 - 0xd0
      12'h98C: dout <= 8'b11000000; // 2444 : 192 - 0xc0
      12'h98D: dout <= 8'b11100000; // 2445 : 224 - 0xe0
      12'h98E: dout <= 8'b01111000; // 2446 : 120 - 0x78
      12'h98F: dout <= 8'b00111000; // 2447 :  56 - 0x38
      12'h990: dout <= 8'b11110110; // 2448 : 246 - 0xf6 -- Background 0x32
      12'h991: dout <= 8'b11110000; // 2449 : 240 - 0xf0
      12'h992: dout <= 8'b00111000; // 2450 :  56 - 0x38
      12'h993: dout <= 8'b11000000; // 2451 : 192 - 0xc0
      12'h994: dout <= 8'b11011000; // 2452 : 216 - 0xd8
      12'h995: dout <= 8'b11111000; // 2453 : 248 - 0xf8
      12'h996: dout <= 8'b01100000; // 2454 :  96 - 0x60
      12'h997: dout <= 8'b00010000; // 2455 :  16 - 0x10
      12'h998: dout <= 8'b00011100; // 2456 :  28 - 0x1c -- Background 0x33
      12'h999: dout <= 8'b00011100; // 2457 :  28 - 0x1c
      12'h99A: dout <= 8'b00011110; // 2458 :  30 - 0x1e
      12'h99B: dout <= 8'b00011111; // 2459 :  31 - 0x1f
      12'h99C: dout <= 8'b00001100; // 2460 :  12 - 0xc
      12'h99D: dout <= 8'b00000000; // 2461 :   0 - 0x0
      12'h99E: dout <= 8'b00000000; // 2462 :   0 - 0x0
      12'h99F: dout <= 8'b00000000; // 2463 :   0 - 0x0
      12'h9A0: dout <= 8'b10000000; // 2464 : 128 - 0x80 -- Background 0x34
      12'h9A1: dout <= 8'b01010000; // 2465 :  80 - 0x50
      12'h9A2: dout <= 8'b10101000; // 2466 : 168 - 0xa8
      12'h9A3: dout <= 8'b00000000; // 2467 :   0 - 0x0
      12'h9A4: dout <= 8'b01011000; // 2468 :  88 - 0x58
      12'h9A5: dout <= 8'b11011000; // 2469 : 216 - 0xd8
      12'h9A6: dout <= 8'b11101100; // 2470 : 236 - 0xec
      12'h9A7: dout <= 8'b00000000; // 2471 :   0 - 0x0
      12'h9A8: dout <= 8'b00011100; // 2472 :  28 - 0x1c -- Background 0x35
      12'h9A9: dout <= 8'b00011100; // 2473 :  28 - 0x1c
      12'h9AA: dout <= 8'b00011110; // 2474 :  30 - 0x1e
      12'h9AB: dout <= 8'b00011111; // 2475 :  31 - 0x1f
      12'h9AC: dout <= 8'b00001100; // 2476 :  12 - 0xc
      12'h9AD: dout <= 8'b00000001; // 2477 :   1 - 0x1
      12'h9AE: dout <= 8'b00000001; // 2478 :   1 - 0x1
      12'h9AF: dout <= 8'b00000000; // 2479 :   0 - 0x0
      12'h9B0: dout <= 8'b10101000; // 2480 : 168 - 0xa8 -- Background 0x36
      12'h9B1: dout <= 8'b01010000; // 2481 :  80 - 0x50
      12'h9B2: dout <= 8'b10101000; // 2482 : 168 - 0xa8
      12'h9B3: dout <= 8'b00000000; // 2483 :   0 - 0x0
      12'h9B4: dout <= 8'b01011000; // 2484 :  88 - 0x58
      12'h9B5: dout <= 8'b11001110; // 2485 : 206 - 0xce
      12'h9B6: dout <= 8'b10000110; // 2486 : 134 - 0x86
      12'h9B7: dout <= 8'b00000000; // 2487 :   0 - 0x0
      12'h9B8: dout <= 8'b10101000; // 2488 : 168 - 0xa8 -- Background 0x37
      12'h9B9: dout <= 8'b01010000; // 2489 :  80 - 0x50
      12'h9BA: dout <= 8'b10101000; // 2490 : 168 - 0xa8
      12'h9BB: dout <= 8'b00000000; // 2491 :   0 - 0x0
      12'h9BC: dout <= 8'b01011000; // 2492 :  88 - 0x58
      12'h9BD: dout <= 8'b11011000; // 2493 : 216 - 0xd8
      12'h9BE: dout <= 8'b11101100; // 2494 : 236 - 0xec
      12'h9BF: dout <= 8'b00000000; // 2495 :   0 - 0x0
      12'h9C0: dout <= 8'b00000000; // 2496 :   0 - 0x0 -- Background 0x38
      12'h9C1: dout <= 8'b00000000; // 2497 :   0 - 0x0
      12'h9C2: dout <= 8'b00000000; // 2498 :   0 - 0x0
      12'h9C3: dout <= 8'b00000000; // 2499 :   0 - 0x0
      12'h9C4: dout <= 8'b00000000; // 2500 :   0 - 0x0
      12'h9C5: dout <= 8'b00000000; // 2501 :   0 - 0x0
      12'h9C6: dout <= 8'b00000000; // 2502 :   0 - 0x0
      12'h9C7: dout <= 8'b00000000; // 2503 :   0 - 0x0
      12'h9C8: dout <= 8'b00000000; // 2504 :   0 - 0x0 -- Background 0x39
      12'h9C9: dout <= 8'b00000000; // 2505 :   0 - 0x0
      12'h9CA: dout <= 8'b00000000; // 2506 :   0 - 0x0
      12'h9CB: dout <= 8'b00000000; // 2507 :   0 - 0x0
      12'h9CC: dout <= 8'b00000000; // 2508 :   0 - 0x0
      12'h9CD: dout <= 8'b00000000; // 2509 :   0 - 0x0
      12'h9CE: dout <= 8'b00000000; // 2510 :   0 - 0x0
      12'h9CF: dout <= 8'b00000000; // 2511 :   0 - 0x0
      12'h9D0: dout <= 8'b00000000; // 2512 :   0 - 0x0 -- Background 0x3a
      12'h9D1: dout <= 8'b00000000; // 2513 :   0 - 0x0
      12'h9D2: dout <= 8'b00000000; // 2514 :   0 - 0x0
      12'h9D3: dout <= 8'b00000000; // 2515 :   0 - 0x0
      12'h9D4: dout <= 8'b00000000; // 2516 :   0 - 0x0
      12'h9D5: dout <= 8'b00000000; // 2517 :   0 - 0x0
      12'h9D6: dout <= 8'b00000000; // 2518 :   0 - 0x0
      12'h9D7: dout <= 8'b00000000; // 2519 :   0 - 0x0
      12'h9D8: dout <= 8'b00000000; // 2520 :   0 - 0x0 -- Background 0x3b
      12'h9D9: dout <= 8'b00000000; // 2521 :   0 - 0x0
      12'h9DA: dout <= 8'b00000000; // 2522 :   0 - 0x0
      12'h9DB: dout <= 8'b00000000; // 2523 :   0 - 0x0
      12'h9DC: dout <= 8'b00000000; // 2524 :   0 - 0x0
      12'h9DD: dout <= 8'b00000000; // 2525 :   0 - 0x0
      12'h9DE: dout <= 8'b00000000; // 2526 :   0 - 0x0
      12'h9DF: dout <= 8'b00000000; // 2527 :   0 - 0x0
      12'h9E0: dout <= 8'b00000000; // 2528 :   0 - 0x0 -- Background 0x3c
      12'h9E1: dout <= 8'b00000000; // 2529 :   0 - 0x0
      12'h9E2: dout <= 8'b00000000; // 2530 :   0 - 0x0
      12'h9E3: dout <= 8'b00000000; // 2531 :   0 - 0x0
      12'h9E4: dout <= 8'b00000000; // 2532 :   0 - 0x0
      12'h9E5: dout <= 8'b00000000; // 2533 :   0 - 0x0
      12'h9E6: dout <= 8'b00000000; // 2534 :   0 - 0x0
      12'h9E7: dout <= 8'b00000000; // 2535 :   0 - 0x0
      12'h9E8: dout <= 8'b00000000; // 2536 :   0 - 0x0 -- Background 0x3d
      12'h9E9: dout <= 8'b00000000; // 2537 :   0 - 0x0
      12'h9EA: dout <= 8'b00000000; // 2538 :   0 - 0x0
      12'h9EB: dout <= 8'b00000000; // 2539 :   0 - 0x0
      12'h9EC: dout <= 8'b00000000; // 2540 :   0 - 0x0
      12'h9ED: dout <= 8'b00000000; // 2541 :   0 - 0x0
      12'h9EE: dout <= 8'b00000000; // 2542 :   0 - 0x0
      12'h9EF: dout <= 8'b00000000; // 2543 :   0 - 0x0
      12'h9F0: dout <= 8'b00000000; // 2544 :   0 - 0x0 -- Background 0x3e
      12'h9F1: dout <= 8'b00000000; // 2545 :   0 - 0x0
      12'h9F2: dout <= 8'b00000000; // 2546 :   0 - 0x0
      12'h9F3: dout <= 8'b00000000; // 2547 :   0 - 0x0
      12'h9F4: dout <= 8'b00000000; // 2548 :   0 - 0x0
      12'h9F5: dout <= 8'b00000000; // 2549 :   0 - 0x0
      12'h9F6: dout <= 8'b00000000; // 2550 :   0 - 0x0
      12'h9F7: dout <= 8'b00000000; // 2551 :   0 - 0x0
      12'h9F8: dout <= 8'b00000000; // 2552 :   0 - 0x0 -- Background 0x3f
      12'h9F9: dout <= 8'b00000000; // 2553 :   0 - 0x0
      12'h9FA: dout <= 8'b00000000; // 2554 :   0 - 0x0
      12'h9FB: dout <= 8'b00000000; // 2555 :   0 - 0x0
      12'h9FC: dout <= 8'b00000000; // 2556 :   0 - 0x0
      12'h9FD: dout <= 8'b00000000; // 2557 :   0 - 0x0
      12'h9FE: dout <= 8'b00000000; // 2558 :   0 - 0x0
      12'h9FF: dout <= 8'b00000000; // 2559 :   0 - 0x0
      12'hA00: dout <= 8'b00111100; // 2560 :  60 - 0x3c -- Background 0x40
      12'hA01: dout <= 8'b01111100; // 2561 : 124 - 0x7c
      12'hA02: dout <= 8'b11100110; // 2562 : 230 - 0xe6
      12'hA03: dout <= 8'b11101110; // 2563 : 238 - 0xee
      12'hA04: dout <= 8'b11110110; // 2564 : 246 - 0xf6
      12'hA05: dout <= 8'b11100110; // 2565 : 230 - 0xe6
      12'hA06: dout <= 8'b00111100; // 2566 :  60 - 0x3c
      12'hA07: dout <= 8'b00000000; // 2567 :   0 - 0x0
      12'hA08: dout <= 8'b00111000; // 2568 :  56 - 0x38 -- Background 0x41
      12'hA09: dout <= 8'b01111000; // 2569 : 120 - 0x78
      12'hA0A: dout <= 8'b00111000; // 2570 :  56 - 0x38
      12'hA0B: dout <= 8'b00111000; // 2571 :  56 - 0x38
      12'hA0C: dout <= 8'b00111000; // 2572 :  56 - 0x38
      12'hA0D: dout <= 8'b00111000; // 2573 :  56 - 0x38
      12'hA0E: dout <= 8'b00111000; // 2574 :  56 - 0x38
      12'hA0F: dout <= 8'b00000000; // 2575 :   0 - 0x0
      12'hA10: dout <= 8'b01111100; // 2576 : 124 - 0x7c -- Background 0x42
      12'hA11: dout <= 8'b11111110; // 2577 : 254 - 0xfe
      12'hA12: dout <= 8'b11100110; // 2578 : 230 - 0xe6
      12'hA13: dout <= 8'b00011110; // 2579 :  30 - 0x1e
      12'hA14: dout <= 8'b01111100; // 2580 : 124 - 0x7c
      12'hA15: dout <= 8'b11100000; // 2581 : 224 - 0xe0
      12'hA16: dout <= 8'b11111110; // 2582 : 254 - 0xfe
      12'hA17: dout <= 8'b00000000; // 2583 :   0 - 0x0
      12'hA18: dout <= 8'b01111100; // 2584 : 124 - 0x7c -- Background 0x43
      12'hA19: dout <= 8'b11111100; // 2585 : 252 - 0xfc
      12'hA1A: dout <= 8'b11100110; // 2586 : 230 - 0xe6
      12'hA1B: dout <= 8'b00011100; // 2587 :  28 - 0x1c
      12'hA1C: dout <= 8'b01100110; // 2588 : 102 - 0x66
      12'hA1D: dout <= 8'b11101110; // 2589 : 238 - 0xee
      12'hA1E: dout <= 8'b11111100; // 2590 : 252 - 0xfc
      12'hA1F: dout <= 8'b00000000; // 2591 :   0 - 0x0
      12'hA20: dout <= 8'b00001100; // 2592 :  12 - 0xc -- Background 0x44
      12'hA21: dout <= 8'b00011100; // 2593 :  28 - 0x1c
      12'hA22: dout <= 8'b00111100; // 2594 :  60 - 0x3c
      12'hA23: dout <= 8'b01111100; // 2595 : 124 - 0x7c
      12'hA24: dout <= 8'b11101100; // 2596 : 236 - 0xec
      12'hA25: dout <= 8'b11111110; // 2597 : 254 - 0xfe
      12'hA26: dout <= 8'b00001100; // 2598 :  12 - 0xc
      12'hA27: dout <= 8'b00000000; // 2599 :   0 - 0x0
      12'hA28: dout <= 8'b11111110; // 2600 : 254 - 0xfe -- Background 0x45
      12'hA29: dout <= 8'b11111110; // 2601 : 254 - 0xfe
      12'hA2A: dout <= 8'b11100000; // 2602 : 224 - 0xe0
      12'hA2B: dout <= 8'b11111110; // 2603 : 254 - 0xfe
      12'hA2C: dout <= 8'b00000110; // 2604 :   6 - 0x6
      12'hA2D: dout <= 8'b11101110; // 2605 : 238 - 0xee
      12'hA2E: dout <= 8'b11111100; // 2606 : 252 - 0xfc
      12'hA2F: dout <= 8'b00000000; // 2607 :   0 - 0x0
      12'hA30: dout <= 8'b00111100; // 2608 :  60 - 0x3c -- Background 0x46
      12'hA31: dout <= 8'b01111100; // 2609 : 124 - 0x7c
      12'hA32: dout <= 8'b11100000; // 2610 : 224 - 0xe0
      12'hA33: dout <= 8'b11111110; // 2611 : 254 - 0xfe
      12'hA34: dout <= 8'b11100110; // 2612 : 230 - 0xe6
      12'hA35: dout <= 8'b11101110; // 2613 : 238 - 0xee
      12'hA36: dout <= 8'b00111100; // 2614 :  60 - 0x3c
      12'hA37: dout <= 8'b00000000; // 2615 :   0 - 0x0
      12'hA38: dout <= 8'b11111110; // 2616 : 254 - 0xfe -- Background 0x47
      12'hA39: dout <= 8'b11111100; // 2617 : 252 - 0xfc
      12'hA3A: dout <= 8'b00001100; // 2618 :  12 - 0xc
      12'hA3B: dout <= 8'b00111000; // 2619 :  56 - 0x38
      12'hA3C: dout <= 8'b00111000; // 2620 :  56 - 0x38
      12'hA3D: dout <= 8'b01110000; // 2621 : 112 - 0x70
      12'hA3E: dout <= 8'b01110000; // 2622 : 112 - 0x70
      12'hA3F: dout <= 8'b00000000; // 2623 :   0 - 0x0
      12'hA40: dout <= 8'b00111110; // 2624 :  62 - 0x3e -- Background 0x48
      12'hA41: dout <= 8'b01111100; // 2625 : 124 - 0x7c
      12'hA42: dout <= 8'b11100110; // 2626 : 230 - 0xe6
      12'hA43: dout <= 8'b10111100; // 2627 : 188 - 0xbc
      12'hA44: dout <= 8'b11100110; // 2628 : 230 - 0xe6
      12'hA45: dout <= 8'b11101110; // 2629 : 238 - 0xee
      12'hA46: dout <= 8'b00111100; // 2630 :  60 - 0x3c
      12'hA47: dout <= 8'b00000000; // 2631 :   0 - 0x0
      12'hA48: dout <= 8'b00111100; // 2632 :  60 - 0x3c -- Background 0x49
      12'hA49: dout <= 8'b01111100; // 2633 : 124 - 0x7c
      12'hA4A: dout <= 8'b11100110; // 2634 : 230 - 0xe6
      12'hA4B: dout <= 8'b11101110; // 2635 : 238 - 0xee
      12'hA4C: dout <= 8'b11111110; // 2636 : 254 - 0xfe
      12'hA4D: dout <= 8'b10000110; // 2637 : 134 - 0x86
      12'hA4E: dout <= 8'b01111100; // 2638 : 124 - 0x7c
      12'hA4F: dout <= 8'b01000000; // 2639 :  64 - 0x40
      12'hA50: dout <= 8'b11101110; // 2640 : 238 - 0xee -- Background 0x4a
      12'hA51: dout <= 8'b11101110; // 2641 : 238 - 0xee
      12'hA52: dout <= 8'b11101110; // 2642 : 238 - 0xee
      12'hA53: dout <= 8'b11101110; // 2643 : 238 - 0xee
      12'hA54: dout <= 8'b11101110; // 2644 : 238 - 0xee
      12'hA55: dout <= 8'b11101110; // 2645 : 238 - 0xee
      12'hA56: dout <= 8'b11101110; // 2646 : 238 - 0xee
      12'hA57: dout <= 8'b10001000; // 2647 : 136 - 0x88
      12'hA58: dout <= 8'b11100000; // 2648 : 224 - 0xe0 -- Background 0x4b
      12'hA59: dout <= 8'b11100000; // 2649 : 224 - 0xe0
      12'hA5A: dout <= 8'b11100000; // 2650 : 224 - 0xe0
      12'hA5B: dout <= 8'b11100000; // 2651 : 224 - 0xe0
      12'hA5C: dout <= 8'b11100000; // 2652 : 224 - 0xe0
      12'hA5D: dout <= 8'b11100000; // 2653 : 224 - 0xe0
      12'hA5E: dout <= 8'b11100000; // 2654 : 224 - 0xe0
      12'hA5F: dout <= 8'b10000000; // 2655 : 128 - 0x80
      12'hA60: dout <= 8'b00000000; // 2656 :   0 - 0x0 -- Background 0x4c
      12'hA61: dout <= 8'b01111111; // 2657 : 127 - 0x7f
      12'hA62: dout <= 8'b01111111; // 2658 : 127 - 0x7f
      12'hA63: dout <= 8'b01111111; // 2659 : 127 - 0x7f
      12'hA64: dout <= 8'b01111111; // 2660 : 127 - 0x7f
      12'hA65: dout <= 8'b01111111; // 2661 : 127 - 0x7f
      12'hA66: dout <= 8'b01111111; // 2662 : 127 - 0x7f
      12'hA67: dout <= 8'b01111111; // 2663 : 127 - 0x7f
      12'hA68: dout <= 8'b01111111; // 2664 : 127 - 0x7f -- Background 0x4d
      12'hA69: dout <= 8'b01111111; // 2665 : 127 - 0x7f
      12'hA6A: dout <= 8'b01111111; // 2666 : 127 - 0x7f
      12'hA6B: dout <= 8'b01111111; // 2667 : 127 - 0x7f
      12'hA6C: dout <= 8'b01111111; // 2668 : 127 - 0x7f
      12'hA6D: dout <= 8'b01111111; // 2669 : 127 - 0x7f
      12'hA6E: dout <= 8'b01111111; // 2670 : 127 - 0x7f
      12'hA6F: dout <= 8'b00000000; // 2671 :   0 - 0x0
      12'hA70: dout <= 8'b00000000; // 2672 :   0 - 0x0 -- Background 0x4e
      12'hA71: dout <= 8'b11111110; // 2673 : 254 - 0xfe
      12'hA72: dout <= 8'b11111110; // 2674 : 254 - 0xfe
      12'hA73: dout <= 8'b11111110; // 2675 : 254 - 0xfe
      12'hA74: dout <= 8'b11111110; // 2676 : 254 - 0xfe
      12'hA75: dout <= 8'b11111110; // 2677 : 254 - 0xfe
      12'hA76: dout <= 8'b11111110; // 2678 : 254 - 0xfe
      12'hA77: dout <= 8'b11111110; // 2679 : 254 - 0xfe
      12'hA78: dout <= 8'b11111110; // 2680 : 254 - 0xfe -- Background 0x4f
      12'hA79: dout <= 8'b11111110; // 2681 : 254 - 0xfe
      12'hA7A: dout <= 8'b11111110; // 2682 : 254 - 0xfe
      12'hA7B: dout <= 8'b11111110; // 2683 : 254 - 0xfe
      12'hA7C: dout <= 8'b11111110; // 2684 : 254 - 0xfe
      12'hA7D: dout <= 8'b11111110; // 2685 : 254 - 0xfe
      12'hA7E: dout <= 8'b11111110; // 2686 : 254 - 0xfe
      12'hA7F: dout <= 8'b00000000; // 2687 :   0 - 0x0
      12'hA80: dout <= 8'b00000000; // 2688 :   0 - 0x0 -- Background 0x50
      12'hA81: dout <= 8'b00000000; // 2689 :   0 - 0x0
      12'hA82: dout <= 8'b00000000; // 2690 :   0 - 0x0
      12'hA83: dout <= 8'b00000000; // 2691 :   0 - 0x0
      12'hA84: dout <= 8'b00000000; // 2692 :   0 - 0x0
      12'hA85: dout <= 8'b00000000; // 2693 :   0 - 0x0
      12'hA86: dout <= 8'b00000000; // 2694 :   0 - 0x0
      12'hA87: dout <= 8'b00000000; // 2695 :   0 - 0x0
      12'hA88: dout <= 8'b00000000; // 2696 :   0 - 0x0 -- Background 0x51
      12'hA89: dout <= 8'b00010000; // 2697 :  16 - 0x10
      12'hA8A: dout <= 8'b00010000; // 2698 :  16 - 0x10
      12'hA8B: dout <= 8'b01111100; // 2699 : 124 - 0x7c
      12'hA8C: dout <= 8'b00111000; // 2700 :  56 - 0x38
      12'hA8D: dout <= 8'b00111000; // 2701 :  56 - 0x38
      12'hA8E: dout <= 8'b01101100; // 2702 : 108 - 0x6c
      12'hA8F: dout <= 8'b00000000; // 2703 :   0 - 0x0
      12'hA90: dout <= 8'b00000000; // 2704 :   0 - 0x0 -- Background 0x52
      12'hA91: dout <= 8'b00010000; // 2705 :  16 - 0x10
      12'hA92: dout <= 8'b00010000; // 2706 :  16 - 0x10
      12'hA93: dout <= 8'b01111100; // 2707 : 124 - 0x7c
      12'hA94: dout <= 8'b00111000; // 2708 :  56 - 0x38
      12'hA95: dout <= 8'b00111000; // 2709 :  56 - 0x38
      12'hA96: dout <= 8'b01101100; // 2710 : 108 - 0x6c
      12'hA97: dout <= 8'b00000000; // 2711 :   0 - 0x0
      12'hA98: dout <= 8'b00000000; // 2712 :   0 - 0x0 -- Background 0x53
      12'hA99: dout <= 8'b00000000; // 2713 :   0 - 0x0
      12'hA9A: dout <= 8'b00000000; // 2714 :   0 - 0x0
      12'hA9B: dout <= 8'b00000000; // 2715 :   0 - 0x0
      12'hA9C: dout <= 8'b00000000; // 2716 :   0 - 0x0
      12'hA9D: dout <= 8'b00000000; // 2717 :   0 - 0x0
      12'hA9E: dout <= 8'b00000000; // 2718 :   0 - 0x0
      12'hA9F: dout <= 8'b00000000; // 2719 :   0 - 0x0
      12'hAA0: dout <= 8'b11111111; // 2720 : 255 - 0xff -- Background 0x54
      12'hAA1: dout <= 8'b11111111; // 2721 : 255 - 0xff
      12'hAA2: dout <= 8'b11111111; // 2722 : 255 - 0xff
      12'hAA3: dout <= 8'b11111111; // 2723 : 255 - 0xff
      12'hAA4: dout <= 8'b11111111; // 2724 : 255 - 0xff
      12'hAA5: dout <= 8'b11111111; // 2725 : 255 - 0xff
      12'hAA6: dout <= 8'b11111111; // 2726 : 255 - 0xff
      12'hAA7: dout <= 8'b11111111; // 2727 : 255 - 0xff
      12'hAA8: dout <= 8'b11111111; // 2728 : 255 - 0xff -- Background 0x55
      12'hAA9: dout <= 8'b11111111; // 2729 : 255 - 0xff
      12'hAAA: dout <= 8'b11111111; // 2730 : 255 - 0xff
      12'hAAB: dout <= 8'b11111111; // 2731 : 255 - 0xff
      12'hAAC: dout <= 8'b11111111; // 2732 : 255 - 0xff
      12'hAAD: dout <= 8'b11111111; // 2733 : 255 - 0xff
      12'hAAE: dout <= 8'b11111111; // 2734 : 255 - 0xff
      12'hAAF: dout <= 8'b11111111; // 2735 : 255 - 0xff
      12'hAB0: dout <= 8'b00000010; // 2736 :   2 - 0x2 -- Background 0x56
      12'hAB1: dout <= 8'b00000101; // 2737 :   5 - 0x5
      12'hAB2: dout <= 8'b10101010; // 2738 : 170 - 0xaa
      12'hAB3: dout <= 8'b01010001; // 2739 :  81 - 0x51
      12'hAB4: dout <= 8'b10101010; // 2740 : 170 - 0xaa
      12'hAB5: dout <= 8'b01010001; // 2741 :  81 - 0x51
      12'hAB6: dout <= 8'b10100010; // 2742 : 162 - 0xa2
      12'hAB7: dout <= 8'b00000100; // 2743 :   4 - 0x4
      12'hAB8: dout <= 8'b00001000; // 2744 :   8 - 0x8 -- Background 0x57
      12'hAB9: dout <= 8'b01010101; // 2745 :  85 - 0x55
      12'hABA: dout <= 8'b00101010; // 2746 :  42 - 0x2a
      12'hABB: dout <= 8'b01010101; // 2747 :  85 - 0x55
      12'hABC: dout <= 8'b00101010; // 2748 :  42 - 0x2a
      12'hABD: dout <= 8'b01000101; // 2749 :  69 - 0x45
      12'hABE: dout <= 8'b00001010; // 2750 :  10 - 0xa
      12'hABF: dout <= 8'b00010000; // 2751 :  16 - 0x10
      12'hAC0: dout <= 8'b00000000; // 2752 :   0 - 0x0 -- Background 0x58
      12'hAC1: dout <= 8'b00111111; // 2753 :  63 - 0x3f
      12'hAC2: dout <= 8'b01011111; // 2754 :  95 - 0x5f
      12'hAC3: dout <= 8'b01101111; // 2755 : 111 - 0x6f
      12'hAC4: dout <= 8'b01110000; // 2756 : 112 - 0x70
      12'hAC5: dout <= 8'b01110111; // 2757 : 119 - 0x77
      12'hAC6: dout <= 8'b01110111; // 2758 : 119 - 0x77
      12'hAC7: dout <= 8'b01110111; // 2759 : 119 - 0x77
      12'hAC8: dout <= 8'b01110111; // 2760 : 119 - 0x77 -- Background 0x59
      12'hAC9: dout <= 8'b01110111; // 2761 : 119 - 0x77
      12'hACA: dout <= 8'b01110111; // 2762 : 119 - 0x77
      12'hACB: dout <= 8'b01110000; // 2763 : 112 - 0x70
      12'hACC: dout <= 8'b01101111; // 2764 : 111 - 0x6f
      12'hACD: dout <= 8'b01011111; // 2765 :  95 - 0x5f
      12'hACE: dout <= 8'b00010101; // 2766 :  21 - 0x15
      12'hACF: dout <= 8'b00000000; // 2767 :   0 - 0x0
      12'hAD0: dout <= 8'b00000000; // 2768 :   0 - 0x0 -- Background 0x5a
      12'hAD1: dout <= 8'b11111100; // 2769 : 252 - 0xfc
      12'hAD2: dout <= 8'b11111000; // 2770 : 248 - 0xf8
      12'hAD3: dout <= 8'b11110110; // 2771 : 246 - 0xf6
      12'hAD4: dout <= 8'b00001100; // 2772 :  12 - 0xc
      12'hAD5: dout <= 8'b11101110; // 2773 : 238 - 0xee
      12'hAD6: dout <= 8'b11101100; // 2774 : 236 - 0xec
      12'hAD7: dout <= 8'b11101110; // 2775 : 238 - 0xee
      12'hAD8: dout <= 8'b11101100; // 2776 : 236 - 0xec -- Background 0x5b
      12'hAD9: dout <= 8'b11101110; // 2777 : 238 - 0xee
      12'hADA: dout <= 8'b11101100; // 2778 : 236 - 0xec
      12'hADB: dout <= 8'b00001110; // 2779 :  14 - 0xe
      12'hADC: dout <= 8'b11110100; // 2780 : 244 - 0xf4
      12'hADD: dout <= 8'b11111010; // 2781 : 250 - 0xfa
      12'hADE: dout <= 8'b01010100; // 2782 :  84 - 0x54
      12'hADF: dout <= 8'b00000000; // 2783 :   0 - 0x0
      12'hAE0: dout <= 8'b00000000; // 2784 :   0 - 0x0 -- Background 0x5c
      12'hAE1: dout <= 8'b00011100; // 2785 :  28 - 0x1c
      12'hAE2: dout <= 8'b00111110; // 2786 :  62 - 0x3e
      12'hAE3: dout <= 8'b00111110; // 2787 :  62 - 0x3e
      12'hAE4: dout <= 8'b00111110; // 2788 :  62 - 0x3e
      12'hAE5: dout <= 8'b00011100; // 2789 :  28 - 0x1c
      12'hAE6: dout <= 8'b00011100; // 2790 :  28 - 0x1c
      12'hAE7: dout <= 8'b00000000; // 2791 :   0 - 0x0
      12'hAE8: dout <= 8'b00000000; // 2792 :   0 - 0x0 -- Background 0x5d
      12'hAE9: dout <= 8'b00000000; // 2793 :   0 - 0x0
      12'hAEA: dout <= 8'b00000000; // 2794 :   0 - 0x0
      12'hAEB: dout <= 8'b00000000; // 2795 :   0 - 0x0
      12'hAEC: dout <= 8'b00000000; // 2796 :   0 - 0x0
      12'hAED: dout <= 8'b00000000; // 2797 :   0 - 0x0
      12'hAEE: dout <= 8'b00000000; // 2798 :   0 - 0x0
      12'hAEF: dout <= 8'b00000000; // 2799 :   0 - 0x0
      12'hAF0: dout <= 8'b00000000; // 2800 :   0 - 0x0 -- Background 0x5e
      12'hAF1: dout <= 8'b00010100; // 2801 :  20 - 0x14
      12'hAF2: dout <= 8'b00110110; // 2802 :  54 - 0x36
      12'hAF3: dout <= 8'b00111110; // 2803 :  62 - 0x3e
      12'hAF4: dout <= 8'b00111110; // 2804 :  62 - 0x3e
      12'hAF5: dout <= 8'b00011100; // 2805 :  28 - 0x1c
      12'hAF6: dout <= 8'b00001000; // 2806 :   8 - 0x8
      12'hAF7: dout <= 8'b00000000; // 2807 :   0 - 0x0
      12'hAF8: dout <= 8'b00000000; // 2808 :   0 - 0x0 -- Background 0x5f
      12'hAF9: dout <= 8'b00010100; // 2809 :  20 - 0x14
      12'hAFA: dout <= 8'b00011100; // 2810 :  28 - 0x1c
      12'hAFB: dout <= 8'b00011100; // 2811 :  28 - 0x1c
      12'hAFC: dout <= 8'b00011100; // 2812 :  28 - 0x1c
      12'hAFD: dout <= 8'b00011100; // 2813 :  28 - 0x1c
      12'hAFE: dout <= 8'b00011100; // 2814 :  28 - 0x1c
      12'hAFF: dout <= 8'b00000000; // 2815 :   0 - 0x0
      12'hB00: dout <= 8'b00000000; // 2816 :   0 - 0x0 -- Background 0x60
      12'hB01: dout <= 8'b01111111; // 2817 : 127 - 0x7f
      12'hB02: dout <= 8'b01111111; // 2818 : 127 - 0x7f
      12'hB03: dout <= 8'b01111111; // 2819 : 127 - 0x7f
      12'hB04: dout <= 8'b01111111; // 2820 : 127 - 0x7f
      12'hB05: dout <= 8'b01111111; // 2821 : 127 - 0x7f
      12'hB06: dout <= 8'b00101010; // 2822 :  42 - 0x2a
      12'hB07: dout <= 8'b00000000; // 2823 :   0 - 0x0
      12'hB08: dout <= 8'b00000000; // 2824 :   0 - 0x0 -- Background 0x61
      12'hB09: dout <= 8'b11111111; // 2825 : 255 - 0xff
      12'hB0A: dout <= 8'b11111111; // 2826 : 255 - 0xff
      12'hB0B: dout <= 8'b11111111; // 2827 : 255 - 0xff
      12'hB0C: dout <= 8'b11111111; // 2828 : 255 - 0xff
      12'hB0D: dout <= 8'b11111111; // 2829 : 255 - 0xff
      12'hB0E: dout <= 8'b10101010; // 2830 : 170 - 0xaa
      12'hB0F: dout <= 8'b00000000; // 2831 :   0 - 0x0
      12'hB10: dout <= 8'b00000000; // 2832 :   0 - 0x0 -- Background 0x62
      12'hB11: dout <= 8'b11111110; // 2833 : 254 - 0xfe
      12'hB12: dout <= 8'b11111110; // 2834 : 254 - 0xfe
      12'hB13: dout <= 8'b11111110; // 2835 : 254 - 0xfe
      12'hB14: dout <= 8'b11111110; // 2836 : 254 - 0xfe
      12'hB15: dout <= 8'b11111110; // 2837 : 254 - 0xfe
      12'hB16: dout <= 8'b10101010; // 2838 : 170 - 0xaa
      12'hB17: dout <= 8'b00000000; // 2839 :   0 - 0x0
      12'hB18: dout <= 8'b00000000; // 2840 :   0 - 0x0 -- Background 0x63
      12'hB19: dout <= 8'b00000000; // 2841 :   0 - 0x0
      12'hB1A: dout <= 8'b00000000; // 2842 :   0 - 0x0
      12'hB1B: dout <= 8'b00000000; // 2843 :   0 - 0x0
      12'hB1C: dout <= 8'b00000000; // 2844 :   0 - 0x0
      12'hB1D: dout <= 8'b00000000; // 2845 :   0 - 0x0
      12'hB1E: dout <= 8'b00000000; // 2846 :   0 - 0x0
      12'hB1F: dout <= 8'b00000000; // 2847 :   0 - 0x0
      12'hB20: dout <= 8'b00000000; // 2848 :   0 - 0x0 -- Background 0x64
      12'hB21: dout <= 8'b00000000; // 2849 :   0 - 0x0
      12'hB22: dout <= 8'b00000001; // 2850 :   1 - 0x1
      12'hB23: dout <= 8'b00000001; // 2851 :   1 - 0x1
      12'hB24: dout <= 8'b00000011; // 2852 :   3 - 0x3
      12'hB25: dout <= 8'b00000011; // 2853 :   3 - 0x3
      12'hB26: dout <= 8'b00000111; // 2854 :   7 - 0x7
      12'hB27: dout <= 8'b00000111; // 2855 :   7 - 0x7
      12'hB28: dout <= 8'b00001111; // 2856 :  15 - 0xf -- Background 0x65
      12'hB29: dout <= 8'b00001111; // 2857 :  15 - 0xf
      12'hB2A: dout <= 8'b00011111; // 2858 :  31 - 0x1f
      12'hB2B: dout <= 8'b00011111; // 2859 :  31 - 0x1f
      12'hB2C: dout <= 8'b00111111; // 2860 :  63 - 0x3f
      12'hB2D: dout <= 8'b00111111; // 2861 :  63 - 0x3f
      12'hB2E: dout <= 8'b01010101; // 2862 :  85 - 0x55
      12'hB2F: dout <= 8'b00000000; // 2863 :   0 - 0x0
      12'hB30: dout <= 8'b00000000; // 2864 :   0 - 0x0 -- Background 0x66
      12'hB31: dout <= 8'b00000000; // 2865 :   0 - 0x0
      12'hB32: dout <= 8'b00000000; // 2866 :   0 - 0x0
      12'hB33: dout <= 8'b10000000; // 2867 : 128 - 0x80
      12'hB34: dout <= 8'b01000000; // 2868 :  64 - 0x40
      12'hB35: dout <= 8'b10000000; // 2869 : 128 - 0x80
      12'hB36: dout <= 8'b11000000; // 2870 : 192 - 0xc0
      12'hB37: dout <= 8'b11100000; // 2871 : 224 - 0xe0
      12'hB38: dout <= 8'b11010000; // 2872 : 208 - 0xd0 -- Background 0x67
      12'hB39: dout <= 8'b11100000; // 2873 : 224 - 0xe0
      12'hB3A: dout <= 8'b11110000; // 2874 : 240 - 0xf0
      12'hB3B: dout <= 8'b11101000; // 2875 : 232 - 0xe8
      12'hB3C: dout <= 8'b11110100; // 2876 : 244 - 0xf4
      12'hB3D: dout <= 8'b11111000; // 2877 : 248 - 0xf8
      12'hB3E: dout <= 8'b01010100; // 2878 :  84 - 0x54
      12'hB3F: dout <= 8'b00000000; // 2879 :   0 - 0x0
      12'hB40: dout <= 8'b00000000; // 2880 :   0 - 0x0 -- Background 0x68
      12'hB41: dout <= 8'b00000000; // 2881 :   0 - 0x0
      12'hB42: dout <= 8'b00000000; // 2882 :   0 - 0x0
      12'hB43: dout <= 8'b00000000; // 2883 :   0 - 0x0
      12'hB44: dout <= 8'b00000000; // 2884 :   0 - 0x0
      12'hB45: dout <= 8'b00000000; // 2885 :   0 - 0x0
      12'hB46: dout <= 8'b00000000; // 2886 :   0 - 0x0
      12'hB47: dout <= 8'b00000000; // 2887 :   0 - 0x0
      12'hB48: dout <= 8'b00000000; // 2888 :   0 - 0x0 -- Background 0x69
      12'hB49: dout <= 8'b00000000; // 2889 :   0 - 0x0
      12'hB4A: dout <= 8'b00000000; // 2890 :   0 - 0x0
      12'hB4B: dout <= 8'b00000000; // 2891 :   0 - 0x0
      12'hB4C: dout <= 8'b00000000; // 2892 :   0 - 0x0
      12'hB4D: dout <= 8'b00000000; // 2893 :   0 - 0x0
      12'hB4E: dout <= 8'b00000000; // 2894 :   0 - 0x0
      12'hB4F: dout <= 8'b00000000; // 2895 :   0 - 0x0
      12'hB50: dout <= 8'b00000000; // 2896 :   0 - 0x0 -- Background 0x6a
      12'hB51: dout <= 8'b00000000; // 2897 :   0 - 0x0
      12'hB52: dout <= 8'b00000000; // 2898 :   0 - 0x0
      12'hB53: dout <= 8'b00000000; // 2899 :   0 - 0x0
      12'hB54: dout <= 8'b00000000; // 2900 :   0 - 0x0
      12'hB55: dout <= 8'b00000000; // 2901 :   0 - 0x0
      12'hB56: dout <= 8'b00000000; // 2902 :   0 - 0x0
      12'hB57: dout <= 8'b00000000; // 2903 :   0 - 0x0
      12'hB58: dout <= 8'b00000000; // 2904 :   0 - 0x0 -- Background 0x6b
      12'hB59: dout <= 8'b00000000; // 2905 :   0 - 0x0
      12'hB5A: dout <= 8'b00000000; // 2906 :   0 - 0x0
      12'hB5B: dout <= 8'b00000000; // 2907 :   0 - 0x0
      12'hB5C: dout <= 8'b00000000; // 2908 :   0 - 0x0
      12'hB5D: dout <= 8'b00000000; // 2909 :   0 - 0x0
      12'hB5E: dout <= 8'b00000000; // 2910 :   0 - 0x0
      12'hB5F: dout <= 8'b00000000; // 2911 :   0 - 0x0
      12'hB60: dout <= 8'b00000000; // 2912 :   0 - 0x0 -- Background 0x6c
      12'hB61: dout <= 8'b00000000; // 2913 :   0 - 0x0
      12'hB62: dout <= 8'b00000000; // 2914 :   0 - 0x0
      12'hB63: dout <= 8'b00000000; // 2915 :   0 - 0x0
      12'hB64: dout <= 8'b00000000; // 2916 :   0 - 0x0
      12'hB65: dout <= 8'b00000000; // 2917 :   0 - 0x0
      12'hB66: dout <= 8'b00000000; // 2918 :   0 - 0x0
      12'hB67: dout <= 8'b00000000; // 2919 :   0 - 0x0
      12'hB68: dout <= 8'b00000000; // 2920 :   0 - 0x0 -- Background 0x6d
      12'hB69: dout <= 8'b00000000; // 2921 :   0 - 0x0
      12'hB6A: dout <= 8'b00000000; // 2922 :   0 - 0x0
      12'hB6B: dout <= 8'b00000000; // 2923 :   0 - 0x0
      12'hB6C: dout <= 8'b00000000; // 2924 :   0 - 0x0
      12'hB6D: dout <= 8'b00000000; // 2925 :   0 - 0x0
      12'hB6E: dout <= 8'b00000000; // 2926 :   0 - 0x0
      12'hB6F: dout <= 8'b00000000; // 2927 :   0 - 0x0
      12'hB70: dout <= 8'b00000000; // 2928 :   0 - 0x0 -- Background 0x6e
      12'hB71: dout <= 8'b00000000; // 2929 :   0 - 0x0
      12'hB72: dout <= 8'b00000000; // 2930 :   0 - 0x0
      12'hB73: dout <= 8'b00000000; // 2931 :   0 - 0x0
      12'hB74: dout <= 8'b00000000; // 2932 :   0 - 0x0
      12'hB75: dout <= 8'b00000000; // 2933 :   0 - 0x0
      12'hB76: dout <= 8'b00000000; // 2934 :   0 - 0x0
      12'hB77: dout <= 8'b00000000; // 2935 :   0 - 0x0
      12'hB78: dout <= 8'b00000000; // 2936 :   0 - 0x0 -- Background 0x6f
      12'hB79: dout <= 8'b00000000; // 2937 :   0 - 0x0
      12'hB7A: dout <= 8'b00000000; // 2938 :   0 - 0x0
      12'hB7B: dout <= 8'b00000000; // 2939 :   0 - 0x0
      12'hB7C: dout <= 8'b00000000; // 2940 :   0 - 0x0
      12'hB7D: dout <= 8'b00000000; // 2941 :   0 - 0x0
      12'hB7E: dout <= 8'b00000000; // 2942 :   0 - 0x0
      12'hB7F: dout <= 8'b00000000; // 2943 :   0 - 0x0
      12'hB80: dout <= 8'b00000000; // 2944 :   0 - 0x0 -- Background 0x70
      12'hB81: dout <= 8'b00000000; // 2945 :   0 - 0x0
      12'hB82: dout <= 8'b00000000; // 2946 :   0 - 0x0
      12'hB83: dout <= 8'b00000000; // 2947 :   0 - 0x0
      12'hB84: dout <= 8'b00000000; // 2948 :   0 - 0x0
      12'hB85: dout <= 8'b00000000; // 2949 :   0 - 0x0
      12'hB86: dout <= 8'b00000000; // 2950 :   0 - 0x0
      12'hB87: dout <= 8'b00000000; // 2951 :   0 - 0x0
      12'hB88: dout <= 8'b00000000; // 2952 :   0 - 0x0 -- Background 0x71
      12'hB89: dout <= 8'b00000000; // 2953 :   0 - 0x0
      12'hB8A: dout <= 8'b00000000; // 2954 :   0 - 0x0
      12'hB8B: dout <= 8'b00000000; // 2955 :   0 - 0x0
      12'hB8C: dout <= 8'b00000000; // 2956 :   0 - 0x0
      12'hB8D: dout <= 8'b00000000; // 2957 :   0 - 0x0
      12'hB8E: dout <= 8'b00000000; // 2958 :   0 - 0x0
      12'hB8F: dout <= 8'b00000000; // 2959 :   0 - 0x0
      12'hB90: dout <= 8'b00000000; // 2960 :   0 - 0x0 -- Background 0x72
      12'hB91: dout <= 8'b00000000; // 2961 :   0 - 0x0
      12'hB92: dout <= 8'b00000000; // 2962 :   0 - 0x0
      12'hB93: dout <= 8'b00000000; // 2963 :   0 - 0x0
      12'hB94: dout <= 8'b00000000; // 2964 :   0 - 0x0
      12'hB95: dout <= 8'b00000000; // 2965 :   0 - 0x0
      12'hB96: dout <= 8'b00000000; // 2966 :   0 - 0x0
      12'hB97: dout <= 8'b00000000; // 2967 :   0 - 0x0
      12'hB98: dout <= 8'b00000000; // 2968 :   0 - 0x0 -- Background 0x73
      12'hB99: dout <= 8'b00000000; // 2969 :   0 - 0x0
      12'hB9A: dout <= 8'b00000000; // 2970 :   0 - 0x0
      12'hB9B: dout <= 8'b00000000; // 2971 :   0 - 0x0
      12'hB9C: dout <= 8'b00000000; // 2972 :   0 - 0x0
      12'hB9D: dout <= 8'b00000000; // 2973 :   0 - 0x0
      12'hB9E: dout <= 8'b00000000; // 2974 :   0 - 0x0
      12'hB9F: dout <= 8'b00000000; // 2975 :   0 - 0x0
      12'hBA0: dout <= 8'b00000000; // 2976 :   0 - 0x0 -- Background 0x74
      12'hBA1: dout <= 8'b00000000; // 2977 :   0 - 0x0
      12'hBA2: dout <= 8'b00000000; // 2978 :   0 - 0x0
      12'hBA3: dout <= 8'b00000000; // 2979 :   0 - 0x0
      12'hBA4: dout <= 8'b00000000; // 2980 :   0 - 0x0
      12'hBA5: dout <= 8'b00000000; // 2981 :   0 - 0x0
      12'hBA6: dout <= 8'b00000000; // 2982 :   0 - 0x0
      12'hBA7: dout <= 8'b00000000; // 2983 :   0 - 0x0
      12'hBA8: dout <= 8'b00000000; // 2984 :   0 - 0x0 -- Background 0x75
      12'hBA9: dout <= 8'b00000000; // 2985 :   0 - 0x0
      12'hBAA: dout <= 8'b00000000; // 2986 :   0 - 0x0
      12'hBAB: dout <= 8'b00000000; // 2987 :   0 - 0x0
      12'hBAC: dout <= 8'b00000000; // 2988 :   0 - 0x0
      12'hBAD: dout <= 8'b00000000; // 2989 :   0 - 0x0
      12'hBAE: dout <= 8'b00000000; // 2990 :   0 - 0x0
      12'hBAF: dout <= 8'b00000000; // 2991 :   0 - 0x0
      12'hBB0: dout <= 8'b00000000; // 2992 :   0 - 0x0 -- Background 0x76
      12'hBB1: dout <= 8'b00000000; // 2993 :   0 - 0x0
      12'hBB2: dout <= 8'b00000000; // 2994 :   0 - 0x0
      12'hBB3: dout <= 8'b00000000; // 2995 :   0 - 0x0
      12'hBB4: dout <= 8'b00000000; // 2996 :   0 - 0x0
      12'hBB5: dout <= 8'b00000000; // 2997 :   0 - 0x0
      12'hBB6: dout <= 8'b00000000; // 2998 :   0 - 0x0
      12'hBB7: dout <= 8'b00000000; // 2999 :   0 - 0x0
      12'hBB8: dout <= 8'b00000000; // 3000 :   0 - 0x0 -- Background 0x77
      12'hBB9: dout <= 8'b00000000; // 3001 :   0 - 0x0
      12'hBBA: dout <= 8'b00000000; // 3002 :   0 - 0x0
      12'hBBB: dout <= 8'b00000000; // 3003 :   0 - 0x0
      12'hBBC: dout <= 8'b00000000; // 3004 :   0 - 0x0
      12'hBBD: dout <= 8'b00000000; // 3005 :   0 - 0x0
      12'hBBE: dout <= 8'b00000000; // 3006 :   0 - 0x0
      12'hBBF: dout <= 8'b00000000; // 3007 :   0 - 0x0
      12'hBC0: dout <= 8'b00000000; // 3008 :   0 - 0x0 -- Background 0x78
      12'hBC1: dout <= 8'b00000000; // 3009 :   0 - 0x0
      12'hBC2: dout <= 8'b00000000; // 3010 :   0 - 0x0
      12'hBC3: dout <= 8'b00000000; // 3011 :   0 - 0x0
      12'hBC4: dout <= 8'b00000000; // 3012 :   0 - 0x0
      12'hBC5: dout <= 8'b00000000; // 3013 :   0 - 0x0
      12'hBC6: dout <= 8'b00000000; // 3014 :   0 - 0x0
      12'hBC7: dout <= 8'b00000000; // 3015 :   0 - 0x0
      12'hBC8: dout <= 8'b00000000; // 3016 :   0 - 0x0 -- Background 0x79
      12'hBC9: dout <= 8'b00000000; // 3017 :   0 - 0x0
      12'hBCA: dout <= 8'b00000000; // 3018 :   0 - 0x0
      12'hBCB: dout <= 8'b00000000; // 3019 :   0 - 0x0
      12'hBCC: dout <= 8'b00000000; // 3020 :   0 - 0x0
      12'hBCD: dout <= 8'b00000000; // 3021 :   0 - 0x0
      12'hBCE: dout <= 8'b00000000; // 3022 :   0 - 0x0
      12'hBCF: dout <= 8'b00000000; // 3023 :   0 - 0x0
      12'hBD0: dout <= 8'b00000000; // 3024 :   0 - 0x0 -- Background 0x7a
      12'hBD1: dout <= 8'b00000000; // 3025 :   0 - 0x0
      12'hBD2: dout <= 8'b00000000; // 3026 :   0 - 0x0
      12'hBD3: dout <= 8'b00000000; // 3027 :   0 - 0x0
      12'hBD4: dout <= 8'b00000000; // 3028 :   0 - 0x0
      12'hBD5: dout <= 8'b00000000; // 3029 :   0 - 0x0
      12'hBD6: dout <= 8'b00000000; // 3030 :   0 - 0x0
      12'hBD7: dout <= 8'b00000000; // 3031 :   0 - 0x0
      12'hBD8: dout <= 8'b00000000; // 3032 :   0 - 0x0 -- Background 0x7b
      12'hBD9: dout <= 8'b00000000; // 3033 :   0 - 0x0
      12'hBDA: dout <= 8'b00000000; // 3034 :   0 - 0x0
      12'hBDB: dout <= 8'b00000000; // 3035 :   0 - 0x0
      12'hBDC: dout <= 8'b00000000; // 3036 :   0 - 0x0
      12'hBDD: dout <= 8'b00000000; // 3037 :   0 - 0x0
      12'hBDE: dout <= 8'b00000000; // 3038 :   0 - 0x0
      12'hBDF: dout <= 8'b00000000; // 3039 :   0 - 0x0
      12'hBE0: dout <= 8'b00000000; // 3040 :   0 - 0x0 -- Background 0x7c
      12'hBE1: dout <= 8'b00000000; // 3041 :   0 - 0x0
      12'hBE2: dout <= 8'b00000000; // 3042 :   0 - 0x0
      12'hBE3: dout <= 8'b00000000; // 3043 :   0 - 0x0
      12'hBE4: dout <= 8'b00000000; // 3044 :   0 - 0x0
      12'hBE5: dout <= 8'b00000000; // 3045 :   0 - 0x0
      12'hBE6: dout <= 8'b00000000; // 3046 :   0 - 0x0
      12'hBE7: dout <= 8'b00000000; // 3047 :   0 - 0x0
      12'hBE8: dout <= 8'b00000000; // 3048 :   0 - 0x0 -- Background 0x7d
      12'hBE9: dout <= 8'b00000000; // 3049 :   0 - 0x0
      12'hBEA: dout <= 8'b00000000; // 3050 :   0 - 0x0
      12'hBEB: dout <= 8'b00000000; // 3051 :   0 - 0x0
      12'hBEC: dout <= 8'b00000000; // 3052 :   0 - 0x0
      12'hBED: dout <= 8'b00000000; // 3053 :   0 - 0x0
      12'hBEE: dout <= 8'b00000000; // 3054 :   0 - 0x0
      12'hBEF: dout <= 8'b00000000; // 3055 :   0 - 0x0
      12'hBF0: dout <= 8'b00000000; // 3056 :   0 - 0x0 -- Background 0x7e
      12'hBF1: dout <= 8'b00000000; // 3057 :   0 - 0x0
      12'hBF2: dout <= 8'b00000000; // 3058 :   0 - 0x0
      12'hBF3: dout <= 8'b00000000; // 3059 :   0 - 0x0
      12'hBF4: dout <= 8'b00000000; // 3060 :   0 - 0x0
      12'hBF5: dout <= 8'b00000000; // 3061 :   0 - 0x0
      12'hBF6: dout <= 8'b00000000; // 3062 :   0 - 0x0
      12'hBF7: dout <= 8'b00000000; // 3063 :   0 - 0x0
      12'hBF8: dout <= 8'b00000000; // 3064 :   0 - 0x0 -- Background 0x7f
      12'hBF9: dout <= 8'b00000000; // 3065 :   0 - 0x0
      12'hBFA: dout <= 8'b00000000; // 3066 :   0 - 0x0
      12'hBFB: dout <= 8'b00000000; // 3067 :   0 - 0x0
      12'hBFC: dout <= 8'b00000000; // 3068 :   0 - 0x0
      12'hBFD: dout <= 8'b00000000; // 3069 :   0 - 0x0
      12'hBFE: dout <= 8'b00000000; // 3070 :   0 - 0x0
      12'hBFF: dout <= 8'b00000000; // 3071 :   0 - 0x0
      12'hC00: dout <= 8'b00000000; // 3072 :   0 - 0x0 -- Background 0x80
      12'hC01: dout <= 8'b00000011; // 3073 :   3 - 0x3
      12'hC02: dout <= 8'b00001111; // 3074 :  15 - 0xf
      12'hC03: dout <= 8'b00011111; // 3075 :  31 - 0x1f
      12'hC04: dout <= 8'b00011111; // 3076 :  31 - 0x1f
      12'hC05: dout <= 8'b00111111; // 3077 :  63 - 0x3f
      12'hC06: dout <= 8'b00111111; // 3078 :  63 - 0x3f
      12'hC07: dout <= 8'b00000000; // 3079 :   0 - 0x0
      12'hC08: dout <= 8'b00000000; // 3080 :   0 - 0x0 -- Background 0x81
      12'hC09: dout <= 8'b00000000; // 3081 :   0 - 0x0
      12'hC0A: dout <= 8'b00000000; // 3082 :   0 - 0x0
      12'hC0B: dout <= 8'b00000000; // 3083 :   0 - 0x0
      12'hC0C: dout <= 8'b00000000; // 3084 :   0 - 0x0
      12'hC0D: dout <= 8'b00000000; // 3085 :   0 - 0x0
      12'hC0E: dout <= 8'b00000000; // 3086 :   0 - 0x0
      12'hC0F: dout <= 8'b00000000; // 3087 :   0 - 0x0
      12'hC10: dout <= 8'b00000000; // 3088 :   0 - 0x0 -- Background 0x82
      12'hC11: dout <= 8'b11000000; // 3089 : 192 - 0xc0
      12'hC12: dout <= 8'b11110000; // 3090 : 240 - 0xf0
      12'hC13: dout <= 8'b11110000; // 3091 : 240 - 0xf0
      12'hC14: dout <= 8'b11101100; // 3092 : 236 - 0xec
      12'hC15: dout <= 8'b11100000; // 3093 : 224 - 0xe0
      12'hC16: dout <= 8'b11111100; // 3094 : 252 - 0xfc
      12'hC17: dout <= 8'b00000000; // 3095 :   0 - 0x0
      12'hC18: dout <= 8'b00000000; // 3096 :   0 - 0x0 -- Background 0x83
      12'hC19: dout <= 8'b00000000; // 3097 :   0 - 0x0
      12'hC1A: dout <= 8'b00000000; // 3098 :   0 - 0x0
      12'hC1B: dout <= 8'b00000000; // 3099 :   0 - 0x0
      12'hC1C: dout <= 8'b00000000; // 3100 :   0 - 0x0
      12'hC1D: dout <= 8'b00000000; // 3101 :   0 - 0x0
      12'hC1E: dout <= 8'b11100000; // 3102 : 224 - 0xe0
      12'hC1F: dout <= 8'b00000000; // 3103 :   0 - 0x0
      12'hC20: dout <= 8'b00000000; // 3104 :   0 - 0x0 -- Background 0x84
      12'hC21: dout <= 8'b00000011; // 3105 :   3 - 0x3
      12'hC22: dout <= 8'b00001111; // 3106 :  15 - 0xf
      12'hC23: dout <= 8'b00011111; // 3107 :  31 - 0x1f
      12'hC24: dout <= 8'b00011111; // 3108 :  31 - 0x1f
      12'hC25: dout <= 8'b00111111; // 3109 :  63 - 0x3f
      12'hC26: dout <= 8'b00111111; // 3110 :  63 - 0x3f
      12'hC27: dout <= 8'b00000000; // 3111 :   0 - 0x0
      12'hC28: dout <= 8'b00000000; // 3112 :   0 - 0x0 -- Background 0x85
      12'hC29: dout <= 8'b00000000; // 3113 :   0 - 0x0
      12'hC2A: dout <= 8'b00000000; // 3114 :   0 - 0x0
      12'hC2B: dout <= 8'b00000000; // 3115 :   0 - 0x0
      12'hC2C: dout <= 8'b00000000; // 3116 :   0 - 0x0
      12'hC2D: dout <= 8'b00001000; // 3117 :   8 - 0x8
      12'hC2E: dout <= 8'b00001110; // 3118 :  14 - 0xe
      12'hC2F: dout <= 8'b00000000; // 3119 :   0 - 0x0
      12'hC30: dout <= 8'b00000000; // 3120 :   0 - 0x0 -- Background 0x86
      12'hC31: dout <= 8'b11000000; // 3121 : 192 - 0xc0
      12'hC32: dout <= 8'b11110000; // 3122 : 240 - 0xf0
      12'hC33: dout <= 8'b11110000; // 3123 : 240 - 0xf0
      12'hC34: dout <= 8'b11101100; // 3124 : 236 - 0xec
      12'hC35: dout <= 8'b11100000; // 3125 : 224 - 0xe0
      12'hC36: dout <= 8'b11111100; // 3126 : 252 - 0xfc
      12'hC37: dout <= 8'b00000000; // 3127 :   0 - 0x0
      12'hC38: dout <= 8'b00000000; // 3128 :   0 - 0x0 -- Background 0x87
      12'hC39: dout <= 8'b00000000; // 3129 :   0 - 0x0
      12'hC3A: dout <= 8'b00000000; // 3130 :   0 - 0x0
      12'hC3B: dout <= 8'b00000000; // 3131 :   0 - 0x0
      12'hC3C: dout <= 8'b00000000; // 3132 :   0 - 0x0
      12'hC3D: dout <= 8'b00000110; // 3133 :   6 - 0x6
      12'hC3E: dout <= 8'b00001100; // 3134 :  12 - 0xc
      12'hC3F: dout <= 8'b00000000; // 3135 :   0 - 0x0
      12'hC40: dout <= 8'b00000000; // 3136 :   0 - 0x0 -- Background 0x88
      12'hC41: dout <= 8'b00000011; // 3137 :   3 - 0x3
      12'hC42: dout <= 8'b00000011; // 3138 :   3 - 0x3
      12'hC43: dout <= 8'b00000100; // 3139 :   4 - 0x4
      12'hC44: dout <= 8'b00001111; // 3140 :  15 - 0xf
      12'hC45: dout <= 8'b00011111; // 3141 :  31 - 0x1f
      12'hC46: dout <= 8'b01101111; // 3142 : 111 - 0x6f
      12'hC47: dout <= 8'b01101111; // 3143 : 111 - 0x6f
      12'hC48: dout <= 8'b01101111; // 3144 : 111 - 0x6f -- Background 0x89
      12'hC49: dout <= 8'b01101111; // 3145 : 111 - 0x6f
      12'hC4A: dout <= 8'b00011111; // 3146 :  31 - 0x1f
      12'hC4B: dout <= 8'b00001111; // 3147 :  15 - 0xf
      12'hC4C: dout <= 8'b00000100; // 3148 :   4 - 0x4
      12'hC4D: dout <= 8'b00000011; // 3149 :   3 - 0x3
      12'hC4E: dout <= 8'b00000011; // 3150 :   3 - 0x3
      12'hC4F: dout <= 8'b00000000; // 3151 :   0 - 0x0
      12'hC50: dout <= 8'b00000000; // 3152 :   0 - 0x0 -- Background 0x8a
      12'hC51: dout <= 8'b00000000; // 3153 :   0 - 0x0
      12'hC52: dout <= 8'b00011000; // 3154 :  24 - 0x18
      12'hC53: dout <= 8'b00110111; // 3155 :  55 - 0x37
      12'hC54: dout <= 8'b00101111; // 3156 :  47 - 0x2f
      12'hC55: dout <= 8'b00011111; // 3157 :  31 - 0x1f
      12'hC56: dout <= 8'b00011111; // 3158 :  31 - 0x1f
      12'hC57: dout <= 8'b00011111; // 3159 :  31 - 0x1f
      12'hC58: dout <= 8'b00011111; // 3160 :  31 - 0x1f -- Background 0x8b
      12'hC59: dout <= 8'b00011111; // 3161 :  31 - 0x1f
      12'hC5A: dout <= 8'b00011111; // 3162 :  31 - 0x1f
      12'hC5B: dout <= 8'b00101111; // 3163 :  47 - 0x2f
      12'hC5C: dout <= 8'b00110111; // 3164 :  55 - 0x37
      12'hC5D: dout <= 8'b00011000; // 3165 :  24 - 0x18
      12'hC5E: dout <= 8'b00000000; // 3166 :   0 - 0x0
      12'hC5F: dout <= 8'b00000000; // 3167 :   0 - 0x0
      12'hC60: dout <= 8'b00000000; // 3168 :   0 - 0x0 -- Background 0x8c
      12'hC61: dout <= 8'b00000011; // 3169 :   3 - 0x3
      12'hC62: dout <= 8'b00000001; // 3170 :   1 - 0x1
      12'hC63: dout <= 8'b00011001; // 3171 :  25 - 0x19
      12'hC64: dout <= 8'b00111001; // 3172 :  57 - 0x39
      12'hC65: dout <= 8'b00011011; // 3173 :  27 - 0x1b
      12'hC66: dout <= 8'b00001111; // 3174 :  15 - 0xf
      12'hC67: dout <= 8'b00001111; // 3175 :  15 - 0xf
      12'hC68: dout <= 8'b01111111; // 3176 : 127 - 0x7f -- Background 0x8d
      12'hC69: dout <= 8'b01111111; // 3177 : 127 - 0x7f
      12'hC6A: dout <= 8'b00111111; // 3178 :  63 - 0x3f
      12'hC6B: dout <= 8'b00010111; // 3179 :  23 - 0x17
      12'hC6C: dout <= 8'b00000110; // 3180 :   6 - 0x6
      12'hC6D: dout <= 8'b00000100; // 3181 :   4 - 0x4
      12'hC6E: dout <= 8'b00000111; // 3182 :   7 - 0x7
      12'hC6F: dout <= 8'b00000000; // 3183 :   0 - 0x0
      12'hC70: dout <= 8'b00000000; // 3184 :   0 - 0x0 -- Background 0x8e
      12'hC71: dout <= 8'b11000000; // 3185 : 192 - 0xc0
      12'hC72: dout <= 8'b11110000; // 3186 : 240 - 0xf0
      12'hC73: dout <= 8'b10111000; // 3187 : 184 - 0xb8
      12'hC74: dout <= 8'b10011100; // 3188 : 156 - 0x9c
      12'hC75: dout <= 8'b11111100; // 3189 : 252 - 0xfc
      12'hC76: dout <= 8'b11111110; // 3190 : 254 - 0xfe
      12'hC77: dout <= 8'b11000000; // 3191 : 192 - 0xc0
      12'hC78: dout <= 8'b11111110; // 3192 : 254 - 0xfe -- Background 0x8f
      12'hC79: dout <= 8'b11111110; // 3193 : 254 - 0xfe
      12'hC7A: dout <= 8'b11111000; // 3194 : 248 - 0xf8
      12'hC7B: dout <= 8'b11110000; // 3195 : 240 - 0xf0
      12'hC7C: dout <= 8'b11000000; // 3196 : 192 - 0xc0
      12'hC7D: dout <= 8'b00000000; // 3197 :   0 - 0x0
      12'hC7E: dout <= 8'b00000000; // 3198 :   0 - 0x0
      12'hC7F: dout <= 8'b10000000; // 3199 : 128 - 0x80
      12'hC80: dout <= 8'b00000000; // 3200 :   0 - 0x0 -- Background 0x90
      12'hC81: dout <= 8'b00000001; // 3201 :   1 - 0x1
      12'hC82: dout <= 8'b00001001; // 3202 :   9 - 0x9
      12'hC83: dout <= 8'b00011001; // 3203 :  25 - 0x19
      12'hC84: dout <= 8'b00011100; // 3204 :  28 - 0x1c
      12'hC85: dout <= 8'b00001101; // 3205 :  13 - 0xd
      12'hC86: dout <= 8'b00001111; // 3206 :  15 - 0xf
      12'hC87: dout <= 8'b00101111; // 3207 :  47 - 0x2f
      12'hC88: dout <= 8'b01111111; // 3208 : 127 - 0x7f -- Background 0x91
      12'hC89: dout <= 8'b01111111; // 3209 : 127 - 0x7f
      12'hC8A: dout <= 8'b00111111; // 3210 :  63 - 0x3f
      12'hC8B: dout <= 8'b00011011; // 3211 :  27 - 0x1b
      12'hC8C: dout <= 8'b00000011; // 3212 :   3 - 0x3
      12'hC8D: dout <= 8'b00000011; // 3213 :   3 - 0x3
      12'hC8E: dout <= 8'b00000001; // 3214 :   1 - 0x1
      12'hC8F: dout <= 8'b00000000; // 3215 :   0 - 0x0
      12'hC90: dout <= 8'b00000000; // 3216 :   0 - 0x0 -- Background 0x92
      12'hC91: dout <= 8'b11000000; // 3217 : 192 - 0xc0
      12'hC92: dout <= 8'b11110000; // 3218 : 240 - 0xf0
      12'hC93: dout <= 8'b11011000; // 3219 : 216 - 0xd8
      12'hC94: dout <= 8'b11001100; // 3220 : 204 - 0xcc
      12'hC95: dout <= 8'b11111100; // 3221 : 252 - 0xfc
      12'hC96: dout <= 8'b11111110; // 3222 : 254 - 0xfe
      12'hC97: dout <= 8'b11100000; // 3223 : 224 - 0xe0
      12'hC98: dout <= 8'b11111110; // 3224 : 254 - 0xfe -- Background 0x93
      12'hC99: dout <= 8'b11111110; // 3225 : 254 - 0xfe
      12'hC9A: dout <= 8'b11111000; // 3226 : 248 - 0xf8
      12'hC9B: dout <= 8'b01110000; // 3227 : 112 - 0x70
      12'hC9C: dout <= 8'b01000000; // 3228 :  64 - 0x40
      12'hC9D: dout <= 8'b00000000; // 3229 :   0 - 0x0
      12'hC9E: dout <= 8'b11000000; // 3230 : 192 - 0xc0
      12'hC9F: dout <= 8'b00100000; // 3231 :  32 - 0x20
      12'hCA0: dout <= 8'b00000000; // 3232 :   0 - 0x0 -- Background 0x94
      12'hCA1: dout <= 8'b00000000; // 3233 :   0 - 0x0
      12'hCA2: dout <= 8'b00001100; // 3234 :  12 - 0xc
      12'hCA3: dout <= 8'b00001110; // 3235 :  14 - 0xe
      12'hCA4: dout <= 8'b00000110; // 3236 :   6 - 0x6
      12'hCA5: dout <= 8'b00100110; // 3237 :  38 - 0x26
      12'hCA6: dout <= 8'b00110111; // 3238 :  55 - 0x37
      12'hCA7: dout <= 8'b00110011; // 3239 :  51 - 0x33
      12'hCA8: dout <= 8'b01111111; // 3240 : 127 - 0x7f -- Background 0x95
      12'hCA9: dout <= 8'b01111111; // 3241 : 127 - 0x7f
      12'hCAA: dout <= 8'b00111111; // 3242 :  63 - 0x3f
      12'hCAB: dout <= 8'b00011111; // 3243 :  31 - 0x1f
      12'hCAC: dout <= 8'b00001110; // 3244 :  14 - 0xe
      12'hCAD: dout <= 8'b00000000; // 3245 :   0 - 0x0
      12'hCAE: dout <= 8'b00000000; // 3246 :   0 - 0x0
      12'hCAF: dout <= 8'b00000000; // 3247 :   0 - 0x0
      12'hCB0: dout <= 8'b00000000; // 3248 :   0 - 0x0 -- Background 0x96
      12'hCB1: dout <= 8'b11000000; // 3249 : 192 - 0xc0
      12'hCB2: dout <= 8'b11110000; // 3250 : 240 - 0xf0
      12'hCB3: dout <= 8'b01101000; // 3251 : 104 - 0x68
      12'hCB4: dout <= 8'b01100100; // 3252 : 100 - 0x64
      12'hCB5: dout <= 8'b11111100; // 3253 : 252 - 0xfc
      12'hCB6: dout <= 8'b11111110; // 3254 : 254 - 0xfe
      12'hCB7: dout <= 8'b11110000; // 3255 : 240 - 0xf0
      12'hCB8: dout <= 8'b11111111; // 3256 : 255 - 0xff -- Background 0x97
      12'hCB9: dout <= 8'b11111110; // 3257 : 254 - 0xfe
      12'hCBA: dout <= 8'b11111100; // 3258 : 252 - 0xfc
      12'hCBB: dout <= 8'b10110000; // 3259 : 176 - 0xb0
      12'hCBC: dout <= 8'b11000000; // 3260 : 192 - 0xc0
      12'hCBD: dout <= 8'b11000000; // 3261 : 192 - 0xc0
      12'hCBE: dout <= 8'b01110000; // 3262 : 112 - 0x70
      12'hCBF: dout <= 8'b00001000; // 3263 :   8 - 0x8
      12'hCC0: dout <= 8'b00000000; // 3264 :   0 - 0x0 -- Background 0x98
      12'hCC1: dout <= 8'b00000001; // 3265 :   1 - 0x1
      12'hCC2: dout <= 8'b00000000; // 3266 :   0 - 0x0
      12'hCC3: dout <= 8'b00000000; // 3267 :   0 - 0x0
      12'hCC4: dout <= 8'b00000000; // 3268 :   0 - 0x0
      12'hCC5: dout <= 8'b00000000; // 3269 :   0 - 0x0
      12'hCC6: dout <= 8'b00000001; // 3270 :   1 - 0x1
      12'hCC7: dout <= 8'b00000011; // 3271 :   3 - 0x3
      12'hCC8: dout <= 8'b00000111; // 3272 :   7 - 0x7 -- Background 0x99
      12'hCC9: dout <= 8'b00010111; // 3273 :  23 - 0x17
      12'hCCA: dout <= 8'b00101111; // 3274 :  47 - 0x2f
      12'hCCB: dout <= 8'b00011110; // 3275 :  30 - 0x1e
      12'hCCC: dout <= 8'b00010001; // 3276 :  17 - 0x11
      12'hCCD: dout <= 8'b00000000; // 3277 :   0 - 0x0
      12'hCCE: dout <= 8'b00000001; // 3278 :   1 - 0x1
      12'hCCF: dout <= 8'b00000000; // 3279 :   0 - 0x0
      12'hCD0: dout <= 8'b00000000; // 3280 :   0 - 0x0 -- Background 0x9a
      12'hCD1: dout <= 8'b00010000; // 3281 :  16 - 0x10
      12'hCD2: dout <= 8'b01111000; // 3282 : 120 - 0x78
      12'hCD3: dout <= 8'b01110100; // 3283 : 116 - 0x74
      12'hCD4: dout <= 8'b11111110; // 3284 : 254 - 0xfe
      12'hCD5: dout <= 8'b11111000; // 3285 : 248 - 0xf8
      12'hCD6: dout <= 8'b11111100; // 3286 : 252 - 0xfc
      12'hCD7: dout <= 8'b11111000; // 3287 : 248 - 0xf8
      12'hCD8: dout <= 8'b11111000; // 3288 : 248 - 0xf8 -- Background 0x9b
      12'hCD9: dout <= 8'b11010000; // 3289 : 208 - 0xd0
      12'hCDA: dout <= 8'b00110000; // 3290 :  48 - 0x30
      12'hCDB: dout <= 8'b01100000; // 3291 :  96 - 0x60
      12'hCDC: dout <= 8'b10000000; // 3292 : 128 - 0x80
      12'hCDD: dout <= 8'b00000000; // 3293 :   0 - 0x0
      12'hCDE: dout <= 8'b00000000; // 3294 :   0 - 0x0
      12'hCDF: dout <= 8'b00000000; // 3295 :   0 - 0x0
      12'hCE0: dout <= 8'b00000000; // 3296 :   0 - 0x0 -- Background 0x9c
      12'hCE1: dout <= 8'b00000001; // 3297 :   1 - 0x1
      12'hCE2: dout <= 8'b00000000; // 3298 :   0 - 0x0
      12'hCE3: dout <= 8'b00000000; // 3299 :   0 - 0x0
      12'hCE4: dout <= 8'b00000000; // 3300 :   0 - 0x0
      12'hCE5: dout <= 8'b00000000; // 3301 :   0 - 0x0
      12'hCE6: dout <= 8'b00000001; // 3302 :   1 - 0x1
      12'hCE7: dout <= 8'b00000011; // 3303 :   3 - 0x3
      12'hCE8: dout <= 8'b00000111; // 3304 :   7 - 0x7 -- Background 0x9d
      12'hCE9: dout <= 8'b00010111; // 3305 :  23 - 0x17
      12'hCEA: dout <= 8'b00101111; // 3306 :  47 - 0x2f
      12'hCEB: dout <= 8'b00011110; // 3307 :  30 - 0x1e
      12'hCEC: dout <= 8'b00010000; // 3308 :  16 - 0x10
      12'hCED: dout <= 8'b00000100; // 3309 :   4 - 0x4
      12'hCEE: dout <= 8'b00000000; // 3310 :   0 - 0x0
      12'hCEF: dout <= 8'b00000000; // 3311 :   0 - 0x0
      12'hCF0: dout <= 8'b00000000; // 3312 :   0 - 0x0 -- Background 0x9e
      12'hCF1: dout <= 8'b00010000; // 3313 :  16 - 0x10
      12'hCF2: dout <= 8'b01111000; // 3314 : 120 - 0x78
      12'hCF3: dout <= 8'b01110100; // 3315 : 116 - 0x74
      12'hCF4: dout <= 8'b11111110; // 3316 : 254 - 0xfe
      12'hCF5: dout <= 8'b11111000; // 3317 : 248 - 0xf8
      12'hCF6: dout <= 8'b11111100; // 3318 : 252 - 0xfc
      12'hCF7: dout <= 8'b11111000; // 3319 : 248 - 0xf8
      12'hCF8: dout <= 8'b11111000; // 3320 : 248 - 0xf8 -- Background 0x9f
      12'hCF9: dout <= 8'b11010000; // 3321 : 208 - 0xd0
      12'hCFA: dout <= 8'b00110000; // 3322 :  48 - 0x30
      12'hCFB: dout <= 8'b11000000; // 3323 : 192 - 0xc0
      12'hCFC: dout <= 8'b00000000; // 3324 :   0 - 0x0
      12'hCFD: dout <= 8'b00000000; // 3325 :   0 - 0x0
      12'hCFE: dout <= 8'b00000000; // 3326 :   0 - 0x0
      12'hCFF: dout <= 8'b00000000; // 3327 :   0 - 0x0
      12'hD00: dout <= 8'b00000000; // 3328 :   0 - 0x0 -- Background 0xa0
      12'hD01: dout <= 8'b00000011; // 3329 :   3 - 0x3
      12'hD02: dout <= 8'b00001111; // 3330 :  15 - 0xf
      12'hD03: dout <= 8'b00011111; // 3331 :  31 - 0x1f
      12'hD04: dout <= 8'b00111111; // 3332 :  63 - 0x3f
      12'hD05: dout <= 8'b00111111; // 3333 :  63 - 0x3f
      12'hD06: dout <= 8'b01111111; // 3334 : 127 - 0x7f
      12'hD07: dout <= 8'b01111111; // 3335 : 127 - 0x7f
      12'hD08: dout <= 8'b01111111; // 3336 : 127 - 0x7f -- Background 0xa1
      12'hD09: dout <= 8'b01111111; // 3337 : 127 - 0x7f
      12'hD0A: dout <= 8'b00111111; // 3338 :  63 - 0x3f
      12'hD0B: dout <= 8'b00111111; // 3339 :  63 - 0x3f
      12'hD0C: dout <= 8'b00011111; // 3340 :  31 - 0x1f
      12'hD0D: dout <= 8'b00000101; // 3341 :   5 - 0x5
      12'hD0E: dout <= 8'b00000010; // 3342 :   2 - 0x2
      12'hD0F: dout <= 8'b00000000; // 3343 :   0 - 0x0
      12'hD10: dout <= 8'b00000000; // 3344 :   0 - 0x0 -- Background 0xa2
      12'hD11: dout <= 8'b11000000; // 3345 : 192 - 0xc0
      12'hD12: dout <= 8'b11110000; // 3346 : 240 - 0xf0
      12'hD13: dout <= 8'b11111000; // 3347 : 248 - 0xf8
      12'hD14: dout <= 8'b11111000; // 3348 : 248 - 0xf8
      12'hD15: dout <= 8'b11111100; // 3349 : 252 - 0xfc
      12'hD16: dout <= 8'b11111010; // 3350 : 250 - 0xfa
      12'hD17: dout <= 8'b11111100; // 3351 : 252 - 0xfc
      12'hD18: dout <= 8'b11111010; // 3352 : 250 - 0xfa -- Background 0xa3
      12'hD19: dout <= 8'b11110100; // 3353 : 244 - 0xf4
      12'hD1A: dout <= 8'b11101000; // 3354 : 232 - 0xe8
      12'hD1B: dout <= 8'b11010100; // 3355 : 212 - 0xd4
      12'hD1C: dout <= 8'b10101000; // 3356 : 168 - 0xa8
      12'hD1D: dout <= 8'b01010000; // 3357 :  80 - 0x50
      12'hD1E: dout <= 8'b10000000; // 3358 : 128 - 0x80
      12'hD1F: dout <= 8'b00000000; // 3359 :   0 - 0x0
      12'hD20: dout <= 8'b00000000; // 3360 :   0 - 0x0 -- Background 0xa4
      12'hD21: dout <= 8'b00000000; // 3361 :   0 - 0x0
      12'hD22: dout <= 8'b00000000; // 3362 :   0 - 0x0
      12'hD23: dout <= 8'b00001110; // 3363 :  14 - 0xe
      12'hD24: dout <= 8'b00000000; // 3364 :   0 - 0x0
      12'hD25: dout <= 8'b00001010; // 3365 :  10 - 0xa
      12'hD26: dout <= 8'b01001010; // 3366 :  74 - 0x4a
      12'hD27: dout <= 8'b01100000; // 3367 :  96 - 0x60
      12'hD28: dout <= 8'b01111111; // 3368 : 127 - 0x7f -- Background 0xa5
      12'hD29: dout <= 8'b01111000; // 3369 : 120 - 0x78
      12'hD2A: dout <= 8'b00110111; // 3370 :  55 - 0x37
      12'hD2B: dout <= 8'b00111011; // 3371 :  59 - 0x3b
      12'hD2C: dout <= 8'b00111100; // 3372 :  60 - 0x3c
      12'hD2D: dout <= 8'b00011111; // 3373 :  31 - 0x1f
      12'hD2E: dout <= 8'b00000111; // 3374 :   7 - 0x7
      12'hD2F: dout <= 8'b00000000; // 3375 :   0 - 0x0
      12'hD30: dout <= 8'b00000000; // 3376 :   0 - 0x0 -- Background 0xa6
      12'hD31: dout <= 8'b00000000; // 3377 :   0 - 0x0
      12'hD32: dout <= 8'b00000000; // 3378 :   0 - 0x0
      12'hD33: dout <= 8'b01110000; // 3379 : 112 - 0x70
      12'hD34: dout <= 8'b00000000; // 3380 :   0 - 0x0
      12'hD35: dout <= 8'b01010000; // 3381 :  80 - 0x50
      12'hD36: dout <= 8'b01010010; // 3382 :  82 - 0x52
      12'hD37: dout <= 8'b00000110; // 3383 :   6 - 0x6
      12'hD38: dout <= 8'b11111100; // 3384 : 252 - 0xfc -- Background 0xa7
      12'hD39: dout <= 8'b00011010; // 3385 :  26 - 0x1a
      12'hD3A: dout <= 8'b11101100; // 3386 : 236 - 0xec
      12'hD3B: dout <= 8'b11011000; // 3387 : 216 - 0xd8
      12'hD3C: dout <= 8'b00110100; // 3388 :  52 - 0x34
      12'hD3D: dout <= 8'b11101000; // 3389 : 232 - 0xe8
      12'hD3E: dout <= 8'b11000000; // 3390 : 192 - 0xc0
      12'hD3F: dout <= 8'b00000000; // 3391 :   0 - 0x0
      12'hD40: dout <= 8'b00000000; // 3392 :   0 - 0x0 -- Background 0xa8
      12'hD41: dout <= 8'b00000000; // 3393 :   0 - 0x0
      12'hD42: dout <= 8'b00000000; // 3394 :   0 - 0x0
      12'hD43: dout <= 8'b00001110; // 3395 :  14 - 0xe
      12'hD44: dout <= 8'b00000000; // 3396 :   0 - 0x0
      12'hD45: dout <= 8'b00001110; // 3397 :  14 - 0xe
      12'hD46: dout <= 8'b01001010; // 3398 :  74 - 0x4a
      12'hD47: dout <= 8'b01100000; // 3399 :  96 - 0x60
      12'hD48: dout <= 8'b01111111; // 3400 : 127 - 0x7f -- Background 0xa9
      12'hD49: dout <= 8'b01111100; // 3401 : 124 - 0x7c
      12'hD4A: dout <= 8'b01111011; // 3402 : 123 - 0x7b
      12'hD4B: dout <= 8'b01110111; // 3403 : 119 - 0x77
      12'hD4C: dout <= 8'b01111000; // 3404 : 120 - 0x78
      12'hD4D: dout <= 8'b01111111; // 3405 : 127 - 0x7f
      12'hD4E: dout <= 8'b01111111; // 3406 : 127 - 0x7f
      12'hD4F: dout <= 8'b00000000; // 3407 :   0 - 0x0
      12'hD50: dout <= 8'b00000000; // 3408 :   0 - 0x0 -- Background 0xaa
      12'hD51: dout <= 8'b00000000; // 3409 :   0 - 0x0
      12'hD52: dout <= 8'b00000000; // 3410 :   0 - 0x0
      12'hD53: dout <= 8'b01110000; // 3411 : 112 - 0x70
      12'hD54: dout <= 8'b00000000; // 3412 :   0 - 0x0
      12'hD55: dout <= 8'b01110000; // 3413 : 112 - 0x70
      12'hD56: dout <= 8'b01010010; // 3414 :  82 - 0x52
      12'hD57: dout <= 8'b00000110; // 3415 :   6 - 0x6
      12'hD58: dout <= 8'b11111100; // 3416 : 252 - 0xfc -- Background 0xab
      12'hD59: dout <= 8'b00111010; // 3417 :  58 - 0x3a
      12'hD5A: dout <= 8'b11011100; // 3418 : 220 - 0xdc
      12'hD5B: dout <= 8'b11101010; // 3419 : 234 - 0xea
      12'hD5C: dout <= 8'b00011100; // 3420 :  28 - 0x1c
      12'hD5D: dout <= 8'b11111010; // 3421 : 250 - 0xfa
      12'hD5E: dout <= 8'b11110100; // 3422 : 244 - 0xf4
      12'hD5F: dout <= 8'b00000000; // 3423 :   0 - 0x0
      12'hD60: dout <= 8'b00000000; // 3424 :   0 - 0x0 -- Background 0xac
      12'hD61: dout <= 8'b00000011; // 3425 :   3 - 0x3
      12'hD62: dout <= 8'b00001111; // 3426 :  15 - 0xf
      12'hD63: dout <= 8'b00001111; // 3427 :  15 - 0xf
      12'hD64: dout <= 8'b00011111; // 3428 :  31 - 0x1f
      12'hD65: dout <= 8'b01011111; // 3429 :  95 - 0x5f
      12'hD66: dout <= 8'b01010000; // 3430 :  80 - 0x50
      12'hD67: dout <= 8'b00010000; // 3431 :  16 - 0x10
      12'hD68: dout <= 8'b00000000; // 3432 :   0 - 0x0 -- Background 0xad
      12'hD69: dout <= 8'b11111010; // 3433 : 250 - 0xfa
      12'hD6A: dout <= 8'b11111010; // 3434 : 250 - 0xfa
      12'hD6B: dout <= 8'b11111010; // 3435 : 250 - 0xfa
      12'hD6C: dout <= 8'b10111010; // 3436 : 186 - 0xba
      12'hD6D: dout <= 8'b10011010; // 3437 : 154 - 0x9a
      12'hD6E: dout <= 8'b00001010; // 3438 :  10 - 0xa
      12'hD6F: dout <= 8'b00000010; // 3439 :   2 - 0x2
      12'hD70: dout <= 8'b00000000; // 3440 :   0 - 0x0 -- Background 0xae
      12'hD71: dout <= 8'b00000011; // 3441 :   3 - 0x3
      12'hD72: dout <= 8'b00001111; // 3442 :  15 - 0xf
      12'hD73: dout <= 8'b00001111; // 3443 :  15 - 0xf
      12'hD74: dout <= 8'b00011111; // 3444 :  31 - 0x1f
      12'hD75: dout <= 8'b01011111; // 3445 :  95 - 0x5f
      12'hD76: dout <= 8'b01010000; // 3446 :  80 - 0x50
      12'hD77: dout <= 8'b00010111; // 3447 :  23 - 0x17
      12'hD78: dout <= 8'b00000000; // 3448 :   0 - 0x0 -- Background 0xaf
      12'hD79: dout <= 8'b11111010; // 3449 : 250 - 0xfa
      12'hD7A: dout <= 8'b11111010; // 3450 : 250 - 0xfa
      12'hD7B: dout <= 8'b11111010; // 3451 : 250 - 0xfa
      12'hD7C: dout <= 8'b00111010; // 3452 :  58 - 0x3a
      12'hD7D: dout <= 8'b01011010; // 3453 :  90 - 0x5a
      12'hD7E: dout <= 8'b01101010; // 3454 : 106 - 0x6a
      12'hD7F: dout <= 8'b11110010; // 3455 : 242 - 0xf2
      12'hD80: dout <= 8'b00000000; // 3456 :   0 - 0x0 -- Background 0xb0
      12'hD81: dout <= 8'b00000000; // 3457 :   0 - 0x0
      12'hD82: dout <= 8'b00000011; // 3458 :   3 - 0x3
      12'hD83: dout <= 8'b00001111; // 3459 :  15 - 0xf
      12'hD84: dout <= 8'b00111011; // 3460 :  59 - 0x3b
      12'hD85: dout <= 8'b00111111; // 3461 :  63 - 0x3f
      12'hD86: dout <= 8'b01101111; // 3462 : 111 - 0x6f
      12'hD87: dout <= 8'b01111101; // 3463 : 125 - 0x7d
      12'hD88: dout <= 8'b00001111; // 3464 :  15 - 0xf -- Background 0xb1
      12'hD89: dout <= 8'b01110000; // 3465 : 112 - 0x70
      12'hD8A: dout <= 8'b01111111; // 3466 : 127 - 0x7f
      12'hD8B: dout <= 8'b00001111; // 3467 :  15 - 0xf
      12'hD8C: dout <= 8'b01110000; // 3468 : 112 - 0x70
      12'hD8D: dout <= 8'b01111111; // 3469 : 127 - 0x7f
      12'hD8E: dout <= 8'b00001111; // 3470 :  15 - 0xf
      12'hD8F: dout <= 8'b00000000; // 3471 :   0 - 0x0
      12'hD90: dout <= 8'b00000000; // 3472 :   0 - 0x0 -- Background 0xb2
      12'hD91: dout <= 8'b00000000; // 3473 :   0 - 0x0
      12'hD92: dout <= 8'b11000000; // 3474 : 192 - 0xc0
      12'hD93: dout <= 8'b11110000; // 3475 : 240 - 0xf0
      12'hD94: dout <= 8'b10111100; // 3476 : 188 - 0xbc
      12'hD95: dout <= 8'b11110100; // 3477 : 244 - 0xf4
      12'hD96: dout <= 8'b11111110; // 3478 : 254 - 0xfe
      12'hD97: dout <= 8'b11011110; // 3479 : 222 - 0xde
      12'hD98: dout <= 8'b11110000; // 3480 : 240 - 0xf0 -- Background 0xb3
      12'hD99: dout <= 8'b00001110; // 3481 :  14 - 0xe
      12'hD9A: dout <= 8'b11111110; // 3482 : 254 - 0xfe
      12'hD9B: dout <= 8'b11110000; // 3483 : 240 - 0xf0
      12'hD9C: dout <= 8'b00001110; // 3484 :  14 - 0xe
      12'hD9D: dout <= 8'b11111110; // 3485 : 254 - 0xfe
      12'hD9E: dout <= 8'b11110000; // 3486 : 240 - 0xf0
      12'hD9F: dout <= 8'b00000000; // 3487 :   0 - 0x0
      12'hDA0: dout <= 8'b00000000; // 3488 :   0 - 0x0 -- Background 0xb4
      12'hDA1: dout <= 8'b00000000; // 3489 :   0 - 0x0
      12'hDA2: dout <= 8'b00000011; // 3490 :   3 - 0x3
      12'hDA3: dout <= 8'b00001111; // 3491 :  15 - 0xf
      12'hDA4: dout <= 8'b00111011; // 3492 :  59 - 0x3b
      12'hDA5: dout <= 8'b00111111; // 3493 :  63 - 0x3f
      12'hDA6: dout <= 8'b01101111; // 3494 : 111 - 0x6f
      12'hDA7: dout <= 8'b01111101; // 3495 : 125 - 0x7d
      12'hDA8: dout <= 8'b00001111; // 3496 :  15 - 0xf -- Background 0xb5
      12'hDA9: dout <= 8'b01110000; // 3497 : 112 - 0x70
      12'hDAA: dout <= 8'b01111111; // 3498 : 127 - 0x7f
      12'hDAB: dout <= 8'b00001111; // 3499 :  15 - 0xf
      12'hDAC: dout <= 8'b01110000; // 3500 : 112 - 0x70
      12'hDAD: dout <= 8'b01111111; // 3501 : 127 - 0x7f
      12'hDAE: dout <= 8'b00001111; // 3502 :  15 - 0xf
      12'hDAF: dout <= 8'b00000000; // 3503 :   0 - 0x0
      12'hDB0: dout <= 8'b00000000; // 3504 :   0 - 0x0 -- Background 0xb6
      12'hDB1: dout <= 8'b00000000; // 3505 :   0 - 0x0
      12'hDB2: dout <= 8'b11000000; // 3506 : 192 - 0xc0
      12'hDB3: dout <= 8'b11110000; // 3507 : 240 - 0xf0
      12'hDB4: dout <= 8'b10111100; // 3508 : 188 - 0xbc
      12'hDB5: dout <= 8'b11110100; // 3509 : 244 - 0xf4
      12'hDB6: dout <= 8'b11111110; // 3510 : 254 - 0xfe
      12'hDB7: dout <= 8'b11011110; // 3511 : 222 - 0xde
      12'hDB8: dout <= 8'b11110000; // 3512 : 240 - 0xf0 -- Background 0xb7
      12'hDB9: dout <= 8'b00001110; // 3513 :  14 - 0xe
      12'hDBA: dout <= 8'b11111110; // 3514 : 254 - 0xfe
      12'hDBB: dout <= 8'b11110000; // 3515 : 240 - 0xf0
      12'hDBC: dout <= 8'b00001110; // 3516 :  14 - 0xe
      12'hDBD: dout <= 8'b11111110; // 3517 : 254 - 0xfe
      12'hDBE: dout <= 8'b11110000; // 3518 : 240 - 0xf0
      12'hDBF: dout <= 8'b00000000; // 3519 :   0 - 0x0
      12'hDC0: dout <= 8'b00000000; // 3520 :   0 - 0x0 -- Background 0xb8
      12'hDC1: dout <= 8'b00000000; // 3521 :   0 - 0x0
      12'hDC2: dout <= 8'b00000011; // 3522 :   3 - 0x3
      12'hDC3: dout <= 8'b00001111; // 3523 :  15 - 0xf
      12'hDC4: dout <= 8'b00111011; // 3524 :  59 - 0x3b
      12'hDC5: dout <= 8'b00111111; // 3525 :  63 - 0x3f
      12'hDC6: dout <= 8'b01101111; // 3526 : 111 - 0x6f
      12'hDC7: dout <= 8'b01111101; // 3527 : 125 - 0x7d
      12'hDC8: dout <= 8'b00001111; // 3528 :  15 - 0xf -- Background 0xb9
      12'hDC9: dout <= 8'b00100000; // 3529 :  32 - 0x20
      12'hDCA: dout <= 8'b01010101; // 3530 :  85 - 0x55
      12'hDCB: dout <= 8'b00001010; // 3531 :  10 - 0xa
      12'hDCC: dout <= 8'b01110000; // 3532 : 112 - 0x70
      12'hDCD: dout <= 8'b01111111; // 3533 : 127 - 0x7f
      12'hDCE: dout <= 8'b00001111; // 3534 :  15 - 0xf
      12'hDCF: dout <= 8'b00000000; // 3535 :   0 - 0x0
      12'hDD0: dout <= 8'b00000000; // 3536 :   0 - 0x0 -- Background 0xba
      12'hDD1: dout <= 8'b00000000; // 3537 :   0 - 0x0
      12'hDD2: dout <= 8'b11000000; // 3538 : 192 - 0xc0
      12'hDD3: dout <= 8'b11110000; // 3539 : 240 - 0xf0
      12'hDD4: dout <= 8'b10111100; // 3540 : 188 - 0xbc
      12'hDD5: dout <= 8'b11110100; // 3541 : 244 - 0xf4
      12'hDD6: dout <= 8'b11111110; // 3542 : 254 - 0xfe
      12'hDD7: dout <= 8'b11011110; // 3543 : 222 - 0xde
      12'hDD8: dout <= 8'b11110000; // 3544 : 240 - 0xf0 -- Background 0xbb
      12'hDD9: dout <= 8'b00001010; // 3545 :  10 - 0xa
      12'hDDA: dout <= 8'b01010100; // 3546 :  84 - 0x54
      12'hDDB: dout <= 8'b10100000; // 3547 : 160 - 0xa0
      12'hDDC: dout <= 8'b00001110; // 3548 :  14 - 0xe
      12'hDDD: dout <= 8'b11111110; // 3549 : 254 - 0xfe
      12'hDDE: dout <= 8'b11110000; // 3550 : 240 - 0xf0
      12'hDDF: dout <= 8'b00000000; // 3551 :   0 - 0x0
      12'hDE0: dout <= 8'b00000000; // 3552 :   0 - 0x0 -- Background 0xbc
      12'hDE1: dout <= 8'b01110011; // 3553 : 115 - 0x73
      12'hDE2: dout <= 8'b01111011; // 3554 : 123 - 0x7b
      12'hDE3: dout <= 8'b01111111; // 3555 : 127 - 0x7f
      12'hDE4: dout <= 8'b00111111; // 3556 :  63 - 0x3f
      12'hDE5: dout <= 8'b00011100; // 3557 :  28 - 0x1c
      12'hDE6: dout <= 8'b01111011; // 3558 : 123 - 0x7b
      12'hDE7: dout <= 8'b01111011; // 3559 : 123 - 0x7b
      12'hDE8: dout <= 8'b01111011; // 3560 : 123 - 0x7b -- Background 0xbd
      12'hDE9: dout <= 8'b01111011; // 3561 : 123 - 0x7b
      12'hDEA: dout <= 8'b00011100; // 3562 :  28 - 0x1c
      12'hDEB: dout <= 8'b00111111; // 3563 :  63 - 0x3f
      12'hDEC: dout <= 8'b01111111; // 3564 : 127 - 0x7f
      12'hDED: dout <= 8'b01111011; // 3565 : 123 - 0x7b
      12'hDEE: dout <= 8'b01110011; // 3566 : 115 - 0x73
      12'hDEF: dout <= 8'b00000000; // 3567 :   0 - 0x0
      12'hDF0: dout <= 8'b00000000; // 3568 :   0 - 0x0 -- Background 0xbe
      12'hDF1: dout <= 8'b11001110; // 3569 : 206 - 0xce
      12'hDF2: dout <= 8'b11011110; // 3570 : 222 - 0xde
      12'hDF3: dout <= 8'b11111110; // 3571 : 254 - 0xfe
      12'hDF4: dout <= 8'b11111100; // 3572 : 252 - 0xfc
      12'hDF5: dout <= 8'b00111000; // 3573 :  56 - 0x38
      12'hDF6: dout <= 8'b11011110; // 3574 : 222 - 0xde
      12'hDF7: dout <= 8'b11011110; // 3575 : 222 - 0xde
      12'hDF8: dout <= 8'b11011110; // 3576 : 222 - 0xde -- Background 0xbf
      12'hDF9: dout <= 8'b11011110; // 3577 : 222 - 0xde
      12'hDFA: dout <= 8'b00111000; // 3578 :  56 - 0x38
      12'hDFB: dout <= 8'b11111100; // 3579 : 252 - 0xfc
      12'hDFC: dout <= 8'b11111110; // 3580 : 254 - 0xfe
      12'hDFD: dout <= 8'b11011110; // 3581 : 222 - 0xde
      12'hDFE: dout <= 8'b11001110; // 3582 : 206 - 0xce
      12'hDFF: dout <= 8'b00000000; // 3583 :   0 - 0x0
      12'hE00: dout <= 8'b00000000; // 3584 :   0 - 0x0 -- Background 0xc0
      12'hE01: dout <= 8'b00000000; // 3585 :   0 - 0x0
      12'hE02: dout <= 8'b01000000; // 3586 :  64 - 0x40
      12'hE03: dout <= 8'b01100000; // 3587 :  96 - 0x60
      12'hE04: dout <= 8'b01100001; // 3588 :  97 - 0x61
      12'hE05: dout <= 8'b00000010; // 3589 :   2 - 0x2
      12'hE06: dout <= 8'b00000010; // 3590 :   2 - 0x2
      12'hE07: dout <= 8'b00000111; // 3591 :   7 - 0x7
      12'hE08: dout <= 8'b00000111; // 3592 :   7 - 0x7 -- Background 0xc1
      12'hE09: dout <= 8'b00000100; // 3593 :   4 - 0x4
      12'hE0A: dout <= 8'b00000111; // 3594 :   7 - 0x7
      12'hE0B: dout <= 8'b00000001; // 3595 :   1 - 0x1
      12'hE0C: dout <= 8'b00000000; // 3596 :   0 - 0x0
      12'hE0D: dout <= 8'b00010000; // 3597 :  16 - 0x10
      12'hE0E: dout <= 8'b00101000; // 3598 :  40 - 0x28
      12'hE0F: dout <= 8'b00000000; // 3599 :   0 - 0x0
      12'hE10: dout <= 8'b00000000; // 3600 :   0 - 0x0 -- Background 0xc2
      12'hE11: dout <= 8'b00000000; // 3601 :   0 - 0x0
      12'hE12: dout <= 8'b00000010; // 3602 :   2 - 0x2
      12'hE13: dout <= 8'b00000110; // 3603 :   6 - 0x6
      12'hE14: dout <= 8'b11100110; // 3604 : 230 - 0xe6
      12'hE15: dout <= 8'b10100000; // 3605 : 160 - 0xa0
      12'hE16: dout <= 8'b10100000; // 3606 : 160 - 0xa0
      12'hE17: dout <= 8'b11110000; // 3607 : 240 - 0xf0
      12'hE18: dout <= 8'b11110000; // 3608 : 240 - 0xf0 -- Background 0xc3
      12'hE19: dout <= 8'b00110000; // 3609 :  48 - 0x30
      12'hE1A: dout <= 8'b11000000; // 3610 : 192 - 0xc0
      12'hE1B: dout <= 8'b10000000; // 3611 : 128 - 0x80
      12'hE1C: dout <= 8'b00000000; // 3612 :   0 - 0x0
      12'hE1D: dout <= 8'b00001000; // 3613 :   8 - 0x8
      12'hE1E: dout <= 8'b00010100; // 3614 :  20 - 0x14
      12'hE1F: dout <= 8'b00000000; // 3615 :   0 - 0x0
      12'hE20: dout <= 8'b00000000; // 3616 :   0 - 0x0 -- Background 0xc4
      12'hE21: dout <= 8'b00000101; // 3617 :   5 - 0x5
      12'hE22: dout <= 8'b00000111; // 3618 :   7 - 0x7
      12'hE23: dout <= 8'b00000000; // 3619 :   0 - 0x0
      12'hE24: dout <= 8'b00000000; // 3620 :   0 - 0x0
      12'hE25: dout <= 8'b00000000; // 3621 :   0 - 0x0
      12'hE26: dout <= 8'b00000000; // 3622 :   0 - 0x0
      12'hE27: dout <= 8'b00000001; // 3623 :   1 - 0x1
      12'hE28: dout <= 8'b00000010; // 3624 :   2 - 0x2 -- Background 0xc5
      12'hE29: dout <= 8'b00000111; // 3625 :   7 - 0x7
      12'hE2A: dout <= 8'b00100111; // 3626 :  39 - 0x27
      12'hE2B: dout <= 8'b01010011; // 3627 :  83 - 0x53
      12'hE2C: dout <= 8'b00000000; // 3628 :   0 - 0x0
      12'hE2D: dout <= 8'b00000010; // 3629 :   2 - 0x2
      12'hE2E: dout <= 8'b00000101; // 3630 :   5 - 0x5
      12'hE2F: dout <= 8'b00000000; // 3631 :   0 - 0x0
      12'hE30: dout <= 8'b00000000; // 3632 :   0 - 0x0 -- Background 0xc6
      12'hE31: dout <= 8'b00000000; // 3633 :   0 - 0x0
      12'hE32: dout <= 8'b00000000; // 3634 :   0 - 0x0
      12'hE33: dout <= 8'b00000000; // 3635 :   0 - 0x0
      12'hE34: dout <= 8'b00000000; // 3636 :   0 - 0x0
      12'hE35: dout <= 8'b01100000; // 3637 :  96 - 0x60
      12'hE36: dout <= 8'b11011000; // 3638 : 216 - 0xd8
      12'hE37: dout <= 8'b10110000; // 3639 : 176 - 0xb0
      12'hE38: dout <= 8'b11101000; // 3640 : 232 - 0xe8 -- Background 0xc7
      12'hE39: dout <= 8'b01111000; // 3641 : 120 - 0x78
      12'hE3A: dout <= 8'b10110110; // 3642 : 182 - 0xb6
      12'hE3B: dout <= 8'b11100100; // 3643 : 228 - 0xe4
      12'hE3C: dout <= 8'b00000110; // 3644 :   6 - 0x6
      12'hE3D: dout <= 8'b00000000; // 3645 :   0 - 0x0
      12'hE3E: dout <= 8'b00000000; // 3646 :   0 - 0x0
      12'hE3F: dout <= 8'b00000000; // 3647 :   0 - 0x0
      12'hE40: dout <= 8'b00000000; // 3648 :   0 - 0x0 -- Background 0xc8
      12'hE41: dout <= 8'b00000000; // 3649 :   0 - 0x0
      12'hE42: dout <= 8'b01000000; // 3650 :  64 - 0x40
      12'hE43: dout <= 8'b00100000; // 3651 :  32 - 0x20
      12'hE44: dout <= 8'b01000000; // 3652 :  64 - 0x40
      12'hE45: dout <= 8'b00000111; // 3653 :   7 - 0x7
      12'hE46: dout <= 8'b00000101; // 3654 :   5 - 0x5
      12'hE47: dout <= 8'b00001101; // 3655 :  13 - 0xd
      12'hE48: dout <= 8'b00001101; // 3656 :  13 - 0xd -- Background 0xc9
      12'hE49: dout <= 8'b00000101; // 3657 :   5 - 0x5
      12'hE4A: dout <= 8'b00000011; // 3658 :   3 - 0x3
      12'hE4B: dout <= 8'b01000011; // 3659 :  67 - 0x43
      12'hE4C: dout <= 8'b00100000; // 3660 :  32 - 0x20
      12'hE4D: dout <= 8'b01000000; // 3661 :  64 - 0x40
      12'hE4E: dout <= 8'b00000000; // 3662 :   0 - 0x0
      12'hE4F: dout <= 8'b00000000; // 3663 :   0 - 0x0
      12'hE50: dout <= 8'b00000000; // 3664 :   0 - 0x0 -- Background 0xca
      12'hE51: dout <= 8'b00011100; // 3665 :  28 - 0x1c
      12'hE52: dout <= 8'b00011000; // 3666 :  24 - 0x18
      12'hE53: dout <= 8'b00000000; // 3667 :   0 - 0x0
      12'hE54: dout <= 8'b00000000; // 3668 :   0 - 0x0
      12'hE55: dout <= 8'b10000000; // 3669 : 128 - 0x80
      12'hE56: dout <= 8'b11100000; // 3670 : 224 - 0xe0
      12'hE57: dout <= 8'b10010000; // 3671 : 144 - 0x90
      12'hE58: dout <= 8'b11110000; // 3672 : 240 - 0xf0 -- Background 0xcb
      12'hE59: dout <= 8'b10010000; // 3673 : 144 - 0x90
      12'hE5A: dout <= 8'b11110000; // 3674 : 240 - 0xf0
      12'hE5B: dout <= 8'b10000000; // 3675 : 128 - 0x80
      12'hE5C: dout <= 8'b00000000; // 3676 :   0 - 0x0
      12'hE5D: dout <= 8'b00011000; // 3677 :  24 - 0x18
      12'hE5E: dout <= 8'b00011100; // 3678 :  28 - 0x1c
      12'hE5F: dout <= 8'b00000000; // 3679 :   0 - 0x0
      12'hE60: dout <= 8'b00000000; // 3680 :   0 - 0x0 -- Background 0xcc
      12'hE61: dout <= 8'b00001000; // 3681 :   8 - 0x8
      12'hE62: dout <= 8'b00000100; // 3682 :   4 - 0x4
      12'hE63: dout <= 8'b00001000; // 3683 :   8 - 0x8
      12'hE64: dout <= 8'b00000000; // 3684 :   0 - 0x0
      12'hE65: dout <= 8'b01000110; // 3685 :  70 - 0x46
      12'hE66: dout <= 8'b00101111; // 3686 :  47 - 0x2f
      12'hE67: dout <= 8'b01001110; // 3687 :  78 - 0x4e
      12'hE68: dout <= 8'b00001101; // 3688 :  13 - 0xd -- Background 0xcd
      12'hE69: dout <= 8'b00001011; // 3689 :  11 - 0xb
      12'hE6A: dout <= 8'b00001111; // 3690 :  15 - 0xf
      12'hE6B: dout <= 8'b00000110; // 3691 :   6 - 0x6
      12'hE6C: dout <= 8'b00000011; // 3692 :   3 - 0x3
      12'hE6D: dout <= 8'b00011100; // 3693 :  28 - 0x1c
      12'hE6E: dout <= 8'b00010100; // 3694 :  20 - 0x14
      12'hE6F: dout <= 8'b00000000; // 3695 :   0 - 0x0
      12'hE70: dout <= 8'b00000000; // 3696 :   0 - 0x0 -- Background 0xce
      12'hE71: dout <= 8'b00000000; // 3697 :   0 - 0x0
      12'hE72: dout <= 8'b00000000; // 3698 :   0 - 0x0
      12'hE73: dout <= 8'b00000000; // 3699 :   0 - 0x0
      12'hE74: dout <= 8'b00000000; // 3700 :   0 - 0x0
      12'hE75: dout <= 8'b00000110; // 3701 :   6 - 0x6
      12'hE76: dout <= 8'b00000100; // 3702 :   4 - 0x4
      12'hE77: dout <= 8'b10000110; // 3703 : 134 - 0x86
      12'hE78: dout <= 8'b11000000; // 3704 : 192 - 0xc0 -- Background 0xcf
      12'hE79: dout <= 8'b01100000; // 3705 :  96 - 0x60
      12'hE7A: dout <= 8'b10100000; // 3706 : 160 - 0xa0
      12'hE7B: dout <= 8'b11000000; // 3707 : 192 - 0xc0
      12'hE7C: dout <= 8'b01000000; // 3708 :  64 - 0x40
      12'hE7D: dout <= 8'b00000000; // 3709 :   0 - 0x0
      12'hE7E: dout <= 8'b00000000; // 3710 :   0 - 0x0
      12'hE7F: dout <= 8'b00000000; // 3711 :   0 - 0x0
      12'hE80: dout <= 8'b00000000; // 3712 :   0 - 0x0 -- Background 0xd0
      12'hE81: dout <= 8'b00000000; // 3713 :   0 - 0x0
      12'hE82: dout <= 8'b00000000; // 3714 :   0 - 0x0
      12'hE83: dout <= 8'b00000000; // 3715 :   0 - 0x0
      12'hE84: dout <= 8'b00000100; // 3716 :   4 - 0x4
      12'hE85: dout <= 8'b00001110; // 3717 :  14 - 0xe
      12'hE86: dout <= 8'b00111111; // 3718 :  63 - 0x3f
      12'hE87: dout <= 8'b00111001; // 3719 :  57 - 0x39
      12'hE88: dout <= 8'b01110000; // 3720 : 112 - 0x70 -- Background 0xd1
      12'hE89: dout <= 8'b01111000; // 3721 : 120 - 0x78
      12'hE8A: dout <= 8'b00111111; // 3722 :  63 - 0x3f
      12'hE8B: dout <= 8'b00111111; // 3723 :  63 - 0x3f
      12'hE8C: dout <= 8'b00000011; // 3724 :   3 - 0x3
      12'hE8D: dout <= 8'b00001100; // 3725 :  12 - 0xc
      12'hE8E: dout <= 8'b00001110; // 3726 :  14 - 0xe
      12'hE8F: dout <= 8'b00000000; // 3727 :   0 - 0x0
      12'hE90: dout <= 8'b00000000; // 3728 :   0 - 0x0 -- Background 0xd2
      12'hE91: dout <= 8'b00000000; // 3729 :   0 - 0x0
      12'hE92: dout <= 8'b00000000; // 3730 :   0 - 0x0
      12'hE93: dout <= 8'b00001000; // 3731 :   8 - 0x8
      12'hE94: dout <= 8'b11011000; // 3732 : 216 - 0xd8
      12'hE95: dout <= 8'b11111100; // 3733 : 252 - 0xfc
      12'hE96: dout <= 8'b11111100; // 3734 : 252 - 0xfc
      12'hE97: dout <= 8'b10011100; // 3735 : 156 - 0x9c
      12'hE98: dout <= 8'b00001100; // 3736 :  12 - 0xc -- Background 0xd3
      12'hE99: dout <= 8'b10011100; // 3737 : 156 - 0x9c
      12'hE9A: dout <= 8'b11111000; // 3738 : 248 - 0xf8
      12'hE9B: dout <= 8'b01111000; // 3739 : 120 - 0x78
      12'hE9C: dout <= 8'b10001000; // 3740 : 136 - 0x88
      12'hE9D: dout <= 8'b00110000; // 3741 :  48 - 0x30
      12'hE9E: dout <= 8'b00111000; // 3742 :  56 - 0x38
      12'hE9F: dout <= 8'b00000000; // 3743 :   0 - 0x0
      12'hEA0: dout <= 8'b00000000; // 3744 :   0 - 0x0 -- Background 0xd4
      12'hEA1: dout <= 8'b00000000; // 3745 :   0 - 0x0
      12'hEA2: dout <= 8'b00000000; // 3746 :   0 - 0x0
      12'hEA3: dout <= 8'b00000000; // 3747 :   0 - 0x0
      12'hEA4: dout <= 8'b00000001; // 3748 :   1 - 0x1
      12'hEA5: dout <= 8'b00001011; // 3749 :  11 - 0xb
      12'hEA6: dout <= 8'b00011111; // 3750 :  31 - 0x1f
      12'hEA7: dout <= 8'b00111001; // 3751 :  57 - 0x39
      12'hEA8: dout <= 8'b01110000; // 3752 : 112 - 0x70 -- Background 0xd5
      12'hEA9: dout <= 8'b01111000; // 3753 : 120 - 0x78
      12'hEAA: dout <= 8'b00111111; // 3754 :  63 - 0x3f
      12'hEAB: dout <= 8'b00111111; // 3755 :  63 - 0x3f
      12'hEAC: dout <= 8'b00000011; // 3756 :   3 - 0x3
      12'hEAD: dout <= 8'b00111000; // 3757 :  56 - 0x38
      12'hEAE: dout <= 8'b00011100; // 3758 :  28 - 0x1c
      12'hEAF: dout <= 8'b00000000; // 3759 :   0 - 0x0
      12'hEB0: dout <= 8'b00000000; // 3760 :   0 - 0x0 -- Background 0xd6
      12'hEB1: dout <= 8'b00000000; // 3761 :   0 - 0x0
      12'hEB2: dout <= 8'b00000000; // 3762 :   0 - 0x0
      12'hEB3: dout <= 8'b11000000; // 3763 : 192 - 0xc0
      12'hEB4: dout <= 8'b11001000; // 3764 : 200 - 0xc8
      12'hEB5: dout <= 8'b11111000; // 3765 : 248 - 0xf8
      12'hEB6: dout <= 8'b11111100; // 3766 : 252 - 0xfc
      12'hEB7: dout <= 8'b10011100; // 3767 : 156 - 0x9c
      12'hEB8: dout <= 8'b00001100; // 3768 :  12 - 0xc -- Background 0xd7
      12'hEB9: dout <= 8'b10011100; // 3769 : 156 - 0x9c
      12'hEBA: dout <= 8'b11111000; // 3770 : 248 - 0xf8
      12'hEBB: dout <= 8'b01111000; // 3771 : 120 - 0x78
      12'hEBC: dout <= 8'b11100010; // 3772 : 226 - 0xe2
      12'hEBD: dout <= 8'b00011110; // 3773 :  30 - 0x1e
      12'hEBE: dout <= 8'b00001100; // 3774 :  12 - 0xc
      12'hEBF: dout <= 8'b00000000; // 3775 :   0 - 0x0
      12'hEC0: dout <= 8'b00000000; // 3776 :   0 - 0x0 -- Background 0xd8
      12'hEC1: dout <= 8'b00110000; // 3777 :  48 - 0x30
      12'hEC2: dout <= 8'b00111100; // 3778 :  60 - 0x3c
      12'hEC3: dout <= 8'b01111100; // 3779 : 124 - 0x7c
      12'hEC4: dout <= 8'b01111100; // 3780 : 124 - 0x7c
      12'hEC5: dout <= 8'b00111110; // 3781 :  62 - 0x3e
      12'hEC6: dout <= 8'b00011100; // 3782 :  28 - 0x1c
      12'hEC7: dout <= 8'b00000000; // 3783 :   0 - 0x0
      12'hEC8: dout <= 8'b00000000; // 3784 :   0 - 0x0 -- Background 0xd9
      12'hEC9: dout <= 8'b00001110; // 3785 :  14 - 0xe
      12'hECA: dout <= 8'b00111110; // 3786 :  62 - 0x3e
      12'hECB: dout <= 8'b01111110; // 3787 : 126 - 0x7e
      12'hECC: dout <= 8'b01111110; // 3788 : 126 - 0x7e
      12'hECD: dout <= 8'b00111100; // 3789 :  60 - 0x3c
      12'hECE: dout <= 8'b00001100; // 3790 :  12 - 0xc
      12'hECF: dout <= 8'b00000000; // 3791 :   0 - 0x0
      12'hED0: dout <= 8'b00000000; // 3792 :   0 - 0x0 -- Background 0xda
      12'hED1: dout <= 8'b00100000; // 3793 :  32 - 0x20
      12'hED2: dout <= 8'b01111110; // 3794 : 126 - 0x7e
      12'hED3: dout <= 8'b01111110; // 3795 : 126 - 0x7e
      12'hED4: dout <= 8'b01111110; // 3796 : 126 - 0x7e
      12'hED5: dout <= 8'b00111100; // 3797 :  60 - 0x3c
      12'hED6: dout <= 8'b00111000; // 3798 :  56 - 0x38
      12'hED7: dout <= 8'b00000000; // 3799 :   0 - 0x0
      12'hED8: dout <= 8'b00000000; // 3800 :   0 - 0x0 -- Background 0xdb
      12'hED9: dout <= 8'b00011100; // 3801 :  28 - 0x1c
      12'hEDA: dout <= 8'b00111110; // 3802 :  62 - 0x3e
      12'hEDB: dout <= 8'b01111110; // 3803 : 126 - 0x7e
      12'hEDC: dout <= 8'b01111110; // 3804 : 126 - 0x7e
      12'hEDD: dout <= 8'b00111100; // 3805 :  60 - 0x3c
      12'hEDE: dout <= 8'b00010000; // 3806 :  16 - 0x10
      12'hEDF: dout <= 8'b00000000; // 3807 :   0 - 0x0
      12'hEE0: dout <= 8'b00000000; // 3808 :   0 - 0x0 -- Background 0xdc
      12'hEE1: dout <= 8'b00000000; // 3809 :   0 - 0x0
      12'hEE2: dout <= 8'b00000000; // 3810 :   0 - 0x0
      12'hEE3: dout <= 8'b00000001; // 3811 :   1 - 0x1
      12'hEE4: dout <= 8'b00000011; // 3812 :   3 - 0x3
      12'hEE5: dout <= 8'b00000001; // 3813 :   1 - 0x1
      12'hEE6: dout <= 8'b00000001; // 3814 :   1 - 0x1
      12'hEE7: dout <= 8'b00001111; // 3815 :  15 - 0xf
      12'hEE8: dout <= 8'b00000111; // 3816 :   7 - 0x7 -- Background 0xdd
      12'hEE9: dout <= 8'b00000111; // 3817 :   7 - 0x7
      12'hEEA: dout <= 8'b00000111; // 3818 :   7 - 0x7
      12'hEEB: dout <= 8'b00011111; // 3819 :  31 - 0x1f
      12'hEEC: dout <= 8'b00001111; // 3820 :  15 - 0xf
      12'hEED: dout <= 8'b00000111; // 3821 :   7 - 0x7
      12'hEEE: dout <= 8'b00000011; // 3822 :   3 - 0x3
      12'hEEF: dout <= 8'b00000000; // 3823 :   0 - 0x0
      12'hEF0: dout <= 8'b00000000; // 3824 :   0 - 0x0 -- Background 0xde
      12'hEF1: dout <= 8'b00000000; // 3825 :   0 - 0x0
      12'hEF2: dout <= 8'b00000000; // 3826 :   0 - 0x0
      12'hEF3: dout <= 8'b00000000; // 3827 :   0 - 0x0
      12'hEF4: dout <= 8'b10000000; // 3828 : 128 - 0x80
      12'hEF5: dout <= 8'b10000000; // 3829 : 128 - 0x80
      12'hEF6: dout <= 8'b10010000; // 3830 : 144 - 0x90
      12'hEF7: dout <= 8'b11110000; // 3831 : 240 - 0xf0
      12'hEF8: dout <= 8'b11100000; // 3832 : 224 - 0xe0 -- Background 0xdf
      12'hEF9: dout <= 8'b11100000; // 3833 : 224 - 0xe0
      12'hEFA: dout <= 8'b11110000; // 3834 : 240 - 0xf0
      12'hEFB: dout <= 8'b11110000; // 3835 : 240 - 0xf0
      12'hEFC: dout <= 8'b11100000; // 3836 : 224 - 0xe0
      12'hEFD: dout <= 8'b11000000; // 3837 : 192 - 0xc0
      12'hEFE: dout <= 8'b11000000; // 3838 : 192 - 0xc0
      12'hEFF: dout <= 8'b00000000; // 3839 :   0 - 0x0
      12'hF00: dout <= 8'b00001111; // 3840 :  15 - 0xf -- Background 0xe0
      12'hF01: dout <= 8'b00011111; // 3841 :  31 - 0x1f
      12'hF02: dout <= 8'b00011111; // 3842 :  31 - 0x1f
      12'hF03: dout <= 8'b00111111; // 3843 :  63 - 0x3f
      12'hF04: dout <= 8'b01111111; // 3844 : 127 - 0x7f
      12'hF05: dout <= 8'b11111111; // 3845 : 255 - 0xff
      12'hF06: dout <= 8'b11111111; // 3846 : 255 - 0xff
      12'hF07: dout <= 8'b11111111; // 3847 : 255 - 0xff
      12'hF08: dout <= 8'b11111111; // 3848 : 255 - 0xff -- Background 0xe1
      12'hF09: dout <= 8'b11111111; // 3849 : 255 - 0xff
      12'hF0A: dout <= 8'b01111111; // 3850 : 127 - 0x7f
      12'hF0B: dout <= 8'b00111111; // 3851 :  63 - 0x3f
      12'hF0C: dout <= 8'b00111111; // 3852 :  63 - 0x3f
      12'hF0D: dout <= 8'b00011111; // 3853 :  31 - 0x1f
      12'hF0E: dout <= 8'b00001111; // 3854 :  15 - 0xf
      12'hF0F: dout <= 8'b00000111; // 3855 :   7 - 0x7
      12'hF10: dout <= 8'b11111110; // 3856 : 254 - 0xfe -- Background 0xe2
      12'hF11: dout <= 8'b11111111; // 3857 : 255 - 0xff
      12'hF12: dout <= 8'b11111111; // 3858 : 255 - 0xff
      12'hF13: dout <= 8'b00001111; // 3859 :  15 - 0xf
      12'hF14: dout <= 8'b10111111; // 3860 : 191 - 0xbf
      12'hF15: dout <= 8'b10100011; // 3861 : 163 - 0xa3
      12'hF16: dout <= 8'b11110111; // 3862 : 247 - 0xf7
      12'hF17: dout <= 8'b11110111; // 3863 : 247 - 0xf7
      12'hF18: dout <= 8'b11111111; // 3864 : 255 - 0xff -- Background 0xe3
      12'hF19: dout <= 8'b11111111; // 3865 : 255 - 0xff
      12'hF1A: dout <= 8'b00111111; // 3866 :  63 - 0x3f
      12'hF1B: dout <= 8'b00011111; // 3867 :  31 - 0x1f
      12'hF1C: dout <= 8'b11111110; // 3868 : 254 - 0xfe
      12'hF1D: dout <= 8'b11111100; // 3869 : 252 - 0xfc
      12'hF1E: dout <= 8'b11111000; // 3870 : 248 - 0xf8
      12'hF1F: dout <= 8'b11110000; // 3871 : 240 - 0xf0
      12'hF20: dout <= 8'b00001111; // 3872 :  15 - 0xf -- Background 0xe4
      12'hF21: dout <= 8'b00011111; // 3873 :  31 - 0x1f
      12'hF22: dout <= 8'b00011111; // 3874 :  31 - 0x1f
      12'hF23: dout <= 8'b00111111; // 3875 :  63 - 0x3f
      12'hF24: dout <= 8'b01111111; // 3876 : 127 - 0x7f
      12'hF25: dout <= 8'b11111111; // 3877 : 255 - 0xff
      12'hF26: dout <= 8'b11111111; // 3878 : 255 - 0xff
      12'hF27: dout <= 8'b11111111; // 3879 : 255 - 0xff
      12'hF28: dout <= 8'b11111111; // 3880 : 255 - 0xff -- Background 0xe5
      12'hF29: dout <= 8'b11111111; // 3881 : 255 - 0xff
      12'hF2A: dout <= 8'b01111110; // 3882 : 126 - 0x7e
      12'hF2B: dout <= 8'b00111111; // 3883 :  63 - 0x3f
      12'hF2C: dout <= 8'b00111111; // 3884 :  63 - 0x3f
      12'hF2D: dout <= 8'b00011111; // 3885 :  31 - 0x1f
      12'hF2E: dout <= 8'b00001111; // 3886 :  15 - 0xf
      12'hF2F: dout <= 8'b00000111; // 3887 :   7 - 0x7
      12'hF30: dout <= 8'b11111110; // 3888 : 254 - 0xfe -- Background 0xe6
      12'hF31: dout <= 8'b11111111; // 3889 : 255 - 0xff
      12'hF32: dout <= 8'b11111111; // 3890 : 255 - 0xff
      12'hF33: dout <= 8'b11100011; // 3891 : 227 - 0xe3
      12'hF34: dout <= 8'b00010111; // 3892 :  23 - 0x17
      12'hF35: dout <= 8'b10110111; // 3893 : 183 - 0xb7
      12'hF36: dout <= 8'b10111111; // 3894 : 191 - 0xbf
      12'hF37: dout <= 8'b11111111; // 3895 : 255 - 0xff
      12'hF38: dout <= 8'b11111111; // 3896 : 255 - 0xff -- Background 0xe7
      12'hF39: dout <= 8'b11111111; // 3897 : 255 - 0xff
      12'hF3A: dout <= 8'b00111111; // 3898 :  63 - 0x3f
      12'hF3B: dout <= 8'b00001111; // 3899 :  15 - 0xf
      12'hF3C: dout <= 8'b00001110; // 3900 :  14 - 0xe
      12'hF3D: dout <= 8'b11111100; // 3901 : 252 - 0xfc
      12'hF3E: dout <= 8'b11111000; // 3902 : 248 - 0xf8
      12'hF3F: dout <= 8'b11110000; // 3903 : 240 - 0xf0
      12'hF40: dout <= 8'b00000000; // 3904 :   0 - 0x0 -- Background 0xe8
      12'hF41: dout <= 8'b00000101; // 3905 :   5 - 0x5
      12'hF42: dout <= 8'b00000111; // 3906 :   7 - 0x7
      12'hF43: dout <= 8'b00000011; // 3907 :   3 - 0x3
      12'hF44: dout <= 8'b00000000; // 3908 :   0 - 0x0
      12'hF45: dout <= 8'b00000000; // 3909 :   0 - 0x0
      12'hF46: dout <= 8'b00000000; // 3910 :   0 - 0x0
      12'hF47: dout <= 8'b00000000; // 3911 :   0 - 0x0
      12'hF48: dout <= 8'b00000000; // 3912 :   0 - 0x0 -- Background 0xe9
      12'hF49: dout <= 8'b00000000; // 3913 :   0 - 0x0
      12'hF4A: dout <= 8'b00000000; // 3914 :   0 - 0x0
      12'hF4B: dout <= 8'b00000000; // 3915 :   0 - 0x0
      12'hF4C: dout <= 8'b00000000; // 3916 :   0 - 0x0
      12'hF4D: dout <= 8'b00000000; // 3917 :   0 - 0x0
      12'hF4E: dout <= 8'b00000000; // 3918 :   0 - 0x0
      12'hF4F: dout <= 8'b00000000; // 3919 :   0 - 0x0
      12'hF50: dout <= 8'b00000011; // 3920 :   3 - 0x3 -- Background 0xea
      12'hF51: dout <= 8'b10011110; // 3921 : 158 - 0x9e
      12'hF52: dout <= 8'b00001110; // 3922 :  14 - 0xe
      12'hF53: dout <= 8'b00000000; // 3923 :   0 - 0x0
      12'hF54: dout <= 8'b00000000; // 3924 :   0 - 0x0
      12'hF55: dout <= 8'b00000000; // 3925 :   0 - 0x0
      12'hF56: dout <= 8'b00000000; // 3926 :   0 - 0x0
      12'hF57: dout <= 8'b00000000; // 3927 :   0 - 0x0
      12'hF58: dout <= 8'b00000000; // 3928 :   0 - 0x0 -- Background 0xeb
      12'hF59: dout <= 8'b00000000; // 3929 :   0 - 0x0
      12'hF5A: dout <= 8'b00000000; // 3930 :   0 - 0x0
      12'hF5B: dout <= 8'b00000000; // 3931 :   0 - 0x0
      12'hF5C: dout <= 8'b00000000; // 3932 :   0 - 0x0
      12'hF5D: dout <= 8'b00000000; // 3933 :   0 - 0x0
      12'hF5E: dout <= 8'b00000000; // 3934 :   0 - 0x0
      12'hF5F: dout <= 8'b00000000; // 3935 :   0 - 0x0
      12'hF60: dout <= 8'b00000000; // 3936 :   0 - 0x0 -- Background 0xec
      12'hF61: dout <= 8'b00000000; // 3937 :   0 - 0x0
      12'hF62: dout <= 8'b00000000; // 3938 :   0 - 0x0
      12'hF63: dout <= 8'b00000000; // 3939 :   0 - 0x0
      12'hF64: dout <= 8'b00000100; // 3940 :   4 - 0x4
      12'hF65: dout <= 8'b00001110; // 3941 :  14 - 0xe
      12'hF66: dout <= 8'b00001111; // 3942 :  15 - 0xf
      12'hF67: dout <= 8'b00001011; // 3943 :  11 - 0xb
      12'hF68: dout <= 8'b00001111; // 3944 :  15 - 0xf -- Background 0xed
      12'hF69: dout <= 8'b00001100; // 3945 :  12 - 0xc
      12'hF6A: dout <= 8'b00001111; // 3946 :  15 - 0xf
      12'hF6B: dout <= 8'b00001111; // 3947 :  15 - 0xf
      12'hF6C: dout <= 8'b00000000; // 3948 :   0 - 0x0
      12'hF6D: dout <= 8'b01111111; // 3949 : 127 - 0x7f
      12'hF6E: dout <= 8'b11010101; // 3950 : 213 - 0xd5
      12'hF6F: dout <= 8'b01111111; // 3951 : 127 - 0x7f
      12'hF70: dout <= 8'b00000000; // 3952 :   0 - 0x0 -- Background 0xee
      12'hF71: dout <= 8'b00000000; // 3953 :   0 - 0x0
      12'hF72: dout <= 8'b00000000; // 3954 :   0 - 0x0
      12'hF73: dout <= 8'b00000000; // 3955 :   0 - 0x0
      12'hF74: dout <= 8'b00100000; // 3956 :  32 - 0x20
      12'hF75: dout <= 8'b01110000; // 3957 : 112 - 0x70
      12'hF76: dout <= 8'b11110000; // 3958 : 240 - 0xf0
      12'hF77: dout <= 8'b11100000; // 3959 : 224 - 0xe0
      12'hF78: dout <= 8'b11110000; // 3960 : 240 - 0xf0 -- Background 0xef
      12'hF79: dout <= 8'b00110000; // 3961 :  48 - 0x30
      12'hF7A: dout <= 8'b11110000; // 3962 : 240 - 0xf0
      12'hF7B: dout <= 8'b11110000; // 3963 : 240 - 0xf0
      12'hF7C: dout <= 8'b00000000; // 3964 :   0 - 0x0
      12'hF7D: dout <= 8'b11111110; // 3965 : 254 - 0xfe
      12'hF7E: dout <= 8'b01010101; // 3966 :  85 - 0x55
      12'hF7F: dout <= 8'b11111110; // 3967 : 254 - 0xfe
      12'hF80: dout <= 8'b00000000; // 3968 :   0 - 0x0 -- Background 0xf0
      12'hF81: dout <= 8'b00000000; // 3969 :   0 - 0x0
      12'hF82: dout <= 8'b00000000; // 3970 :   0 - 0x0
      12'hF83: dout <= 8'b00000000; // 3971 :   0 - 0x0
      12'hF84: dout <= 8'b00000100; // 3972 :   4 - 0x4
      12'hF85: dout <= 8'b00001110; // 3973 :  14 - 0xe
      12'hF86: dout <= 8'b00001111; // 3974 :  15 - 0xf
      12'hF87: dout <= 8'b00001011; // 3975 :  11 - 0xb
      12'hF88: dout <= 8'b00001111; // 3976 :  15 - 0xf -- Background 0xf1
      12'hF89: dout <= 8'b00001100; // 3977 :  12 - 0xc
      12'hF8A: dout <= 8'b00001111; // 3978 :  15 - 0xf
      12'hF8B: dout <= 8'b00001111; // 3979 :  15 - 0xf
      12'hF8C: dout <= 8'b00000000; // 3980 :   0 - 0x0
      12'hF8D: dout <= 8'b01111111; // 3981 : 127 - 0x7f
      12'hF8E: dout <= 8'b10101010; // 3982 : 170 - 0xaa
      12'hF8F: dout <= 8'b01111111; // 3983 : 127 - 0x7f
      12'hF90: dout <= 8'b00000000; // 3984 :   0 - 0x0 -- Background 0xf2
      12'hF91: dout <= 8'b00000000; // 3985 :   0 - 0x0
      12'hF92: dout <= 8'b00000000; // 3986 :   0 - 0x0
      12'hF93: dout <= 8'b00000000; // 3987 :   0 - 0x0
      12'hF94: dout <= 8'b00100000; // 3988 :  32 - 0x20
      12'hF95: dout <= 8'b01110000; // 3989 : 112 - 0x70
      12'hF96: dout <= 8'b11110000; // 3990 : 240 - 0xf0
      12'hF97: dout <= 8'b11100000; // 3991 : 224 - 0xe0
      12'hF98: dout <= 8'b11110000; // 3992 : 240 - 0xf0 -- Background 0xf3
      12'hF99: dout <= 8'b00110000; // 3993 :  48 - 0x30
      12'hF9A: dout <= 8'b11110000; // 3994 : 240 - 0xf0
      12'hF9B: dout <= 8'b11110000; // 3995 : 240 - 0xf0
      12'hF9C: dout <= 8'b00000000; // 3996 :   0 - 0x0
      12'hF9D: dout <= 8'b11111110; // 3997 : 254 - 0xfe
      12'hF9E: dout <= 8'b10101011; // 3998 : 171 - 0xab
      12'hF9F: dout <= 8'b11111110; // 3999 : 254 - 0xfe
      12'hFA0: dout <= 8'b00000000; // 4000 :   0 - 0x0 -- Background 0xf4
      12'hFA1: dout <= 8'b00010101; // 4001 :  21 - 0x15
      12'hFA2: dout <= 8'b00001010; // 4002 :  10 - 0xa
      12'hFA3: dout <= 8'b00000101; // 4003 :   5 - 0x5
      12'hFA4: dout <= 8'b00000010; // 4004 :   2 - 0x2
      12'hFA5: dout <= 8'b00000101; // 4005 :   5 - 0x5
      12'hFA6: dout <= 8'b00000111; // 4006 :   7 - 0x7
      12'hFA7: dout <= 8'b00000111; // 4007 :   7 - 0x7
      12'hFA8: dout <= 8'b00111100; // 4008 :  60 - 0x3c -- Background 0xf5
      12'hFA9: dout <= 8'b01111011; // 4009 : 123 - 0x7b
      12'hFAA: dout <= 8'b01111011; // 4010 : 123 - 0x7b
      12'hFAB: dout <= 8'b01111111; // 4011 : 127 - 0x7f
      12'hFAC: dout <= 8'b01111110; // 4012 : 126 - 0x7e
      12'hFAD: dout <= 8'b01111111; // 4013 : 127 - 0x7f
      12'hFAE: dout <= 8'b00111110; // 4014 :  62 - 0x3e
      12'hFAF: dout <= 8'b00000000; // 4015 :   0 - 0x0
      12'hFB0: dout <= 8'b00000000; // 4016 :   0 - 0x0 -- Background 0xf6
      12'hFB1: dout <= 8'b01010000; // 4017 :  80 - 0x50
      12'hFB2: dout <= 8'b10100000; // 4018 : 160 - 0xa0
      12'hFB3: dout <= 8'b01000000; // 4019 :  64 - 0x40
      12'hFB4: dout <= 8'b10100000; // 4020 : 160 - 0xa0
      12'hFB5: dout <= 8'b01000000; // 4021 :  64 - 0x40
      12'hFB6: dout <= 8'b11100000; // 4022 : 224 - 0xe0
      12'hFB7: dout <= 8'b11100000; // 4023 : 224 - 0xe0
      12'hFB8: dout <= 8'b01111000; // 4024 : 120 - 0x78 -- Background 0xf7
      12'hFB9: dout <= 8'b10111100; // 4025 : 188 - 0xbc
      12'hFBA: dout <= 8'b10111000; // 4026 : 184 - 0xb8
      12'hFBB: dout <= 8'b10111110; // 4027 : 190 - 0xbe
      12'hFBC: dout <= 8'b01111100; // 4028 : 124 - 0x7c
      12'hFBD: dout <= 8'b11111110; // 4029 : 254 - 0xfe
      12'hFBE: dout <= 8'b01111000; // 4030 : 120 - 0x78
      12'hFBF: dout <= 8'b00000000; // 4031 :   0 - 0x0
      12'hFC0: dout <= 8'b00000011; // 4032 :   3 - 0x3 -- Background 0xf8
      12'hFC1: dout <= 8'b00000011; // 4033 :   3 - 0x3
      12'hFC2: dout <= 8'b00000000; // 4034 :   0 - 0x0
      12'hFC3: dout <= 8'b00000011; // 4035 :   3 - 0x3
      12'hFC4: dout <= 8'b00000111; // 4036 :   7 - 0x7
      12'hFC5: dout <= 8'b00000110; // 4037 :   6 - 0x6
      12'hFC6: dout <= 8'b00000111; // 4038 :   7 - 0x7
      12'hFC7: dout <= 8'b00000000; // 4039 :   0 - 0x0
      12'hFC8: dout <= 8'b00000000; // 4040 :   0 - 0x0 -- Background 0xf9
      12'hFC9: dout <= 8'b00011111; // 4041 :  31 - 0x1f
      12'hFCA: dout <= 8'b00011111; // 4042 :  31 - 0x1f
      12'hFCB: dout <= 8'b00001111; // 4043 :  15 - 0xf
      12'hFCC: dout <= 8'b00000011; // 4044 :   3 - 0x3
      12'hFCD: dout <= 8'b00000000; // 4045 :   0 - 0x0
      12'hFCE: dout <= 8'b00000000; // 4046 :   0 - 0x0
      12'hFCF: dout <= 8'b00000000; // 4047 :   0 - 0x0
      12'hFD0: dout <= 8'b11100000; // 4048 : 224 - 0xe0 -- Background 0xfa
      12'hFD1: dout <= 8'b11100000; // 4049 : 224 - 0xe0
      12'hFD2: dout <= 8'b00000000; // 4050 :   0 - 0x0
      12'hFD3: dout <= 8'b00110000; // 4051 :  48 - 0x30
      12'hFD4: dout <= 8'b01110000; // 4052 : 112 - 0x70
      12'hFD5: dout <= 8'b01100000; // 4053 :  96 - 0x60
      12'hFD6: dout <= 8'b01110000; // 4054 : 112 - 0x70
      12'hFD7: dout <= 8'b00000000; // 4055 :   0 - 0x0
      12'hFD8: dout <= 8'b00000000; // 4056 :   0 - 0x0 -- Background 0xfb
      12'hFD9: dout <= 8'b11111000; // 4057 : 248 - 0xf8
      12'hFDA: dout <= 8'b11111000; // 4058 : 248 - 0xf8
      12'hFDB: dout <= 8'b11110000; // 4059 : 240 - 0xf0
      12'hFDC: dout <= 8'b11000000; // 4060 : 192 - 0xc0
      12'hFDD: dout <= 8'b00000000; // 4061 :   0 - 0x0
      12'hFDE: dout <= 8'b00000000; // 4062 :   0 - 0x0
      12'hFDF: dout <= 8'b00000000; // 4063 :   0 - 0x0
      12'hFE0: dout <= 8'b00111000; // 4064 :  56 - 0x38 -- Background 0xfc
      12'hFE1: dout <= 8'b00111000; // 4065 :  56 - 0x38
      12'hFE2: dout <= 8'b00000000; // 4066 :   0 - 0x0
      12'hFE3: dout <= 8'b01111100; // 4067 : 124 - 0x7c
      12'hFE4: dout <= 8'b00000000; // 4068 :   0 - 0x0
      12'hFE5: dout <= 8'b00111000; // 4069 :  56 - 0x38
      12'hFE6: dout <= 8'b00111000; // 4070 :  56 - 0x38
      12'hFE7: dout <= 8'b01111100; // 4071 : 124 - 0x7c
      12'hFE8: dout <= 8'b01111100; // 4072 : 124 - 0x7c -- Background 0xfd
      12'hFE9: dout <= 8'b01111100; // 4073 : 124 - 0x7c
      12'hFEA: dout <= 8'b01111100; // 4074 : 124 - 0x7c
      12'hFEB: dout <= 8'b00111000; // 4075 :  56 - 0x38
      12'hFEC: dout <= 8'b00000000; // 4076 :   0 - 0x0
      12'hFED: dout <= 8'b01111100; // 4077 : 124 - 0x7c
      12'hFEE: dout <= 8'b01111100; // 4078 : 124 - 0x7c
      12'hFEF: dout <= 8'b00000000; // 4079 :   0 - 0x0
      12'hFF0: dout <= 8'b00000000; // 4080 :   0 - 0x0 -- Background 0xfe
      12'hFF1: dout <= 8'b00000000; // 4081 :   0 - 0x0
      12'hFF2: dout <= 8'b00010001; // 4082 :  17 - 0x11
      12'hFF3: dout <= 8'b11010111; // 4083 : 215 - 0xd7
      12'hFF4: dout <= 8'b11010111; // 4084 : 215 - 0xd7
      12'hFF5: dout <= 8'b11010111; // 4085 : 215 - 0xd7
      12'hFF6: dout <= 8'b00010001; // 4086 :  17 - 0x11
      12'hFF7: dout <= 8'b00000000; // 4087 :   0 - 0x0
      12'hFF8: dout <= 8'b00000000; // 4088 :   0 - 0x0 -- Background 0xff
      12'hFF9: dout <= 8'b00000000; // 4089 :   0 - 0x0
      12'hFFA: dout <= 8'b11100110; // 4090 : 230 - 0xe6
      12'hFFB: dout <= 8'b11110110; // 4091 : 246 - 0xf6
      12'hFFC: dout <= 8'b11110110; // 4092 : 246 - 0xf6
      12'hFFD: dout <= 8'b11110110; // 4093 : 246 - 0xf6
      12'hFFE: dout <= 8'b11100110; // 4094 : 230 - 0xe6
      12'hFFF: dout <= 8'b00000000; // 4095 :   0 - 0x0
    endcase
  end

endmodule
