//---- Felipe Machado -------------------------------
//---- Area de Tecnologia Electronica ---------------
//---- Universidad Rey Juan Carlos ------------------
//---- https://github.com/felipe-m ------------------
//---------------------------------------------------
//---- Autcmatically generated verilog ROM blockfrom a VHDL file----
//  Original VHDL file name: rom_red_square_80x60_rgb_8b.vhd
//  Constant VHDL name: filaimg
//  Memory with blocking assignments (=)

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module rom_red_square_80x60_rgb_8b
  (
     //input     clk,   // clock
     input      [13-1:0] addr,  //4800 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


//  Memory without clock

  always @(*)
  begin
    case(addr)
            //"RRRGGGBB"
      13'h0: dout = 8'b10111011;
      13'h1: dout = 8'b10111011;
      13'h2: dout = 8'b10111011;
      13'h3: dout = 8'b10111011;
      13'h4: dout = 8'b10111011;
      13'h5: dout = 8'b10111011;
      13'h6: dout = 8'b10111011;
      13'h7: dout = 8'b10111011;
      13'h8: dout = 8'b10111011;
      13'h9: dout = 8'b10111011;
      13'hA: dout = 8'b10111011;
      13'hB: dout = 8'b10111011;
      13'hC: dout = 8'b10111011;
      13'hD: dout = 8'b10111011;
      13'hE: dout = 8'b10111011;
      13'hF: dout = 8'b10111011;
      13'h10: dout = 8'b10111011;
      13'h11: dout = 8'b10111011;
      13'h12: dout = 8'b10111011;
      13'h13: dout = 8'b10111011;
      13'h14: dout = 8'b10111011;
      13'h15: dout = 8'b10111011;
      13'h16: dout = 8'b10111011;
      13'h17: dout = 8'b10111011;
      13'h18: dout = 8'b10111011;
      13'h19: dout = 8'b10111011;
      13'h1A: dout = 8'b10111011;
      13'h1B: dout = 8'b10111011;
      13'h1C: dout = 8'b10111011;
      13'h1D: dout = 8'b10111011;
      13'h1E: dout = 8'b10111011;
      13'h1F: dout = 8'b10111011;
      13'h20: dout = 8'b10111011;
      13'h21: dout = 8'b10111011;
      13'h22: dout = 8'b10111011;
      13'h23: dout = 8'b10111011;
      13'h24: dout = 8'b10111011;
      13'h25: dout = 8'b10111011;
      13'h26: dout = 8'b10111011;
      13'h27: dout = 8'b10111011;
      13'h28: dout = 8'b10111011;
      13'h29: dout = 8'b10111011;
      13'h2A: dout = 8'b10111011;
      13'h2B: dout = 8'b10111011;
      13'h2C: dout = 8'b10111011;
      13'h2D: dout = 8'b10111011;
      13'h2E: dout = 8'b10111011;
      13'h2F: dout = 8'b10111011;
      13'h30: dout = 8'b10111011;
      13'h31: dout = 8'b10111011;
      13'h32: dout = 8'b10111011;
      13'h33: dout = 8'b10111011;
      13'h34: dout = 8'b10111011;
      13'h35: dout = 8'b10111011;
      13'h36: dout = 8'b10111011;
      13'h37: dout = 8'b10111011;
      13'h38: dout = 8'b10111011;
      13'h39: dout = 8'b10111011;
      13'h3A: dout = 8'b10111011;
      13'h3B: dout = 8'b10111011;
      13'h3C: dout = 8'b10111011;
      13'h3D: dout = 8'b10111011;
      13'h3E: dout = 8'b10111011;
      13'h3F: dout = 8'b10111011;
      13'h40: dout = 8'b10111011;
      13'h41: dout = 8'b10111011;
      13'h42: dout = 8'b10111011;
      13'h43: dout = 8'b10111011;
      13'h44: dout = 8'b10111011;
      13'h45: dout = 8'b10111011;
      13'h46: dout = 8'b10111011;
      13'h47: dout = 8'b10111011;
      13'h48: dout = 8'b10111011;
      13'h49: dout = 8'b10111011;
      13'h4A: dout = 8'b10111011;
      13'h4B: dout = 8'b10111011;
      13'h4C: dout = 8'b10111011;
      13'h4D: dout = 8'b10111011;
      13'h4E: dout = 8'b10111011;
      13'h4F: dout = 8'b10111011;
      13'h50: dout = 8'b10111011;
      13'h51: dout = 8'b10111011;
      13'h52: dout = 8'b10111011;
      13'h53: dout = 8'b10111011;
      13'h54: dout = 8'b10111011;
      13'h55: dout = 8'b10111011;
      13'h56: dout = 8'b10111011;
      13'h57: dout = 8'b10111011;
      13'h58: dout = 8'b10111011;
      13'h59: dout = 8'b10111011;
      13'h5A: dout = 8'b10111011;
      13'h5B: dout = 8'b10111011;
      13'h5C: dout = 8'b10111011;
      13'h5D: dout = 8'b10111011;
      13'h5E: dout = 8'b10111011;
      13'h5F: dout = 8'b10111011;
      13'h60: dout = 8'b10111011;
      13'h61: dout = 8'b10111011;
      13'h62: dout = 8'b10111011;
      13'h63: dout = 8'b10111011;
      13'h64: dout = 8'b10111011;
      13'h65: dout = 8'b10111011;
      13'h66: dout = 8'b10111011;
      13'h67: dout = 8'b10111011;
      13'h68: dout = 8'b10111011;
      13'h69: dout = 8'b10111011;
      13'h6A: dout = 8'b10111011;
      13'h6B: dout = 8'b10111011;
      13'h6C: dout = 8'b10111011;
      13'h6D: dout = 8'b10111011;
      13'h6E: dout = 8'b10111011;
      13'h6F: dout = 8'b10111011;
      13'h70: dout = 8'b10111011;
      13'h71: dout = 8'b10111011;
      13'h72: dout = 8'b10111011;
      13'h73: dout = 8'b10111011;
      13'h74: dout = 8'b10111011;
      13'h75: dout = 8'b10111011;
      13'h76: dout = 8'b10111011;
      13'h77: dout = 8'b10111011;
      13'h78: dout = 8'b10111011;
      13'h79: dout = 8'b10111011;
      13'h7A: dout = 8'b10111011;
      13'h7B: dout = 8'b10111011;
      13'h7C: dout = 8'b10111011;
      13'h7D: dout = 8'b10111011;
      13'h7E: dout = 8'b10111011;
      13'h7F: dout = 8'b10111011;
      13'h80: dout = 8'b10111011;
      13'h81: dout = 8'b10111011;
      13'h82: dout = 8'b10111011;
      13'h83: dout = 8'b10111011;
      13'h84: dout = 8'b10111011;
      13'h85: dout = 8'b10111011;
      13'h86: dout = 8'b10111011;
      13'h87: dout = 8'b10111011;
      13'h88: dout = 8'b10111011;
      13'h89: dout = 8'b10111011;
      13'h8A: dout = 8'b10111011;
      13'h8B: dout = 8'b10111011;
      13'h8C: dout = 8'b10111011;
      13'h8D: dout = 8'b10111011;
      13'h8E: dout = 8'b10111011;
      13'h8F: dout = 8'b10111011;
      13'h90: dout = 8'b10111011;
      13'h91: dout = 8'b10111011;
      13'h92: dout = 8'b10111011;
      13'h93: dout = 8'b10111011;
      13'h94: dout = 8'b10111011;
      13'h95: dout = 8'b10111011;
      13'h96: dout = 8'b10111011;
      13'h97: dout = 8'b10111011;
      13'h98: dout = 8'b10111011;
      13'h99: dout = 8'b10111011;
      13'h9A: dout = 8'b10111011;
      13'h9B: dout = 8'b10111011;
      13'h9C: dout = 8'b10111011;
      13'h9D: dout = 8'b10111011;
      13'h9E: dout = 8'b10111011;
      13'h9F: dout = 8'b10111011;
      13'hA0: dout = 8'b10111011;
      13'hA1: dout = 8'b10111011;
      13'hA2: dout = 8'b10111011;
      13'hA3: dout = 8'b10111011;
      13'hA4: dout = 8'b10111011;
      13'hA5: dout = 8'b10111011;
      13'hA6: dout = 8'b10111011;
      13'hA7: dout = 8'b10111011;
      13'hA8: dout = 8'b10111011;
      13'hA9: dout = 8'b10111011;
      13'hAA: dout = 8'b10111011;
      13'hAB: dout = 8'b10111011;
      13'hAC: dout = 8'b10111011;
      13'hAD: dout = 8'b10111011;
      13'hAE: dout = 8'b10111011;
      13'hAF: dout = 8'b10111011;
      13'hB0: dout = 8'b10111011;
      13'hB1: dout = 8'b10111011;
      13'hB2: dout = 8'b10111011;
      13'hB3: dout = 8'b10111011;
      13'hB4: dout = 8'b10111011;
      13'hB5: dout = 8'b10111011;
      13'hB6: dout = 8'b10111011;
      13'hB7: dout = 8'b10111011;
      13'hB8: dout = 8'b10111011;
      13'hB9: dout = 8'b10111011;
      13'hBA: dout = 8'b10111011;
      13'hBB: dout = 8'b10111011;
      13'hBC: dout = 8'b10111011;
      13'hBD: dout = 8'b10111011;
      13'hBE: dout = 8'b10111011;
      13'hBF: dout = 8'b10111011;
      13'hC0: dout = 8'b10111011;
      13'hC1: dout = 8'b10111011;
      13'hC2: dout = 8'b10111011;
      13'hC3: dout = 8'b10111011;
      13'hC4: dout = 8'b10111011;
      13'hC5: dout = 8'b10111011;
      13'hC6: dout = 8'b10111011;
      13'hC7: dout = 8'b10111011;
      13'hC8: dout = 8'b10111011;
      13'hC9: dout = 8'b10111011;
      13'hCA: dout = 8'b10111011;
      13'hCB: dout = 8'b10111011;
      13'hCC: dout = 8'b10111011;
      13'hCD: dout = 8'b10111011;
      13'hCE: dout = 8'b10111011;
      13'hCF: dout = 8'b10111011;
      13'hD0: dout = 8'b10111011;
      13'hD1: dout = 8'b10111011;
      13'hD2: dout = 8'b10111011;
      13'hD3: dout = 8'b10111011;
      13'hD4: dout = 8'b10111011;
      13'hD5: dout = 8'b10111011;
      13'hD6: dout = 8'b10111011;
      13'hD7: dout = 8'b10111011;
      13'hD8: dout = 8'b10111011;
      13'hD9: dout = 8'b10111011;
      13'hDA: dout = 8'b10111011;
      13'hDB: dout = 8'b10111011;
      13'hDC: dout = 8'b10111011;
      13'hDD: dout = 8'b10111011;
      13'hDE: dout = 8'b10111011;
      13'hDF: dout = 8'b10111011;
      13'hE0: dout = 8'b10111011;
      13'hE1: dout = 8'b10111011;
      13'hE2: dout = 8'b10111011;
      13'hE3: dout = 8'b10111011;
      13'hE4: dout = 8'b10111011;
      13'hE5: dout = 8'b10111011;
      13'hE6: dout = 8'b10111011;
      13'hE7: dout = 8'b10111011;
      13'hE8: dout = 8'b10111011;
      13'hE9: dout = 8'b10111011;
      13'hEA: dout = 8'b10111011;
      13'hEB: dout = 8'b10111011;
      13'hEC: dout = 8'b10111011;
      13'hED: dout = 8'b10111011;
      13'hEE: dout = 8'b10111011;
      13'hEF: dout = 8'b10111011;
      13'hF0: dout = 8'b10111011;
      13'hF1: dout = 8'b10111011;
      13'hF2: dout = 8'b10111011;
      13'hF3: dout = 8'b10111011;
      13'hF4: dout = 8'b10111011;
      13'hF5: dout = 8'b10111011;
      13'hF6: dout = 8'b10111011;
      13'hF7: dout = 8'b10111011;
      13'hF8: dout = 8'b10111011;
      13'hF9: dout = 8'b10111011;
      13'hFA: dout = 8'b10111011;
      13'hFB: dout = 8'b10111011;
      13'hFC: dout = 8'b10111011;
      13'hFD: dout = 8'b10111011;
      13'hFE: dout = 8'b10111011;
      13'hFF: dout = 8'b10111011;
      13'h100: dout = 8'b10111011;
      13'h101: dout = 8'b10111011;
      13'h102: dout = 8'b10111011;
      13'h103: dout = 8'b10111011;
      13'h104: dout = 8'b10111011;
      13'h105: dout = 8'b10111011;
      13'h106: dout = 8'b10111011;
      13'h107: dout = 8'b10111011;
      13'h108: dout = 8'b10111011;
      13'h109: dout = 8'b10111011;
      13'h10A: dout = 8'b10111011;
      13'h10B: dout = 8'b10111011;
      13'h10C: dout = 8'b10111011;
      13'h10D: dout = 8'b10111011;
      13'h10E: dout = 8'b10111011;
      13'h10F: dout = 8'b10111011;
      13'h110: dout = 8'b10111011;
      13'h111: dout = 8'b10111011;
      13'h112: dout = 8'b10111011;
      13'h113: dout = 8'b10111011;
      13'h114: dout = 8'b10111011;
      13'h115: dout = 8'b10111011;
      13'h116: dout = 8'b10111011;
      13'h117: dout = 8'b10111011;
      13'h118: dout = 8'b10111011;
      13'h119: dout = 8'b10111011;
      13'h11A: dout = 8'b10111011;
      13'h11B: dout = 8'b10111011;
      13'h11C: dout = 8'b10111011;
      13'h11D: dout = 8'b10111011;
      13'h11E: dout = 8'b10111011;
      13'h11F: dout = 8'b10111011;
      13'h120: dout = 8'b10111011;
      13'h121: dout = 8'b10111011;
      13'h122: dout = 8'b10111011;
      13'h123: dout = 8'b10111011;
      13'h124: dout = 8'b10111011;
      13'h125: dout = 8'b10111011;
      13'h126: dout = 8'b10111011;
      13'h127: dout = 8'b10111011;
      13'h128: dout = 8'b10111011;
      13'h129: dout = 8'b10111011;
      13'h12A: dout = 8'b10111011;
      13'h12B: dout = 8'b10111011;
      13'h12C: dout = 8'b10111011;
      13'h12D: dout = 8'b10111011;
      13'h12E: dout = 8'b10111011;
      13'h12F: dout = 8'b10111011;
      13'h130: dout = 8'b10111011;
      13'h131: dout = 8'b10111011;
      13'h132: dout = 8'b10111011;
      13'h133: dout = 8'b10111011;
      13'h134: dout = 8'b10111011;
      13'h135: dout = 8'b10111011;
      13'h136: dout = 8'b10111011;
      13'h137: dout = 8'b10111011;
      13'h138: dout = 8'b10111011;
      13'h139: dout = 8'b10111011;
      13'h13A: dout = 8'b10111011;
      13'h13B: dout = 8'b10111011;
      13'h13C: dout = 8'b10111011;
      13'h13D: dout = 8'b10111011;
      13'h13E: dout = 8'b10111011;
      13'h13F: dout = 8'b10111011;
      13'h140: dout = 8'b10111011;
      13'h141: dout = 8'b10111011;
      13'h142: dout = 8'b10111011;
      13'h143: dout = 8'b10111011;
      13'h144: dout = 8'b10111011;
      13'h145: dout = 8'b10111011;
      13'h146: dout = 8'b10111011;
      13'h147: dout = 8'b10111011;
      13'h148: dout = 8'b10111011;
      13'h149: dout = 8'b10111011;
      13'h14A: dout = 8'b10111011;
      13'h14B: dout = 8'b10111011;
      13'h14C: dout = 8'b10111011;
      13'h14D: dout = 8'b10111011;
      13'h14E: dout = 8'b10111011;
      13'h14F: dout = 8'b10111011;
      13'h150: dout = 8'b10111011;
      13'h151: dout = 8'b10111011;
      13'h152: dout = 8'b10111011;
      13'h153: dout = 8'b10111011;
      13'h154: dout = 8'b10111011;
      13'h155: dout = 8'b10111011;
      13'h156: dout = 8'b10111011;
      13'h157: dout = 8'b10111011;
      13'h158: dout = 8'b10111011;
      13'h159: dout = 8'b10111011;
      13'h15A: dout = 8'b10111011;
      13'h15B: dout = 8'b10111011;
      13'h15C: dout = 8'b10111011;
      13'h15D: dout = 8'b10111011;
      13'h15E: dout = 8'b10111011;
      13'h15F: dout = 8'b10111011;
      13'h160: dout = 8'b10111011;
      13'h161: dout = 8'b10111011;
      13'h162: dout = 8'b10111011;
      13'h163: dout = 8'b10111011;
      13'h164: dout = 8'b10111011;
      13'h165: dout = 8'b10111011;
      13'h166: dout = 8'b10111011;
      13'h167: dout = 8'b10111011;
      13'h168: dout = 8'b10111011;
      13'h169: dout = 8'b10111011;
      13'h16A: dout = 8'b10111011;
      13'h16B: dout = 8'b10111011;
      13'h16C: dout = 8'b10111011;
      13'h16D: dout = 8'b10111011;
      13'h16E: dout = 8'b10111011;
      13'h16F: dout = 8'b10111011;
      13'h170: dout = 8'b10111011;
      13'h171: dout = 8'b10111011;
      13'h172: dout = 8'b10111011;
      13'h173: dout = 8'b10111011;
      13'h174: dout = 8'b10111011;
      13'h175: dout = 8'b10111011;
      13'h176: dout = 8'b10111011;
      13'h177: dout = 8'b10111011;
      13'h178: dout = 8'b10111011;
      13'h179: dout = 8'b10111011;
      13'h17A: dout = 8'b10111011;
      13'h17B: dout = 8'b10111011;
      13'h17C: dout = 8'b10111011;
      13'h17D: dout = 8'b10111011;
      13'h17E: dout = 8'b10111011;
      13'h17F: dout = 8'b10111011;
      13'h180: dout = 8'b10111011;
      13'h181: dout = 8'b10111011;
      13'h182: dout = 8'b10111011;
      13'h183: dout = 8'b10111011;
      13'h184: dout = 8'b10111011;
      13'h185: dout = 8'b10111011;
      13'h186: dout = 8'b10111011;
      13'h187: dout = 8'b10111011;
      13'h188: dout = 8'b10111011;
      13'h189: dout = 8'b10111011;
      13'h18A: dout = 8'b10111011;
      13'h18B: dout = 8'b10111011;
      13'h18C: dout = 8'b10111011;
      13'h18D: dout = 8'b10111011;
      13'h18E: dout = 8'b10111011;
      13'h18F: dout = 8'b10111011;
      13'h190: dout = 8'b10111011;
      13'h191: dout = 8'b10111011;
      13'h192: dout = 8'b10111011;
      13'h193: dout = 8'b10111011;
      13'h194: dout = 8'b10111011;
      13'h195: dout = 8'b10111011;
      13'h196: dout = 8'b10111011;
      13'h197: dout = 8'b10111011;
      13'h198: dout = 8'b10111011;
      13'h199: dout = 8'b10111011;
      13'h19A: dout = 8'b10111011;
      13'h19B: dout = 8'b10111011;
      13'h19C: dout = 8'b10111011;
      13'h19D: dout = 8'b10111011;
      13'h19E: dout = 8'b10111011;
      13'h19F: dout = 8'b10111011;
      13'h1A0: dout = 8'b10111011;
      13'h1A1: dout = 8'b10111011;
      13'h1A2: dout = 8'b10111011;
      13'h1A3: dout = 8'b10111011;
      13'h1A4: dout = 8'b10111011;
      13'h1A5: dout = 8'b10111011;
      13'h1A6: dout = 8'b10111011;
      13'h1A7: dout = 8'b10111011;
      13'h1A8: dout = 8'b10111011;
      13'h1A9: dout = 8'b10111011;
      13'h1AA: dout = 8'b10111011;
      13'h1AB: dout = 8'b10111011;
      13'h1AC: dout = 8'b10111011;
      13'h1AD: dout = 8'b10111011;
      13'h1AE: dout = 8'b10111011;
      13'h1AF: dout = 8'b10111011;
      13'h1B0: dout = 8'b10111011;
      13'h1B1: dout = 8'b10111011;
      13'h1B2: dout = 8'b10111011;
      13'h1B3: dout = 8'b10111011;
      13'h1B4: dout = 8'b10111011;
      13'h1B5: dout = 8'b10111011;
      13'h1B6: dout = 8'b10111011;
      13'h1B7: dout = 8'b10111011;
      13'h1B8: dout = 8'b10111011;
      13'h1B9: dout = 8'b10111011;
      13'h1BA: dout = 8'b10111011;
      13'h1BB: dout = 8'b10111011;
      13'h1BC: dout = 8'b10111011;
      13'h1BD: dout = 8'b10111011;
      13'h1BE: dout = 8'b10111011;
      13'h1BF: dout = 8'b10111011;
      13'h1C0: dout = 8'b10111011;
      13'h1C1: dout = 8'b10111011;
      13'h1C2: dout = 8'b10111011;
      13'h1C3: dout = 8'b10111011;
      13'h1C4: dout = 8'b10111011;
      13'h1C5: dout = 8'b10111011;
      13'h1C6: dout = 8'b10111011;
      13'h1C7: dout = 8'b10111011;
      13'h1C8: dout = 8'b10111011;
      13'h1C9: dout = 8'b10111011;
      13'h1CA: dout = 8'b10111011;
      13'h1CB: dout = 8'b10111011;
      13'h1CC: dout = 8'b10111011;
      13'h1CD: dout = 8'b10111011;
      13'h1CE: dout = 8'b10111011;
      13'h1CF: dout = 8'b10111011;
      13'h1D0: dout = 8'b10111011;
      13'h1D1: dout = 8'b10111011;
      13'h1D2: dout = 8'b10111011;
      13'h1D3: dout = 8'b10111011;
      13'h1D4: dout = 8'b10111011;
      13'h1D5: dout = 8'b10111011;
      13'h1D6: dout = 8'b10111011;
      13'h1D7: dout = 8'b10111011;
      13'h1D8: dout = 8'b10111011;
      13'h1D9: dout = 8'b10111011;
      13'h1DA: dout = 8'b10111011;
      13'h1DB: dout = 8'b10111011;
      13'h1DC: dout = 8'b10111011;
      13'h1DD: dout = 8'b10111011;
      13'h1DE: dout = 8'b10111011;
      13'h1DF: dout = 8'b10111011;
      13'h1E0: dout = 8'b10111011;
      13'h1E1: dout = 8'b10111011;
      13'h1E2: dout = 8'b10111011;
      13'h1E3: dout = 8'b10111011;
      13'h1E4: dout = 8'b10111011;
      13'h1E5: dout = 8'b10111011;
      13'h1E6: dout = 8'b10111011;
      13'h1E7: dout = 8'b10111011;
      13'h1E8: dout = 8'b10111011;
      13'h1E9: dout = 8'b10111011;
      13'h1EA: dout = 8'b10111011;
      13'h1EB: dout = 8'b10111011;
      13'h1EC: dout = 8'b10111011;
      13'h1ED: dout = 8'b10111011;
      13'h1EE: dout = 8'b10111011;
      13'h1EF: dout = 8'b10111011;
      13'h1F0: dout = 8'b10111011;
      13'h1F1: dout = 8'b10111011;
      13'h1F2: dout = 8'b10111011;
      13'h1F3: dout = 8'b10111011;
      13'h1F4: dout = 8'b10111011;
      13'h1F5: dout = 8'b10111011;
      13'h1F6: dout = 8'b10111011;
      13'h1F7: dout = 8'b10111011;
      13'h1F8: dout = 8'b10111011;
      13'h1F9: dout = 8'b10111011;
      13'h1FA: dout = 8'b10111011;
      13'h1FB: dout = 8'b10111011;
      13'h1FC: dout = 8'b10111011;
      13'h1FD: dout = 8'b10111011;
      13'h1FE: dout = 8'b10111011;
      13'h1FF: dout = 8'b10111011;
      13'h200: dout = 8'b10111011;
      13'h201: dout = 8'b10111011;
      13'h202: dout = 8'b10111011;
      13'h203: dout = 8'b10111011;
      13'h204: dout = 8'b10111011;
      13'h205: dout = 8'b10111011;
      13'h206: dout = 8'b10111011;
      13'h207: dout = 8'b10111011;
      13'h208: dout = 8'b10111011;
      13'h209: dout = 8'b10111011;
      13'h20A: dout = 8'b10111011;
      13'h20B: dout = 8'b10111011;
      13'h20C: dout = 8'b10111011;
      13'h20D: dout = 8'b10111011;
      13'h20E: dout = 8'b10111011;
      13'h20F: dout = 8'b10111011;
      13'h210: dout = 8'b10111011;
      13'h211: dout = 8'b10111011;
      13'h212: dout = 8'b10111011;
      13'h213: dout = 8'b10111011;
      13'h214: dout = 8'b10111011;
      13'h215: dout = 8'b10111011;
      13'h216: dout = 8'b10111011;
      13'h217: dout = 8'b10111011;
      13'h218: dout = 8'b10111011;
      13'h219: dout = 8'b10111011;
      13'h21A: dout = 8'b10111011;
      13'h21B: dout = 8'b10111011;
      13'h21C: dout = 8'b10111011;
      13'h21D: dout = 8'b10111011;
      13'h21E: dout = 8'b10111011;
      13'h21F: dout = 8'b10111011;
      13'h220: dout = 8'b10111011;
      13'h221: dout = 8'b10111011;
      13'h222: dout = 8'b10111011;
      13'h223: dout = 8'b10111011;
      13'h224: dout = 8'b10111011;
      13'h225: dout = 8'b10111011;
      13'h226: dout = 8'b10111011;
      13'h227: dout = 8'b10111011;
      13'h228: dout = 8'b10111011;
      13'h229: dout = 8'b10111011;
      13'h22A: dout = 8'b10111011;
      13'h22B: dout = 8'b10111011;
      13'h22C: dout = 8'b10111011;
      13'h22D: dout = 8'b10111011;
      13'h22E: dout = 8'b10111011;
      13'h22F: dout = 8'b10111011;
      13'h230: dout = 8'b10111011;
      13'h231: dout = 8'b10111011;
      13'h232: dout = 8'b10111011;
      13'h233: dout = 8'b10111011;
      13'h234: dout = 8'b10111011;
      13'h235: dout = 8'b10111011;
      13'h236: dout = 8'b10111011;
      13'h237: dout = 8'b10111011;
      13'h238: dout = 8'b10111011;
      13'h239: dout = 8'b10111011;
      13'h23A: dout = 8'b10111011;
      13'h23B: dout = 8'b10111011;
      13'h23C: dout = 8'b10111011;
      13'h23D: dout = 8'b10111011;
      13'h23E: dout = 8'b10111011;
      13'h23F: dout = 8'b10111011;
      13'h240: dout = 8'b10111011;
      13'h241: dout = 8'b10111011;
      13'h242: dout = 8'b10111011;
      13'h243: dout = 8'b10111011;
      13'h244: dout = 8'b10111011;
      13'h245: dout = 8'b10111011;
      13'h246: dout = 8'b10111011;
      13'h247: dout = 8'b10111011;
      13'h248: dout = 8'b10111011;
      13'h249: dout = 8'b10111011;
      13'h24A: dout = 8'b10111011;
      13'h24B: dout = 8'b10111011;
      13'h24C: dout = 8'b10111011;
      13'h24D: dout = 8'b10111011;
      13'h24E: dout = 8'b10111011;
      13'h24F: dout = 8'b10111011;
      13'h250: dout = 8'b10111011;
      13'h251: dout = 8'b10111011;
      13'h252: dout = 8'b10111011;
      13'h253: dout = 8'b10111011;
      13'h254: dout = 8'b10111011;
      13'h255: dout = 8'b10111011;
      13'h256: dout = 8'b10111011;
      13'h257: dout = 8'b10111011;
      13'h258: dout = 8'b10111011;
      13'h259: dout = 8'b10111011;
      13'h25A: dout = 8'b10111011;
      13'h25B: dout = 8'b10111011;
      13'h25C: dout = 8'b10111011;
      13'h25D: dout = 8'b10111011;
      13'h25E: dout = 8'b10111011;
      13'h25F: dout = 8'b10111011;
      13'h260: dout = 8'b10111011;
      13'h261: dout = 8'b10111011;
      13'h262: dout = 8'b10111011;
      13'h263: dout = 8'b10111011;
      13'h264: dout = 8'b10111011;
      13'h265: dout = 8'b10111011;
      13'h266: dout = 8'b10111011;
      13'h267: dout = 8'b10111011;
      13'h268: dout = 8'b10111011;
      13'h269: dout = 8'b10111011;
      13'h26A: dout = 8'b10111011;
      13'h26B: dout = 8'b10111011;
      13'h26C: dout = 8'b10111011;
      13'h26D: dout = 8'b10111011;
      13'h26E: dout = 8'b10111011;
      13'h26F: dout = 8'b10111011;
      13'h270: dout = 8'b10111011;
      13'h271: dout = 8'b10111011;
      13'h272: dout = 8'b10111011;
      13'h273: dout = 8'b10111011;
      13'h274: dout = 8'b10111011;
      13'h275: dout = 8'b10111011;
      13'h276: dout = 8'b10111011;
      13'h277: dout = 8'b10111011;
      13'h278: dout = 8'b10111011;
      13'h279: dout = 8'b10111011;
      13'h27A: dout = 8'b10111011;
      13'h27B: dout = 8'b10111011;
      13'h27C: dout = 8'b10111011;
      13'h27D: dout = 8'b10111011;
      13'h27E: dout = 8'b10111011;
      13'h27F: dout = 8'b10111011;
      13'h280: dout = 8'b10111011;
      13'h281: dout = 8'b10111011;
      13'h282: dout = 8'b10111011;
      13'h283: dout = 8'b10111011;
      13'h284: dout = 8'b10111011;
      13'h285: dout = 8'b10111011;
      13'h286: dout = 8'b10111011;
      13'h287: dout = 8'b10111011;
      13'h288: dout = 8'b10111011;
      13'h289: dout = 8'b10111011;
      13'h28A: dout = 8'b10111011;
      13'h28B: dout = 8'b10111011;
      13'h28C: dout = 8'b10111011;
      13'h28D: dout = 8'b10111011;
      13'h28E: dout = 8'b10111011;
      13'h28F: dout = 8'b10111011;
      13'h290: dout = 8'b10111011;
      13'h291: dout = 8'b10111011;
      13'h292: dout = 8'b10111011;
      13'h293: dout = 8'b10111011;
      13'h294: dout = 8'b10111011;
      13'h295: dout = 8'b10111011;
      13'h296: dout = 8'b10111011;
      13'h297: dout = 8'b10111011;
      13'h298: dout = 8'b10111011;
      13'h299: dout = 8'b10111011;
      13'h29A: dout = 8'b10111011;
      13'h29B: dout = 8'b10111011;
      13'h29C: dout = 8'b10111011;
      13'h29D: dout = 8'b10111011;
      13'h29E: dout = 8'b10111011;
      13'h29F: dout = 8'b10111011;
      13'h2A0: dout = 8'b10111011;
      13'h2A1: dout = 8'b10111011;
      13'h2A2: dout = 8'b10111011;
      13'h2A3: dout = 8'b10111011;
      13'h2A4: dout = 8'b10111011;
      13'h2A5: dout = 8'b10111011;
      13'h2A6: dout = 8'b10111011;
      13'h2A7: dout = 8'b10111011;
      13'h2A8: dout = 8'b10111011;
      13'h2A9: dout = 8'b10111011;
      13'h2AA: dout = 8'b10111011;
      13'h2AB: dout = 8'b10111011;
      13'h2AC: dout = 8'b10111011;
      13'h2AD: dout = 8'b10111011;
      13'h2AE: dout = 8'b10111011;
      13'h2AF: dout = 8'b10111011;
      13'h2B0: dout = 8'b10111011;
      13'h2B1: dout = 8'b10111011;
      13'h2B2: dout = 8'b10111011;
      13'h2B3: dout = 8'b10111011;
      13'h2B4: dout = 8'b10111011;
      13'h2B5: dout = 8'b10111011;
      13'h2B6: dout = 8'b10111011;
      13'h2B7: dout = 8'b10111011;
      13'h2B8: dout = 8'b10111011;
      13'h2B9: dout = 8'b10111011;
      13'h2BA: dout = 8'b10111011;
      13'h2BB: dout = 8'b10111011;
      13'h2BC: dout = 8'b10111011;
      13'h2BD: dout = 8'b10111011;
      13'h2BE: dout = 8'b10111011;
      13'h2BF: dout = 8'b10111011;
      13'h2C0: dout = 8'b10111011;
      13'h2C1: dout = 8'b10111011;
      13'h2C2: dout = 8'b10111011;
      13'h2C3: dout = 8'b10111011;
      13'h2C4: dout = 8'b10111011;
      13'h2C5: dout = 8'b10111011;
      13'h2C6: dout = 8'b10111011;
      13'h2C7: dout = 8'b10111011;
      13'h2C8: dout = 8'b10111011;
      13'h2C9: dout = 8'b10111011;
      13'h2CA: dout = 8'b10111011;
      13'h2CB: dout = 8'b10111011;
      13'h2CC: dout = 8'b10111011;
      13'h2CD: dout = 8'b10111011;
      13'h2CE: dout = 8'b10111011;
      13'h2CF: dout = 8'b10111011;
      13'h2D0: dout = 8'b10111011;
      13'h2D1: dout = 8'b10111011;
      13'h2D2: dout = 8'b10111011;
      13'h2D3: dout = 8'b10111011;
      13'h2D4: dout = 8'b10111011;
      13'h2D5: dout = 8'b10111011;
      13'h2D6: dout = 8'b10111011;
      13'h2D7: dout = 8'b10111011;
      13'h2D8: dout = 8'b10111011;
      13'h2D9: dout = 8'b10111011;
      13'h2DA: dout = 8'b10111011;
      13'h2DB: dout = 8'b10111011;
      13'h2DC: dout = 8'b10111011;
      13'h2DD: dout = 8'b10111011;
      13'h2DE: dout = 8'b10111011;
      13'h2DF: dout = 8'b10111011;
      13'h2E0: dout = 8'b10111011;
      13'h2E1: dout = 8'b10111011;
      13'h2E2: dout = 8'b10111011;
      13'h2E3: dout = 8'b10111011;
      13'h2E4: dout = 8'b10111011;
      13'h2E5: dout = 8'b10111011;
      13'h2E6: dout = 8'b10111011;
      13'h2E7: dout = 8'b10111011;
      13'h2E8: dout = 8'b10111011;
      13'h2E9: dout = 8'b10111011;
      13'h2EA: dout = 8'b10111011;
      13'h2EB: dout = 8'b10111011;
      13'h2EC: dout = 8'b10111011;
      13'h2ED: dout = 8'b10111011;
      13'h2EE: dout = 8'b10111011;
      13'h2EF: dout = 8'b10111011;
      13'h2F0: dout = 8'b10111011;
      13'h2F1: dout = 8'b10111011;
      13'h2F2: dout = 8'b10111011;
      13'h2F3: dout = 8'b10111011;
      13'h2F4: dout = 8'b10111011;
      13'h2F5: dout = 8'b10111011;
      13'h2F6: dout = 8'b10111011;
      13'h2F7: dout = 8'b10111011;
      13'h2F8: dout = 8'b10111011;
      13'h2F9: dout = 8'b10111011;
      13'h2FA: dout = 8'b10111011;
      13'h2FB: dout = 8'b10111011;
      13'h2FC: dout = 8'b10111011;
      13'h2FD: dout = 8'b10111011;
      13'h2FE: dout = 8'b10111011;
      13'h2FF: dout = 8'b10111011;
      13'h300: dout = 8'b10111011;
      13'h301: dout = 8'b10111011;
      13'h302: dout = 8'b10111011;
      13'h303: dout = 8'b10111011;
      13'h304: dout = 8'b10111011;
      13'h305: dout = 8'b10111011;
      13'h306: dout = 8'b10111011;
      13'h307: dout = 8'b10111011;
      13'h308: dout = 8'b10111011;
      13'h309: dout = 8'b10111011;
      13'h30A: dout = 8'b10111011;
      13'h30B: dout = 8'b10111011;
      13'h30C: dout = 8'b10111011;
      13'h30D: dout = 8'b10111011;
      13'h30E: dout = 8'b10111011;
      13'h30F: dout = 8'b10111011;
      13'h310: dout = 8'b10111011;
      13'h311: dout = 8'b10111011;
      13'h312: dout = 8'b10111011;
      13'h313: dout = 8'b10111011;
      13'h314: dout = 8'b10111011;
      13'h315: dout = 8'b10111011;
      13'h316: dout = 8'b10111011;
      13'h317: dout = 8'b10111011;
      13'h318: dout = 8'b10111011;
      13'h319: dout = 8'b10111011;
      13'h31A: dout = 8'b10111011;
      13'h31B: dout = 8'b10111011;
      13'h31C: dout = 8'b10111011;
      13'h31D: dout = 8'b10111011;
      13'h31E: dout = 8'b10111011;
      13'h31F: dout = 8'b10111011;
      13'h320: dout = 8'b10111011;
      13'h321: dout = 8'b10111011;
      13'h322: dout = 8'b10111011;
      13'h323: dout = 8'b10111011;
      13'h324: dout = 8'b10111011;
      13'h325: dout = 8'b10111011;
      13'h326: dout = 8'b10111011;
      13'h327: dout = 8'b10111011;
      13'h328: dout = 8'b10111011;
      13'h329: dout = 8'b10111011;
      13'h32A: dout = 8'b10111011;
      13'h32B: dout = 8'b10111011;
      13'h32C: dout = 8'b10111011;
      13'h32D: dout = 8'b10111011;
      13'h32E: dout = 8'b10111011;
      13'h32F: dout = 8'b10111011;
      13'h330: dout = 8'b10111011;
      13'h331: dout = 8'b10111011;
      13'h332: dout = 8'b10111011;
      13'h333: dout = 8'b10111011;
      13'h334: dout = 8'b10111011;
      13'h335: dout = 8'b10111011;
      13'h336: dout = 8'b10111011;
      13'h337: dout = 8'b10111011;
      13'h338: dout = 8'b10111011;
      13'h339: dout = 8'b10111011;
      13'h33A: dout = 8'b10111011;
      13'h33B: dout = 8'b10111011;
      13'h33C: dout = 8'b10111011;
      13'h33D: dout = 8'b10111011;
      13'h33E: dout = 8'b10111011;
      13'h33F: dout = 8'b10111011;
      13'h340: dout = 8'b10111011;
      13'h341: dout = 8'b10111011;
      13'h342: dout = 8'b10111011;
      13'h343: dout = 8'b10111011;
      13'h344: dout = 8'b10111011;
      13'h345: dout = 8'b10111011;
      13'h346: dout = 8'b10111011;
      13'h347: dout = 8'b10111011;
      13'h348: dout = 8'b10111011;
      13'h349: dout = 8'b10111011;
      13'h34A: dout = 8'b10111011;
      13'h34B: dout = 8'b10111011;
      13'h34C: dout = 8'b10111011;
      13'h34D: dout = 8'b10111011;
      13'h34E: dout = 8'b10111011;
      13'h34F: dout = 8'b10111011;
      13'h350: dout = 8'b10111011;
      13'h351: dout = 8'b10111011;
      13'h352: dout = 8'b10111011;
      13'h353: dout = 8'b10111011;
      13'h354: dout = 8'b10111011;
      13'h355: dout = 8'b10111011;
      13'h356: dout = 8'b10111011;
      13'h357: dout = 8'b10111011;
      13'h358: dout = 8'b10111011;
      13'h359: dout = 8'b10111011;
      13'h35A: dout = 8'b10111011;
      13'h35B: dout = 8'b10111011;
      13'h35C: dout = 8'b10111011;
      13'h35D: dout = 8'b10111011;
      13'h35E: dout = 8'b10111011;
      13'h35F: dout = 8'b10111011;
      13'h360: dout = 8'b10111011;
      13'h361: dout = 8'b10111011;
      13'h362: dout = 8'b10111011;
      13'h363: dout = 8'b10111011;
      13'h364: dout = 8'b10111011;
      13'h365: dout = 8'b10111011;
      13'h366: dout = 8'b10111011;
      13'h367: dout = 8'b10111011;
      13'h368: dout = 8'b10111011;
      13'h369: dout = 8'b10111011;
      13'h36A: dout = 8'b10111011;
      13'h36B: dout = 8'b10111011;
      13'h36C: dout = 8'b10111011;
      13'h36D: dout = 8'b10111011;
      13'h36E: dout = 8'b10111011;
      13'h36F: dout = 8'b10111011;
      13'h370: dout = 8'b10111011;
      13'h371: dout = 8'b10111011;
      13'h372: dout = 8'b10111011;
      13'h373: dout = 8'b10111011;
      13'h374: dout = 8'b10111011;
      13'h375: dout = 8'b10111011;
      13'h376: dout = 8'b10111011;
      13'h377: dout = 8'b10111011;
      13'h378: dout = 8'b10111011;
      13'h379: dout = 8'b10111011;
      13'h37A: dout = 8'b10111011;
      13'h37B: dout = 8'b10111011;
      13'h37C: dout = 8'b10111011;
      13'h37D: dout = 8'b10111011;
      13'h37E: dout = 8'b10111011;
      13'h37F: dout = 8'b10111011;
      13'h380: dout = 8'b10111011;
      13'h381: dout = 8'b10111011;
      13'h382: dout = 8'b10111011;
      13'h383: dout = 8'b10111011;
      13'h384: dout = 8'b10111011;
      13'h385: dout = 8'b10111011;
      13'h386: dout = 8'b10111011;
      13'h387: dout = 8'b10111011;
      13'h388: dout = 8'b10111011;
      13'h389: dout = 8'b10111011;
      13'h38A: dout = 8'b10111011;
      13'h38B: dout = 8'b10111011;
      13'h38C: dout = 8'b10111011;
      13'h38D: dout = 8'b10111011;
      13'h38E: dout = 8'b10111011;
      13'h38F: dout = 8'b10111011;
      13'h390: dout = 8'b10111011;
      13'h391: dout = 8'b10111011;
      13'h392: dout = 8'b10111011;
      13'h393: dout = 8'b10111011;
      13'h394: dout = 8'b10111011;
      13'h395: dout = 8'b10111011;
      13'h396: dout = 8'b10111011;
      13'h397: dout = 8'b10111011;
      13'h398: dout = 8'b10111011;
      13'h399: dout = 8'b10111011;
      13'h39A: dout = 8'b10111011;
      13'h39B: dout = 8'b10111011;
      13'h39C: dout = 8'b10111011;
      13'h39D: dout = 8'b10111011;
      13'h39E: dout = 8'b10111011;
      13'h39F: dout = 8'b10111011;
      13'h3A0: dout = 8'b10111011;
      13'h3A1: dout = 8'b10111011;
      13'h3A2: dout = 8'b10111011;
      13'h3A3: dout = 8'b10111011;
      13'h3A4: dout = 8'b10111011;
      13'h3A5: dout = 8'b10111011;
      13'h3A6: dout = 8'b10111011;
      13'h3A7: dout = 8'b10111011;
      13'h3A8: dout = 8'b10111011;
      13'h3A9: dout = 8'b10111011;
      13'h3AA: dout = 8'b10111011;
      13'h3AB: dout = 8'b10111011;
      13'h3AC: dout = 8'b10111011;
      13'h3AD: dout = 8'b10111011;
      13'h3AE: dout = 8'b10111011;
      13'h3AF: dout = 8'b10111011;
      13'h3B0: dout = 8'b10111011;
      13'h3B1: dout = 8'b10111011;
      13'h3B2: dout = 8'b10111011;
      13'h3B3: dout = 8'b10111011;
      13'h3B4: dout = 8'b10111011;
      13'h3B5: dout = 8'b10111011;
      13'h3B6: dout = 8'b10111011;
      13'h3B7: dout = 8'b10111011;
      13'h3B8: dout = 8'b10111011;
      13'h3B9: dout = 8'b10111011;
      13'h3BA: dout = 8'b10111011;
      13'h3BB: dout = 8'b10111011;
      13'h3BC: dout = 8'b10111011;
      13'h3BD: dout = 8'b10111011;
      13'h3BE: dout = 8'b10111011;
      13'h3BF: dout = 8'b10111011;
      13'h3C0: dout = 8'b10111011;
      13'h3C1: dout = 8'b10111011;
      13'h3C2: dout = 8'b10111011;
      13'h3C3: dout = 8'b10111011;
      13'h3C4: dout = 8'b10111011;
      13'h3C5: dout = 8'b10111011;
      13'h3C6: dout = 8'b10111011;
      13'h3C7: dout = 8'b10111011;
      13'h3C8: dout = 8'b10111011;
      13'h3C9: dout = 8'b10111011;
      13'h3CA: dout = 8'b10111011;
      13'h3CB: dout = 8'b10111011;
      13'h3CC: dout = 8'b10111011;
      13'h3CD: dout = 8'b10111011;
      13'h3CE: dout = 8'b10111011;
      13'h3CF: dout = 8'b10111011;
      13'h3D0: dout = 8'b10111011;
      13'h3D1: dout = 8'b10111011;
      13'h3D2: dout = 8'b10111011;
      13'h3D3: dout = 8'b10111011;
      13'h3D4: dout = 8'b10111011;
      13'h3D5: dout = 8'b10111011;
      13'h3D6: dout = 8'b10111011;
      13'h3D7: dout = 8'b10111011;
      13'h3D8: dout = 8'b10111011;
      13'h3D9: dout = 8'b10111011;
      13'h3DA: dout = 8'b10111011;
      13'h3DB: dout = 8'b10111011;
      13'h3DC: dout = 8'b10111011;
      13'h3DD: dout = 8'b10111011;
      13'h3DE: dout = 8'b10111011;
      13'h3DF: dout = 8'b10111011;
      13'h3E0: dout = 8'b10111011;
      13'h3E1: dout = 8'b10111011;
      13'h3E2: dout = 8'b10111011;
      13'h3E3: dout = 8'b10111011;
      13'h3E4: dout = 8'b10111011;
      13'h3E5: dout = 8'b10111011;
      13'h3E6: dout = 8'b10111011;
      13'h3E7: dout = 8'b10111011;
      13'h3E8: dout = 8'b10111011;
      13'h3E9: dout = 8'b10111011;
      13'h3EA: dout = 8'b10111011;
      13'h3EB: dout = 8'b10111011;
      13'h3EC: dout = 8'b10111011;
      13'h3ED: dout = 8'b10111011;
      13'h3EE: dout = 8'b10111011;
      13'h3EF: dout = 8'b10111011;
      13'h3F0: dout = 8'b10111011;
      13'h3F1: dout = 8'b10111011;
      13'h3F2: dout = 8'b10111011;
      13'h3F3: dout = 8'b10111011;
      13'h3F4: dout = 8'b10111011;
      13'h3F5: dout = 8'b10111011;
      13'h3F6: dout = 8'b10111011;
      13'h3F7: dout = 8'b10111011;
      13'h3F8: dout = 8'b10111011;
      13'h3F9: dout = 8'b10111011;
      13'h3FA: dout = 8'b10111011;
      13'h3FB: dout = 8'b10111011;
      13'h3FC: dout = 8'b10111011;
      13'h3FD: dout = 8'b10111011;
      13'h3FE: dout = 8'b10111011;
      13'h3FF: dout = 8'b10111011;
      13'h400: dout = 8'b10111011;
      13'h401: dout = 8'b10111011;
      13'h402: dout = 8'b10111011;
      13'h403: dout = 8'b10111011;
      13'h404: dout = 8'b10111011;
      13'h405: dout = 8'b10111011;
      13'h406: dout = 8'b10111011;
      13'h407: dout = 8'b10111011;
      13'h408: dout = 8'b10111011;
      13'h409: dout = 8'b10111011;
      13'h40A: dout = 8'b10111011;
      13'h40B: dout = 8'b10111011;
      13'h40C: dout = 8'b10111011;
      13'h40D: dout = 8'b10111011;
      13'h40E: dout = 8'b10111011;
      13'h40F: dout = 8'b10111011;
      13'h410: dout = 8'b10111011;
      13'h411: dout = 8'b10111011;
      13'h412: dout = 8'b10111011;
      13'h413: dout = 8'b10111011;
      13'h414: dout = 8'b10111011;
      13'h415: dout = 8'b10111011;
      13'h416: dout = 8'b10111011;
      13'h417: dout = 8'b10111011;
      13'h418: dout = 8'b10111011;
      13'h419: dout = 8'b10111011;
      13'h41A: dout = 8'b10111011;
      13'h41B: dout = 8'b10111011;
      13'h41C: dout = 8'b10111011;
      13'h41D: dout = 8'b10111011;
      13'h41E: dout = 8'b10111011;
      13'h41F: dout = 8'b10111011;
      13'h420: dout = 8'b10111011;
      13'h421: dout = 8'b10111011;
      13'h422: dout = 8'b10111011;
      13'h423: dout = 8'b10111011;
      13'h424: dout = 8'b10111011;
      13'h425: dout = 8'b10111011;
      13'h426: dout = 8'b10111011;
      13'h427: dout = 8'b10111011;
      13'h428: dout = 8'b10111011;
      13'h429: dout = 8'b10111011;
      13'h42A: dout = 8'b10111011;
      13'h42B: dout = 8'b10111011;
      13'h42C: dout = 8'b10111011;
      13'h42D: dout = 8'b10111011;
      13'h42E: dout = 8'b10111011;
      13'h42F: dout = 8'b10111011;
      13'h430: dout = 8'b10111011;
      13'h431: dout = 8'b10111011;
      13'h432: dout = 8'b10111011;
      13'h433: dout = 8'b10111011;
      13'h434: dout = 8'b10111011;
      13'h435: dout = 8'b10111011;
      13'h436: dout = 8'b10111011;
      13'h437: dout = 8'b10111011;
      13'h438: dout = 8'b10111011;
      13'h439: dout = 8'b10111011;
      13'h43A: dout = 8'b10111011;
      13'h43B: dout = 8'b10111011;
      13'h43C: dout = 8'b10111011;
      13'h43D: dout = 8'b10111011;
      13'h43E: dout = 8'b10111011;
      13'h43F: dout = 8'b10111011;
      13'h440: dout = 8'b10111011;
      13'h441: dout = 8'b10111011;
      13'h442: dout = 8'b10111011;
      13'h443: dout = 8'b10111011;
      13'h444: dout = 8'b10111011;
      13'h445: dout = 8'b10111011;
      13'h446: dout = 8'b10111011;
      13'h447: dout = 8'b10111011;
      13'h448: dout = 8'b10111011;
      13'h449: dout = 8'b10111011;
      13'h44A: dout = 8'b10111011;
      13'h44B: dout = 8'b10111011;
      13'h44C: dout = 8'b10111011;
      13'h44D: dout = 8'b10111011;
      13'h44E: dout = 8'b10111011;
      13'h44F: dout = 8'b10111011;
      13'h450: dout = 8'b10111011;
      13'h451: dout = 8'b10111011;
      13'h452: dout = 8'b10111011;
      13'h453: dout = 8'b10111011;
      13'h454: dout = 8'b10111011;
      13'h455: dout = 8'b10111011;
      13'h456: dout = 8'b10111011;
      13'h457: dout = 8'b10111011;
      13'h458: dout = 8'b10111011;
      13'h459: dout = 8'b10111011;
      13'h45A: dout = 8'b10111011;
      13'h45B: dout = 8'b10111011;
      13'h45C: dout = 8'b10111011;
      13'h45D: dout = 8'b10111011;
      13'h45E: dout = 8'b10111011;
      13'h45F: dout = 8'b10111011;
      13'h460: dout = 8'b10111011;
      13'h461: dout = 8'b10111011;
      13'h462: dout = 8'b10111011;
      13'h463: dout = 8'b10111011;
      13'h464: dout = 8'b10111011;
      13'h465: dout = 8'b10111011;
      13'h466: dout = 8'b10111011;
      13'h467: dout = 8'b10111011;
      13'h468: dout = 8'b10111011;
      13'h469: dout = 8'b10111011;
      13'h46A: dout = 8'b10111011;
      13'h46B: dout = 8'b10111011;
      13'h46C: dout = 8'b10111011;
      13'h46D: dout = 8'b10111011;
      13'h46E: dout = 8'b10111011;
      13'h46F: dout = 8'b10111011;
      13'h470: dout = 8'b10111011;
      13'h471: dout = 8'b10111011;
      13'h472: dout = 8'b10111011;
      13'h473: dout = 8'b10111011;
      13'h474: dout = 8'b10111011;
      13'h475: dout = 8'b10111011;
      13'h476: dout = 8'b10111011;
      13'h477: dout = 8'b10111011;
      13'h478: dout = 8'b10111011;
      13'h479: dout = 8'b10111011;
      13'h47A: dout = 8'b10111011;
      13'h47B: dout = 8'b10111011;
      13'h47C: dout = 8'b10111011;
      13'h47D: dout = 8'b10111011;
      13'h47E: dout = 8'b10111011;
      13'h47F: dout = 8'b10111011;
      13'h480: dout = 8'b10111011;
      13'h481: dout = 8'b10111011;
      13'h482: dout = 8'b10111011;
      13'h483: dout = 8'b10111011;
      13'h484: dout = 8'b10111011;
      13'h485: dout = 8'b10111011;
      13'h486: dout = 8'b10111011;
      13'h487: dout = 8'b10111011;
      13'h488: dout = 8'b10111011;
      13'h489: dout = 8'b10111011;
      13'h48A: dout = 8'b10111011;
      13'h48B: dout = 8'b10111011;
      13'h48C: dout = 8'b10111011;
      13'h48D: dout = 8'b10111011;
      13'h48E: dout = 8'b10111011;
      13'h48F: dout = 8'b10111011;
      13'h490: dout = 8'b10111011;
      13'h491: dout = 8'b10111011;
      13'h492: dout = 8'b10111011;
      13'h493: dout = 8'b10111011;
      13'h494: dout = 8'b10111011;
      13'h495: dout = 8'b10111011;
      13'h496: dout = 8'b10111011;
      13'h497: dout = 8'b10111011;
      13'h498: dout = 8'b10111011;
      13'h499: dout = 8'b10111011;
      13'h49A: dout = 8'b10111011;
      13'h49B: dout = 8'b10111011;
      13'h49C: dout = 8'b10111011;
      13'h49D: dout = 8'b10111011;
      13'h49E: dout = 8'b10111011;
      13'h49F: dout = 8'b10111011;
      13'h4A0: dout = 8'b10111011;
      13'h4A1: dout = 8'b10111011;
      13'h4A2: dout = 8'b10111011;
      13'h4A3: dout = 8'b10111011;
      13'h4A4: dout = 8'b10111011;
      13'h4A5: dout = 8'b10111011;
      13'h4A6: dout = 8'b10111011;
      13'h4A7: dout = 8'b10111011;
      13'h4A8: dout = 8'b10111011;
      13'h4A9: dout = 8'b10111011;
      13'h4AA: dout = 8'b10111011;
      13'h4AB: dout = 8'b10111011;
      13'h4AC: dout = 8'b10111011;
      13'h4AD: dout = 8'b10111011;
      13'h4AE: dout = 8'b10111011;
      13'h4AF: dout = 8'b10111011;
      13'h4B0: dout = 8'b10111011;
      13'h4B1: dout = 8'b10111011;
      13'h4B2: dout = 8'b10111011;
      13'h4B3: dout = 8'b10111011;
      13'h4B4: dout = 8'b10111011;
      13'h4B5: dout = 8'b10111011;
      13'h4B6: dout = 8'b10111011;
      13'h4B7: dout = 8'b10111011;
      13'h4B8: dout = 8'b10111011;
      13'h4B9: dout = 8'b10111011;
      13'h4BA: dout = 8'b10111011;
      13'h4BB: dout = 8'b10111011;
      13'h4BC: dout = 8'b10111011;
      13'h4BD: dout = 8'b10111011;
      13'h4BE: dout = 8'b10111011;
      13'h4BF: dout = 8'b10111011;
      13'h4C0: dout = 8'b10111011;
      13'h4C1: dout = 8'b10111011;
      13'h4C2: dout = 8'b10111011;
      13'h4C3: dout = 8'b10111011;
      13'h4C4: dout = 8'b10111011;
      13'h4C5: dout = 8'b10111011;
      13'h4C6: dout = 8'b10111011;
      13'h4C7: dout = 8'b10111011;
      13'h4C8: dout = 8'b10111011;
      13'h4C9: dout = 8'b10111011;
      13'h4CA: dout = 8'b10111011;
      13'h4CB: dout = 8'b10111011;
      13'h4CC: dout = 8'b10111011;
      13'h4CD: dout = 8'b10111011;
      13'h4CE: dout = 8'b10111011;
      13'h4CF: dout = 8'b10111011;
      13'h4D0: dout = 8'b10111011;
      13'h4D1: dout = 8'b10111011;
      13'h4D2: dout = 8'b10111011;
      13'h4D3: dout = 8'b10111011;
      13'h4D4: dout = 8'b10111011;
      13'h4D5: dout = 8'b10111011;
      13'h4D6: dout = 8'b10111011;
      13'h4D7: dout = 8'b10111011;
      13'h4D8: dout = 8'b10111011;
      13'h4D9: dout = 8'b10111011;
      13'h4DA: dout = 8'b10111011;
      13'h4DB: dout = 8'b10111011;
      13'h4DC: dout = 8'b10111011;
      13'h4DD: dout = 8'b10111011;
      13'h4DE: dout = 8'b10111011;
      13'h4DF: dout = 8'b10111011;
      13'h4E0: dout = 8'b10111011;
      13'h4E1: dout = 8'b10111011;
      13'h4E2: dout = 8'b10111011;
      13'h4E3: dout = 8'b10111011;
      13'h4E4: dout = 8'b10111011;
      13'h4E5: dout = 8'b10111011;
      13'h4E6: dout = 8'b10111011;
      13'h4E7: dout = 8'b10111011;
      13'h4E8: dout = 8'b10111011;
      13'h4E9: dout = 8'b10111011;
      13'h4EA: dout = 8'b10111011;
      13'h4EB: dout = 8'b10111011;
      13'h4EC: dout = 8'b10111011;
      13'h4ED: dout = 8'b10111011;
      13'h4EE: dout = 8'b10111011;
      13'h4EF: dout = 8'b10111011;
      13'h4F0: dout = 8'b10111011;
      13'h4F1: dout = 8'b10111011;
      13'h4F2: dout = 8'b10111011;
      13'h4F3: dout = 8'b10111011;
      13'h4F4: dout = 8'b10111011;
      13'h4F5: dout = 8'b10111011;
      13'h4F6: dout = 8'b10111011;
      13'h4F7: dout = 8'b10111011;
      13'h4F8: dout = 8'b10111011;
      13'h4F9: dout = 8'b10111011;
      13'h4FA: dout = 8'b10111011;
      13'h4FB: dout = 8'b10111011;
      13'h4FC: dout = 8'b10111011;
      13'h4FD: dout = 8'b10111011;
      13'h4FE: dout = 8'b10111011;
      13'h4FF: dout = 8'b10111011;
      13'h500: dout = 8'b10111011;
      13'h501: dout = 8'b10111011;
      13'h502: dout = 8'b10111011;
      13'h503: dout = 8'b10111011;
      13'h504: dout = 8'b10111011;
      13'h505: dout = 8'b10111011;
      13'h506: dout = 8'b10111011;
      13'h507: dout = 8'b10111011;
      13'h508: dout = 8'b10111011;
      13'h509: dout = 8'b10111011;
      13'h50A: dout = 8'b10111011;
      13'h50B: dout = 8'b10111011;
      13'h50C: dout = 8'b10111011;
      13'h50D: dout = 8'b10111011;
      13'h50E: dout = 8'b10111011;
      13'h50F: dout = 8'b10111011;
      13'h510: dout = 8'b10111011;
      13'h511: dout = 8'b10111011;
      13'h512: dout = 8'b10111011;
      13'h513: dout = 8'b10111011;
      13'h514: dout = 8'b10111011;
      13'h515: dout = 8'b10111011;
      13'h516: dout = 8'b10111011;
      13'h517: dout = 8'b10111011;
      13'h518: dout = 8'b10111011;
      13'h519: dout = 8'b10111011;
      13'h51A: dout = 8'b10111011;
      13'h51B: dout = 8'b10111011;
      13'h51C: dout = 8'b10111011;
      13'h51D: dout = 8'b10111011;
      13'h51E: dout = 8'b10111011;
      13'h51F: dout = 8'b10111011;
      13'h520: dout = 8'b10111011;
      13'h521: dout = 8'b10111011;
      13'h522: dout = 8'b10111011;
      13'h523: dout = 8'b10111011;
      13'h524: dout = 8'b10111011;
      13'h525: dout = 8'b10111011;
      13'h526: dout = 8'b10111011;
      13'h527: dout = 8'b10111011;
      13'h528: dout = 8'b10111011;
      13'h529: dout = 8'b10111011;
      13'h52A: dout = 8'b10111011;
      13'h52B: dout = 8'b10111011;
      13'h52C: dout = 8'b10111011;
      13'h52D: dout = 8'b10111011;
      13'h52E: dout = 8'b10111011;
      13'h52F: dout = 8'b10111011;
      13'h530: dout = 8'b10111011;
      13'h531: dout = 8'b10111011;
      13'h532: dout = 8'b10111011;
      13'h533: dout = 8'b10111011;
      13'h534: dout = 8'b10111011;
      13'h535: dout = 8'b10111011;
      13'h536: dout = 8'b10111011;
      13'h537: dout = 8'b10111011;
      13'h538: dout = 8'b10111011;
      13'h539: dout = 8'b10111011;
      13'h53A: dout = 8'b10111011;
      13'h53B: dout = 8'b10111011;
      13'h53C: dout = 8'b10111011;
      13'h53D: dout = 8'b10111011;
      13'h53E: dout = 8'b10111011;
      13'h53F: dout = 8'b10111011;
      13'h540: dout = 8'b10111011;
      13'h541: dout = 8'b10111011;
      13'h542: dout = 8'b10111011;
      13'h543: dout = 8'b10111011;
      13'h544: dout = 8'b10111011;
      13'h545: dout = 8'b10111011;
      13'h546: dout = 8'b10111011;
      13'h547: dout = 8'b10111011;
      13'h548: dout = 8'b10111011;
      13'h549: dout = 8'b10111011;
      13'h54A: dout = 8'b10111011;
      13'h54B: dout = 8'b10111011;
      13'h54C: dout = 8'b10111011;
      13'h54D: dout = 8'b10111011;
      13'h54E: dout = 8'b10111011;
      13'h54F: dout = 8'b10111011;
      13'h550: dout = 8'b10111011;
      13'h551: dout = 8'b10111011;
      13'h552: dout = 8'b10111011;
      13'h553: dout = 8'b10111011;
      13'h554: dout = 8'b10111011;
      13'h555: dout = 8'b10111011;
      13'h556: dout = 8'b10111011;
      13'h557: dout = 8'b10111011;
      13'h558: dout = 8'b10111011;
      13'h559: dout = 8'b10111011;
      13'h55A: dout = 8'b10111011;
      13'h55B: dout = 8'b10111011;
      13'h55C: dout = 8'b10111011;
      13'h55D: dout = 8'b10111011;
      13'h55E: dout = 8'b10111011;
      13'h55F: dout = 8'b10111011;
      13'h560: dout = 8'b10111011;
      13'h561: dout = 8'b10111011;
      13'h562: dout = 8'b10111011;
      13'h563: dout = 8'b10111011;
      13'h564: dout = 8'b10111011;
      13'h565: dout = 8'b10111011;
      13'h566: dout = 8'b10111011;
      13'h567: dout = 8'b10111011;
      13'h568: dout = 8'b10111011;
      13'h569: dout = 8'b10111011;
      13'h56A: dout = 8'b10111011;
      13'h56B: dout = 8'b10111011;
      13'h56C: dout = 8'b10111011;
      13'h56D: dout = 8'b10111011;
      13'h56E: dout = 8'b10111011;
      13'h56F: dout = 8'b10111011;
      13'h570: dout = 8'b10111011;
      13'h571: dout = 8'b10111011;
      13'h572: dout = 8'b10111011;
      13'h573: dout = 8'b10111011;
      13'h574: dout = 8'b10111011;
      13'h575: dout = 8'b10111011;
      13'h576: dout = 8'b10111011;
      13'h577: dout = 8'b10111011;
      13'h578: dout = 8'b10111011;
      13'h579: dout = 8'b10111011;
      13'h57A: dout = 8'b10111011;
      13'h57B: dout = 8'b10111011;
      13'h57C: dout = 8'b10111011;
      13'h57D: dout = 8'b10111011;
      13'h57E: dout = 8'b10111011;
      13'h57F: dout = 8'b10111011;
      13'h580: dout = 8'b10111011;
      13'h581: dout = 8'b10111011;
      13'h582: dout = 8'b10111011;
      13'h583: dout = 8'b10111011;
      13'h584: dout = 8'b10111011;
      13'h585: dout = 8'b10111011;
      13'h586: dout = 8'b10111011;
      13'h587: dout = 8'b10111011;
      13'h588: dout = 8'b10111011;
      13'h589: dout = 8'b10111011;
      13'h58A: dout = 8'b10111011;
      13'h58B: dout = 8'b10111011;
      13'h58C: dout = 8'b10111011;
      13'h58D: dout = 8'b10111011;
      13'h58E: dout = 8'b10111011;
      13'h58F: dout = 8'b10111011;
      13'h590: dout = 8'b10111011;
      13'h591: dout = 8'b10111011;
      13'h592: dout = 8'b10111011;
      13'h593: dout = 8'b10111011;
      13'h594: dout = 8'b10111011;
      13'h595: dout = 8'b10111011;
      13'h596: dout = 8'b10111011;
      13'h597: dout = 8'b10111011;
      13'h598: dout = 8'b10111011;
      13'h599: dout = 8'b10111011;
      13'h59A: dout = 8'b10111011;
      13'h59B: dout = 8'b10111011;
      13'h59C: dout = 8'b10111011;
      13'h59D: dout = 8'b10111011;
      13'h59E: dout = 8'b10111011;
      13'h59F: dout = 8'b10111011;
      13'h5A0: dout = 8'b10111011;
      13'h5A1: dout = 8'b10111011;
      13'h5A2: dout = 8'b10111011;
      13'h5A3: dout = 8'b10111011;
      13'h5A4: dout = 8'b10111011;
      13'h5A5: dout = 8'b10111011;
      13'h5A6: dout = 8'b10111011;
      13'h5A7: dout = 8'b10111011;
      13'h5A8: dout = 8'b10111011;
      13'h5A9: dout = 8'b10111011;
      13'h5AA: dout = 8'b10111011;
      13'h5AB: dout = 8'b10111011;
      13'h5AC: dout = 8'b10111011;
      13'h5AD: dout = 8'b10111011;
      13'h5AE: dout = 8'b10111011;
      13'h5AF: dout = 8'b10111011;
      13'h5B0: dout = 8'b10111011;
      13'h5B1: dout = 8'b10111011;
      13'h5B2: dout = 8'b10111011;
      13'h5B3: dout = 8'b10111011;
      13'h5B4: dout = 8'b10111011;
      13'h5B5: dout = 8'b10111011;
      13'h5B6: dout = 8'b10111011;
      13'h5B7: dout = 8'b10111011;
      13'h5B8: dout = 8'b10111011;
      13'h5B9: dout = 8'b10111011;
      13'h5BA: dout = 8'b10111011;
      13'h5BB: dout = 8'b10111011;
      13'h5BC: dout = 8'b10111011;
      13'h5BD: dout = 8'b10111011;
      13'h5BE: dout = 8'b10111011;
      13'h5BF: dout = 8'b10111011;
      13'h5C0: dout = 8'b10111011;
      13'h5C1: dout = 8'b10111011;
      13'h5C2: dout = 8'b10111011;
      13'h5C3: dout = 8'b10111011;
      13'h5C4: dout = 8'b10111011;
      13'h5C5: dout = 8'b10111011;
      13'h5C6: dout = 8'b10111011;
      13'h5C7: dout = 8'b10111011;
      13'h5C8: dout = 8'b10111011;
      13'h5C9: dout = 8'b10111011;
      13'h5CA: dout = 8'b10111011;
      13'h5CB: dout = 8'b10111011;
      13'h5CC: dout = 8'b10111011;
      13'h5CD: dout = 8'b10111011;
      13'h5CE: dout = 8'b10111011;
      13'h5CF: dout = 8'b10111011;
      13'h5D0: dout = 8'b10111011;
      13'h5D1: dout = 8'b10111011;
      13'h5D2: dout = 8'b10111011;
      13'h5D3: dout = 8'b10111011;
      13'h5D4: dout = 8'b10111011;
      13'h5D5: dout = 8'b10111011;
      13'h5D6: dout = 8'b10111011;
      13'h5D7: dout = 8'b10111011;
      13'h5D8: dout = 8'b10111011;
      13'h5D9: dout = 8'b10111011;
      13'h5DA: dout = 8'b10111011;
      13'h5DB: dout = 8'b10111011;
      13'h5DC: dout = 8'b10111011;
      13'h5DD: dout = 8'b10111011;
      13'h5DE: dout = 8'b10111011;
      13'h5DF: dout = 8'b10111011;
      13'h5E0: dout = 8'b10111011;
      13'h5E1: dout = 8'b10111011;
      13'h5E2: dout = 8'b10111011;
      13'h5E3: dout = 8'b10111011;
      13'h5E4: dout = 8'b10111011;
      13'h5E5: dout = 8'b10111011;
      13'h5E6: dout = 8'b10111011;
      13'h5E7: dout = 8'b10111011;
      13'h5E8: dout = 8'b10111011;
      13'h5E9: dout = 8'b10111011;
      13'h5EA: dout = 8'b10111011;
      13'h5EB: dout = 8'b10111011;
      13'h5EC: dout = 8'b10111011;
      13'h5ED: dout = 8'b10111011;
      13'h5EE: dout = 8'b10111011;
      13'h5EF: dout = 8'b10111011;
      13'h5F0: dout = 8'b10111011;
      13'h5F1: dout = 8'b10111011;
      13'h5F2: dout = 8'b10111011;
      13'h5F3: dout = 8'b10111011;
      13'h5F4: dout = 8'b10111011;
      13'h5F5: dout = 8'b10111011;
      13'h5F6: dout = 8'b10111011;
      13'h5F7: dout = 8'b10111011;
      13'h5F8: dout = 8'b10111011;
      13'h5F9: dout = 8'b10111011;
      13'h5FA: dout = 8'b10111011;
      13'h5FB: dout = 8'b10111011;
      13'h5FC: dout = 8'b10111011;
      13'h5FD: dout = 8'b10111011;
      13'h5FE: dout = 8'b10111011;
      13'h5FF: dout = 8'b10111011;
      13'h600: dout = 8'b10111011;
      13'h601: dout = 8'b10111011;
      13'h602: dout = 8'b10111011;
      13'h603: dout = 8'b10111011;
      13'h604: dout = 8'b10111011;
      13'h605: dout = 8'b10111011;
      13'h606: dout = 8'b10111011;
      13'h607: dout = 8'b10111011;
      13'h608: dout = 8'b10111011;
      13'h609: dout = 8'b10111011;
      13'h60A: dout = 8'b10111011;
      13'h60B: dout = 8'b10111011;
      13'h60C: dout = 8'b10111011;
      13'h60D: dout = 8'b10111011;
      13'h60E: dout = 8'b10111011;
      13'h60F: dout = 8'b10111011;
      13'h610: dout = 8'b10111011;
      13'h611: dout = 8'b10111011;
      13'h612: dout = 8'b10111011;
      13'h613: dout = 8'b10111011;
      13'h614: dout = 8'b10111011;
      13'h615: dout = 8'b10111011;
      13'h616: dout = 8'b10111011;
      13'h617: dout = 8'b10111011;
      13'h618: dout = 8'b10111011;
      13'h619: dout = 8'b10111011;
      13'h61A: dout = 8'b10111011;
      13'h61B: dout = 8'b10111011;
      13'h61C: dout = 8'b10111011;
      13'h61D: dout = 8'b10111011;
      13'h61E: dout = 8'b10111011;
      13'h61F: dout = 8'b10111011;
      13'h620: dout = 8'b10111011;
      13'h621: dout = 8'b10111011;
      13'h622: dout = 8'b10111011;
      13'h623: dout = 8'b10111011;
      13'h624: dout = 8'b10111011;
      13'h625: dout = 8'b10111011;
      13'h626: dout = 8'b10111011;
      13'h627: dout = 8'b10111011;
      13'h628: dout = 8'b10111011;
      13'h629: dout = 8'b10111011;
      13'h62A: dout = 8'b10111011;
      13'h62B: dout = 8'b10111011;
      13'h62C: dout = 8'b10111011;
      13'h62D: dout = 8'b10111011;
      13'h62E: dout = 8'b10111011;
      13'h62F: dout = 8'b10111011;
      13'h630: dout = 8'b10111011;
      13'h631: dout = 8'b10111011;
      13'h632: dout = 8'b10111011;
      13'h633: dout = 8'b10111011;
      13'h634: dout = 8'b10111011;
      13'h635: dout = 8'b10111011;
      13'h636: dout = 8'b10111011;
      13'h637: dout = 8'b10111011;
      13'h638: dout = 8'b10111011;
      13'h639: dout = 8'b10111011;
      13'h63A: dout = 8'b10111011;
      13'h63B: dout = 8'b10111011;
      13'h63C: dout = 8'b10111011;
      13'h63D: dout = 8'b10111011;
      13'h63E: dout = 8'b10111011;
      13'h63F: dout = 8'b10111011;
      13'h640: dout = 8'b10111011;
      13'h641: dout = 8'b10111011;
      13'h642: dout = 8'b10111011;
      13'h643: dout = 8'b10111011;
      13'h644: dout = 8'b10111011;
      13'h645: dout = 8'b10111011;
      13'h646: dout = 8'b10111011;
      13'h647: dout = 8'b10111011;
      13'h648: dout = 8'b10111011;
      13'h649: dout = 8'b10111011;
      13'h64A: dout = 8'b10111011;
      13'h64B: dout = 8'b10111011;
      13'h64C: dout = 8'b10111011;
      13'h64D: dout = 8'b10111011;
      13'h64E: dout = 8'b10111011;
      13'h64F: dout = 8'b10111011;
      13'h650: dout = 8'b10111011;
      13'h651: dout = 8'b10111011;
      13'h652: dout = 8'b10111011;
      13'h653: dout = 8'b10111011;
      13'h654: dout = 8'b10111011;
      13'h655: dout = 8'b10111011;
      13'h656: dout = 8'b10111011;
      13'h657: dout = 8'b10111011;
      13'h658: dout = 8'b10111011;
      13'h659: dout = 8'b10111011;
      13'h65A: dout = 8'b10111011;
      13'h65B: dout = 8'b10111011;
      13'h65C: dout = 8'b10111011;
      13'h65D: dout = 8'b10111011;
      13'h65E: dout = 8'b10111011;
      13'h65F: dout = 8'b10111011;
      13'h660: dout = 8'b10111011;
      13'h661: dout = 8'b10111011;
      13'h662: dout = 8'b10111011;
      13'h663: dout = 8'b10111011;
      13'h664: dout = 8'b10111011;
      13'h665: dout = 8'b10111011;
      13'h666: dout = 8'b10111011;
      13'h667: dout = 8'b10111011;
      13'h668: dout = 8'b10111011;
      13'h669: dout = 8'b10111011;
      13'h66A: dout = 8'b10111011;
      13'h66B: dout = 8'b10111011;
      13'h66C: dout = 8'b10111011;
      13'h66D: dout = 8'b10111011;
      13'h66E: dout = 8'b10111011;
      13'h66F: dout = 8'b10111011;
      13'h670: dout = 8'b10111011;
      13'h671: dout = 8'b10111011;
      13'h672: dout = 8'b10111011;
      13'h673: dout = 8'b10111011;
      13'h674: dout = 8'b10111011;
      13'h675: dout = 8'b10111011;
      13'h676: dout = 8'b10111011;
      13'h677: dout = 8'b10111011;
      13'h678: dout = 8'b10111011;
      13'h679: dout = 8'b10111011;
      13'h67A: dout = 8'b10111011;
      13'h67B: dout = 8'b10111011;
      13'h67C: dout = 8'b10111011;
      13'h67D: dout = 8'b10111011;
      13'h67E: dout = 8'b10111011;
      13'h67F: dout = 8'b10111011;
      13'h680: dout = 8'b10111011;
      13'h681: dout = 8'b10111011;
      13'h682: dout = 8'b10111011;
      13'h683: dout = 8'b10111011;
      13'h684: dout = 8'b10111011;
      13'h685: dout = 8'b10111011;
      13'h686: dout = 8'b10111011;
      13'h687: dout = 8'b10111011;
      13'h688: dout = 8'b10111011;
      13'h689: dout = 8'b10111011;
      13'h68A: dout = 8'b10111011;
      13'h68B: dout = 8'b10111011;
      13'h68C: dout = 8'b10111011;
      13'h68D: dout = 8'b10111011;
      13'h68E: dout = 8'b10111011;
      13'h68F: dout = 8'b10111011;
      13'h690: dout = 8'b10111011;
      13'h691: dout = 8'b10111011;
      13'h692: dout = 8'b10111011;
      13'h693: dout = 8'b10111011;
      13'h694: dout = 8'b10111011;
      13'h695: dout = 8'b10111011;
      13'h696: dout = 8'b10111011;
      13'h697: dout = 8'b10111011;
      13'h698: dout = 8'b10111011;
      13'h699: dout = 8'b10111011;
      13'h69A: dout = 8'b10111011;
      13'h69B: dout = 8'b10111011;
      13'h69C: dout = 8'b10111011;
      13'h69D: dout = 8'b10111011;
      13'h69E: dout = 8'b10111011;
      13'h69F: dout = 8'b10111011;
      13'h6A0: dout = 8'b10111011;
      13'h6A1: dout = 8'b10111011;
      13'h6A2: dout = 8'b10111011;
      13'h6A3: dout = 8'b10111011;
      13'h6A4: dout = 8'b10111011;
      13'h6A5: dout = 8'b10111011;
      13'h6A6: dout = 8'b10111011;
      13'h6A7: dout = 8'b10111011;
      13'h6A8: dout = 8'b10111011;
      13'h6A9: dout = 8'b10111011;
      13'h6AA: dout = 8'b10111011;
      13'h6AB: dout = 8'b10111011;
      13'h6AC: dout = 8'b10111011;
      13'h6AD: dout = 8'b10111011;
      13'h6AE: dout = 8'b10111011;
      13'h6AF: dout = 8'b10111011;
      13'h6B0: dout = 8'b10111011;
      13'h6B1: dout = 8'b10111011;
      13'h6B2: dout = 8'b10111011;
      13'h6B3: dout = 8'b10111011;
      13'h6B4: dout = 8'b10111011;
      13'h6B5: dout = 8'b10111011;
      13'h6B6: dout = 8'b10111011;
      13'h6B7: dout = 8'b10111011;
      13'h6B8: dout = 8'b10111011;
      13'h6B9: dout = 8'b10111011;
      13'h6BA: dout = 8'b10111011;
      13'h6BB: dout = 8'b10111011;
      13'h6BC: dout = 8'b10111011;
      13'h6BD: dout = 8'b10111011;
      13'h6BE: dout = 8'b10111011;
      13'h6BF: dout = 8'b10111011;
      13'h6C0: dout = 8'b10111011;
      13'h6C1: dout = 8'b10111011;
      13'h6C2: dout = 8'b10111011;
      13'h6C3: dout = 8'b10111011;
      13'h6C4: dout = 8'b10111011;
      13'h6C5: dout = 8'b10111011;
      13'h6C6: dout = 8'b10111011;
      13'h6C7: dout = 8'b10111011;
      13'h6C8: dout = 8'b10111011;
      13'h6C9: dout = 8'b10111011;
      13'h6CA: dout = 8'b10111011;
      13'h6CB: dout = 8'b10111011;
      13'h6CC: dout = 8'b10111011;
      13'h6CD: dout = 8'b10111011;
      13'h6CE: dout = 8'b10111011;
      13'h6CF: dout = 8'b10111011;
      13'h6D0: dout = 8'b10111011;
      13'h6D1: dout = 8'b10111011;
      13'h6D2: dout = 8'b10111011;
      13'h6D3: dout = 8'b10111011;
      13'h6D4: dout = 8'b10111011;
      13'h6D5: dout = 8'b10111011;
      13'h6D6: dout = 8'b10111011;
      13'h6D7: dout = 8'b10111011;
      13'h6D8: dout = 8'b10111011;
      13'h6D9: dout = 8'b10111011;
      13'h6DA: dout = 8'b10111011;
      13'h6DB: dout = 8'b10111011;
      13'h6DC: dout = 8'b10111011;
      13'h6DD: dout = 8'b10111011;
      13'h6DE: dout = 8'b10111011;
      13'h6DF: dout = 8'b10111011;
      13'h6E0: dout = 8'b10111011;
      13'h6E1: dout = 8'b10111011;
      13'h6E2: dout = 8'b10111011;
      13'h6E3: dout = 8'b10111011;
      13'h6E4: dout = 8'b10111011;
      13'h6E5: dout = 8'b10111011;
      13'h6E6: dout = 8'b10111011;
      13'h6E7: dout = 8'b10111011;
      13'h6E8: dout = 8'b10111011;
      13'h6E9: dout = 8'b10111011;
      13'h6EA: dout = 8'b10111011;
      13'h6EB: dout = 8'b10111011;
      13'h6EC: dout = 8'b10111011;
      13'h6ED: dout = 8'b10111011;
      13'h6EE: dout = 8'b10111011;
      13'h6EF: dout = 8'b10111011;
      13'h6F0: dout = 8'b10111011;
      13'h6F1: dout = 8'b10111011;
      13'h6F2: dout = 8'b10111011;
      13'h6F3: dout = 8'b10111011;
      13'h6F4: dout = 8'b10111011;
      13'h6F5: dout = 8'b11100000;
      13'h6F6: dout = 8'b11100000;
      13'h6F7: dout = 8'b11100000;
      13'h6F8: dout = 8'b11100000;
      13'h6F9: dout = 8'b11100000;
      13'h6FA: dout = 8'b11100000;
      13'h6FB: dout = 8'b11100000;
      13'h6FC: dout = 8'b11100000;
      13'h6FD: dout = 8'b11100000;
      13'h6FE: dout = 8'b11100000;
      13'h6FF: dout = 8'b11100000;
      13'h700: dout = 8'b11100000;
      13'h701: dout = 8'b11100000;
      13'h702: dout = 8'b11100000;
      13'h703: dout = 8'b11100000;
      13'h704: dout = 8'b11100000;
      13'h705: dout = 8'b11100000;
      13'h706: dout = 8'b11100000;
      13'h707: dout = 8'b11100000;
      13'h708: dout = 8'b11100000;
      13'h709: dout = 8'b11100000;
      13'h70A: dout = 8'b11100000;
      13'h70B: dout = 8'b10111011;
      13'h70C: dout = 8'b10111011;
      13'h70D: dout = 8'b10111011;
      13'h70E: dout = 8'b10111011;
      13'h70F: dout = 8'b10111011;
      13'h710: dout = 8'b10111011;
      13'h711: dout = 8'b10111011;
      13'h712: dout = 8'b10111011;
      13'h713: dout = 8'b10111011;
      13'h714: dout = 8'b10111011;
      13'h715: dout = 8'b10111011;
      13'h716: dout = 8'b10111011;
      13'h717: dout = 8'b10111011;
      13'h718: dout = 8'b10111011;
      13'h719: dout = 8'b10111011;
      13'h71A: dout = 8'b10111011;
      13'h71B: dout = 8'b10111011;
      13'h71C: dout = 8'b10111011;
      13'h71D: dout = 8'b10111011;
      13'h71E: dout = 8'b10111011;
      13'h71F: dout = 8'b10111011;
      13'h720: dout = 8'b10111011;
      13'h721: dout = 8'b10111011;
      13'h722: dout = 8'b10111011;
      13'h723: dout = 8'b10111011;
      13'h724: dout = 8'b10111011;
      13'h725: dout = 8'b10111011;
      13'h726: dout = 8'b10111011;
      13'h727: dout = 8'b10111011;
      13'h728: dout = 8'b10111011;
      13'h729: dout = 8'b10111011;
      13'h72A: dout = 8'b10111011;
      13'h72B: dout = 8'b10111011;
      13'h72C: dout = 8'b10111011;
      13'h72D: dout = 8'b10111011;
      13'h72E: dout = 8'b10111011;
      13'h72F: dout = 8'b10111011;
      13'h730: dout = 8'b10111011;
      13'h731: dout = 8'b10111011;
      13'h732: dout = 8'b10111011;
      13'h733: dout = 8'b10111011;
      13'h734: dout = 8'b10111011;
      13'h735: dout = 8'b10111011;
      13'h736: dout = 8'b10111011;
      13'h737: dout = 8'b10111011;
      13'h738: dout = 8'b10111011;
      13'h739: dout = 8'b10111011;
      13'h73A: dout = 8'b10111011;
      13'h73B: dout = 8'b10111011;
      13'h73C: dout = 8'b10111011;
      13'h73D: dout = 8'b10111011;
      13'h73E: dout = 8'b10111011;
      13'h73F: dout = 8'b10111011;
      13'h740: dout = 8'b10111011;
      13'h741: dout = 8'b10111011;
      13'h742: dout = 8'b10111011;
      13'h743: dout = 8'b10111011;
      13'h744: dout = 8'b10111011;
      13'h745: dout = 8'b11100000;
      13'h746: dout = 8'b11100000;
      13'h747: dout = 8'b11100000;
      13'h748: dout = 8'b11100000;
      13'h749: dout = 8'b11100000;
      13'h74A: dout = 8'b11100000;
      13'h74B: dout = 8'b11100000;
      13'h74C: dout = 8'b11100000;
      13'h74D: dout = 8'b11100000;
      13'h74E: dout = 8'b11100000;
      13'h74F: dout = 8'b11100000;
      13'h750: dout = 8'b11100000;
      13'h751: dout = 8'b11100000;
      13'h752: dout = 8'b11100000;
      13'h753: dout = 8'b11100000;
      13'h754: dout = 8'b11100000;
      13'h755: dout = 8'b11100000;
      13'h756: dout = 8'b11100000;
      13'h757: dout = 8'b11100000;
      13'h758: dout = 8'b11100000;
      13'h759: dout = 8'b11100000;
      13'h75A: dout = 8'b11100000;
      13'h75B: dout = 8'b10111011;
      13'h75C: dout = 8'b10111011;
      13'h75D: dout = 8'b10111011;
      13'h75E: dout = 8'b10111011;
      13'h75F: dout = 8'b10111011;
      13'h760: dout = 8'b10111011;
      13'h761: dout = 8'b10111011;
      13'h762: dout = 8'b10111011;
      13'h763: dout = 8'b10111011;
      13'h764: dout = 8'b10111011;
      13'h765: dout = 8'b10111011;
      13'h766: dout = 8'b10111011;
      13'h767: dout = 8'b10111011;
      13'h768: dout = 8'b10111011;
      13'h769: dout = 8'b10111011;
      13'h76A: dout = 8'b10111011;
      13'h76B: dout = 8'b10111011;
      13'h76C: dout = 8'b10111011;
      13'h76D: dout = 8'b10111011;
      13'h76E: dout = 8'b10111011;
      13'h76F: dout = 8'b10111011;
      13'h770: dout = 8'b10111011;
      13'h771: dout = 8'b10111011;
      13'h772: dout = 8'b10111011;
      13'h773: dout = 8'b10111011;
      13'h774: dout = 8'b10111011;
      13'h775: dout = 8'b10111011;
      13'h776: dout = 8'b10111011;
      13'h777: dout = 8'b10111011;
      13'h778: dout = 8'b10111011;
      13'h779: dout = 8'b10111011;
      13'h77A: dout = 8'b10111011;
      13'h77B: dout = 8'b10111011;
      13'h77C: dout = 8'b10111011;
      13'h77D: dout = 8'b10111011;
      13'h77E: dout = 8'b10111011;
      13'h77F: dout = 8'b10111011;
      13'h780: dout = 8'b10111011;
      13'h781: dout = 8'b10111011;
      13'h782: dout = 8'b10111011;
      13'h783: dout = 8'b10111011;
      13'h784: dout = 8'b10111011;
      13'h785: dout = 8'b10111011;
      13'h786: dout = 8'b10111011;
      13'h787: dout = 8'b10111011;
      13'h788: dout = 8'b10111011;
      13'h789: dout = 8'b10111011;
      13'h78A: dout = 8'b10111011;
      13'h78B: dout = 8'b10111011;
      13'h78C: dout = 8'b10111011;
      13'h78D: dout = 8'b10111011;
      13'h78E: dout = 8'b10111011;
      13'h78F: dout = 8'b10111011;
      13'h790: dout = 8'b10111011;
      13'h791: dout = 8'b10111011;
      13'h792: dout = 8'b10111011;
      13'h793: dout = 8'b10111011;
      13'h794: dout = 8'b10111011;
      13'h795: dout = 8'b11100000;
      13'h796: dout = 8'b11100000;
      13'h797: dout = 8'b11100000;
      13'h798: dout = 8'b11100000;
      13'h799: dout = 8'b11100000;
      13'h79A: dout = 8'b11100000;
      13'h79B: dout = 8'b11100000;
      13'h79C: dout = 8'b11100000;
      13'h79D: dout = 8'b11100000;
      13'h79E: dout = 8'b11100000;
      13'h79F: dout = 8'b11100000;
      13'h7A0: dout = 8'b11100000;
      13'h7A1: dout = 8'b11100000;
      13'h7A2: dout = 8'b11100000;
      13'h7A3: dout = 8'b11100000;
      13'h7A4: dout = 8'b11100000;
      13'h7A5: dout = 8'b11100000;
      13'h7A6: dout = 8'b11100000;
      13'h7A7: dout = 8'b11100000;
      13'h7A8: dout = 8'b11100000;
      13'h7A9: dout = 8'b11100000;
      13'h7AA: dout = 8'b11100000;
      13'h7AB: dout = 8'b10111011;
      13'h7AC: dout = 8'b10111011;
      13'h7AD: dout = 8'b10111011;
      13'h7AE: dout = 8'b10111011;
      13'h7AF: dout = 8'b10111011;
      13'h7B0: dout = 8'b10111011;
      13'h7B1: dout = 8'b10111011;
      13'h7B2: dout = 8'b10111011;
      13'h7B3: dout = 8'b10111011;
      13'h7B4: dout = 8'b10111011;
      13'h7B5: dout = 8'b10111011;
      13'h7B6: dout = 8'b10111011;
      13'h7B7: dout = 8'b10111011;
      13'h7B8: dout = 8'b10111011;
      13'h7B9: dout = 8'b10111011;
      13'h7BA: dout = 8'b10111011;
      13'h7BB: dout = 8'b10111011;
      13'h7BC: dout = 8'b10111011;
      13'h7BD: dout = 8'b10111011;
      13'h7BE: dout = 8'b10111011;
      13'h7BF: dout = 8'b10111011;
      13'h7C0: dout = 8'b10111011;
      13'h7C1: dout = 8'b10111011;
      13'h7C2: dout = 8'b10111011;
      13'h7C3: dout = 8'b10111011;
      13'h7C4: dout = 8'b10111011;
      13'h7C5: dout = 8'b10111011;
      13'h7C6: dout = 8'b10111011;
      13'h7C7: dout = 8'b10111011;
      13'h7C8: dout = 8'b10111011;
      13'h7C9: dout = 8'b10111011;
      13'h7CA: dout = 8'b10111011;
      13'h7CB: dout = 8'b10111011;
      13'h7CC: dout = 8'b10111011;
      13'h7CD: dout = 8'b10111011;
      13'h7CE: dout = 8'b10111011;
      13'h7CF: dout = 8'b10111011;
      13'h7D0: dout = 8'b10111011;
      13'h7D1: dout = 8'b10111011;
      13'h7D2: dout = 8'b10111011;
      13'h7D3: dout = 8'b10111011;
      13'h7D4: dout = 8'b10111011;
      13'h7D5: dout = 8'b10111011;
      13'h7D6: dout = 8'b10111011;
      13'h7D7: dout = 8'b10111011;
      13'h7D8: dout = 8'b10111011;
      13'h7D9: dout = 8'b10111011;
      13'h7DA: dout = 8'b10111011;
      13'h7DB: dout = 8'b10111011;
      13'h7DC: dout = 8'b10111011;
      13'h7DD: dout = 8'b10111011;
      13'h7DE: dout = 8'b10111011;
      13'h7DF: dout = 8'b10111011;
      13'h7E0: dout = 8'b10111011;
      13'h7E1: dout = 8'b10111011;
      13'h7E2: dout = 8'b10111011;
      13'h7E3: dout = 8'b10111011;
      13'h7E4: dout = 8'b10111011;
      13'h7E5: dout = 8'b11100000;
      13'h7E6: dout = 8'b11100000;
      13'h7E7: dout = 8'b11100000;
      13'h7E8: dout = 8'b11100000;
      13'h7E9: dout = 8'b11100000;
      13'h7EA: dout = 8'b11100000;
      13'h7EB: dout = 8'b11100000;
      13'h7EC: dout = 8'b11100000;
      13'h7ED: dout = 8'b11100000;
      13'h7EE: dout = 8'b11100000;
      13'h7EF: dout = 8'b11100000;
      13'h7F0: dout = 8'b11100000;
      13'h7F1: dout = 8'b11100000;
      13'h7F2: dout = 8'b11100000;
      13'h7F3: dout = 8'b11100000;
      13'h7F4: dout = 8'b11100000;
      13'h7F5: dout = 8'b11100000;
      13'h7F6: dout = 8'b11100000;
      13'h7F7: dout = 8'b11100000;
      13'h7F8: dout = 8'b11100000;
      13'h7F9: dout = 8'b11100000;
      13'h7FA: dout = 8'b11100000;
      13'h7FB: dout = 8'b10111011;
      13'h7FC: dout = 8'b10111011;
      13'h7FD: dout = 8'b10111011;
      13'h7FE: dout = 8'b10111011;
      13'h7FF: dout = 8'b10111011;
      13'h800: dout = 8'b10111011;
      13'h801: dout = 8'b10111011;
      13'h802: dout = 8'b10111011;
      13'h803: dout = 8'b10111011;
      13'h804: dout = 8'b10111011;
      13'h805: dout = 8'b10111011;
      13'h806: dout = 8'b10111011;
      13'h807: dout = 8'b10111011;
      13'h808: dout = 8'b10111011;
      13'h809: dout = 8'b10111011;
      13'h80A: dout = 8'b10111011;
      13'h80B: dout = 8'b10111011;
      13'h80C: dout = 8'b10111011;
      13'h80D: dout = 8'b10111011;
      13'h80E: dout = 8'b10111011;
      13'h80F: dout = 8'b10111011;
      13'h810: dout = 8'b10111011;
      13'h811: dout = 8'b10111011;
      13'h812: dout = 8'b10111011;
      13'h813: dout = 8'b10111011;
      13'h814: dout = 8'b10111011;
      13'h815: dout = 8'b10111011;
      13'h816: dout = 8'b10111011;
      13'h817: dout = 8'b10111011;
      13'h818: dout = 8'b10111011;
      13'h819: dout = 8'b10111011;
      13'h81A: dout = 8'b10111011;
      13'h81B: dout = 8'b10111011;
      13'h81C: dout = 8'b10111011;
      13'h81D: dout = 8'b10111011;
      13'h81E: dout = 8'b10111011;
      13'h81F: dout = 8'b10111011;
      13'h820: dout = 8'b10111011;
      13'h821: dout = 8'b10111011;
      13'h822: dout = 8'b10111011;
      13'h823: dout = 8'b10111011;
      13'h824: dout = 8'b10111011;
      13'h825: dout = 8'b10111011;
      13'h826: dout = 8'b10111011;
      13'h827: dout = 8'b10111011;
      13'h828: dout = 8'b10111011;
      13'h829: dout = 8'b10111011;
      13'h82A: dout = 8'b10111011;
      13'h82B: dout = 8'b10111011;
      13'h82C: dout = 8'b10111011;
      13'h82D: dout = 8'b10111011;
      13'h82E: dout = 8'b10111011;
      13'h82F: dout = 8'b10111011;
      13'h830: dout = 8'b10111011;
      13'h831: dout = 8'b10111011;
      13'h832: dout = 8'b10111011;
      13'h833: dout = 8'b10111011;
      13'h834: dout = 8'b10111011;
      13'h835: dout = 8'b11100000;
      13'h836: dout = 8'b11100000;
      13'h837: dout = 8'b11100000;
      13'h838: dout = 8'b11100000;
      13'h839: dout = 8'b11100000;
      13'h83A: dout = 8'b11100000;
      13'h83B: dout = 8'b11100000;
      13'h83C: dout = 8'b11100000;
      13'h83D: dout = 8'b11100000;
      13'h83E: dout = 8'b11100000;
      13'h83F: dout = 8'b11100000;
      13'h840: dout = 8'b11100000;
      13'h841: dout = 8'b11100000;
      13'h842: dout = 8'b11100000;
      13'h843: dout = 8'b11100000;
      13'h844: dout = 8'b11100000;
      13'h845: dout = 8'b11100000;
      13'h846: dout = 8'b11100000;
      13'h847: dout = 8'b11100000;
      13'h848: dout = 8'b11100000;
      13'h849: dout = 8'b11100000;
      13'h84A: dout = 8'b11100000;
      13'h84B: dout = 8'b10111011;
      13'h84C: dout = 8'b10111011;
      13'h84D: dout = 8'b10111011;
      13'h84E: dout = 8'b10111011;
      13'h84F: dout = 8'b10111011;
      13'h850: dout = 8'b10111011;
      13'h851: dout = 8'b10111011;
      13'h852: dout = 8'b10111011;
      13'h853: dout = 8'b10111011;
      13'h854: dout = 8'b10111011;
      13'h855: dout = 8'b10111011;
      13'h856: dout = 8'b10111011;
      13'h857: dout = 8'b10111011;
      13'h858: dout = 8'b10111011;
      13'h859: dout = 8'b10111011;
      13'h85A: dout = 8'b10111011;
      13'h85B: dout = 8'b10111011;
      13'h85C: dout = 8'b10111011;
      13'h85D: dout = 8'b10111011;
      13'h85E: dout = 8'b10111011;
      13'h85F: dout = 8'b10111011;
      13'h860: dout = 8'b10111011;
      13'h861: dout = 8'b10111011;
      13'h862: dout = 8'b10111011;
      13'h863: dout = 8'b10111011;
      13'h864: dout = 8'b10111011;
      13'h865: dout = 8'b10111011;
      13'h866: dout = 8'b10111011;
      13'h867: dout = 8'b10111011;
      13'h868: dout = 8'b10111011;
      13'h869: dout = 8'b10111011;
      13'h86A: dout = 8'b10111011;
      13'h86B: dout = 8'b10111011;
      13'h86C: dout = 8'b10111011;
      13'h86D: dout = 8'b10111011;
      13'h86E: dout = 8'b10111011;
      13'h86F: dout = 8'b10111011;
      13'h870: dout = 8'b10111011;
      13'h871: dout = 8'b10111011;
      13'h872: dout = 8'b10111011;
      13'h873: dout = 8'b10111011;
      13'h874: dout = 8'b10111011;
      13'h875: dout = 8'b10111011;
      13'h876: dout = 8'b10111011;
      13'h877: dout = 8'b10111011;
      13'h878: dout = 8'b10111011;
      13'h879: dout = 8'b10111011;
      13'h87A: dout = 8'b10111011;
      13'h87B: dout = 8'b10111011;
      13'h87C: dout = 8'b10111011;
      13'h87D: dout = 8'b10111011;
      13'h87E: dout = 8'b10111011;
      13'h87F: dout = 8'b10111011;
      13'h880: dout = 8'b10111011;
      13'h881: dout = 8'b10111011;
      13'h882: dout = 8'b10111011;
      13'h883: dout = 8'b10111011;
      13'h884: dout = 8'b10111011;
      13'h885: dout = 8'b11100000;
      13'h886: dout = 8'b11100000;
      13'h887: dout = 8'b11100000;
      13'h888: dout = 8'b11100000;
      13'h889: dout = 8'b11100000;
      13'h88A: dout = 8'b11100000;
      13'h88B: dout = 8'b11100000;
      13'h88C: dout = 8'b11100000;
      13'h88D: dout = 8'b11100000;
      13'h88E: dout = 8'b11100000;
      13'h88F: dout = 8'b11100000;
      13'h890: dout = 8'b11100000;
      13'h891: dout = 8'b11100000;
      13'h892: dout = 8'b11100000;
      13'h893: dout = 8'b11100000;
      13'h894: dout = 8'b11100000;
      13'h895: dout = 8'b11100000;
      13'h896: dout = 8'b11100000;
      13'h897: dout = 8'b11100000;
      13'h898: dout = 8'b11100000;
      13'h899: dout = 8'b11100000;
      13'h89A: dout = 8'b11100000;
      13'h89B: dout = 8'b10111011;
      13'h89C: dout = 8'b10111011;
      13'h89D: dout = 8'b10111011;
      13'h89E: dout = 8'b10111011;
      13'h89F: dout = 8'b10111011;
      13'h8A0: dout = 8'b10111011;
      13'h8A1: dout = 8'b10111011;
      13'h8A2: dout = 8'b10111011;
      13'h8A3: dout = 8'b10111011;
      13'h8A4: dout = 8'b10111011;
      13'h8A5: dout = 8'b10111011;
      13'h8A6: dout = 8'b10111011;
      13'h8A7: dout = 8'b10111011;
      13'h8A8: dout = 8'b10111011;
      13'h8A9: dout = 8'b10111011;
      13'h8AA: dout = 8'b10111011;
      13'h8AB: dout = 8'b10111011;
      13'h8AC: dout = 8'b10111011;
      13'h8AD: dout = 8'b10111011;
      13'h8AE: dout = 8'b10111011;
      13'h8AF: dout = 8'b10111011;
      13'h8B0: dout = 8'b10111011;
      13'h8B1: dout = 8'b10111011;
      13'h8B2: dout = 8'b10111011;
      13'h8B3: dout = 8'b10111011;
      13'h8B4: dout = 8'b10111011;
      13'h8B5: dout = 8'b10111011;
      13'h8B6: dout = 8'b10111011;
      13'h8B7: dout = 8'b10111011;
      13'h8B8: dout = 8'b10111011;
      13'h8B9: dout = 8'b10111011;
      13'h8BA: dout = 8'b10111011;
      13'h8BB: dout = 8'b10111011;
      13'h8BC: dout = 8'b10111011;
      13'h8BD: dout = 8'b10111011;
      13'h8BE: dout = 8'b10111011;
      13'h8BF: dout = 8'b10111011;
      13'h8C0: dout = 8'b10111011;
      13'h8C1: dout = 8'b10111011;
      13'h8C2: dout = 8'b10111011;
      13'h8C3: dout = 8'b10111011;
      13'h8C4: dout = 8'b10111011;
      13'h8C5: dout = 8'b10111011;
      13'h8C6: dout = 8'b10111011;
      13'h8C7: dout = 8'b10111011;
      13'h8C8: dout = 8'b10111011;
      13'h8C9: dout = 8'b10111011;
      13'h8CA: dout = 8'b10111011;
      13'h8CB: dout = 8'b10111011;
      13'h8CC: dout = 8'b10111011;
      13'h8CD: dout = 8'b10111011;
      13'h8CE: dout = 8'b10111011;
      13'h8CF: dout = 8'b10111011;
      13'h8D0: dout = 8'b10111011;
      13'h8D1: dout = 8'b10111011;
      13'h8D2: dout = 8'b10111011;
      13'h8D3: dout = 8'b10111011;
      13'h8D4: dout = 8'b10111011;
      13'h8D5: dout = 8'b11100000;
      13'h8D6: dout = 8'b11100000;
      13'h8D7: dout = 8'b11100000;
      13'h8D8: dout = 8'b11100000;
      13'h8D9: dout = 8'b11100000;
      13'h8DA: dout = 8'b11100000;
      13'h8DB: dout = 8'b11100000;
      13'h8DC: dout = 8'b11100000;
      13'h8DD: dout = 8'b11100000;
      13'h8DE: dout = 8'b11100000;
      13'h8DF: dout = 8'b11100000;
      13'h8E0: dout = 8'b11100000;
      13'h8E1: dout = 8'b11100000;
      13'h8E2: dout = 8'b11100000;
      13'h8E3: dout = 8'b11100000;
      13'h8E4: dout = 8'b11100000;
      13'h8E5: dout = 8'b11100000;
      13'h8E6: dout = 8'b11100000;
      13'h8E7: dout = 8'b11100000;
      13'h8E8: dout = 8'b11100000;
      13'h8E9: dout = 8'b11100000;
      13'h8EA: dout = 8'b11100000;
      13'h8EB: dout = 8'b10111011;
      13'h8EC: dout = 8'b10111011;
      13'h8ED: dout = 8'b10111011;
      13'h8EE: dout = 8'b10111011;
      13'h8EF: dout = 8'b10111011;
      13'h8F0: dout = 8'b10111011;
      13'h8F1: dout = 8'b10111011;
      13'h8F2: dout = 8'b10111011;
      13'h8F3: dout = 8'b10111011;
      13'h8F4: dout = 8'b10111011;
      13'h8F5: dout = 8'b10111011;
      13'h8F6: dout = 8'b10111011;
      13'h8F7: dout = 8'b10111011;
      13'h8F8: dout = 8'b10111011;
      13'h8F9: dout = 8'b10111011;
      13'h8FA: dout = 8'b10111011;
      13'h8FB: dout = 8'b10111011;
      13'h8FC: dout = 8'b10111011;
      13'h8FD: dout = 8'b10111011;
      13'h8FE: dout = 8'b10111011;
      13'h8FF: dout = 8'b10111011;
      13'h900: dout = 8'b10111011;
      13'h901: dout = 8'b10111011;
      13'h902: dout = 8'b10111011;
      13'h903: dout = 8'b10111011;
      13'h904: dout = 8'b10111011;
      13'h905: dout = 8'b10111011;
      13'h906: dout = 8'b10111011;
      13'h907: dout = 8'b10111011;
      13'h908: dout = 8'b10111011;
      13'h909: dout = 8'b10111011;
      13'h90A: dout = 8'b10111011;
      13'h90B: dout = 8'b10111011;
      13'h90C: dout = 8'b10111011;
      13'h90D: dout = 8'b10111011;
      13'h90E: dout = 8'b10111011;
      13'h90F: dout = 8'b10111011;
      13'h910: dout = 8'b10111011;
      13'h911: dout = 8'b10111011;
      13'h912: dout = 8'b10111011;
      13'h913: dout = 8'b10111011;
      13'h914: dout = 8'b10111011;
      13'h915: dout = 8'b10111011;
      13'h916: dout = 8'b10111011;
      13'h917: dout = 8'b10111011;
      13'h918: dout = 8'b10111011;
      13'h919: dout = 8'b10111011;
      13'h91A: dout = 8'b10111011;
      13'h91B: dout = 8'b10111011;
      13'h91C: dout = 8'b10111011;
      13'h91D: dout = 8'b10111011;
      13'h91E: dout = 8'b10111011;
      13'h91F: dout = 8'b10111011;
      13'h920: dout = 8'b10111011;
      13'h921: dout = 8'b10111011;
      13'h922: dout = 8'b10111011;
      13'h923: dout = 8'b10111011;
      13'h924: dout = 8'b10111011;
      13'h925: dout = 8'b11100000;
      13'h926: dout = 8'b11100000;
      13'h927: dout = 8'b11100000;
      13'h928: dout = 8'b11100000;
      13'h929: dout = 8'b11100000;
      13'h92A: dout = 8'b11100000;
      13'h92B: dout = 8'b11100000;
      13'h92C: dout = 8'b11100000;
      13'h92D: dout = 8'b11100000;
      13'h92E: dout = 8'b11100000;
      13'h92F: dout = 8'b11100000;
      13'h930: dout = 8'b11100000;
      13'h931: dout = 8'b11100000;
      13'h932: dout = 8'b11100000;
      13'h933: dout = 8'b11100000;
      13'h934: dout = 8'b11100000;
      13'h935: dout = 8'b11100000;
      13'h936: dout = 8'b11100000;
      13'h937: dout = 8'b11100000;
      13'h938: dout = 8'b11100000;
      13'h939: dout = 8'b11100000;
      13'h93A: dout = 8'b11100000;
      13'h93B: dout = 8'b10111011;
      13'h93C: dout = 8'b10111011;
      13'h93D: dout = 8'b10111011;
      13'h93E: dout = 8'b10111011;
      13'h93F: dout = 8'b10111011;
      13'h940: dout = 8'b10111011;
      13'h941: dout = 8'b10111011;
      13'h942: dout = 8'b10111011;
      13'h943: dout = 8'b10111011;
      13'h944: dout = 8'b10111011;
      13'h945: dout = 8'b10111011;
      13'h946: dout = 8'b10111011;
      13'h947: dout = 8'b10111011;
      13'h948: dout = 8'b10111011;
      13'h949: dout = 8'b10111011;
      13'h94A: dout = 8'b10111011;
      13'h94B: dout = 8'b10111011;
      13'h94C: dout = 8'b10111011;
      13'h94D: dout = 8'b10111011;
      13'h94E: dout = 8'b10111011;
      13'h94F: dout = 8'b10111011;
      13'h950: dout = 8'b10111011;
      13'h951: dout = 8'b10111011;
      13'h952: dout = 8'b10111011;
      13'h953: dout = 8'b10111011;
      13'h954: dout = 8'b10111011;
      13'h955: dout = 8'b10111011;
      13'h956: dout = 8'b10111011;
      13'h957: dout = 8'b10111011;
      13'h958: dout = 8'b10111011;
      13'h959: dout = 8'b10111011;
      13'h95A: dout = 8'b10111011;
      13'h95B: dout = 8'b10111011;
      13'h95C: dout = 8'b10111011;
      13'h95D: dout = 8'b10111011;
      13'h95E: dout = 8'b10111011;
      13'h95F: dout = 8'b10111011;
      13'h960: dout = 8'b10111011;
      13'h961: dout = 8'b10111011;
      13'h962: dout = 8'b10111011;
      13'h963: dout = 8'b10111011;
      13'h964: dout = 8'b10111011;
      13'h965: dout = 8'b10111011;
      13'h966: dout = 8'b10111011;
      13'h967: dout = 8'b10111011;
      13'h968: dout = 8'b10111011;
      13'h969: dout = 8'b10111011;
      13'h96A: dout = 8'b10111011;
      13'h96B: dout = 8'b10111011;
      13'h96C: dout = 8'b10111011;
      13'h96D: dout = 8'b10111011;
      13'h96E: dout = 8'b10111011;
      13'h96F: dout = 8'b10111011;
      13'h970: dout = 8'b10111011;
      13'h971: dout = 8'b10111011;
      13'h972: dout = 8'b10111011;
      13'h973: dout = 8'b10111011;
      13'h974: dout = 8'b10111011;
      13'h975: dout = 8'b11100000;
      13'h976: dout = 8'b11100000;
      13'h977: dout = 8'b11100000;
      13'h978: dout = 8'b11100000;
      13'h979: dout = 8'b11100000;
      13'h97A: dout = 8'b11100000;
      13'h97B: dout = 8'b11100000;
      13'h97C: dout = 8'b11100000;
      13'h97D: dout = 8'b11100000;
      13'h97E: dout = 8'b11100000;
      13'h97F: dout = 8'b11100000;
      13'h980: dout = 8'b11100000;
      13'h981: dout = 8'b11100000;
      13'h982: dout = 8'b11100000;
      13'h983: dout = 8'b11100000;
      13'h984: dout = 8'b11100000;
      13'h985: dout = 8'b11100000;
      13'h986: dout = 8'b11100000;
      13'h987: dout = 8'b11100000;
      13'h988: dout = 8'b11100000;
      13'h989: dout = 8'b11100000;
      13'h98A: dout = 8'b11100000;
      13'h98B: dout = 8'b10111011;
      13'h98C: dout = 8'b10111011;
      13'h98D: dout = 8'b10111011;
      13'h98E: dout = 8'b10111011;
      13'h98F: dout = 8'b10111011;
      13'h990: dout = 8'b10111011;
      13'h991: dout = 8'b10111011;
      13'h992: dout = 8'b10111011;
      13'h993: dout = 8'b10111011;
      13'h994: dout = 8'b10111011;
      13'h995: dout = 8'b10111011;
      13'h996: dout = 8'b10111011;
      13'h997: dout = 8'b10111011;
      13'h998: dout = 8'b10111011;
      13'h999: dout = 8'b10111011;
      13'h99A: dout = 8'b10111011;
      13'h99B: dout = 8'b10111011;
      13'h99C: dout = 8'b10111011;
      13'h99D: dout = 8'b10111011;
      13'h99E: dout = 8'b10111011;
      13'h99F: dout = 8'b10111011;
      13'h9A0: dout = 8'b10111011;
      13'h9A1: dout = 8'b10111011;
      13'h9A2: dout = 8'b10111011;
      13'h9A3: dout = 8'b10111011;
      13'h9A4: dout = 8'b10111011;
      13'h9A5: dout = 8'b10111011;
      13'h9A6: dout = 8'b10111011;
      13'h9A7: dout = 8'b10111011;
      13'h9A8: dout = 8'b10111011;
      13'h9A9: dout = 8'b10111011;
      13'h9AA: dout = 8'b10111011;
      13'h9AB: dout = 8'b10111011;
      13'h9AC: dout = 8'b10111011;
      13'h9AD: dout = 8'b10111011;
      13'h9AE: dout = 8'b10111011;
      13'h9AF: dout = 8'b10111011;
      13'h9B0: dout = 8'b10111011;
      13'h9B1: dout = 8'b10111011;
      13'h9B2: dout = 8'b10111011;
      13'h9B3: dout = 8'b10111011;
      13'h9B4: dout = 8'b10111011;
      13'h9B5: dout = 8'b10111011;
      13'h9B6: dout = 8'b10111011;
      13'h9B7: dout = 8'b10111011;
      13'h9B8: dout = 8'b10111011;
      13'h9B9: dout = 8'b10111011;
      13'h9BA: dout = 8'b10111011;
      13'h9BB: dout = 8'b10111011;
      13'h9BC: dout = 8'b10111011;
      13'h9BD: dout = 8'b10111011;
      13'h9BE: dout = 8'b10111011;
      13'h9BF: dout = 8'b10111011;
      13'h9C0: dout = 8'b10111011;
      13'h9C1: dout = 8'b10111011;
      13'h9C2: dout = 8'b10111011;
      13'h9C3: dout = 8'b10111011;
      13'h9C4: dout = 8'b10111011;
      13'h9C5: dout = 8'b11100000;
      13'h9C6: dout = 8'b11100000;
      13'h9C7: dout = 8'b11100000;
      13'h9C8: dout = 8'b11100000;
      13'h9C9: dout = 8'b11100000;
      13'h9CA: dout = 8'b11100000;
      13'h9CB: dout = 8'b11100000;
      13'h9CC: dout = 8'b11100000;
      13'h9CD: dout = 8'b11100000;
      13'h9CE: dout = 8'b11100000;
      13'h9CF: dout = 8'b11100000;
      13'h9D0: dout = 8'b11100000;
      13'h9D1: dout = 8'b11100000;
      13'h9D2: dout = 8'b11100000;
      13'h9D3: dout = 8'b11100000;
      13'h9D4: dout = 8'b11100000;
      13'h9D5: dout = 8'b11100000;
      13'h9D6: dout = 8'b11100000;
      13'h9D7: dout = 8'b11100000;
      13'h9D8: dout = 8'b11100000;
      13'h9D9: dout = 8'b11100000;
      13'h9DA: dout = 8'b11100000;
      13'h9DB: dout = 8'b10111011;
      13'h9DC: dout = 8'b10111011;
      13'h9DD: dout = 8'b10111011;
      13'h9DE: dout = 8'b10111011;
      13'h9DF: dout = 8'b10111011;
      13'h9E0: dout = 8'b10111011;
      13'h9E1: dout = 8'b10111011;
      13'h9E2: dout = 8'b10111011;
      13'h9E3: dout = 8'b10111011;
      13'h9E4: dout = 8'b10111011;
      13'h9E5: dout = 8'b10111011;
      13'h9E6: dout = 8'b10111011;
      13'h9E7: dout = 8'b10111011;
      13'h9E8: dout = 8'b10111011;
      13'h9E9: dout = 8'b10111011;
      13'h9EA: dout = 8'b10111011;
      13'h9EB: dout = 8'b10111011;
      13'h9EC: dout = 8'b10111011;
      13'h9ED: dout = 8'b10111011;
      13'h9EE: dout = 8'b10111011;
      13'h9EF: dout = 8'b10111011;
      13'h9F0: dout = 8'b10111011;
      13'h9F1: dout = 8'b10111011;
      13'h9F2: dout = 8'b10111011;
      13'h9F3: dout = 8'b10111011;
      13'h9F4: dout = 8'b10111011;
      13'h9F5: dout = 8'b10111011;
      13'h9F6: dout = 8'b10111011;
      13'h9F7: dout = 8'b10111011;
      13'h9F8: dout = 8'b10111011;
      13'h9F9: dout = 8'b10111011;
      13'h9FA: dout = 8'b10111011;
      13'h9FB: dout = 8'b10111011;
      13'h9FC: dout = 8'b10111011;
      13'h9FD: dout = 8'b10111011;
      13'h9FE: dout = 8'b10111011;
      13'h9FF: dout = 8'b10111011;
      13'hA00: dout = 8'b10111011;
      13'hA01: dout = 8'b10111011;
      13'hA02: dout = 8'b10111011;
      13'hA03: dout = 8'b10111011;
      13'hA04: dout = 8'b10111011;
      13'hA05: dout = 8'b10111011;
      13'hA06: dout = 8'b10111011;
      13'hA07: dout = 8'b10111011;
      13'hA08: dout = 8'b10111011;
      13'hA09: dout = 8'b10111011;
      13'hA0A: dout = 8'b10111011;
      13'hA0B: dout = 8'b10111011;
      13'hA0C: dout = 8'b10111011;
      13'hA0D: dout = 8'b10111011;
      13'hA0E: dout = 8'b10111011;
      13'hA0F: dout = 8'b10111011;
      13'hA10: dout = 8'b10111011;
      13'hA11: dout = 8'b10111011;
      13'hA12: dout = 8'b10111011;
      13'hA13: dout = 8'b10111011;
      13'hA14: dout = 8'b10111011;
      13'hA15: dout = 8'b11100000;
      13'hA16: dout = 8'b11100000;
      13'hA17: dout = 8'b11100000;
      13'hA18: dout = 8'b11100000;
      13'hA19: dout = 8'b11100000;
      13'hA1A: dout = 8'b11100000;
      13'hA1B: dout = 8'b11100000;
      13'hA1C: dout = 8'b11100000;
      13'hA1D: dout = 8'b11100000;
      13'hA1E: dout = 8'b11100000;
      13'hA1F: dout = 8'b11100000;
      13'hA20: dout = 8'b11100000;
      13'hA21: dout = 8'b11100000;
      13'hA22: dout = 8'b11100000;
      13'hA23: dout = 8'b11100000;
      13'hA24: dout = 8'b11100000;
      13'hA25: dout = 8'b11100000;
      13'hA26: dout = 8'b11100000;
      13'hA27: dout = 8'b11100000;
      13'hA28: dout = 8'b11100000;
      13'hA29: dout = 8'b11100000;
      13'hA2A: dout = 8'b11100000;
      13'hA2B: dout = 8'b10111011;
      13'hA2C: dout = 8'b10111011;
      13'hA2D: dout = 8'b10111011;
      13'hA2E: dout = 8'b10111011;
      13'hA2F: dout = 8'b10111011;
      13'hA30: dout = 8'b10111011;
      13'hA31: dout = 8'b10111011;
      13'hA32: dout = 8'b10111011;
      13'hA33: dout = 8'b10111011;
      13'hA34: dout = 8'b10111011;
      13'hA35: dout = 8'b10111011;
      13'hA36: dout = 8'b10111011;
      13'hA37: dout = 8'b10111011;
      13'hA38: dout = 8'b10111011;
      13'hA39: dout = 8'b10111011;
      13'hA3A: dout = 8'b10111011;
      13'hA3B: dout = 8'b10111011;
      13'hA3C: dout = 8'b10111011;
      13'hA3D: dout = 8'b10111011;
      13'hA3E: dout = 8'b10111011;
      13'hA3F: dout = 8'b10111011;
      13'hA40: dout = 8'b10111011;
      13'hA41: dout = 8'b10111011;
      13'hA42: dout = 8'b10111011;
      13'hA43: dout = 8'b10111011;
      13'hA44: dout = 8'b10111011;
      13'hA45: dout = 8'b10111011;
      13'hA46: dout = 8'b10111011;
      13'hA47: dout = 8'b10111011;
      13'hA48: dout = 8'b10111011;
      13'hA49: dout = 8'b10111011;
      13'hA4A: dout = 8'b10111011;
      13'hA4B: dout = 8'b10111011;
      13'hA4C: dout = 8'b10111011;
      13'hA4D: dout = 8'b10111011;
      13'hA4E: dout = 8'b10111011;
      13'hA4F: dout = 8'b10111011;
      13'hA50: dout = 8'b10111011;
      13'hA51: dout = 8'b10111011;
      13'hA52: dout = 8'b10111011;
      13'hA53: dout = 8'b10111011;
      13'hA54: dout = 8'b10111011;
      13'hA55: dout = 8'b10111011;
      13'hA56: dout = 8'b10111011;
      13'hA57: dout = 8'b10111011;
      13'hA58: dout = 8'b10111011;
      13'hA59: dout = 8'b10111011;
      13'hA5A: dout = 8'b10111011;
      13'hA5B: dout = 8'b10111011;
      13'hA5C: dout = 8'b10111011;
      13'hA5D: dout = 8'b10111011;
      13'hA5E: dout = 8'b10111011;
      13'hA5F: dout = 8'b10111011;
      13'hA60: dout = 8'b10111011;
      13'hA61: dout = 8'b10111011;
      13'hA62: dout = 8'b10111011;
      13'hA63: dout = 8'b10111011;
      13'hA64: dout = 8'b10111011;
      13'hA65: dout = 8'b11100000;
      13'hA66: dout = 8'b11100000;
      13'hA67: dout = 8'b11100000;
      13'hA68: dout = 8'b11100000;
      13'hA69: dout = 8'b11100000;
      13'hA6A: dout = 8'b11100000;
      13'hA6B: dout = 8'b11100000;
      13'hA6C: dout = 8'b11100000;
      13'hA6D: dout = 8'b11100000;
      13'hA6E: dout = 8'b11100000;
      13'hA6F: dout = 8'b11100000;
      13'hA70: dout = 8'b11100000;
      13'hA71: dout = 8'b11100000;
      13'hA72: dout = 8'b11100000;
      13'hA73: dout = 8'b11100000;
      13'hA74: dout = 8'b11100000;
      13'hA75: dout = 8'b11100000;
      13'hA76: dout = 8'b11100000;
      13'hA77: dout = 8'b11100000;
      13'hA78: dout = 8'b11100000;
      13'hA79: dout = 8'b11100000;
      13'hA7A: dout = 8'b11100000;
      13'hA7B: dout = 8'b10111011;
      13'hA7C: dout = 8'b10111011;
      13'hA7D: dout = 8'b10111011;
      13'hA7E: dout = 8'b10111011;
      13'hA7F: dout = 8'b10111011;
      13'hA80: dout = 8'b10111011;
      13'hA81: dout = 8'b10111011;
      13'hA82: dout = 8'b10111011;
      13'hA83: dout = 8'b10111011;
      13'hA84: dout = 8'b10111011;
      13'hA85: dout = 8'b10111011;
      13'hA86: dout = 8'b10111011;
      13'hA87: dout = 8'b10111011;
      13'hA88: dout = 8'b10111011;
      13'hA89: dout = 8'b10111011;
      13'hA8A: dout = 8'b10111011;
      13'hA8B: dout = 8'b10111011;
      13'hA8C: dout = 8'b10111011;
      13'hA8D: dout = 8'b10111011;
      13'hA8E: dout = 8'b10111011;
      13'hA8F: dout = 8'b10111011;
      13'hA90: dout = 8'b10111011;
      13'hA91: dout = 8'b10111011;
      13'hA92: dout = 8'b10111011;
      13'hA93: dout = 8'b10111011;
      13'hA94: dout = 8'b10111011;
      13'hA95: dout = 8'b10111011;
      13'hA96: dout = 8'b10111011;
      13'hA97: dout = 8'b10111011;
      13'hA98: dout = 8'b10111011;
      13'hA99: dout = 8'b10111011;
      13'hA9A: dout = 8'b10111011;
      13'hA9B: dout = 8'b10111011;
      13'hA9C: dout = 8'b10111011;
      13'hA9D: dout = 8'b10111011;
      13'hA9E: dout = 8'b10111011;
      13'hA9F: dout = 8'b10111011;
      13'hAA0: dout = 8'b10111011;
      13'hAA1: dout = 8'b10111011;
      13'hAA2: dout = 8'b10111011;
      13'hAA3: dout = 8'b10111011;
      13'hAA4: dout = 8'b10111011;
      13'hAA5: dout = 8'b10111011;
      13'hAA6: dout = 8'b10111011;
      13'hAA7: dout = 8'b10111011;
      13'hAA8: dout = 8'b10111011;
      13'hAA9: dout = 8'b10111011;
      13'hAAA: dout = 8'b10111011;
      13'hAAB: dout = 8'b10111011;
      13'hAAC: dout = 8'b10111011;
      13'hAAD: dout = 8'b10111011;
      13'hAAE: dout = 8'b10111011;
      13'hAAF: dout = 8'b10111011;
      13'hAB0: dout = 8'b10111011;
      13'hAB1: dout = 8'b10111011;
      13'hAB2: dout = 8'b10111011;
      13'hAB3: dout = 8'b10111011;
      13'hAB4: dout = 8'b10111011;
      13'hAB5: dout = 8'b11100000;
      13'hAB6: dout = 8'b11100000;
      13'hAB7: dout = 8'b11100000;
      13'hAB8: dout = 8'b11100000;
      13'hAB9: dout = 8'b11100000;
      13'hABA: dout = 8'b11100000;
      13'hABB: dout = 8'b11100000;
      13'hABC: dout = 8'b11100000;
      13'hABD: dout = 8'b11100000;
      13'hABE: dout = 8'b11100000;
      13'hABF: dout = 8'b11100000;
      13'hAC0: dout = 8'b11100000;
      13'hAC1: dout = 8'b11100000;
      13'hAC2: dout = 8'b11100000;
      13'hAC3: dout = 8'b11100000;
      13'hAC4: dout = 8'b11100000;
      13'hAC5: dout = 8'b11100000;
      13'hAC6: dout = 8'b11100000;
      13'hAC7: dout = 8'b11100000;
      13'hAC8: dout = 8'b11100000;
      13'hAC9: dout = 8'b11100000;
      13'hACA: dout = 8'b11100000;
      13'hACB: dout = 8'b10111011;
      13'hACC: dout = 8'b10111011;
      13'hACD: dout = 8'b10111011;
      13'hACE: dout = 8'b10111011;
      13'hACF: dout = 8'b10111011;
      13'hAD0: dout = 8'b10111011;
      13'hAD1: dout = 8'b10111011;
      13'hAD2: dout = 8'b10111011;
      13'hAD3: dout = 8'b10111011;
      13'hAD4: dout = 8'b10111011;
      13'hAD5: dout = 8'b10111011;
      13'hAD6: dout = 8'b10111011;
      13'hAD7: dout = 8'b10111011;
      13'hAD8: dout = 8'b10111011;
      13'hAD9: dout = 8'b10111011;
      13'hADA: dout = 8'b10111011;
      13'hADB: dout = 8'b10111011;
      13'hADC: dout = 8'b10111011;
      13'hADD: dout = 8'b10111011;
      13'hADE: dout = 8'b10111011;
      13'hADF: dout = 8'b10111011;
      13'hAE0: dout = 8'b10111011;
      13'hAE1: dout = 8'b10111011;
      13'hAE2: dout = 8'b10111011;
      13'hAE3: dout = 8'b10111011;
      13'hAE4: dout = 8'b10111011;
      13'hAE5: dout = 8'b10111011;
      13'hAE6: dout = 8'b10111011;
      13'hAE7: dout = 8'b10111011;
      13'hAE8: dout = 8'b10111011;
      13'hAE9: dout = 8'b10111011;
      13'hAEA: dout = 8'b10111011;
      13'hAEB: dout = 8'b10111011;
      13'hAEC: dout = 8'b10111011;
      13'hAED: dout = 8'b10111011;
      13'hAEE: dout = 8'b10111011;
      13'hAEF: dout = 8'b10111011;
      13'hAF0: dout = 8'b10111011;
      13'hAF1: dout = 8'b10111011;
      13'hAF2: dout = 8'b10111011;
      13'hAF3: dout = 8'b10111011;
      13'hAF4: dout = 8'b10111011;
      13'hAF5: dout = 8'b10111011;
      13'hAF6: dout = 8'b10111011;
      13'hAF7: dout = 8'b10111011;
      13'hAF8: dout = 8'b10111011;
      13'hAF9: dout = 8'b10111011;
      13'hAFA: dout = 8'b10111011;
      13'hAFB: dout = 8'b10111011;
      13'hAFC: dout = 8'b10111011;
      13'hAFD: dout = 8'b10111011;
      13'hAFE: dout = 8'b10111011;
      13'hAFF: dout = 8'b10111011;
      13'hB00: dout = 8'b10111011;
      13'hB01: dout = 8'b10111011;
      13'hB02: dout = 8'b10111011;
      13'hB03: dout = 8'b10111011;
      13'hB04: dout = 8'b10111011;
      13'hB05: dout = 8'b11100000;
      13'hB06: dout = 8'b11100000;
      13'hB07: dout = 8'b11100000;
      13'hB08: dout = 8'b11100000;
      13'hB09: dout = 8'b11100000;
      13'hB0A: dout = 8'b11100000;
      13'hB0B: dout = 8'b11100000;
      13'hB0C: dout = 8'b11100000;
      13'hB0D: dout = 8'b11100000;
      13'hB0E: dout = 8'b11100000;
      13'hB0F: dout = 8'b11100000;
      13'hB10: dout = 8'b11100000;
      13'hB11: dout = 8'b11100000;
      13'hB12: dout = 8'b11100000;
      13'hB13: dout = 8'b11100000;
      13'hB14: dout = 8'b11100000;
      13'hB15: dout = 8'b11100000;
      13'hB16: dout = 8'b11100000;
      13'hB17: dout = 8'b11100000;
      13'hB18: dout = 8'b11100000;
      13'hB19: dout = 8'b11100000;
      13'hB1A: dout = 8'b11100000;
      13'hB1B: dout = 8'b10111011;
      13'hB1C: dout = 8'b10111011;
      13'hB1D: dout = 8'b10111011;
      13'hB1E: dout = 8'b10111011;
      13'hB1F: dout = 8'b10111011;
      13'hB20: dout = 8'b10111011;
      13'hB21: dout = 8'b10111011;
      13'hB22: dout = 8'b10111011;
      13'hB23: dout = 8'b10111011;
      13'hB24: dout = 8'b10111011;
      13'hB25: dout = 8'b10111011;
      13'hB26: dout = 8'b10111011;
      13'hB27: dout = 8'b10111011;
      13'hB28: dout = 8'b10111011;
      13'hB29: dout = 8'b10111011;
      13'hB2A: dout = 8'b10111011;
      13'hB2B: dout = 8'b10111011;
      13'hB2C: dout = 8'b10111011;
      13'hB2D: dout = 8'b10111011;
      13'hB2E: dout = 8'b10111011;
      13'hB2F: dout = 8'b10111011;
      13'hB30: dout = 8'b10111011;
      13'hB31: dout = 8'b10111011;
      13'hB32: dout = 8'b10111011;
      13'hB33: dout = 8'b10111011;
      13'hB34: dout = 8'b10111011;
      13'hB35: dout = 8'b10111011;
      13'hB36: dout = 8'b10111011;
      13'hB37: dout = 8'b10111011;
      13'hB38: dout = 8'b10111011;
      13'hB39: dout = 8'b10111011;
      13'hB3A: dout = 8'b10111011;
      13'hB3B: dout = 8'b10111011;
      13'hB3C: dout = 8'b10111011;
      13'hB3D: dout = 8'b10111011;
      13'hB3E: dout = 8'b10111011;
      13'hB3F: dout = 8'b10111011;
      13'hB40: dout = 8'b10111011;
      13'hB41: dout = 8'b10111011;
      13'hB42: dout = 8'b10111011;
      13'hB43: dout = 8'b10111011;
      13'hB44: dout = 8'b10111011;
      13'hB45: dout = 8'b10111011;
      13'hB46: dout = 8'b10111011;
      13'hB47: dout = 8'b10111011;
      13'hB48: dout = 8'b10111011;
      13'hB49: dout = 8'b10111011;
      13'hB4A: dout = 8'b10111011;
      13'hB4B: dout = 8'b10111011;
      13'hB4C: dout = 8'b10111011;
      13'hB4D: dout = 8'b10111011;
      13'hB4E: dout = 8'b10111011;
      13'hB4F: dout = 8'b10111011;
      13'hB50: dout = 8'b10111011;
      13'hB51: dout = 8'b10111011;
      13'hB52: dout = 8'b10111011;
      13'hB53: dout = 8'b10111011;
      13'hB54: dout = 8'b10111011;
      13'hB55: dout = 8'b11100000;
      13'hB56: dout = 8'b11100000;
      13'hB57: dout = 8'b11100000;
      13'hB58: dout = 8'b11100000;
      13'hB59: dout = 8'b11100000;
      13'hB5A: dout = 8'b11100000;
      13'hB5B: dout = 8'b11100000;
      13'hB5C: dout = 8'b11100000;
      13'hB5D: dout = 8'b11100000;
      13'hB5E: dout = 8'b11100000;
      13'hB5F: dout = 8'b11100000;
      13'hB60: dout = 8'b11100000;
      13'hB61: dout = 8'b11100000;
      13'hB62: dout = 8'b11100000;
      13'hB63: dout = 8'b11100000;
      13'hB64: dout = 8'b11100000;
      13'hB65: dout = 8'b11100000;
      13'hB66: dout = 8'b11100000;
      13'hB67: dout = 8'b11100000;
      13'hB68: dout = 8'b11100000;
      13'hB69: dout = 8'b11100000;
      13'hB6A: dout = 8'b11100000;
      13'hB6B: dout = 8'b10111011;
      13'hB6C: dout = 8'b10111011;
      13'hB6D: dout = 8'b10111011;
      13'hB6E: dout = 8'b10111011;
      13'hB6F: dout = 8'b10111011;
      13'hB70: dout = 8'b10111011;
      13'hB71: dout = 8'b10111011;
      13'hB72: dout = 8'b10111011;
      13'hB73: dout = 8'b10111011;
      13'hB74: dout = 8'b10111011;
      13'hB75: dout = 8'b10111011;
      13'hB76: dout = 8'b10111011;
      13'hB77: dout = 8'b10111011;
      13'hB78: dout = 8'b10111011;
      13'hB79: dout = 8'b10111011;
      13'hB7A: dout = 8'b10111011;
      13'hB7B: dout = 8'b10111011;
      13'hB7C: dout = 8'b10111011;
      13'hB7D: dout = 8'b10111011;
      13'hB7E: dout = 8'b10111011;
      13'hB7F: dout = 8'b10111011;
      13'hB80: dout = 8'b10111011;
      13'hB81: dout = 8'b10111011;
      13'hB82: dout = 8'b10111011;
      13'hB83: dout = 8'b10111011;
      13'hB84: dout = 8'b10111011;
      13'hB85: dout = 8'b10111011;
      13'hB86: dout = 8'b10111011;
      13'hB87: dout = 8'b10111011;
      13'hB88: dout = 8'b10111011;
      13'hB89: dout = 8'b10111011;
      13'hB8A: dout = 8'b10111011;
      13'hB8B: dout = 8'b10111011;
      13'hB8C: dout = 8'b10111011;
      13'hB8D: dout = 8'b10111011;
      13'hB8E: dout = 8'b10111011;
      13'hB8F: dout = 8'b10111011;
      13'hB90: dout = 8'b10111011;
      13'hB91: dout = 8'b10111011;
      13'hB92: dout = 8'b10111011;
      13'hB93: dout = 8'b10111011;
      13'hB94: dout = 8'b10111011;
      13'hB95: dout = 8'b10111011;
      13'hB96: dout = 8'b10111011;
      13'hB97: dout = 8'b10111011;
      13'hB98: dout = 8'b10111011;
      13'hB99: dout = 8'b10111011;
      13'hB9A: dout = 8'b10111011;
      13'hB9B: dout = 8'b10111011;
      13'hB9C: dout = 8'b10111011;
      13'hB9D: dout = 8'b10111011;
      13'hB9E: dout = 8'b10111011;
      13'hB9F: dout = 8'b10111011;
      13'hBA0: dout = 8'b10111011;
      13'hBA1: dout = 8'b10111011;
      13'hBA2: dout = 8'b10111011;
      13'hBA3: dout = 8'b10111011;
      13'hBA4: dout = 8'b10111011;
      13'hBA5: dout = 8'b11100000;
      13'hBA6: dout = 8'b11100000;
      13'hBA7: dout = 8'b11100000;
      13'hBA8: dout = 8'b11100000;
      13'hBA9: dout = 8'b11100000;
      13'hBAA: dout = 8'b11100000;
      13'hBAB: dout = 8'b11100000;
      13'hBAC: dout = 8'b11100000;
      13'hBAD: dout = 8'b11100000;
      13'hBAE: dout = 8'b11100000;
      13'hBAF: dout = 8'b11100000;
      13'hBB0: dout = 8'b11100000;
      13'hBB1: dout = 8'b11100000;
      13'hBB2: dout = 8'b11100000;
      13'hBB3: dout = 8'b11100000;
      13'hBB4: dout = 8'b11100000;
      13'hBB5: dout = 8'b11100000;
      13'hBB6: dout = 8'b11100000;
      13'hBB7: dout = 8'b11100000;
      13'hBB8: dout = 8'b11100000;
      13'hBB9: dout = 8'b11100000;
      13'hBBA: dout = 8'b11100000;
      13'hBBB: dout = 8'b10111011;
      13'hBBC: dout = 8'b10111011;
      13'hBBD: dout = 8'b10111011;
      13'hBBE: dout = 8'b10111011;
      13'hBBF: dout = 8'b10111011;
      13'hBC0: dout = 8'b10111011;
      13'hBC1: dout = 8'b10111011;
      13'hBC2: dout = 8'b10111011;
      13'hBC3: dout = 8'b10111011;
      13'hBC4: dout = 8'b10111011;
      13'hBC5: dout = 8'b10111011;
      13'hBC6: dout = 8'b10111011;
      13'hBC7: dout = 8'b10111011;
      13'hBC8: dout = 8'b10111011;
      13'hBC9: dout = 8'b10111011;
      13'hBCA: dout = 8'b10111011;
      13'hBCB: dout = 8'b10111011;
      13'hBCC: dout = 8'b10111011;
      13'hBCD: dout = 8'b10111011;
      13'hBCE: dout = 8'b10111011;
      13'hBCF: dout = 8'b10111011;
      13'hBD0: dout = 8'b10111011;
      13'hBD1: dout = 8'b10111011;
      13'hBD2: dout = 8'b10111011;
      13'hBD3: dout = 8'b10111011;
      13'hBD4: dout = 8'b10111011;
      13'hBD5: dout = 8'b10111011;
      13'hBD6: dout = 8'b10111011;
      13'hBD7: dout = 8'b10111011;
      13'hBD8: dout = 8'b10111011;
      13'hBD9: dout = 8'b10111011;
      13'hBDA: dout = 8'b10111011;
      13'hBDB: dout = 8'b10111011;
      13'hBDC: dout = 8'b10111011;
      13'hBDD: dout = 8'b10111011;
      13'hBDE: dout = 8'b10111011;
      13'hBDF: dout = 8'b10111011;
      13'hBE0: dout = 8'b10111011;
      13'hBE1: dout = 8'b10111011;
      13'hBE2: dout = 8'b10111011;
      13'hBE3: dout = 8'b10111011;
      13'hBE4: dout = 8'b10111011;
      13'hBE5: dout = 8'b10111011;
      13'hBE6: dout = 8'b10111011;
      13'hBE7: dout = 8'b10111011;
      13'hBE8: dout = 8'b10111011;
      13'hBE9: dout = 8'b10111011;
      13'hBEA: dout = 8'b10111011;
      13'hBEB: dout = 8'b10111011;
      13'hBEC: dout = 8'b10111011;
      13'hBED: dout = 8'b10111011;
      13'hBEE: dout = 8'b10111011;
      13'hBEF: dout = 8'b10111011;
      13'hBF0: dout = 8'b10111011;
      13'hBF1: dout = 8'b10111011;
      13'hBF2: dout = 8'b10111011;
      13'hBF3: dout = 8'b10111011;
      13'hBF4: dout = 8'b10111011;
      13'hBF5: dout = 8'b11100000;
      13'hBF6: dout = 8'b11100000;
      13'hBF7: dout = 8'b11100000;
      13'hBF8: dout = 8'b11100000;
      13'hBF9: dout = 8'b11100000;
      13'hBFA: dout = 8'b11100000;
      13'hBFB: dout = 8'b11100000;
      13'hBFC: dout = 8'b11100000;
      13'hBFD: dout = 8'b11100000;
      13'hBFE: dout = 8'b11100000;
      13'hBFF: dout = 8'b11100000;
      13'hC00: dout = 8'b11100000;
      13'hC01: dout = 8'b11100000;
      13'hC02: dout = 8'b11100000;
      13'hC03: dout = 8'b11100000;
      13'hC04: dout = 8'b11100000;
      13'hC05: dout = 8'b11100000;
      13'hC06: dout = 8'b11100000;
      13'hC07: dout = 8'b11100000;
      13'hC08: dout = 8'b11100000;
      13'hC09: dout = 8'b11100000;
      13'hC0A: dout = 8'b11100000;
      13'hC0B: dout = 8'b10111011;
      13'hC0C: dout = 8'b10111011;
      13'hC0D: dout = 8'b10111011;
      13'hC0E: dout = 8'b10111011;
      13'hC0F: dout = 8'b10111011;
      13'hC10: dout = 8'b10111011;
      13'hC11: dout = 8'b10111011;
      13'hC12: dout = 8'b10111011;
      13'hC13: dout = 8'b10111011;
      13'hC14: dout = 8'b10111011;
      13'hC15: dout = 8'b10111011;
      13'hC16: dout = 8'b10111011;
      13'hC17: dout = 8'b10111011;
      13'hC18: dout = 8'b10111011;
      13'hC19: dout = 8'b10111011;
      13'hC1A: dout = 8'b10111011;
      13'hC1B: dout = 8'b10111011;
      13'hC1C: dout = 8'b10111011;
      13'hC1D: dout = 8'b10111011;
      13'hC1E: dout = 8'b10111011;
      13'hC1F: dout = 8'b10111011;
      13'hC20: dout = 8'b10111011;
      13'hC21: dout = 8'b10111011;
      13'hC22: dout = 8'b10111011;
      13'hC23: dout = 8'b10111011;
      13'hC24: dout = 8'b10111011;
      13'hC25: dout = 8'b10111011;
      13'hC26: dout = 8'b10111011;
      13'hC27: dout = 8'b10111011;
      13'hC28: dout = 8'b10111011;
      13'hC29: dout = 8'b10111011;
      13'hC2A: dout = 8'b10111011;
      13'hC2B: dout = 8'b10111011;
      13'hC2C: dout = 8'b10111011;
      13'hC2D: dout = 8'b10111011;
      13'hC2E: dout = 8'b10111011;
      13'hC2F: dout = 8'b10111011;
      13'hC30: dout = 8'b10111011;
      13'hC31: dout = 8'b10111011;
      13'hC32: dout = 8'b10111011;
      13'hC33: dout = 8'b10111011;
      13'hC34: dout = 8'b10111011;
      13'hC35: dout = 8'b10111011;
      13'hC36: dout = 8'b10111011;
      13'hC37: dout = 8'b10111011;
      13'hC38: dout = 8'b10111011;
      13'hC39: dout = 8'b10111011;
      13'hC3A: dout = 8'b10111011;
      13'hC3B: dout = 8'b10111011;
      13'hC3C: dout = 8'b10111011;
      13'hC3D: dout = 8'b10111011;
      13'hC3E: dout = 8'b10111011;
      13'hC3F: dout = 8'b10111011;
      13'hC40: dout = 8'b10111011;
      13'hC41: dout = 8'b10111011;
      13'hC42: dout = 8'b10111011;
      13'hC43: dout = 8'b10111011;
      13'hC44: dout = 8'b10111011;
      13'hC45: dout = 8'b10111011;
      13'hC46: dout = 8'b10111011;
      13'hC47: dout = 8'b10111011;
      13'hC48: dout = 8'b10111011;
      13'hC49: dout = 8'b10111011;
      13'hC4A: dout = 8'b10111011;
      13'hC4B: dout = 8'b10111011;
      13'hC4C: dout = 8'b10111011;
      13'hC4D: dout = 8'b10111011;
      13'hC4E: dout = 8'b10111011;
      13'hC4F: dout = 8'b10111011;
      13'hC50: dout = 8'b10111011;
      13'hC51: dout = 8'b10111011;
      13'hC52: dout = 8'b10111011;
      13'hC53: dout = 8'b10111011;
      13'hC54: dout = 8'b10111011;
      13'hC55: dout = 8'b10111011;
      13'hC56: dout = 8'b10111011;
      13'hC57: dout = 8'b10111011;
      13'hC58: dout = 8'b10111011;
      13'hC59: dout = 8'b10111011;
      13'hC5A: dout = 8'b10111011;
      13'hC5B: dout = 8'b10111011;
      13'hC5C: dout = 8'b10111011;
      13'hC5D: dout = 8'b10111011;
      13'hC5E: dout = 8'b10111011;
      13'hC5F: dout = 8'b10111011;
      13'hC60: dout = 8'b10111011;
      13'hC61: dout = 8'b10111011;
      13'hC62: dout = 8'b10111011;
      13'hC63: dout = 8'b10111011;
      13'hC64: dout = 8'b10111011;
      13'hC65: dout = 8'b10111011;
      13'hC66: dout = 8'b10111011;
      13'hC67: dout = 8'b10111011;
      13'hC68: dout = 8'b10111011;
      13'hC69: dout = 8'b10111011;
      13'hC6A: dout = 8'b10111011;
      13'hC6B: dout = 8'b10111011;
      13'hC6C: dout = 8'b10111011;
      13'hC6D: dout = 8'b10111011;
      13'hC6E: dout = 8'b10111011;
      13'hC6F: dout = 8'b10111011;
      13'hC70: dout = 8'b10111011;
      13'hC71: dout = 8'b10111011;
      13'hC72: dout = 8'b10111011;
      13'hC73: dout = 8'b10111011;
      13'hC74: dout = 8'b10111011;
      13'hC75: dout = 8'b10111011;
      13'hC76: dout = 8'b10111011;
      13'hC77: dout = 8'b10111011;
      13'hC78: dout = 8'b10111011;
      13'hC79: dout = 8'b10111011;
      13'hC7A: dout = 8'b10111011;
      13'hC7B: dout = 8'b10111011;
      13'hC7C: dout = 8'b10111011;
      13'hC7D: dout = 8'b10111011;
      13'hC7E: dout = 8'b10111011;
      13'hC7F: dout = 8'b10111011;
      13'hC80: dout = 8'b10111011;
      13'hC81: dout = 8'b10111011;
      13'hC82: dout = 8'b10111011;
      13'hC83: dout = 8'b10111011;
      13'hC84: dout = 8'b10111011;
      13'hC85: dout = 8'b10111011;
      13'hC86: dout = 8'b10111011;
      13'hC87: dout = 8'b10111011;
      13'hC88: dout = 8'b10111011;
      13'hC89: dout = 8'b10111011;
      13'hC8A: dout = 8'b10111011;
      13'hC8B: dout = 8'b10111011;
      13'hC8C: dout = 8'b10111011;
      13'hC8D: dout = 8'b10111011;
      13'hC8E: dout = 8'b10111011;
      13'hC8F: dout = 8'b10111011;
      13'hC90: dout = 8'b10111011;
      13'hC91: dout = 8'b10111011;
      13'hC92: dout = 8'b10111011;
      13'hC93: dout = 8'b10111011;
      13'hC94: dout = 8'b10111011;
      13'hC95: dout = 8'b10111011;
      13'hC96: dout = 8'b10111011;
      13'hC97: dout = 8'b10111011;
      13'hC98: dout = 8'b10111011;
      13'hC99: dout = 8'b10111011;
      13'hC9A: dout = 8'b10111011;
      13'hC9B: dout = 8'b10111011;
      13'hC9C: dout = 8'b10111011;
      13'hC9D: dout = 8'b10111011;
      13'hC9E: dout = 8'b10111011;
      13'hC9F: dout = 8'b10111011;
      13'hCA0: dout = 8'b10111011;
      13'hCA1: dout = 8'b10111011;
      13'hCA2: dout = 8'b10111011;
      13'hCA3: dout = 8'b10111011;
      13'hCA4: dout = 8'b10111011;
      13'hCA5: dout = 8'b10111011;
      13'hCA6: dout = 8'b10111011;
      13'hCA7: dout = 8'b10111011;
      13'hCA8: dout = 8'b10111011;
      13'hCA9: dout = 8'b10111011;
      13'hCAA: dout = 8'b10111011;
      13'hCAB: dout = 8'b10111011;
      13'hCAC: dout = 8'b10111011;
      13'hCAD: dout = 8'b10111011;
      13'hCAE: dout = 8'b10111011;
      13'hCAF: dout = 8'b10111011;
      13'hCB0: dout = 8'b10111011;
      13'hCB1: dout = 8'b10111011;
      13'hCB2: dout = 8'b10111011;
      13'hCB3: dout = 8'b10111011;
      13'hCB4: dout = 8'b10111011;
      13'hCB5: dout = 8'b10111011;
      13'hCB6: dout = 8'b10111011;
      13'hCB7: dout = 8'b10111011;
      13'hCB8: dout = 8'b10111011;
      13'hCB9: dout = 8'b10111011;
      13'hCBA: dout = 8'b10111011;
      13'hCBB: dout = 8'b10111011;
      13'hCBC: dout = 8'b10111011;
      13'hCBD: dout = 8'b10111011;
      13'hCBE: dout = 8'b10111011;
      13'hCBF: dout = 8'b10111011;
      13'hCC0: dout = 8'b10111011;
      13'hCC1: dout = 8'b10111011;
      13'hCC2: dout = 8'b10111011;
      13'hCC3: dout = 8'b10111011;
      13'hCC4: dout = 8'b10111011;
      13'hCC5: dout = 8'b10111011;
      13'hCC6: dout = 8'b10111011;
      13'hCC7: dout = 8'b10111011;
      13'hCC8: dout = 8'b10111011;
      13'hCC9: dout = 8'b10111011;
      13'hCCA: dout = 8'b10111011;
      13'hCCB: dout = 8'b10111011;
      13'hCCC: dout = 8'b10111011;
      13'hCCD: dout = 8'b10111011;
      13'hCCE: dout = 8'b10111011;
      13'hCCF: dout = 8'b10111011;
      13'hCD0: dout = 8'b10111011;
      13'hCD1: dout = 8'b10111011;
      13'hCD2: dout = 8'b10111011;
      13'hCD3: dout = 8'b10111011;
      13'hCD4: dout = 8'b10111011;
      13'hCD5: dout = 8'b10111011;
      13'hCD6: dout = 8'b10111011;
      13'hCD7: dout = 8'b10111011;
      13'hCD8: dout = 8'b10111011;
      13'hCD9: dout = 8'b10111011;
      13'hCDA: dout = 8'b10111011;
      13'hCDB: dout = 8'b10111011;
      13'hCDC: dout = 8'b10111011;
      13'hCDD: dout = 8'b10111011;
      13'hCDE: dout = 8'b10111011;
      13'hCDF: dout = 8'b10111011;
      13'hCE0: dout = 8'b10111011;
      13'hCE1: dout = 8'b10111011;
      13'hCE2: dout = 8'b10111011;
      13'hCE3: dout = 8'b10111011;
      13'hCE4: dout = 8'b10111011;
      13'hCE5: dout = 8'b10111011;
      13'hCE6: dout = 8'b10111011;
      13'hCE7: dout = 8'b10111011;
      13'hCE8: dout = 8'b10111011;
      13'hCE9: dout = 8'b10111011;
      13'hCEA: dout = 8'b10111011;
      13'hCEB: dout = 8'b10111011;
      13'hCEC: dout = 8'b10111011;
      13'hCED: dout = 8'b10111011;
      13'hCEE: dout = 8'b10111011;
      13'hCEF: dout = 8'b10111011;
      13'hCF0: dout = 8'b10111011;
      13'hCF1: dout = 8'b10111011;
      13'hCF2: dout = 8'b10111011;
      13'hCF3: dout = 8'b10111011;
      13'hCF4: dout = 8'b10111011;
      13'hCF5: dout = 8'b10111011;
      13'hCF6: dout = 8'b10111011;
      13'hCF7: dout = 8'b10111011;
      13'hCF8: dout = 8'b10111011;
      13'hCF9: dout = 8'b10111011;
      13'hCFA: dout = 8'b10111011;
      13'hCFB: dout = 8'b10111011;
      13'hCFC: dout = 8'b10111011;
      13'hCFD: dout = 8'b10111011;
      13'hCFE: dout = 8'b10111011;
      13'hCFF: dout = 8'b10111011;
      13'hD00: dout = 8'b10111011;
      13'hD01: dout = 8'b10111011;
      13'hD02: dout = 8'b10111011;
      13'hD03: dout = 8'b10111011;
      13'hD04: dout = 8'b10111011;
      13'hD05: dout = 8'b10111011;
      13'hD06: dout = 8'b10111011;
      13'hD07: dout = 8'b10111011;
      13'hD08: dout = 8'b10111011;
      13'hD09: dout = 8'b10111011;
      13'hD0A: dout = 8'b10111011;
      13'hD0B: dout = 8'b10111011;
      13'hD0C: dout = 8'b10111011;
      13'hD0D: dout = 8'b10111011;
      13'hD0E: dout = 8'b10111011;
      13'hD0F: dout = 8'b10111011;
      13'hD10: dout = 8'b10111011;
      13'hD11: dout = 8'b10111011;
      13'hD12: dout = 8'b10111011;
      13'hD13: dout = 8'b10111011;
      13'hD14: dout = 8'b10111011;
      13'hD15: dout = 8'b10111011;
      13'hD16: dout = 8'b10111011;
      13'hD17: dout = 8'b10111011;
      13'hD18: dout = 8'b10111011;
      13'hD19: dout = 8'b10111011;
      13'hD1A: dout = 8'b10111011;
      13'hD1B: dout = 8'b10111011;
      13'hD1C: dout = 8'b10111011;
      13'hD1D: dout = 8'b10111011;
      13'hD1E: dout = 8'b10111011;
      13'hD1F: dout = 8'b10111011;
      13'hD20: dout = 8'b10111011;
      13'hD21: dout = 8'b10111011;
      13'hD22: dout = 8'b10111011;
      13'hD23: dout = 8'b10111011;
      13'hD24: dout = 8'b10111011;
      13'hD25: dout = 8'b10111011;
      13'hD26: dout = 8'b10111011;
      13'hD27: dout = 8'b10111011;
      13'hD28: dout = 8'b10111011;
      13'hD29: dout = 8'b10111011;
      13'hD2A: dout = 8'b10111011;
      13'hD2B: dout = 8'b10111011;
      13'hD2C: dout = 8'b10111011;
      13'hD2D: dout = 8'b10111011;
      13'hD2E: dout = 8'b10111011;
      13'hD2F: dout = 8'b10111011;
      13'hD30: dout = 8'b10111011;
      13'hD31: dout = 8'b10111011;
      13'hD32: dout = 8'b10111011;
      13'hD33: dout = 8'b10111011;
      13'hD34: dout = 8'b10111011;
      13'hD35: dout = 8'b10111011;
      13'hD36: dout = 8'b10111011;
      13'hD37: dout = 8'b10111011;
      13'hD38: dout = 8'b10111011;
      13'hD39: dout = 8'b10111011;
      13'hD3A: dout = 8'b10111011;
      13'hD3B: dout = 8'b10111011;
      13'hD3C: dout = 8'b10111011;
      13'hD3D: dout = 8'b10111011;
      13'hD3E: dout = 8'b10111011;
      13'hD3F: dout = 8'b10111011;
      13'hD40: dout = 8'b10111011;
      13'hD41: dout = 8'b10111011;
      13'hD42: dout = 8'b10111011;
      13'hD43: dout = 8'b10111011;
      13'hD44: dout = 8'b10111011;
      13'hD45: dout = 8'b10111011;
      13'hD46: dout = 8'b10111011;
      13'hD47: dout = 8'b10111011;
      13'hD48: dout = 8'b10111011;
      13'hD49: dout = 8'b10111011;
      13'hD4A: dout = 8'b10111011;
      13'hD4B: dout = 8'b10111011;
      13'hD4C: dout = 8'b10111011;
      13'hD4D: dout = 8'b10111011;
      13'hD4E: dout = 8'b10111011;
      13'hD4F: dout = 8'b10111011;
      13'hD50: dout = 8'b10111011;
      13'hD51: dout = 8'b10111011;
      13'hD52: dout = 8'b10111011;
      13'hD53: dout = 8'b10111011;
      13'hD54: dout = 8'b10111011;
      13'hD55: dout = 8'b10111011;
      13'hD56: dout = 8'b10111011;
      13'hD57: dout = 8'b10111011;
      13'hD58: dout = 8'b10111011;
      13'hD59: dout = 8'b10111011;
      13'hD5A: dout = 8'b10111011;
      13'hD5B: dout = 8'b10111011;
      13'hD5C: dout = 8'b10111011;
      13'hD5D: dout = 8'b10111011;
      13'hD5E: dout = 8'b10111011;
      13'hD5F: dout = 8'b10111011;
      13'hD60: dout = 8'b10111011;
      13'hD61: dout = 8'b10111011;
      13'hD62: dout = 8'b10111011;
      13'hD63: dout = 8'b10111011;
      13'hD64: dout = 8'b10111011;
      13'hD65: dout = 8'b10111011;
      13'hD66: dout = 8'b10111011;
      13'hD67: dout = 8'b10111011;
      13'hD68: dout = 8'b10111011;
      13'hD69: dout = 8'b10111011;
      13'hD6A: dout = 8'b10111011;
      13'hD6B: dout = 8'b10111011;
      13'hD6C: dout = 8'b10111011;
      13'hD6D: dout = 8'b10111011;
      13'hD6E: dout = 8'b10111011;
      13'hD6F: dout = 8'b10111011;
      13'hD70: dout = 8'b10111011;
      13'hD71: dout = 8'b10111011;
      13'hD72: dout = 8'b10111011;
      13'hD73: dout = 8'b10111011;
      13'hD74: dout = 8'b10111011;
      13'hD75: dout = 8'b10111011;
      13'hD76: dout = 8'b10111011;
      13'hD77: dout = 8'b10111011;
      13'hD78: dout = 8'b10111011;
      13'hD79: dout = 8'b10111011;
      13'hD7A: dout = 8'b10111011;
      13'hD7B: dout = 8'b10111011;
      13'hD7C: dout = 8'b10111011;
      13'hD7D: dout = 8'b10111011;
      13'hD7E: dout = 8'b10111011;
      13'hD7F: dout = 8'b10111011;
      13'hD80: dout = 8'b10111011;
      13'hD81: dout = 8'b10111011;
      13'hD82: dout = 8'b10111011;
      13'hD83: dout = 8'b10111011;
      13'hD84: dout = 8'b10111011;
      13'hD85: dout = 8'b10111011;
      13'hD86: dout = 8'b10111011;
      13'hD87: dout = 8'b10111011;
      13'hD88: dout = 8'b10111011;
      13'hD89: dout = 8'b10111011;
      13'hD8A: dout = 8'b10111011;
      13'hD8B: dout = 8'b10111011;
      13'hD8C: dout = 8'b10111011;
      13'hD8D: dout = 8'b10111011;
      13'hD8E: dout = 8'b10111011;
      13'hD8F: dout = 8'b10111011;
      13'hD90: dout = 8'b10111011;
      13'hD91: dout = 8'b10111011;
      13'hD92: dout = 8'b10111011;
      13'hD93: dout = 8'b10111011;
      13'hD94: dout = 8'b10111011;
      13'hD95: dout = 8'b10111011;
      13'hD96: dout = 8'b10111011;
      13'hD97: dout = 8'b10111011;
      13'hD98: dout = 8'b10111011;
      13'hD99: dout = 8'b10111011;
      13'hD9A: dout = 8'b10111011;
      13'hD9B: dout = 8'b10111011;
      13'hD9C: dout = 8'b10111011;
      13'hD9D: dout = 8'b10111011;
      13'hD9E: dout = 8'b10111011;
      13'hD9F: dout = 8'b10111011;
      13'hDA0: dout = 8'b10111011;
      13'hDA1: dout = 8'b10111011;
      13'hDA2: dout = 8'b10111011;
      13'hDA3: dout = 8'b10111011;
      13'hDA4: dout = 8'b10111011;
      13'hDA5: dout = 8'b10111011;
      13'hDA6: dout = 8'b10111011;
      13'hDA7: dout = 8'b10111011;
      13'hDA8: dout = 8'b10111011;
      13'hDA9: dout = 8'b10111011;
      13'hDAA: dout = 8'b10111011;
      13'hDAB: dout = 8'b10111011;
      13'hDAC: dout = 8'b10111011;
      13'hDAD: dout = 8'b10111011;
      13'hDAE: dout = 8'b10111011;
      13'hDAF: dout = 8'b10111011;
      13'hDB0: dout = 8'b10111011;
      13'hDB1: dout = 8'b10111011;
      13'hDB2: dout = 8'b10111011;
      13'hDB3: dout = 8'b10111011;
      13'hDB4: dout = 8'b10111011;
      13'hDB5: dout = 8'b10111011;
      13'hDB6: dout = 8'b10111011;
      13'hDB7: dout = 8'b10111011;
      13'hDB8: dout = 8'b10111011;
      13'hDB9: dout = 8'b10111011;
      13'hDBA: dout = 8'b10111011;
      13'hDBB: dout = 8'b10111011;
      13'hDBC: dout = 8'b10111011;
      13'hDBD: dout = 8'b10111011;
      13'hDBE: dout = 8'b10111011;
      13'hDBF: dout = 8'b10111011;
      13'hDC0: dout = 8'b10111011;
      13'hDC1: dout = 8'b10111011;
      13'hDC2: dout = 8'b10111011;
      13'hDC3: dout = 8'b10111011;
      13'hDC4: dout = 8'b10111011;
      13'hDC5: dout = 8'b10111011;
      13'hDC6: dout = 8'b10111011;
      13'hDC7: dout = 8'b10111011;
      13'hDC8: dout = 8'b10111011;
      13'hDC9: dout = 8'b10111011;
      13'hDCA: dout = 8'b10111011;
      13'hDCB: dout = 8'b10111011;
      13'hDCC: dout = 8'b10111011;
      13'hDCD: dout = 8'b10111011;
      13'hDCE: dout = 8'b10111011;
      13'hDCF: dout = 8'b10111011;
      13'hDD0: dout = 8'b10111011;
      13'hDD1: dout = 8'b10111011;
      13'hDD2: dout = 8'b10111011;
      13'hDD3: dout = 8'b10111011;
      13'hDD4: dout = 8'b10111011;
      13'hDD5: dout = 8'b10111011;
      13'hDD6: dout = 8'b10111011;
      13'hDD7: dout = 8'b10111011;
      13'hDD8: dout = 8'b10111011;
      13'hDD9: dout = 8'b10111011;
      13'hDDA: dout = 8'b10111011;
      13'hDDB: dout = 8'b10111011;
      13'hDDC: dout = 8'b10111011;
      13'hDDD: dout = 8'b10111011;
      13'hDDE: dout = 8'b10111011;
      13'hDDF: dout = 8'b10111011;
      13'hDE0: dout = 8'b10111011;
      13'hDE1: dout = 8'b10111011;
      13'hDE2: dout = 8'b10111011;
      13'hDE3: dout = 8'b10111011;
      13'hDE4: dout = 8'b10111011;
      13'hDE5: dout = 8'b10111011;
      13'hDE6: dout = 8'b10111011;
      13'hDE7: dout = 8'b10111011;
      13'hDE8: dout = 8'b10111011;
      13'hDE9: dout = 8'b10111011;
      13'hDEA: dout = 8'b10111011;
      13'hDEB: dout = 8'b10111011;
      13'hDEC: dout = 8'b10111011;
      13'hDED: dout = 8'b10111011;
      13'hDEE: dout = 8'b10111011;
      13'hDEF: dout = 8'b10111011;
      13'hDF0: dout = 8'b10111011;
      13'hDF1: dout = 8'b10111011;
      13'hDF2: dout = 8'b10111011;
      13'hDF3: dout = 8'b10111011;
      13'hDF4: dout = 8'b10111011;
      13'hDF5: dout = 8'b10111011;
      13'hDF6: dout = 8'b10111011;
      13'hDF7: dout = 8'b10111011;
      13'hDF8: dout = 8'b10111011;
      13'hDF9: dout = 8'b10111011;
      13'hDFA: dout = 8'b10111011;
      13'hDFB: dout = 8'b10111011;
      13'hDFC: dout = 8'b10111011;
      13'hDFD: dout = 8'b10111011;
      13'hDFE: dout = 8'b10111011;
      13'hDFF: dout = 8'b10111011;
      13'hE00: dout = 8'b10111011;
      13'hE01: dout = 8'b10111011;
      13'hE02: dout = 8'b10111011;
      13'hE03: dout = 8'b10111011;
      13'hE04: dout = 8'b10111011;
      13'hE05: dout = 8'b10111011;
      13'hE06: dout = 8'b10111011;
      13'hE07: dout = 8'b10111011;
      13'hE08: dout = 8'b10111011;
      13'hE09: dout = 8'b10111011;
      13'hE0A: dout = 8'b10111011;
      13'hE0B: dout = 8'b10111011;
      13'hE0C: dout = 8'b10111011;
      13'hE0D: dout = 8'b10111011;
      13'hE0E: dout = 8'b10111011;
      13'hE0F: dout = 8'b10111011;
      13'hE10: dout = 8'b10111011;
      13'hE11: dout = 8'b10111011;
      13'hE12: dout = 8'b10111011;
      13'hE13: dout = 8'b10111011;
      13'hE14: dout = 8'b10111011;
      13'hE15: dout = 8'b10111011;
      13'hE16: dout = 8'b10111011;
      13'hE17: dout = 8'b10111011;
      13'hE18: dout = 8'b10111011;
      13'hE19: dout = 8'b10111011;
      13'hE1A: dout = 8'b10111011;
      13'hE1B: dout = 8'b10111011;
      13'hE1C: dout = 8'b10111011;
      13'hE1D: dout = 8'b10111011;
      13'hE1E: dout = 8'b10111011;
      13'hE1F: dout = 8'b10111011;
      13'hE20: dout = 8'b10111011;
      13'hE21: dout = 8'b10111011;
      13'hE22: dout = 8'b10111011;
      13'hE23: dout = 8'b10111011;
      13'hE24: dout = 8'b10111011;
      13'hE25: dout = 8'b10111011;
      13'hE26: dout = 8'b10111011;
      13'hE27: dout = 8'b10111011;
      13'hE28: dout = 8'b10111011;
      13'hE29: dout = 8'b10111011;
      13'hE2A: dout = 8'b10111011;
      13'hE2B: dout = 8'b10111011;
      13'hE2C: dout = 8'b10111011;
      13'hE2D: dout = 8'b10111011;
      13'hE2E: dout = 8'b10111011;
      13'hE2F: dout = 8'b10111011;
      13'hE30: dout = 8'b10111011;
      13'hE31: dout = 8'b10111011;
      13'hE32: dout = 8'b10111011;
      13'hE33: dout = 8'b10111011;
      13'hE34: dout = 8'b10111011;
      13'hE35: dout = 8'b10111011;
      13'hE36: dout = 8'b10111011;
      13'hE37: dout = 8'b10111011;
      13'hE38: dout = 8'b10111011;
      13'hE39: dout = 8'b10111011;
      13'hE3A: dout = 8'b10111011;
      13'hE3B: dout = 8'b10111011;
      13'hE3C: dout = 8'b10111011;
      13'hE3D: dout = 8'b10111011;
      13'hE3E: dout = 8'b10111011;
      13'hE3F: dout = 8'b10111011;
      13'hE40: dout = 8'b10111011;
      13'hE41: dout = 8'b10111011;
      13'hE42: dout = 8'b10111011;
      13'hE43: dout = 8'b10111011;
      13'hE44: dout = 8'b10111011;
      13'hE45: dout = 8'b10111011;
      13'hE46: dout = 8'b10111011;
      13'hE47: dout = 8'b10111011;
      13'hE48: dout = 8'b10111011;
      13'hE49: dout = 8'b10111011;
      13'hE4A: dout = 8'b10111011;
      13'hE4B: dout = 8'b10111011;
      13'hE4C: dout = 8'b10111011;
      13'hE4D: dout = 8'b10111011;
      13'hE4E: dout = 8'b10111011;
      13'hE4F: dout = 8'b10111011;
      13'hE50: dout = 8'b10111011;
      13'hE51: dout = 8'b10111011;
      13'hE52: dout = 8'b10111011;
      13'hE53: dout = 8'b10111011;
      13'hE54: dout = 8'b10111011;
      13'hE55: dout = 8'b10111011;
      13'hE56: dout = 8'b10111011;
      13'hE57: dout = 8'b10111011;
      13'hE58: dout = 8'b10111011;
      13'hE59: dout = 8'b10111011;
      13'hE5A: dout = 8'b10111011;
      13'hE5B: dout = 8'b10111011;
      13'hE5C: dout = 8'b10111011;
      13'hE5D: dout = 8'b10111011;
      13'hE5E: dout = 8'b10111011;
      13'hE5F: dout = 8'b10111011;
      13'hE60: dout = 8'b10111011;
      13'hE61: dout = 8'b10111011;
      13'hE62: dout = 8'b10111011;
      13'hE63: dout = 8'b10111011;
      13'hE64: dout = 8'b10111011;
      13'hE65: dout = 8'b10111011;
      13'hE66: dout = 8'b10111011;
      13'hE67: dout = 8'b10111011;
      13'hE68: dout = 8'b10111011;
      13'hE69: dout = 8'b10111011;
      13'hE6A: dout = 8'b10111011;
      13'hE6B: dout = 8'b10111011;
      13'hE6C: dout = 8'b10111011;
      13'hE6D: dout = 8'b10111011;
      13'hE6E: dout = 8'b10111011;
      13'hE6F: dout = 8'b10111011;
      13'hE70: dout = 8'b10111011;
      13'hE71: dout = 8'b10111011;
      13'hE72: dout = 8'b10111011;
      13'hE73: dout = 8'b10111011;
      13'hE74: dout = 8'b10111011;
      13'hE75: dout = 8'b10111011;
      13'hE76: dout = 8'b10111011;
      13'hE77: dout = 8'b10111011;
      13'hE78: dout = 8'b10111011;
      13'hE79: dout = 8'b10111011;
      13'hE7A: dout = 8'b10111011;
      13'hE7B: dout = 8'b10111011;
      13'hE7C: dout = 8'b10111011;
      13'hE7D: dout = 8'b10111011;
      13'hE7E: dout = 8'b10111011;
      13'hE7F: dout = 8'b10111011;
      13'hE80: dout = 8'b10111011;
      13'hE81: dout = 8'b10111011;
      13'hE82: dout = 8'b10111011;
      13'hE83: dout = 8'b10111011;
      13'hE84: dout = 8'b10111011;
      13'hE85: dout = 8'b10111011;
      13'hE86: dout = 8'b10111011;
      13'hE87: dout = 8'b10111011;
      13'hE88: dout = 8'b10111011;
      13'hE89: dout = 8'b10111011;
      13'hE8A: dout = 8'b10111011;
      13'hE8B: dout = 8'b10111011;
      13'hE8C: dout = 8'b10111011;
      13'hE8D: dout = 8'b10111011;
      13'hE8E: dout = 8'b10111011;
      13'hE8F: dout = 8'b10111011;
      13'hE90: dout = 8'b10111011;
      13'hE91: dout = 8'b10111011;
      13'hE92: dout = 8'b10111011;
      13'hE93: dout = 8'b10111011;
      13'hE94: dout = 8'b10111011;
      13'hE95: dout = 8'b10111011;
      13'hE96: dout = 8'b10111011;
      13'hE97: dout = 8'b10111011;
      13'hE98: dout = 8'b10111011;
      13'hE99: dout = 8'b10111011;
      13'hE9A: dout = 8'b10111011;
      13'hE9B: dout = 8'b10111011;
      13'hE9C: dout = 8'b10111011;
      13'hE9D: dout = 8'b10111011;
      13'hE9E: dout = 8'b10111011;
      13'hE9F: dout = 8'b10111011;
      13'hEA0: dout = 8'b10111011;
      13'hEA1: dout = 8'b10111011;
      13'hEA2: dout = 8'b10111011;
      13'hEA3: dout = 8'b10111011;
      13'hEA4: dout = 8'b10111011;
      13'hEA5: dout = 8'b10111011;
      13'hEA6: dout = 8'b10111011;
      13'hEA7: dout = 8'b10111011;
      13'hEA8: dout = 8'b10111011;
      13'hEA9: dout = 8'b10111011;
      13'hEAA: dout = 8'b10111011;
      13'hEAB: dout = 8'b10111011;
      13'hEAC: dout = 8'b10111011;
      13'hEAD: dout = 8'b10111011;
      13'hEAE: dout = 8'b10111011;
      13'hEAF: dout = 8'b10111011;
      13'hEB0: dout = 8'b10111011;
      13'hEB1: dout = 8'b10111011;
      13'hEB2: dout = 8'b10111011;
      13'hEB3: dout = 8'b10111011;
      13'hEB4: dout = 8'b10111011;
      13'hEB5: dout = 8'b10111011;
      13'hEB6: dout = 8'b10111011;
      13'hEB7: dout = 8'b10111011;
      13'hEB8: dout = 8'b10111011;
      13'hEB9: dout = 8'b10111011;
      13'hEBA: dout = 8'b10111011;
      13'hEBB: dout = 8'b10111011;
      13'hEBC: dout = 8'b10111011;
      13'hEBD: dout = 8'b10111011;
      13'hEBE: dout = 8'b10111011;
      13'hEBF: dout = 8'b10111011;
      13'hEC0: dout = 8'b10111011;
      13'hEC1: dout = 8'b10111011;
      13'hEC2: dout = 8'b10111011;
      13'hEC3: dout = 8'b10111011;
      13'hEC4: dout = 8'b10111011;
      13'hEC5: dout = 8'b10111011;
      13'hEC6: dout = 8'b10111011;
      13'hEC7: dout = 8'b10111011;
      13'hEC8: dout = 8'b10111011;
      13'hEC9: dout = 8'b10111011;
      13'hECA: dout = 8'b10111011;
      13'hECB: dout = 8'b10111011;
      13'hECC: dout = 8'b10111011;
      13'hECD: dout = 8'b10111011;
      13'hECE: dout = 8'b10111011;
      13'hECF: dout = 8'b10111011;
      13'hED0: dout = 8'b10111011;
      13'hED1: dout = 8'b10111011;
      13'hED2: dout = 8'b10111011;
      13'hED3: dout = 8'b10111011;
      13'hED4: dout = 8'b10111011;
      13'hED5: dout = 8'b10111011;
      13'hED6: dout = 8'b10111011;
      13'hED7: dout = 8'b10111011;
      13'hED8: dout = 8'b10111011;
      13'hED9: dout = 8'b10111011;
      13'hEDA: dout = 8'b10111011;
      13'hEDB: dout = 8'b10111011;
      13'hEDC: dout = 8'b10111011;
      13'hEDD: dout = 8'b10111011;
      13'hEDE: dout = 8'b10111011;
      13'hEDF: dout = 8'b10111011;
      13'hEE0: dout = 8'b10111011;
      13'hEE1: dout = 8'b10111011;
      13'hEE2: dout = 8'b10111011;
      13'hEE3: dout = 8'b10111011;
      13'hEE4: dout = 8'b10111011;
      13'hEE5: dout = 8'b10111011;
      13'hEE6: dout = 8'b10111011;
      13'hEE7: dout = 8'b10111011;
      13'hEE8: dout = 8'b10111011;
      13'hEE9: dout = 8'b10111011;
      13'hEEA: dout = 8'b10111011;
      13'hEEB: dout = 8'b10111011;
      13'hEEC: dout = 8'b10111011;
      13'hEED: dout = 8'b10111011;
      13'hEEE: dout = 8'b10111011;
      13'hEEF: dout = 8'b10111011;
      13'hEF0: dout = 8'b10111011;
      13'hEF1: dout = 8'b10111011;
      13'hEF2: dout = 8'b10111011;
      13'hEF3: dout = 8'b10111011;
      13'hEF4: dout = 8'b10111011;
      13'hEF5: dout = 8'b10111011;
      13'hEF6: dout = 8'b10111011;
      13'hEF7: dout = 8'b10111011;
      13'hEF8: dout = 8'b10111011;
      13'hEF9: dout = 8'b10111011;
      13'hEFA: dout = 8'b10111011;
      13'hEFB: dout = 8'b10111011;
      13'hEFC: dout = 8'b10111011;
      13'hEFD: dout = 8'b10111011;
      13'hEFE: dout = 8'b10111011;
      13'hEFF: dout = 8'b10111011;
      13'hF00: dout = 8'b10111011;
      13'hF01: dout = 8'b10111011;
      13'hF02: dout = 8'b10111011;
      13'hF03: dout = 8'b10111011;
      13'hF04: dout = 8'b10111011;
      13'hF05: dout = 8'b10111011;
      13'hF06: dout = 8'b10111011;
      13'hF07: dout = 8'b10111011;
      13'hF08: dout = 8'b10111011;
      13'hF09: dout = 8'b10111011;
      13'hF0A: dout = 8'b10111011;
      13'hF0B: dout = 8'b10111011;
      13'hF0C: dout = 8'b10111011;
      13'hF0D: dout = 8'b10111011;
      13'hF0E: dout = 8'b10111011;
      13'hF0F: dout = 8'b10111011;
      13'hF10: dout = 8'b10111011;
      13'hF11: dout = 8'b10111011;
      13'hF12: dout = 8'b10111011;
      13'hF13: dout = 8'b10111011;
      13'hF14: dout = 8'b10111011;
      13'hF15: dout = 8'b10111011;
      13'hF16: dout = 8'b10111011;
      13'hF17: dout = 8'b10111011;
      13'hF18: dout = 8'b10111011;
      13'hF19: dout = 8'b10111011;
      13'hF1A: dout = 8'b10111011;
      13'hF1B: dout = 8'b10111011;
      13'hF1C: dout = 8'b10111011;
      13'hF1D: dout = 8'b10111011;
      13'hF1E: dout = 8'b10111011;
      13'hF1F: dout = 8'b10111011;
      13'hF20: dout = 8'b10111011;
      13'hF21: dout = 8'b10111011;
      13'hF22: dout = 8'b10111011;
      13'hF23: dout = 8'b10111011;
      13'hF24: dout = 8'b10111011;
      13'hF25: dout = 8'b10111011;
      13'hF26: dout = 8'b10111011;
      13'hF27: dout = 8'b10111011;
      13'hF28: dout = 8'b10111011;
      13'hF29: dout = 8'b10111011;
      13'hF2A: dout = 8'b10111011;
      13'hF2B: dout = 8'b10111011;
      13'hF2C: dout = 8'b10111011;
      13'hF2D: dout = 8'b10111011;
      13'hF2E: dout = 8'b10111011;
      13'hF2F: dout = 8'b10111011;
      13'hF30: dout = 8'b10111011;
      13'hF31: dout = 8'b10111011;
      13'hF32: dout = 8'b10111011;
      13'hF33: dout = 8'b10111011;
      13'hF34: dout = 8'b10111011;
      13'hF35: dout = 8'b10111011;
      13'hF36: dout = 8'b10111011;
      13'hF37: dout = 8'b10111011;
      13'hF38: dout = 8'b10111011;
      13'hF39: dout = 8'b10111011;
      13'hF3A: dout = 8'b10111011;
      13'hF3B: dout = 8'b10111011;
      13'hF3C: dout = 8'b10111011;
      13'hF3D: dout = 8'b10111011;
      13'hF3E: dout = 8'b10111011;
      13'hF3F: dout = 8'b10111011;
      13'hF40: dout = 8'b10111011;
      13'hF41: dout = 8'b10111011;
      13'hF42: dout = 8'b10111011;
      13'hF43: dout = 8'b10111011;
      13'hF44: dout = 8'b10111011;
      13'hF45: dout = 8'b10111011;
      13'hF46: dout = 8'b10111011;
      13'hF47: dout = 8'b10111011;
      13'hF48: dout = 8'b10111011;
      13'hF49: dout = 8'b10111011;
      13'hF4A: dout = 8'b10111011;
      13'hF4B: dout = 8'b10111011;
      13'hF4C: dout = 8'b10111011;
      13'hF4D: dout = 8'b10111011;
      13'hF4E: dout = 8'b10111011;
      13'hF4F: dout = 8'b10111011;
      13'hF50: dout = 8'b10111011;
      13'hF51: dout = 8'b10111011;
      13'hF52: dout = 8'b10111011;
      13'hF53: dout = 8'b10111011;
      13'hF54: dout = 8'b10111011;
      13'hF55: dout = 8'b10111011;
      13'hF56: dout = 8'b10111011;
      13'hF57: dout = 8'b10111011;
      13'hF58: dout = 8'b10111011;
      13'hF59: dout = 8'b10111011;
      13'hF5A: dout = 8'b10111011;
      13'hF5B: dout = 8'b10111011;
      13'hF5C: dout = 8'b10111011;
      13'hF5D: dout = 8'b10111011;
      13'hF5E: dout = 8'b10111011;
      13'hF5F: dout = 8'b10111011;
      13'hF60: dout = 8'b10111011;
      13'hF61: dout = 8'b10111011;
      13'hF62: dout = 8'b10111011;
      13'hF63: dout = 8'b10111011;
      13'hF64: dout = 8'b10111011;
      13'hF65: dout = 8'b10111011;
      13'hF66: dout = 8'b10111011;
      13'hF67: dout = 8'b10111011;
      13'hF68: dout = 8'b10111011;
      13'hF69: dout = 8'b10111011;
      13'hF6A: dout = 8'b10111011;
      13'hF6B: dout = 8'b10111011;
      13'hF6C: dout = 8'b10111011;
      13'hF6D: dout = 8'b10111011;
      13'hF6E: dout = 8'b10111011;
      13'hF6F: dout = 8'b10111011;
      13'hF70: dout = 8'b10111011;
      13'hF71: dout = 8'b10111011;
      13'hF72: dout = 8'b10111011;
      13'hF73: dout = 8'b10111011;
      13'hF74: dout = 8'b10111011;
      13'hF75: dout = 8'b10111011;
      13'hF76: dout = 8'b10111011;
      13'hF77: dout = 8'b10111011;
      13'hF78: dout = 8'b10111011;
      13'hF79: dout = 8'b10111011;
      13'hF7A: dout = 8'b10111011;
      13'hF7B: dout = 8'b10111011;
      13'hF7C: dout = 8'b10111011;
      13'hF7D: dout = 8'b10111011;
      13'hF7E: dout = 8'b10111011;
      13'hF7F: dout = 8'b10111011;
      13'hF80: dout = 8'b10111011;
      13'hF81: dout = 8'b10111011;
      13'hF82: dout = 8'b10111011;
      13'hF83: dout = 8'b10111011;
      13'hF84: dout = 8'b10111011;
      13'hF85: dout = 8'b10111011;
      13'hF86: dout = 8'b10111011;
      13'hF87: dout = 8'b10111011;
      13'hF88: dout = 8'b10111011;
      13'hF89: dout = 8'b10111011;
      13'hF8A: dout = 8'b10111011;
      13'hF8B: dout = 8'b10111011;
      13'hF8C: dout = 8'b10111011;
      13'hF8D: dout = 8'b10111011;
      13'hF8E: dout = 8'b10111011;
      13'hF8F: dout = 8'b10111011;
      13'hF90: dout = 8'b10111011;
      13'hF91: dout = 8'b10111011;
      13'hF92: dout = 8'b10111011;
      13'hF93: dout = 8'b10111011;
      13'hF94: dout = 8'b10111011;
      13'hF95: dout = 8'b10111011;
      13'hF96: dout = 8'b10111011;
      13'hF97: dout = 8'b10111011;
      13'hF98: dout = 8'b10111011;
      13'hF99: dout = 8'b10111011;
      13'hF9A: dout = 8'b10111011;
      13'hF9B: dout = 8'b10111011;
      13'hF9C: dout = 8'b10111011;
      13'hF9D: dout = 8'b10111011;
      13'hF9E: dout = 8'b10111011;
      13'hF9F: dout = 8'b10111011;
      13'hFA0: dout = 8'b10111011;
      13'hFA1: dout = 8'b10111011;
      13'hFA2: dout = 8'b10111011;
      13'hFA3: dout = 8'b10111011;
      13'hFA4: dout = 8'b10111011;
      13'hFA5: dout = 8'b10111011;
      13'hFA6: dout = 8'b10111011;
      13'hFA7: dout = 8'b10111011;
      13'hFA8: dout = 8'b10111011;
      13'hFA9: dout = 8'b10111011;
      13'hFAA: dout = 8'b10111011;
      13'hFAB: dout = 8'b10111011;
      13'hFAC: dout = 8'b10111011;
      13'hFAD: dout = 8'b10111011;
      13'hFAE: dout = 8'b10111011;
      13'hFAF: dout = 8'b10111011;
      13'hFB0: dout = 8'b10111011;
      13'hFB1: dout = 8'b10111011;
      13'hFB2: dout = 8'b10111011;
      13'hFB3: dout = 8'b10111011;
      13'hFB4: dout = 8'b10111011;
      13'hFB5: dout = 8'b10111011;
      13'hFB6: dout = 8'b10111011;
      13'hFB7: dout = 8'b10111011;
      13'hFB8: dout = 8'b10111011;
      13'hFB9: dout = 8'b10111011;
      13'hFBA: dout = 8'b10111011;
      13'hFBB: dout = 8'b10111011;
      13'hFBC: dout = 8'b10111011;
      13'hFBD: dout = 8'b10111011;
      13'hFBE: dout = 8'b10111011;
      13'hFBF: dout = 8'b10111011;
      13'hFC0: dout = 8'b10111011;
      13'hFC1: dout = 8'b10111011;
      13'hFC2: dout = 8'b10111011;
      13'hFC3: dout = 8'b10111011;
      13'hFC4: dout = 8'b10111011;
      13'hFC5: dout = 8'b10111011;
      13'hFC6: dout = 8'b10111011;
      13'hFC7: dout = 8'b10111011;
      13'hFC8: dout = 8'b10111011;
      13'hFC9: dout = 8'b10111011;
      13'hFCA: dout = 8'b10111011;
      13'hFCB: dout = 8'b10111011;
      13'hFCC: dout = 8'b10111011;
      13'hFCD: dout = 8'b10111011;
      13'hFCE: dout = 8'b10111011;
      13'hFCF: dout = 8'b10111011;
      13'hFD0: dout = 8'b10111011;
      13'hFD1: dout = 8'b10111011;
      13'hFD2: dout = 8'b10111011;
      13'hFD3: dout = 8'b10111011;
      13'hFD4: dout = 8'b10111011;
      13'hFD5: dout = 8'b10111011;
      13'hFD6: dout = 8'b10111011;
      13'hFD7: dout = 8'b10111011;
      13'hFD8: dout = 8'b10111011;
      13'hFD9: dout = 8'b10111011;
      13'hFDA: dout = 8'b10111011;
      13'hFDB: dout = 8'b10111011;
      13'hFDC: dout = 8'b10111011;
      13'hFDD: dout = 8'b10111011;
      13'hFDE: dout = 8'b10111011;
      13'hFDF: dout = 8'b10111011;
      13'hFE0: dout = 8'b10111011;
      13'hFE1: dout = 8'b10111011;
      13'hFE2: dout = 8'b10111011;
      13'hFE3: dout = 8'b10111011;
      13'hFE4: dout = 8'b10111011;
      13'hFE5: dout = 8'b10111011;
      13'hFE6: dout = 8'b10111011;
      13'hFE7: dout = 8'b10111011;
      13'hFE8: dout = 8'b10111011;
      13'hFE9: dout = 8'b10111011;
      13'hFEA: dout = 8'b10111011;
      13'hFEB: dout = 8'b10111011;
      13'hFEC: dout = 8'b10111011;
      13'hFED: dout = 8'b10111011;
      13'hFEE: dout = 8'b10111011;
      13'hFEF: dout = 8'b10111011;
      13'hFF0: dout = 8'b10111011;
      13'hFF1: dout = 8'b10111011;
      13'hFF2: dout = 8'b10111011;
      13'hFF3: dout = 8'b10111011;
      13'hFF4: dout = 8'b10111011;
      13'hFF5: dout = 8'b10111011;
      13'hFF6: dout = 8'b10111011;
      13'hFF7: dout = 8'b10111011;
      13'hFF8: dout = 8'b10111011;
      13'hFF9: dout = 8'b10111011;
      13'hFFA: dout = 8'b10111011;
      13'hFFB: dout = 8'b10111011;
      13'hFFC: dout = 8'b10111011;
      13'hFFD: dout = 8'b10111011;
      13'hFFE: dout = 8'b10111011;
      13'hFFF: dout = 8'b10111011;
      13'h1000: dout = 8'b10111011;
      13'h1001: dout = 8'b10111011;
      13'h1002: dout = 8'b10111011;
      13'h1003: dout = 8'b10111011;
      13'h1004: dout = 8'b10111011;
      13'h1005: dout = 8'b10111011;
      13'h1006: dout = 8'b10111011;
      13'h1007: dout = 8'b10111011;
      13'h1008: dout = 8'b10111011;
      13'h1009: dout = 8'b10111011;
      13'h100A: dout = 8'b10111011;
      13'h100B: dout = 8'b10111011;
      13'h100C: dout = 8'b10111011;
      13'h100D: dout = 8'b10111011;
      13'h100E: dout = 8'b10111011;
      13'h100F: dout = 8'b10111011;
      13'h1010: dout = 8'b10111011;
      13'h1011: dout = 8'b10111011;
      13'h1012: dout = 8'b10111011;
      13'h1013: dout = 8'b10111011;
      13'h1014: dout = 8'b10111011;
      13'h1015: dout = 8'b10111011;
      13'h1016: dout = 8'b10111011;
      13'h1017: dout = 8'b10111011;
      13'h1018: dout = 8'b10111011;
      13'h1019: dout = 8'b10111011;
      13'h101A: dout = 8'b10111011;
      13'h101B: dout = 8'b10111011;
      13'h101C: dout = 8'b10111011;
      13'h101D: dout = 8'b10111011;
      13'h101E: dout = 8'b10111011;
      13'h101F: dout = 8'b10111011;
      13'h1020: dout = 8'b10111011;
      13'h1021: dout = 8'b10111011;
      13'h1022: dout = 8'b10111011;
      13'h1023: dout = 8'b10111011;
      13'h1024: dout = 8'b10111011;
      13'h1025: dout = 8'b10111011;
      13'h1026: dout = 8'b10111011;
      13'h1027: dout = 8'b10111011;
      13'h1028: dout = 8'b10111011;
      13'h1029: dout = 8'b10111011;
      13'h102A: dout = 8'b10111011;
      13'h102B: dout = 8'b10111011;
      13'h102C: dout = 8'b10111011;
      13'h102D: dout = 8'b10111011;
      13'h102E: dout = 8'b10111011;
      13'h102F: dout = 8'b10111011;
      13'h1030: dout = 8'b10111011;
      13'h1031: dout = 8'b10111011;
      13'h1032: dout = 8'b10111011;
      13'h1033: dout = 8'b10111011;
      13'h1034: dout = 8'b10111011;
      13'h1035: dout = 8'b10111011;
      13'h1036: dout = 8'b10111011;
      13'h1037: dout = 8'b10111011;
      13'h1038: dout = 8'b10111011;
      13'h1039: dout = 8'b10111011;
      13'h103A: dout = 8'b10111011;
      13'h103B: dout = 8'b10111011;
      13'h103C: dout = 8'b10111011;
      13'h103D: dout = 8'b10111011;
      13'h103E: dout = 8'b10111011;
      13'h103F: dout = 8'b10111011;
      13'h1040: dout = 8'b10111011;
      13'h1041: dout = 8'b10111011;
      13'h1042: dout = 8'b10111011;
      13'h1043: dout = 8'b10111011;
      13'h1044: dout = 8'b10111011;
      13'h1045: dout = 8'b10111011;
      13'h1046: dout = 8'b10111011;
      13'h1047: dout = 8'b10111011;
      13'h1048: dout = 8'b10111011;
      13'h1049: dout = 8'b10111011;
      13'h104A: dout = 8'b10111011;
      13'h104B: dout = 8'b10111011;
      13'h104C: dout = 8'b10111011;
      13'h104D: dout = 8'b10111011;
      13'h104E: dout = 8'b10111011;
      13'h104F: dout = 8'b10111011;
      13'h1050: dout = 8'b10111011;
      13'h1051: dout = 8'b10111011;
      13'h1052: dout = 8'b10111011;
      13'h1053: dout = 8'b10111011;
      13'h1054: dout = 8'b10111011;
      13'h1055: dout = 8'b10111011;
      13'h1056: dout = 8'b10111011;
      13'h1057: dout = 8'b10111011;
      13'h1058: dout = 8'b10111011;
      13'h1059: dout = 8'b10111011;
      13'h105A: dout = 8'b10111011;
      13'h105B: dout = 8'b10111011;
      13'h105C: dout = 8'b10111011;
      13'h105D: dout = 8'b10111011;
      13'h105E: dout = 8'b10111011;
      13'h105F: dout = 8'b10111011;
      13'h1060: dout = 8'b10111011;
      13'h1061: dout = 8'b10111011;
      13'h1062: dout = 8'b10111011;
      13'h1063: dout = 8'b10111011;
      13'h1064: dout = 8'b10111011;
      13'h1065: dout = 8'b10111011;
      13'h1066: dout = 8'b10111011;
      13'h1067: dout = 8'b10111011;
      13'h1068: dout = 8'b10111011;
      13'h1069: dout = 8'b10111011;
      13'h106A: dout = 8'b10111011;
      13'h106B: dout = 8'b10111011;
      13'h106C: dout = 8'b10111011;
      13'h106D: dout = 8'b10111011;
      13'h106E: dout = 8'b10111011;
      13'h106F: dout = 8'b10111011;
      13'h1070: dout = 8'b10111011;
      13'h1071: dout = 8'b10111011;
      13'h1072: dout = 8'b10111011;
      13'h1073: dout = 8'b10111011;
      13'h1074: dout = 8'b10111011;
      13'h1075: dout = 8'b10111011;
      13'h1076: dout = 8'b10111011;
      13'h1077: dout = 8'b10111011;
      13'h1078: dout = 8'b10111011;
      13'h1079: dout = 8'b10111011;
      13'h107A: dout = 8'b10111011;
      13'h107B: dout = 8'b10111011;
      13'h107C: dout = 8'b10111011;
      13'h107D: dout = 8'b10111011;
      13'h107E: dout = 8'b10111011;
      13'h107F: dout = 8'b10111011;
      13'h1080: dout = 8'b10111011;
      13'h1081: dout = 8'b10111011;
      13'h1082: dout = 8'b10111011;
      13'h1083: dout = 8'b10111011;
      13'h1084: dout = 8'b10111011;
      13'h1085: dout = 8'b10111011;
      13'h1086: dout = 8'b10111011;
      13'h1087: dout = 8'b10111011;
      13'h1088: dout = 8'b10111011;
      13'h1089: dout = 8'b10111011;
      13'h108A: dout = 8'b10111011;
      13'h108B: dout = 8'b10111011;
      13'h108C: dout = 8'b10111011;
      13'h108D: dout = 8'b10111011;
      13'h108E: dout = 8'b10111011;
      13'h108F: dout = 8'b10111011;
      13'h1090: dout = 8'b10111011;
      13'h1091: dout = 8'b10111011;
      13'h1092: dout = 8'b10111011;
      13'h1093: dout = 8'b10111011;
      13'h1094: dout = 8'b10111011;
      13'h1095: dout = 8'b10111011;
      13'h1096: dout = 8'b10111011;
      13'h1097: dout = 8'b10111011;
      13'h1098: dout = 8'b10111011;
      13'h1099: dout = 8'b10111011;
      13'h109A: dout = 8'b10111011;
      13'h109B: dout = 8'b10111011;
      13'h109C: dout = 8'b10111011;
      13'h109D: dout = 8'b10111011;
      13'h109E: dout = 8'b10111011;
      13'h109F: dout = 8'b10111011;
      13'h10A0: dout = 8'b10111011;
      13'h10A1: dout = 8'b10111011;
      13'h10A2: dout = 8'b10111011;
      13'h10A3: dout = 8'b10111011;
      13'h10A4: dout = 8'b10111011;
      13'h10A5: dout = 8'b10111011;
      13'h10A6: dout = 8'b10111011;
      13'h10A7: dout = 8'b10111011;
      13'h10A8: dout = 8'b10111011;
      13'h10A9: dout = 8'b10111011;
      13'h10AA: dout = 8'b10111011;
      13'h10AB: dout = 8'b10111011;
      13'h10AC: dout = 8'b10111011;
      13'h10AD: dout = 8'b10111011;
      13'h10AE: dout = 8'b10111011;
      13'h10AF: dout = 8'b10111011;
      13'h10B0: dout = 8'b10111011;
      13'h10B1: dout = 8'b10111011;
      13'h10B2: dout = 8'b10111011;
      13'h10B3: dout = 8'b10111011;
      13'h10B4: dout = 8'b10111011;
      13'h10B5: dout = 8'b10111011;
      13'h10B6: dout = 8'b10111011;
      13'h10B7: dout = 8'b10111011;
      13'h10B8: dout = 8'b10111011;
      13'h10B9: dout = 8'b10111011;
      13'h10BA: dout = 8'b10111011;
      13'h10BB: dout = 8'b10111011;
      13'h10BC: dout = 8'b10111011;
      13'h10BD: dout = 8'b10111011;
      13'h10BE: dout = 8'b10111011;
      13'h10BF: dout = 8'b10111011;
      13'h10C0: dout = 8'b10111011;
      13'h10C1: dout = 8'b10111011;
      13'h10C2: dout = 8'b10111011;
      13'h10C3: dout = 8'b10111011;
      13'h10C4: dout = 8'b10111011;
      13'h10C5: dout = 8'b10111011;
      13'h10C6: dout = 8'b10111011;
      13'h10C7: dout = 8'b10111011;
      13'h10C8: dout = 8'b10111011;
      13'h10C9: dout = 8'b10111011;
      13'h10CA: dout = 8'b10111011;
      13'h10CB: dout = 8'b10111011;
      13'h10CC: dout = 8'b10111011;
      13'h10CD: dout = 8'b10111011;
      13'h10CE: dout = 8'b10111011;
      13'h10CF: dout = 8'b10111011;
      13'h10D0: dout = 8'b10111011;
      13'h10D1: dout = 8'b10111011;
      13'h10D2: dout = 8'b10111011;
      13'h10D3: dout = 8'b10111011;
      13'h10D4: dout = 8'b10111011;
      13'h10D5: dout = 8'b10111011;
      13'h10D6: dout = 8'b10111011;
      13'h10D7: dout = 8'b10111011;
      13'h10D8: dout = 8'b10111011;
      13'h10D9: dout = 8'b10111011;
      13'h10DA: dout = 8'b10111011;
      13'h10DB: dout = 8'b10111011;
      13'h10DC: dout = 8'b10111011;
      13'h10DD: dout = 8'b10111011;
      13'h10DE: dout = 8'b10111011;
      13'h10DF: dout = 8'b10111011;
      13'h10E0: dout = 8'b10111011;
      13'h10E1: dout = 8'b10111011;
      13'h10E2: dout = 8'b10111011;
      13'h10E3: dout = 8'b10111011;
      13'h10E4: dout = 8'b10111011;
      13'h10E5: dout = 8'b10111011;
      13'h10E6: dout = 8'b10111011;
      13'h10E7: dout = 8'b10111011;
      13'h10E8: dout = 8'b10111011;
      13'h10E9: dout = 8'b10111011;
      13'h10EA: dout = 8'b10111011;
      13'h10EB: dout = 8'b10111011;
      13'h10EC: dout = 8'b10111011;
      13'h10ED: dout = 8'b10111011;
      13'h10EE: dout = 8'b10111011;
      13'h10EF: dout = 8'b10111011;
      13'h10F0: dout = 8'b10111011;
      13'h10F1: dout = 8'b10111011;
      13'h10F2: dout = 8'b10111011;
      13'h10F3: dout = 8'b10111011;
      13'h10F4: dout = 8'b10111011;
      13'h10F5: dout = 8'b10111011;
      13'h10F6: dout = 8'b10111011;
      13'h10F7: dout = 8'b10111011;
      13'h10F8: dout = 8'b10111011;
      13'h10F9: dout = 8'b10111011;
      13'h10FA: dout = 8'b10111011;
      13'h10FB: dout = 8'b10111011;
      13'h10FC: dout = 8'b10111011;
      13'h10FD: dout = 8'b10111011;
      13'h10FE: dout = 8'b10111011;
      13'h10FF: dout = 8'b10111011;
      13'h1100: dout = 8'b10111011;
      13'h1101: dout = 8'b10111011;
      13'h1102: dout = 8'b10111011;
      13'h1103: dout = 8'b10111011;
      13'h1104: dout = 8'b10111011;
      13'h1105: dout = 8'b10111011;
      13'h1106: dout = 8'b10111011;
      13'h1107: dout = 8'b10111011;
      13'h1108: dout = 8'b10111011;
      13'h1109: dout = 8'b10111011;
      13'h110A: dout = 8'b10111011;
      13'h110B: dout = 8'b10111011;
      13'h110C: dout = 8'b10111011;
      13'h110D: dout = 8'b10111011;
      13'h110E: dout = 8'b10111011;
      13'h110F: dout = 8'b10111011;
      13'h1110: dout = 8'b10111011;
      13'h1111: dout = 8'b10111011;
      13'h1112: dout = 8'b10111011;
      13'h1113: dout = 8'b10111011;
      13'h1114: dout = 8'b10111011;
      13'h1115: dout = 8'b10111011;
      13'h1116: dout = 8'b10111011;
      13'h1117: dout = 8'b10111011;
      13'h1118: dout = 8'b10111011;
      13'h1119: dout = 8'b10111011;
      13'h111A: dout = 8'b10111011;
      13'h111B: dout = 8'b10111011;
      13'h111C: dout = 8'b10111011;
      13'h111D: dout = 8'b10111011;
      13'h111E: dout = 8'b10111011;
      13'h111F: dout = 8'b10111011;
      13'h1120: dout = 8'b10111011;
      13'h1121: dout = 8'b10111011;
      13'h1122: dout = 8'b10111011;
      13'h1123: dout = 8'b10111011;
      13'h1124: dout = 8'b10111011;
      13'h1125: dout = 8'b10111011;
      13'h1126: dout = 8'b10111011;
      13'h1127: dout = 8'b10111011;
      13'h1128: dout = 8'b10111011;
      13'h1129: dout = 8'b10111011;
      13'h112A: dout = 8'b10111011;
      13'h112B: dout = 8'b10111011;
      13'h112C: dout = 8'b10111011;
      13'h112D: dout = 8'b10111011;
      13'h112E: dout = 8'b10111011;
      13'h112F: dout = 8'b10111011;
      13'h1130: dout = 8'b10111011;
      13'h1131: dout = 8'b10111011;
      13'h1132: dout = 8'b10111011;
      13'h1133: dout = 8'b10111011;
      13'h1134: dout = 8'b10111011;
      13'h1135: dout = 8'b10111011;
      13'h1136: dout = 8'b10111011;
      13'h1137: dout = 8'b10111011;
      13'h1138: dout = 8'b10111011;
      13'h1139: dout = 8'b10111011;
      13'h113A: dout = 8'b10111011;
      13'h113B: dout = 8'b10111011;
      13'h113C: dout = 8'b10111011;
      13'h113D: dout = 8'b10111011;
      13'h113E: dout = 8'b10111011;
      13'h113F: dout = 8'b10111011;
      13'h1140: dout = 8'b10111011;
      13'h1141: dout = 8'b10111011;
      13'h1142: dout = 8'b10111011;
      13'h1143: dout = 8'b10111011;
      13'h1144: dout = 8'b10111011;
      13'h1145: dout = 8'b10111011;
      13'h1146: dout = 8'b10111011;
      13'h1147: dout = 8'b10111011;
      13'h1148: dout = 8'b10111011;
      13'h1149: dout = 8'b10111011;
      13'h114A: dout = 8'b10111011;
      13'h114B: dout = 8'b10111011;
      13'h114C: dout = 8'b10111011;
      13'h114D: dout = 8'b10111011;
      13'h114E: dout = 8'b10111011;
      13'h114F: dout = 8'b10111011;
      13'h1150: dout = 8'b10111011;
      13'h1151: dout = 8'b10111011;
      13'h1152: dout = 8'b10111011;
      13'h1153: dout = 8'b10111011;
      13'h1154: dout = 8'b10111011;
      13'h1155: dout = 8'b10111011;
      13'h1156: dout = 8'b10111011;
      13'h1157: dout = 8'b10111011;
      13'h1158: dout = 8'b10111011;
      13'h1159: dout = 8'b10111011;
      13'h115A: dout = 8'b10111011;
      13'h115B: dout = 8'b10111011;
      13'h115C: dout = 8'b10111011;
      13'h115D: dout = 8'b10111011;
      13'h115E: dout = 8'b10111011;
      13'h115F: dout = 8'b10111011;
      13'h1160: dout = 8'b10111011;
      13'h1161: dout = 8'b10111011;
      13'h1162: dout = 8'b10111011;
      13'h1163: dout = 8'b10111011;
      13'h1164: dout = 8'b10111011;
      13'h1165: dout = 8'b10111011;
      13'h1166: dout = 8'b10111011;
      13'h1167: dout = 8'b10111011;
      13'h1168: dout = 8'b10111011;
      13'h1169: dout = 8'b10111011;
      13'h116A: dout = 8'b10111011;
      13'h116B: dout = 8'b10111011;
      13'h116C: dout = 8'b10111011;
      13'h116D: dout = 8'b10111011;
      13'h116E: dout = 8'b10111011;
      13'h116F: dout = 8'b10111011;
      13'h1170: dout = 8'b10111011;
      13'h1171: dout = 8'b10111011;
      13'h1172: dout = 8'b10111011;
      13'h1173: dout = 8'b10111011;
      13'h1174: dout = 8'b10111011;
      13'h1175: dout = 8'b10111011;
      13'h1176: dout = 8'b10111011;
      13'h1177: dout = 8'b10111011;
      13'h1178: dout = 8'b10111011;
      13'h1179: dout = 8'b10111011;
      13'h117A: dout = 8'b10111011;
      13'h117B: dout = 8'b10111011;
      13'h117C: dout = 8'b10111011;
      13'h117D: dout = 8'b10111011;
      13'h117E: dout = 8'b10111011;
      13'h117F: dout = 8'b10111011;
      13'h1180: dout = 8'b10111011;
      13'h1181: dout = 8'b10111011;
      13'h1182: dout = 8'b10111011;
      13'h1183: dout = 8'b10111011;
      13'h1184: dout = 8'b10111011;
      13'h1185: dout = 8'b10111011;
      13'h1186: dout = 8'b10111011;
      13'h1187: dout = 8'b10111011;
      13'h1188: dout = 8'b10111011;
      13'h1189: dout = 8'b10111011;
      13'h118A: dout = 8'b10111011;
      13'h118B: dout = 8'b10111011;
      13'h118C: dout = 8'b10111011;
      13'h118D: dout = 8'b10111011;
      13'h118E: dout = 8'b10111011;
      13'h118F: dout = 8'b10111011;
      13'h1190: dout = 8'b10111011;
      13'h1191: dout = 8'b10111011;
      13'h1192: dout = 8'b10111011;
      13'h1193: dout = 8'b10111011;
      13'h1194: dout = 8'b10111011;
      13'h1195: dout = 8'b10111011;
      13'h1196: dout = 8'b10111011;
      13'h1197: dout = 8'b10111011;
      13'h1198: dout = 8'b10111011;
      13'h1199: dout = 8'b10111011;
      13'h119A: dout = 8'b10111011;
      13'h119B: dout = 8'b10111011;
      13'h119C: dout = 8'b10111011;
      13'h119D: dout = 8'b10111011;
      13'h119E: dout = 8'b10111011;
      13'h119F: dout = 8'b10111011;
      13'h11A0: dout = 8'b10111011;
      13'h11A1: dout = 8'b10111011;
      13'h11A2: dout = 8'b10111011;
      13'h11A3: dout = 8'b10111011;
      13'h11A4: dout = 8'b10111011;
      13'h11A5: dout = 8'b10111011;
      13'h11A6: dout = 8'b10111011;
      13'h11A7: dout = 8'b10111011;
      13'h11A8: dout = 8'b10111011;
      13'h11A9: dout = 8'b10111011;
      13'h11AA: dout = 8'b10111011;
      13'h11AB: dout = 8'b10111011;
      13'h11AC: dout = 8'b10111011;
      13'h11AD: dout = 8'b10111011;
      13'h11AE: dout = 8'b10111011;
      13'h11AF: dout = 8'b10111011;
      13'h11B0: dout = 8'b10111011;
      13'h11B1: dout = 8'b10111011;
      13'h11B2: dout = 8'b10111011;
      13'h11B3: dout = 8'b10111011;
      13'h11B4: dout = 8'b10111011;
      13'h11B5: dout = 8'b10111011;
      13'h11B6: dout = 8'b10111011;
      13'h11B7: dout = 8'b10111011;
      13'h11B8: dout = 8'b10111011;
      13'h11B9: dout = 8'b10111011;
      13'h11BA: dout = 8'b10111011;
      13'h11BB: dout = 8'b10111011;
      13'h11BC: dout = 8'b10111011;
      13'h11BD: dout = 8'b10111011;
      13'h11BE: dout = 8'b10111011;
      13'h11BF: dout = 8'b10111011;
      13'h11C0: dout = 8'b10111011;
      13'h11C1: dout = 8'b10111011;
      13'h11C2: dout = 8'b10111011;
      13'h11C3: dout = 8'b10111011;
      13'h11C4: dout = 8'b10111011;
      13'h11C5: dout = 8'b10111011;
      13'h11C6: dout = 8'b10111011;
      13'h11C7: dout = 8'b10111011;
      13'h11C8: dout = 8'b10111011;
      13'h11C9: dout = 8'b10111011;
      13'h11CA: dout = 8'b10111011;
      13'h11CB: dout = 8'b10111011;
      13'h11CC: dout = 8'b10111011;
      13'h11CD: dout = 8'b10111011;
      13'h11CE: dout = 8'b10111011;
      13'h11CF: dout = 8'b10111011;
      13'h11D0: dout = 8'b10111011;
      13'h11D1: dout = 8'b10111011;
      13'h11D2: dout = 8'b10111011;
      13'h11D3: dout = 8'b10111011;
      13'h11D4: dout = 8'b10111011;
      13'h11D5: dout = 8'b10111011;
      13'h11D6: dout = 8'b10111011;
      13'h11D7: dout = 8'b10111011;
      13'h11D8: dout = 8'b10111011;
      13'h11D9: dout = 8'b10111011;
      13'h11DA: dout = 8'b10111011;
      13'h11DB: dout = 8'b10111011;
      13'h11DC: dout = 8'b10111011;
      13'h11DD: dout = 8'b10111011;
      13'h11DE: dout = 8'b10111011;
      13'h11DF: dout = 8'b10111011;
      13'h11E0: dout = 8'b10111011;
      13'h11E1: dout = 8'b10111011;
      13'h11E2: dout = 8'b10111011;
      13'h11E3: dout = 8'b10111011;
      13'h11E4: dout = 8'b10111011;
      13'h11E5: dout = 8'b10111011;
      13'h11E6: dout = 8'b10111011;
      13'h11E7: dout = 8'b10111011;
      13'h11E8: dout = 8'b10111011;
      13'h11E9: dout = 8'b10111011;
      13'h11EA: dout = 8'b10111011;
      13'h11EB: dout = 8'b10111011;
      13'h11EC: dout = 8'b10111011;
      13'h11ED: dout = 8'b10111011;
      13'h11EE: dout = 8'b10111011;
      13'h11EF: dout = 8'b10111011;
      13'h11F0: dout = 8'b10111011;
      13'h11F1: dout = 8'b10111011;
      13'h11F2: dout = 8'b10111011;
      13'h11F3: dout = 8'b10111011;
      13'h11F4: dout = 8'b10111011;
      13'h11F5: dout = 8'b10111011;
      13'h11F6: dout = 8'b10111011;
      13'h11F7: dout = 8'b10111011;
      13'h11F8: dout = 8'b10111011;
      13'h11F9: dout = 8'b10111011;
      13'h11FA: dout = 8'b10111011;
      13'h11FB: dout = 8'b10111011;
      13'h11FC: dout = 8'b10111011;
      13'h11FD: dout = 8'b10111011;
      13'h11FE: dout = 8'b10111011;
      13'h11FF: dout = 8'b10111011;
      13'h1200: dout = 8'b10111011;
      13'h1201: dout = 8'b10111011;
      13'h1202: dout = 8'b10111011;
      13'h1203: dout = 8'b10111011;
      13'h1204: dout = 8'b10111011;
      13'h1205: dout = 8'b10111011;
      13'h1206: dout = 8'b10111011;
      13'h1207: dout = 8'b10111011;
      13'h1208: dout = 8'b10111011;
      13'h1209: dout = 8'b10111011;
      13'h120A: dout = 8'b10111011;
      13'h120B: dout = 8'b10111011;
      13'h120C: dout = 8'b10111011;
      13'h120D: dout = 8'b10111011;
      13'h120E: dout = 8'b10111011;
      13'h120F: dout = 8'b10111011;
      13'h1210: dout = 8'b10111011;
      13'h1211: dout = 8'b10111011;
      13'h1212: dout = 8'b10111011;
      13'h1213: dout = 8'b10111011;
      13'h1214: dout = 8'b10111011;
      13'h1215: dout = 8'b10111011;
      13'h1216: dout = 8'b10111011;
      13'h1217: dout = 8'b10111011;
      13'h1218: dout = 8'b10111011;
      13'h1219: dout = 8'b10111011;
      13'h121A: dout = 8'b10111011;
      13'h121B: dout = 8'b10111011;
      13'h121C: dout = 8'b10111011;
      13'h121D: dout = 8'b10111011;
      13'h121E: dout = 8'b10111011;
      13'h121F: dout = 8'b10111011;
      13'h1220: dout = 8'b10111011;
      13'h1221: dout = 8'b10111011;
      13'h1222: dout = 8'b10111011;
      13'h1223: dout = 8'b10111011;
      13'h1224: dout = 8'b10111011;
      13'h1225: dout = 8'b10111011;
      13'h1226: dout = 8'b10111011;
      13'h1227: dout = 8'b10111011;
      13'h1228: dout = 8'b10111011;
      13'h1229: dout = 8'b10111011;
      13'h122A: dout = 8'b10111011;
      13'h122B: dout = 8'b10111011;
      13'h122C: dout = 8'b10111011;
      13'h122D: dout = 8'b10111011;
      13'h122E: dout = 8'b10111011;
      13'h122F: dout = 8'b10111011;
      13'h1230: dout = 8'b10111011;
      13'h1231: dout = 8'b10111011;
      13'h1232: dout = 8'b10111011;
      13'h1233: dout = 8'b10111011;
      13'h1234: dout = 8'b10111011;
      13'h1235: dout = 8'b10111011;
      13'h1236: dout = 8'b10111011;
      13'h1237: dout = 8'b10111011;
      13'h1238: dout = 8'b10111011;
      13'h1239: dout = 8'b10111011;
      13'h123A: dout = 8'b10111011;
      13'h123B: dout = 8'b10111011;
      13'h123C: dout = 8'b10111011;
      13'h123D: dout = 8'b10111011;
      13'h123E: dout = 8'b10111011;
      13'h123F: dout = 8'b10111011;
      13'h1240: dout = 8'b10111011;
      13'h1241: dout = 8'b10111011;
      13'h1242: dout = 8'b10111011;
      13'h1243: dout = 8'b10111011;
      13'h1244: dout = 8'b10111011;
      13'h1245: dout = 8'b10111011;
      13'h1246: dout = 8'b10111011;
      13'h1247: dout = 8'b10111011;
      13'h1248: dout = 8'b10111011;
      13'h1249: dout = 8'b10111011;
      13'h124A: dout = 8'b10111011;
      13'h124B: dout = 8'b10111011;
      13'h124C: dout = 8'b10111011;
      13'h124D: dout = 8'b10111011;
      13'h124E: dout = 8'b10111011;
      13'h124F: dout = 8'b10111011;
      13'h1250: dout = 8'b10111011;
      13'h1251: dout = 8'b10111011;
      13'h1252: dout = 8'b10111011;
      13'h1253: dout = 8'b10111011;
      13'h1254: dout = 8'b10111011;
      13'h1255: dout = 8'b10111011;
      13'h1256: dout = 8'b10111011;
      13'h1257: dout = 8'b10111011;
      13'h1258: dout = 8'b10111011;
      13'h1259: dout = 8'b10111011;
      13'h125A: dout = 8'b10111011;
      13'h125B: dout = 8'b10111011;
      13'h125C: dout = 8'b10111011;
      13'h125D: dout = 8'b10111011;
      13'h125E: dout = 8'b10111011;
      13'h125F: dout = 8'b10111011;
      13'h1260: dout = 8'b10111011;
      13'h1261: dout = 8'b10111011;
      13'h1262: dout = 8'b10111011;
      13'h1263: dout = 8'b10111011;
      13'h1264: dout = 8'b10111011;
      13'h1265: dout = 8'b10111011;
      13'h1266: dout = 8'b10111011;
      13'h1267: dout = 8'b10111011;
      13'h1268: dout = 8'b10111011;
      13'h1269: dout = 8'b10111011;
      13'h126A: dout = 8'b10111011;
      13'h126B: dout = 8'b10111011;
      13'h126C: dout = 8'b10111011;
      13'h126D: dout = 8'b10111011;
      13'h126E: dout = 8'b10111011;
      13'h126F: dout = 8'b10111011;
      13'h1270: dout = 8'b10111011;
      13'h1271: dout = 8'b10111011;
      13'h1272: dout = 8'b10111011;
      13'h1273: dout = 8'b10111011;
      13'h1274: dout = 8'b10111011;
      13'h1275: dout = 8'b10111011;
      13'h1276: dout = 8'b10111011;
      13'h1277: dout = 8'b10111011;
      13'h1278: dout = 8'b10111011;
      13'h1279: dout = 8'b10111011;
      13'h127A: dout = 8'b10111011;
      13'h127B: dout = 8'b10111011;
      13'h127C: dout = 8'b10111011;
      13'h127D: dout = 8'b10111011;
      13'h127E: dout = 8'b10111011;
      13'h127F: dout = 8'b10111011;
      13'h1280: dout = 8'b10111011;
      13'h1281: dout = 8'b10111011;
      13'h1282: dout = 8'b10111011;
      13'h1283: dout = 8'b10111011;
      13'h1284: dout = 8'b10111011;
      13'h1285: dout = 8'b10111011;
      13'h1286: dout = 8'b10111011;
      13'h1287: dout = 8'b10111011;
      13'h1288: dout = 8'b10111011;
      13'h1289: dout = 8'b10111011;
      13'h128A: dout = 8'b10111011;
      13'h128B: dout = 8'b10111011;
      13'h128C: dout = 8'b10111011;
      13'h128D: dout = 8'b10111011;
      13'h128E: dout = 8'b10111011;
      13'h128F: dout = 8'b10111011;
      13'h1290: dout = 8'b10111011;
      13'h1291: dout = 8'b10111011;
      13'h1292: dout = 8'b10111011;
      13'h1293: dout = 8'b10111011;
      13'h1294: dout = 8'b10111011;
      13'h1295: dout = 8'b10111011;
      13'h1296: dout = 8'b10111011;
      13'h1297: dout = 8'b10111011;
      13'h1298: dout = 8'b10111011;
      13'h1299: dout = 8'b10111011;
      13'h129A: dout = 8'b10111011;
      13'h129B: dout = 8'b10111011;
      13'h129C: dout = 8'b10111011;
      13'h129D: dout = 8'b10111011;
      13'h129E: dout = 8'b10111011;
      13'h129F: dout = 8'b10111011;
      13'h12A0: dout = 8'b10111011;
      13'h12A1: dout = 8'b10111011;
      13'h12A2: dout = 8'b10111011;
      13'h12A3: dout = 8'b10111011;
      13'h12A4: dout = 8'b10111011;
      13'h12A5: dout = 8'b10111011;
      13'h12A6: dout = 8'b10111011;
      13'h12A7: dout = 8'b10111011;
      13'h12A8: dout = 8'b10111011;
      13'h12A9: dout = 8'b10111011;
      13'h12AA: dout = 8'b10111011;
      13'h12AB: dout = 8'b10111011;
      13'h12AC: dout = 8'b10111011;
      13'h12AD: dout = 8'b10111011;
      13'h12AE: dout = 8'b10111011;
      13'h12AF: dout = 8'b10111011;
      13'h12B0: dout = 8'b10111011;
      13'h12B1: dout = 8'b10111011;
      13'h12B2: dout = 8'b10111011;
      13'h12B3: dout = 8'b10111011;
      13'h12B4: dout = 8'b10111011;
      13'h12B5: dout = 8'b10111011;
      13'h12B6: dout = 8'b10111011;
      13'h12B7: dout = 8'b10111011;
      13'h12B8: dout = 8'b10111011;
      13'h12B9: dout = 8'b10111011;
      13'h12BA: dout = 8'b10111011;
      13'h12BB: dout = 8'b10111011;
      13'h12BC: dout = 8'b10111011;
      13'h12BD: dout = 8'b10111011;
      13'h12BE: dout = 8'b10111011;
      13'h12BF: dout = 8'b10111011;
      default: dout = 8'b10111011;
    endcase
  end

endmodule
