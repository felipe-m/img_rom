//-   Background Pattern table COLOR PLANE 0
// https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
//- Autcmatically generated verilog ROM from a NES memory file----


//-  Original memory dump file name: donkeykong_ptable.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory without clock -----

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//   // clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (no clock: in the same clock cycle)




module ROM_PTABLE_DONKEYKONG_BG_PLN0
  (
     //input     clk,   // clock
     input      [11-1:0] addr,  //2048 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @*
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
          // Background pattern Table COLOR PLANE 0
      11'h0: dout  = 8'b00111000; //    0 :  56 - 0x38 -- Background 0x0
      11'h1: dout  = 8'b01001100; //    1 :  76 - 0x4c
      11'h2: dout  = 8'b11000110; //    2 : 198 - 0xc6
      11'h3: dout  = 8'b11000110; //    3 : 198 - 0xc6
      11'h4: dout  = 8'b11000110; //    4 : 198 - 0xc6
      11'h5: dout  = 8'b01100100; //    5 : 100 - 0x64
      11'h6: dout  = 8'b00111000; //    6 :  56 - 0x38
      11'h7: dout  = 8'b00000000; //    7 :   0 - 0x0
      11'h8: dout  = 8'b00011000; //    8 :  24 - 0x18 -- Background 0x1
      11'h9: dout  = 8'b00111000; //    9 :  56 - 0x38
      11'hA: dout  = 8'b00011000; //   10 :  24 - 0x18
      11'hB: dout  = 8'b00011000; //   11 :  24 - 0x18
      11'hC: dout  = 8'b00011000; //   12 :  24 - 0x18
      11'hD: dout  = 8'b00011000; //   13 :  24 - 0x18
      11'hE: dout  = 8'b01111110; //   14 : 126 - 0x7e
      11'hF: dout  = 8'b00000000; //   15 :   0 - 0x0
      11'h10: dout  = 8'b01111100; //   16 : 124 - 0x7c -- Background 0x2
      11'h11: dout  = 8'b11000110; //   17 : 198 - 0xc6
      11'h12: dout  = 8'b00001110; //   18 :  14 - 0xe
      11'h13: dout  = 8'b00111100; //   19 :  60 - 0x3c
      11'h14: dout  = 8'b01111000; //   20 : 120 - 0x78
      11'h15: dout  = 8'b11100000; //   21 : 224 - 0xe0
      11'h16: dout  = 8'b11111110; //   22 : 254 - 0xfe
      11'h17: dout  = 8'b00000000; //   23 :   0 - 0x0
      11'h18: dout  = 8'b01111110; //   24 : 126 - 0x7e -- Background 0x3
      11'h19: dout  = 8'b00001100; //   25 :  12 - 0xc
      11'h1A: dout  = 8'b00011000; //   26 :  24 - 0x18
      11'h1B: dout  = 8'b00111100; //   27 :  60 - 0x3c
      11'h1C: dout  = 8'b00000110; //   28 :   6 - 0x6
      11'h1D: dout  = 8'b11000110; //   29 : 198 - 0xc6
      11'h1E: dout  = 8'b01111100; //   30 : 124 - 0x7c
      11'h1F: dout  = 8'b00000000; //   31 :   0 - 0x0
      11'h20: dout  = 8'b00011100; //   32 :  28 - 0x1c -- Background 0x4
      11'h21: dout  = 8'b00111100; //   33 :  60 - 0x3c
      11'h22: dout  = 8'b01101100; //   34 : 108 - 0x6c
      11'h23: dout  = 8'b11001100; //   35 : 204 - 0xcc
      11'h24: dout  = 8'b11111110; //   36 : 254 - 0xfe
      11'h25: dout  = 8'b00001100; //   37 :  12 - 0xc
      11'h26: dout  = 8'b00001100; //   38 :  12 - 0xc
      11'h27: dout  = 8'b00000000; //   39 :   0 - 0x0
      11'h28: dout  = 8'b11111100; //   40 : 252 - 0xfc -- Background 0x5
      11'h29: dout  = 8'b11000000; //   41 : 192 - 0xc0
      11'h2A: dout  = 8'b11111100; //   42 : 252 - 0xfc
      11'h2B: dout  = 8'b00000110; //   43 :   6 - 0x6
      11'h2C: dout  = 8'b00000110; //   44 :   6 - 0x6
      11'h2D: dout  = 8'b11000110; //   45 : 198 - 0xc6
      11'h2E: dout  = 8'b01111100; //   46 : 124 - 0x7c
      11'h2F: dout  = 8'b00000000; //   47 :   0 - 0x0
      11'h30: dout  = 8'b00111100; //   48 :  60 - 0x3c -- Background 0x6
      11'h31: dout  = 8'b01100000; //   49 :  96 - 0x60
      11'h32: dout  = 8'b11000000; //   50 : 192 - 0xc0
      11'h33: dout  = 8'b11111100; //   51 : 252 - 0xfc
      11'h34: dout  = 8'b11000110; //   52 : 198 - 0xc6
      11'h35: dout  = 8'b11000110; //   53 : 198 - 0xc6
      11'h36: dout  = 8'b01111100; //   54 : 124 - 0x7c
      11'h37: dout  = 8'b00000000; //   55 :   0 - 0x0
      11'h38: dout  = 8'b11111110; //   56 : 254 - 0xfe -- Background 0x7
      11'h39: dout  = 8'b11000110; //   57 : 198 - 0xc6
      11'h3A: dout  = 8'b00001100; //   58 :  12 - 0xc
      11'h3B: dout  = 8'b00011000; //   59 :  24 - 0x18
      11'h3C: dout  = 8'b00110000; //   60 :  48 - 0x30
      11'h3D: dout  = 8'b00110000; //   61 :  48 - 0x30
      11'h3E: dout  = 8'b00110000; //   62 :  48 - 0x30
      11'h3F: dout  = 8'b00000000; //   63 :   0 - 0x0
      11'h40: dout  = 8'b01111000; //   64 : 120 - 0x78 -- Background 0x8
      11'h41: dout  = 8'b11000100; //   65 : 196 - 0xc4
      11'h42: dout  = 8'b11100100; //   66 : 228 - 0xe4
      11'h43: dout  = 8'b01111000; //   67 : 120 - 0x78
      11'h44: dout  = 8'b10000110; //   68 : 134 - 0x86
      11'h45: dout  = 8'b10000110; //   69 : 134 - 0x86
      11'h46: dout  = 8'b01111100; //   70 : 124 - 0x7c
      11'h47: dout  = 8'b00000000; //   71 :   0 - 0x0
      11'h48: dout  = 8'b01111100; //   72 : 124 - 0x7c -- Background 0x9
      11'h49: dout  = 8'b11000110; //   73 : 198 - 0xc6
      11'h4A: dout  = 8'b11000110; //   74 : 198 - 0xc6
      11'h4B: dout  = 8'b01111110; //   75 : 126 - 0x7e
      11'h4C: dout  = 8'b00000110; //   76 :   6 - 0x6
      11'h4D: dout  = 8'b00001100; //   77 :  12 - 0xc
      11'h4E: dout  = 8'b01111000; //   78 : 120 - 0x78
      11'h4F: dout  = 8'b00000000; //   79 :   0 - 0x0
      11'h50: dout  = 8'b00111000; //   80 :  56 - 0x38 -- Background 0xa
      11'h51: dout  = 8'b01101100; //   81 : 108 - 0x6c
      11'h52: dout  = 8'b11000110; //   82 : 198 - 0xc6
      11'h53: dout  = 8'b11000110; //   83 : 198 - 0xc6
      11'h54: dout  = 8'b11111110; //   84 : 254 - 0xfe
      11'h55: dout  = 8'b11000110; //   85 : 198 - 0xc6
      11'h56: dout  = 8'b11000110; //   86 : 198 - 0xc6
      11'h57: dout  = 8'b00000000; //   87 :   0 - 0x0
      11'h58: dout  = 8'b11111100; //   88 : 252 - 0xfc -- Background 0xb
      11'h59: dout  = 8'b11000110; //   89 : 198 - 0xc6
      11'h5A: dout  = 8'b11000110; //   90 : 198 - 0xc6
      11'h5B: dout  = 8'b11111100; //   91 : 252 - 0xfc
      11'h5C: dout  = 8'b11000110; //   92 : 198 - 0xc6
      11'h5D: dout  = 8'b11000110; //   93 : 198 - 0xc6
      11'h5E: dout  = 8'b11111100; //   94 : 252 - 0xfc
      11'h5F: dout  = 8'b00000000; //   95 :   0 - 0x0
      11'h60: dout  = 8'b00111100; //   96 :  60 - 0x3c -- Background 0xc
      11'h61: dout  = 8'b01100110; //   97 : 102 - 0x66
      11'h62: dout  = 8'b11000000; //   98 : 192 - 0xc0
      11'h63: dout  = 8'b11000000; //   99 : 192 - 0xc0
      11'h64: dout  = 8'b11000000; //  100 : 192 - 0xc0
      11'h65: dout  = 8'b01100110; //  101 : 102 - 0x66
      11'h66: dout  = 8'b00111100; //  102 :  60 - 0x3c
      11'h67: dout  = 8'b00000000; //  103 :   0 - 0x0
      11'h68: dout  = 8'b11111000; //  104 : 248 - 0xf8 -- Background 0xd
      11'h69: dout  = 8'b11001100; //  105 : 204 - 0xcc
      11'h6A: dout  = 8'b11000110; //  106 : 198 - 0xc6
      11'h6B: dout  = 8'b11000110; //  107 : 198 - 0xc6
      11'h6C: dout  = 8'b11000110; //  108 : 198 - 0xc6
      11'h6D: dout  = 8'b11001100; //  109 : 204 - 0xcc
      11'h6E: dout  = 8'b11111000; //  110 : 248 - 0xf8
      11'h6F: dout  = 8'b00000000; //  111 :   0 - 0x0
      11'h70: dout  = 8'b11111110; //  112 : 254 - 0xfe -- Background 0xe
      11'h71: dout  = 8'b11000000; //  113 : 192 - 0xc0
      11'h72: dout  = 8'b11000000; //  114 : 192 - 0xc0
      11'h73: dout  = 8'b11111100; //  115 : 252 - 0xfc
      11'h74: dout  = 8'b11000000; //  116 : 192 - 0xc0
      11'h75: dout  = 8'b11000000; //  117 : 192 - 0xc0
      11'h76: dout  = 8'b11111110; //  118 : 254 - 0xfe
      11'h77: dout  = 8'b00000000; //  119 :   0 - 0x0
      11'h78: dout  = 8'b11111110; //  120 : 254 - 0xfe -- Background 0xf
      11'h79: dout  = 8'b11000000; //  121 : 192 - 0xc0
      11'h7A: dout  = 8'b11000000; //  122 : 192 - 0xc0
      11'h7B: dout  = 8'b11111100; //  123 : 252 - 0xfc
      11'h7C: dout  = 8'b11000000; //  124 : 192 - 0xc0
      11'h7D: dout  = 8'b11000000; //  125 : 192 - 0xc0
      11'h7E: dout  = 8'b11000000; //  126 : 192 - 0xc0
      11'h7F: dout  = 8'b00000000; //  127 :   0 - 0x0
      11'h80: dout  = 8'b00111110; //  128 :  62 - 0x3e -- Background 0x10
      11'h81: dout  = 8'b01100000; //  129 :  96 - 0x60
      11'h82: dout  = 8'b11000000; //  130 : 192 - 0xc0
      11'h83: dout  = 8'b11011110; //  131 : 222 - 0xde
      11'h84: dout  = 8'b11000110; //  132 : 198 - 0xc6
      11'h85: dout  = 8'b01100110; //  133 : 102 - 0x66
      11'h86: dout  = 8'b01111110; //  134 : 126 - 0x7e
      11'h87: dout  = 8'b00000000; //  135 :   0 - 0x0
      11'h88: dout  = 8'b11000110; //  136 : 198 - 0xc6 -- Background 0x11
      11'h89: dout  = 8'b11000110; //  137 : 198 - 0xc6
      11'h8A: dout  = 8'b11000110; //  138 : 198 - 0xc6
      11'h8B: dout  = 8'b11111110; //  139 : 254 - 0xfe
      11'h8C: dout  = 8'b11000110; //  140 : 198 - 0xc6
      11'h8D: dout  = 8'b11000110; //  141 : 198 - 0xc6
      11'h8E: dout  = 8'b11000110; //  142 : 198 - 0xc6
      11'h8F: dout  = 8'b00000000; //  143 :   0 - 0x0
      11'h90: dout  = 8'b01111110; //  144 : 126 - 0x7e -- Background 0x12
      11'h91: dout  = 8'b00011000; //  145 :  24 - 0x18
      11'h92: dout  = 8'b00011000; //  146 :  24 - 0x18
      11'h93: dout  = 8'b00011000; //  147 :  24 - 0x18
      11'h94: dout  = 8'b00011000; //  148 :  24 - 0x18
      11'h95: dout  = 8'b00011000; //  149 :  24 - 0x18
      11'h96: dout  = 8'b01111110; //  150 : 126 - 0x7e
      11'h97: dout  = 8'b00000000; //  151 :   0 - 0x0
      11'h98: dout  = 8'b00011110; //  152 :  30 - 0x1e -- Background 0x13
      11'h99: dout  = 8'b00000110; //  153 :   6 - 0x6
      11'h9A: dout  = 8'b00000110; //  154 :   6 - 0x6
      11'h9B: dout  = 8'b00000110; //  155 :   6 - 0x6
      11'h9C: dout  = 8'b11000110; //  156 : 198 - 0xc6
      11'h9D: dout  = 8'b11000110; //  157 : 198 - 0xc6
      11'h9E: dout  = 8'b01111100; //  158 : 124 - 0x7c
      11'h9F: dout  = 8'b00000000; //  159 :   0 - 0x0
      11'hA0: dout  = 8'b11000110; //  160 : 198 - 0xc6 -- Background 0x14
      11'hA1: dout  = 8'b11001100; //  161 : 204 - 0xcc
      11'hA2: dout  = 8'b11011000; //  162 : 216 - 0xd8
      11'hA3: dout  = 8'b11110000; //  163 : 240 - 0xf0
      11'hA4: dout  = 8'b11111000; //  164 : 248 - 0xf8
      11'hA5: dout  = 8'b11011100; //  165 : 220 - 0xdc
      11'hA6: dout  = 8'b11001110; //  166 : 206 - 0xce
      11'hA7: dout  = 8'b00000000; //  167 :   0 - 0x0
      11'hA8: dout  = 8'b01100000; //  168 :  96 - 0x60 -- Background 0x15
      11'hA9: dout  = 8'b01100000; //  169 :  96 - 0x60
      11'hAA: dout  = 8'b01100000; //  170 :  96 - 0x60
      11'hAB: dout  = 8'b01100000; //  171 :  96 - 0x60
      11'hAC: dout  = 8'b01100000; //  172 :  96 - 0x60
      11'hAD: dout  = 8'b01100000; //  173 :  96 - 0x60
      11'hAE: dout  = 8'b01111110; //  174 : 126 - 0x7e
      11'hAF: dout  = 8'b00000000; //  175 :   0 - 0x0
      11'hB0: dout  = 8'b11000110; //  176 : 198 - 0xc6 -- Background 0x16
      11'hB1: dout  = 8'b11101110; //  177 : 238 - 0xee
      11'hB2: dout  = 8'b11111110; //  178 : 254 - 0xfe
      11'hB3: dout  = 8'b11111110; //  179 : 254 - 0xfe
      11'hB4: dout  = 8'b11010110; //  180 : 214 - 0xd6
      11'hB5: dout  = 8'b11000110; //  181 : 198 - 0xc6
      11'hB6: dout  = 8'b11000110; //  182 : 198 - 0xc6
      11'hB7: dout  = 8'b00000000; //  183 :   0 - 0x0
      11'hB8: dout  = 8'b11000110; //  184 : 198 - 0xc6 -- Background 0x17
      11'hB9: dout  = 8'b11100110; //  185 : 230 - 0xe6
      11'hBA: dout  = 8'b11110110; //  186 : 246 - 0xf6
      11'hBB: dout  = 8'b11111110; //  187 : 254 - 0xfe
      11'hBC: dout  = 8'b11011110; //  188 : 222 - 0xde
      11'hBD: dout  = 8'b11001110; //  189 : 206 - 0xce
      11'hBE: dout  = 8'b11000110; //  190 : 198 - 0xc6
      11'hBF: dout  = 8'b00000000; //  191 :   0 - 0x0
      11'hC0: dout  = 8'b01111100; //  192 : 124 - 0x7c -- Background 0x18
      11'hC1: dout  = 8'b11000110; //  193 : 198 - 0xc6
      11'hC2: dout  = 8'b11000110; //  194 : 198 - 0xc6
      11'hC3: dout  = 8'b11000110; //  195 : 198 - 0xc6
      11'hC4: dout  = 8'b11000110; //  196 : 198 - 0xc6
      11'hC5: dout  = 8'b11000110; //  197 : 198 - 0xc6
      11'hC6: dout  = 8'b01111100; //  198 : 124 - 0x7c
      11'hC7: dout  = 8'b00000000; //  199 :   0 - 0x0
      11'hC8: dout  = 8'b11111100; //  200 : 252 - 0xfc -- Background 0x19
      11'hC9: dout  = 8'b11000110; //  201 : 198 - 0xc6
      11'hCA: dout  = 8'b11000110; //  202 : 198 - 0xc6
      11'hCB: dout  = 8'b11000110; //  203 : 198 - 0xc6
      11'hCC: dout  = 8'b11111100; //  204 : 252 - 0xfc
      11'hCD: dout  = 8'b11000000; //  205 : 192 - 0xc0
      11'hCE: dout  = 8'b11000000; //  206 : 192 - 0xc0
      11'hCF: dout  = 8'b00000000; //  207 :   0 - 0x0
      11'hD0: dout  = 8'b01111100; //  208 : 124 - 0x7c -- Background 0x1a
      11'hD1: dout  = 8'b11000110; //  209 : 198 - 0xc6
      11'hD2: dout  = 8'b11000110; //  210 : 198 - 0xc6
      11'hD3: dout  = 8'b11000110; //  211 : 198 - 0xc6
      11'hD4: dout  = 8'b11011110; //  212 : 222 - 0xde
      11'hD5: dout  = 8'b11001100; //  213 : 204 - 0xcc
      11'hD6: dout  = 8'b01111010; //  214 : 122 - 0x7a
      11'hD7: dout  = 8'b00000000; //  215 :   0 - 0x0
      11'hD8: dout  = 8'b11111100; //  216 : 252 - 0xfc -- Background 0x1b
      11'hD9: dout  = 8'b11000110; //  217 : 198 - 0xc6
      11'hDA: dout  = 8'b11000110; //  218 : 198 - 0xc6
      11'hDB: dout  = 8'b11001110; //  219 : 206 - 0xce
      11'hDC: dout  = 8'b11111000; //  220 : 248 - 0xf8
      11'hDD: dout  = 8'b11011100; //  221 : 220 - 0xdc
      11'hDE: dout  = 8'b11001110; //  222 : 206 - 0xce
      11'hDF: dout  = 8'b00000000; //  223 :   0 - 0x0
      11'hE0: dout  = 8'b01111000; //  224 : 120 - 0x78 -- Background 0x1c
      11'hE1: dout  = 8'b11001100; //  225 : 204 - 0xcc
      11'hE2: dout  = 8'b11000000; //  226 : 192 - 0xc0
      11'hE3: dout  = 8'b01111100; //  227 : 124 - 0x7c
      11'hE4: dout  = 8'b00000110; //  228 :   6 - 0x6
      11'hE5: dout  = 8'b11000110; //  229 : 198 - 0xc6
      11'hE6: dout  = 8'b01111100; //  230 : 124 - 0x7c
      11'hE7: dout  = 8'b00000000; //  231 :   0 - 0x0
      11'hE8: dout  = 8'b01111110; //  232 : 126 - 0x7e -- Background 0x1d
      11'hE9: dout  = 8'b00011000; //  233 :  24 - 0x18
      11'hEA: dout  = 8'b00011000; //  234 :  24 - 0x18
      11'hEB: dout  = 8'b00011000; //  235 :  24 - 0x18
      11'hEC: dout  = 8'b00011000; //  236 :  24 - 0x18
      11'hED: dout  = 8'b00011000; //  237 :  24 - 0x18
      11'hEE: dout  = 8'b00011000; //  238 :  24 - 0x18
      11'hEF: dout  = 8'b00000000; //  239 :   0 - 0x0
      11'hF0: dout  = 8'b11000110; //  240 : 198 - 0xc6 -- Background 0x1e
      11'hF1: dout  = 8'b11000110; //  241 : 198 - 0xc6
      11'hF2: dout  = 8'b11000110; //  242 : 198 - 0xc6
      11'hF3: dout  = 8'b11000110; //  243 : 198 - 0xc6
      11'hF4: dout  = 8'b11000110; //  244 : 198 - 0xc6
      11'hF5: dout  = 8'b11000110; //  245 : 198 - 0xc6
      11'hF6: dout  = 8'b01111100; //  246 : 124 - 0x7c
      11'hF7: dout  = 8'b00000000; //  247 :   0 - 0x0
      11'hF8: dout  = 8'b11000110; //  248 : 198 - 0xc6 -- Background 0x1f
      11'hF9: dout  = 8'b11000110; //  249 : 198 - 0xc6
      11'hFA: dout  = 8'b11000110; //  250 : 198 - 0xc6
      11'hFB: dout  = 8'b11101110; //  251 : 238 - 0xee
      11'hFC: dout  = 8'b01111100; //  252 : 124 - 0x7c
      11'hFD: dout  = 8'b00111000; //  253 :  56 - 0x38
      11'hFE: dout  = 8'b00010000; //  254 :  16 - 0x10
      11'hFF: dout  = 8'b00000000; //  255 :   0 - 0x0
      11'h100: dout  = 8'b11000110; //  256 : 198 - 0xc6 -- Background 0x20
      11'h101: dout  = 8'b11000110; //  257 : 198 - 0xc6
      11'h102: dout  = 8'b11010110; //  258 : 214 - 0xd6
      11'h103: dout  = 8'b11111110; //  259 : 254 - 0xfe
      11'h104: dout  = 8'b11111110; //  260 : 254 - 0xfe
      11'h105: dout  = 8'b11101110; //  261 : 238 - 0xee
      11'h106: dout  = 8'b11000110; //  262 : 198 - 0xc6
      11'h107: dout  = 8'b00000000; //  263 :   0 - 0x0
      11'h108: dout  = 8'b11000110; //  264 : 198 - 0xc6 -- Background 0x21
      11'h109: dout  = 8'b11101110; //  265 : 238 - 0xee
      11'h10A: dout  = 8'b01111100; //  266 : 124 - 0x7c
      11'h10B: dout  = 8'b00111000; //  267 :  56 - 0x38
      11'h10C: dout  = 8'b01111100; //  268 : 124 - 0x7c
      11'h10D: dout  = 8'b11101110; //  269 : 238 - 0xee
      11'h10E: dout  = 8'b11000110; //  270 : 198 - 0xc6
      11'h10F: dout  = 8'b00000000; //  271 :   0 - 0x0
      11'h110: dout  = 8'b01100110; //  272 : 102 - 0x66 -- Background 0x22
      11'h111: dout  = 8'b01100110; //  273 : 102 - 0x66
      11'h112: dout  = 8'b01100110; //  274 : 102 - 0x66
      11'h113: dout  = 8'b00111100; //  275 :  60 - 0x3c
      11'h114: dout  = 8'b00011000; //  276 :  24 - 0x18
      11'h115: dout  = 8'b00011000; //  277 :  24 - 0x18
      11'h116: dout  = 8'b00011000; //  278 :  24 - 0x18
      11'h117: dout  = 8'b00000000; //  279 :   0 - 0x0
      11'h118: dout  = 8'b11111110; //  280 : 254 - 0xfe -- Background 0x23
      11'h119: dout  = 8'b00001110; //  281 :  14 - 0xe
      11'h11A: dout  = 8'b00011100; //  282 :  28 - 0x1c
      11'h11B: dout  = 8'b00111000; //  283 :  56 - 0x38
      11'h11C: dout  = 8'b01110000; //  284 : 112 - 0x70
      11'h11D: dout  = 8'b11100000; //  285 : 224 - 0xe0
      11'h11E: dout  = 8'b11111110; //  286 : 254 - 0xfe
      11'h11F: dout  = 8'b00000000; //  287 :   0 - 0x0
      11'h120: dout  = 8'b00000000; //  288 :   0 - 0x0 -- Background 0x24
      11'h121: dout  = 8'b00000000; //  289 :   0 - 0x0
      11'h122: dout  = 8'b00000000; //  290 :   0 - 0x0
      11'h123: dout  = 8'b00000000; //  291 :   0 - 0x0
      11'h124: dout  = 8'b00000000; //  292 :   0 - 0x0
      11'h125: dout  = 8'b00000000; //  293 :   0 - 0x0
      11'h126: dout  = 8'b00000000; //  294 :   0 - 0x0
      11'h127: dout  = 8'b00000000; //  295 :   0 - 0x0
      11'h128: dout  = 8'b00000000; //  296 :   0 - 0x0 -- Background 0x25
      11'h129: dout  = 8'b00000000; //  297 :   0 - 0x0
      11'h12A: dout  = 8'b00000110; //  298 :   6 - 0x6
      11'h12B: dout  = 8'b00001110; //  299 :  14 - 0xe
      11'h12C: dout  = 8'b00001000; //  300 :   8 - 0x8
      11'h12D: dout  = 8'b00001000; //  301 :   8 - 0x8
      11'h12E: dout  = 8'b00001000; //  302 :   8 - 0x8
      11'h12F: dout  = 8'b00001000; //  303 :   8 - 0x8
      11'h130: dout  = 8'b00000000; //  304 :   0 - 0x0 -- Background 0x26
      11'h131: dout  = 8'b01111000; //  305 : 120 - 0x78
      11'h132: dout  = 8'b01100101; //  306 : 101 - 0x65
      11'h133: dout  = 8'b01111001; //  307 : 121 - 0x79
      11'h134: dout  = 8'b01100101; //  308 : 101 - 0x65
      11'h135: dout  = 8'b01100101; //  309 : 101 - 0x65
      11'h136: dout  = 8'b01111000; //  310 : 120 - 0x78
      11'h137: dout  = 8'b00000000; //  311 :   0 - 0x0
      11'h138: dout  = 8'b00000000; //  312 :   0 - 0x0 -- Background 0x27
      11'h139: dout  = 8'b11100100; //  313 : 228 - 0xe4
      11'h13A: dout  = 8'b10010110; //  314 : 150 - 0x96
      11'h13B: dout  = 8'b10010110; //  315 : 150 - 0x96
      11'h13C: dout  = 8'b10010111; //  316 : 151 - 0x97
      11'h13D: dout  = 8'b10010110; //  317 : 150 - 0x96
      11'h13E: dout  = 8'b11100110; //  318 : 230 - 0xe6
      11'h13F: dout  = 8'b00000000; //  319 :   0 - 0x0
      11'h140: dout  = 8'b00000000; //  320 :   0 - 0x0 -- Background 0x28
      11'h141: dout  = 8'b01011001; //  321 :  89 - 0x59
      11'h142: dout  = 8'b01011001; //  322 :  89 - 0x59
      11'h143: dout  = 8'b01011001; //  323 :  89 - 0x59
      11'h144: dout  = 8'b01011001; //  324 :  89 - 0x59
      11'h145: dout  = 8'b11011001; //  325 : 217 - 0xd9
      11'h146: dout  = 8'b01001110; //  326 :  78 - 0x4e
      11'h147: dout  = 8'b00000000; //  327 :   0 - 0x0
      11'h148: dout  = 8'b00000000; //  328 :   0 - 0x0 -- Background 0x29
      11'h149: dout  = 8'b00111100; //  329 :  60 - 0x3c
      11'h14A: dout  = 8'b01110000; //  330 : 112 - 0x70
      11'h14B: dout  = 8'b01110000; //  331 : 112 - 0x70
      11'h14C: dout  = 8'b00111100; //  332 :  60 - 0x3c
      11'h14D: dout  = 8'b00001100; //  333 :  12 - 0xc
      11'h14E: dout  = 8'b01111000; //  334 : 120 - 0x78
      11'h14F: dout  = 8'b00000000; //  335 :   0 - 0x0
      11'h150: dout  = 8'b00000000; //  336 :   0 - 0x0 -- Background 0x2a
      11'h151: dout  = 8'b00000000; //  337 :   0 - 0x0
      11'h152: dout  = 8'b11000110; //  338 : 198 - 0xc6
      11'h153: dout  = 8'b11101110; //  339 : 238 - 0xee
      11'h154: dout  = 8'b00101000; //  340 :  40 - 0x28
      11'h155: dout  = 8'b00101000; //  341 :  40 - 0x28
      11'h156: dout  = 8'b00101000; //  342 :  40 - 0x28
      11'h157: dout  = 8'b00101000; //  343 :  40 - 0x28
      11'h158: dout  = 8'b00001000; //  344 :   8 - 0x8 -- Background 0x2b
      11'h159: dout  = 8'b00001000; //  345 :   8 - 0x8
      11'h15A: dout  = 8'b00001000; //  346 :   8 - 0x8
      11'h15B: dout  = 8'b00001000; //  347 :   8 - 0x8
      11'h15C: dout  = 8'b00001110; //  348 :  14 - 0xe
      11'h15D: dout  = 8'b00000110; //  349 :   6 - 0x6
      11'h15E: dout  = 8'b00000000; //  350 :   0 - 0x0
      11'h15F: dout  = 8'b00000000; //  351 :   0 - 0x0
      11'h160: dout  = 8'b00101000; //  352 :  40 - 0x28 -- Background 0x2c
      11'h161: dout  = 8'b00101000; //  353 :  40 - 0x28
      11'h162: dout  = 8'b00101000; //  354 :  40 - 0x28
      11'h163: dout  = 8'b00101000; //  355 :  40 - 0x28
      11'h164: dout  = 8'b11101110; //  356 : 238 - 0xee
      11'h165: dout  = 8'b11000110; //  357 : 198 - 0xc6
      11'h166: dout  = 8'b00000000; //  358 :   0 - 0x0
      11'h167: dout  = 8'b00000000; //  359 :   0 - 0x0
      11'h168: dout  = 8'b00000000; //  360 :   0 - 0x0 -- Background 0x2d
      11'h169: dout  = 8'b00000000; //  361 :   0 - 0x0
      11'h16A: dout  = 8'b01100000; //  362 :  96 - 0x60
      11'h16B: dout  = 8'b01110000; //  363 : 112 - 0x70
      11'h16C: dout  = 8'b00010000; //  364 :  16 - 0x10
      11'h16D: dout  = 8'b00010000; //  365 :  16 - 0x10
      11'h16E: dout  = 8'b00010000; //  366 :  16 - 0x10
      11'h16F: dout  = 8'b00010000; //  367 :  16 - 0x10
      11'h170: dout  = 8'b00011100; //  368 :  28 - 0x1c -- Background 0x2e
      11'h171: dout  = 8'b00111110; //  369 :  62 - 0x3e
      11'h172: dout  = 8'b00111100; //  370 :  60 - 0x3c
      11'h173: dout  = 8'b00111000; //  371 :  56 - 0x38
      11'h174: dout  = 8'b00110000; //  372 :  48 - 0x30
      11'h175: dout  = 8'b00000000; //  373 :   0 - 0x0
      11'h176: dout  = 8'b01100000; //  374 :  96 - 0x60
      11'h177: dout  = 8'b00000000; //  375 :   0 - 0x0
      11'h178: dout  = 8'b00010000; //  376 :  16 - 0x10 -- Background 0x2f
      11'h179: dout  = 8'b00010000; //  377 :  16 - 0x10
      11'h17A: dout  = 8'b00010000; //  378 :  16 - 0x10
      11'h17B: dout  = 8'b00010000; //  379 :  16 - 0x10
      11'h17C: dout  = 8'b01110000; //  380 : 112 - 0x70
      11'h17D: dout  = 8'b01100000; //  381 :  96 - 0x60
      11'h17E: dout  = 8'b00000000; //  382 :   0 - 0x0
      11'h17F: dout  = 8'b00000000; //  383 :   0 - 0x0
      11'h180: dout  = 8'b11111111; //  384 : 255 - 0xff -- Background 0x30
      11'h181: dout  = 8'b11111111; //  385 : 255 - 0xff
      11'h182: dout  = 8'b00111000; //  386 :  56 - 0x38
      11'h183: dout  = 8'b01101100; //  387 : 108 - 0x6c
      11'h184: dout  = 8'b11000110; //  388 : 198 - 0xc6
      11'h185: dout  = 8'b10000011; //  389 : 131 - 0x83
      11'h186: dout  = 8'b11111111; //  390 : 255 - 0xff
      11'h187: dout  = 8'b11111111; //  391 : 255 - 0xff
      11'h188: dout  = 8'b11111111; //  392 : 255 - 0xff -- Background 0x31
      11'h189: dout  = 8'b00111000; //  393 :  56 - 0x38
      11'h18A: dout  = 8'b01101100; //  394 : 108 - 0x6c
      11'h18B: dout  = 8'b11000110; //  395 : 198 - 0xc6
      11'h18C: dout  = 8'b10000011; //  396 : 131 - 0x83
      11'h18D: dout  = 8'b11111111; //  397 : 255 - 0xff
      11'h18E: dout  = 8'b11111111; //  398 : 255 - 0xff
      11'h18F: dout  = 8'b00000000; //  399 :   0 - 0x0
      11'h190: dout  = 8'b00111000; //  400 :  56 - 0x38 -- Background 0x32
      11'h191: dout  = 8'b01101100; //  401 : 108 - 0x6c
      11'h192: dout  = 8'b11000110; //  402 : 198 - 0xc6
      11'h193: dout  = 8'b10000011; //  403 : 131 - 0x83
      11'h194: dout  = 8'b11111111; //  404 : 255 - 0xff
      11'h195: dout  = 8'b11111111; //  405 : 255 - 0xff
      11'h196: dout  = 8'b00000000; //  406 :   0 - 0x0
      11'h197: dout  = 8'b00000000; //  407 :   0 - 0x0
      11'h198: dout  = 8'b01101100; //  408 : 108 - 0x6c -- Background 0x33
      11'h199: dout  = 8'b11000110; //  409 : 198 - 0xc6
      11'h19A: dout  = 8'b10000011; //  410 : 131 - 0x83
      11'h19B: dout  = 8'b11111111; //  411 : 255 - 0xff
      11'h19C: dout  = 8'b11111111; //  412 : 255 - 0xff
      11'h19D: dout  = 8'b00000000; //  413 :   0 - 0x0
      11'h19E: dout  = 8'b00000000; //  414 :   0 - 0x0
      11'h19F: dout  = 8'b00000000; //  415 :   0 - 0x0
      11'h1A0: dout  = 8'b11000110; //  416 : 198 - 0xc6 -- Background 0x34
      11'h1A1: dout  = 8'b10000011; //  417 : 131 - 0x83
      11'h1A2: dout  = 8'b11111111; //  418 : 255 - 0xff
      11'h1A3: dout  = 8'b11111111; //  419 : 255 - 0xff
      11'h1A4: dout  = 8'b00000000; //  420 :   0 - 0x0
      11'h1A5: dout  = 8'b00000000; //  421 :   0 - 0x0
      11'h1A6: dout  = 8'b00000000; //  422 :   0 - 0x0
      11'h1A7: dout  = 8'b00000000; //  423 :   0 - 0x0
      11'h1A8: dout  = 8'b10000011; //  424 : 131 - 0x83 -- Background 0x35
      11'h1A9: dout  = 8'b11111111; //  425 : 255 - 0xff
      11'h1AA: dout  = 8'b11111111; //  426 : 255 - 0xff
      11'h1AB: dout  = 8'b00000000; //  427 :   0 - 0x0
      11'h1AC: dout  = 8'b00000000; //  428 :   0 - 0x0
      11'h1AD: dout  = 8'b00000000; //  429 :   0 - 0x0
      11'h1AE: dout  = 8'b00000000; //  430 :   0 - 0x0
      11'h1AF: dout  = 8'b00000000; //  431 :   0 - 0x0
      11'h1B0: dout  = 8'b11111111; //  432 : 255 - 0xff -- Background 0x36
      11'h1B1: dout  = 8'b11111111; //  433 : 255 - 0xff
      11'h1B2: dout  = 8'b00000000; //  434 :   0 - 0x0
      11'h1B3: dout  = 8'b00000000; //  435 :   0 - 0x0
      11'h1B4: dout  = 8'b00000000; //  436 :   0 - 0x0
      11'h1B5: dout  = 8'b00000000; //  437 :   0 - 0x0
      11'h1B6: dout  = 8'b00000000; //  438 :   0 - 0x0
      11'h1B7: dout  = 8'b00000000; //  439 :   0 - 0x0
      11'h1B8: dout  = 8'b11111111; //  440 : 255 - 0xff -- Background 0x37
      11'h1B9: dout  = 8'b00000000; //  441 :   0 - 0x0
      11'h1BA: dout  = 8'b00000000; //  442 :   0 - 0x0
      11'h1BB: dout  = 8'b00000000; //  443 :   0 - 0x0
      11'h1BC: dout  = 8'b00000000; //  444 :   0 - 0x0
      11'h1BD: dout  = 8'b00000000; //  445 :   0 - 0x0
      11'h1BE: dout  = 8'b00000000; //  446 :   0 - 0x0
      11'h1BF: dout  = 8'b00000000; //  447 :   0 - 0x0
      11'h1C0: dout  = 8'b00000000; //  448 :   0 - 0x0 -- Background 0x38
      11'h1C1: dout  = 8'b00000000; //  449 :   0 - 0x0
      11'h1C2: dout  = 8'b00000000; //  450 :   0 - 0x0
      11'h1C3: dout  = 8'b00000000; //  451 :   0 - 0x0
      11'h1C4: dout  = 8'b00000000; //  452 :   0 - 0x0
      11'h1C5: dout  = 8'b00000000; //  453 :   0 - 0x0
      11'h1C6: dout  = 8'b00000000; //  454 :   0 - 0x0
      11'h1C7: dout  = 8'b11111111; //  455 : 255 - 0xff
      11'h1C8: dout  = 8'b00000000; //  456 :   0 - 0x0 -- Background 0x39
      11'h1C9: dout  = 8'b00000000; //  457 :   0 - 0x0
      11'h1CA: dout  = 8'b00000000; //  458 :   0 - 0x0
      11'h1CB: dout  = 8'b00000000; //  459 :   0 - 0x0
      11'h1CC: dout  = 8'b00000000; //  460 :   0 - 0x0
      11'h1CD: dout  = 8'b00000000; //  461 :   0 - 0x0
      11'h1CE: dout  = 8'b11111111; //  462 : 255 - 0xff
      11'h1CF: dout  = 8'b11111111; //  463 : 255 - 0xff
      11'h1D0: dout  = 8'b00000000; //  464 :   0 - 0x0 -- Background 0x3a
      11'h1D1: dout  = 8'b00000000; //  465 :   0 - 0x0
      11'h1D2: dout  = 8'b00000000; //  466 :   0 - 0x0
      11'h1D3: dout  = 8'b00000000; //  467 :   0 - 0x0
      11'h1D4: dout  = 8'b00000000; //  468 :   0 - 0x0
      11'h1D5: dout  = 8'b11111111; //  469 : 255 - 0xff
      11'h1D6: dout  = 8'b11111111; //  470 : 255 - 0xff
      11'h1D7: dout  = 8'b00111000; //  471 :  56 - 0x38
      11'h1D8: dout  = 8'b00000000; //  472 :   0 - 0x0 -- Background 0x3b
      11'h1D9: dout  = 8'b00000000; //  473 :   0 - 0x0
      11'h1DA: dout  = 8'b00000000; //  474 :   0 - 0x0
      11'h1DB: dout  = 8'b00000000; //  475 :   0 - 0x0
      11'h1DC: dout  = 8'b11111111; //  476 : 255 - 0xff
      11'h1DD: dout  = 8'b11111111; //  477 : 255 - 0xff
      11'h1DE: dout  = 8'b00111000; //  478 :  56 - 0x38
      11'h1DF: dout  = 8'b01101100; //  479 : 108 - 0x6c
      11'h1E0: dout  = 8'b00000000; //  480 :   0 - 0x0 -- Background 0x3c
      11'h1E1: dout  = 8'b00000000; //  481 :   0 - 0x0
      11'h1E2: dout  = 8'b00000000; //  482 :   0 - 0x0
      11'h1E3: dout  = 8'b11111111; //  483 : 255 - 0xff
      11'h1E4: dout  = 8'b11111111; //  484 : 255 - 0xff
      11'h1E5: dout  = 8'b00111000; //  485 :  56 - 0x38
      11'h1E6: dout  = 8'b01101100; //  486 : 108 - 0x6c
      11'h1E7: dout  = 8'b11000110; //  487 : 198 - 0xc6
      11'h1E8: dout  = 8'b00000000; //  488 :   0 - 0x0 -- Background 0x3d
      11'h1E9: dout  = 8'b00000000; //  489 :   0 - 0x0
      11'h1EA: dout  = 8'b11111111; //  490 : 255 - 0xff
      11'h1EB: dout  = 8'b11111111; //  491 : 255 - 0xff
      11'h1EC: dout  = 8'b00111000; //  492 :  56 - 0x38
      11'h1ED: dout  = 8'b01101100; //  493 : 108 - 0x6c
      11'h1EE: dout  = 8'b11000110; //  494 : 198 - 0xc6
      11'h1EF: dout  = 8'b10000011; //  495 : 131 - 0x83
      11'h1F0: dout  = 8'b00000000; //  496 :   0 - 0x0 -- Background 0x3e
      11'h1F1: dout  = 8'b11111111; //  497 : 255 - 0xff
      11'h1F2: dout  = 8'b11111111; //  498 : 255 - 0xff
      11'h1F3: dout  = 8'b00111000; //  499 :  56 - 0x38
      11'h1F4: dout  = 8'b01101100; //  500 : 108 - 0x6c
      11'h1F5: dout  = 8'b11000110; //  501 : 198 - 0xc6
      11'h1F6: dout  = 8'b10000011; //  502 : 131 - 0x83
      11'h1F7: dout  = 8'b11111111; //  503 : 255 - 0xff
      11'h1F8: dout  = 8'b00000000; //  504 :   0 - 0x0 -- Background 0x3f
      11'h1F9: dout  = 8'b00000000; //  505 :   0 - 0x0
      11'h1FA: dout  = 8'b00000000; //  506 :   0 - 0x0
      11'h1FB: dout  = 8'b00000000; //  507 :   0 - 0x0
      11'h1FC: dout  = 8'b00000000; //  508 :   0 - 0x0
      11'h1FD: dout  = 8'b00000000; //  509 :   0 - 0x0
      11'h1FE: dout  = 8'b00000000; //  510 :   0 - 0x0
      11'h1FF: dout  = 8'b00000000; //  511 :   0 - 0x0
      11'h200: dout  = 8'b00000000; //  512 :   0 - 0x0 -- Background 0x40
      11'h201: dout  = 8'b00000000; //  513 :   0 - 0x0
      11'h202: dout  = 8'b00000000; //  514 :   0 - 0x0
      11'h203: dout  = 8'b00000000; //  515 :   0 - 0x0
      11'h204: dout  = 8'b00000000; //  516 :   0 - 0x0
      11'h205: dout  = 8'b00000000; //  517 :   0 - 0x0
      11'h206: dout  = 8'b00000000; //  518 :   0 - 0x0
      11'h207: dout  = 8'b11111111; //  519 : 255 - 0xff
      11'h208: dout  = 8'b00000000; //  520 :   0 - 0x0 -- Background 0x41
      11'h209: dout  = 8'b00000000; //  521 :   0 - 0x0
      11'h20A: dout  = 8'b00000000; //  522 :   0 - 0x0
      11'h20B: dout  = 8'b00000000; //  523 :   0 - 0x0
      11'h20C: dout  = 8'b00000000; //  524 :   0 - 0x0
      11'h20D: dout  = 8'b11111111; //  525 : 255 - 0xff
      11'h20E: dout  = 8'b11111111; //  526 : 255 - 0xff
      11'h20F: dout  = 8'b00111000; //  527 :  56 - 0x38
      11'h210: dout  = 8'b00000000; //  528 :   0 - 0x0 -- Background 0x42
      11'h211: dout  = 8'b00000000; //  529 :   0 - 0x0
      11'h212: dout  = 8'b00000000; //  530 :   0 - 0x0
      11'h213: dout  = 8'b00000000; //  531 :   0 - 0x0
      11'h214: dout  = 8'b11111111; //  532 : 255 - 0xff
      11'h215: dout  = 8'b11111111; //  533 : 255 - 0xff
      11'h216: dout  = 8'b00111000; //  534 :  56 - 0x38
      11'h217: dout  = 8'b01101100; //  535 : 108 - 0x6c
      11'h218: dout  = 8'b00000000; //  536 :   0 - 0x0 -- Background 0x43
      11'h219: dout  = 8'b00000000; //  537 :   0 - 0x0
      11'h21A: dout  = 8'b00000000; //  538 :   0 - 0x0
      11'h21B: dout  = 8'b11111111; //  539 : 255 - 0xff
      11'h21C: dout  = 8'b11111111; //  540 : 255 - 0xff
      11'h21D: dout  = 8'b00111000; //  541 :  56 - 0x38
      11'h21E: dout  = 8'b01101100; //  542 : 108 - 0x6c
      11'h21F: dout  = 8'b11000110; //  543 : 198 - 0xc6
      11'h220: dout  = 8'b00000000; //  544 :   0 - 0x0 -- Background 0x44
      11'h221: dout  = 8'b00000000; //  545 :   0 - 0x0
      11'h222: dout  = 8'b11111111; //  546 : 255 - 0xff
      11'h223: dout  = 8'b11111111; //  547 : 255 - 0xff
      11'h224: dout  = 8'b00111000; //  548 :  56 - 0x38
      11'h225: dout  = 8'b01101100; //  549 : 108 - 0x6c
      11'h226: dout  = 8'b11000110; //  550 : 198 - 0xc6
      11'h227: dout  = 8'b10000011; //  551 : 131 - 0x83
      11'h228: dout  = 8'b00000000; //  552 :   0 - 0x0 -- Background 0x45
      11'h229: dout  = 8'b11111111; //  553 : 255 - 0xff
      11'h22A: dout  = 8'b11111111; //  554 : 255 - 0xff
      11'h22B: dout  = 8'b00111000; //  555 :  56 - 0x38
      11'h22C: dout  = 8'b01101100; //  556 : 108 - 0x6c
      11'h22D: dout  = 8'b11000110; //  557 : 198 - 0xc6
      11'h22E: dout  = 8'b10000011; //  558 : 131 - 0x83
      11'h22F: dout  = 8'b11111111; //  559 : 255 - 0xff
      11'h230: dout  = 8'b11111111; //  560 : 255 - 0xff -- Background 0x46
      11'h231: dout  = 8'b00111000; //  561 :  56 - 0x38
      11'h232: dout  = 8'b01101100; //  562 : 108 - 0x6c
      11'h233: dout  = 8'b11000110; //  563 : 198 - 0xc6
      11'h234: dout  = 8'b10000011; //  564 : 131 - 0x83
      11'h235: dout  = 8'b11111111; //  565 : 255 - 0xff
      11'h236: dout  = 8'b11111111; //  566 : 255 - 0xff
      11'h237: dout  = 8'b00000000; //  567 :   0 - 0x0
      11'h238: dout  = 8'b00111000; //  568 :  56 - 0x38 -- Background 0x47
      11'h239: dout  = 8'b01101100; //  569 : 108 - 0x6c
      11'h23A: dout  = 8'b11000110; //  570 : 198 - 0xc6
      11'h23B: dout  = 8'b10000011; //  571 : 131 - 0x83
      11'h23C: dout  = 8'b11111111; //  572 : 255 - 0xff
      11'h23D: dout  = 8'b11111111; //  573 : 255 - 0xff
      11'h23E: dout  = 8'b00000000; //  574 :   0 - 0x0
      11'h23F: dout  = 8'b00000000; //  575 :   0 - 0x0
      11'h240: dout  = 8'b01101100; //  576 : 108 - 0x6c -- Background 0x48
      11'h241: dout  = 8'b11000110; //  577 : 198 - 0xc6
      11'h242: dout  = 8'b10000011; //  578 : 131 - 0x83
      11'h243: dout  = 8'b11111111; //  579 : 255 - 0xff
      11'h244: dout  = 8'b11111111; //  580 : 255 - 0xff
      11'h245: dout  = 8'b00000000; //  581 :   0 - 0x0
      11'h246: dout  = 8'b00000000; //  582 :   0 - 0x0
      11'h247: dout  = 8'b00000000; //  583 :   0 - 0x0
      11'h248: dout  = 8'b11000110; //  584 : 198 - 0xc6 -- Background 0x49
      11'h249: dout  = 8'b10000011; //  585 : 131 - 0x83
      11'h24A: dout  = 8'b11111111; //  586 : 255 - 0xff
      11'h24B: dout  = 8'b11111111; //  587 : 255 - 0xff
      11'h24C: dout  = 8'b00000000; //  588 :   0 - 0x0
      11'h24D: dout  = 8'b00000000; //  589 :   0 - 0x0
      11'h24E: dout  = 8'b00000000; //  590 :   0 - 0x0
      11'h24F: dout  = 8'b00000000; //  591 :   0 - 0x0
      11'h250: dout  = 8'b10000011; //  592 : 131 - 0x83 -- Background 0x4a
      11'h251: dout  = 8'b11111111; //  593 : 255 - 0xff
      11'h252: dout  = 8'b11111111; //  594 : 255 - 0xff
      11'h253: dout  = 8'b00000000; //  595 :   0 - 0x0
      11'h254: dout  = 8'b00000000; //  596 :   0 - 0x0
      11'h255: dout  = 8'b00000000; //  597 :   0 - 0x0
      11'h256: dout  = 8'b00000000; //  598 :   0 - 0x0
      11'h257: dout  = 8'b00000000; //  599 :   0 - 0x0
      11'h258: dout  = 8'b11111111; //  600 : 255 - 0xff -- Background 0x4b
      11'h259: dout  = 8'b11111111; //  601 : 255 - 0xff
      11'h25A: dout  = 8'b00000000; //  602 :   0 - 0x0
      11'h25B: dout  = 8'b00000000; //  603 :   0 - 0x0
      11'h25C: dout  = 8'b00000000; //  604 :   0 - 0x0
      11'h25D: dout  = 8'b00000000; //  605 :   0 - 0x0
      11'h25E: dout  = 8'b00000000; //  606 :   0 - 0x0
      11'h25F: dout  = 8'b00000000; //  607 :   0 - 0x0
      11'h260: dout  = 8'b10111111; //  608 : 191 - 0xbf -- Background 0x4c
      11'h261: dout  = 8'b01011111; //  609 :  95 - 0x5f
      11'h262: dout  = 8'b01011111; //  610 :  95 - 0x5f
      11'h263: dout  = 8'b01011111; //  611 :  95 - 0x5f
      11'h264: dout  = 8'b00000000; //  612 :   0 - 0x0
      11'h265: dout  = 8'b01011111; //  613 :  95 - 0x5f
      11'h266: dout  = 8'b01010001; //  614 :  81 - 0x51
      11'h267: dout  = 8'b01010101; //  615 :  85 - 0x55
      11'h268: dout  = 8'b01010001; //  616 :  81 - 0x51 -- Background 0x4d
      11'h269: dout  = 8'b01011111; //  617 :  95 - 0x5f
      11'h26A: dout  = 8'b00000000; //  618 :   0 - 0x0
      11'h26B: dout  = 8'b01011111; //  619 :  95 - 0x5f
      11'h26C: dout  = 8'b01011111; //  620 :  95 - 0x5f
      11'h26D: dout  = 8'b01011111; //  621 :  95 - 0x5f
      11'h26E: dout  = 8'b01011111; //  622 :  95 - 0x5f
      11'h26F: dout  = 8'b10111111; //  623 : 191 - 0xbf
      11'h270: dout  = 8'b11111111; //  624 : 255 - 0xff -- Background 0x4e
      11'h271: dout  = 8'b11111110; //  625 : 254 - 0xfe
      11'h272: dout  = 8'b11111110; //  626 : 254 - 0xfe
      11'h273: dout  = 8'b11111110; //  627 : 254 - 0xfe
      11'h274: dout  = 8'b00000000; //  628 :   0 - 0x0
      11'h275: dout  = 8'b11111110; //  629 : 254 - 0xfe
      11'h276: dout  = 8'b00100110; //  630 :  38 - 0x26
      11'h277: dout  = 8'b00100110; //  631 :  38 - 0x26
      11'h278: dout  = 8'b00100010; //  632 :  34 - 0x22 -- Background 0x4f
      11'h279: dout  = 8'b11111110; //  633 : 254 - 0xfe
      11'h27A: dout  = 8'b00000000; //  634 :   0 - 0x0
      11'h27B: dout  = 8'b11111110; //  635 : 254 - 0xfe
      11'h27C: dout  = 8'b11111110; //  636 : 254 - 0xfe
      11'h27D: dout  = 8'b11111110; //  637 : 254 - 0xfe
      11'h27E: dout  = 8'b11111110; //  638 : 254 - 0xfe
      11'h27F: dout  = 8'b11111111; //  639 : 255 - 0xff
      11'h280: dout  = 8'b00000111; //  640 :   7 - 0x7 -- Background 0x50
      11'h281: dout  = 8'b00000000; //  641 :   0 - 0x0
      11'h282: dout  = 8'b00001111; //  642 :  15 - 0xf
      11'h283: dout  = 8'b00011111; //  643 :  31 - 0x1f
      11'h284: dout  = 8'b00011111; //  644 :  31 - 0x1f
      11'h285: dout  = 8'b00011111; //  645 :  31 - 0x1f
      11'h286: dout  = 8'b00011111; //  646 :  31 - 0x1f
      11'h287: dout  = 8'b00011111; //  647 :  31 - 0x1f
      11'h288: dout  = 8'b00011111; //  648 :  31 - 0x1f -- Background 0x51
      11'h289: dout  = 8'b00011111; //  649 :  31 - 0x1f
      11'h28A: dout  = 8'b00011111; //  650 :  31 - 0x1f
      11'h28B: dout  = 8'b00011111; //  651 :  31 - 0x1f
      11'h28C: dout  = 8'b00011111; //  652 :  31 - 0x1f
      11'h28D: dout  = 8'b00001111; //  653 :  15 - 0xf
      11'h28E: dout  = 8'b00000000; //  654 :   0 - 0x0
      11'h28F: dout  = 8'b00000111; //  655 :   7 - 0x7
      11'h290: dout  = 8'b00000111; //  656 :   7 - 0x7 -- Background 0x52
      11'h291: dout  = 8'b00000000; //  657 :   0 - 0x0
      11'h292: dout  = 8'b00001111; //  658 :  15 - 0xf
      11'h293: dout  = 8'b00011111; //  659 :  31 - 0x1f
      11'h294: dout  = 8'b00011111; //  660 :  31 - 0x1f
      11'h295: dout  = 8'b00011111; //  661 :  31 - 0x1f
      11'h296: dout  = 8'b00011111; //  662 :  31 - 0x1f
      11'h297: dout  = 8'b00011111; //  663 :  31 - 0x1f
      11'h298: dout  = 8'b00011111; //  664 :  31 - 0x1f -- Background 0x53
      11'h299: dout  = 8'b00011111; //  665 :  31 - 0x1f
      11'h29A: dout  = 8'b00011111; //  666 :  31 - 0x1f
      11'h29B: dout  = 8'b00011111; //  667 :  31 - 0x1f
      11'h29C: dout  = 8'b00011111; //  668 :  31 - 0x1f
      11'h29D: dout  = 8'b00001111; //  669 :  15 - 0xf
      11'h29E: dout  = 8'b00000000; //  670 :   0 - 0x0
      11'h29F: dout  = 8'b00000111; //  671 :   7 - 0x7
      11'h2A0: dout  = 8'b11100000; //  672 : 224 - 0xe0 -- Background 0x54
      11'h2A1: dout  = 8'b00000000; //  673 :   0 - 0x0
      11'h2A2: dout  = 8'b11110001; //  674 : 241 - 0xf1
      11'h2A3: dout  = 8'b11111011; //  675 : 251 - 0xfb
      11'h2A4: dout  = 8'b11111011; //  676 : 251 - 0xfb
      11'h2A5: dout  = 8'b11111011; //  677 : 251 - 0xfb
      11'h2A6: dout  = 8'b11111011; //  678 : 251 - 0xfb
      11'h2A7: dout  = 8'b11111011; //  679 : 251 - 0xfb
      11'h2A8: dout  = 8'b11111011; //  680 : 251 - 0xfb -- Background 0x55
      11'h2A9: dout  = 8'b11111011; //  681 : 251 - 0xfb
      11'h2AA: dout  = 8'b11111011; //  682 : 251 - 0xfb
      11'h2AB: dout  = 8'b11111011; //  683 : 251 - 0xfb
      11'h2AC: dout  = 8'b11111011; //  684 : 251 - 0xfb
      11'h2AD: dout  = 8'b11110001; //  685 : 241 - 0xf1
      11'h2AE: dout  = 8'b00000000; //  686 :   0 - 0x0
      11'h2AF: dout  = 8'b11100000; //  687 : 224 - 0xe0
      11'h2B0: dout  = 8'b11100000; //  688 : 224 - 0xe0 -- Background 0x56
      11'h2B1: dout  = 8'b00000000; //  689 :   0 - 0x0
      11'h2B2: dout  = 8'b11110001; //  690 : 241 - 0xf1
      11'h2B3: dout  = 8'b11111011; //  691 : 251 - 0xfb
      11'h2B4: dout  = 8'b11111011; //  692 : 251 - 0xfb
      11'h2B5: dout  = 8'b11111011; //  693 : 251 - 0xfb
      11'h2B6: dout  = 8'b11111011; //  694 : 251 - 0xfb
      11'h2B7: dout  = 8'b11111011; //  695 : 251 - 0xfb
      11'h2B8: dout  = 8'b11111011; //  696 : 251 - 0xfb -- Background 0x57
      11'h2B9: dout  = 8'b11111011; //  697 : 251 - 0xfb
      11'h2BA: dout  = 8'b11111011; //  698 : 251 - 0xfb
      11'h2BB: dout  = 8'b11111011; //  699 : 251 - 0xfb
      11'h2BC: dout  = 8'b11111011; //  700 : 251 - 0xfb
      11'h2BD: dout  = 8'b11110001; //  701 : 241 - 0xf1
      11'h2BE: dout  = 8'b00000000; //  702 :   0 - 0x0
      11'h2BF: dout  = 8'b11100000; //  703 : 224 - 0xe0
      11'h2C0: dout  = 8'b11111100; //  704 : 252 - 0xfc -- Background 0x58
      11'h2C1: dout  = 8'b00000000; //  705 :   0 - 0x0
      11'h2C2: dout  = 8'b11111110; //  706 : 254 - 0xfe
      11'h2C3: dout  = 8'b11111111; //  707 : 255 - 0xff
      11'h2C4: dout  = 8'b11111111; //  708 : 255 - 0xff
      11'h2C5: dout  = 8'b11111111; //  709 : 255 - 0xff
      11'h2C6: dout  = 8'b11111111; //  710 : 255 - 0xff
      11'h2C7: dout  = 8'b11111111; //  711 : 255 - 0xff
      11'h2C8: dout  = 8'b11111111; //  712 : 255 - 0xff -- Background 0x59
      11'h2C9: dout  = 8'b11111111; //  713 : 255 - 0xff
      11'h2CA: dout  = 8'b11111111; //  714 : 255 - 0xff
      11'h2CB: dout  = 8'b11111111; //  715 : 255 - 0xff
      11'h2CC: dout  = 8'b11111111; //  716 : 255 - 0xff
      11'h2CD: dout  = 8'b11111110; //  717 : 254 - 0xfe
      11'h2CE: dout  = 8'b00000000; //  718 :   0 - 0x0
      11'h2CF: dout  = 8'b11111100; //  719 : 252 - 0xfc
      11'h2D0: dout  = 8'b11111100; //  720 : 252 - 0xfc -- Background 0x5a
      11'h2D1: dout  = 8'b00000000; //  721 :   0 - 0x0
      11'h2D2: dout  = 8'b11111110; //  722 : 254 - 0xfe
      11'h2D3: dout  = 8'b11111111; //  723 : 255 - 0xff
      11'h2D4: dout  = 8'b11111111; //  724 : 255 - 0xff
      11'h2D5: dout  = 8'b11111111; //  725 : 255 - 0xff
      11'h2D6: dout  = 8'b11111111; //  726 : 255 - 0xff
      11'h2D7: dout  = 8'b11111111; //  727 : 255 - 0xff
      11'h2D8: dout  = 8'b11111111; //  728 : 255 - 0xff -- Background 0x5b
      11'h2D9: dout  = 8'b11111111; //  729 : 255 - 0xff
      11'h2DA: dout  = 8'b11111111; //  730 : 255 - 0xff
      11'h2DB: dout  = 8'b11111111; //  731 : 255 - 0xff
      11'h2DC: dout  = 8'b11111111; //  732 : 255 - 0xff
      11'h2DD: dout  = 8'b11111110; //  733 : 254 - 0xfe
      11'h2DE: dout  = 8'b00000000; //  734 :   0 - 0x0
      11'h2DF: dout  = 8'b11111100; //  735 : 252 - 0xfc
      11'h2E0: dout  = 8'b00000000; //  736 :   0 - 0x0 -- Background 0x5c
      11'h2E1: dout  = 8'b00000000; //  737 :   0 - 0x0
      11'h2E2: dout  = 8'b00011111; //  738 :  31 - 0x1f
      11'h2E3: dout  = 8'b00010000; //  739 :  16 - 0x10
      11'h2E4: dout  = 8'b00010000; //  740 :  16 - 0x10
      11'h2E5: dout  = 8'b00011111; //  741 :  31 - 0x1f
      11'h2E6: dout  = 8'b00000000; //  742 :   0 - 0x0
      11'h2E7: dout  = 8'b00000000; //  743 :   0 - 0x0
      11'h2E8: dout  = 8'b00000000; //  744 :   0 - 0x0 -- Background 0x5d
      11'h2E9: dout  = 8'b00000000; //  745 :   0 - 0x0
      11'h2EA: dout  = 8'b11111000; //  746 : 248 - 0xf8
      11'h2EB: dout  = 8'b00001000; //  747 :   8 - 0x8
      11'h2EC: dout  = 8'b00001000; //  748 :   8 - 0x8
      11'h2ED: dout  = 8'b11111000; //  749 : 248 - 0xf8
      11'h2EE: dout  = 8'b00000000; //  750 :   0 - 0x0
      11'h2EF: dout  = 8'b00000000; //  751 :   0 - 0x0
      11'h2F0: dout  = 8'b00000000; //  752 :   0 - 0x0 -- Background 0x5e
      11'h2F1: dout  = 8'b00000001; //  753 :   1 - 0x1
      11'h2F2: dout  = 8'b00000010; //  754 :   2 - 0x2
      11'h2F3: dout  = 8'b00000010; //  755 :   2 - 0x2
      11'h2F4: dout  = 8'b11110001; //  756 : 241 - 0xf1
      11'h2F5: dout  = 8'b00001000; //  757 :   8 - 0x8
      11'h2F6: dout  = 8'b00000100; //  758 :   4 - 0x4
      11'h2F7: dout  = 8'b00000011; //  759 :   3 - 0x3
      11'h2F8: dout  = 8'b00000000; //  760 :   0 - 0x0 -- Background 0x5f
      11'h2F9: dout  = 8'b10000000; //  761 : 128 - 0x80
      11'h2FA: dout  = 8'b01000000; //  762 :  64 - 0x40
      11'h2FB: dout  = 8'b01000000; //  763 :  64 - 0x40
      11'h2FC: dout  = 8'b10001111; //  764 : 143 - 0x8f
      11'h2FD: dout  = 8'b00010000; //  765 :  16 - 0x10
      11'h2FE: dout  = 8'b00100000; //  766 :  32 - 0x20
      11'h2FF: dout  = 8'b11000000; //  767 : 192 - 0xc0
      11'h300: dout  = 8'b00000011; //  768 :   3 - 0x3 -- Background 0x60
      11'h301: dout  = 8'b00000100; //  769 :   4 - 0x4
      11'h302: dout  = 8'b00001000; //  770 :   8 - 0x8
      11'h303: dout  = 8'b11110001; //  771 : 241 - 0xf1
      11'h304: dout  = 8'b00000010; //  772 :   2 - 0x2
      11'h305: dout  = 8'b00000010; //  773 :   2 - 0x2
      11'h306: dout  = 8'b00000001; //  774 :   1 - 0x1
      11'h307: dout  = 8'b00000000; //  775 :   0 - 0x0
      11'h308: dout  = 8'b11000000; //  776 : 192 - 0xc0 -- Background 0x61
      11'h309: dout  = 8'b00100000; //  777 :  32 - 0x20
      11'h30A: dout  = 8'b00010000; //  778 :  16 - 0x10
      11'h30B: dout  = 8'b10001111; //  779 : 143 - 0x8f
      11'h30C: dout  = 8'b01000000; //  780 :  64 - 0x40
      11'h30D: dout  = 8'b01000000; //  781 :  64 - 0x40
      11'h30E: dout  = 8'b10000000; //  782 : 128 - 0x80
      11'h30F: dout  = 8'b00000000; //  783 :   0 - 0x0
      11'h310: dout  = 8'b11111111; //  784 : 255 - 0xff -- Background 0x62
      11'h311: dout  = 8'b11111111; //  785 : 255 - 0xff
      11'h312: dout  = 8'b11000011; //  786 : 195 - 0xc3
      11'h313: dout  = 8'b10000001; //  787 : 129 - 0x81
      11'h314: dout  = 8'b10000001; //  788 : 129 - 0x81
      11'h315: dout  = 8'b11000011; //  789 : 195 - 0xc3
      11'h316: dout  = 8'b11111111; //  790 : 255 - 0xff
      11'h317: dout  = 8'b11111111; //  791 : 255 - 0xff
      11'h318: dout  = 8'b11111111; //  792 : 255 - 0xff -- Background 0x63
      11'h319: dout  = 8'b10011001; //  793 : 153 - 0x99
      11'h31A: dout  = 8'b00000000; //  794 :   0 - 0x0
      11'h31B: dout  = 8'b00000000; //  795 :   0 - 0x0
      11'h31C: dout  = 8'b00000000; //  796 :   0 - 0x0
      11'h31D: dout  = 8'b10000001; //  797 : 129 - 0x81
      11'h31E: dout  = 8'b10000001; //  798 : 129 - 0x81
      11'h31F: dout  = 8'b10000001; //  799 : 129 - 0x81
      11'h320: dout  = 8'b00000000; //  800 :   0 - 0x0 -- Background 0x64
      11'h321: dout  = 8'b00000000; //  801 :   0 - 0x0
      11'h322: dout  = 8'b00000000; //  802 :   0 - 0x0
      11'h323: dout  = 8'b00000000; //  803 :   0 - 0x0
      11'h324: dout  = 8'b01100000; //  804 :  96 - 0x60
      11'h325: dout  = 8'b01100000; //  805 :  96 - 0x60
      11'h326: dout  = 8'b00000000; //  806 :   0 - 0x0
      11'h327: dout  = 8'b00000000; //  807 :   0 - 0x0
      11'h328: dout  = 8'b00000000; //  808 :   0 - 0x0 -- Background 0x65
      11'h329: dout  = 8'b00000000; //  809 :   0 - 0x0
      11'h32A: dout  = 8'b00000000; //  810 :   0 - 0x0
      11'h32B: dout  = 8'b00000000; //  811 :   0 - 0x0
      11'h32C: dout  = 8'b01101100; //  812 : 108 - 0x6c
      11'h32D: dout  = 8'b01101100; //  813 : 108 - 0x6c
      11'h32E: dout  = 8'b00001000; //  814 :   8 - 0x8
      11'h32F: dout  = 8'b00000000; //  815 :   0 - 0x0
      11'h330: dout  = 8'b00111100; //  816 :  60 - 0x3c -- Background 0x66
      11'h331: dout  = 8'b00011000; //  817 :  24 - 0x18
      11'h332: dout  = 8'b00011000; //  818 :  24 - 0x18
      11'h333: dout  = 8'b00011000; //  819 :  24 - 0x18
      11'h334: dout  = 8'b00011000; //  820 :  24 - 0x18
      11'h335: dout  = 8'b00011000; //  821 :  24 - 0x18
      11'h336: dout  = 8'b00111100; //  822 :  60 - 0x3c
      11'h337: dout  = 8'b00000000; //  823 :   0 - 0x0
      11'h338: dout  = 8'b11111111; //  824 : 255 - 0xff -- Background 0x67
      11'h339: dout  = 8'b01100110; //  825 : 102 - 0x66
      11'h33A: dout  = 8'b01100110; //  826 : 102 - 0x66
      11'h33B: dout  = 8'b01100110; //  827 : 102 - 0x66
      11'h33C: dout  = 8'b01100110; //  828 : 102 - 0x66
      11'h33D: dout  = 8'b01100110; //  829 : 102 - 0x66
      11'h33E: dout  = 8'b01100110; //  830 : 102 - 0x66
      11'h33F: dout  = 8'b11111111; //  831 : 255 - 0xff
      11'h340: dout  = 8'b00000011; //  832 :   3 - 0x3 -- Background 0x68
      11'h341: dout  = 8'b00000001; //  833 :   1 - 0x1
      11'h342: dout  = 8'b00000000; //  834 :   0 - 0x0
      11'h343: dout  = 8'b00000000; //  835 :   0 - 0x0
      11'h344: dout  = 8'b00000000; //  836 :   0 - 0x0
      11'h345: dout  = 8'b00000000; //  837 :   0 - 0x0
      11'h346: dout  = 8'b00000000; //  838 :   0 - 0x0
      11'h347: dout  = 8'b00000000; //  839 :   0 - 0x0
      11'h348: dout  = 8'b10000011; //  840 : 131 - 0x83 -- Background 0x69
      11'h349: dout  = 8'b11010001; //  841 : 209 - 0xd1
      11'h34A: dout  = 8'b11100001; //  842 : 225 - 0xe1
      11'h34B: dout  = 8'b11010001; //  843 : 209 - 0xd1
      11'h34C: dout  = 8'b00000010; //  844 :   2 - 0x2
      11'h34D: dout  = 8'b10000100; //  845 : 132 - 0x84
      11'h34E: dout  = 8'b11110000; //  846 : 240 - 0xf0
      11'h34F: dout  = 8'b11001110; //  847 : 206 - 0xce
      11'h350: dout  = 8'b11000000; //  848 : 192 - 0xc0 -- Background 0x6a
      11'h351: dout  = 8'b10000000; //  849 : 128 - 0x80
      11'h352: dout  = 8'b00000000; //  850 :   0 - 0x0
      11'h353: dout  = 8'b00000000; //  851 :   0 - 0x0
      11'h354: dout  = 8'b00000000; //  852 :   0 - 0x0
      11'h355: dout  = 8'b00000000; //  853 :   0 - 0x0
      11'h356: dout  = 8'b00000000; //  854 :   0 - 0x0
      11'h357: dout  = 8'b00000000; //  855 :   0 - 0x0
      11'h358: dout  = 8'b11000001; //  856 : 193 - 0xc1 -- Background 0x6b
      11'h359: dout  = 8'b10001011; //  857 : 139 - 0x8b
      11'h35A: dout  = 8'b10000111; //  858 : 135 - 0x87
      11'h35B: dout  = 8'b10001011; //  859 : 139 - 0x8b
      11'h35C: dout  = 8'b01000000; //  860 :  64 - 0x40
      11'h35D: dout  = 8'b00100001; //  861 :  33 - 0x21
      11'h35E: dout  = 8'b00001111; //  862 :  15 - 0xf
      11'h35F: dout  = 8'b11010011; //  863 : 211 - 0xd3
      11'h360: dout  = 8'b11111111; //  864 : 255 - 0xff -- Background 0x6c
      11'h361: dout  = 8'b11111111; //  865 : 255 - 0xff
      11'h362: dout  = 8'b11111111; //  866 : 255 - 0xff
      11'h363: dout  = 8'b00011111; //  867 :  31 - 0x1f
      11'h364: dout  = 8'b00001111; //  868 :  15 - 0xf
      11'h365: dout  = 8'b00011110; //  869 :  30 - 0x1e
      11'h366: dout  = 8'b00111111; //  870 :  63 - 0x3f
      11'h367: dout  = 8'b01111111; //  871 : 127 - 0x7f
      11'h368: dout  = 8'b11111111; //  872 : 255 - 0xff -- Background 0x6d
      11'h369: dout  = 8'b11111111; //  873 : 255 - 0xff
      11'h36A: dout  = 8'b11111111; //  874 : 255 - 0xff
      11'h36B: dout  = 8'b11111000; //  875 : 248 - 0xf8
      11'h36C: dout  = 8'b11110000; //  876 : 240 - 0xf0
      11'h36D: dout  = 8'b01111000; //  877 : 120 - 0x78
      11'h36E: dout  = 8'b11111100; //  878 : 252 - 0xfc
      11'h36F: dout  = 8'b11111110; //  879 : 254 - 0xfe
      11'h370: dout  = 8'b00000000; //  880 :   0 - 0x0 -- Background 0x6e
      11'h371: dout  = 8'b00000000; //  881 :   0 - 0x0
      11'h372: dout  = 8'b00000000; //  882 :   0 - 0x0
      11'h373: dout  = 8'b00000000; //  883 :   0 - 0x0
      11'h374: dout  = 8'b00000000; //  884 :   0 - 0x0
      11'h375: dout  = 8'b00111100; //  885 :  60 - 0x3c
      11'h376: dout  = 8'b01000010; //  886 :  66 - 0x42
      11'h377: dout  = 8'b10000001; //  887 : 129 - 0x81
      11'h378: dout  = 8'b10000001; //  888 : 129 - 0x81 -- Background 0x6f
      11'h379: dout  = 8'b10111101; //  889 : 189 - 0xbd
      11'h37A: dout  = 8'b01111110; //  890 : 126 - 0x7e
      11'h37B: dout  = 8'b11111111; //  891 : 255 - 0xff
      11'h37C: dout  = 8'b11100111; //  892 : 231 - 0xe7
      11'h37D: dout  = 8'b11111111; //  893 : 255 - 0xff
      11'h37E: dout  = 8'b11111111; //  894 : 255 - 0xff
      11'h37F: dout  = 8'b11111111; //  895 : 255 - 0xff
      11'h380: dout  = 8'b00000001; //  896 :   1 - 0x1 -- Background 0x70
      11'h381: dout  = 8'b00000111; //  897 :   7 - 0x7
      11'h382: dout  = 8'b00011111; //  898 :  31 - 0x1f
      11'h383: dout  = 8'b00111111; //  899 :  63 - 0x3f
      11'h384: dout  = 8'b01111111; //  900 : 127 - 0x7f
      11'h385: dout  = 8'b11111111; //  901 : 255 - 0xff
      11'h386: dout  = 8'b11111111; //  902 : 255 - 0xff
      11'h387: dout  = 8'b11011101; //  903 : 221 - 0xdd
      11'h388: dout  = 8'b10001001; //  904 : 137 - 0x89 -- Background 0x71
      11'h389: dout  = 8'b00000001; //  905 :   1 - 0x1
      11'h38A: dout  = 8'b00000001; //  906 :   1 - 0x1
      11'h38B: dout  = 8'b00000001; //  907 :   1 - 0x1
      11'h38C: dout  = 8'b00000001; //  908 :   1 - 0x1
      11'h38D: dout  = 8'b00000001; //  909 :   1 - 0x1
      11'h38E: dout  = 8'b00000000; //  910 :   0 - 0x0
      11'h38F: dout  = 8'b00000000; //  911 :   0 - 0x0
      11'h390: dout  = 8'b10000000; //  912 : 128 - 0x80 -- Background 0x72
      11'h391: dout  = 8'b11100000; //  913 : 224 - 0xe0
      11'h392: dout  = 8'b11111000; //  914 : 248 - 0xf8
      11'h393: dout  = 8'b11111100; //  915 : 252 - 0xfc
      11'h394: dout  = 8'b11111110; //  916 : 254 - 0xfe
      11'h395: dout  = 8'b11111111; //  917 : 255 - 0xff
      11'h396: dout  = 8'b11111111; //  918 : 255 - 0xff
      11'h397: dout  = 8'b00111011; //  919 :  59 - 0x3b
      11'h398: dout  = 8'b00010001; //  920 :  17 - 0x11 -- Background 0x73
      11'h399: dout  = 8'b00000000; //  921 :   0 - 0x0
      11'h39A: dout  = 8'b00000000; //  922 :   0 - 0x0
      11'h39B: dout  = 8'b00000000; //  923 :   0 - 0x0
      11'h39C: dout  = 8'b00000000; //  924 :   0 - 0x0
      11'h39D: dout  = 8'b01000000; //  925 :  64 - 0x40
      11'h39E: dout  = 8'b10000000; //  926 : 128 - 0x80
      11'h39F: dout  = 8'b00000000; //  927 :   0 - 0x0
      11'h3A0: dout  = 8'b00000001; //  928 :   1 - 0x1 -- Background 0x74
      11'h3A1: dout  = 8'b00000001; //  929 :   1 - 0x1
      11'h3A2: dout  = 8'b00000001; //  930 :   1 - 0x1
      11'h3A3: dout  = 8'b00000001; //  931 :   1 - 0x1
      11'h3A4: dout  = 8'b00000001; //  932 :   1 - 0x1
      11'h3A5: dout  = 8'b00000001; //  933 :   1 - 0x1
      11'h3A6: dout  = 8'b00000001; //  934 :   1 - 0x1
      11'h3A7: dout  = 8'b00000001; //  935 :   1 - 0x1
      11'h3A8: dout  = 8'b10000000; //  936 : 128 - 0x80 -- Background 0x75
      11'h3A9: dout  = 8'b10000000; //  937 : 128 - 0x80
      11'h3AA: dout  = 8'b10000000; //  938 : 128 - 0x80
      11'h3AB: dout  = 8'b10000000; //  939 : 128 - 0x80
      11'h3AC: dout  = 8'b10000000; //  940 : 128 - 0x80
      11'h3AD: dout  = 8'b10000000; //  941 : 128 - 0x80
      11'h3AE: dout  = 8'b10000000; //  942 : 128 - 0x80
      11'h3AF: dout  = 8'b10000000; //  943 : 128 - 0x80
      11'h3B0: dout  = 8'b00000001; //  944 :   1 - 0x1 -- Background 0x76
      11'h3B1: dout  = 8'b00000011; //  945 :   3 - 0x3
      11'h3B2: dout  = 8'b00000000; //  946 :   0 - 0x0
      11'h3B3: dout  = 8'b00000000; //  947 :   0 - 0x0
      11'h3B4: dout  = 8'b00000011; //  948 :   3 - 0x3
      11'h3B5: dout  = 8'b00011001; //  949 :  25 - 0x19
      11'h3B6: dout  = 8'b00000000; //  950 :   0 - 0x0
      11'h3B7: dout  = 8'b00000000; //  951 :   0 - 0x0
      11'h3B8: dout  = 8'b00000000; //  952 :   0 - 0x0 -- Background 0x77
      11'h3B9: dout  = 8'b00000000; //  953 :   0 - 0x0
      11'h3BA: dout  = 8'b01111100; //  954 : 124 - 0x7c
      11'h3BB: dout  = 8'b00000010; //  955 :   2 - 0x2
      11'h3BC: dout  = 8'b00000001; //  956 :   1 - 0x1
      11'h3BD: dout  = 8'b00000000; //  957 :   0 - 0x0
      11'h3BE: dout  = 8'b00000000; //  958 :   0 - 0x0
      11'h3BF: dout  = 8'b00000000; //  959 :   0 - 0x0
      11'h3C0: dout  = 8'b00000000; //  960 :   0 - 0x0 -- Background 0x78
      11'h3C1: dout  = 8'b00000000; //  961 :   0 - 0x0
      11'h3C2: dout  = 8'b00000001; //  962 :   1 - 0x1
      11'h3C3: dout  = 8'b00000001; //  963 :   1 - 0x1
      11'h3C4: dout  = 8'b00000011; //  964 :   3 - 0x3
      11'h3C5: dout  = 8'b00000111; //  965 :   7 - 0x7
      11'h3C6: dout  = 8'b00000111; //  966 :   7 - 0x7
      11'h3C7: dout  = 8'b00001111; //  967 :  15 - 0xf
      11'h3C8: dout  = 8'b00001111; //  968 :  15 - 0xf -- Background 0x79
      11'h3C9: dout  = 8'b00000111; //  969 :   7 - 0x7
      11'h3CA: dout  = 8'b00001111; //  970 :  15 - 0xf
      11'h3CB: dout  = 8'b00000111; //  971 :   7 - 0x7
      11'h3CC: dout  = 8'b00000001; //  972 :   1 - 0x1
      11'h3CD: dout  = 8'b00010000; //  973 :  16 - 0x10
      11'h3CE: dout  = 8'b00100000; //  974 :  32 - 0x20
      11'h3CF: dout  = 8'b00000000; //  975 :   0 - 0x0
      11'h3D0: dout  = 8'b11111000; //  976 : 248 - 0xf8 -- Background 0x7a
      11'h3D1: dout  = 8'b11111110; //  977 : 254 - 0xfe
      11'h3D2: dout  = 8'b01111111; //  978 : 127 - 0x7f
      11'h3D3: dout  = 8'b00011111; //  979 :  31 - 0x1f
      11'h3D4: dout  = 8'b00001111; //  980 :  15 - 0xf
      11'h3D5: dout  = 8'b00011001; //  981 :  25 - 0x19
      11'h3D6: dout  = 8'b00110000; //  982 :  48 - 0x30
      11'h3D7: dout  = 8'b01110000; //  983 : 112 - 0x70
      11'h3D8: dout  = 8'b11111011; //  984 : 251 - 0xfb -- Background 0x7b
      11'h3D9: dout  = 8'b01110011; //  985 : 115 - 0x73
      11'h3DA: dout  = 8'b00100111; //  986 :  39 - 0x27
      11'h3DB: dout  = 8'b00001111; //  987 :  15 - 0xf
      11'h3DC: dout  = 8'b00011111; //  988 :  31 - 0x1f
      11'h3DD: dout  = 8'b00011111; //  989 :  31 - 0x1f
      11'h3DE: dout  = 8'b00111111; //  990 :  63 - 0x3f
      11'h3DF: dout  = 8'b01111111; //  991 : 127 - 0x7f
      11'h3E0: dout  = 8'b11111111; //  992 : 255 - 0xff -- Background 0x7c
      11'h3E1: dout  = 8'b11111111; //  993 : 255 - 0xff
      11'h3E2: dout  = 8'b11111111; //  994 : 255 - 0xff
      11'h3E3: dout  = 8'b11111111; //  995 : 255 - 0xff
      11'h3E4: dout  = 8'b11111110; //  996 : 254 - 0xfe
      11'h3E5: dout  = 8'b11111101; //  997 : 253 - 0xfd
      11'h3E6: dout  = 8'b11111000; //  998 : 248 - 0xf8
      11'h3E7: dout  = 8'b11110110; //  999 : 246 - 0xf6
      11'h3E8: dout  = 8'b11101111; // 1000 : 239 - 0xef -- Background 0x7d
      11'h3E9: dout  = 8'b11001111; // 1001 : 207 - 0xcf
      11'h3EA: dout  = 8'b10011111; // 1002 : 159 - 0x9f
      11'h3EB: dout  = 8'b00011111; // 1003 :  31 - 0x1f
      11'h3EC: dout  = 8'b00001111; // 1004 :  15 - 0xf
      11'h3ED: dout  = 8'b00101101; // 1005 :  45 - 0x2d
      11'h3EE: dout  = 8'b01010000; // 1006 :  80 - 0x50
      11'h3EF: dout  = 8'b01000000; // 1007 :  64 - 0x40
      11'h3F0: dout  = 8'b00000000; // 1008 :   0 - 0x0 -- Background 0x7e
      11'h3F1: dout  = 8'b00000000; // 1009 :   0 - 0x0
      11'h3F2: dout  = 8'b00000000; // 1010 :   0 - 0x0
      11'h3F3: dout  = 8'b00000000; // 1011 :   0 - 0x0
      11'h3F4: dout  = 8'b11100000; // 1012 : 224 - 0xe0
      11'h3F5: dout  = 8'b11111110; // 1013 : 254 - 0xfe
      11'h3F6: dout  = 8'b11111111; // 1014 : 255 - 0xff
      11'h3F7: dout  = 8'b11110011; // 1015 : 243 - 0xf3
      11'h3F8: dout  = 8'b11111011; // 1016 : 251 - 0xfb -- Background 0x7f
      11'h3F9: dout  = 8'b11111011; // 1017 : 251 - 0xfb
      11'h3FA: dout  = 8'b11111011; // 1018 : 251 - 0xfb
      11'h3FB: dout  = 8'b11111011; // 1019 : 251 - 0xfb
      11'h3FC: dout  = 8'b11111011; // 1020 : 251 - 0xfb
      11'h3FD: dout  = 8'b11110011; // 1021 : 243 - 0xf3
      11'h3FE: dout  = 8'b11110111; // 1022 : 247 - 0xf7
      11'h3FF: dout  = 8'b11100111; // 1023 : 231 - 0xe7
      11'h400: dout  = 8'b11001111; // 1024 : 207 - 0xcf -- Background 0x80
      11'h401: dout  = 8'b10011111; // 1025 : 159 - 0x9f
      11'h402: dout  = 8'b00111111; // 1026 :  63 - 0x3f
      11'h403: dout  = 8'b00111111; // 1027 :  63 - 0x3f
      11'h404: dout  = 8'b00111111; // 1028 :  63 - 0x3f
      11'h405: dout  = 8'b00001111; // 1029 :  15 - 0xf
      11'h406: dout  = 8'b00000011; // 1030 :   3 - 0x3
      11'h407: dout  = 8'b00000000; // 1031 :   0 - 0x0
      11'h408: dout  = 8'b11000000; // 1032 : 192 - 0xc0 -- Background 0x81
      11'h409: dout  = 8'b11110000; // 1033 : 240 - 0xf0
      11'h40A: dout  = 8'b11111100; // 1034 : 252 - 0xfc
      11'h40B: dout  = 8'b11110000; // 1035 : 240 - 0xf0
      11'h40C: dout  = 8'b11110000; // 1036 : 240 - 0xf0
      11'h40D: dout  = 8'b10011000; // 1037 : 152 - 0x98
      11'h40E: dout  = 8'b00001000; // 1038 :   8 - 0x8
      11'h40F: dout  = 8'b00000000; // 1039 :   0 - 0x0
      11'h410: dout  = 8'b00000000; // 1040 :   0 - 0x0 -- Background 0x82
      11'h411: dout  = 8'b00000000; // 1041 :   0 - 0x0
      11'h412: dout  = 8'b00000000; // 1042 :   0 - 0x0
      11'h413: dout  = 8'b00000000; // 1043 :   0 - 0x0
      11'h414: dout  = 8'b00000000; // 1044 :   0 - 0x0
      11'h415: dout  = 8'b00000000; // 1045 :   0 - 0x0
      11'h416: dout  = 8'b10000000; // 1046 : 128 - 0x80
      11'h417: dout  = 8'b11000000; // 1047 : 192 - 0xc0
      11'h418: dout  = 8'b11100000; // 1048 : 224 - 0xe0 -- Background 0x83
      11'h419: dout  = 8'b11100000; // 1049 : 224 - 0xe0
      11'h41A: dout  = 8'b11110000; // 1050 : 240 - 0xf0
      11'h41B: dout  = 8'b11110000; // 1051 : 240 - 0xf0
      11'h41C: dout  = 8'b11110000; // 1052 : 240 - 0xf0
      11'h41D: dout  = 8'b11110000; // 1053 : 240 - 0xf0
      11'h41E: dout  = 8'b11111000; // 1054 : 248 - 0xf8
      11'h41F: dout  = 8'b11111000; // 1055 : 248 - 0xf8
      11'h420: dout  = 8'b11111110; // 1056 : 254 - 0xfe -- Background 0x84
      11'h421: dout  = 8'b11111111; // 1057 : 255 - 0xff
      11'h422: dout  = 8'b11111111; // 1058 : 255 - 0xff
      11'h423: dout  = 8'b11111111; // 1059 : 255 - 0xff
      11'h424: dout  = 8'b11111111; // 1060 : 255 - 0xff
      11'h425: dout  = 8'b11111111; // 1061 : 255 - 0xff
      11'h426: dout  = 8'b11111111; // 1062 : 255 - 0xff
      11'h427: dout  = 8'b11111111; // 1063 : 255 - 0xff
      11'h428: dout  = 8'b00111111; // 1064 :  63 - 0x3f -- Background 0x85
      11'h429: dout  = 8'b00011111; // 1065 :  31 - 0x1f
      11'h42A: dout  = 8'b00011111; // 1066 :  31 - 0x1f
      11'h42B: dout  = 8'b00001111; // 1067 :  15 - 0xf
      11'h42C: dout  = 8'b00000111; // 1068 :   7 - 0x7
      11'h42D: dout  = 8'b00000000; // 1069 :   0 - 0x0
      11'h42E: dout  = 8'b00000000; // 1070 :   0 - 0x0
      11'h42F: dout  = 8'b00000000; // 1071 :   0 - 0x0
      11'h430: dout  = 8'b00000000; // 1072 :   0 - 0x0 -- Background 0x86
      11'h431: dout  = 8'b00000000; // 1073 :   0 - 0x0
      11'h432: dout  = 8'b11000000; // 1074 : 192 - 0xc0
      11'h433: dout  = 8'b11100000; // 1075 : 224 - 0xe0
      11'h434: dout  = 8'b11110000; // 1076 : 240 - 0xf0
      11'h435: dout  = 8'b11110000; // 1077 : 240 - 0xf0
      11'h436: dout  = 8'b11110000; // 1078 : 240 - 0xf0
      11'h437: dout  = 8'b11111000; // 1079 : 248 - 0xf8
      11'h438: dout  = 8'b11111001; // 1080 : 249 - 0xf9 -- Background 0x87
      11'h439: dout  = 8'b11111111; // 1081 : 255 - 0xff
      11'h43A: dout  = 8'b11111111; // 1082 : 255 - 0xff
      11'h43B: dout  = 8'b11111111; // 1083 : 255 - 0xff
      11'h43C: dout  = 8'b11111111; // 1084 : 255 - 0xff
      11'h43D: dout  = 8'b00001110; // 1085 :  14 - 0xe
      11'h43E: dout  = 8'b00000010; // 1086 :   2 - 0x2
      11'h43F: dout  = 8'b00010100; // 1087 :  20 - 0x14
      11'h440: dout  = 8'b10000000; // 1088 : 128 - 0x80 -- Background 0x88
      11'h441: dout  = 8'b10100000; // 1089 : 160 - 0xa0
      11'h442: dout  = 8'b00100000; // 1090 :  32 - 0x20
      11'h443: dout  = 8'b00100000; // 1091 :  32 - 0x20
      11'h444: dout  = 8'b10100000; // 1092 : 160 - 0xa0
      11'h445: dout  = 8'b10000000; // 1093 : 128 - 0x80
      11'h446: dout  = 8'b00000000; // 1094 :   0 - 0x0
      11'h447: dout  = 8'b00000000; // 1095 :   0 - 0x0
      11'h448: dout  = 8'b00000001; // 1096 :   1 - 0x1 -- Background 0x89
      11'h449: dout  = 8'b00000101; // 1097 :   5 - 0x5
      11'h44A: dout  = 8'b00000100; // 1098 :   4 - 0x4
      11'h44B: dout  = 8'b00000100; // 1099 :   4 - 0x4
      11'h44C: dout  = 8'b00000101; // 1100 :   5 - 0x5
      11'h44D: dout  = 8'b00000001; // 1101 :   1 - 0x1
      11'h44E: dout  = 8'b00000000; // 1102 :   0 - 0x0
      11'h44F: dout  = 8'b00000000; // 1103 :   0 - 0x0
      11'h450: dout  = 8'b00000000; // 1104 :   0 - 0x0 -- Background 0x8a
      11'h451: dout  = 8'b00000000; // 1105 :   0 - 0x0
      11'h452: dout  = 8'b00000011; // 1106 :   3 - 0x3
      11'h453: dout  = 8'b00000111; // 1107 :   7 - 0x7
      11'h454: dout  = 8'b00001111; // 1108 :  15 - 0xf
      11'h455: dout  = 8'b00001111; // 1109 :  15 - 0xf
      11'h456: dout  = 8'b00001111; // 1110 :  15 - 0xf
      11'h457: dout  = 8'b00001111; // 1111 :  15 - 0xf
      11'h458: dout  = 8'b10011111; // 1112 : 159 - 0x9f -- Background 0x8b
      11'h459: dout  = 8'b11111111; // 1113 : 255 - 0xff
      11'h45A: dout  = 8'b11111111; // 1114 : 255 - 0xff
      11'h45B: dout  = 8'b11111111; // 1115 : 255 - 0xff
      11'h45C: dout  = 8'b11111111; // 1116 : 255 - 0xff
      11'h45D: dout  = 8'b01110000; // 1117 : 112 - 0x70
      11'h45E: dout  = 8'b01000000; // 1118 :  64 - 0x40
      11'h45F: dout  = 8'b00101000; // 1119 :  40 - 0x28
      11'h460: dout  = 8'b00000000; // 1120 :   0 - 0x0 -- Background 0x8c
      11'h461: dout  = 8'b00000000; // 1121 :   0 - 0x0
      11'h462: dout  = 8'b00000000; // 1122 :   0 - 0x0
      11'h463: dout  = 8'b00000000; // 1123 :   0 - 0x0
      11'h464: dout  = 8'b00000000; // 1124 :   0 - 0x0
      11'h465: dout  = 8'b00000000; // 1125 :   0 - 0x0
      11'h466: dout  = 8'b00000001; // 1126 :   1 - 0x1
      11'h467: dout  = 8'b00000011; // 1127 :   3 - 0x3
      11'h468: dout  = 8'b00000111; // 1128 :   7 - 0x7 -- Background 0x8d
      11'h469: dout  = 8'b00000111; // 1129 :   7 - 0x7
      11'h46A: dout  = 8'b00001111; // 1130 :  15 - 0xf
      11'h46B: dout  = 8'b00001111; // 1131 :  15 - 0xf
      11'h46C: dout  = 8'b00001111; // 1132 :  15 - 0xf
      11'h46D: dout  = 8'b00001111; // 1133 :  15 - 0xf
      11'h46E: dout  = 8'b00011111; // 1134 :  31 - 0x1f
      11'h46F: dout  = 8'b00011111; // 1135 :  31 - 0x1f
      11'h470: dout  = 8'b01111111; // 1136 : 127 - 0x7f -- Background 0x8e
      11'h471: dout  = 8'b11111111; // 1137 : 255 - 0xff
      11'h472: dout  = 8'b11111111; // 1138 : 255 - 0xff
      11'h473: dout  = 8'b11111111; // 1139 : 255 - 0xff
      11'h474: dout  = 8'b11111111; // 1140 : 255 - 0xff
      11'h475: dout  = 8'b11111111; // 1141 : 255 - 0xff
      11'h476: dout  = 8'b11111111; // 1142 : 255 - 0xff
      11'h477: dout  = 8'b11111111; // 1143 : 255 - 0xff
      11'h478: dout  = 8'b11111100; // 1144 : 252 - 0xfc -- Background 0x8f
      11'h479: dout  = 8'b11111000; // 1145 : 248 - 0xf8
      11'h47A: dout  = 8'b11111000; // 1146 : 248 - 0xf8
      11'h47B: dout  = 8'b11110000; // 1147 : 240 - 0xf0
      11'h47C: dout  = 8'b11100000; // 1148 : 224 - 0xe0
      11'h47D: dout  = 8'b00000000; // 1149 :   0 - 0x0
      11'h47E: dout  = 8'b00000000; // 1150 :   0 - 0x0
      11'h47F: dout  = 8'b00000000; // 1151 :   0 - 0x0
      11'h480: dout  = 8'b00000000; // 1152 :   0 - 0x0 -- Background 0x90
      11'h481: dout  = 8'b00000000; // 1153 :   0 - 0x0
      11'h482: dout  = 8'b00000000; // 1154 :   0 - 0x0
      11'h483: dout  = 8'b00000000; // 1155 :   0 - 0x0
      11'h484: dout  = 8'b00000111; // 1156 :   7 - 0x7
      11'h485: dout  = 8'b01111111; // 1157 : 127 - 0x7f
      11'h486: dout  = 8'b11111111; // 1158 : 255 - 0xff
      11'h487: dout  = 8'b11001111; // 1159 : 207 - 0xcf
      11'h488: dout  = 8'b11011111; // 1160 : 223 - 0xdf -- Background 0x91
      11'h489: dout  = 8'b11011111; // 1161 : 223 - 0xdf
      11'h48A: dout  = 8'b11011111; // 1162 : 223 - 0xdf
      11'h48B: dout  = 8'b11011111; // 1163 : 223 - 0xdf
      11'h48C: dout  = 8'b11011111; // 1164 : 223 - 0xdf
      11'h48D: dout  = 8'b11001111; // 1165 : 207 - 0xcf
      11'h48E: dout  = 8'b11101111; // 1166 : 239 - 0xef
      11'h48F: dout  = 8'b11100111; // 1167 : 231 - 0xe7
      11'h490: dout  = 8'b11110011; // 1168 : 243 - 0xf3 -- Background 0x92
      11'h491: dout  = 8'b11111001; // 1169 : 249 - 0xf9
      11'h492: dout  = 8'b11111100; // 1170 : 252 - 0xfc
      11'h493: dout  = 8'b11111100; // 1171 : 252 - 0xfc
      11'h494: dout  = 8'b11111100; // 1172 : 252 - 0xfc
      11'h495: dout  = 8'b11110000; // 1173 : 240 - 0xf0
      11'h496: dout  = 8'b11000000; // 1174 : 192 - 0xc0
      11'h497: dout  = 8'b00000000; // 1175 :   0 - 0x0
      11'h498: dout  = 8'b00000011; // 1176 :   3 - 0x3 -- Background 0x93
      11'h499: dout  = 8'b00001111; // 1177 :  15 - 0xf
      11'h49A: dout  = 8'b00111111; // 1178 :  63 - 0x3f
      11'h49B: dout  = 8'b00001111; // 1179 :  15 - 0xf
      11'h49C: dout  = 8'b00001111; // 1180 :  15 - 0xf
      11'h49D: dout  = 8'b00011001; // 1181 :  25 - 0x19
      11'h49E: dout  = 8'b00010000; // 1182 :  16 - 0x10
      11'h49F: dout  = 8'b00000000; // 1183 :   0 - 0x0
      11'h4A0: dout  = 8'b00011111; // 1184 :  31 - 0x1f -- Background 0x94
      11'h4A1: dout  = 8'b01111111; // 1185 : 127 - 0x7f
      11'h4A2: dout  = 8'b11111110; // 1186 : 254 - 0xfe
      11'h4A3: dout  = 8'b11111000; // 1187 : 248 - 0xf8
      11'h4A4: dout  = 8'b11110000; // 1188 : 240 - 0xf0
      11'h4A5: dout  = 8'b10011000; // 1189 : 152 - 0x98
      11'h4A6: dout  = 8'b00001100; // 1190 :  12 - 0xc
      11'h4A7: dout  = 8'b00001110; // 1191 :  14 - 0xe
      11'h4A8: dout  = 8'b11011111; // 1192 : 223 - 0xdf -- Background 0x95
      11'h4A9: dout  = 8'b11001110; // 1193 : 206 - 0xce
      11'h4AA: dout  = 8'b11100100; // 1194 : 228 - 0xe4
      11'h4AB: dout  = 8'b11110000; // 1195 : 240 - 0xf0
      11'h4AC: dout  = 8'b11111000; // 1196 : 248 - 0xf8
      11'h4AD: dout  = 8'b11111000; // 1197 : 248 - 0xf8
      11'h4AE: dout  = 8'b11111100; // 1198 : 252 - 0xfc
      11'h4AF: dout  = 8'b11111110; // 1199 : 254 - 0xfe
      11'h4B0: dout  = 8'b11111111; // 1200 : 255 - 0xff -- Background 0x96
      11'h4B1: dout  = 8'b11111111; // 1201 : 255 - 0xff
      11'h4B2: dout  = 8'b11111111; // 1202 : 255 - 0xff
      11'h4B3: dout  = 8'b11111111; // 1203 : 255 - 0xff
      11'h4B4: dout  = 8'b01111111; // 1204 : 127 - 0x7f
      11'h4B5: dout  = 8'b10111111; // 1205 : 191 - 0xbf
      11'h4B6: dout  = 8'b00011111; // 1206 :  31 - 0x1f
      11'h4B7: dout  = 8'b01101111; // 1207 : 111 - 0x6f
      11'h4B8: dout  = 8'b11110111; // 1208 : 247 - 0xf7 -- Background 0x97
      11'h4B9: dout  = 8'b11110011; // 1209 : 243 - 0xf3
      11'h4BA: dout  = 8'b11111001; // 1210 : 249 - 0xf9
      11'h4BB: dout  = 8'b11111000; // 1211 : 248 - 0xf8
      11'h4BC: dout  = 8'b11110000; // 1212 : 240 - 0xf0
      11'h4BD: dout  = 8'b10110100; // 1213 : 180 - 0xb4
      11'h4BE: dout  = 8'b00001010; // 1214 :  10 - 0xa
      11'h4BF: dout  = 8'b00000010; // 1215 :   2 - 0x2
      11'h4C0: dout  = 8'b10000000; // 1216 : 128 - 0x80 -- Background 0x98
      11'h4C1: dout  = 8'b11000000; // 1217 : 192 - 0xc0
      11'h4C2: dout  = 8'b00000000; // 1218 :   0 - 0x0
      11'h4C3: dout  = 8'b00000000; // 1219 :   0 - 0x0
      11'h4C4: dout  = 8'b11000000; // 1220 : 192 - 0xc0
      11'h4C5: dout  = 8'b10011000; // 1221 : 152 - 0x98
      11'h4C6: dout  = 8'b00000000; // 1222 :   0 - 0x0
      11'h4C7: dout  = 8'b00000000; // 1223 :   0 - 0x0
      11'h4C8: dout  = 8'b00000000; // 1224 :   0 - 0x0 -- Background 0x99
      11'h4C9: dout  = 8'b00000000; // 1225 :   0 - 0x0
      11'h4CA: dout  = 8'b00111110; // 1226 :  62 - 0x3e
      11'h4CB: dout  = 8'b01000000; // 1227 :  64 - 0x40
      11'h4CC: dout  = 8'b10000000; // 1228 : 128 - 0x80
      11'h4CD: dout  = 8'b00000000; // 1229 :   0 - 0x0
      11'h4CE: dout  = 8'b00000000; // 1230 :   0 - 0x0
      11'h4CF: dout  = 8'b00000000; // 1231 :   0 - 0x0
      11'h4D0: dout  = 8'b00000000; // 1232 :   0 - 0x0 -- Background 0x9a
      11'h4D1: dout  = 8'b00000000; // 1233 :   0 - 0x0
      11'h4D2: dout  = 8'b10000000; // 1234 : 128 - 0x80
      11'h4D3: dout  = 8'b10000000; // 1235 : 128 - 0x80
      11'h4D4: dout  = 8'b11000000; // 1236 : 192 - 0xc0
      11'h4D5: dout  = 8'b11100000; // 1237 : 224 - 0xe0
      11'h4D6: dout  = 8'b11100000; // 1238 : 224 - 0xe0
      11'h4D7: dout  = 8'b11110000; // 1239 : 240 - 0xf0
      11'h4D8: dout  = 8'b11110000; // 1240 : 240 - 0xf0 -- Background 0x9b
      11'h4D9: dout  = 8'b11100000; // 1241 : 224 - 0xe0
      11'h4DA: dout  = 8'b11110000; // 1242 : 240 - 0xf0
      11'h4DB: dout  = 8'b11100000; // 1243 : 224 - 0xe0
      11'h4DC: dout  = 8'b10000000; // 1244 : 128 - 0x80
      11'h4DD: dout  = 8'b00001000; // 1245 :   8 - 0x8
      11'h4DE: dout  = 8'b00000100; // 1246 :   4 - 0x4
      11'h4DF: dout  = 8'b00000000; // 1247 :   0 - 0x0
      11'h4E0: dout  = 8'b00000000; // 1248 :   0 - 0x0 -- Background 0x9c
      11'h4E1: dout  = 8'b00000000; // 1249 :   0 - 0x0
      11'h4E2: dout  = 8'b00000001; // 1250 :   1 - 0x1
      11'h4E3: dout  = 8'b00000011; // 1251 :   3 - 0x3
      11'h4E4: dout  = 8'b00000011; // 1252 :   3 - 0x3
      11'h4E5: dout  = 8'b00000011; // 1253 :   3 - 0x3
      11'h4E6: dout  = 8'b00000111; // 1254 :   7 - 0x7
      11'h4E7: dout  = 8'b00000111; // 1255 :   7 - 0x7
      11'h4E8: dout  = 8'b00000111; // 1256 :   7 - 0x7 -- Background 0x9d
      11'h4E9: dout  = 8'b00000011; // 1257 :   3 - 0x3
      11'h4EA: dout  = 8'b00000011; // 1258 :   3 - 0x3
      11'h4EB: dout  = 8'b00000011; // 1259 :   3 - 0x3
      11'h4EC: dout  = 8'b00000011; // 1260 :   3 - 0x3
      11'h4ED: dout  = 8'b00000011; // 1261 :   3 - 0x3
      11'h4EE: dout  = 8'b00000011; // 1262 :   3 - 0x3
      11'h4EF: dout  = 8'b00000001; // 1263 :   1 - 0x1
      11'h4F0: dout  = 8'b00000000; // 1264 :   0 - 0x0 -- Background 0x9e
      11'h4F1: dout  = 8'b00000000; // 1265 :   0 - 0x0
      11'h4F2: dout  = 8'b00000000; // 1266 :   0 - 0x0
      11'h4F3: dout  = 8'b00000000; // 1267 :   0 - 0x0
      11'h4F4: dout  = 8'b00000000; // 1268 :   0 - 0x0
      11'h4F5: dout  = 8'b00000001; // 1269 :   1 - 0x1
      11'h4F6: dout  = 8'b00000010; // 1270 :   2 - 0x2
      11'h4F7: dout  = 8'b00000100; // 1271 :   4 - 0x4
      11'h4F8: dout  = 8'b00000000; // 1272 :   0 - 0x0 -- Background 0x9f
      11'h4F9: dout  = 8'b00000000; // 1273 :   0 - 0x0
      11'h4FA: dout  = 8'b00000000; // 1274 :   0 - 0x0
      11'h4FB: dout  = 8'b00000000; // 1275 :   0 - 0x0
      11'h4FC: dout  = 8'b00000000; // 1276 :   0 - 0x0
      11'h4FD: dout  = 8'b00000000; // 1277 :   0 - 0x0
      11'h4FE: dout  = 8'b00011100; // 1278 :  28 - 0x1c
      11'h4FF: dout  = 8'b00111011; // 1279 :  59 - 0x3b
      11'h500: dout  = 8'b01111110; // 1280 : 126 - 0x7e -- Background 0xa0
      11'h501: dout  = 8'b11111110; // 1281 : 254 - 0xfe
      11'h502: dout  = 8'b11111111; // 1282 : 255 - 0xff
      11'h503: dout  = 8'b11111111; // 1283 : 255 - 0xff
      11'h504: dout  = 8'b11111111; // 1284 : 255 - 0xff
      11'h505: dout  = 8'b11111111; // 1285 : 255 - 0xff
      11'h506: dout  = 8'b11111101; // 1286 : 253 - 0xfd
      11'h507: dout  = 8'b11111001; // 1287 : 249 - 0xf9
      11'h508: dout  = 8'b11110011; // 1288 : 243 - 0xf3 -- Background 0xa1
      11'h509: dout  = 8'b11110111; // 1289 : 247 - 0xf7
      11'h50A: dout  = 8'b11110110; // 1290 : 246 - 0xf6
      11'h50B: dout  = 8'b11101110; // 1291 : 238 - 0xee
      11'h50C: dout  = 8'b11111101; // 1292 : 253 - 0xfd
      11'h50D: dout  = 8'b11111100; // 1293 : 252 - 0xfc
      11'h50E: dout  = 8'b11111000; // 1294 : 248 - 0xf8
      11'h50F: dout  = 8'b11100001; // 1295 : 225 - 0xe1
      11'h510: dout  = 8'b11010011; // 1296 : 211 - 0xd3 -- Background 0xa2
      11'h511: dout  = 8'b11001011; // 1297 : 203 - 0xcb
      11'h512: dout  = 8'b11000011; // 1298 : 195 - 0xc3
      11'h513: dout  = 8'b11100001; // 1299 : 225 - 0xe1
      11'h514: dout  = 8'b11111001; // 1300 : 249 - 0xf9
      11'h515: dout  = 8'b00111001; // 1301 :  57 - 0x39
      11'h516: dout  = 8'b01000010; // 1302 :  66 - 0x42
      11'h517: dout  = 8'b00000000; // 1303 :   0 - 0x0
      11'h518: dout  = 8'b00000111; // 1304 :   7 - 0x7 -- Background 0xa3
      11'h519: dout  = 8'b00001111; // 1305 :  15 - 0xf
      11'h51A: dout  = 8'b00011001; // 1306 :  25 - 0x19
      11'h51B: dout  = 8'b00110000; // 1307 :  48 - 0x30
      11'h51C: dout  = 8'b01100011; // 1308 :  99 - 0x63
      11'h51D: dout  = 8'b01110010; // 1309 : 114 - 0x72
      11'h51E: dout  = 8'b01110000; // 1310 : 112 - 0x70
      11'h51F: dout  = 8'b00000001; // 1311 :   1 - 0x1
      11'h520: dout  = 8'b00000000; // 1312 :   0 - 0x0 -- Background 0xa4
      11'h521: dout  = 8'b00011111; // 1313 :  31 - 0x1f
      11'h522: dout  = 8'b00100000; // 1314 :  32 - 0x20
      11'h523: dout  = 8'b11000000; // 1315 : 192 - 0xc0
      11'h524: dout  = 8'b11000000; // 1316 : 192 - 0xc0
      11'h525: dout  = 8'b11110000; // 1317 : 240 - 0xf0
      11'h526: dout  = 8'b11111111; // 1318 : 255 - 0xff
      11'h527: dout  = 8'b11111111; // 1319 : 255 - 0xff
      11'h528: dout  = 8'b10101011; // 1320 : 171 - 0xab -- Background 0xa5
      11'h529: dout  = 8'b11000001; // 1321 : 193 - 0xc1
      11'h52A: dout  = 8'b10000001; // 1322 : 129 - 0x81
      11'h52B: dout  = 8'b10010001; // 1323 : 145 - 0x91
      11'h52C: dout  = 8'b10000010; // 1324 : 130 - 0x82
      11'h52D: dout  = 8'b11111100; // 1325 : 252 - 0xfc
      11'h52E: dout  = 8'b11100000; // 1326 : 224 - 0xe0
      11'h52F: dout  = 8'b11001110; // 1327 : 206 - 0xce
      11'h530: dout  = 8'b11100101; // 1328 : 229 - 0xe5 -- Background 0xa6
      11'h531: dout  = 8'b11011010; // 1329 : 218 - 0xda
      11'h532: dout  = 8'b11110000; // 1330 : 240 - 0xf0
      11'h533: dout  = 8'b11100000; // 1331 : 224 - 0xe0
      11'h534: dout  = 8'b11000000; // 1332 : 192 - 0xc0
      11'h535: dout  = 8'b00000000; // 1333 :   0 - 0x0
      11'h536: dout  = 8'b00000000; // 1334 :   0 - 0x0
      11'h537: dout  = 8'b00000000; // 1335 :   0 - 0x0
      11'h538: dout  = 8'b11110000; // 1336 : 240 - 0xf0 -- Background 0xa7
      11'h539: dout  = 8'b11111000; // 1337 : 248 - 0xf8
      11'h53A: dout  = 8'b11001100; // 1338 : 204 - 0xcc
      11'h53B: dout  = 8'b10000110; // 1339 : 134 - 0x86
      11'h53C: dout  = 8'b01100010; // 1340 :  98 - 0x62
      11'h53D: dout  = 8'b00100110; // 1341 :  38 - 0x26
      11'h53E: dout  = 8'b00000110; // 1342 :   6 - 0x6
      11'h53F: dout  = 8'b11000000; // 1343 : 192 - 0xc0
      11'h540: dout  = 8'b00000000; // 1344 :   0 - 0x0 -- Background 0xa8
      11'h541: dout  = 8'b11111100; // 1345 : 252 - 0xfc
      11'h542: dout  = 8'b00000110; // 1346 :   6 - 0x6
      11'h543: dout  = 8'b00000011; // 1347 :   3 - 0x3
      11'h544: dout  = 8'b00000001; // 1348 :   1 - 0x1
      11'h545: dout  = 8'b00000111; // 1349 :   7 - 0x7
      11'h546: dout  = 8'b11111111; // 1350 : 255 - 0xff
      11'h547: dout  = 8'b11111111; // 1351 : 255 - 0xff
      11'h548: dout  = 8'b11010101; // 1352 : 213 - 0xd5 -- Background 0xa9
      11'h549: dout  = 8'b10000011; // 1353 : 131 - 0x83
      11'h54A: dout  = 8'b10000001; // 1354 : 129 - 0x81
      11'h54B: dout  = 8'b10001001; // 1355 : 137 - 0x89
      11'h54C: dout  = 8'b01000001; // 1356 :  65 - 0x41
      11'h54D: dout  = 8'b00111111; // 1357 :  63 - 0x3f
      11'h54E: dout  = 8'b00000111; // 1358 :   7 - 0x7
      11'h54F: dout  = 8'b11010011; // 1359 : 211 - 0xd3
      11'h550: dout  = 8'b01101111; // 1360 : 111 - 0x6f -- Background 0xaa
      11'h551: dout  = 8'b11011011; // 1361 : 219 - 0xdb
      11'h552: dout  = 8'b00001111; // 1362 :  15 - 0xf
      11'h553: dout  = 8'b00000111; // 1363 :   7 - 0x7
      11'h554: dout  = 8'b00000011; // 1364 :   3 - 0x3
      11'h555: dout  = 8'b00000000; // 1365 :   0 - 0x0
      11'h556: dout  = 8'b00000000; // 1366 :   0 - 0x0
      11'h557: dout  = 8'b00000000; // 1367 :   0 - 0x0
      11'h558: dout  = 8'b00000000; // 1368 :   0 - 0x0 -- Background 0xab
      11'h559: dout  = 8'b00000000; // 1369 :   0 - 0x0
      11'h55A: dout  = 8'b00000000; // 1370 :   0 - 0x0
      11'h55B: dout  = 8'b00000000; // 1371 :   0 - 0x0
      11'h55C: dout  = 8'b00000000; // 1372 :   0 - 0x0
      11'h55D: dout  = 8'b00000000; // 1373 :   0 - 0x0
      11'h55E: dout  = 8'b00111000; // 1374 :  56 - 0x38
      11'h55F: dout  = 8'b11011100; // 1375 : 220 - 0xdc
      11'h560: dout  = 8'b01111110; // 1376 : 126 - 0x7e -- Background 0xac
      11'h561: dout  = 8'b01111111; // 1377 : 127 - 0x7f
      11'h562: dout  = 8'b01111111; // 1378 : 127 - 0x7f
      11'h563: dout  = 8'b11111111; // 1379 : 255 - 0xff
      11'h564: dout  = 8'b11111111; // 1380 : 255 - 0xff
      11'h565: dout  = 8'b11111111; // 1381 : 255 - 0xff
      11'h566: dout  = 8'b10111111; // 1382 : 191 - 0xbf
      11'h567: dout  = 8'b10011111; // 1383 : 159 - 0x9f
      11'h568: dout  = 8'b11001111; // 1384 : 207 - 0xcf -- Background 0xad
      11'h569: dout  = 8'b11101111; // 1385 : 239 - 0xef
      11'h56A: dout  = 8'b01101111; // 1386 : 111 - 0x6f
      11'h56B: dout  = 8'b01110111; // 1387 : 119 - 0x77
      11'h56C: dout  = 8'b10111111; // 1388 : 191 - 0xbf
      11'h56D: dout  = 8'b00111111; // 1389 :  63 - 0x3f
      11'h56E: dout  = 8'b00011111; // 1390 :  31 - 0x1f
      11'h56F: dout  = 8'b10000111; // 1391 : 135 - 0x87
      11'h570: dout  = 8'b11001011; // 1392 : 203 - 0xcb -- Background 0xae
      11'h571: dout  = 8'b11010011; // 1393 : 211 - 0xd3
      11'h572: dout  = 8'b11000011; // 1394 : 195 - 0xc3
      11'h573: dout  = 8'b10000111; // 1395 : 135 - 0x87
      11'h574: dout  = 8'b10011111; // 1396 : 159 - 0x9f
      11'h575: dout  = 8'b10011100; // 1397 : 156 - 0x9c
      11'h576: dout  = 8'b01000010; // 1398 :  66 - 0x42
      11'h577: dout  = 8'b00000000; // 1399 :   0 - 0x0
      11'h578: dout  = 8'b00000000; // 1400 :   0 - 0x0 -- Background 0xaf
      11'h579: dout  = 8'b00000000; // 1401 :   0 - 0x0
      11'h57A: dout  = 8'b10000000; // 1402 : 128 - 0x80
      11'h57B: dout  = 8'b11000000; // 1403 : 192 - 0xc0
      11'h57C: dout  = 8'b11000000; // 1404 : 192 - 0xc0
      11'h57D: dout  = 8'b11000000; // 1405 : 192 - 0xc0
      11'h57E: dout  = 8'b11100000; // 1406 : 224 - 0xe0
      11'h57F: dout  = 8'b11100000; // 1407 : 224 - 0xe0
      11'h580: dout  = 8'b11100000; // 1408 : 224 - 0xe0 -- Background 0xb0
      11'h581: dout  = 8'b11000000; // 1409 : 192 - 0xc0
      11'h582: dout  = 8'b11000000; // 1410 : 192 - 0xc0
      11'h583: dout  = 8'b11000000; // 1411 : 192 - 0xc0
      11'h584: dout  = 8'b11000000; // 1412 : 192 - 0xc0
      11'h585: dout  = 8'b11000000; // 1413 : 192 - 0xc0
      11'h586: dout  = 8'b11000000; // 1414 : 192 - 0xc0
      11'h587: dout  = 8'b10000000; // 1415 : 128 - 0x80
      11'h588: dout  = 8'b00000000; // 1416 :   0 - 0x0 -- Background 0xb1
      11'h589: dout  = 8'b00000000; // 1417 :   0 - 0x0
      11'h58A: dout  = 8'b00000000; // 1418 :   0 - 0x0
      11'h58B: dout  = 8'b00000000; // 1419 :   0 - 0x0
      11'h58C: dout  = 8'b00000000; // 1420 :   0 - 0x0
      11'h58D: dout  = 8'b10000000; // 1421 : 128 - 0x80
      11'h58E: dout  = 8'b01000000; // 1422 :  64 - 0x40
      11'h58F: dout  = 8'b00100000; // 1423 :  32 - 0x20
      11'h590: dout  = 8'b00000000; // 1424 :   0 - 0x0 -- Background 0xb2
      11'h591: dout  = 8'b00000000; // 1425 :   0 - 0x0
      11'h592: dout  = 8'b00000000; // 1426 :   0 - 0x0
      11'h593: dout  = 8'b00000001; // 1427 :   1 - 0x1
      11'h594: dout  = 8'b00000011; // 1428 :   3 - 0x3
      11'h595: dout  = 8'b00000111; // 1429 :   7 - 0x7
      11'h596: dout  = 8'b00000111; // 1430 :   7 - 0x7
      11'h597: dout  = 8'b00000111; // 1431 :   7 - 0x7
      11'h598: dout  = 8'b00000011; // 1432 :   3 - 0x3 -- Background 0xb3
      11'h599: dout  = 8'b00000001; // 1433 :   1 - 0x1
      11'h59A: dout  = 8'b00000000; // 1434 :   0 - 0x0
      11'h59B: dout  = 8'b00000000; // 1435 :   0 - 0x0
      11'h59C: dout  = 8'b00000000; // 1436 :   0 - 0x0
      11'h59D: dout  = 8'b00000000; // 1437 :   0 - 0x0
      11'h59E: dout  = 8'b00000001; // 1438 :   1 - 0x1
      11'h59F: dout  = 8'b00000001; // 1439 :   1 - 0x1
      11'h5A0: dout  = 8'b00000001; // 1440 :   1 - 0x1 -- Background 0xb4
      11'h5A1: dout  = 8'b00000001; // 1441 :   1 - 0x1
      11'h5A2: dout  = 8'b00000111; // 1442 :   7 - 0x7
      11'h5A3: dout  = 8'b00000011; // 1443 :   3 - 0x3
      11'h5A4: dout  = 8'b00000100; // 1444 :   4 - 0x4
      11'h5A5: dout  = 8'b00000000; // 1445 :   0 - 0x0
      11'h5A6: dout  = 8'b00000000; // 1446 :   0 - 0x0
      11'h5A7: dout  = 8'b00000000; // 1447 :   0 - 0x0
      11'h5A8: dout  = 8'b00000000; // 1448 :   0 - 0x0 -- Background 0xb5
      11'h5A9: dout  = 8'b00000000; // 1449 :   0 - 0x0
      11'h5AA: dout  = 8'b00000000; // 1450 :   0 - 0x0
      11'h5AB: dout  = 8'b00000000; // 1451 :   0 - 0x0
      11'h5AC: dout  = 8'b00000000; // 1452 :   0 - 0x0
      11'h5AD: dout  = 8'b00000000; // 1453 :   0 - 0x0
      11'h5AE: dout  = 8'b00000000; // 1454 :   0 - 0x0
      11'h5AF: dout  = 8'b00000111; // 1455 :   7 - 0x7
      11'h5B0: dout  = 8'b00001110; // 1456 :  14 - 0xe -- Background 0xb6
      11'h5B1: dout  = 8'b00111110; // 1457 :  62 - 0x3e
      11'h5B2: dout  = 8'b01111111; // 1458 : 127 - 0x7f
      11'h5B3: dout  = 8'b11111111; // 1459 : 255 - 0xff
      11'h5B4: dout  = 8'b11111111; // 1460 : 255 - 0xff
      11'h5B5: dout  = 8'b11101111; // 1461 : 239 - 0xef
      11'h5B6: dout  = 8'b11110111; // 1462 : 247 - 0xf7
      11'h5B7: dout  = 8'b11111000; // 1463 : 248 - 0xf8
      11'h5B8: dout  = 8'b11111111; // 1464 : 255 - 0xff -- Background 0xb7
      11'h5B9: dout  = 8'b11111111; // 1465 : 255 - 0xff
      11'h5BA: dout  = 8'b11111111; // 1466 : 255 - 0xff
      11'h5BB: dout  = 8'b00011111; // 1467 :  31 - 0x1f
      11'h5BC: dout  = 8'b00011111; // 1468 :  31 - 0x1f
      11'h5BD: dout  = 8'b01111111; // 1469 : 127 - 0x7f
      11'h5BE: dout  = 8'b11111111; // 1470 : 255 - 0xff
      11'h5BF: dout  = 8'b11111110; // 1471 : 254 - 0xfe
      11'h5C0: dout  = 8'b11111111; // 1472 : 255 - 0xff -- Background 0xb8
      11'h5C1: dout  = 8'b11111111; // 1473 : 255 - 0xff
      11'h5C2: dout  = 8'b11111111; // 1474 : 255 - 0xff
      11'h5C3: dout  = 8'b11111100; // 1475 : 252 - 0xfc
      11'h5C4: dout  = 8'b11111000; // 1476 : 248 - 0xf8
      11'h5C5: dout  = 8'b10000000; // 1477 : 128 - 0x80
      11'h5C6: dout  = 8'b00000000; // 1478 :   0 - 0x0
      11'h5C7: dout  = 8'b00000000; // 1479 :   0 - 0x0
      11'h5C8: dout  = 8'b00110000; // 1480 :  48 - 0x30 -- Background 0xb9
      11'h5C9: dout  = 8'b01111111; // 1481 : 127 - 0x7f
      11'h5CA: dout  = 8'b01111111; // 1482 : 127 - 0x7f
      11'h5CB: dout  = 8'b00111111; // 1483 :  63 - 0x3f
      11'h5CC: dout  = 8'b10000111; // 1484 : 135 - 0x87
      11'h5CD: dout  = 8'b11110000; // 1485 : 240 - 0xf0
      11'h5CE: dout  = 8'b11111111; // 1486 : 255 - 0xff
      11'h5CF: dout  = 8'b11111111; // 1487 : 255 - 0xff
      11'h5D0: dout  = 8'b11100101; // 1488 : 229 - 0xe5 -- Background 0xba
      11'h5D1: dout  = 8'b11011010; // 1489 : 218 - 0xda
      11'h5D2: dout  = 8'b11000000; // 1490 : 192 - 0xc0
      11'h5D3: dout  = 8'b00000000; // 1491 :   0 - 0x0
      11'h5D4: dout  = 8'b00000000; // 1492 :   0 - 0x0
      11'h5D5: dout  = 8'b00000000; // 1493 :   0 - 0x0
      11'h5D6: dout  = 8'b00000000; // 1494 :   0 - 0x0
      11'h5D7: dout  = 8'b00000000; // 1495 :   0 - 0x0
      11'h5D8: dout  = 8'b00000110; // 1496 :   6 - 0x6 -- Background 0xbb
      11'h5D9: dout  = 8'b11111111; // 1497 : 255 - 0xff
      11'h5DA: dout  = 8'b11111111; // 1498 : 255 - 0xff
      11'h5DB: dout  = 8'b11111110; // 1499 : 254 - 0xfe
      11'h5DC: dout  = 8'b11110001; // 1500 : 241 - 0xf1
      11'h5DD: dout  = 8'b00000111; // 1501 :   7 - 0x7
      11'h5DE: dout  = 8'b11111111; // 1502 : 255 - 0xff
      11'h5DF: dout  = 8'b11111111; // 1503 : 255 - 0xff
      11'h5E0: dout  = 8'b00000000; // 1504 :   0 - 0x0 -- Background 0xbc
      11'h5E1: dout  = 8'b00000001; // 1505 :   1 - 0x1
      11'h5E2: dout  = 8'b00000010; // 1506 :   2 - 0x2
      11'h5E3: dout  = 8'b00000111; // 1507 :   7 - 0x7
      11'h5E4: dout  = 8'b00000000; // 1508 :   0 - 0x0
      11'h5E5: dout  = 8'b00000000; // 1509 :   0 - 0x0
      11'h5E6: dout  = 8'b00100000; // 1510 :  32 - 0x20
      11'h5E7: dout  = 8'b11111111; // 1511 : 255 - 0xff
      11'h5E8: dout  = 8'b01111111; // 1512 : 127 - 0x7f -- Background 0xbd
      11'h5E9: dout  = 8'b01111111; // 1513 : 127 - 0x7f
      11'h5EA: dout  = 8'b01111111; // 1514 : 127 - 0x7f
      11'h5EB: dout  = 8'b11111111; // 1515 : 255 - 0xff
      11'h5EC: dout  = 8'b11111111; // 1516 : 255 - 0xff
      11'h5ED: dout  = 8'b11111111; // 1517 : 255 - 0xff
      11'h5EE: dout  = 8'b11111111; // 1518 : 255 - 0xff
      11'h5EF: dout  = 8'b11111110; // 1519 : 254 - 0xfe
      11'h5F0: dout  = 8'b11111100; // 1520 : 252 - 0xfc -- Background 0xbe
      11'h5F1: dout  = 8'b10111000; // 1521 : 184 - 0xb8
      11'h5F2: dout  = 8'b01111000; // 1522 : 120 - 0x78
      11'h5F3: dout  = 8'b01111000; // 1523 : 120 - 0x78
      11'h5F4: dout  = 8'b10110000; // 1524 : 176 - 0xb0
      11'h5F5: dout  = 8'b01111000; // 1525 : 120 - 0x78
      11'h5F6: dout  = 8'b11111100; // 1526 : 252 - 0xfc
      11'h5F7: dout  = 8'b11111110; // 1527 : 254 - 0xfe
      11'h5F8: dout  = 8'b11111111; // 1528 : 255 - 0xff -- Background 0xbf
      11'h5F9: dout  = 8'b11111111; // 1529 : 255 - 0xff
      11'h5FA: dout  = 8'b11111111; // 1530 : 255 - 0xff
      11'h5FB: dout  = 8'b11111111; // 1531 : 255 - 0xff
      11'h5FC: dout  = 8'b11111111; // 1532 : 255 - 0xff
      11'h5FD: dout  = 8'b10011100; // 1533 : 156 - 0x9c
      11'h5FE: dout  = 8'b01000010; // 1534 :  66 - 0x42
      11'h5FF: dout  = 8'b00000000; // 1535 :   0 - 0x0
      11'h600: dout  = 8'b00000000; // 1536 :   0 - 0x0 -- Background 0xc0
      11'h601: dout  = 8'b00000000; // 1537 :   0 - 0x0
      11'h602: dout  = 8'b00100000; // 1538 :  32 - 0x20
      11'h603: dout  = 8'b01000000; // 1539 :  64 - 0x40
      11'h604: dout  = 8'b10001010; // 1540 : 138 - 0x8a
      11'h605: dout  = 8'b00011110; // 1541 :  30 - 0x1e
      11'h606: dout  = 8'b01111110; // 1542 : 126 - 0x7e
      11'h607: dout  = 8'b10111110; // 1543 : 190 - 0xbe
      11'h608: dout  = 8'b11011111; // 1544 : 223 - 0xdf -- Background 0xc1
      11'h609: dout  = 8'b11111111; // 1545 : 255 - 0xff
      11'h60A: dout  = 8'b11111110; // 1546 : 254 - 0xfe
      11'h60B: dout  = 8'b11111100; // 1547 : 252 - 0xfc
      11'h60C: dout  = 8'b11110000; // 1548 : 240 - 0xf0
      11'h60D: dout  = 8'b11100000; // 1549 : 224 - 0xe0
      11'h60E: dout  = 8'b10000000; // 1550 : 128 - 0x80
      11'h60F: dout  = 8'b00000000; // 1551 :   0 - 0x0
      11'h610: dout  = 8'b00000000; // 1552 :   0 - 0x0 -- Background 0xc2
      11'h611: dout  = 8'b00000000; // 1553 :   0 - 0x0
      11'h612: dout  = 8'b00000100; // 1554 :   4 - 0x4
      11'h613: dout  = 8'b00000010; // 1555 :   2 - 0x2
      11'h614: dout  = 8'b01010001; // 1556 :  81 - 0x51
      11'h615: dout  = 8'b01111000; // 1557 : 120 - 0x78
      11'h616: dout  = 8'b01111110; // 1558 : 126 - 0x7e
      11'h617: dout  = 8'b11111101; // 1559 : 253 - 0xfd
      11'h618: dout  = 8'b11111011; // 1560 : 251 - 0xfb -- Background 0xc3
      11'h619: dout  = 8'b11111111; // 1561 : 255 - 0xff
      11'h61A: dout  = 8'b01111111; // 1562 : 127 - 0x7f
      11'h61B: dout  = 8'b00111111; // 1563 :  63 - 0x3f
      11'h61C: dout  = 8'b00001111; // 1564 :  15 - 0xf
      11'h61D: dout  = 8'b00000111; // 1565 :   7 - 0x7
      11'h61E: dout  = 8'b00000001; // 1566 :   1 - 0x1
      11'h61F: dout  = 8'b00000000; // 1567 :   0 - 0x0
      11'h620: dout  = 8'b00000000; // 1568 :   0 - 0x0 -- Background 0xc4
      11'h621: dout  = 8'b10000000; // 1569 : 128 - 0x80
      11'h622: dout  = 8'b01000000; // 1570 :  64 - 0x40
      11'h623: dout  = 8'b11100000; // 1571 : 224 - 0xe0
      11'h624: dout  = 8'b00000000; // 1572 :   0 - 0x0
      11'h625: dout  = 8'b00000000; // 1573 :   0 - 0x0
      11'h626: dout  = 8'b00000100; // 1574 :   4 - 0x4
      11'h627: dout  = 8'b11111111; // 1575 : 255 - 0xff
      11'h628: dout  = 8'b11111110; // 1576 : 254 - 0xfe -- Background 0xc5
      11'h629: dout  = 8'b11111110; // 1577 : 254 - 0xfe
      11'h62A: dout  = 8'b11111110; // 1578 : 254 - 0xfe
      11'h62B: dout  = 8'b11111111; // 1579 : 255 - 0xff
      11'h62C: dout  = 8'b11111111; // 1580 : 255 - 0xff
      11'h62D: dout  = 8'b11111111; // 1581 : 255 - 0xff
      11'h62E: dout  = 8'b11111111; // 1582 : 255 - 0xff
      11'h62F: dout  = 8'b01111111; // 1583 : 127 - 0x7f
      11'h630: dout  = 8'b00111111; // 1584 :  63 - 0x3f -- Background 0xc6
      11'h631: dout  = 8'b00011101; // 1585 :  29 - 0x1d
      11'h632: dout  = 8'b00011110; // 1586 :  30 - 0x1e
      11'h633: dout  = 8'b00011110; // 1587 :  30 - 0x1e
      11'h634: dout  = 8'b00001101; // 1588 :  13 - 0xd
      11'h635: dout  = 8'b00011110; // 1589 :  30 - 0x1e
      11'h636: dout  = 8'b00111111; // 1590 :  63 - 0x3f
      11'h637: dout  = 8'b01111111; // 1591 : 127 - 0x7f
      11'h638: dout  = 8'b11111111; // 1592 : 255 - 0xff -- Background 0xc7
      11'h639: dout  = 8'b11111111; // 1593 : 255 - 0xff
      11'h63A: dout  = 8'b11111111; // 1594 : 255 - 0xff
      11'h63B: dout  = 8'b11111111; // 1595 : 255 - 0xff
      11'h63C: dout  = 8'b11111111; // 1596 : 255 - 0xff
      11'h63D: dout  = 8'b00111001; // 1597 :  57 - 0x39
      11'h63E: dout  = 8'b01000010; // 1598 :  66 - 0x42
      11'h63F: dout  = 8'b00000000; // 1599 :   0 - 0x0
      11'h640: dout  = 8'b01101111; // 1600 : 111 - 0x6f -- Background 0xc8
      11'h641: dout  = 8'b11011011; // 1601 : 219 - 0xdb
      11'h642: dout  = 8'b00000011; // 1602 :   3 - 0x3
      11'h643: dout  = 8'b00000000; // 1603 :   0 - 0x0
      11'h644: dout  = 8'b00000000; // 1604 :   0 - 0x0
      11'h645: dout  = 8'b00000000; // 1605 :   0 - 0x0
      11'h646: dout  = 8'b00000000; // 1606 :   0 - 0x0
      11'h647: dout  = 8'b00000000; // 1607 :   0 - 0x0
      11'h648: dout  = 8'b00000000; // 1608 :   0 - 0x0 -- Background 0xc9
      11'h649: dout  = 8'b00000000; // 1609 :   0 - 0x0
      11'h64A: dout  = 8'b00000000; // 1610 :   0 - 0x0
      11'h64B: dout  = 8'b00000000; // 1611 :   0 - 0x0
      11'h64C: dout  = 8'b00000000; // 1612 :   0 - 0x0
      11'h64D: dout  = 8'b00000000; // 1613 :   0 - 0x0
      11'h64E: dout  = 8'b00000000; // 1614 :   0 - 0x0
      11'h64F: dout  = 8'b11100000; // 1615 : 224 - 0xe0
      11'h650: dout  = 8'b01110000; // 1616 : 112 - 0x70 -- Background 0xca
      11'h651: dout  = 8'b01111100; // 1617 : 124 - 0x7c
      11'h652: dout  = 8'b01111110; // 1618 : 126 - 0x7e
      11'h653: dout  = 8'b11111111; // 1619 : 255 - 0xff
      11'h654: dout  = 8'b11111111; // 1620 : 255 - 0xff
      11'h655: dout  = 8'b11110111; // 1621 : 247 - 0xf7
      11'h656: dout  = 8'b11101111; // 1622 : 239 - 0xef
      11'h657: dout  = 8'b00011111; // 1623 :  31 - 0x1f
      11'h658: dout  = 8'b11111111; // 1624 : 255 - 0xff -- Background 0xcb
      11'h659: dout  = 8'b11111111; // 1625 : 255 - 0xff
      11'h65A: dout  = 8'b11111111; // 1626 : 255 - 0xff
      11'h65B: dout  = 8'b11111000; // 1627 : 248 - 0xf8
      11'h65C: dout  = 8'b11111000; // 1628 : 248 - 0xf8
      11'h65D: dout  = 8'b11111110; // 1629 : 254 - 0xfe
      11'h65E: dout  = 8'b11111111; // 1630 : 255 - 0xff
      11'h65F: dout  = 8'b11111111; // 1631 : 255 - 0xff
      11'h660: dout  = 8'b11111111; // 1632 : 255 - 0xff -- Background 0xcc
      11'h661: dout  = 8'b11111111; // 1633 : 255 - 0xff
      11'h662: dout  = 8'b11111111; // 1634 : 255 - 0xff
      11'h663: dout  = 8'b00111111; // 1635 :  63 - 0x3f
      11'h664: dout  = 8'b00011110; // 1636 :  30 - 0x1e
      11'h665: dout  = 8'b00000001; // 1637 :   1 - 0x1
      11'h666: dout  = 8'b00000000; // 1638 :   0 - 0x0
      11'h667: dout  = 8'b00000000; // 1639 :   0 - 0x0
      11'h668: dout  = 8'b00000000; // 1640 :   0 - 0x0 -- Background 0xcd
      11'h669: dout  = 8'b00000000; // 1641 :   0 - 0x0
      11'h66A: dout  = 8'b00000000; // 1642 :   0 - 0x0
      11'h66B: dout  = 8'b10000000; // 1643 : 128 - 0x80
      11'h66C: dout  = 8'b11000000; // 1644 : 192 - 0xc0
      11'h66D: dout  = 8'b11100000; // 1645 : 224 - 0xe0
      11'h66E: dout  = 8'b11100000; // 1646 : 224 - 0xe0
      11'h66F: dout  = 8'b11100000; // 1647 : 224 - 0xe0
      11'h670: dout  = 8'b11000000; // 1648 : 192 - 0xc0 -- Background 0xce
      11'h671: dout  = 8'b10000000; // 1649 : 128 - 0x80
      11'h672: dout  = 8'b00000000; // 1650 :   0 - 0x0
      11'h673: dout  = 8'b00000000; // 1651 :   0 - 0x0
      11'h674: dout  = 8'b00000000; // 1652 :   0 - 0x0
      11'h675: dout  = 8'b00000000; // 1653 :   0 - 0x0
      11'h676: dout  = 8'b10000000; // 1654 : 128 - 0x80
      11'h677: dout  = 8'b10000000; // 1655 : 128 - 0x80
      11'h678: dout  = 8'b10000000; // 1656 : 128 - 0x80 -- Background 0xcf
      11'h679: dout  = 8'b10000000; // 1657 : 128 - 0x80
      11'h67A: dout  = 8'b11100000; // 1658 : 224 - 0xe0
      11'h67B: dout  = 8'b11000000; // 1659 : 192 - 0xc0
      11'h67C: dout  = 8'b00100000; // 1660 :  32 - 0x20
      11'h67D: dout  = 8'b00000000; // 1661 :   0 - 0x0
      11'h67E: dout  = 8'b00000000; // 1662 :   0 - 0x0
      11'h67F: dout  = 8'b00000000; // 1663 :   0 - 0x0
      11'h680: dout  = 8'b00011111; // 1664 :  31 - 0x1f -- Background 0xd0
      11'h681: dout  = 8'b00000110; // 1665 :   6 - 0x6
      11'h682: dout  = 8'b00000110; // 1666 :   6 - 0x6
      11'h683: dout  = 8'b00000110; // 1667 :   6 - 0x6
      11'h684: dout  = 8'b00000110; // 1668 :   6 - 0x6
      11'h685: dout  = 8'b00000110; // 1669 :   6 - 0x6
      11'h686: dout  = 8'b00000110; // 1670 :   6 - 0x6
      11'h687: dout  = 8'b00000000; // 1671 :   0 - 0x0
      11'h688: dout  = 8'b00111001; // 1672 :  57 - 0x39 -- Background 0xd1
      11'h689: dout  = 8'b01100101; // 1673 : 101 - 0x65
      11'h68A: dout  = 8'b01100101; // 1674 : 101 - 0x65
      11'h68B: dout  = 8'b01100101; // 1675 : 101 - 0x65
      11'h68C: dout  = 8'b01100101; // 1676 : 101 - 0x65
      11'h68D: dout  = 8'b01100101; // 1677 : 101 - 0x65
      11'h68E: dout  = 8'b00111001; // 1678 :  57 - 0x39
      11'h68F: dout  = 8'b00000000; // 1679 :   0 - 0x0
      11'h690: dout  = 8'b11100000; // 1680 : 224 - 0xe0 -- Background 0xd2
      11'h691: dout  = 8'b10110000; // 1681 : 176 - 0xb0
      11'h692: dout  = 8'b10110000; // 1682 : 176 - 0xb0
      11'h693: dout  = 8'b10110110; // 1683 : 182 - 0xb6
      11'h694: dout  = 8'b11100110; // 1684 : 230 - 0xe6
      11'h695: dout  = 8'b10000000; // 1685 : 128 - 0x80
      11'h696: dout  = 8'b10000000; // 1686 : 128 - 0x80
      11'h697: dout  = 8'b00000000; // 1687 :   0 - 0x0
      11'h698: dout  = 8'b00111100; // 1688 :  60 - 0x3c -- Background 0xd3
      11'h699: dout  = 8'b01000010; // 1689 :  66 - 0x42
      11'h69A: dout  = 8'b10011001; // 1690 : 153 - 0x99
      11'h69B: dout  = 8'b10100001; // 1691 : 161 - 0xa1
      11'h69C: dout  = 8'b10100001; // 1692 : 161 - 0xa1
      11'h69D: dout  = 8'b10011001; // 1693 : 153 - 0x99
      11'h69E: dout  = 8'b01000010; // 1694 :  66 - 0x42
      11'h69F: dout  = 8'b00111100; // 1695 :  60 - 0x3c
      11'h6A0: dout  = 8'b00000000; // 1696 :   0 - 0x0 -- Background 0xd4
      11'h6A1: dout  = 8'b00000000; // 1697 :   0 - 0x0
      11'h6A2: dout  = 8'b00000000; // 1698 :   0 - 0x0
      11'h6A3: dout  = 8'b00000011; // 1699 :   3 - 0x3
      11'h6A4: dout  = 8'b00000110; // 1700 :   6 - 0x6
      11'h6A5: dout  = 8'b00000000; // 1701 :   0 - 0x0
      11'h6A6: dout  = 8'b00000001; // 1702 :   1 - 0x1
      11'h6A7: dout  = 8'b00000111; // 1703 :   7 - 0x7
      11'h6A8: dout  = 8'b00001111; // 1704 :  15 - 0xf -- Background 0xd5
      11'h6A9: dout  = 8'b00011111; // 1705 :  31 - 0x1f
      11'h6AA: dout  = 8'b00111111; // 1706 :  63 - 0x3f
      11'h6AB: dout  = 8'b01111111; // 1707 : 127 - 0x7f
      11'h6AC: dout  = 8'b01111111; // 1708 : 127 - 0x7f
      11'h6AD: dout  = 8'b01111111; // 1709 : 127 - 0x7f
      11'h6AE: dout  = 8'b11111111; // 1710 : 255 - 0xff
      11'h6AF: dout  = 8'b01111111; // 1711 : 127 - 0x7f
      11'h6B0: dout  = 8'b00000000; // 1712 :   0 - 0x0 -- Background 0xd6
      11'h6B1: dout  = 8'b00000000; // 1713 :   0 - 0x0
      11'h6B2: dout  = 8'b00000000; // 1714 :   0 - 0x0
      11'h6B3: dout  = 8'b10000000; // 1715 : 128 - 0x80
      11'h6B4: dout  = 8'b00000000; // 1716 :   0 - 0x0
      11'h6B5: dout  = 8'b00000000; // 1717 :   0 - 0x0
      11'h6B6: dout  = 8'b00000000; // 1718 :   0 - 0x0
      11'h6B7: dout  = 8'b10100000; // 1719 : 160 - 0xa0
      11'h6B8: dout  = 8'b11100000; // 1720 : 224 - 0xe0 -- Background 0xd7
      11'h6B9: dout  = 8'b11110000; // 1721 : 240 - 0xf0
      11'h6BA: dout  = 8'b11100000; // 1722 : 224 - 0xe0
      11'h6BB: dout  = 8'b11011101; // 1723 : 221 - 0xdd
      11'h6BC: dout  = 8'b11111010; // 1724 : 250 - 0xfa
      11'h6BD: dout  = 8'b11101011; // 1725 : 235 - 0xeb
      11'h6BE: dout  = 8'b10000000; // 1726 : 128 - 0x80
      11'h6BF: dout  = 8'b00000000; // 1727 :   0 - 0x0
      11'h6C0: dout  = 8'b00000000; // 1728 :   0 - 0x0 -- Background 0xd8
      11'h6C1: dout  = 8'b00000000; // 1729 :   0 - 0x0
      11'h6C2: dout  = 8'b00000000; // 1730 :   0 - 0x0
      11'h6C3: dout  = 8'b00000011; // 1731 :   3 - 0x3
      11'h6C4: dout  = 8'b00000110; // 1732 :   6 - 0x6
      11'h6C5: dout  = 8'b00000000; // 1733 :   0 - 0x0
      11'h6C6: dout  = 8'b00000001; // 1734 :   1 - 0x1
      11'h6C7: dout  = 8'b00000001; // 1735 :   1 - 0x1
      11'h6C8: dout  = 8'b00001011; // 1736 :  11 - 0xb -- Background 0xd9
      11'h6C9: dout  = 8'b00000111; // 1737 :   7 - 0x7
      11'h6CA: dout  = 8'b00000011; // 1738 :   3 - 0x3
      11'h6CB: dout  = 8'b01011101; // 1739 :  93 - 0x5d
      11'h6CC: dout  = 8'b10101111; // 1740 : 175 - 0xaf
      11'h6CD: dout  = 8'b01010011; // 1741 :  83 - 0x53
      11'h6CE: dout  = 8'b00000000; // 1742 :   0 - 0x0
      11'h6CF: dout  = 8'b00000000; // 1743 :   0 - 0x0
      11'h6D0: dout  = 8'b00000000; // 1744 :   0 - 0x0 -- Background 0xda
      11'h6D1: dout  = 8'b00000000; // 1745 :   0 - 0x0
      11'h6D2: dout  = 8'b00000000; // 1746 :   0 - 0x0
      11'h6D3: dout  = 8'b10000000; // 1747 : 128 - 0x80
      11'h6D4: dout  = 8'b00000000; // 1748 :   0 - 0x0
      11'h6D5: dout  = 8'b00000000; // 1749 :   0 - 0x0
      11'h6D6: dout  = 8'b01100000; // 1750 :  96 - 0x60
      11'h6D7: dout  = 8'b11110000; // 1751 : 240 - 0xf0
      11'h6D8: dout  = 8'b11111000; // 1752 : 248 - 0xf8 -- Background 0xdb
      11'h6D9: dout  = 8'b11111100; // 1753 : 252 - 0xfc
      11'h6DA: dout  = 8'b11111100; // 1754 : 252 - 0xfc
      11'h6DB: dout  = 8'b11111110; // 1755 : 254 - 0xfe
      11'h6DC: dout  = 8'b11111110; // 1756 : 254 - 0xfe
      11'h6DD: dout  = 8'b11111111; // 1757 : 255 - 0xff
      11'h6DE: dout  = 8'b11111111; // 1758 : 255 - 0xff
      11'h6DF: dout  = 8'b01111110; // 1759 : 126 - 0x7e
      11'h6E0: dout  = 8'b00000000; // 1760 :   0 - 0x0 -- Background 0xdc
      11'h6E1: dout  = 8'b00000000; // 1761 :   0 - 0x0
      11'h6E2: dout  = 8'b00000000; // 1762 :   0 - 0x0
      11'h6E3: dout  = 8'b00000000; // 1763 :   0 - 0x0
      11'h6E4: dout  = 8'b00000000; // 1764 :   0 - 0x0
      11'h6E5: dout  = 8'b00000000; // 1765 :   0 - 0x0
      11'h6E6: dout  = 8'b00100001; // 1766 :  33 - 0x21
      11'h6E7: dout  = 8'b00111111; // 1767 :  63 - 0x3f
      11'h6E8: dout  = 8'b00111111; // 1768 :  63 - 0x3f -- Background 0xdd
      11'h6E9: dout  = 8'b00011111; // 1769 :  31 - 0x1f
      11'h6EA: dout  = 8'b00011111; // 1770 :  31 - 0x1f
      11'h6EB: dout  = 8'b00001111; // 1771 :  15 - 0xf
      11'h6EC: dout  = 8'b00000111; // 1772 :   7 - 0x7
      11'h6ED: dout  = 8'b00000011; // 1773 :   3 - 0x3
      11'h6EE: dout  = 8'b00000000; // 1774 :   0 - 0x0
      11'h6EF: dout  = 8'b00000000; // 1775 :   0 - 0x0
      11'h6F0: dout  = 8'b00111110; // 1776 :  62 - 0x3e -- Background 0xde
      11'h6F1: dout  = 8'b00011110; // 1777 :  30 - 0x1e
      11'h6F2: dout  = 8'b00011110; // 1778 :  30 - 0x1e
      11'h6F3: dout  = 8'b00001110; // 1779 :  14 - 0xe
      11'h6F4: dout  = 8'b00001111; // 1780 :  15 - 0xf
      11'h6F5: dout  = 8'b00011111; // 1781 :  31 - 0x1f
      11'h6F6: dout  = 8'b10011111; // 1782 : 159 - 0x9f
      11'h6F7: dout  = 8'b10011111; // 1783 : 159 - 0x9f
      11'h6F8: dout  = 8'b11011111; // 1784 : 223 - 0xdf -- Background 0xdf
      11'h6F9: dout  = 8'b11111111; // 1785 : 255 - 0xff
      11'h6FA: dout  = 8'b11111111; // 1786 : 255 - 0xff
      11'h6FB: dout  = 8'b11111111; // 1787 : 255 - 0xff
      11'h6FC: dout  = 8'b11111111; // 1788 : 255 - 0xff
      11'h6FD: dout  = 8'b11011111; // 1789 : 223 - 0xdf
      11'h6FE: dout  = 8'b11100111; // 1790 : 231 - 0xe7
      11'h6FF: dout  = 8'b00000000; // 1791 :   0 - 0x0
      11'h700: dout  = 8'b00100000; // 1792 :  32 - 0x20 -- Background 0xe0
      11'h701: dout  = 8'b00001111; // 1793 :  15 - 0xf
      11'h702: dout  = 8'b00110000; // 1794 :  48 - 0x30
      11'h703: dout  = 8'b01000000; // 1795 :  64 - 0x40
      11'h704: dout  = 8'b10011000; // 1796 : 152 - 0x98
      11'h705: dout  = 8'b00111110; // 1797 :  62 - 0x3e
      11'h706: dout  = 8'b00011111; // 1798 :  31 - 0x1f
      11'h707: dout  = 8'b00000000; // 1799 :   0 - 0x0
      11'h708: dout  = 8'b10000001; // 1800 : 129 - 0x81 -- Background 0xe1
      11'h709: dout  = 8'b00110110; // 1801 :  54 - 0x36
      11'h70A: dout  = 8'b00101110; // 1802 :  46 - 0x2e
      11'h70B: dout  = 8'b10101111; // 1803 : 175 - 0xaf
      11'h70C: dout  = 8'b10101110; // 1804 : 174 - 0xae
      11'h70D: dout  = 8'b11010001; // 1805 : 209 - 0xd1
      11'h70E: dout  = 8'b11101111; // 1806 : 239 - 0xef
      11'h70F: dout  = 8'b10000111; // 1807 : 135 - 0x87
      11'h710: dout  = 8'b00000010; // 1808 :   2 - 0x2 -- Background 0xe2
      11'h711: dout  = 8'b11111000; // 1809 : 248 - 0xf8
      11'h712: dout  = 8'b00000110; // 1810 :   6 - 0x6
      11'h713: dout  = 8'b00000001; // 1811 :   1 - 0x1
      11'h714: dout  = 8'b00001100; // 1812 :  12 - 0xc
      11'h715: dout  = 8'b00111110; // 1813 :  62 - 0x3e
      11'h716: dout  = 8'b11111100; // 1814 : 252 - 0xfc
      11'h717: dout  = 8'b00000000; // 1815 :   0 - 0x0
      11'h718: dout  = 8'b11000000; // 1816 : 192 - 0xc0 -- Background 0xe3
      11'h719: dout  = 8'b00110110; // 1817 :  54 - 0x36
      11'h71A: dout  = 8'b00111110; // 1818 :  62 - 0x3e
      11'h71B: dout  = 8'b01111010; // 1819 : 122 - 0x7a
      11'h71C: dout  = 8'b10110110; // 1820 : 182 - 0xb6
      11'h71D: dout  = 8'b11001101; // 1821 : 205 - 0xcd
      11'h71E: dout  = 8'b11111011; // 1822 : 251 - 0xfb
      11'h71F: dout  = 8'b11110000; // 1823 : 240 - 0xf0
      11'h720: dout  = 8'b00111110; // 1824 :  62 - 0x3e -- Background 0xe4
      11'h721: dout  = 8'b00111100; // 1825 :  60 - 0x3c
      11'h722: dout  = 8'b00111100; // 1826 :  60 - 0x3c
      11'h723: dout  = 8'b00111000; // 1827 :  56 - 0x38
      11'h724: dout  = 8'b11111000; // 1828 : 248 - 0xf8
      11'h725: dout  = 8'b01111100; // 1829 : 124 - 0x7c
      11'h726: dout  = 8'b01111110; // 1830 : 126 - 0x7e
      11'h727: dout  = 8'b01111000; // 1831 : 120 - 0x78
      11'h728: dout  = 8'b11111000; // 1832 : 248 - 0xf8 -- Background 0xe5
      11'h729: dout  = 8'b01111111; // 1833 : 127 - 0x7f
      11'h72A: dout  = 8'b01111111; // 1834 : 127 - 0x7f
      11'h72B: dout  = 8'b11111110; // 1835 : 254 - 0xfe
      11'h72C: dout  = 8'b11111111; // 1836 : 255 - 0xff
      11'h72D: dout  = 8'b11111111; // 1837 : 255 - 0xff
      11'h72E: dout  = 8'b11110011; // 1838 : 243 - 0xf3
      11'h72F: dout  = 8'b10000001; // 1839 : 129 - 0x81
      11'h730: dout  = 8'b00000000; // 1840 :   0 - 0x0 -- Background 0xe6
      11'h731: dout  = 8'b00000000; // 1841 :   0 - 0x0
      11'h732: dout  = 8'b00000000; // 1842 :   0 - 0x0
      11'h733: dout  = 8'b00010000; // 1843 :  16 - 0x10
      11'h734: dout  = 8'b01000000; // 1844 :  64 - 0x40
      11'h735: dout  = 8'b00100000; // 1845 :  32 - 0x20
      11'h736: dout  = 8'b00000000; // 1846 :   0 - 0x0
      11'h737: dout  = 8'b00000000; // 1847 :   0 - 0x0
      11'h738: dout  = 8'b00000110; // 1848 :   6 - 0x6 -- Background 0xe7
      11'h739: dout  = 8'b00001110; // 1849 :  14 - 0xe
      11'h73A: dout  = 8'b01111110; // 1850 : 126 - 0x7e
      11'h73B: dout  = 8'b11111110; // 1851 : 254 - 0xfe
      11'h73C: dout  = 8'b11111110; // 1852 : 254 - 0xfe
      11'h73D: dout  = 8'b11111100; // 1853 : 252 - 0xfc
      11'h73E: dout  = 8'b11111000; // 1854 : 248 - 0xf8
      11'h73F: dout  = 8'b11110000; // 1855 : 240 - 0xf0
      11'h740: dout  = 8'b00000000; // 1856 :   0 - 0x0 -- Background 0xe8
      11'h741: dout  = 8'b00000000; // 1857 :   0 - 0x0
      11'h742: dout  = 8'b00000000; // 1858 :   0 - 0x0
      11'h743: dout  = 8'b00000000; // 1859 :   0 - 0x0
      11'h744: dout  = 8'b00000000; // 1860 :   0 - 0x0
      11'h745: dout  = 8'b00000000; // 1861 :   0 - 0x0
      11'h746: dout  = 8'b00000000; // 1862 :   0 - 0x0
      11'h747: dout  = 8'b00000001; // 1863 :   1 - 0x1
      11'h748: dout  = 8'b00000010; // 1864 :   2 - 0x2 -- Background 0xe9
      11'h749: dout  = 8'b00000000; // 1865 :   0 - 0x0
      11'h74A: dout  = 8'b00001000; // 1866 :   8 - 0x8
      11'h74B: dout  = 8'b00000001; // 1867 :   1 - 0x1
      11'h74C: dout  = 8'b00010011; // 1868 :  19 - 0x13
      11'h74D: dout  = 8'b00000001; // 1869 :   1 - 0x1
      11'h74E: dout  = 8'b00000000; // 1870 :   0 - 0x0
      11'h74F: dout  = 8'b00000000; // 1871 :   0 - 0x0
      11'h750: dout  = 8'b00000000; // 1872 :   0 - 0x0 -- Background 0xea
      11'h751: dout  = 8'b00000000; // 1873 :   0 - 0x0
      11'h752: dout  = 8'b00000000; // 1874 :   0 - 0x0
      11'h753: dout  = 8'b00000000; // 1875 :   0 - 0x0
      11'h754: dout  = 8'b00000000; // 1876 :   0 - 0x0
      11'h755: dout  = 8'b00000000; // 1877 :   0 - 0x0
      11'h756: dout  = 8'b00000000; // 1878 :   0 - 0x0
      11'h757: dout  = 8'b00000000; // 1879 :   0 - 0x0
      11'h758: dout  = 8'b00000000; // 1880 :   0 - 0x0 -- Background 0xeb
      11'h759: dout  = 8'b01000011; // 1881 :  67 - 0x43
      11'h75A: dout  = 8'b01111111; // 1882 : 127 - 0x7f
      11'h75B: dout  = 8'b01111111; // 1883 : 127 - 0x7f
      11'h75C: dout  = 8'b01111111; // 1884 : 127 - 0x7f
      11'h75D: dout  = 8'b00111111; // 1885 :  63 - 0x3f
      11'h75E: dout  = 8'b00011111; // 1886 :  31 - 0x1f
      11'h75F: dout  = 8'b00000111; // 1887 :   7 - 0x7
      11'h760: dout  = 8'b00000000; // 1888 :   0 - 0x0 -- Background 0xec
      11'h761: dout  = 8'b00000000; // 1889 :   0 - 0x0
      11'h762: dout  = 8'b00000000; // 1890 :   0 - 0x0
      11'h763: dout  = 8'b00000000; // 1891 :   0 - 0x0
      11'h764: dout  = 8'b00000000; // 1892 :   0 - 0x0
      11'h765: dout  = 8'b00000000; // 1893 :   0 - 0x0
      11'h766: dout  = 8'b11000000; // 1894 : 192 - 0xc0
      11'h767: dout  = 8'b00000000; // 1895 :   0 - 0x0
      11'h768: dout  = 8'b00010000; // 1896 :  16 - 0x10 -- Background 0xed
      11'h769: dout  = 8'b00111000; // 1897 :  56 - 0x38
      11'h76A: dout  = 8'b10111111; // 1898 : 191 - 0xbf
      11'h76B: dout  = 8'b11111111; // 1899 : 255 - 0xff
      11'h76C: dout  = 8'b11111111; // 1900 : 255 - 0xff
      11'h76D: dout  = 8'b11111111; // 1901 : 255 - 0xff
      11'h76E: dout  = 8'b11111111; // 1902 : 255 - 0xff
      11'h76F: dout  = 8'b11111111; // 1903 : 255 - 0xff
      11'h770: dout  = 8'b01111110; // 1904 : 126 - 0x7e -- Background 0xee
      11'h771: dout  = 8'b00011110; // 1905 :  30 - 0x1e
      11'h772: dout  = 8'b00011110; // 1906 :  30 - 0x1e
      11'h773: dout  = 8'b00001110; // 1907 :  14 - 0xe
      11'h774: dout  = 8'b00001111; // 1908 :  15 - 0xf
      11'h775: dout  = 8'b00011110; // 1909 :  30 - 0x1e
      11'h776: dout  = 8'b00011110; // 1910 :  30 - 0x1e
      11'h777: dout  = 8'b00111110; // 1911 :  62 - 0x3e
      11'h778: dout  = 8'b01111111; // 1912 : 127 - 0x7f -- Background 0xef
      11'h779: dout  = 8'b01111111; // 1913 : 127 - 0x7f
      11'h77A: dout  = 8'b10111111; // 1914 : 191 - 0xbf
      11'h77B: dout  = 8'b11111111; // 1915 : 255 - 0xff
      11'h77C: dout  = 8'b11111111; // 1916 : 255 - 0xff
      11'h77D: dout  = 8'b11111111; // 1917 : 255 - 0xff
      11'h77E: dout  = 8'b11100111; // 1918 : 231 - 0xe7
      11'h77F: dout  = 8'b11000000; // 1919 : 192 - 0xc0
      11'h780: dout  = 8'b00000000; // 1920 :   0 - 0x0 -- Background 0xf0
      11'h781: dout  = 8'b00000000; // 1921 :   0 - 0x0
      11'h782: dout  = 8'b00010000; // 1922 :  16 - 0x10
      11'h783: dout  = 8'b11111101; // 1923 : 253 - 0xfd
      11'h784: dout  = 8'b11111010; // 1924 : 250 - 0xfa
      11'h785: dout  = 8'b11101011; // 1925 : 235 - 0xeb
      11'h786: dout  = 8'b10000000; // 1926 : 128 - 0x80
      11'h787: dout  = 8'b00000000; // 1927 :   0 - 0x0
      11'h788: dout  = 8'b00100000; // 1928 :  32 - 0x20 -- Background 0xf1
      11'h789: dout  = 8'b00011111; // 1929 :  31 - 0x1f
      11'h78A: dout  = 8'b01100000; // 1930 :  96 - 0x60
      11'h78B: dout  = 8'b10001110; // 1931 : 142 - 0x8e
      11'h78C: dout  = 8'b00111111; // 1932 :  63 - 0x3f
      11'h78D: dout  = 8'b01111111; // 1933 : 127 - 0x7f
      11'h78E: dout  = 8'b01111111; // 1934 : 127 - 0x7f
      11'h78F: dout  = 8'b01111100; // 1935 : 124 - 0x7c
      11'h790: dout  = 8'b00111001; // 1936 :  57 - 0x39 -- Background 0xf2
      11'h791: dout  = 8'b00110110; // 1937 :  54 - 0x36
      11'h792: dout  = 8'b00101110; // 1938 :  46 - 0x2e
      11'h793: dout  = 8'b10101111; // 1939 : 175 - 0xaf
      11'h794: dout  = 8'b10101110; // 1940 : 174 - 0xae
      11'h795: dout  = 8'b11010001; // 1941 : 209 - 0xd1
      11'h796: dout  = 8'b11101111; // 1942 : 239 - 0xef
      11'h797: dout  = 8'b10000111; // 1943 : 135 - 0x87
      11'h798: dout  = 8'b00000000; // 1944 :   0 - 0x0 -- Background 0xf3
      11'h799: dout  = 8'b00000000; // 1945 :   0 - 0x0
      11'h79A: dout  = 8'b00000100; // 1946 :   4 - 0x4
      11'h79B: dout  = 8'b01011111; // 1947 :  95 - 0x5f
      11'h79C: dout  = 8'b10101111; // 1948 : 175 - 0xaf
      11'h79D: dout  = 8'b01010011; // 1949 :  83 - 0x53
      11'h79E: dout  = 8'b00000000; // 1950 :   0 - 0x0
      11'h79F: dout  = 8'b00000000; // 1951 :   0 - 0x0
      11'h7A0: dout  = 8'b00000010; // 1952 :   2 - 0x2 -- Background 0xf4
      11'h7A1: dout  = 8'b11111100; // 1953 : 252 - 0xfc
      11'h7A2: dout  = 8'b00000011; // 1954 :   3 - 0x3
      11'h7A3: dout  = 8'b00111000; // 1955 :  56 - 0x38
      11'h7A4: dout  = 8'b11111110; // 1956 : 254 - 0xfe
      11'h7A5: dout  = 8'b11111111; // 1957 : 255 - 0xff
      11'h7A6: dout  = 8'b11111111; // 1958 : 255 - 0xff
      11'h7A7: dout  = 8'b00011110; // 1959 :  30 - 0x1e
      11'h7A8: dout  = 8'b11000000; // 1960 : 192 - 0xc0 -- Background 0xf5
      11'h7A9: dout  = 8'b00110110; // 1961 :  54 - 0x36
      11'h7AA: dout  = 8'b00111110; // 1962 :  62 - 0x3e
      11'h7AB: dout  = 8'b01111010; // 1963 : 122 - 0x7a
      11'h7AC: dout  = 8'b10110110; // 1964 : 182 - 0xb6
      11'h7AD: dout  = 8'b11001101; // 1965 : 205 - 0xcd
      11'h7AE: dout  = 8'b11111011; // 1966 : 251 - 0xfb
      11'h7AF: dout  = 8'b11110000; // 1967 : 240 - 0xf0
      11'h7B0: dout  = 8'b00000000; // 1968 :   0 - 0x0 -- Background 0xf6
      11'h7B1: dout  = 8'b00000000; // 1969 :   0 - 0x0
      11'h7B2: dout  = 8'b00000000; // 1970 :   0 - 0x0
      11'h7B3: dout  = 8'b00000000; // 1971 :   0 - 0x0
      11'h7B4: dout  = 8'b00000000; // 1972 :   0 - 0x0
      11'h7B5: dout  = 8'b00001110; // 1973 :  14 - 0xe
      11'h7B6: dout  = 8'b00001000; // 1974 :   8 - 0x8
      11'h7B7: dout  = 8'b00001000; // 1975 :   8 - 0x8
      11'h7B8: dout  = 8'b00011111; // 1976 :  31 - 0x1f -- Background 0xf7
      11'h7B9: dout  = 8'b00111111; // 1977 :  63 - 0x3f
      11'h7BA: dout  = 8'b11111111; // 1978 : 255 - 0xff
      11'h7BB: dout  = 8'b11111111; // 1979 : 255 - 0xff
      11'h7BC: dout  = 8'b11111111; // 1980 : 255 - 0xff
      11'h7BD: dout  = 8'b11111111; // 1981 : 255 - 0xff
      11'h7BE: dout  = 8'b11111111; // 1982 : 255 - 0xff
      11'h7BF: dout  = 8'b01111111; // 1983 : 127 - 0x7f
      11'h7C0: dout  = 8'b00111111; // 1984 :  63 - 0x3f -- Background 0xf8
      11'h7C1: dout  = 8'b00111110; // 1985 :  62 - 0x3e
      11'h7C2: dout  = 8'b00111100; // 1986 :  60 - 0x3c
      11'h7C3: dout  = 8'b10111000; // 1987 : 184 - 0xb8
      11'h7C4: dout  = 8'b01111000; // 1988 : 120 - 0x78
      11'h7C5: dout  = 8'b01111000; // 1989 : 120 - 0x78
      11'h7C6: dout  = 8'b01111110; // 1990 : 126 - 0x7e
      11'h7C7: dout  = 8'b01111110; // 1991 : 126 - 0x7e
      11'h7C8: dout  = 8'b11111101; // 1992 : 253 - 0xfd -- Background 0xf9
      11'h7C9: dout  = 8'b01111001; // 1993 : 121 - 0x79
      11'h7CA: dout  = 8'b01111011; // 1994 : 123 - 0x7b
      11'h7CB: dout  = 8'b11111111; // 1995 : 255 - 0xff
      11'h7CC: dout  = 8'b11111111; // 1996 : 255 - 0xff
      11'h7CD: dout  = 8'b11111111; // 1997 : 255 - 0xff
      11'h7CE: dout  = 8'b11110011; // 1998 : 243 - 0xf3
      11'h7CF: dout  = 8'b10000000; // 1999 : 128 - 0x80
      11'h7D0: dout  = 8'b00000000; // 2000 :   0 - 0x0 -- Background 0xfa
      11'h7D1: dout  = 8'b00000000; // 2001 :   0 - 0x0
      11'h7D2: dout  = 8'b00000000; // 2002 :   0 - 0x0
      11'h7D3: dout  = 8'b00000000; // 2003 :   0 - 0x0
      11'h7D4: dout  = 8'b00000000; // 2004 :   0 - 0x0
      11'h7D5: dout  = 8'b00000000; // 2005 :   0 - 0x0
      11'h7D6: dout  = 8'b00000000; // 2006 :   0 - 0x0
      11'h7D7: dout  = 8'b00000000; // 2007 :   0 - 0x0
      11'h7D8: dout  = 8'b00010000; // 2008 :  16 - 0x10 -- Background 0xfb
      11'h7D9: dout  = 8'b10000100; // 2009 : 132 - 0x84
      11'h7DA: dout  = 8'b11100000; // 2010 : 224 - 0xe0
      11'h7DB: dout  = 8'b11000000; // 2011 : 192 - 0xc0
      11'h7DC: dout  = 8'b10000000; // 2012 : 128 - 0x80
      11'h7DD: dout  = 8'b10000000; // 2013 : 128 - 0x80
      11'h7DE: dout  = 8'b00000000; // 2014 :   0 - 0x0
      11'h7DF: dout  = 8'b00000000; // 2015 :   0 - 0x0
      11'h7E0: dout  = 8'b00000000; // 2016 :   0 - 0x0 -- Background 0xfc
      11'h7E1: dout  = 8'b01001000; // 2017 :  72 - 0x48
      11'h7E2: dout  = 8'b00100000; // 2018 :  32 - 0x20
      11'h7E3: dout  = 8'b00000000; // 2019 :   0 - 0x0
      11'h7E4: dout  = 8'b00000000; // 2020 :   0 - 0x0
      11'h7E5: dout  = 8'b00000100; // 2021 :   4 - 0x4
      11'h7E6: dout  = 8'b00001110; // 2022 :  14 - 0xe
      11'h7E7: dout  = 8'b11111110; // 2023 : 254 - 0xfe
      11'h7E8: dout  = 8'b11111110; // 2024 : 254 - 0xfe -- Background 0xfd
      11'h7E9: dout  = 8'b11111100; // 2025 : 252 - 0xfc
      11'h7EA: dout  = 8'b11111100; // 2026 : 252 - 0xfc
      11'h7EB: dout  = 8'b11111000; // 2027 : 248 - 0xf8
      11'h7EC: dout  = 8'b11110000; // 2028 : 240 - 0xf0
      11'h7ED: dout  = 8'b11100000; // 2029 : 224 - 0xe0
      11'h7EE: dout  = 8'b10000000; // 2030 : 128 - 0x80
      11'h7EF: dout  = 8'b00000000; // 2031 :   0 - 0x0
      11'h7F0: dout  = 8'b00001111; // 2032 :  15 - 0xf -- Background 0xfe
      11'h7F1: dout  = 8'b00000110; // 2033 :   6 - 0x6
      11'h7F2: dout  = 8'b00000110; // 2034 :   6 - 0x6
      11'h7F3: dout  = 8'b00000110; // 2035 :   6 - 0x6
      11'h7F4: dout  = 8'b00000110; // 2036 :   6 - 0x6
      11'h7F5: dout  = 8'b00000110; // 2037 :   6 - 0x6
      11'h7F6: dout  = 8'b00001111; // 2038 :  15 - 0xf
      11'h7F7: dout  = 8'b00000000; // 2039 :   0 - 0x0
      11'h7F8: dout  = 8'b11110000; // 2040 : 240 - 0xf0 -- Background 0xff
      11'h7F9: dout  = 8'b01100000; // 2041 :  96 - 0x60
      11'h7FA: dout  = 8'b01100000; // 2042 :  96 - 0x60
      11'h7FB: dout  = 8'b01100110; // 2043 : 102 - 0x66
      11'h7FC: dout  = 8'b01100110; // 2044 : 102 - 0x66
      11'h7FD: dout  = 8'b01100000; // 2045 :  96 - 0x60
      11'h7FE: dout  = 8'b11110000; // 2046 : 240 - 0xf0
      11'h7FF: dout  = 8'b00000000; // 2047 :   0 - 0x0
    endcase
  end

endmodule
