//- Autcmatically generated verilog ROM from a NES memory file----
//-   NAME TABLE
// https://wiki.nesdev.com/w/index.php/PPU_nametables
//- Only the first Name Table: 1KiB


//-  Original memory dump file name: sprilo_menuscr.bin --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_NTABLE0_SPRILO_MENU
  (
     input     clk,   // clock
     input      [10-1:0] addr,  //1024 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
     //----- Name Table 0---------
      10'h0: dout <= 8'b11111010; //    0 : 250 - 0xfa -- line 0x0
      10'h1: dout <= 8'b11111010; //    1 : 250 - 0xfa
      10'h2: dout <= 8'b11111010; //    2 : 250 - 0xfa
      10'h3: dout <= 8'b11111010; //    3 : 250 - 0xfa
      10'h4: dout <= 8'b11111010; //    4 : 250 - 0xfa
      10'h5: dout <= 8'b11111010; //    5 : 250 - 0xfa
      10'h6: dout <= 8'b11111010; //    6 : 250 - 0xfa
      10'h7: dout <= 8'b11111010; //    7 : 250 - 0xfa
      10'h8: dout <= 8'b11111010; //    8 : 250 - 0xfa
      10'h9: dout <= 8'b11111010; //    9 : 250 - 0xfa
      10'hA: dout <= 8'b11111010; //   10 : 250 - 0xfa
      10'hB: dout <= 8'b11111010; //   11 : 250 - 0xfa
      10'hC: dout <= 8'b11111010; //   12 : 250 - 0xfa
      10'hD: dout <= 8'b11111010; //   13 : 250 - 0xfa
      10'hE: dout <= 8'b11111010; //   14 : 250 - 0xfa
      10'hF: dout <= 8'b11111010; //   15 : 250 - 0xfa
      10'h10: dout <= 8'b11111010; //   16 : 250 - 0xfa
      10'h11: dout <= 8'b11111010; //   17 : 250 - 0xfa
      10'h12: dout <= 8'b11111010; //   18 : 250 - 0xfa
      10'h13: dout <= 8'b11111010; //   19 : 250 - 0xfa
      10'h14: dout <= 8'b11111010; //   20 : 250 - 0xfa
      10'h15: dout <= 8'b11111010; //   21 : 250 - 0xfa
      10'h16: dout <= 8'b11111010; //   22 : 250 - 0xfa
      10'h17: dout <= 8'b11111010; //   23 : 250 - 0xfa
      10'h18: dout <= 8'b11111010; //   24 : 250 - 0xfa
      10'h19: dout <= 8'b11111010; //   25 : 250 - 0xfa
      10'h1A: dout <= 8'b11111010; //   26 : 250 - 0xfa
      10'h1B: dout <= 8'b11111010; //   27 : 250 - 0xfa
      10'h1C: dout <= 8'b11111010; //   28 : 250 - 0xfa
      10'h1D: dout <= 8'b11111010; //   29 : 250 - 0xfa
      10'h1E: dout <= 8'b11111010; //   30 : 250 - 0xfa
      10'h1F: dout <= 8'b11111010; //   31 : 250 - 0xfa
      10'h20: dout <= 8'b11111010; //   32 : 250 - 0xfa -- line 0x1
      10'h21: dout <= 8'b11111010; //   33 : 250 - 0xfa
      10'h22: dout <= 8'b11111010; //   34 : 250 - 0xfa
      10'h23: dout <= 8'b11111010; //   35 : 250 - 0xfa
      10'h24: dout <= 8'b11111010; //   36 : 250 - 0xfa
      10'h25: dout <= 8'b11111010; //   37 : 250 - 0xfa
      10'h26: dout <= 8'b11111010; //   38 : 250 - 0xfa
      10'h27: dout <= 8'b11111001; //   39 : 249 - 0xf9
      10'h28: dout <= 8'b11111010; //   40 : 250 - 0xfa
      10'h29: dout <= 8'b11111010; //   41 : 250 - 0xfa
      10'h2A: dout <= 8'b11111010; //   42 : 250 - 0xfa
      10'h2B: dout <= 8'b11111010; //   43 : 250 - 0xfa
      10'h2C: dout <= 8'b11111010; //   44 : 250 - 0xfa
      10'h2D: dout <= 8'b11111010; //   45 : 250 - 0xfa
      10'h2E: dout <= 8'b11111010; //   46 : 250 - 0xfa
      10'h2F: dout <= 8'b11111010; //   47 : 250 - 0xfa
      10'h30: dout <= 8'b11111010; //   48 : 250 - 0xfa
      10'h31: dout <= 8'b11111001; //   49 : 249 - 0xf9
      10'h32: dout <= 8'b11111010; //   50 : 250 - 0xfa
      10'h33: dout <= 8'b11111010; //   51 : 250 - 0xfa
      10'h34: dout <= 8'b11111010; //   52 : 250 - 0xfa
      10'h35: dout <= 8'b11111010; //   53 : 250 - 0xfa
      10'h36: dout <= 8'b11111010; //   54 : 250 - 0xfa
      10'h37: dout <= 8'b11111010; //   55 : 250 - 0xfa
      10'h38: dout <= 8'b11111010; //   56 : 250 - 0xfa
      10'h39: dout <= 8'b11111010; //   57 : 250 - 0xfa
      10'h3A: dout <= 8'b11111010; //   58 : 250 - 0xfa
      10'h3B: dout <= 8'b11111010; //   59 : 250 - 0xfa
      10'h3C: dout <= 8'b11111001; //   60 : 249 - 0xf9
      10'h3D: dout <= 8'b11111010; //   61 : 250 - 0xfa
      10'h3E: dout <= 8'b11111010; //   62 : 250 - 0xfa
      10'h3F: dout <= 8'b11111010; //   63 : 250 - 0xfa
      10'h40: dout <= 8'b11111010; //   64 : 250 - 0xfa -- line 0x2
      10'h41: dout <= 8'b11111010; //   65 : 250 - 0xfa
      10'h42: dout <= 8'b11111010; //   66 : 250 - 0xfa
      10'h43: dout <= 8'b11111010; //   67 : 250 - 0xfa
      10'h44: dout <= 8'b11111010; //   68 : 250 - 0xfa
      10'h45: dout <= 8'b11111010; //   69 : 250 - 0xfa
      10'h46: dout <= 8'b11111010; //   70 : 250 - 0xfa
      10'h47: dout <= 8'b11111010; //   71 : 250 - 0xfa
      10'h48: dout <= 8'b11111010; //   72 : 250 - 0xfa
      10'h49: dout <= 8'b11111010; //   73 : 250 - 0xfa
      10'h4A: dout <= 8'b11111001; //   74 : 249 - 0xf9
      10'h4B: dout <= 8'b11111010; //   75 : 250 - 0xfa
      10'h4C: dout <= 8'b11111010; //   76 : 250 - 0xfa
      10'h4D: dout <= 8'b11111010; //   77 : 250 - 0xfa
      10'h4E: dout <= 8'b11101010; //   78 : 234 - 0xea
      10'h4F: dout <= 8'b11111010; //   79 : 250 - 0xfa
      10'h50: dout <= 8'b11111010; //   80 : 250 - 0xfa
      10'h51: dout <= 8'b11111010; //   81 : 250 - 0xfa
      10'h52: dout <= 8'b11111010; //   82 : 250 - 0xfa
      10'h53: dout <= 8'b11111010; //   83 : 250 - 0xfa
      10'h54: dout <= 8'b11111010; //   84 : 250 - 0xfa
      10'h55: dout <= 8'b11111010; //   85 : 250 - 0xfa
      10'h56: dout <= 8'b11111010; //   86 : 250 - 0xfa
      10'h57: dout <= 8'b11111010; //   87 : 250 - 0xfa
      10'h58: dout <= 8'b11111010; //   88 : 250 - 0xfa
      10'h59: dout <= 8'b11111010; //   89 : 250 - 0xfa
      10'h5A: dout <= 8'b11111010; //   90 : 250 - 0xfa
      10'h5B: dout <= 8'b11111010; //   91 : 250 - 0xfa
      10'h5C: dout <= 8'b11111010; //   92 : 250 - 0xfa
      10'h5D: dout <= 8'b11111010; //   93 : 250 - 0xfa
      10'h5E: dout <= 8'b11111010; //   94 : 250 - 0xfa
      10'h5F: dout <= 8'b11111010; //   95 : 250 - 0xfa
      10'h60: dout <= 8'b11111010; //   96 : 250 - 0xfa -- line 0x3
      10'h61: dout <= 8'b11111010; //   97 : 250 - 0xfa
      10'h62: dout <= 8'b11111010; //   98 : 250 - 0xfa
      10'h63: dout <= 8'b11111010; //   99 : 250 - 0xfa
      10'h64: dout <= 8'b11111010; //  100 : 250 - 0xfa
      10'h65: dout <= 8'b11111010; //  101 : 250 - 0xfa
      10'h66: dout <= 8'b11111010; //  102 : 250 - 0xfa
      10'h67: dout <= 8'b11111010; //  103 : 250 - 0xfa
      10'h68: dout <= 8'b11111010; //  104 : 250 - 0xfa
      10'h69: dout <= 8'b11111010; //  105 : 250 - 0xfa
      10'h6A: dout <= 8'b11111010; //  106 : 250 - 0xfa
      10'h6B: dout <= 8'b11111010; //  107 : 250 - 0xfa
      10'h6C: dout <= 8'b11111010; //  108 : 250 - 0xfa
      10'h6D: dout <= 8'b11111010; //  109 : 250 - 0xfa
      10'h6E: dout <= 8'b11111010; //  110 : 250 - 0xfa
      10'h6F: dout <= 8'b11111010; //  111 : 250 - 0xfa
      10'h70: dout <= 8'b11111010; //  112 : 250 - 0xfa
      10'h71: dout <= 8'b11111010; //  113 : 250 - 0xfa
      10'h72: dout <= 8'b11111010; //  114 : 250 - 0xfa
      10'h73: dout <= 8'b11111010; //  115 : 250 - 0xfa
      10'h74: dout <= 8'b11111010; //  116 : 250 - 0xfa
      10'h75: dout <= 8'b11111010; //  117 : 250 - 0xfa
      10'h76: dout <= 8'b11111010; //  118 : 250 - 0xfa
      10'h77: dout <= 8'b11111010; //  119 : 250 - 0xfa
      10'h78: dout <= 8'b11111010; //  120 : 250 - 0xfa
      10'h79: dout <= 8'b11101010; //  121 : 234 - 0xea
      10'h7A: dout <= 8'b11111010; //  122 : 250 - 0xfa
      10'h7B: dout <= 8'b11111010; //  123 : 250 - 0xfa
      10'h7C: dout <= 8'b11111010; //  124 : 250 - 0xfa
      10'h7D: dout <= 8'b11101010; //  125 : 234 - 0xea
      10'h7E: dout <= 8'b11111010; //  126 : 250 - 0xfa
      10'h7F: dout <= 8'b11111010; //  127 : 250 - 0xfa
      10'h80: dout <= 8'b11111010; //  128 : 250 - 0xfa -- line 0x4
      10'h81: dout <= 8'b11111010; //  129 : 250 - 0xfa
      10'h82: dout <= 8'b11111010; //  130 : 250 - 0xfa
      10'h83: dout <= 8'b11111010; //  131 : 250 - 0xfa
      10'h84: dout <= 8'b11101010; //  132 : 234 - 0xea
      10'h85: dout <= 8'b11111010; //  133 : 250 - 0xfa
      10'h86: dout <= 8'b11111010; //  134 : 250 - 0xfa
      10'h87: dout <= 8'b11111001; //  135 : 249 - 0xf9
      10'h88: dout <= 8'b11111010; //  136 : 250 - 0xfa
      10'h89: dout <= 8'b11111010; //  137 : 250 - 0xfa
      10'h8A: dout <= 8'b11111010; //  138 : 250 - 0xfa
      10'h8B: dout <= 8'b11111010; //  139 : 250 - 0xfa
      10'h8C: dout <= 8'b11111010; //  140 : 250 - 0xfa
      10'h8D: dout <= 8'b11111010; //  141 : 250 - 0xfa
      10'h8E: dout <= 8'b11111010; //  142 : 250 - 0xfa
      10'h8F: dout <= 8'b11111010; //  143 : 250 - 0xfa
      10'h90: dout <= 8'b11111010; //  144 : 250 - 0xfa
      10'h91: dout <= 8'b11111010; //  145 : 250 - 0xfa
      10'h92: dout <= 8'b11111010; //  146 : 250 - 0xfa
      10'h93: dout <= 8'b11111010; //  147 : 250 - 0xfa
      10'h94: dout <= 8'b11111010; //  148 : 250 - 0xfa
      10'h95: dout <= 8'b11111001; //  149 : 249 - 0xf9
      10'h96: dout <= 8'b11111010; //  150 : 250 - 0xfa
      10'h97: dout <= 8'b11111010; //  151 : 250 - 0xfa
      10'h98: dout <= 8'b11111010; //  152 : 250 - 0xfa
      10'h99: dout <= 8'b11111010; //  153 : 250 - 0xfa
      10'h9A: dout <= 8'b11111010; //  154 : 250 - 0xfa
      10'h9B: dout <= 8'b11111010; //  155 : 250 - 0xfa
      10'h9C: dout <= 8'b11111010; //  156 : 250 - 0xfa
      10'h9D: dout <= 8'b11111010; //  157 : 250 - 0xfa
      10'h9E: dout <= 8'b11111010; //  158 : 250 - 0xfa
      10'h9F: dout <= 8'b11111010; //  159 : 250 - 0xfa
      10'hA0: dout <= 8'b11111010; //  160 : 250 - 0xfa -- line 0x5
      10'hA1: dout <= 8'b11111010; //  161 : 250 - 0xfa
      10'hA2: dout <= 8'b11111010; //  162 : 250 - 0xfa
      10'hA3: dout <= 8'b11111010; //  163 : 250 - 0xfa
      10'hA4: dout <= 8'b11111010; //  164 : 250 - 0xfa
      10'hA5: dout <= 8'b11111010; //  165 : 250 - 0xfa
      10'hA6: dout <= 8'b11111010; //  166 : 250 - 0xfa
      10'hA7: dout <= 8'b11111010; //  167 : 250 - 0xfa
      10'hA8: dout <= 8'b11111010; //  168 : 250 - 0xfa
      10'hA9: dout <= 8'b11111010; //  169 : 250 - 0xfa
      10'hAA: dout <= 8'b11111010; //  170 : 250 - 0xfa
      10'hAB: dout <= 8'b11001101; //  171 : 205 - 0xcd
      10'hAC: dout <= 8'b11101101; //  172 : 237 - 0xed
      10'hAD: dout <= 8'b11101101; //  173 : 237 - 0xed
      10'hAE: dout <= 8'b11101101; //  174 : 237 - 0xed
      10'hAF: dout <= 8'b11101101; //  175 : 237 - 0xed
      10'hB0: dout <= 8'b11101101; //  176 : 237 - 0xed
      10'hB1: dout <= 8'b11101101; //  177 : 237 - 0xed
      10'hB2: dout <= 8'b11101101; //  178 : 237 - 0xed
      10'hB3: dout <= 8'b11101101; //  179 : 237 - 0xed
      10'hB4: dout <= 8'b11001110; //  180 : 206 - 0xce
      10'hB5: dout <= 8'b11111010; //  181 : 250 - 0xfa
      10'hB6: dout <= 8'b11111010; //  182 : 250 - 0xfa
      10'hB7: dout <= 8'b11111010; //  183 : 250 - 0xfa
      10'hB8: dout <= 8'b11111010; //  184 : 250 - 0xfa
      10'hB9: dout <= 8'b11111010; //  185 : 250 - 0xfa
      10'hBA: dout <= 8'b11111010; //  186 : 250 - 0xfa
      10'hBB: dout <= 8'b11111010; //  187 : 250 - 0xfa
      10'hBC: dout <= 8'b11111010; //  188 : 250 - 0xfa
      10'hBD: dout <= 8'b11111010; //  189 : 250 - 0xfa
      10'hBE: dout <= 8'b11111010; //  190 : 250 - 0xfa
      10'hBF: dout <= 8'b11111010; //  191 : 250 - 0xfa
      10'hC0: dout <= 8'b11111001; //  192 : 249 - 0xf9 -- line 0x6
      10'hC1: dout <= 8'b11111010; //  193 : 250 - 0xfa
      10'hC2: dout <= 8'b11111010; //  194 : 250 - 0xfa
      10'hC3: dout <= 8'b11111010; //  195 : 250 - 0xfa
      10'hC4: dout <= 8'b11111010; //  196 : 250 - 0xfa
      10'hC5: dout <= 8'b11111010; //  197 : 250 - 0xfa
      10'hC6: dout <= 8'b11111010; //  198 : 250 - 0xfa
      10'hC7: dout <= 8'b11111010; //  199 : 250 - 0xfa
      10'hC8: dout <= 8'b11111010; //  200 : 250 - 0xfa
      10'hC9: dout <= 8'b11111010; //  201 : 250 - 0xfa
      10'hCA: dout <= 8'b11111010; //  202 : 250 - 0xfa
      10'hCB: dout <= 8'b11101110; //  203 : 238 - 0xee
      10'hCC: dout <= 8'b11111010; //  204 : 250 - 0xfa
      10'hCD: dout <= 8'b11111010; //  205 : 250 - 0xfa
      10'hCE: dout <= 8'b11111010; //  206 : 250 - 0xfa
      10'hCF: dout <= 8'b11111010; //  207 : 250 - 0xfa
      10'hD0: dout <= 8'b11111010; //  208 : 250 - 0xfa
      10'hD1: dout <= 8'b11111010; //  209 : 250 - 0xfa
      10'hD2: dout <= 8'b11111010; //  210 : 250 - 0xfa
      10'hD3: dout <= 8'b11111010; //  211 : 250 - 0xfa
      10'hD4: dout <= 8'b11101110; //  212 : 238 - 0xee
      10'hD5: dout <= 8'b11111010; //  213 : 250 - 0xfa
      10'hD6: dout <= 8'b11111010; //  214 : 250 - 0xfa
      10'hD7: dout <= 8'b11111010; //  215 : 250 - 0xfa
      10'hD8: dout <= 8'b11111010; //  216 : 250 - 0xfa
      10'hD9: dout <= 8'b11111010; //  217 : 250 - 0xfa
      10'hDA: dout <= 8'b11111010; //  218 : 250 - 0xfa
      10'hDB: dout <= 8'b11111001; //  219 : 249 - 0xf9
      10'hDC: dout <= 8'b11111010; //  220 : 250 - 0xfa
      10'hDD: dout <= 8'b11111010; //  221 : 250 - 0xfa
      10'hDE: dout <= 8'b11111010; //  222 : 250 - 0xfa
      10'hDF: dout <= 8'b11111010; //  223 : 250 - 0xfa
      10'hE0: dout <= 8'b11111010; //  224 : 250 - 0xfa -- line 0x7
      10'hE1: dout <= 8'b11111010; //  225 : 250 - 0xfa
      10'hE2: dout <= 8'b11111010; //  226 : 250 - 0xfa
      10'hE3: dout <= 8'b11111010; //  227 : 250 - 0xfa
      10'hE4: dout <= 8'b11111001; //  228 : 249 - 0xf9
      10'hE5: dout <= 8'b11111010; //  229 : 250 - 0xfa
      10'hE6: dout <= 8'b11111010; //  230 : 250 - 0xfa
      10'hE7: dout <= 8'b11111010; //  231 : 250 - 0xfa
      10'hE8: dout <= 8'b11111010; //  232 : 250 - 0xfa
      10'hE9: dout <= 8'b11111010; //  233 : 250 - 0xfa
      10'hEA: dout <= 8'b11111010; //  234 : 250 - 0xfa
      10'hEB: dout <= 8'b11101110; //  235 : 238 - 0xee
      10'hEC: dout <= 8'b11111010; //  236 : 250 - 0xfa
      10'hED: dout <= 8'b00100011; //  237 :  35 - 0x23
      10'hEE: dout <= 8'b00100000; //  238 :  32 - 0x20
      10'hEF: dout <= 8'b00100010; //  239 :  34 - 0x22
      10'hF0: dout <= 8'b00011001; //  240 :  25 - 0x19
      10'hF1: dout <= 8'b00011100; //  241 :  28 - 0x1c
      10'hF2: dout <= 8'b00011111; //  242 :  31 - 0x1f
      10'hF3: dout <= 8'b11111010; //  243 : 250 - 0xfa
      10'hF4: dout <= 8'b11101110; //  244 : 238 - 0xee
      10'hF5: dout <= 8'b11111010; //  245 : 250 - 0xfa
      10'hF6: dout <= 8'b11111010; //  246 : 250 - 0xfa
      10'hF7: dout <= 8'b11111010; //  247 : 250 - 0xfa
      10'hF8: dout <= 8'b11111010; //  248 : 250 - 0xfa
      10'hF9: dout <= 8'b11111010; //  249 : 250 - 0xfa
      10'hFA: dout <= 8'b11111010; //  250 : 250 - 0xfa
      10'hFB: dout <= 8'b11111010; //  251 : 250 - 0xfa
      10'hFC: dout <= 8'b11111010; //  252 : 250 - 0xfa
      10'hFD: dout <= 8'b11111010; //  253 : 250 - 0xfa
      10'hFE: dout <= 8'b11111010; //  254 : 250 - 0xfa
      10'hFF: dout <= 8'b11111010; //  255 : 250 - 0xfa
      10'h100: dout <= 8'b11111010; //  256 : 250 - 0xfa -- line 0x8
      10'h101: dout <= 8'b11111010; //  257 : 250 - 0xfa
      10'h102: dout <= 8'b11111010; //  258 : 250 - 0xfa
      10'h103: dout <= 8'b11111010; //  259 : 250 - 0xfa
      10'h104: dout <= 8'b11111010; //  260 : 250 - 0xfa
      10'h105: dout <= 8'b11111010; //  261 : 250 - 0xfa
      10'h106: dout <= 8'b11111010; //  262 : 250 - 0xfa
      10'h107: dout <= 8'b11111010; //  263 : 250 - 0xfa
      10'h108: dout <= 8'b11111010; //  264 : 250 - 0xfa
      10'h109: dout <= 8'b11111010; //  265 : 250 - 0xfa
      10'h10A: dout <= 8'b11111010; //  266 : 250 - 0xfa
      10'h10B: dout <= 8'b11101110; //  267 : 238 - 0xee
      10'h10C: dout <= 8'b11111010; //  268 : 250 - 0xfa
      10'h10D: dout <= 8'b11111010; //  269 : 250 - 0xfa
      10'h10E: dout <= 8'b11111010; //  270 : 250 - 0xfa
      10'h10F: dout <= 8'b11111010; //  271 : 250 - 0xfa
      10'h110: dout <= 8'b11111010; //  272 : 250 - 0xfa
      10'h111: dout <= 8'b11111010; //  273 : 250 - 0xfa
      10'h112: dout <= 8'b11111010; //  274 : 250 - 0xfa
      10'h113: dout <= 8'b11111010; //  275 : 250 - 0xfa
      10'h114: dout <= 8'b11101110; //  276 : 238 - 0xee
      10'h115: dout <= 8'b11111010; //  277 : 250 - 0xfa
      10'h116: dout <= 8'b11111010; //  278 : 250 - 0xfa
      10'h117: dout <= 8'b11111010; //  279 : 250 - 0xfa
      10'h118: dout <= 8'b11111010; //  280 : 250 - 0xfa
      10'h119: dout <= 8'b11111010; //  281 : 250 - 0xfa
      10'h11A: dout <= 8'b11111010; //  282 : 250 - 0xfa
      10'h11B: dout <= 8'b11111010; //  283 : 250 - 0xfa
      10'h11C: dout <= 8'b11111010; //  284 : 250 - 0xfa
      10'h11D: dout <= 8'b11111001; //  285 : 249 - 0xf9
      10'h11E: dout <= 8'b11111010; //  286 : 250 - 0xfa
      10'h11F: dout <= 8'b11111010; //  287 : 250 - 0xfa
      10'h120: dout <= 8'b11111010; //  288 : 250 - 0xfa -- line 0x9
      10'h121: dout <= 8'b11111010; //  289 : 250 - 0xfa
      10'h122: dout <= 8'b11111010; //  290 : 250 - 0xfa
      10'h123: dout <= 8'b11111010; //  291 : 250 - 0xfa
      10'h124: dout <= 8'b11111010; //  292 : 250 - 0xfa
      10'h125: dout <= 8'b11111010; //  293 : 250 - 0xfa
      10'h126: dout <= 8'b11111010; //  294 : 250 - 0xfa
      10'h127: dout <= 8'b11111010; //  295 : 250 - 0xfa
      10'h128: dout <= 8'b11111010; //  296 : 250 - 0xfa
      10'h129: dout <= 8'b11111010; //  297 : 250 - 0xfa
      10'h12A: dout <= 8'b11111010; //  298 : 250 - 0xfa
      10'h12B: dout <= 8'b11011101; //  299 : 221 - 0xdd
      10'h12C: dout <= 8'b11101101; //  300 : 237 - 0xed
      10'h12D: dout <= 8'b11101101; //  301 : 237 - 0xed
      10'h12E: dout <= 8'b11101101; //  302 : 237 - 0xed
      10'h12F: dout <= 8'b11101101; //  303 : 237 - 0xed
      10'h130: dout <= 8'b11101101; //  304 : 237 - 0xed
      10'h131: dout <= 8'b11101101; //  305 : 237 - 0xed
      10'h132: dout <= 8'b11101101; //  306 : 237 - 0xed
      10'h133: dout <= 8'b11101101; //  307 : 237 - 0xed
      10'h134: dout <= 8'b11011110; //  308 : 222 - 0xde
      10'h135: dout <= 8'b11111010; //  309 : 250 - 0xfa
      10'h136: dout <= 8'b11101010; //  310 : 234 - 0xea
      10'h137: dout <= 8'b11111010; //  311 : 250 - 0xfa
      10'h138: dout <= 8'b11111010; //  312 : 250 - 0xfa
      10'h139: dout <= 8'b11111010; //  313 : 250 - 0xfa
      10'h13A: dout <= 8'b11111010; //  314 : 250 - 0xfa
      10'h13B: dout <= 8'b11111010; //  315 : 250 - 0xfa
      10'h13C: dout <= 8'b11111010; //  316 : 250 - 0xfa
      10'h13D: dout <= 8'b11111010; //  317 : 250 - 0xfa
      10'h13E: dout <= 8'b11111010; //  318 : 250 - 0xfa
      10'h13F: dout <= 8'b11111010; //  319 : 250 - 0xfa
      10'h140: dout <= 8'b11111010; //  320 : 250 - 0xfa -- line 0xa
      10'h141: dout <= 8'b11111010; //  321 : 250 - 0xfa
      10'h142: dout <= 8'b11111010; //  322 : 250 - 0xfa
      10'h143: dout <= 8'b11111010; //  323 : 250 - 0xfa
      10'h144: dout <= 8'b11111010; //  324 : 250 - 0xfa
      10'h145: dout <= 8'b11111010; //  325 : 250 - 0xfa
      10'h146: dout <= 8'b11111010; //  326 : 250 - 0xfa
      10'h147: dout <= 8'b11111010; //  327 : 250 - 0xfa
      10'h148: dout <= 8'b11111010; //  328 : 250 - 0xfa
      10'h149: dout <= 8'b11111010; //  329 : 250 - 0xfa
      10'h14A: dout <= 8'b11111010; //  330 : 250 - 0xfa
      10'h14B: dout <= 8'b11111010; //  331 : 250 - 0xfa
      10'h14C: dout <= 8'b11111010; //  332 : 250 - 0xfa
      10'h14D: dout <= 8'b11111010; //  333 : 250 - 0xfa
      10'h14E: dout <= 8'b11111010; //  334 : 250 - 0xfa
      10'h14F: dout <= 8'b11111010; //  335 : 250 - 0xfa
      10'h150: dout <= 8'b11111010; //  336 : 250 - 0xfa
      10'h151: dout <= 8'b11111010; //  337 : 250 - 0xfa
      10'h152: dout <= 8'b11111010; //  338 : 250 - 0xfa
      10'h153: dout <= 8'b11111010; //  339 : 250 - 0xfa
      10'h154: dout <= 8'b11111010; //  340 : 250 - 0xfa
      10'h155: dout <= 8'b11111010; //  341 : 250 - 0xfa
      10'h156: dout <= 8'b11111010; //  342 : 250 - 0xfa
      10'h157: dout <= 8'b11111010; //  343 : 250 - 0xfa
      10'h158: dout <= 8'b11111010; //  344 : 250 - 0xfa
      10'h159: dout <= 8'b11111010; //  345 : 250 - 0xfa
      10'h15A: dout <= 8'b11111010; //  346 : 250 - 0xfa
      10'h15B: dout <= 8'b11111010; //  347 : 250 - 0xfa
      10'h15C: dout <= 8'b11111010; //  348 : 250 - 0xfa
      10'h15D: dout <= 8'b11111010; //  349 : 250 - 0xfa
      10'h15E: dout <= 8'b11111010; //  350 : 250 - 0xfa
      10'h15F: dout <= 8'b11111010; //  351 : 250 - 0xfa
      10'h160: dout <= 8'b11111010; //  352 : 250 - 0xfa -- line 0xb
      10'h161: dout <= 8'b11111010; //  353 : 250 - 0xfa
      10'h162: dout <= 8'b11111010; //  354 : 250 - 0xfa
      10'h163: dout <= 8'b11111010; //  355 : 250 - 0xfa
      10'h164: dout <= 8'b11111010; //  356 : 250 - 0xfa
      10'h165: dout <= 8'b11111010; //  357 : 250 - 0xfa
      10'h166: dout <= 8'b11111001; //  358 : 249 - 0xf9
      10'h167: dout <= 8'b11111010; //  359 : 250 - 0xfa
      10'h168: dout <= 8'b11111010; //  360 : 250 - 0xfa
      10'h169: dout <= 8'b11101010; //  361 : 234 - 0xea
      10'h16A: dout <= 8'b11111010; //  362 : 250 - 0xfa
      10'h16B: dout <= 8'b11111010; //  363 : 250 - 0xfa
      10'h16C: dout <= 8'b11111010; //  364 : 250 - 0xfa
      10'h16D: dout <= 8'b11111010; //  365 : 250 - 0xfa
      10'h16E: dout <= 8'b11111010; //  366 : 250 - 0xfa
      10'h16F: dout <= 8'b11111010; //  367 : 250 - 0xfa
      10'h170: dout <= 8'b11111010; //  368 : 250 - 0xfa
      10'h171: dout <= 8'b11111010; //  369 : 250 - 0xfa
      10'h172: dout <= 8'b11111010; //  370 : 250 - 0xfa
      10'h173: dout <= 8'b11111010; //  371 : 250 - 0xfa
      10'h174: dout <= 8'b11111010; //  372 : 250 - 0xfa
      10'h175: dout <= 8'b11111010; //  373 : 250 - 0xfa
      10'h176: dout <= 8'b11111010; //  374 : 250 - 0xfa
      10'h177: dout <= 8'b11111010; //  375 : 250 - 0xfa
      10'h178: dout <= 8'b11111010; //  376 : 250 - 0xfa
      10'h179: dout <= 8'b11111010; //  377 : 250 - 0xfa
      10'h17A: dout <= 8'b11111010; //  378 : 250 - 0xfa
      10'h17B: dout <= 8'b11111010; //  379 : 250 - 0xfa
      10'h17C: dout <= 8'b11111010; //  380 : 250 - 0xfa
      10'h17D: dout <= 8'b11111010; //  381 : 250 - 0xfa
      10'h17E: dout <= 8'b11111010; //  382 : 250 - 0xfa
      10'h17F: dout <= 8'b11111010; //  383 : 250 - 0xfa
      10'h180: dout <= 8'b11111010; //  384 : 250 - 0xfa -- line 0xc
      10'h181: dout <= 8'b11111010; //  385 : 250 - 0xfa
      10'h182: dout <= 8'b11101010; //  386 : 234 - 0xea
      10'h183: dout <= 8'b11111010; //  387 : 250 - 0xfa
      10'h184: dout <= 8'b11111010; //  388 : 250 - 0xfa
      10'h185: dout <= 8'b11111010; //  389 : 250 - 0xfa
      10'h186: dout <= 8'b11111010; //  390 : 250 - 0xfa
      10'h187: dout <= 8'b11111010; //  391 : 250 - 0xfa
      10'h188: dout <= 8'b11111010; //  392 : 250 - 0xfa
      10'h189: dout <= 8'b11111010; //  393 : 250 - 0xfa
      10'h18A: dout <= 8'b00100000; //  394 :  32 - 0x20
      10'h18B: dout <= 8'b00100010; //  395 :  34 - 0x22
      10'h18C: dout <= 8'b00010101; //  396 :  21 - 0x15
      10'h18D: dout <= 8'b00100011; //  397 :  35 - 0x23
      10'h18E: dout <= 8'b00100011; //  398 :  35 - 0x23
      10'h18F: dout <= 8'b11111010; //  399 : 250 - 0xfa
      10'h190: dout <= 8'b11111010; //  400 : 250 - 0xfa
      10'h191: dout <= 8'b00100011; //  401 :  35 - 0x23
      10'h192: dout <= 8'b00100100; //  402 :  36 - 0x24
      10'h193: dout <= 8'b00010001; //  403 :  17 - 0x11
      10'h194: dout <= 8'b00100010; //  404 :  34 - 0x22
      10'h195: dout <= 8'b00100100; //  405 :  36 - 0x24
      10'h196: dout <= 8'b11111010; //  406 : 250 - 0xfa
      10'h197: dout <= 8'b11111010; //  407 : 250 - 0xfa
      10'h198: dout <= 8'b11111010; //  408 : 250 - 0xfa
      10'h199: dout <= 8'b11111010; //  409 : 250 - 0xfa
      10'h19A: dout <= 8'b11111010; //  410 : 250 - 0xfa
      10'h19B: dout <= 8'b11101010; //  411 : 234 - 0xea
      10'h19C: dout <= 8'b11111010; //  412 : 250 - 0xfa
      10'h19D: dout <= 8'b11111010; //  413 : 250 - 0xfa
      10'h19E: dout <= 8'b11111010; //  414 : 250 - 0xfa
      10'h19F: dout <= 8'b11111010; //  415 : 250 - 0xfa
      10'h1A0: dout <= 8'b11111010; //  416 : 250 - 0xfa -- line 0xd
      10'h1A1: dout <= 8'b11111010; //  417 : 250 - 0xfa
      10'h1A2: dout <= 8'b11111010; //  418 : 250 - 0xfa
      10'h1A3: dout <= 8'b11111010; //  419 : 250 - 0xfa
      10'h1A4: dout <= 8'b11111010; //  420 : 250 - 0xfa
      10'h1A5: dout <= 8'b11111010; //  421 : 250 - 0xfa
      10'h1A6: dout <= 8'b11111010; //  422 : 250 - 0xfa
      10'h1A7: dout <= 8'b11111010; //  423 : 250 - 0xfa
      10'h1A8: dout <= 8'b11111010; //  424 : 250 - 0xfa
      10'h1A9: dout <= 8'b11111010; //  425 : 250 - 0xfa
      10'h1AA: dout <= 8'b11111010; //  426 : 250 - 0xfa
      10'h1AB: dout <= 8'b11111010; //  427 : 250 - 0xfa
      10'h1AC: dout <= 8'b11111010; //  428 : 250 - 0xfa
      10'h1AD: dout <= 8'b11111010; //  429 : 250 - 0xfa
      10'h1AE: dout <= 8'b11101010; //  430 : 234 - 0xea
      10'h1AF: dout <= 8'b11111010; //  431 : 250 - 0xfa
      10'h1B0: dout <= 8'b11111010; //  432 : 250 - 0xfa
      10'h1B1: dout <= 8'b11111010; //  433 : 250 - 0xfa
      10'h1B2: dout <= 8'b11111010; //  434 : 250 - 0xfa
      10'h1B3: dout <= 8'b11111010; //  435 : 250 - 0xfa
      10'h1B4: dout <= 8'b11111010; //  436 : 250 - 0xfa
      10'h1B5: dout <= 8'b11111010; //  437 : 250 - 0xfa
      10'h1B6: dout <= 8'b11111010; //  438 : 250 - 0xfa
      10'h1B7: dout <= 8'b11111010; //  439 : 250 - 0xfa
      10'h1B8: dout <= 8'b11111010; //  440 : 250 - 0xfa
      10'h1B9: dout <= 8'b11111010; //  441 : 250 - 0xfa
      10'h1BA: dout <= 8'b11111010; //  442 : 250 - 0xfa
      10'h1BB: dout <= 8'b11111010; //  443 : 250 - 0xfa
      10'h1BC: dout <= 8'b11111010; //  444 : 250 - 0xfa
      10'h1BD: dout <= 8'b11111010; //  445 : 250 - 0xfa
      10'h1BE: dout <= 8'b11111010; //  446 : 250 - 0xfa
      10'h1BF: dout <= 8'b11111010; //  447 : 250 - 0xfa
      10'h1C0: dout <= 8'b11111010; //  448 : 250 - 0xfa -- line 0xe
      10'h1C1: dout <= 8'b11111010; //  449 : 250 - 0xfa
      10'h1C2: dout <= 8'b11111010; //  450 : 250 - 0xfa
      10'h1C3: dout <= 8'b11111010; //  451 : 250 - 0xfa
      10'h1C4: dout <= 8'b11111010; //  452 : 250 - 0xfa
      10'h1C5: dout <= 8'b11111010; //  453 : 250 - 0xfa
      10'h1C6: dout <= 8'b11111010; //  454 : 250 - 0xfa
      10'h1C7: dout <= 8'b11111010; //  455 : 250 - 0xfa
      10'h1C8: dout <= 8'b11111001; //  456 : 249 - 0xf9
      10'h1C9: dout <= 8'b11111010; //  457 : 250 - 0xfa
      10'h1CA: dout <= 8'b11111010; //  458 : 250 - 0xfa
      10'h1CB: dout <= 8'b11111010; //  459 : 250 - 0xfa
      10'h1CC: dout <= 8'b00100100; //  460 :  36 - 0x24
      10'h1CD: dout <= 8'b00011111; //  461 :  31 - 0x1f
      10'h1CE: dout <= 8'b11111010; //  462 : 250 - 0xfa
      10'h1CF: dout <= 8'b11111010; //  463 : 250 - 0xfa
      10'h1D0: dout <= 8'b00100010; //  464 :  34 - 0x22
      10'h1D1: dout <= 8'b00010001; //  465 :  17 - 0x11
      10'h1D2: dout <= 8'b00010011; //  466 :  19 - 0x13
      10'h1D3: dout <= 8'b00010101; //  467 :  21 - 0x15
      10'h1D4: dout <= 8'b11111010; //  468 : 250 - 0xfa
      10'h1D5: dout <= 8'b11111010; //  469 : 250 - 0xfa
      10'h1D6: dout <= 8'b11111010; //  470 : 250 - 0xfa
      10'h1D7: dout <= 8'b11111010; //  471 : 250 - 0xfa
      10'h1D8: dout <= 8'b11111001; //  472 : 249 - 0xf9
      10'h1D9: dout <= 8'b11111010; //  473 : 250 - 0xfa
      10'h1DA: dout <= 8'b11111010; //  474 : 250 - 0xfa
      10'h1DB: dout <= 8'b11111010; //  475 : 250 - 0xfa
      10'h1DC: dout <= 8'b11111010; //  476 : 250 - 0xfa
      10'h1DD: dout <= 8'b11111010; //  477 : 250 - 0xfa
      10'h1DE: dout <= 8'b11111010; //  478 : 250 - 0xfa
      10'h1DF: dout <= 8'b11111010; //  479 : 250 - 0xfa
      10'h1E0: dout <= 8'b11111010; //  480 : 250 - 0xfa -- line 0xf
      10'h1E1: dout <= 8'b11111010; //  481 : 250 - 0xfa
      10'h1E2: dout <= 8'b11111010; //  482 : 250 - 0xfa
      10'h1E3: dout <= 8'b11111010; //  483 : 250 - 0xfa
      10'h1E4: dout <= 8'b11111010; //  484 : 250 - 0xfa
      10'h1E5: dout <= 8'b11111010; //  485 : 250 - 0xfa
      10'h1E6: dout <= 8'b11111010; //  486 : 250 - 0xfa
      10'h1E7: dout <= 8'b11111010; //  487 : 250 - 0xfa
      10'h1E8: dout <= 8'b11111010; //  488 : 250 - 0xfa
      10'h1E9: dout <= 8'b11111010; //  489 : 250 - 0xfa
      10'h1EA: dout <= 8'b11111010; //  490 : 250 - 0xfa
      10'h1EB: dout <= 8'b11111010; //  491 : 250 - 0xfa
      10'h1EC: dout <= 8'b11111010; //  492 : 250 - 0xfa
      10'h1ED: dout <= 8'b11111010; //  493 : 250 - 0xfa
      10'h1EE: dout <= 8'b11111010; //  494 : 250 - 0xfa
      10'h1EF: dout <= 8'b11111010; //  495 : 250 - 0xfa
      10'h1F0: dout <= 8'b11111010; //  496 : 250 - 0xfa
      10'h1F1: dout <= 8'b11111010; //  497 : 250 - 0xfa
      10'h1F2: dout <= 8'b11111010; //  498 : 250 - 0xfa
      10'h1F3: dout <= 8'b11111010; //  499 : 250 - 0xfa
      10'h1F4: dout <= 8'b11111010; //  500 : 250 - 0xfa
      10'h1F5: dout <= 8'b11111010; //  501 : 250 - 0xfa
      10'h1F6: dout <= 8'b11111010; //  502 : 250 - 0xfa
      10'h1F7: dout <= 8'b11111010; //  503 : 250 - 0xfa
      10'h1F8: dout <= 8'b11111010; //  504 : 250 - 0xfa
      10'h1F9: dout <= 8'b11111010; //  505 : 250 - 0xfa
      10'h1FA: dout <= 8'b11111010; //  506 : 250 - 0xfa
      10'h1FB: dout <= 8'b11111010; //  507 : 250 - 0xfa
      10'h1FC: dout <= 8'b11111010; //  508 : 250 - 0xfa
      10'h1FD: dout <= 8'b11111010; //  509 : 250 - 0xfa
      10'h1FE: dout <= 8'b11111010; //  510 : 250 - 0xfa
      10'h1FF: dout <= 8'b11111010; //  511 : 250 - 0xfa
      10'h200: dout <= 8'b11111010; //  512 : 250 - 0xfa -- line 0x10
      10'h201: dout <= 8'b11111010; //  513 : 250 - 0xfa
      10'h202: dout <= 8'b11111010; //  514 : 250 - 0xfa
      10'h203: dout <= 8'b11111010; //  515 : 250 - 0xfa
      10'h204: dout <= 8'b11111010; //  516 : 250 - 0xfa
      10'h205: dout <= 8'b11111010; //  517 : 250 - 0xfa
      10'h206: dout <= 8'b11111010; //  518 : 250 - 0xfa
      10'h207: dout <= 8'b11111010; //  519 : 250 - 0xfa
      10'h208: dout <= 8'b11111010; //  520 : 250 - 0xfa
      10'h209: dout <= 8'b11111010; //  521 : 250 - 0xfa
      10'h20A: dout <= 8'b11111010; //  522 : 250 - 0xfa
      10'h20B: dout <= 8'b11111010; //  523 : 250 - 0xfa
      10'h20C: dout <= 8'b11111010; //  524 : 250 - 0xfa
      10'h20D: dout <= 8'b11111010; //  525 : 250 - 0xfa
      10'h20E: dout <= 8'b11111010; //  526 : 250 - 0xfa
      10'h20F: dout <= 8'b11111010; //  527 : 250 - 0xfa
      10'h210: dout <= 8'b11111010; //  528 : 250 - 0xfa
      10'h211: dout <= 8'b11111010; //  529 : 250 - 0xfa
      10'h212: dout <= 8'b11111010; //  530 : 250 - 0xfa
      10'h213: dout <= 8'b11111010; //  531 : 250 - 0xfa
      10'h214: dout <= 8'b11111010; //  532 : 250 - 0xfa
      10'h215: dout <= 8'b11111010; //  533 : 250 - 0xfa
      10'h216: dout <= 8'b11111010; //  534 : 250 - 0xfa
      10'h217: dout <= 8'b11111010; //  535 : 250 - 0xfa
      10'h218: dout <= 8'b11101001; //  536 : 233 - 0xe9
      10'h219: dout <= 8'b11111010; //  537 : 250 - 0xfa
      10'h21A: dout <= 8'b11111010; //  538 : 250 - 0xfa
      10'h21B: dout <= 8'b11111001; //  539 : 249 - 0xf9
      10'h21C: dout <= 8'b11111010; //  540 : 250 - 0xfa
      10'h21D: dout <= 8'b11111010; //  541 : 250 - 0xfa
      10'h21E: dout <= 8'b11111010; //  542 : 250 - 0xfa
      10'h21F: dout <= 8'b11111010; //  543 : 250 - 0xfa
      10'h220: dout <= 8'b11111010; //  544 : 250 - 0xfa -- line 0x11
      10'h221: dout <= 8'b11111010; //  545 : 250 - 0xfa
      10'h222: dout <= 8'b11111010; //  546 : 250 - 0xfa
      10'h223: dout <= 8'b11111010; //  547 : 250 - 0xfa
      10'h224: dout <= 8'b11111001; //  548 : 249 - 0xf9
      10'h225: dout <= 8'b11111010; //  549 : 250 - 0xfa
      10'h226: dout <= 8'b00101100; //  550 :  44 - 0x2c
      10'h227: dout <= 8'b00100100; //  551 :  36 - 0x24
      10'h228: dout <= 8'b00100010; //  552 :  34 - 0x22
      10'h229: dout <= 8'b00010001; //  553 :  17 - 0x11
      10'h22A: dout <= 8'b00010011; //  554 :  19 - 0x13
      10'h22B: dout <= 8'b00011011; //  555 :  27 - 0x1b
      10'h22C: dout <= 8'b00101101; //  556 :  45 - 0x2d
      10'h22D: dout <= 8'b11111010; //  557 : 250 - 0xfa
      10'h22E: dout <= 8'b11111001; //  558 : 249 - 0xf9
      10'h22F: dout <= 8'b11111010; //  559 : 250 - 0xfa
      10'h230: dout <= 8'b11111010; //  560 : 250 - 0xfa
      10'h231: dout <= 8'b11111010; //  561 : 250 - 0xfa
      10'h232: dout <= 8'b11111010; //  562 : 250 - 0xfa
      10'h233: dout <= 8'b00000001; //  563 :   1 - 0x1
      10'h234: dout <= 8'b11111010; //  564 : 250 - 0xfa
      10'h235: dout <= 8'b11111010; //  565 : 250 - 0xfa
      10'h236: dout <= 8'b11111010; //  566 : 250 - 0xfa
      10'h237: dout <= 8'b11111010; //  567 : 250 - 0xfa
      10'h238: dout <= 8'b11111010; //  568 : 250 - 0xfa
      10'h239: dout <= 8'b11111010; //  569 : 250 - 0xfa
      10'h23A: dout <= 8'b11111010; //  570 : 250 - 0xfa
      10'h23B: dout <= 8'b11111010; //  571 : 250 - 0xfa
      10'h23C: dout <= 8'b11111010; //  572 : 250 - 0xfa
      10'h23D: dout <= 8'b11111010; //  573 : 250 - 0xfa
      10'h23E: dout <= 8'b11111010; //  574 : 250 - 0xfa
      10'h23F: dout <= 8'b11111010; //  575 : 250 - 0xfa
      10'h240: dout <= 8'b11111010; //  576 : 250 - 0xfa -- line 0x12
      10'h241: dout <= 8'b11111010; //  577 : 250 - 0xfa
      10'h242: dout <= 8'b11111010; //  578 : 250 - 0xfa
      10'h243: dout <= 8'b11111010; //  579 : 250 - 0xfa
      10'h244: dout <= 8'b11111010; //  580 : 250 - 0xfa
      10'h245: dout <= 8'b11111010; //  581 : 250 - 0xfa
      10'h246: dout <= 8'b11101001; //  582 : 233 - 0xe9
      10'h247: dout <= 8'b11111010; //  583 : 250 - 0xfa
      10'h248: dout <= 8'b11111010; //  584 : 250 - 0xfa
      10'h249: dout <= 8'b11111001; //  585 : 249 - 0xf9
      10'h24A: dout <= 8'b11111010; //  586 : 250 - 0xfa
      10'h24B: dout <= 8'b11111010; //  587 : 250 - 0xfa
      10'h24C: dout <= 8'b11111010; //  588 : 250 - 0xfa
      10'h24D: dout <= 8'b11111010; //  589 : 250 - 0xfa
      10'h24E: dout <= 8'b11111010; //  590 : 250 - 0xfa
      10'h24F: dout <= 8'b11111010; //  591 : 250 - 0xfa
      10'h250: dout <= 8'b11111010; //  592 : 250 - 0xfa
      10'h251: dout <= 8'b11111010; //  593 : 250 - 0xfa
      10'h252: dout <= 8'b11111010; //  594 : 250 - 0xfa
      10'h253: dout <= 8'b11111010; //  595 : 250 - 0xfa
      10'h254: dout <= 8'b11111010; //  596 : 250 - 0xfa
      10'h255: dout <= 8'b11111010; //  597 : 250 - 0xfa
      10'h256: dout <= 8'b11111010; //  598 : 250 - 0xfa
      10'h257: dout <= 8'b11111010; //  599 : 250 - 0xfa
      10'h258: dout <= 8'b11111010; //  600 : 250 - 0xfa
      10'h259: dout <= 8'b11111010; //  601 : 250 - 0xfa
      10'h25A: dout <= 8'b11111010; //  602 : 250 - 0xfa
      10'h25B: dout <= 8'b11111010; //  603 : 250 - 0xfa
      10'h25C: dout <= 8'b11111010; //  604 : 250 - 0xfa
      10'h25D: dout <= 8'b11111010; //  605 : 250 - 0xfa
      10'h25E: dout <= 8'b11111010; //  606 : 250 - 0xfa
      10'h25F: dout <= 8'b11111010; //  607 : 250 - 0xfa
      10'h260: dout <= 8'b11111010; //  608 : 250 - 0xfa -- line 0x13
      10'h261: dout <= 8'b11111010; //  609 : 250 - 0xfa
      10'h262: dout <= 8'b11111010; //  610 : 250 - 0xfa
      10'h263: dout <= 8'b11111010; //  611 : 250 - 0xfa
      10'h264: dout <= 8'b11111010; //  612 : 250 - 0xfa
      10'h265: dout <= 8'b11111010; //  613 : 250 - 0xfa
      10'h266: dout <= 8'b11111010; //  614 : 250 - 0xfa
      10'h267: dout <= 8'b00010100; //  615 :  20 - 0x14
      10'h268: dout <= 8'b00011001; //  616 :  25 - 0x19
      10'h269: dout <= 8'b00010110; //  617 :  22 - 0x16
      10'h26A: dout <= 8'b00010110; //  618 :  22 - 0x16
      10'h26B: dout <= 8'b00011001; //  619 :  25 - 0x19
      10'h26C: dout <= 8'b00010011; //  620 :  19 - 0x13
      10'h26D: dout <= 8'b00100101; //  621 :  37 - 0x25
      10'h26E: dout <= 8'b00011100; //  622 :  28 - 0x1c
      10'h26F: dout <= 8'b00100100; //  623 :  36 - 0x24
      10'h270: dout <= 8'b00101001; //  624 :  41 - 0x29
      10'h271: dout <= 8'b00101101; //  625 :  45 - 0x2d
      10'h272: dout <= 8'b11111010; //  626 : 250 - 0xfa
      10'h273: dout <= 8'b00011000; //  627 :  24 - 0x18
      10'h274: dout <= 8'b00010001; //  628 :  17 - 0x11
      10'h275: dout <= 8'b00100010; //  629 :  34 - 0x22
      10'h276: dout <= 8'b00010100; //  630 :  20 - 0x14
      10'h277: dout <= 8'b11111010; //  631 : 250 - 0xfa
      10'h278: dout <= 8'b11111010; //  632 : 250 - 0xfa
      10'h279: dout <= 8'b11111010; //  633 : 250 - 0xfa
      10'h27A: dout <= 8'b11111010; //  634 : 250 - 0xfa
      10'h27B: dout <= 8'b11111010; //  635 : 250 - 0xfa
      10'h27C: dout <= 8'b11111010; //  636 : 250 - 0xfa
      10'h27D: dout <= 8'b11111010; //  637 : 250 - 0xfa
      10'h27E: dout <= 8'b11111001; //  638 : 249 - 0xf9
      10'h27F: dout <= 8'b11111010; //  639 : 250 - 0xfa
      10'h280: dout <= 8'b11111010; //  640 : 250 - 0xfa -- line 0x14
      10'h281: dout <= 8'b11111010; //  641 : 250 - 0xfa
      10'h282: dout <= 8'b11101001; //  642 : 233 - 0xe9
      10'h283: dout <= 8'b11111010; //  643 : 250 - 0xfa
      10'h284: dout <= 8'b11111010; //  644 : 250 - 0xfa
      10'h285: dout <= 8'b11111010; //  645 : 250 - 0xfa
      10'h286: dout <= 8'b11111010; //  646 : 250 - 0xfa
      10'h287: dout <= 8'b11111001; //  647 : 249 - 0xf9
      10'h288: dout <= 8'b11111001; //  648 : 249 - 0xf9
      10'h289: dout <= 8'b11111010; //  649 : 250 - 0xfa
      10'h28A: dout <= 8'b11111010; //  650 : 250 - 0xfa
      10'h28B: dout <= 8'b11111010; //  651 : 250 - 0xfa
      10'h28C: dout <= 8'b11111010; //  652 : 250 - 0xfa
      10'h28D: dout <= 8'b11111010; //  653 : 250 - 0xfa
      10'h28E: dout <= 8'b11111010; //  654 : 250 - 0xfa
      10'h28F: dout <= 8'b11111010; //  655 : 250 - 0xfa
      10'h290: dout <= 8'b11111010; //  656 : 250 - 0xfa
      10'h291: dout <= 8'b11111010; //  657 : 250 - 0xfa
      10'h292: dout <= 8'b11111010; //  658 : 250 - 0xfa
      10'h293: dout <= 8'b11101001; //  659 : 233 - 0xe9
      10'h294: dout <= 8'b11111010; //  660 : 250 - 0xfa
      10'h295: dout <= 8'b11111010; //  661 : 250 - 0xfa
      10'h296: dout <= 8'b11111010; //  662 : 250 - 0xfa
      10'h297: dout <= 8'b11111010; //  663 : 250 - 0xfa
      10'h298: dout <= 8'b11101010; //  664 : 234 - 0xea
      10'h299: dout <= 8'b11111010; //  665 : 250 - 0xfa
      10'h29A: dout <= 8'b11111010; //  666 : 250 - 0xfa
      10'h29B: dout <= 8'b11111010; //  667 : 250 - 0xfa
      10'h29C: dout <= 8'b11111010; //  668 : 250 - 0xfa
      10'h29D: dout <= 8'b11111010; //  669 : 250 - 0xfa
      10'h29E: dout <= 8'b11111010; //  670 : 250 - 0xfa
      10'h29F: dout <= 8'b11111010; //  671 : 250 - 0xfa
      10'h2A0: dout <= 8'b11111010; //  672 : 250 - 0xfa -- line 0x15
      10'h2A1: dout <= 8'b11111010; //  673 : 250 - 0xfa
      10'h2A2: dout <= 8'b11111010; //  674 : 250 - 0xfa
      10'h2A3: dout <= 8'b11111010; //  675 : 250 - 0xfa
      10'h2A4: dout <= 8'b11111010; //  676 : 250 - 0xfa
      10'h2A5: dout <= 8'b11111010; //  677 : 250 - 0xfa
      10'h2A6: dout <= 8'b11111010; //  678 : 250 - 0xfa
      10'h2A7: dout <= 8'b00011100; //  679 :  28 - 0x1c
      10'h2A8: dout <= 8'b00010001; //  680 :  17 - 0x11
      10'h2A9: dout <= 8'b00100000; //  681 :  32 - 0x20
      10'h2AA: dout <= 8'b00100011; //  682 :  35 - 0x23
      10'h2AB: dout <= 8'b00101101; //  683 :  45 - 0x2d
      10'h2AC: dout <= 8'b11111010; //  684 : 250 - 0xfa
      10'h2AD: dout <= 8'b11111010; //  685 : 250 - 0xfa
      10'h2AE: dout <= 8'b11111010; //  686 : 250 - 0xfa
      10'h2AF: dout <= 8'b11101010; //  687 : 234 - 0xea
      10'h2B0: dout <= 8'b11111010; //  688 : 250 - 0xfa
      10'h2B1: dout <= 8'b11111010; //  689 : 250 - 0xfa
      10'h2B2: dout <= 8'b11111010; //  690 : 250 - 0xfa
      10'h2B3: dout <= 8'b00000011; //  691 :   3 - 0x3
      10'h2B4: dout <= 8'b11111010; //  692 : 250 - 0xfa
      10'h2B5: dout <= 8'b11111010; //  693 : 250 - 0xfa
      10'h2B6: dout <= 8'b11111010; //  694 : 250 - 0xfa
      10'h2B7: dout <= 8'b11111010; //  695 : 250 - 0xfa
      10'h2B8: dout <= 8'b11111010; //  696 : 250 - 0xfa
      10'h2B9: dout <= 8'b11111010; //  697 : 250 - 0xfa
      10'h2BA: dout <= 8'b11111010; //  698 : 250 - 0xfa
      10'h2BB: dout <= 8'b11111010; //  699 : 250 - 0xfa
      10'h2BC: dout <= 8'b11111010; //  700 : 250 - 0xfa
      10'h2BD: dout <= 8'b11111010; //  701 : 250 - 0xfa
      10'h2BE: dout <= 8'b11111010; //  702 : 250 - 0xfa
      10'h2BF: dout <= 8'b11111010; //  703 : 250 - 0xfa
      10'h2C0: dout <= 8'b11111010; //  704 : 250 - 0xfa -- line 0x16
      10'h2C1: dout <= 8'b11111010; //  705 : 250 - 0xfa
      10'h2C2: dout <= 8'b11111010; //  706 : 250 - 0xfa
      10'h2C3: dout <= 8'b11111010; //  707 : 250 - 0xfa
      10'h2C4: dout <= 8'b11111010; //  708 : 250 - 0xfa
      10'h2C5: dout <= 8'b11111010; //  709 : 250 - 0xfa
      10'h2C6: dout <= 8'b11111010; //  710 : 250 - 0xfa
      10'h2C7: dout <= 8'b11111010; //  711 : 250 - 0xfa
      10'h2C8: dout <= 8'b11111010; //  712 : 250 - 0xfa
      10'h2C9: dout <= 8'b11111010; //  713 : 250 - 0xfa
      10'h2CA: dout <= 8'b11111010; //  714 : 250 - 0xfa
      10'h2CB: dout <= 8'b11111010; //  715 : 250 - 0xfa
      10'h2CC: dout <= 8'b11111010; //  716 : 250 - 0xfa
      10'h2CD: dout <= 8'b11111010; //  717 : 250 - 0xfa
      10'h2CE: dout <= 8'b11111010; //  718 : 250 - 0xfa
      10'h2CF: dout <= 8'b11111010; //  719 : 250 - 0xfa
      10'h2D0: dout <= 8'b11111010; //  720 : 250 - 0xfa
      10'h2D1: dout <= 8'b11111010; //  721 : 250 - 0xfa
      10'h2D2: dout <= 8'b11111010; //  722 : 250 - 0xfa
      10'h2D3: dout <= 8'b11111010; //  723 : 250 - 0xfa
      10'h2D4: dout <= 8'b11111010; //  724 : 250 - 0xfa
      10'h2D5: dout <= 8'b11111010; //  725 : 250 - 0xfa
      10'h2D6: dout <= 8'b11111010; //  726 : 250 - 0xfa
      10'h2D7: dout <= 8'b11111010; //  727 : 250 - 0xfa
      10'h2D8: dout <= 8'b11111010; //  728 : 250 - 0xfa
      10'h2D9: dout <= 8'b11111010; //  729 : 250 - 0xfa
      10'h2DA: dout <= 8'b11111010; //  730 : 250 - 0xfa
      10'h2DB: dout <= 8'b11111010; //  731 : 250 - 0xfa
      10'h2DC: dout <= 8'b11111010; //  732 : 250 - 0xfa
      10'h2DD: dout <= 8'b11101010; //  733 : 234 - 0xea
      10'h2DE: dout <= 8'b11111010; //  734 : 250 - 0xfa
      10'h2DF: dout <= 8'b11111010; //  735 : 250 - 0xfa
      10'h2E0: dout <= 8'b11111011; //  736 : 251 - 0xfb -- line 0x17
      10'h2E1: dout <= 8'b11111011; //  737 : 251 - 0xfb
      10'h2E2: dout <= 8'b11111011; //  738 : 251 - 0xfb
      10'h2E3: dout <= 8'b11111011; //  739 : 251 - 0xfb
      10'h2E4: dout <= 8'b11111011; //  740 : 251 - 0xfb
      10'h2E5: dout <= 8'b11111011; //  741 : 251 - 0xfb
      10'h2E6: dout <= 8'b11111011; //  742 : 251 - 0xfb
      10'h2E7: dout <= 8'b11111011; //  743 : 251 - 0xfb
      10'h2E8: dout <= 8'b11111011; //  744 : 251 - 0xfb
      10'h2E9: dout <= 8'b11111011; //  745 : 251 - 0xfb
      10'h2EA: dout <= 8'b11111011; //  746 : 251 - 0xfb
      10'h2EB: dout <= 8'b11111011; //  747 : 251 - 0xfb
      10'h2EC: dout <= 8'b11111011; //  748 : 251 - 0xfb
      10'h2ED: dout <= 8'b11111011; //  749 : 251 - 0xfb
      10'h2EE: dout <= 8'b11111011; //  750 : 251 - 0xfb
      10'h2EF: dout <= 8'b11111011; //  751 : 251 - 0xfb
      10'h2F0: dout <= 8'b11111011; //  752 : 251 - 0xfb
      10'h2F1: dout <= 8'b11111011; //  753 : 251 - 0xfb
      10'h2F2: dout <= 8'b11111011; //  754 : 251 - 0xfb
      10'h2F3: dout <= 8'b11111011; //  755 : 251 - 0xfb
      10'h2F4: dout <= 8'b11111011; //  756 : 251 - 0xfb
      10'h2F5: dout <= 8'b11111011; //  757 : 251 - 0xfb
      10'h2F6: dout <= 8'b11111011; //  758 : 251 - 0xfb
      10'h2F7: dout <= 8'b11111011; //  759 : 251 - 0xfb
      10'h2F8: dout <= 8'b11111011; //  760 : 251 - 0xfb
      10'h2F9: dout <= 8'b11111011; //  761 : 251 - 0xfb
      10'h2FA: dout <= 8'b11111011; //  762 : 251 - 0xfb
      10'h2FB: dout <= 8'b11111011; //  763 : 251 - 0xfb
      10'h2FC: dout <= 8'b11111011; //  764 : 251 - 0xfb
      10'h2FD: dout <= 8'b11111011; //  765 : 251 - 0xfb
      10'h2FE: dout <= 8'b11111011; //  766 : 251 - 0xfb
      10'h2FF: dout <= 8'b11111011; //  767 : 251 - 0xfb
      10'h300: dout <= 8'b11111111; //  768 : 255 - 0xff -- line 0x18
      10'h301: dout <= 8'b11111111; //  769 : 255 - 0xff
      10'h302: dout <= 8'b11111111; //  770 : 255 - 0xff
      10'h303: dout <= 8'b11111111; //  771 : 255 - 0xff
      10'h304: dout <= 8'b11111111; //  772 : 255 - 0xff
      10'h305: dout <= 8'b11111111; //  773 : 255 - 0xff
      10'h306: dout <= 8'b11111111; //  774 : 255 - 0xff
      10'h307: dout <= 8'b11111111; //  775 : 255 - 0xff
      10'h308: dout <= 8'b11111111; //  776 : 255 - 0xff
      10'h309: dout <= 8'b11111111; //  777 : 255 - 0xff
      10'h30A: dout <= 8'b11111111; //  778 : 255 - 0xff
      10'h30B: dout <= 8'b11111111; //  779 : 255 - 0xff
      10'h30C: dout <= 8'b11111111; //  780 : 255 - 0xff
      10'h30D: dout <= 8'b11111111; //  781 : 255 - 0xff
      10'h30E: dout <= 8'b11111111; //  782 : 255 - 0xff
      10'h30F: dout <= 8'b11111111; //  783 : 255 - 0xff
      10'h310: dout <= 8'b11111111; //  784 : 255 - 0xff
      10'h311: dout <= 8'b11111111; //  785 : 255 - 0xff
      10'h312: dout <= 8'b11111111; //  786 : 255 - 0xff
      10'h313: dout <= 8'b11111111; //  787 : 255 - 0xff
      10'h314: dout <= 8'b11111111; //  788 : 255 - 0xff
      10'h315: dout <= 8'b11111111; //  789 : 255 - 0xff
      10'h316: dout <= 8'b11111111; //  790 : 255 - 0xff
      10'h317: dout <= 8'b11111111; //  791 : 255 - 0xff
      10'h318: dout <= 8'b11111111; //  792 : 255 - 0xff
      10'h319: dout <= 8'b11111111; //  793 : 255 - 0xff
      10'h31A: dout <= 8'b11111111; //  794 : 255 - 0xff
      10'h31B: dout <= 8'b11111111; //  795 : 255 - 0xff
      10'h31C: dout <= 8'b11111111; //  796 : 255 - 0xff
      10'h31D: dout <= 8'b11111111; //  797 : 255 - 0xff
      10'h31E: dout <= 8'b11111111; //  798 : 255 - 0xff
      10'h31F: dout <= 8'b11111111; //  799 : 255 - 0xff
      10'h320: dout <= 8'b11111111; //  800 : 255 - 0xff -- line 0x19
      10'h321: dout <= 8'b11111101; //  801 : 253 - 0xfd
      10'h322: dout <= 8'b11111111; //  802 : 255 - 0xff
      10'h323: dout <= 8'b11111101; //  803 : 253 - 0xfd
      10'h324: dout <= 8'b11111111; //  804 : 255 - 0xff
      10'h325: dout <= 8'b11111101; //  805 : 253 - 0xfd
      10'h326: dout <= 8'b11111111; //  806 : 255 - 0xff
      10'h327: dout <= 8'b11111101; //  807 : 253 - 0xfd
      10'h328: dout <= 8'b11111111; //  808 : 255 - 0xff
      10'h329: dout <= 8'b11111101; //  809 : 253 - 0xfd
      10'h32A: dout <= 8'b11111111; //  810 : 255 - 0xff
      10'h32B: dout <= 8'b11111101; //  811 : 253 - 0xfd
      10'h32C: dout <= 8'b11111111; //  812 : 255 - 0xff
      10'h32D: dout <= 8'b11111101; //  813 : 253 - 0xfd
      10'h32E: dout <= 8'b11111111; //  814 : 255 - 0xff
      10'h32F: dout <= 8'b11111101; //  815 : 253 - 0xfd
      10'h330: dout <= 8'b11111111; //  816 : 255 - 0xff
      10'h331: dout <= 8'b11111101; //  817 : 253 - 0xfd
      10'h332: dout <= 8'b11111111; //  818 : 255 - 0xff
      10'h333: dout <= 8'b11111101; //  819 : 253 - 0xfd
      10'h334: dout <= 8'b11111111; //  820 : 255 - 0xff
      10'h335: dout <= 8'b11111101; //  821 : 253 - 0xfd
      10'h336: dout <= 8'b11111111; //  822 : 255 - 0xff
      10'h337: dout <= 8'b11111101; //  823 : 253 - 0xfd
      10'h338: dout <= 8'b11111111; //  824 : 255 - 0xff
      10'h339: dout <= 8'b11111101; //  825 : 253 - 0xfd
      10'h33A: dout <= 8'b11111111; //  826 : 255 - 0xff
      10'h33B: dout <= 8'b11111101; //  827 : 253 - 0xfd
      10'h33C: dout <= 8'b11111111; //  828 : 255 - 0xff
      10'h33D: dout <= 8'b11111101; //  829 : 253 - 0xfd
      10'h33E: dout <= 8'b11111111; //  830 : 255 - 0xff
      10'h33F: dout <= 8'b11111101; //  831 : 253 - 0xfd
      10'h340: dout <= 8'b11111111; //  832 : 255 - 0xff -- line 0x1a
      10'h341: dout <= 8'b11111101; //  833 : 253 - 0xfd
      10'h342: dout <= 8'b11111111; //  834 : 255 - 0xff
      10'h343: dout <= 8'b11111101; //  835 : 253 - 0xfd
      10'h344: dout <= 8'b11111111; //  836 : 255 - 0xff
      10'h345: dout <= 8'b11111101; //  837 : 253 - 0xfd
      10'h346: dout <= 8'b11111111; //  838 : 255 - 0xff
      10'h347: dout <= 8'b11111101; //  839 : 253 - 0xfd
      10'h348: dout <= 8'b11111111; //  840 : 255 - 0xff
      10'h349: dout <= 8'b11111101; //  841 : 253 - 0xfd
      10'h34A: dout <= 8'b11111111; //  842 : 255 - 0xff
      10'h34B: dout <= 8'b11111101; //  843 : 253 - 0xfd
      10'h34C: dout <= 8'b11111111; //  844 : 255 - 0xff
      10'h34D: dout <= 8'b11111101; //  845 : 253 - 0xfd
      10'h34E: dout <= 8'b11111111; //  846 : 255 - 0xff
      10'h34F: dout <= 8'b11111101; //  847 : 253 - 0xfd
      10'h350: dout <= 8'b11111111; //  848 : 255 - 0xff
      10'h351: dout <= 8'b11111101; //  849 : 253 - 0xfd
      10'h352: dout <= 8'b11111111; //  850 : 255 - 0xff
      10'h353: dout <= 8'b11111101; //  851 : 253 - 0xfd
      10'h354: dout <= 8'b11111111; //  852 : 255 - 0xff
      10'h355: dout <= 8'b11111101; //  853 : 253 - 0xfd
      10'h356: dout <= 8'b11111111; //  854 : 255 - 0xff
      10'h357: dout <= 8'b11111101; //  855 : 253 - 0xfd
      10'h358: dout <= 8'b11111111; //  856 : 255 - 0xff
      10'h359: dout <= 8'b11111101; //  857 : 253 - 0xfd
      10'h35A: dout <= 8'b11111111; //  858 : 255 - 0xff
      10'h35B: dout <= 8'b11111101; //  859 : 253 - 0xfd
      10'h35C: dout <= 8'b11111111; //  860 : 255 - 0xff
      10'h35D: dout <= 8'b11111101; //  861 : 253 - 0xfd
      10'h35E: dout <= 8'b11111111; //  862 : 255 - 0xff
      10'h35F: dout <= 8'b11111101; //  863 : 253 - 0xfd
      10'h360: dout <= 8'b11111111; //  864 : 255 - 0xff -- line 0x1b
      10'h361: dout <= 8'b11111111; //  865 : 255 - 0xff
      10'h362: dout <= 8'b11111111; //  866 : 255 - 0xff
      10'h363: dout <= 8'b11111111; //  867 : 255 - 0xff
      10'h364: dout <= 8'b11111111; //  868 : 255 - 0xff
      10'h365: dout <= 8'b11111111; //  869 : 255 - 0xff
      10'h366: dout <= 8'b11111111; //  870 : 255 - 0xff
      10'h367: dout <= 8'b11111111; //  871 : 255 - 0xff
      10'h368: dout <= 8'b11111111; //  872 : 255 - 0xff
      10'h369: dout <= 8'b11111111; //  873 : 255 - 0xff
      10'h36A: dout <= 8'b11111111; //  874 : 255 - 0xff
      10'h36B: dout <= 8'b11111111; //  875 : 255 - 0xff
      10'h36C: dout <= 8'b11111111; //  876 : 255 - 0xff
      10'h36D: dout <= 8'b11111111; //  877 : 255 - 0xff
      10'h36E: dout <= 8'b11111111; //  878 : 255 - 0xff
      10'h36F: dout <= 8'b11111111; //  879 : 255 - 0xff
      10'h370: dout <= 8'b11111111; //  880 : 255 - 0xff
      10'h371: dout <= 8'b11111111; //  881 : 255 - 0xff
      10'h372: dout <= 8'b11111111; //  882 : 255 - 0xff
      10'h373: dout <= 8'b11111111; //  883 : 255 - 0xff
      10'h374: dout <= 8'b11111111; //  884 : 255 - 0xff
      10'h375: dout <= 8'b11111111; //  885 : 255 - 0xff
      10'h376: dout <= 8'b11111111; //  886 : 255 - 0xff
      10'h377: dout <= 8'b11111111; //  887 : 255 - 0xff
      10'h378: dout <= 8'b11111111; //  888 : 255 - 0xff
      10'h379: dout <= 8'b11111111; //  889 : 255 - 0xff
      10'h37A: dout <= 8'b11111111; //  890 : 255 - 0xff
      10'h37B: dout <= 8'b11111111; //  891 : 255 - 0xff
      10'h37C: dout <= 8'b11111111; //  892 : 255 - 0xff
      10'h37D: dout <= 8'b11111111; //  893 : 255 - 0xff
      10'h37E: dout <= 8'b11111111; //  894 : 255 - 0xff
      10'h37F: dout <= 8'b11111111; //  895 : 255 - 0xff
      10'h380: dout <= 8'b11101011; //  896 : 235 - 0xeb -- line 0x1c
      10'h381: dout <= 8'b11101011; //  897 : 235 - 0xeb
      10'h382: dout <= 8'b11101011; //  898 : 235 - 0xeb
      10'h383: dout <= 8'b11101011; //  899 : 235 - 0xeb
      10'h384: dout <= 8'b11101011; //  900 : 235 - 0xeb
      10'h385: dout <= 8'b11101011; //  901 : 235 - 0xeb
      10'h386: dout <= 8'b11101011; //  902 : 235 - 0xeb
      10'h387: dout <= 8'b11101011; //  903 : 235 - 0xeb
      10'h388: dout <= 8'b11101011; //  904 : 235 - 0xeb
      10'h389: dout <= 8'b11101011; //  905 : 235 - 0xeb
      10'h38A: dout <= 8'b11101011; //  906 : 235 - 0xeb
      10'h38B: dout <= 8'b11101011; //  907 : 235 - 0xeb
      10'h38C: dout <= 8'b11101011; //  908 : 235 - 0xeb
      10'h38D: dout <= 8'b11101011; //  909 : 235 - 0xeb
      10'h38E: dout <= 8'b11101011; //  910 : 235 - 0xeb
      10'h38F: dout <= 8'b11101011; //  911 : 235 - 0xeb
      10'h390: dout <= 8'b11101011; //  912 : 235 - 0xeb
      10'h391: dout <= 8'b11101011; //  913 : 235 - 0xeb
      10'h392: dout <= 8'b11101011; //  914 : 235 - 0xeb
      10'h393: dout <= 8'b11101011; //  915 : 235 - 0xeb
      10'h394: dout <= 8'b11101011; //  916 : 235 - 0xeb
      10'h395: dout <= 8'b11101011; //  917 : 235 - 0xeb
      10'h396: dout <= 8'b11101011; //  918 : 235 - 0xeb
      10'h397: dout <= 8'b11101011; //  919 : 235 - 0xeb
      10'h398: dout <= 8'b11101011; //  920 : 235 - 0xeb
      10'h399: dout <= 8'b11101011; //  921 : 235 - 0xeb
      10'h39A: dout <= 8'b11101011; //  922 : 235 - 0xeb
      10'h39B: dout <= 8'b11101011; //  923 : 235 - 0xeb
      10'h39C: dout <= 8'b11101011; //  924 : 235 - 0xeb
      10'h39D: dout <= 8'b11101011; //  925 : 235 - 0xeb
      10'h39E: dout <= 8'b11101011; //  926 : 235 - 0xeb
      10'h39F: dout <= 8'b11101011; //  927 : 235 - 0xeb
      10'h3A0: dout <= 8'b11111010; //  928 : 250 - 0xfa -- line 0x1d
      10'h3A1: dout <= 8'b11111010; //  929 : 250 - 0xfa
      10'h3A2: dout <= 8'b11111010; //  930 : 250 - 0xfa
      10'h3A3: dout <= 8'b11111010; //  931 : 250 - 0xfa
      10'h3A4: dout <= 8'b11111010; //  932 : 250 - 0xfa
      10'h3A5: dout <= 8'b11111010; //  933 : 250 - 0xfa
      10'h3A6: dout <= 8'b11111010; //  934 : 250 - 0xfa
      10'h3A7: dout <= 8'b11111010; //  935 : 250 - 0xfa
      10'h3A8: dout <= 8'b11111010; //  936 : 250 - 0xfa
      10'h3A9: dout <= 8'b11111010; //  937 : 250 - 0xfa
      10'h3AA: dout <= 8'b11111010; //  938 : 250 - 0xfa
      10'h3AB: dout <= 8'b11111010; //  939 : 250 - 0xfa
      10'h3AC: dout <= 8'b11111010; //  940 : 250 - 0xfa
      10'h3AD: dout <= 8'b11111010; //  941 : 250 - 0xfa
      10'h3AE: dout <= 8'b11111010; //  942 : 250 - 0xfa
      10'h3AF: dout <= 8'b11101010; //  943 : 234 - 0xea
      10'h3B0: dout <= 8'b11111010; //  944 : 250 - 0xfa
      10'h3B1: dout <= 8'b11111010; //  945 : 250 - 0xfa
      10'h3B2: dout <= 8'b11111010; //  946 : 250 - 0xfa
      10'h3B3: dout <= 8'b11111010; //  947 : 250 - 0xfa
      10'h3B4: dout <= 8'b11111010; //  948 : 250 - 0xfa
      10'h3B5: dout <= 8'b11111010; //  949 : 250 - 0xfa
      10'h3B6: dout <= 8'b11111010; //  950 : 250 - 0xfa
      10'h3B7: dout <= 8'b11111010; //  951 : 250 - 0xfa
      10'h3B8: dout <= 8'b11111010; //  952 : 250 - 0xfa
      10'h3B9: dout <= 8'b11111010; //  953 : 250 - 0xfa
      10'h3BA: dout <= 8'b11111010; //  954 : 250 - 0xfa
      10'h3BB: dout <= 8'b11111010; //  955 : 250 - 0xfa
      10'h3BC: dout <= 8'b11111010; //  956 : 250 - 0xfa
      10'h3BD: dout <= 8'b11111010; //  957 : 250 - 0xfa
      10'h3BE: dout <= 8'b11111010; //  958 : 250 - 0xfa
      10'h3BF: dout <= 8'b11111001; //  959 : 249 - 0xf9
        //-- Attribute Table 0----
      10'h3C0: dout <= 8'b01010101; //  960 :  85 - 0x55
      10'h3C1: dout <= 8'b01010101; //  961 :  85 - 0x55
      10'h3C2: dout <= 8'b01010101; //  962 :  85 - 0x55
      10'h3C3: dout <= 8'b01010101; //  963 :  85 - 0x55
      10'h3C4: dout <= 8'b01010101; //  964 :  85 - 0x55
      10'h3C5: dout <= 8'b01010101; //  965 :  85 - 0x55
      10'h3C6: dout <= 8'b01010101; //  966 :  85 - 0x55
      10'h3C7: dout <= 8'b01010101; //  967 :  85 - 0x55
      10'h3C8: dout <= 8'b01010101; //  968 :  85 - 0x55
      10'h3C9: dout <= 8'b01010101; //  969 :  85 - 0x55
      10'h3CA: dout <= 8'b01010101; //  970 :  85 - 0x55
      10'h3CB: dout <= 8'b01010101; //  971 :  85 - 0x55
      10'h3CC: dout <= 8'b01010101; //  972 :  85 - 0x55
      10'h3CD: dout <= 8'b01010101; //  973 :  85 - 0x55
      10'h3CE: dout <= 8'b01010101; //  974 :  85 - 0x55
      10'h3CF: dout <= 8'b01010101; //  975 :  85 - 0x55
      10'h3D0: dout <= 8'b01010101; //  976 :  85 - 0x55
      10'h3D1: dout <= 8'b01010101; //  977 :  85 - 0x55
      10'h3D2: dout <= 8'b01010101; //  978 :  85 - 0x55
      10'h3D3: dout <= 8'b01010101; //  979 :  85 - 0x55
      10'h3D4: dout <= 8'b01010101; //  980 :  85 - 0x55
      10'h3D5: dout <= 8'b01010101; //  981 :  85 - 0x55
      10'h3D6: dout <= 8'b01010101; //  982 :  85 - 0x55
      10'h3D7: dout <= 8'b01010101; //  983 :  85 - 0x55
      10'h3D8: dout <= 8'b01010101; //  984 :  85 - 0x55
      10'h3D9: dout <= 8'b01010101; //  985 :  85 - 0x55
      10'h3DA: dout <= 8'b01010101; //  986 :  85 - 0x55
      10'h3DB: dout <= 8'b01010101; //  987 :  85 - 0x55
      10'h3DC: dout <= 8'b01010101; //  988 :  85 - 0x55
      10'h3DD: dout <= 8'b01010101; //  989 :  85 - 0x55
      10'h3DE: dout <= 8'b01010101; //  990 :  85 - 0x55
      10'h3DF: dout <= 8'b01010101; //  991 :  85 - 0x55
      10'h3E0: dout <= 8'b01010101; //  992 :  85 - 0x55
      10'h3E1: dout <= 8'b01010101; //  993 :  85 - 0x55
      10'h3E2: dout <= 8'b01010101; //  994 :  85 - 0x55
      10'h3E3: dout <= 8'b01010101; //  995 :  85 - 0x55
      10'h3E4: dout <= 8'b01010101; //  996 :  85 - 0x55
      10'h3E5: dout <= 8'b01010101; //  997 :  85 - 0x55
      10'h3E6: dout <= 8'b01010101; //  998 :  85 - 0x55
      10'h3E7: dout <= 8'b01010101; //  999 :  85 - 0x55
      10'h3E8: dout <= 8'b01010101; // 1000 :  85 - 0x55
      10'h3E9: dout <= 8'b01010101; // 1001 :  85 - 0x55
      10'h3EA: dout <= 8'b01010101; // 1002 :  85 - 0x55
      10'h3EB: dout <= 8'b01010101; // 1003 :  85 - 0x55
      10'h3EC: dout <= 8'b01010101; // 1004 :  85 - 0x55
      10'h3ED: dout <= 8'b01010101; // 1005 :  85 - 0x55
      10'h3EE: dout <= 8'b01010101; // 1006 :  85 - 0x55
      10'h3EF: dout <= 8'b01010101; // 1007 :  85 - 0x55
      10'h3F0: dout <= 8'b00000000; // 1008 :   0 - 0x0
      10'h3F1: dout <= 8'b00000000; // 1009 :   0 - 0x0
      10'h3F2: dout <= 8'b00000000; // 1010 :   0 - 0x0
      10'h3F3: dout <= 8'b00000000; // 1011 :   0 - 0x0
      10'h3F4: dout <= 8'b00000000; // 1012 :   0 - 0x0
      10'h3F5: dout <= 8'b00000000; // 1013 :   0 - 0x0
      10'h3F6: dout <= 8'b00000000; // 1014 :   0 - 0x0
      10'h3F7: dout <= 8'b00000000; // 1015 :   0 - 0x0
      10'h3F8: dout <= 8'b00000101; // 1016 :   5 - 0x5
      10'h3F9: dout <= 8'b00000101; // 1017 :   5 - 0x5
      10'h3FA: dout <= 8'b00000101; // 1018 :   5 - 0x5
      10'h3FB: dout <= 8'b00000101; // 1019 :   5 - 0x5
      10'h3FC: dout <= 8'b00000101; // 1020 :   5 - 0x5
      10'h3FD: dout <= 8'b00000101; // 1021 :   5 - 0x5
      10'h3FE: dout <= 8'b00000101; // 1022 :   5 - 0x5
      10'h3FF: dout <= 8'b00000101; // 1023 :   5 - 0x5
    endcase
  end

endmodule
