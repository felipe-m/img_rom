--- Autcmatically generated VHDL ROM from a NES memory file----
---   NAME TABLE
-- https://wiki.nesdev.com/w/index.php/PPU_nametables
--- Only the first Name Table: 1KiB


---  Original memory dump file name: sprilo_racet2.bin --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory with clock ------

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--    clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (a clock cycle later)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_NTABLE_SPRILO_RACE2 is
  port (
    clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(10-1 downto 0);  --1024 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_NTABLE_SPRILO_RACE2;

architecture BEHAVIORAL of ROM_NTABLE_SPRILO_RACE2 is
  signal addr_int  : natural range 0 to 2**10-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
     ------- Name Table 0---------
    "11111010", --    0 -  0x0  :  250 - 0xfa -- line 0x0
    "11111010", --    1 -  0x1  :  250 - 0xfa
    "11111010", --    2 -  0x2  :  250 - 0xfa
    "11101010", --    3 -  0x3  :  234 - 0xea
    "11111010", --    4 -  0x4  :  250 - 0xfa
    "11111010", --    5 -  0x5  :  250 - 0xfa
    "11111010", --    6 -  0x6  :  250 - 0xfa
    "11111010", --    7 -  0x7  :  250 - 0xfa
    "11111010", --    8 -  0x8  :  250 - 0xfa
    "11111010", --    9 -  0x9  :  250 - 0xfa
    "11111010", --   10 -  0xa  :  250 - 0xfa
    "11111010", --   11 -  0xb  :  250 - 0xfa
    "11111010", --   12 -  0xc  :  250 - 0xfa
    "11111010", --   13 -  0xd  :  250 - 0xfa
    "11101010", --   14 -  0xe  :  234 - 0xea
    "11111010", --   15 -  0xf  :  250 - 0xfa
    "11111010", --   16 - 0x10  :  250 - 0xfa
    "11111010", --   17 - 0x11  :  250 - 0xfa
    "11111010", --   18 - 0x12  :  250 - 0xfa
    "11111010", --   19 - 0x13  :  250 - 0xfa
    "11111010", --   20 - 0x14  :  250 - 0xfa
    "11111010", --   21 - 0x15  :  250 - 0xfa
    "11111010", --   22 - 0x16  :  250 - 0xfa
    "11111010", --   23 - 0x17  :  250 - 0xfa
    "11111010", --   24 - 0x18  :  250 - 0xfa
    "11111010", --   25 - 0x19  :  250 - 0xfa
    "11111010", --   26 - 0x1a  :  250 - 0xfa
    "11111010", --   27 - 0x1b  :  250 - 0xfa
    "11101010", --   28 - 0x1c  :  234 - 0xea
    "11111010", --   29 - 0x1d  :  250 - 0xfa
    "11111010", --   30 - 0x1e  :  250 - 0xfa
    "11111010", --   31 - 0x1f  :  250 - 0xfa
    "11111010", --   32 - 0x20  :  250 - 0xfa -- line 0x1
    "11100111", --   33 - 0x21  :  231 - 0xe7
    "11111011", --   34 - 0x22  :  251 - 0xfb
    "11111011", --   35 - 0x23  :  251 - 0xfb
    "11111011", --   36 - 0x24  :  251 - 0xfb
    "11111011", --   37 - 0x25  :  251 - 0xfb
    "11111011", --   38 - 0x26  :  251 - 0xfb
    "11111011", --   39 - 0x27  :  251 - 0xfb
    "11111011", --   40 - 0x28  :  251 - 0xfb
    "11111011", --   41 - 0x29  :  251 - 0xfb
    "11111011", --   42 - 0x2a  :  251 - 0xfb
    "11111011", --   43 - 0x2b  :  251 - 0xfb
    "11111011", --   44 - 0x2c  :  251 - 0xfb
    "11111011", --   45 - 0x2d  :  251 - 0xfb
    "11111011", --   46 - 0x2e  :  251 - 0xfb
    "11111011", --   47 - 0x2f  :  251 - 0xfb
    "11111011", --   48 - 0x30  :  251 - 0xfb
    "11111011", --   49 - 0x31  :  251 - 0xfb
    "11111011", --   50 - 0x32  :  251 - 0xfb
    "11111011", --   51 - 0x33  :  251 - 0xfb
    "11111011", --   52 - 0x34  :  251 - 0xfb
    "11111011", --   53 - 0x35  :  251 - 0xfb
    "11111011", --   54 - 0x36  :  251 - 0xfb
    "11111011", --   55 - 0x37  :  251 - 0xfb
    "11111011", --   56 - 0x38  :  251 - 0xfb
    "11111011", --   57 - 0x39  :  251 - 0xfb
    "11101000", --   58 - 0x3a  :  232 - 0xe8
    "11111010", --   59 - 0x3b  :  250 - 0xfa
    "11111010", --   60 - 0x3c  :  250 - 0xfa
    "11111001", --   61 - 0x3d  :  249 - 0xf9
    "11111010", --   62 - 0x3e  :  250 - 0xfa
    "11111010", --   63 - 0x3f  :  250 - 0xfa
    "11101010", --   64 - 0x40  :  234 - 0xea -- line 0x2
    "11111100", --   65 - 0x41  :  252 - 0xfc
    "11111111", --   66 - 0x42  :  255 - 0xff
    "11111111", --   67 - 0x43  :  255 - 0xff
    "11111111", --   68 - 0x44  :  255 - 0xff
    "11111111", --   69 - 0x45  :  255 - 0xff
    "11111111", --   70 - 0x46  :  255 - 0xff
    "11111111", --   71 - 0x47  :  255 - 0xff
    "11111111", --   72 - 0x48  :  255 - 0xff
    "11111111", --   73 - 0x49  :  255 - 0xff
    "11111111", --   74 - 0x4a  :  255 - 0xff
    "11111111", --   75 - 0x4b  :  255 - 0xff
    "11111111", --   76 - 0x4c  :  255 - 0xff
    "11111111", --   77 - 0x4d  :  255 - 0xff
    "11111111", --   78 - 0x4e  :  255 - 0xff
    "11111111", --   79 - 0x4f  :  255 - 0xff
    "11101111", --   80 - 0x50  :  239 - 0xef
    "11111111", --   81 - 0x51  :  255 - 0xff
    "11111111", --   82 - 0x52  :  255 - 0xff
    "11111111", --   83 - 0x53  :  255 - 0xff
    "11111111", --   84 - 0x54  :  255 - 0xff
    "11111111", --   85 - 0x55  :  255 - 0xff
    "11111111", --   86 - 0x56  :  255 - 0xff
    "11111111", --   87 - 0x57  :  255 - 0xff
    "11111111", --   88 - 0x58  :  255 - 0xff
    "11111111", --   89 - 0x59  :  255 - 0xff
    "11101100", --   90 - 0x5a  :  236 - 0xec
    "11111010", --   91 - 0x5b  :  250 - 0xfa
    "11111010", --   92 - 0x5c  :  250 - 0xfa
    "11111010", --   93 - 0x5d  :  250 - 0xfa
    "11111010", --   94 - 0x5e  :  250 - 0xfa
    "11111010", --   95 - 0x5f  :  250 - 0xfa
    "11111010", --   96 - 0x60  :  250 - 0xfa -- line 0x3
    "11111100", --   97 - 0x61  :  252 - 0xfc
    "11111111", --   98 - 0x62  :  255 - 0xff
    "11111111", --   99 - 0x63  :  255 - 0xff
    "11111111", --  100 - 0x64  :  255 - 0xff
    "11111111", --  101 - 0x65  :  255 - 0xff
    "11111101", --  102 - 0x66  :  253 - 0xfd
    "11111111", --  103 - 0x67  :  255 - 0xff
    "11111101", --  104 - 0x68  :  253 - 0xfd
    "11111111", --  105 - 0x69  :  255 - 0xff
    "11111101", --  106 - 0x6a  :  253 - 0xfd
    "11111111", --  107 - 0x6b  :  255 - 0xff
    "11111101", --  108 - 0x6c  :  253 - 0xfd
    "11111111", --  109 - 0x6d  :  255 - 0xff
    "11111101", --  110 - 0x6e  :  253 - 0xfd
    "11111111", --  111 - 0x6f  :  255 - 0xff
    "11101111", --  112 - 0x70  :  239 - 0xef
    "11111111", --  113 - 0x71  :  255 - 0xff
    "11111101", --  114 - 0x72  :  253 - 0xfd
    "11111111", --  115 - 0x73  :  255 - 0xff
    "11111101", --  116 - 0x74  :  253 - 0xfd
    "11111111", --  117 - 0x75  :  255 - 0xff
    "11111101", --  118 - 0x76  :  253 - 0xfd
    "11111111", --  119 - 0x77  :  255 - 0xff
    "11111101", --  120 - 0x78  :  253 - 0xfd
    "11111111", --  121 - 0x79  :  255 - 0xff
    "11110101", --  122 - 0x7a  :  245 - 0xf5
    "11111011", --  123 - 0x7b  :  251 - 0xfb
    "11111011", --  124 - 0x7c  :  251 - 0xfb
    "11111011", --  125 - 0x7d  :  251 - 0xfb
    "11101000", --  126 - 0x7e  :  232 - 0xe8
    "11111010", --  127 - 0x7f  :  250 - 0xfa
    "11101001", --  128 - 0x80  :  233 - 0xe9 -- line 0x4
    "11111100", --  129 - 0x81  :  252 - 0xfc
    "11111111", --  130 - 0x82  :  255 - 0xff
    "11111111", --  131 - 0x83  :  255 - 0xff
    "11111111", --  132 - 0x84  :  255 - 0xff
    "11111111", --  133 - 0x85  :  255 - 0xff
    "11111101", --  134 - 0x86  :  253 - 0xfd
    "11111111", --  135 - 0x87  :  255 - 0xff
    "11111101", --  136 - 0x88  :  253 - 0xfd
    "11111111", --  137 - 0x89  :  255 - 0xff
    "11111101", --  138 - 0x8a  :  253 - 0xfd
    "11111111", --  139 - 0x8b  :  255 - 0xff
    "11111101", --  140 - 0x8c  :  253 - 0xfd
    "11111111", --  141 - 0x8d  :  255 - 0xff
    "11111101", --  142 - 0x8e  :  253 - 0xfd
    "11111111", --  143 - 0x8f  :  255 - 0xff
    "11101111", --  144 - 0x90  :  239 - 0xef
    "11111111", --  145 - 0x91  :  255 - 0xff
    "11111101", --  146 - 0x92  :  253 - 0xfd
    "11111111", --  147 - 0x93  :  255 - 0xff
    "11111101", --  148 - 0x94  :  253 - 0xfd
    "11111111", --  149 - 0x95  :  255 - 0xff
    "11111101", --  150 - 0x96  :  253 - 0xfd
    "11111111", --  151 - 0x97  :  255 - 0xff
    "11111101", --  152 - 0x98  :  253 - 0xfd
    "11111111", --  153 - 0x99  :  255 - 0xff
    "11111111", --  154 - 0x9a  :  255 - 0xff
    "11111111", --  155 - 0x9b  :  255 - 0xff
    "11111111", --  156 - 0x9c  :  255 - 0xff
    "11111111", --  157 - 0x9d  :  255 - 0xff
    "11101100", --  158 - 0x9e  :  236 - 0xec
    "11111010", --  159 - 0x9f  :  250 - 0xfa
    "11111010", --  160 - 0xa0  :  250 - 0xfa -- line 0x5
    "11111100", --  161 - 0xa1  :  252 - 0xfc
    "11111111", --  162 - 0xa2  :  255 - 0xff
    "11111110", --  163 - 0xa3  :  254 - 0xfe
    "11111110", --  164 - 0xa4  :  254 - 0xfe
    "11111111", --  165 - 0xa5  :  255 - 0xff
    "11111111", --  166 - 0xa6  :  255 - 0xff
    "11111111", --  167 - 0xa7  :  255 - 0xff
    "11111111", --  168 - 0xa8  :  255 - 0xff
    "11111111", --  169 - 0xa9  :  255 - 0xff
    "11111111", --  170 - 0xaa  :  255 - 0xff
    "11111111", --  171 - 0xab  :  255 - 0xff
    "11111111", --  172 - 0xac  :  255 - 0xff
    "11111111", --  173 - 0xad  :  255 - 0xff
    "11111111", --  174 - 0xae  :  255 - 0xff
    "11111111", --  175 - 0xaf  :  255 - 0xff
    "11101111", --  176 - 0xb0  :  239 - 0xef
    "11111111", --  177 - 0xb1  :  255 - 0xff
    "11111111", --  178 - 0xb2  :  255 - 0xff
    "11111111", --  179 - 0xb3  :  255 - 0xff
    "11111111", --  180 - 0xb4  :  255 - 0xff
    "11111111", --  181 - 0xb5  :  255 - 0xff
    "11111111", --  182 - 0xb6  :  255 - 0xff
    "11111111", --  183 - 0xb7  :  255 - 0xff
    "11111111", --  184 - 0xb8  :  255 - 0xff
    "11111111", --  185 - 0xb9  :  255 - 0xff
    "11111101", --  186 - 0xba  :  253 - 0xfd
    "11111111", --  187 - 0xbb  :  255 - 0xff
    "11111111", --  188 - 0xbc  :  255 - 0xff
    "11111111", --  189 - 0xbd  :  255 - 0xff
    "11101100", --  190 - 0xbe  :  236 - 0xec
    "11111010", --  191 - 0xbf  :  250 - 0xfa
    "11111010", --  192 - 0xc0  :  250 - 0xfa -- line 0x6
    "11111100", --  193 - 0xc1  :  252 - 0xfc
    "11111111", --  194 - 0xc2  :  255 - 0xff
    "11111111", --  195 - 0xc3  :  255 - 0xff
    "11111111", --  196 - 0xc4  :  255 - 0xff
    "11111111", --  197 - 0xc5  :  255 - 0xff
    "11100101", --  198 - 0xc6  :  229 - 0xe5
    "11101011", --  199 - 0xc7  :  235 - 0xeb
    "11101011", --  200 - 0xc8  :  235 - 0xeb
    "11101011", --  201 - 0xc9  :  235 - 0xeb
    "11101011", --  202 - 0xca  :  235 - 0xeb
    "11101011", --  203 - 0xcb  :  235 - 0xeb
    "11101011", --  204 - 0xcc  :  235 - 0xeb
    "11101011", --  205 - 0xcd  :  235 - 0xeb
    "11101011", --  206 - 0xce  :  235 - 0xeb
    "11101011", --  207 - 0xcf  :  235 - 0xeb
    "11101011", --  208 - 0xd0  :  235 - 0xeb
    "11101011", --  209 - 0xd1  :  235 - 0xeb
    "11101011", --  210 - 0xd2  :  235 - 0xeb
    "11101011", --  211 - 0xd3  :  235 - 0xeb
    "11101011", --  212 - 0xd4  :  235 - 0xeb
    "11101011", --  213 - 0xd5  :  235 - 0xeb
    "11101011", --  214 - 0xd6  :  235 - 0xeb
    "11100110", --  215 - 0xd7  :  230 - 0xe6
    "11111111", --  216 - 0xd8  :  255 - 0xff
    "11111111", --  217 - 0xd9  :  255 - 0xff
    "11111101", --  218 - 0xda  :  253 - 0xfd
    "11111111", --  219 - 0xdb  :  255 - 0xff
    "11111111", --  220 - 0xdc  :  255 - 0xff
    "11111111", --  221 - 0xdd  :  255 - 0xff
    "11101100", --  222 - 0xde  :  236 - 0xec
    "11111010", --  223 - 0xdf  :  250 - 0xfa
    "11111010", --  224 - 0xe0  :  250 - 0xfa -- line 0x7
    "11111100", --  225 - 0xe1  :  252 - 0xfc
    "11111111", --  226 - 0xe2  :  255 - 0xff
    "11111110", --  227 - 0xe3  :  254 - 0xfe
    "11111110", --  228 - 0xe4  :  254 - 0xfe
    "11111111", --  229 - 0xe5  :  255 - 0xff
    "11101100", --  230 - 0xe6  :  236 - 0xec
    "11100111", --  231 - 0xe7  :  231 - 0xe7
    "11111011", --  232 - 0xe8  :  251 - 0xfb
    "11111011", --  233 - 0xe9  :  251 - 0xfb
    "11111011", --  234 - 0xea  :  251 - 0xfb
    "11111011", --  235 - 0xeb  :  251 - 0xfb
    "11111011", --  236 - 0xec  :  251 - 0xfb
    "11111011", --  237 - 0xed  :  251 - 0xfb
    "11111011", --  238 - 0xee  :  251 - 0xfb
    "11111011", --  239 - 0xef  :  251 - 0xfb
    "11111011", --  240 - 0xf0  :  251 - 0xfb
    "11111011", --  241 - 0xf1  :  251 - 0xfb
    "11111011", --  242 - 0xf2  :  251 - 0xfb
    "11111011", --  243 - 0xf3  :  251 - 0xfb
    "11111011", --  244 - 0xf4  :  251 - 0xfb
    "11111011", --  245 - 0xf5  :  251 - 0xfb
    "11101000", --  246 - 0xf6  :  232 - 0xe8
    "11111100", --  247 - 0xf7  :  252 - 0xfc
    "11111111", --  248 - 0xf8  :  255 - 0xff
    "11111111", --  249 - 0xf9  :  255 - 0xff
    "11111111", --  250 - 0xfa  :  255 - 0xff
    "11111111", --  251 - 0xfb  :  255 - 0xff
    "11111111", --  252 - 0xfc  :  255 - 0xff
    "11111111", --  253 - 0xfd  :  255 - 0xff
    "11101100", --  254 - 0xfe  :  236 - 0xec
    "11111010", --  255 - 0xff  :  250 - 0xfa
    "11111010", --  256 - 0x100  :  250 - 0xfa -- line 0x8
    "11111100", --  257 - 0x101  :  252 - 0xfc
    "11111111", --  258 - 0x102  :  255 - 0xff
    "11111111", --  259 - 0x103  :  255 - 0xff
    "11111111", --  260 - 0x104  :  255 - 0xff
    "11111111", --  261 - 0x105  :  255 - 0xff
    "11101100", --  262 - 0x106  :  236 - 0xec
    "11111100", --  263 - 0x107  :  252 - 0xfc
    "11111111", --  264 - 0x108  :  255 - 0xff
    "11111111", --  265 - 0x109  :  255 - 0xff
    "11111111", --  266 - 0x10a  :  255 - 0xff
    "11111111", --  267 - 0x10b  :  255 - 0xff
    "11111111", --  268 - 0x10c  :  255 - 0xff
    "11111111", --  269 - 0x10d  :  255 - 0xff
    "11111111", --  270 - 0x10e  :  255 - 0xff
    "11111111", --  271 - 0x10f  :  255 - 0xff
    "11111111", --  272 - 0x110  :  255 - 0xff
    "11111111", --  273 - 0x111  :  255 - 0xff
    "11111111", --  274 - 0x112  :  255 - 0xff
    "11111111", --  275 - 0x113  :  255 - 0xff
    "11111111", --  276 - 0x114  :  255 - 0xff
    "11111111", --  277 - 0x115  :  255 - 0xff
    "11101100", --  278 - 0x116  :  236 - 0xec
    "11110111", --  279 - 0x117  :  247 - 0xf7
    "11101011", --  280 - 0x118  :  235 - 0xeb
    "11100110", --  281 - 0x119  :  230 - 0xe6
    "11111111", --  282 - 0x11a  :  255 - 0xff
    "11111110", --  283 - 0x11b  :  254 - 0xfe
    "11111110", --  284 - 0x11c  :  254 - 0xfe
    "11111111", --  285 - 0x11d  :  255 - 0xff
    "11101100", --  286 - 0x11e  :  236 - 0xec
    "11111010", --  287 - 0x11f  :  250 - 0xfa
    "11111010", --  288 - 0x120  :  250 - 0xfa -- line 0x9
    "11111100", --  289 - 0x121  :  252 - 0xfc
    "11111111", --  290 - 0x122  :  255 - 0xff
    "11111110", --  291 - 0x123  :  254 - 0xfe
    "11111110", --  292 - 0x124  :  254 - 0xfe
    "11111111", --  293 - 0x125  :  255 - 0xff
    "11101100", --  294 - 0x126  :  236 - 0xec
    "11111100", --  295 - 0x127  :  252 - 0xfc
    "11111111", --  296 - 0x128  :  255 - 0xff
    "11111111", --  297 - 0x129  :  255 - 0xff
    "11111111", --  298 - 0x12a  :  255 - 0xff
    "11111111", --  299 - 0x12b  :  255 - 0xff
    "11111101", --  300 - 0x12c  :  253 - 0xfd
    "11111111", --  301 - 0x12d  :  255 - 0xff
    "11111101", --  302 - 0x12e  :  253 - 0xfd
    "11111111", --  303 - 0x12f  :  255 - 0xff
    "11111101", --  304 - 0x130  :  253 - 0xfd
    "11111111", --  305 - 0x131  :  255 - 0xff
    "11111101", --  306 - 0x132  :  253 - 0xfd
    "11111111", --  307 - 0x133  :  255 - 0xff
    "11111111", --  308 - 0x134  :  255 - 0xff
    "11111111", --  309 - 0x135  :  255 - 0xff
    "11101100", --  310 - 0x136  :  236 - 0xec
    "11111010", --  311 - 0x137  :  250 - 0xfa
    "11111010", --  312 - 0x138  :  250 - 0xfa
    "11111100", --  313 - 0x139  :  252 - 0xfc
    "11111111", --  314 - 0x13a  :  255 - 0xff
    "11111111", --  315 - 0x13b  :  255 - 0xff
    "11111111", --  316 - 0x13c  :  255 - 0xff
    "11111111", --  317 - 0x13d  :  255 - 0xff
    "11101100", --  318 - 0x13e  :  236 - 0xec
    "11111010", --  319 - 0x13f  :  250 - 0xfa
    "11111010", --  320 - 0x140  :  250 - 0xfa -- line 0xa
    "11111100", --  321 - 0x141  :  252 - 0xfc
    "11111111", --  322 - 0x142  :  255 - 0xff
    "11111111", --  323 - 0x143  :  255 - 0xff
    "11111111", --  324 - 0x144  :  255 - 0xff
    "11111111", --  325 - 0x145  :  255 - 0xff
    "11101100", --  326 - 0x146  :  236 - 0xec
    "11111100", --  327 - 0x147  :  252 - 0xfc
    "11111111", --  328 - 0x148  :  255 - 0xff
    "11111111", --  329 - 0x149  :  255 - 0xff
    "11111111", --  330 - 0x14a  :  255 - 0xff
    "11111111", --  331 - 0x14b  :  255 - 0xff
    "11111101", --  332 - 0x14c  :  253 - 0xfd
    "11111111", --  333 - 0x14d  :  255 - 0xff
    "11111101", --  334 - 0x14e  :  253 - 0xfd
    "11111111", --  335 - 0x14f  :  255 - 0xff
    "11111101", --  336 - 0x150  :  253 - 0xfd
    "11111111", --  337 - 0x151  :  255 - 0xff
    "11111101", --  338 - 0x152  :  253 - 0xfd
    "11111111", --  339 - 0x153  :  255 - 0xff
    "11111111", --  340 - 0x154  :  255 - 0xff
    "11111111", --  341 - 0x155  :  255 - 0xff
    "11101100", --  342 - 0x156  :  236 - 0xec
    "11111010", --  343 - 0x157  :  250 - 0xfa
    "11111010", --  344 - 0x158  :  250 - 0xfa
    "11111100", --  345 - 0x159  :  252 - 0xfc
    "11111111", --  346 - 0x15a  :  255 - 0xff
    "11111110", --  347 - 0x15b  :  254 - 0xfe
    "11111110", --  348 - 0x15c  :  254 - 0xfe
    "11111111", --  349 - 0x15d  :  255 - 0xff
    "11101100", --  350 - 0x15e  :  236 - 0xec
    "11111010", --  351 - 0x15f  :  250 - 0xfa
    "11111010", --  352 - 0x160  :  250 - 0xfa -- line 0xb
    "11111100", --  353 - 0x161  :  252 - 0xfc
    "11111111", --  354 - 0x162  :  255 - 0xff
    "11111110", --  355 - 0x163  :  254 - 0xfe
    "11111110", --  356 - 0x164  :  254 - 0xfe
    "11111111", --  357 - 0x165  :  255 - 0xff
    "11101100", --  358 - 0x166  :  236 - 0xec
    "11111100", --  359 - 0x167  :  252 - 0xfc
    "11111111", --  360 - 0x168  :  255 - 0xff
    "11111111", --  361 - 0x169  :  255 - 0xff
    "11111111", --  362 - 0x16a  :  255 - 0xff
    "11111111", --  363 - 0x16b  :  255 - 0xff
    "11111111", --  364 - 0x16c  :  255 - 0xff
    "11111111", --  365 - 0x16d  :  255 - 0xff
    "11111111", --  366 - 0x16e  :  255 - 0xff
    "11111111", --  367 - 0x16f  :  255 - 0xff
    "11111111", --  368 - 0x170  :  255 - 0xff
    "11111111", --  369 - 0x171  :  255 - 0xff
    "11111111", --  370 - 0x172  :  255 - 0xff
    "11111111", --  371 - 0x173  :  255 - 0xff
    "11111111", --  372 - 0x174  :  255 - 0xff
    "11111111", --  373 - 0x175  :  255 - 0xff
    "11101100", --  374 - 0x176  :  236 - 0xec
    "11111010", --  375 - 0x177  :  250 - 0xfa
    "11101010", --  376 - 0x178  :  234 - 0xea
    "11111100", --  377 - 0x179  :  252 - 0xfc
    "11111111", --  378 - 0x17a  :  255 - 0xff
    "11111111", --  379 - 0x17b  :  255 - 0xff
    "11111111", --  380 - 0x17c  :  255 - 0xff
    "11111111", --  381 - 0x17d  :  255 - 0xff
    "11101100", --  382 - 0x17e  :  236 - 0xec
    "11111010", --  383 - 0x17f  :  250 - 0xfa
    "11101001", --  384 - 0x180  :  233 - 0xe9 -- line 0xc
    "11111100", --  385 - 0x181  :  252 - 0xfc
    "11111111", --  386 - 0x182  :  255 - 0xff
    "11111111", --  387 - 0x183  :  255 - 0xff
    "11111111", --  388 - 0x184  :  255 - 0xff
    "11111111", --  389 - 0x185  :  255 - 0xff
    "11101100", --  390 - 0x186  :  236 - 0xec
    "11111100", --  391 - 0x187  :  252 - 0xfc
    "11111111", --  392 - 0x188  :  255 - 0xff
    "11111110", --  393 - 0x189  :  254 - 0xfe
    "11111110", --  394 - 0x18a  :  254 - 0xfe
    "11111111", --  395 - 0x18b  :  255 - 0xff
    "11100101", --  396 - 0x18c  :  229 - 0xe5
    "11101011", --  397 - 0x18d  :  235 - 0xeb
    "11101011", --  398 - 0x18e  :  235 - 0xeb
    "11101011", --  399 - 0x18f  :  235 - 0xeb
    "11101011", --  400 - 0x190  :  235 - 0xeb
    "11100110", --  401 - 0x191  :  230 - 0xe6
    "11111111", --  402 - 0x192  :  255 - 0xff
    "11111110", --  403 - 0x193  :  254 - 0xfe
    "11111110", --  404 - 0x194  :  254 - 0xfe
    "11111111", --  405 - 0x195  :  255 - 0xff
    "11101100", --  406 - 0x196  :  236 - 0xec
    "11101010", --  407 - 0x197  :  234 - 0xea
    "11111010", --  408 - 0x198  :  250 - 0xfa
    "11111100", --  409 - 0x199  :  252 - 0xfc
    "11111111", --  410 - 0x19a  :  255 - 0xff
    "11111110", --  411 - 0x19b  :  254 - 0xfe
    "11111110", --  412 - 0x19c  :  254 - 0xfe
    "11111111", --  413 - 0x19d  :  255 - 0xff
    "11101100", --  414 - 0x19e  :  236 - 0xec
    "11111010", --  415 - 0x19f  :  250 - 0xfa
    "11111010", --  416 - 0x1a0  :  250 - 0xfa -- line 0xd
    "11111100", --  417 - 0x1a1  :  252 - 0xfc
    "11111111", --  418 - 0x1a2  :  255 - 0xff
    "11111110", --  419 - 0x1a3  :  254 - 0xfe
    "11111110", --  420 - 0x1a4  :  254 - 0xfe
    "11111111", --  421 - 0x1a5  :  255 - 0xff
    "11101100", --  422 - 0x1a6  :  236 - 0xec
    "11111100", --  423 - 0x1a7  :  252 - 0xfc
    "11111111", --  424 - 0x1a8  :  255 - 0xff
    "11111111", --  425 - 0x1a9  :  255 - 0xff
    "11111111", --  426 - 0x1aa  :  255 - 0xff
    "11111111", --  427 - 0x1ab  :  255 - 0xff
    "11101100", --  428 - 0x1ac  :  236 - 0xec
    "11100111", --  429 - 0x1ad  :  231 - 0xe7
    "11111011", --  430 - 0x1ae  :  251 - 0xfb
    "11111011", --  431 - 0x1af  :  251 - 0xfb
    "11111011", --  432 - 0x1b0  :  251 - 0xfb
    "11110110", --  433 - 0x1b1  :  246 - 0xf6
    "11111111", --  434 - 0x1b2  :  255 - 0xff
    "11111111", --  435 - 0x1b3  :  255 - 0xff
    "11111111", --  436 - 0x1b4  :  255 - 0xff
    "11111111", --  437 - 0x1b5  :  255 - 0xff
    "11101100", --  438 - 0x1b6  :  236 - 0xec
    "11111010", --  439 - 0x1b7  :  250 - 0xfa
    "11111010", --  440 - 0x1b8  :  250 - 0xfa
    "11111100", --  441 - 0x1b9  :  252 - 0xfc
    "11111111", --  442 - 0x1ba  :  255 - 0xff
    "11111111", --  443 - 0x1bb  :  255 - 0xff
    "11111111", --  444 - 0x1bc  :  255 - 0xff
    "11111111", --  445 - 0x1bd  :  255 - 0xff
    "11101100", --  446 - 0x1be  :  236 - 0xec
    "11101001", --  447 - 0x1bf  :  233 - 0xe9
    "11111010", --  448 - 0x1c0  :  250 - 0xfa -- line 0xe
    "11111100", --  449 - 0x1c1  :  252 - 0xfc
    "11111111", --  450 - 0x1c2  :  255 - 0xff
    "11111111", --  451 - 0x1c3  :  255 - 0xff
    "11111111", --  452 - 0x1c4  :  255 - 0xff
    "11111111", --  453 - 0x1c5  :  255 - 0xff
    "11101100", --  454 - 0x1c6  :  236 - 0xec
    "11111100", --  455 - 0x1c7  :  252 - 0xfc
    "11111111", --  456 - 0x1c8  :  255 - 0xff
    "11111110", --  457 - 0x1c9  :  254 - 0xfe
    "11111110", --  458 - 0x1ca  :  254 - 0xfe
    "11111111", --  459 - 0x1cb  :  255 - 0xff
    "11101100", --  460 - 0x1cc  :  236 - 0xec
    "11111100", --  461 - 0x1cd  :  252 - 0xfc
    "11111111", --  462 - 0x1ce  :  255 - 0xff
    "11111111", --  463 - 0x1cf  :  255 - 0xff
    "11111111", --  464 - 0x1d0  :  255 - 0xff
    "11111111", --  465 - 0x1d1  :  255 - 0xff
    "11111111", --  466 - 0x1d2  :  255 - 0xff
    "11111110", --  467 - 0x1d3  :  254 - 0xfe
    "11111110", --  468 - 0x1d4  :  254 - 0xfe
    "11111111", --  469 - 0x1d5  :  255 - 0xff
    "11101100", --  470 - 0x1d6  :  236 - 0xec
    "11111010", --  471 - 0x1d7  :  250 - 0xfa
    "11111010", --  472 - 0x1d8  :  250 - 0xfa
    "11111100", --  473 - 0x1d9  :  252 - 0xfc
    "11111111", --  474 - 0x1da  :  255 - 0xff
    "11111110", --  475 - 0x1db  :  254 - 0xfe
    "11111110", --  476 - 0x1dc  :  254 - 0xfe
    "11111111", --  477 - 0x1dd  :  255 - 0xff
    "11101100", --  478 - 0x1de  :  236 - 0xec
    "11111010", --  479 - 0x1df  :  250 - 0xfa
    "11101010", --  480 - 0x1e0  :  234 - 0xea -- line 0xf
    "11111100", --  481 - 0x1e1  :  252 - 0xfc
    "11111111", --  482 - 0x1e2  :  255 - 0xff
    "11111110", --  483 - 0x1e3  :  254 - 0xfe
    "11111110", --  484 - 0x1e4  :  254 - 0xfe
    "11111111", --  485 - 0x1e5  :  255 - 0xff
    "11101100", --  486 - 0x1e6  :  236 - 0xec
    "11111100", --  487 - 0x1e7  :  252 - 0xfc
    "11111111", --  488 - 0x1e8  :  255 - 0xff
    "11111111", --  489 - 0x1e9  :  255 - 0xff
    "11111111", --  490 - 0x1ea  :  255 - 0xff
    "11111111", --  491 - 0x1eb  :  255 - 0xff
    "11101100", --  492 - 0x1ec  :  236 - 0xec
    "11111100", --  493 - 0x1ed  :  252 - 0xfc
    "11111111", --  494 - 0x1ee  :  255 - 0xff
    "11111111", --  495 - 0x1ef  :  255 - 0xff
    "11111111", --  496 - 0x1f0  :  255 - 0xff
    "11111101", --  497 - 0x1f1  :  253 - 0xfd
    "11111111", --  498 - 0x1f2  :  255 - 0xff
    "11111111", --  499 - 0x1f3  :  255 - 0xff
    "11111111", --  500 - 0x1f4  :  255 - 0xff
    "11111111", --  501 - 0x1f5  :  255 - 0xff
    "11101100", --  502 - 0x1f6  :  236 - 0xec
    "11100111", --  503 - 0x1f7  :  231 - 0xe7
    "11111011", --  504 - 0x1f8  :  251 - 0xfb
    "11110110", --  505 - 0x1f9  :  246 - 0xf6
    "11111111", --  506 - 0x1fa  :  255 - 0xff
    "11111111", --  507 - 0x1fb  :  255 - 0xff
    "11111111", --  508 - 0x1fc  :  255 - 0xff
    "11111111", --  509 - 0x1fd  :  255 - 0xff
    "11101100", --  510 - 0x1fe  :  236 - 0xec
    "11111010", --  511 - 0x1ff  :  250 - 0xfa
    "11111010", --  512 - 0x200  :  250 - 0xfa -- line 0x10
    "11111100", --  513 - 0x201  :  252 - 0xfc
    "11111111", --  514 - 0x202  :  255 - 0xff
    "11111111", --  515 - 0x203  :  255 - 0xff
    "11111111", --  516 - 0x204  :  255 - 0xff
    "11111111", --  517 - 0x205  :  255 - 0xff
    "11101100", --  518 - 0x206  :  236 - 0xec
    "11111100", --  519 - 0x207  :  252 - 0xfc
    "11111111", --  520 - 0x208  :  255 - 0xff
    "11111110", --  521 - 0x209  :  254 - 0xfe
    "11111110", --  522 - 0x20a  :  254 - 0xfe
    "11111111", --  523 - 0x20b  :  255 - 0xff
    "11101100", --  524 - 0x20c  :  236 - 0xec
    "11111100", --  525 - 0x20d  :  252 - 0xfc
    "11111111", --  526 - 0x20e  :  255 - 0xff
    "11111111", --  527 - 0x20f  :  255 - 0xff
    "11111111", --  528 - 0x210  :  255 - 0xff
    "11111101", --  529 - 0x211  :  253 - 0xfd
    "11111111", --  530 - 0x212  :  255 - 0xff
    "11111111", --  531 - 0x213  :  255 - 0xff
    "11111111", --  532 - 0x214  :  255 - 0xff
    "11111111", --  533 - 0x215  :  255 - 0xff
    "11101100", --  534 - 0x216  :  236 - 0xec
    "11111100", --  535 - 0x217  :  252 - 0xfc
    "11111111", --  536 - 0x218  :  255 - 0xff
    "11111111", --  537 - 0x219  :  255 - 0xff
    "11111111", --  538 - 0x21a  :  255 - 0xff
    "11111111", --  539 - 0x21b  :  255 - 0xff
    "11111111", --  540 - 0x21c  :  255 - 0xff
    "11111111", --  541 - 0x21d  :  255 - 0xff
    "11101100", --  542 - 0x21e  :  236 - 0xec
    "11101010", --  543 - 0x21f  :  234 - 0xea
    "11111010", --  544 - 0x220  :  250 - 0xfa -- line 0x11
    "11111100", --  545 - 0x221  :  252 - 0xfc
    "11111111", --  546 - 0x222  :  255 - 0xff
    "11111110", --  547 - 0x223  :  254 - 0xfe
    "11111110", --  548 - 0x224  :  254 - 0xfe
    "11111111", --  549 - 0x225  :  255 - 0xff
    "11110101", --  550 - 0x226  :  245 - 0xf5
    "11110110", --  551 - 0x227  :  246 - 0xf6
    "11111111", --  552 - 0x228  :  255 - 0xff
    "11111111", --  553 - 0x229  :  255 - 0xff
    "11111111", --  554 - 0x22a  :  255 - 0xff
    "11111111", --  555 - 0x22b  :  255 - 0xff
    "11101100", --  556 - 0x22c  :  236 - 0xec
    "11111100", --  557 - 0x22d  :  252 - 0xfc
    "11111111", --  558 - 0x22e  :  255 - 0xff
    "11111111", --  559 - 0x22f  :  255 - 0xff
    "11111111", --  560 - 0x230  :  255 - 0xff
    "11111111", --  561 - 0x231  :  255 - 0xff
    "11111111", --  562 - 0x232  :  255 - 0xff
    "11111111", --  563 - 0x233  :  255 - 0xff
    "11111111", --  564 - 0x234  :  255 - 0xff
    "11111111", --  565 - 0x235  :  255 - 0xff
    "11101100", --  566 - 0x236  :  236 - 0xec
    "11111100", --  567 - 0x237  :  252 - 0xfc
    "11111111", --  568 - 0x238  :  255 - 0xff
    "11111111", --  569 - 0x239  :  255 - 0xff
    "11111101", --  570 - 0x23a  :  253 - 0xfd
    "11111111", --  571 - 0x23b  :  255 - 0xff
    "11111111", --  572 - 0x23c  :  255 - 0xff
    "11111111", --  573 - 0x23d  :  255 - 0xff
    "11101100", --  574 - 0x23e  :  236 - 0xec
    "11111010", --  575 - 0x23f  :  250 - 0xfa
    "11111010", --  576 - 0x240  :  250 - 0xfa -- line 0x12
    "11111100", --  577 - 0x241  :  252 - 0xfc
    "11111111", --  578 - 0x242  :  255 - 0xff
    "11111111", --  579 - 0x243  :  255 - 0xff
    "11111111", --  580 - 0x244  :  255 - 0xff
    "11111111", --  581 - 0x245  :  255 - 0xff
    "11111111", --  582 - 0x246  :  255 - 0xff
    "11111111", --  583 - 0x247  :  255 - 0xff
    "11111111", --  584 - 0x248  :  255 - 0xff
    "11111110", --  585 - 0x249  :  254 - 0xfe
    "11111110", --  586 - 0x24a  :  254 - 0xfe
    "11111111", --  587 - 0x24b  :  255 - 0xff
    "11101100", --  588 - 0x24c  :  236 - 0xec
    "11111100", --  589 - 0x24d  :  252 - 0xfc
    "11111111", --  590 - 0x24e  :  255 - 0xff
    "11111111", --  591 - 0x24f  :  255 - 0xff
    "11111111", --  592 - 0x250  :  255 - 0xff
    "11111111", --  593 - 0x251  :  255 - 0xff
    "11100101", --  594 - 0x252  :  229 - 0xe5
    "11101011", --  595 - 0x253  :  235 - 0xeb
    "11101011", --  596 - 0x254  :  235 - 0xeb
    "11101011", --  597 - 0x255  :  235 - 0xeb
    "11111000", --  598 - 0x256  :  248 - 0xf8
    "11111100", --  599 - 0x257  :  252 - 0xfc
    "11111111", --  600 - 0x258  :  255 - 0xff
    "11111111", --  601 - 0x259  :  255 - 0xff
    "11111101", --  602 - 0x25a  :  253 - 0xfd
    "11111111", --  603 - 0x25b  :  255 - 0xff
    "11100101", --  604 - 0x25c  :  229 - 0xe5
    "11101011", --  605 - 0x25d  :  235 - 0xeb
    "11111000", --  606 - 0x25e  :  248 - 0xf8
    "11111010", --  607 - 0x25f  :  250 - 0xfa
    "11111001", --  608 - 0x260  :  249 - 0xf9 -- line 0x13
    "11111100", --  609 - 0x261  :  252 - 0xfc
    "11111111", --  610 - 0x262  :  255 - 0xff
    "11111111", --  611 - 0x263  :  255 - 0xff
    "11111111", --  612 - 0x264  :  255 - 0xff
    "11111101", --  613 - 0x265  :  253 - 0xfd
    "11111111", --  614 - 0x266  :  255 - 0xff
    "11111101", --  615 - 0x267  :  253 - 0xfd
    "11111111", --  616 - 0x268  :  255 - 0xff
    "11111111", --  617 - 0x269  :  255 - 0xff
    "11111111", --  618 - 0x26a  :  255 - 0xff
    "11111111", --  619 - 0x26b  :  255 - 0xff
    "11101100", --  620 - 0x26c  :  236 - 0xec
    "11111100", --  621 - 0x26d  :  252 - 0xfc
    "11111111", --  622 - 0x26e  :  255 - 0xff
    "11111110", --  623 - 0x26f  :  254 - 0xfe
    "11111110", --  624 - 0x270  :  254 - 0xfe
    "11111111", --  625 - 0x271  :  255 - 0xff
    "11101100", --  626 - 0x272  :  236 - 0xec
    "11111001", --  627 - 0x273  :  249 - 0xf9
    "11111010", --  628 - 0x274  :  250 - 0xfa
    "11100111", --  629 - 0x275  :  231 - 0xe7
    "11111011", --  630 - 0x276  :  251 - 0xfb
    "11110110", --  631 - 0x277  :  246 - 0xf6
    "11111111", --  632 - 0x278  :  255 - 0xff
    "11111111", --  633 - 0x279  :  255 - 0xff
    "11111111", --  634 - 0x27a  :  255 - 0xff
    "11111111", --  635 - 0x27b  :  255 - 0xff
    "11101100", --  636 - 0x27c  :  236 - 0xec
    "11111001", --  637 - 0x27d  :  249 - 0xf9
    "11111010", --  638 - 0x27e  :  250 - 0xfa
    "11111010", --  639 - 0x27f  :  250 - 0xfa
    "11111010", --  640 - 0x280  :  250 - 0xfa -- line 0x14
    "11111100", --  641 - 0x281  :  252 - 0xfc
    "11111111", --  642 - 0x282  :  255 - 0xff
    "11111111", --  643 - 0x283  :  255 - 0xff
    "11111111", --  644 - 0x284  :  255 - 0xff
    "11111101", --  645 - 0x285  :  253 - 0xfd
    "11111111", --  646 - 0x286  :  255 - 0xff
    "11111101", --  647 - 0x287  :  253 - 0xfd
    "11111111", --  648 - 0x288  :  255 - 0xff
    "11111111", --  649 - 0x289  :  255 - 0xff
    "11111111", --  650 - 0x28a  :  255 - 0xff
    "11111111", --  651 - 0x28b  :  255 - 0xff
    "11101100", --  652 - 0x28c  :  236 - 0xec
    "11111100", --  653 - 0x28d  :  252 - 0xfc
    "11111111", --  654 - 0x28e  :  255 - 0xff
    "11111111", --  655 - 0x28f  :  255 - 0xff
    "11111111", --  656 - 0x290  :  255 - 0xff
    "11111111", --  657 - 0x291  :  255 - 0xff
    "11101100", --  658 - 0x292  :  236 - 0xec
    "11111010", --  659 - 0x293  :  250 - 0xfa
    "11111010", --  660 - 0x294  :  250 - 0xfa
    "11111100", --  661 - 0x295  :  252 - 0xfc
    "11111111", --  662 - 0x296  :  255 - 0xff
    "11111111", --  663 - 0x297  :  255 - 0xff
    "11111111", --  664 - 0x298  :  255 - 0xff
    "11111111", --  665 - 0x299  :  255 - 0xff
    "11111111", --  666 - 0x29a  :  255 - 0xff
    "11111111", --  667 - 0x29b  :  255 - 0xff
    "11101100", --  668 - 0x29c  :  236 - 0xec
    "11111010", --  669 - 0x29d  :  250 - 0xfa
    "11111010", --  670 - 0x29e  :  250 - 0xfa
    "11101010", --  671 - 0x29f  :  234 - 0xea
    "11111010", --  672 - 0x2a0  :  250 - 0xfa -- line 0x15
    "11111100", --  673 - 0x2a1  :  252 - 0xfc
    "11111111", --  674 - 0x2a2  :  255 - 0xff
    "11111111", --  675 - 0x2a3  :  255 - 0xff
    "11111111", --  676 - 0x2a4  :  255 - 0xff
    "11111111", --  677 - 0x2a5  :  255 - 0xff
    "11111111", --  678 - 0x2a6  :  255 - 0xff
    "11111111", --  679 - 0x2a7  :  255 - 0xff
    "11111111", --  680 - 0x2a8  :  255 - 0xff
    "11111111", --  681 - 0x2a9  :  255 - 0xff
    "11111111", --  682 - 0x2aa  :  255 - 0xff
    "11111111", --  683 - 0x2ab  :  255 - 0xff
    "11101100", --  684 - 0x2ac  :  236 - 0xec
    "11111100", --  685 - 0x2ad  :  252 - 0xfc
    "11111111", --  686 - 0x2ae  :  255 - 0xff
    "11111110", --  687 - 0x2af  :  254 - 0xfe
    "11111110", --  688 - 0x2b0  :  254 - 0xfe
    "11111111", --  689 - 0x2b1  :  255 - 0xff
    "11101100", --  690 - 0x2b2  :  236 - 0xec
    "11111010", --  691 - 0x2b3  :  250 - 0xfa
    "11111001", --  692 - 0x2b4  :  249 - 0xf9
    "11111100", --  693 - 0x2b5  :  252 - 0xfc
    "11111111", --  694 - 0x2b6  :  255 - 0xff
    "11111111", --  695 - 0x2b7  :  255 - 0xff
    "11111111", --  696 - 0x2b8  :  255 - 0xff
    "11111101", --  697 - 0x2b9  :  253 - 0xfd
    "11111111", --  698 - 0x2ba  :  255 - 0xff
    "11111111", --  699 - 0x2bb  :  255 - 0xff
    "11101100", --  700 - 0x2bc  :  236 - 0xec
    "11111010", --  701 - 0x2bd  :  250 - 0xfa
    "11111010", --  702 - 0x2be  :  250 - 0xfa
    "11111010", --  703 - 0x2bf  :  250 - 0xfa
    "11111010", --  704 - 0x2c0  :  250 - 0xfa -- line 0x16
    "11110111", --  705 - 0x2c1  :  247 - 0xf7
    "11101011", --  706 - 0x2c2  :  235 - 0xeb
    "11101011", --  707 - 0x2c3  :  235 - 0xeb
    "11101011", --  708 - 0x2c4  :  235 - 0xeb
    "11101011", --  709 - 0x2c5  :  235 - 0xeb
    "11101011", --  710 - 0x2c6  :  235 - 0xeb
    "11101011", --  711 - 0x2c7  :  235 - 0xeb
    "11101011", --  712 - 0x2c8  :  235 - 0xeb
    "11101011", --  713 - 0x2c9  :  235 - 0xeb
    "11101011", --  714 - 0x2ca  :  235 - 0xeb
    "11101011", --  715 - 0x2cb  :  235 - 0xeb
    "11111000", --  716 - 0x2cc  :  248 - 0xf8
    "11111100", --  717 - 0x2cd  :  252 - 0xfc
    "11111111", --  718 - 0x2ce  :  255 - 0xff
    "11111111", --  719 - 0x2cf  :  255 - 0xff
    "11111111", --  720 - 0x2d0  :  255 - 0xff
    "11111111", --  721 - 0x2d1  :  255 - 0xff
    "11101100", --  722 - 0x2d2  :  236 - 0xec
    "11111010", --  723 - 0x2d3  :  250 - 0xfa
    "11111010", --  724 - 0x2d4  :  250 - 0xfa
    "11111100", --  725 - 0x2d5  :  252 - 0xfc
    "11111111", --  726 - 0x2d6  :  255 - 0xff
    "11111111", --  727 - 0x2d7  :  255 - 0xff
    "11111111", --  728 - 0x2d8  :  255 - 0xff
    "11111101", --  729 - 0x2d9  :  253 - 0xfd
    "11111111", --  730 - 0x2da  :  255 - 0xff
    "11111111", --  731 - 0x2db  :  255 - 0xff
    "11101100", --  732 - 0x2dc  :  236 - 0xec
    "11111010", --  733 - 0x2dd  :  250 - 0xfa
    "11111010", --  734 - 0x2de  :  250 - 0xfa
    "11111010", --  735 - 0x2df  :  250 - 0xfa
    "11111010", --  736 - 0x2e0  :  250 - 0xfa -- line 0x17
    "11111010", --  737 - 0x2e1  :  250 - 0xfa
    "11111010", --  738 - 0x2e2  :  250 - 0xfa
    "11111010", --  739 - 0x2e3  :  250 - 0xfa
    "11111010", --  740 - 0x2e4  :  250 - 0xfa
    "11111010", --  741 - 0x2e5  :  250 - 0xfa
    "11111010", --  742 - 0x2e6  :  250 - 0xfa
    "11111010", --  743 - 0x2e7  :  250 - 0xfa
    "11111010", --  744 - 0x2e8  :  250 - 0xfa
    "11111010", --  745 - 0x2e9  :  250 - 0xfa
    "11111001", --  746 - 0x2ea  :  249 - 0xf9
    "11111010", --  747 - 0x2eb  :  250 - 0xfa
    "11111010", --  748 - 0x2ec  :  250 - 0xfa
    "11111100", --  749 - 0x2ed  :  252 - 0xfc
    "11111111", --  750 - 0x2ee  :  255 - 0xff
    "11111110", --  751 - 0x2ef  :  254 - 0xfe
    "11111110", --  752 - 0x2f0  :  254 - 0xfe
    "11111111", --  753 - 0x2f1  :  255 - 0xff
    "11110101", --  754 - 0x2f2  :  245 - 0xf5
    "11111011", --  755 - 0x2f3  :  251 - 0xfb
    "11111011", --  756 - 0x2f4  :  251 - 0xfb
    "11110110", --  757 - 0x2f5  :  246 - 0xf6
    "11111111", --  758 - 0x2f6  :  255 - 0xff
    "11111111", --  759 - 0x2f7  :  255 - 0xff
    "11111111", --  760 - 0x2f8  :  255 - 0xff
    "11111111", --  761 - 0x2f9  :  255 - 0xff
    "11111111", --  762 - 0x2fa  :  255 - 0xff
    "11111111", --  763 - 0x2fb  :  255 - 0xff
    "11101100", --  764 - 0x2fc  :  236 - 0xec
    "11111001", --  765 - 0x2fd  :  249 - 0xf9
    "11111010", --  766 - 0x2fe  :  250 - 0xfa
    "11111010", --  767 - 0x2ff  :  250 - 0xfa
    "11111010", --  768 - 0x300  :  250 - 0xfa -- line 0x18
    "11111010", --  769 - 0x301  :  250 - 0xfa
    "11111010", --  770 - 0x302  :  250 - 0xfa
    "11111010", --  771 - 0x303  :  250 - 0xfa
    "11111001", --  772 - 0x304  :  249 - 0xf9
    "11111010", --  773 - 0x305  :  250 - 0xfa
    "11111010", --  774 - 0x306  :  250 - 0xfa
    "11111010", --  775 - 0x307  :  250 - 0xfa
    "11111010", --  776 - 0x308  :  250 - 0xfa
    "11111010", --  777 - 0x309  :  250 - 0xfa
    "11111010", --  778 - 0x30a  :  250 - 0xfa
    "11111001", --  779 - 0x30b  :  249 - 0xf9
    "11111010", --  780 - 0x30c  :  250 - 0xfa
    "11111100", --  781 - 0x30d  :  252 - 0xfc
    "11111111", --  782 - 0x30e  :  255 - 0xff
    "11111111", --  783 - 0x30f  :  255 - 0xff
    "11111111", --  784 - 0x310  :  255 - 0xff
    "11111111", --  785 - 0x311  :  255 - 0xff
    "11111111", --  786 - 0x312  :  255 - 0xff
    "11111111", --  787 - 0x313  :  255 - 0xff
    "11111111", --  788 - 0x314  :  255 - 0xff
    "11111111", --  789 - 0x315  :  255 - 0xff
    "11111111", --  790 - 0x316  :  255 - 0xff
    "11111110", --  791 - 0x317  :  254 - 0xfe
    "11111110", --  792 - 0x318  :  254 - 0xfe
    "11111111", --  793 - 0x319  :  255 - 0xff
    "11100101", --  794 - 0x31a  :  229 - 0xe5
    "11101011", --  795 - 0x31b  :  235 - 0xeb
    "11111000", --  796 - 0x31c  :  248 - 0xf8
    "11111010", --  797 - 0x31d  :  250 - 0xfa
    "11111010", --  798 - 0x31e  :  250 - 0xfa
    "11101001", --  799 - 0x31f  :  233 - 0xe9
    "11101010", --  800 - 0x320  :  234 - 0xea -- line 0x19
    "11111010", --  801 - 0x321  :  250 - 0xfa
    "11111010", --  802 - 0x322  :  250 - 0xfa
    "11111010", --  803 - 0x323  :  250 - 0xfa
    "11111010", --  804 - 0x324  :  250 - 0xfa
    "11111010", --  805 - 0x325  :  250 - 0xfa
    "11111001", --  806 - 0x326  :  249 - 0xf9
    "11111001", --  807 - 0x327  :  249 - 0xf9
    "11111010", --  808 - 0x328  :  250 - 0xfa
    "11111010", --  809 - 0x329  :  250 - 0xfa
    "11111010", --  810 - 0x32a  :  250 - 0xfa
    "11101010", --  811 - 0x32b  :  234 - 0xea
    "11111010", --  812 - 0x32c  :  250 - 0xfa
    "11111100", --  813 - 0x32d  :  252 - 0xfc
    "11111111", --  814 - 0x32e  :  255 - 0xff
    "11111111", --  815 - 0x32f  :  255 - 0xff
    "11111111", --  816 - 0x330  :  255 - 0xff
    "11111101", --  817 - 0x331  :  253 - 0xfd
    "11111111", --  818 - 0x332  :  255 - 0xff
    "11111101", --  819 - 0x333  :  253 - 0xfd
    "11111111", --  820 - 0x334  :  255 - 0xff
    "11111101", --  821 - 0x335  :  253 - 0xfd
    "11111111", --  822 - 0x336  :  255 - 0xff
    "11111111", --  823 - 0x337  :  255 - 0xff
    "11111111", --  824 - 0x338  :  255 - 0xff
    "11111111", --  825 - 0x339  :  255 - 0xff
    "11101100", --  826 - 0x33a  :  236 - 0xec
    "11111010", --  827 - 0x33b  :  250 - 0xfa
    "11111010", --  828 - 0x33c  :  250 - 0xfa
    "11111010", --  829 - 0x33d  :  250 - 0xfa
    "11111010", --  830 - 0x33e  :  250 - 0xfa
    "11111010", --  831 - 0x33f  :  250 - 0xfa
    "11111010", --  832 - 0x340  :  250 - 0xfa -- line 0x1a
    "11111010", --  833 - 0x341  :  250 - 0xfa
    "11111010", --  834 - 0x342  :  250 - 0xfa
    "11111010", --  835 - 0x343  :  250 - 0xfa
    "11101010", --  836 - 0x344  :  234 - 0xea
    "11111010", --  837 - 0x345  :  250 - 0xfa
    "11111010", --  838 - 0x346  :  250 - 0xfa
    "11111010", --  839 - 0x347  :  250 - 0xfa
    "11111010", --  840 - 0x348  :  250 - 0xfa
    "11111001", --  841 - 0x349  :  249 - 0xf9
    "11111010", --  842 - 0x34a  :  250 - 0xfa
    "11111010", --  843 - 0x34b  :  250 - 0xfa
    "11111010", --  844 - 0x34c  :  250 - 0xfa
    "11111100", --  845 - 0x34d  :  252 - 0xfc
    "11111111", --  846 - 0x34e  :  255 - 0xff
    "11111111", --  847 - 0x34f  :  255 - 0xff
    "11111111", --  848 - 0x350  :  255 - 0xff
    "11111101", --  849 - 0x351  :  253 - 0xfd
    "11111111", --  850 - 0x352  :  255 - 0xff
    "11111101", --  851 - 0x353  :  253 - 0xfd
    "11111111", --  852 - 0x354  :  255 - 0xff
    "11111101", --  853 - 0x355  :  253 - 0xfd
    "11111111", --  854 - 0x356  :  255 - 0xff
    "11111111", --  855 - 0x357  :  255 - 0xff
    "11111111", --  856 - 0x358  :  255 - 0xff
    "11111111", --  857 - 0x359  :  255 - 0xff
    "11101100", --  858 - 0x35a  :  236 - 0xec
    "11111010", --  859 - 0x35b  :  250 - 0xfa
    "11111010", --  860 - 0x35c  :  250 - 0xfa
    "11101010", --  861 - 0x35d  :  234 - 0xea
    "11111010", --  862 - 0x35e  :  250 - 0xfa
    "11111010", --  863 - 0x35f  :  250 - 0xfa
    "11111010", --  864 - 0x360  :  250 - 0xfa -- line 0x1b
    "11111010", --  865 - 0x361  :  250 - 0xfa
    "11111010", --  866 - 0x362  :  250 - 0xfa
    "11111010", --  867 - 0x363  :  250 - 0xfa
    "11111010", --  868 - 0x364  :  250 - 0xfa
    "11111010", --  869 - 0x365  :  250 - 0xfa
    "11111010", --  870 - 0x366  :  250 - 0xfa
    "11111010", --  871 - 0x367  :  250 - 0xfa
    "11111010", --  872 - 0x368  :  250 - 0xfa
    "11111010", --  873 - 0x369  :  250 - 0xfa
    "11111010", --  874 - 0x36a  :  250 - 0xfa
    "11111010", --  875 - 0x36b  :  250 - 0xfa
    "11111010", --  876 - 0x36c  :  250 - 0xfa
    "11111100", --  877 - 0x36d  :  252 - 0xfc
    "11111111", --  878 - 0x36e  :  255 - 0xff
    "11111111", --  879 - 0x36f  :  255 - 0xff
    "11111111", --  880 - 0x370  :  255 - 0xff
    "11111111", --  881 - 0x371  :  255 - 0xff
    "11111111", --  882 - 0x372  :  255 - 0xff
    "11111111", --  883 - 0x373  :  255 - 0xff
    "11111111", --  884 - 0x374  :  255 - 0xff
    "11111111", --  885 - 0x375  :  255 - 0xff
    "11111111", --  886 - 0x376  :  255 - 0xff
    "11111111", --  887 - 0x377  :  255 - 0xff
    "11111111", --  888 - 0x378  :  255 - 0xff
    "11111111", --  889 - 0x379  :  255 - 0xff
    "11101100", --  890 - 0x37a  :  236 - 0xec
    "11111010", --  891 - 0x37b  :  250 - 0xfa
    "11111010", --  892 - 0x37c  :  250 - 0xfa
    "11111010", --  893 - 0x37d  :  250 - 0xfa
    "11111010", --  894 - 0x37e  :  250 - 0xfa
    "11111001", --  895 - 0x37f  :  249 - 0xf9
    "11111010", --  896 - 0x380  :  250 - 0xfa -- line 0x1c
    "11111010", --  897 - 0x381  :  250 - 0xfa
    "11111010", --  898 - 0x382  :  250 - 0xfa
    "11111010", --  899 - 0x383  :  250 - 0xfa
    "11111010", --  900 - 0x384  :  250 - 0xfa
    "11111010", --  901 - 0x385  :  250 - 0xfa
    "11111001", --  902 - 0x386  :  249 - 0xf9
    "11111010", --  903 - 0x387  :  250 - 0xfa
    "11111010", --  904 - 0x388  :  250 - 0xfa
    "11111010", --  905 - 0x389  :  250 - 0xfa
    "11111001", --  906 - 0x38a  :  249 - 0xf9
    "11111010", --  907 - 0x38b  :  250 - 0xfa
    "11111010", --  908 - 0x38c  :  250 - 0xfa
    "11110111", --  909 - 0x38d  :  247 - 0xf7
    "11101011", --  910 - 0x38e  :  235 - 0xeb
    "11101011", --  911 - 0x38f  :  235 - 0xeb
    "11101011", --  912 - 0x390  :  235 - 0xeb
    "11101011", --  913 - 0x391  :  235 - 0xeb
    "11101011", --  914 - 0x392  :  235 - 0xeb
    "11101011", --  915 - 0x393  :  235 - 0xeb
    "11101011", --  916 - 0x394  :  235 - 0xeb
    "11101011", --  917 - 0x395  :  235 - 0xeb
    "11101011", --  918 - 0x396  :  235 - 0xeb
    "11101011", --  919 - 0x397  :  235 - 0xeb
    "11101011", --  920 - 0x398  :  235 - 0xeb
    "11101011", --  921 - 0x399  :  235 - 0xeb
    "11111000", --  922 - 0x39a  :  248 - 0xf8
    "11111010", --  923 - 0x39b  :  250 - 0xfa
    "11111010", --  924 - 0x39c  :  250 - 0xfa
    "11111010", --  925 - 0x39d  :  250 - 0xfa
    "11111010", --  926 - 0x39e  :  250 - 0xfa
    "11111010", --  927 - 0x39f  :  250 - 0xfa
    "11111010", --  928 - 0x3a0  :  250 - 0xfa -- line 0x1d
    "11111001", --  929 - 0x3a1  :  249 - 0xf9
    "11111010", --  930 - 0x3a2  :  250 - 0xfa
    "11111010", --  931 - 0x3a3  :  250 - 0xfa
    "11111010", --  932 - 0x3a4  :  250 - 0xfa
    "11111010", --  933 - 0x3a5  :  250 - 0xfa
    "11111010", --  934 - 0x3a6  :  250 - 0xfa
    "11111010", --  935 - 0x3a7  :  250 - 0xfa
    "11111010", --  936 - 0x3a8  :  250 - 0xfa
    "11111010", --  937 - 0x3a9  :  250 - 0xfa
    "11111010", --  938 - 0x3aa  :  250 - 0xfa
    "11111010", --  939 - 0x3ab  :  250 - 0xfa
    "11111010", --  940 - 0x3ac  :  250 - 0xfa
    "11111010", --  941 - 0x3ad  :  250 - 0xfa
    "11111010", --  942 - 0x3ae  :  250 - 0xfa
    "11111010", --  943 - 0x3af  :  250 - 0xfa
    "11111010", --  944 - 0x3b0  :  250 - 0xfa
    "11111010", --  945 - 0x3b1  :  250 - 0xfa
    "11111010", --  946 - 0x3b2  :  250 - 0xfa
    "11111010", --  947 - 0x3b3  :  250 - 0xfa
    "11111010", --  948 - 0x3b4  :  250 - 0xfa
    "11101001", --  949 - 0x3b5  :  233 - 0xe9
    "11111010", --  950 - 0x3b6  :  250 - 0xfa
    "11111010", --  951 - 0x3b7  :  250 - 0xfa
    "11111010", --  952 - 0x3b8  :  250 - 0xfa
    "11111010", --  953 - 0x3b9  :  250 - 0xfa
    "11111010", --  954 - 0x3ba  :  250 - 0xfa
    "11111010", --  955 - 0x3bb  :  250 - 0xfa
    "11101010", --  956 - 0x3bc  :  234 - 0xea
    "11111010", --  957 - 0x3bd  :  250 - 0xfa
    "11111010", --  958 - 0x3be  :  250 - 0xfa
    "11111010", --  959 - 0x3bf  :  250 - 0xfa
        ---- Attribute Table 0----
    "00010101", --  960 - 0x3c0  :   21 - 0x15
    "00000101", --  961 - 0x3c1  :    5 - 0x5
    "00000101", --  962 - 0x3c2  :    5 - 0x5
    "00000101", --  963 - 0x3c3  :    5 - 0x5
    "00000101", --  964 - 0x3c4  :    5 - 0x5
    "00000101", --  965 - 0x3c5  :    5 - 0x5
    "01000101", --  966 - 0x3c6  :   69 - 0x45
    "01010101", --  967 - 0x3c7  :   85 - 0x55
    "00010001", --  968 - 0x3c8  :   17 - 0x11
    "01000000", --  969 - 0x3c9  :   64 - 0x40
    "01010000", --  970 - 0x3ca  :   80 - 0x50
    "01010000", --  971 - 0x3cb  :   80 - 0x50
    "01010000", --  972 - 0x3cc  :   80 - 0x50
    "01010000", --  973 - 0x3cd  :   80 - 0x50
    "00000000", --  974 - 0x3ce  :    0 - 0x0
    "01000100", --  975 - 0x3cf  :   68 - 0x44
    "00010001", --  976 - 0x3d0  :   17 - 0x11
    "01000100", --  977 - 0x3d1  :   68 - 0x44
    "00000000", --  978 - 0x3d2  :    0 - 0x0
    "00000000", --  979 - 0x3d3  :    0 - 0x0
    "00000000", --  980 - 0x3d4  :    0 - 0x0
    "01000100", --  981 - 0x3d5  :   68 - 0x44
    "00010001", --  982 - 0x3d6  :   17 - 0x11
    "01000100", --  983 - 0x3d7  :   68 - 0x44
    "00010001", --  984 - 0x3d8  :   17 - 0x11
    "01000100", --  985 - 0x3d9  :   68 - 0x44
    "00000000", --  986 - 0x3da  :    0 - 0x0
    "00010101", --  987 - 0x3db  :   21 - 0x15
    "00000001", --  988 - 0x3dc  :    1 - 0x1
    "01000100", --  989 - 0x3dd  :   68 - 0x44
    "00010001", --  990 - 0x3de  :   17 - 0x11
    "01000100", --  991 - 0x3df  :   68 - 0x44
    "00010001", --  992 - 0x3e0  :   17 - 0x11
    "00000100", --  993 - 0x3e1  :    4 - 0x4
    "00000000", --  994 - 0x3e2  :    0 - 0x0
    "00010001", --  995 - 0x3e3  :   17 - 0x11
    "01000000", --  996 - 0x3e4  :   64 - 0x40
    "01010100", --  997 - 0x3e5  :   84 - 0x54
    "00000000", --  998 - 0x3e6  :    0 - 0x0
    "01010100", --  999 - 0x3e7  :   84 - 0x54
    "01010001", -- 1000 - 0x3e8  :   81 - 0x51
    "01010000", -- 1001 - 0x3e9  :   80 - 0x50
    "01010000", -- 1002 - 0x3ea  :   80 - 0x50
    "00010001", -- 1003 - 0x3eb  :   17 - 0x11
    "01000100", -- 1004 - 0x3ec  :   68 - 0x44
    "00010001", -- 1005 - 0x3ed  :   17 - 0x11
    "00000000", -- 1006 - 0x3ee  :    0 - 0x0
    "01010101", -- 1007 - 0x3ef  :   85 - 0x55
    "01010101", -- 1008 - 0x3f0  :   85 - 0x55
    "01010101", -- 1009 - 0x3f1  :   85 - 0x55
    "01010101", -- 1010 - 0x3f2  :   85 - 0x55
    "00010001", -- 1011 - 0x3f3  :   17 - 0x11
    "00000000", -- 1012 - 0x3f4  :    0 - 0x0
    "00000000", -- 1013 - 0x3f5  :    0 - 0x0
    "01000100", -- 1014 - 0x3f6  :   68 - 0x44
    "01010101", -- 1015 - 0x3f7  :   85 - 0x55
    "00000101", -- 1016 - 0x3f8  :    5 - 0x5
    "00000101", -- 1017 - 0x3f9  :    5 - 0x5
    "00000101", -- 1018 - 0x3fa  :    5 - 0x5
    "00000101", -- 1019 - 0x3fb  :    5 - 0x5
    "00000101", -- 1020 - 0x3fc  :    5 - 0x5
    "00000101", -- 1021 - 0x3fd  :    5 - 0x5
    "00000101", -- 1022 - 0x3fe  :    5 - 0x5
    "00000101"  -- 1023 - 0x3ff  :    5 - 0x5
    );
begin
  addr_int <= to_integer(unsigned(addr));
  P_ROM: process(clk)
  begin
    if clk'event and clk='1' then
      dout <= table_mem(addr_int);
    end if;
  end process;
end BEHAVIORAL;
