//- Autcmatically generated verilog ROM from a NES memory file----
//-   NAME TABLE
// https://wiki.nesdev.com/w/index.php/PPU_nametables


//-  Original memory dump file name: smario_ntable_01.dmp --
//---- Felipe Machado -----------------------------------
//---- Area de Tecnologia Electronica -----------
//---- Universidad Rey Juan Carlos ----------------------
//---- https://github.com/felipe-m ----------------------
//-------------------------------------------------------
//--- Memory with clock ------

//--- Ports ---------------------------------------------
// Inputs   ---------------------------------------------
//    clk  :  clock signal
//    addr :  memory address
// Outputs  ---------------------------------------------
//    dout :  memory data out  (a clock cycle later)




module ROM_NTABLE_SMARIO_01
  (
     input     clk,   // clock
     input      [11-1:0] addr,  //2048 memory positions
     output reg  [8-1:0] dout  // memory data width
  );


  always @(posedge clk)
  begin
    case (addr)
                               //  address:   value 
                               //    dec  : dec - hex
     //----- Name Table 0---------
      11'h0: dout <= 8'b00100100; //    0 :  36 - 0x24 -- line 0x0
      11'h1: dout <= 8'b00100100; //    1 :  36 - 0x24
      11'h2: dout <= 8'b00100100; //    2 :  36 - 0x24
      11'h3: dout <= 8'b00100100; //    3 :  36 - 0x24
      11'h4: dout <= 8'b00100100; //    4 :  36 - 0x24
      11'h5: dout <= 8'b00100100; //    5 :  36 - 0x24
      11'h6: dout <= 8'b00100100; //    6 :  36 - 0x24
      11'h7: dout <= 8'b00100100; //    7 :  36 - 0x24
      11'h8: dout <= 8'b00100100; //    8 :  36 - 0x24
      11'h9: dout <= 8'b00100100; //    9 :  36 - 0x24
      11'hA: dout <= 8'b00100100; //   10 :  36 - 0x24
      11'hB: dout <= 8'b00100100; //   11 :  36 - 0x24
      11'hC: dout <= 8'b00100100; //   12 :  36 - 0x24
      11'hD: dout <= 8'b00100100; //   13 :  36 - 0x24
      11'hE: dout <= 8'b00100100; //   14 :  36 - 0x24
      11'hF: dout <= 8'b00100100; //   15 :  36 - 0x24
      11'h10: dout <= 8'b00100100; //   16 :  36 - 0x24
      11'h11: dout <= 8'b00100100; //   17 :  36 - 0x24
      11'h12: dout <= 8'b00100100; //   18 :  36 - 0x24
      11'h13: dout <= 8'b00100100; //   19 :  36 - 0x24
      11'h14: dout <= 8'b00100100; //   20 :  36 - 0x24
      11'h15: dout <= 8'b00100100; //   21 :  36 - 0x24
      11'h16: dout <= 8'b00100100; //   22 :  36 - 0x24
      11'h17: dout <= 8'b00100100; //   23 :  36 - 0x24
      11'h18: dout <= 8'b00100100; //   24 :  36 - 0x24
      11'h19: dout <= 8'b00100100; //   25 :  36 - 0x24
      11'h1A: dout <= 8'b00100100; //   26 :  36 - 0x24
      11'h1B: dout <= 8'b00100100; //   27 :  36 - 0x24
      11'h1C: dout <= 8'b00100100; //   28 :  36 - 0x24
      11'h1D: dout <= 8'b00100100; //   29 :  36 - 0x24
      11'h1E: dout <= 8'b00100100; //   30 :  36 - 0x24
      11'h1F: dout <= 8'b00100100; //   31 :  36 - 0x24
      11'h20: dout <= 8'b00100100; //   32 :  36 - 0x24 -- line 0x1
      11'h21: dout <= 8'b00100100; //   33 :  36 - 0x24
      11'h22: dout <= 8'b00100100; //   34 :  36 - 0x24
      11'h23: dout <= 8'b00100100; //   35 :  36 - 0x24
      11'h24: dout <= 8'b00100100; //   36 :  36 - 0x24
      11'h25: dout <= 8'b00100100; //   37 :  36 - 0x24
      11'h26: dout <= 8'b00100100; //   38 :  36 - 0x24
      11'h27: dout <= 8'b00100100; //   39 :  36 - 0x24
      11'h28: dout <= 8'b00100100; //   40 :  36 - 0x24
      11'h29: dout <= 8'b00100100; //   41 :  36 - 0x24
      11'h2A: dout <= 8'b00100100; //   42 :  36 - 0x24
      11'h2B: dout <= 8'b00100100; //   43 :  36 - 0x24
      11'h2C: dout <= 8'b00100100; //   44 :  36 - 0x24
      11'h2D: dout <= 8'b00100100; //   45 :  36 - 0x24
      11'h2E: dout <= 8'b00100100; //   46 :  36 - 0x24
      11'h2F: dout <= 8'b00100100; //   47 :  36 - 0x24
      11'h30: dout <= 8'b00100100; //   48 :  36 - 0x24
      11'h31: dout <= 8'b00100100; //   49 :  36 - 0x24
      11'h32: dout <= 8'b00100100; //   50 :  36 - 0x24
      11'h33: dout <= 8'b00100100; //   51 :  36 - 0x24
      11'h34: dout <= 8'b00100100; //   52 :  36 - 0x24
      11'h35: dout <= 8'b00100100; //   53 :  36 - 0x24
      11'h36: dout <= 8'b00100100; //   54 :  36 - 0x24
      11'h37: dout <= 8'b00100100; //   55 :  36 - 0x24
      11'h38: dout <= 8'b00100100; //   56 :  36 - 0x24
      11'h39: dout <= 8'b00100100; //   57 :  36 - 0x24
      11'h3A: dout <= 8'b00100100; //   58 :  36 - 0x24
      11'h3B: dout <= 8'b00100100; //   59 :  36 - 0x24
      11'h3C: dout <= 8'b00100100; //   60 :  36 - 0x24
      11'h3D: dout <= 8'b00100100; //   61 :  36 - 0x24
      11'h3E: dout <= 8'b00100100; //   62 :  36 - 0x24
      11'h3F: dout <= 8'b00100100; //   63 :  36 - 0x24
      11'h40: dout <= 8'b00100100; //   64 :  36 - 0x24 -- line 0x2
      11'h41: dout <= 8'b00100100; //   65 :  36 - 0x24
      11'h42: dout <= 8'b00100100; //   66 :  36 - 0x24
      11'h43: dout <= 8'b00010110; //   67 :  22 - 0x16
      11'h44: dout <= 8'b00001010; //   68 :  10 - 0xa
      11'h45: dout <= 8'b00011011; //   69 :  27 - 0x1b
      11'h46: dout <= 8'b00010010; //   70 :  18 - 0x12
      11'h47: dout <= 8'b00011000; //   71 :  24 - 0x18
      11'h48: dout <= 8'b00100100; //   72 :  36 - 0x24
      11'h49: dout <= 8'b00100100; //   73 :  36 - 0x24
      11'h4A: dout <= 8'b00100100; //   74 :  36 - 0x24
      11'h4B: dout <= 8'b00100100; //   75 :  36 - 0x24
      11'h4C: dout <= 8'b00100100; //   76 :  36 - 0x24
      11'h4D: dout <= 8'b00100100; //   77 :  36 - 0x24
      11'h4E: dout <= 8'b00100100; //   78 :  36 - 0x24
      11'h4F: dout <= 8'b00100100; //   79 :  36 - 0x24
      11'h50: dout <= 8'b00100100; //   80 :  36 - 0x24
      11'h51: dout <= 8'b00100100; //   81 :  36 - 0x24
      11'h52: dout <= 8'b00100000; //   82 :  32 - 0x20
      11'h53: dout <= 8'b00011000; //   83 :  24 - 0x18
      11'h54: dout <= 8'b00011011; //   84 :  27 - 0x1b
      11'h55: dout <= 8'b00010101; //   85 :  21 - 0x15
      11'h56: dout <= 8'b00001101; //   86 :  13 - 0xd
      11'h57: dout <= 8'b00100100; //   87 :  36 - 0x24
      11'h58: dout <= 8'b00100100; //   88 :  36 - 0x24
      11'h59: dout <= 8'b00011101; //   89 :  29 - 0x1d
      11'h5A: dout <= 8'b00010010; //   90 :  18 - 0x12
      11'h5B: dout <= 8'b00010110; //   91 :  22 - 0x16
      11'h5C: dout <= 8'b00001110; //   92 :  14 - 0xe
      11'h5D: dout <= 8'b00100100; //   93 :  36 - 0x24
      11'h5E: dout <= 8'b00100100; //   94 :  36 - 0x24
      11'h5F: dout <= 8'b00100100; //   95 :  36 - 0x24
      11'h60: dout <= 8'b00100100; //   96 :  36 - 0x24 -- line 0x3
      11'h61: dout <= 8'b00100100; //   97 :  36 - 0x24
      11'h62: dout <= 8'b00100100; //   98 :  36 - 0x24
      11'h63: dout <= 8'b00000000; //   99 :   0 - 0x0
      11'h64: dout <= 8'b00000000; //  100 :   0 - 0x0
      11'h65: dout <= 8'b00000000; //  101 :   0 - 0x0
      11'h66: dout <= 8'b00000000; //  102 :   0 - 0x0
      11'h67: dout <= 8'b00000000; //  103 :   0 - 0x0
      11'h68: dout <= 8'b00000000; //  104 :   0 - 0x0
      11'h69: dout <= 8'b00100100; //  105 :  36 - 0x24
      11'h6A: dout <= 8'b00100100; //  106 :  36 - 0x24
      11'h6B: dout <= 8'b00101110; //  107 :  46 - 0x2e
      11'h6C: dout <= 8'b00101001; //  108 :  41 - 0x29
      11'h6D: dout <= 8'b00000000; //  109 :   0 - 0x0
      11'h6E: dout <= 8'b00000000; //  110 :   0 - 0x0
      11'h6F: dout <= 8'b00100100; //  111 :  36 - 0x24
      11'h70: dout <= 8'b00100100; //  112 :  36 - 0x24
      11'h71: dout <= 8'b00100100; //  113 :  36 - 0x24
      11'h72: dout <= 8'b00100100; //  114 :  36 - 0x24
      11'h73: dout <= 8'b00000001; //  115 :   1 - 0x1
      11'h74: dout <= 8'b00101000; //  116 :  40 - 0x28
      11'h75: dout <= 8'b00000001; //  117 :   1 - 0x1
      11'h76: dout <= 8'b00100100; //  118 :  36 - 0x24
      11'h77: dout <= 8'b00100100; //  119 :  36 - 0x24
      11'h78: dout <= 8'b00100100; //  120 :  36 - 0x24
      11'h79: dout <= 8'b00100100; //  121 :  36 - 0x24
      11'h7A: dout <= 8'b00100100; //  122 :  36 - 0x24
      11'h7B: dout <= 8'b00100100; //  123 :  36 - 0x24
      11'h7C: dout <= 8'b00100100; //  124 :  36 - 0x24
      11'h7D: dout <= 8'b00100100; //  125 :  36 - 0x24
      11'h7E: dout <= 8'b00100100; //  126 :  36 - 0x24
      11'h7F: dout <= 8'b00100100; //  127 :  36 - 0x24
      11'h80: dout <= 8'b00100100; //  128 :  36 - 0x24 -- line 0x4
      11'h81: dout <= 8'b00100100; //  129 :  36 - 0x24
      11'h82: dout <= 8'b00100100; //  130 :  36 - 0x24
      11'h83: dout <= 8'b00100100; //  131 :  36 - 0x24
      11'h84: dout <= 8'b00100100; //  132 :  36 - 0x24
      11'h85: dout <= 8'b01000100; //  133 :  68 - 0x44
      11'h86: dout <= 8'b01001000; //  134 :  72 - 0x48
      11'h87: dout <= 8'b01001000; //  135 :  72 - 0x48
      11'h88: dout <= 8'b01001000; //  136 :  72 - 0x48
      11'h89: dout <= 8'b01001000; //  137 :  72 - 0x48
      11'h8A: dout <= 8'b01001000; //  138 :  72 - 0x48
      11'h8B: dout <= 8'b01001000; //  139 :  72 - 0x48
      11'h8C: dout <= 8'b01001000; //  140 :  72 - 0x48
      11'h8D: dout <= 8'b01001000; //  141 :  72 - 0x48
      11'h8E: dout <= 8'b01001000; //  142 :  72 - 0x48
      11'h8F: dout <= 8'b01001000; //  143 :  72 - 0x48
      11'h90: dout <= 8'b01001000; //  144 :  72 - 0x48
      11'h91: dout <= 8'b01001000; //  145 :  72 - 0x48
      11'h92: dout <= 8'b01001000; //  146 :  72 - 0x48
      11'h93: dout <= 8'b01001000; //  147 :  72 - 0x48
      11'h94: dout <= 8'b01001000; //  148 :  72 - 0x48
      11'h95: dout <= 8'b01001000; //  149 :  72 - 0x48
      11'h96: dout <= 8'b01001000; //  150 :  72 - 0x48
      11'h97: dout <= 8'b01001000; //  151 :  72 - 0x48
      11'h98: dout <= 8'b01001000; //  152 :  72 - 0x48
      11'h99: dout <= 8'b01001000; //  153 :  72 - 0x48
      11'h9A: dout <= 8'b01001001; //  154 :  73 - 0x49
      11'h9B: dout <= 8'b00100100; //  155 :  36 - 0x24
      11'h9C: dout <= 8'b00100100; //  156 :  36 - 0x24
      11'h9D: dout <= 8'b00100100; //  157 :  36 - 0x24
      11'h9E: dout <= 8'b00100100; //  158 :  36 - 0x24
      11'h9F: dout <= 8'b00100100; //  159 :  36 - 0x24
      11'hA0: dout <= 8'b00100100; //  160 :  36 - 0x24 -- line 0x5
      11'hA1: dout <= 8'b00100100; //  161 :  36 - 0x24
      11'hA2: dout <= 8'b00100100; //  162 :  36 - 0x24
      11'hA3: dout <= 8'b00100100; //  163 :  36 - 0x24
      11'hA4: dout <= 8'b00100100; //  164 :  36 - 0x24
      11'hA5: dout <= 8'b01000110; //  165 :  70 - 0x46
      11'hA6: dout <= 8'b11010000; //  166 : 208 - 0xd0
      11'hA7: dout <= 8'b11010001; //  167 : 209 - 0xd1
      11'hA8: dout <= 8'b11011000; //  168 : 216 - 0xd8
      11'hA9: dout <= 8'b11011000; //  169 : 216 - 0xd8
      11'hAA: dout <= 8'b11011110; //  170 : 222 - 0xde
      11'hAB: dout <= 8'b11010001; //  171 : 209 - 0xd1
      11'hAC: dout <= 8'b11010000; //  172 : 208 - 0xd0
      11'hAD: dout <= 8'b11011010; //  173 : 218 - 0xda
      11'hAE: dout <= 8'b11011110; //  174 : 222 - 0xde
      11'hAF: dout <= 8'b11010001; //  175 : 209 - 0xd1
      11'hB0: dout <= 8'b00100110; //  176 :  38 - 0x26
      11'hB1: dout <= 8'b00100110; //  177 :  38 - 0x26
      11'hB2: dout <= 8'b00100110; //  178 :  38 - 0x26
      11'hB3: dout <= 8'b00100110; //  179 :  38 - 0x26
      11'hB4: dout <= 8'b00100110; //  180 :  38 - 0x26
      11'hB5: dout <= 8'b00100110; //  181 :  38 - 0x26
      11'hB6: dout <= 8'b00100110; //  182 :  38 - 0x26
      11'hB7: dout <= 8'b00100110; //  183 :  38 - 0x26
      11'hB8: dout <= 8'b00100110; //  184 :  38 - 0x26
      11'hB9: dout <= 8'b00100110; //  185 :  38 - 0x26
      11'hBA: dout <= 8'b01001010; //  186 :  74 - 0x4a
      11'hBB: dout <= 8'b00100100; //  187 :  36 - 0x24
      11'hBC: dout <= 8'b00100100; //  188 :  36 - 0x24
      11'hBD: dout <= 8'b00100100; //  189 :  36 - 0x24
      11'hBE: dout <= 8'b00100100; //  190 :  36 - 0x24
      11'hBF: dout <= 8'b00100100; //  191 :  36 - 0x24
      11'hC0: dout <= 8'b00100100; //  192 :  36 - 0x24 -- line 0x6
      11'hC1: dout <= 8'b00100100; //  193 :  36 - 0x24
      11'hC2: dout <= 8'b00100100; //  194 :  36 - 0x24
      11'hC3: dout <= 8'b00100100; //  195 :  36 - 0x24
      11'hC4: dout <= 8'b00100100; //  196 :  36 - 0x24
      11'hC5: dout <= 8'b01000110; //  197 :  70 - 0x46
      11'hC6: dout <= 8'b11010010; //  198 : 210 - 0xd2
      11'hC7: dout <= 8'b11010011; //  199 : 211 - 0xd3
      11'hC8: dout <= 8'b11011011; //  200 : 219 - 0xdb
      11'hC9: dout <= 8'b11011011; //  201 : 219 - 0xdb
      11'hCA: dout <= 8'b11011011; //  202 : 219 - 0xdb
      11'hCB: dout <= 8'b11011001; //  203 : 217 - 0xd9
      11'hCC: dout <= 8'b11011011; //  204 : 219 - 0xdb
      11'hCD: dout <= 8'b11011100; //  205 : 220 - 0xdc
      11'hCE: dout <= 8'b11011011; //  206 : 219 - 0xdb
      11'hCF: dout <= 8'b11011111; //  207 : 223 - 0xdf
      11'hD0: dout <= 8'b00100110; //  208 :  38 - 0x26
      11'hD1: dout <= 8'b00100110; //  209 :  38 - 0x26
      11'hD2: dout <= 8'b00100110; //  210 :  38 - 0x26
      11'hD3: dout <= 8'b00100110; //  211 :  38 - 0x26
      11'hD4: dout <= 8'b00100110; //  212 :  38 - 0x26
      11'hD5: dout <= 8'b00100110; //  213 :  38 - 0x26
      11'hD6: dout <= 8'b00100110; //  214 :  38 - 0x26
      11'hD7: dout <= 8'b00100110; //  215 :  38 - 0x26
      11'hD8: dout <= 8'b00100110; //  216 :  38 - 0x26
      11'hD9: dout <= 8'b00100110; //  217 :  38 - 0x26
      11'hDA: dout <= 8'b01001010; //  218 :  74 - 0x4a
      11'hDB: dout <= 8'b00100100; //  219 :  36 - 0x24
      11'hDC: dout <= 8'b00100100; //  220 :  36 - 0x24
      11'hDD: dout <= 8'b00100100; //  221 :  36 - 0x24
      11'hDE: dout <= 8'b00100100; //  222 :  36 - 0x24
      11'hDF: dout <= 8'b00100100; //  223 :  36 - 0x24
      11'hE0: dout <= 8'b00100100; //  224 :  36 - 0x24 -- line 0x7
      11'hE1: dout <= 8'b00100100; //  225 :  36 - 0x24
      11'hE2: dout <= 8'b00100100; //  226 :  36 - 0x24
      11'hE3: dout <= 8'b00100100; //  227 :  36 - 0x24
      11'hE4: dout <= 8'b00100100; //  228 :  36 - 0x24
      11'hE5: dout <= 8'b01000110; //  229 :  70 - 0x46
      11'hE6: dout <= 8'b11010100; //  230 : 212 - 0xd4
      11'hE7: dout <= 8'b11010101; //  231 : 213 - 0xd5
      11'hE8: dout <= 8'b11010100; //  232 : 212 - 0xd4
      11'hE9: dout <= 8'b11011001; //  233 : 217 - 0xd9
      11'hEA: dout <= 8'b11011011; //  234 : 219 - 0xdb
      11'hEB: dout <= 8'b11100010; //  235 : 226 - 0xe2
      11'hEC: dout <= 8'b11010100; //  236 : 212 - 0xd4
      11'hED: dout <= 8'b11011010; //  237 : 218 - 0xda
      11'hEE: dout <= 8'b11011011; //  238 : 219 - 0xdb
      11'hEF: dout <= 8'b11100000; //  239 : 224 - 0xe0
      11'hF0: dout <= 8'b00100110; //  240 :  38 - 0x26
      11'hF1: dout <= 8'b00100110; //  241 :  38 - 0x26
      11'hF2: dout <= 8'b00100110; //  242 :  38 - 0x26
      11'hF3: dout <= 8'b00100110; //  243 :  38 - 0x26
      11'hF4: dout <= 8'b00100110; //  244 :  38 - 0x26
      11'hF5: dout <= 8'b00100110; //  245 :  38 - 0x26
      11'hF6: dout <= 8'b00100110; //  246 :  38 - 0x26
      11'hF7: dout <= 8'b00100110; //  247 :  38 - 0x26
      11'hF8: dout <= 8'b00100110; //  248 :  38 - 0x26
      11'hF9: dout <= 8'b00100110; //  249 :  38 - 0x26
      11'hFA: dout <= 8'b01001010; //  250 :  74 - 0x4a
      11'hFB: dout <= 8'b00100100; //  251 :  36 - 0x24
      11'hFC: dout <= 8'b00100100; //  252 :  36 - 0x24
      11'hFD: dout <= 8'b00100100; //  253 :  36 - 0x24
      11'hFE: dout <= 8'b00100100; //  254 :  36 - 0x24
      11'hFF: dout <= 8'b00100100; //  255 :  36 - 0x24
      11'h100: dout <= 8'b00100100; //  256 :  36 - 0x24 -- line 0x8
      11'h101: dout <= 8'b00100100; //  257 :  36 - 0x24
      11'h102: dout <= 8'b00100100; //  258 :  36 - 0x24
      11'h103: dout <= 8'b00100100; //  259 :  36 - 0x24
      11'h104: dout <= 8'b00100100; //  260 :  36 - 0x24
      11'h105: dout <= 8'b01000110; //  261 :  70 - 0x46
      11'h106: dout <= 8'b11010110; //  262 : 214 - 0xd6
      11'h107: dout <= 8'b11010111; //  263 : 215 - 0xd7
      11'h108: dout <= 8'b11010110; //  264 : 214 - 0xd6
      11'h109: dout <= 8'b11010111; //  265 : 215 - 0xd7
      11'h10A: dout <= 8'b11100001; //  266 : 225 - 0xe1
      11'h10B: dout <= 8'b00100110; //  267 :  38 - 0x26
      11'h10C: dout <= 8'b11010110; //  268 : 214 - 0xd6
      11'h10D: dout <= 8'b11011101; //  269 : 221 - 0xdd
      11'h10E: dout <= 8'b11100001; //  270 : 225 - 0xe1
      11'h10F: dout <= 8'b11100001; //  271 : 225 - 0xe1
      11'h110: dout <= 8'b00100110; //  272 :  38 - 0x26
      11'h111: dout <= 8'b00100110; //  273 :  38 - 0x26
      11'h112: dout <= 8'b00100110; //  274 :  38 - 0x26
      11'h113: dout <= 8'b00100110; //  275 :  38 - 0x26
      11'h114: dout <= 8'b00100110; //  276 :  38 - 0x26
      11'h115: dout <= 8'b00100110; //  277 :  38 - 0x26
      11'h116: dout <= 8'b00100110; //  278 :  38 - 0x26
      11'h117: dout <= 8'b00100110; //  279 :  38 - 0x26
      11'h118: dout <= 8'b00100110; //  280 :  38 - 0x26
      11'h119: dout <= 8'b00100110; //  281 :  38 - 0x26
      11'h11A: dout <= 8'b01001010; //  282 :  74 - 0x4a
      11'h11B: dout <= 8'b00100100; //  283 :  36 - 0x24
      11'h11C: dout <= 8'b00100100; //  284 :  36 - 0x24
      11'h11D: dout <= 8'b00100100; //  285 :  36 - 0x24
      11'h11E: dout <= 8'b00100100; //  286 :  36 - 0x24
      11'h11F: dout <= 8'b00100100; //  287 :  36 - 0x24
      11'h120: dout <= 8'b00100100; //  288 :  36 - 0x24 -- line 0x9
      11'h121: dout <= 8'b00100100; //  289 :  36 - 0x24
      11'h122: dout <= 8'b00100100; //  290 :  36 - 0x24
      11'h123: dout <= 8'b00100100; //  291 :  36 - 0x24
      11'h124: dout <= 8'b00100100; //  292 :  36 - 0x24
      11'h125: dout <= 8'b01000110; //  293 :  70 - 0x46
      11'h126: dout <= 8'b11010000; //  294 : 208 - 0xd0
      11'h127: dout <= 8'b11101000; //  295 : 232 - 0xe8
      11'h128: dout <= 8'b11010001; //  296 : 209 - 0xd1
      11'h129: dout <= 8'b11010000; //  297 : 208 - 0xd0
      11'h12A: dout <= 8'b11010001; //  298 : 209 - 0xd1
      11'h12B: dout <= 8'b11011110; //  299 : 222 - 0xde
      11'h12C: dout <= 8'b11010001; //  300 : 209 - 0xd1
      11'h12D: dout <= 8'b11011000; //  301 : 216 - 0xd8
      11'h12E: dout <= 8'b11010000; //  302 : 208 - 0xd0
      11'h12F: dout <= 8'b11010001; //  303 : 209 - 0xd1
      11'h130: dout <= 8'b00100110; //  304 :  38 - 0x26
      11'h131: dout <= 8'b11011110; //  305 : 222 - 0xde
      11'h132: dout <= 8'b11010001; //  306 : 209 - 0xd1
      11'h133: dout <= 8'b11011110; //  307 : 222 - 0xde
      11'h134: dout <= 8'b11010001; //  308 : 209 - 0xd1
      11'h135: dout <= 8'b11010000; //  309 : 208 - 0xd0
      11'h136: dout <= 8'b11010001; //  310 : 209 - 0xd1
      11'h137: dout <= 8'b11010000; //  311 : 208 - 0xd0
      11'h138: dout <= 8'b11010001; //  312 : 209 - 0xd1
      11'h139: dout <= 8'b00100110; //  313 :  38 - 0x26
      11'h13A: dout <= 8'b01001010; //  314 :  74 - 0x4a
      11'h13B: dout <= 8'b00100100; //  315 :  36 - 0x24
      11'h13C: dout <= 8'b00100100; //  316 :  36 - 0x24
      11'h13D: dout <= 8'b00100100; //  317 :  36 - 0x24
      11'h13E: dout <= 8'b00100100; //  318 :  36 - 0x24
      11'h13F: dout <= 8'b00100100; //  319 :  36 - 0x24
      11'h140: dout <= 8'b00100100; //  320 :  36 - 0x24 -- line 0xa
      11'h141: dout <= 8'b00100100; //  321 :  36 - 0x24
      11'h142: dout <= 8'b00100100; //  322 :  36 - 0x24
      11'h143: dout <= 8'b00100100; //  323 :  36 - 0x24
      11'h144: dout <= 8'b00100100; //  324 :  36 - 0x24
      11'h145: dout <= 8'b01000110; //  325 :  70 - 0x46
      11'h146: dout <= 8'b11011011; //  326 : 219 - 0xdb
      11'h147: dout <= 8'b01000010; //  327 :  66 - 0x42
      11'h148: dout <= 8'b01000010; //  328 :  66 - 0x42
      11'h149: dout <= 8'b11011011; //  329 : 219 - 0xdb
      11'h14A: dout <= 8'b01000010; //  330 :  66 - 0x42
      11'h14B: dout <= 8'b11011011; //  331 : 219 - 0xdb
      11'h14C: dout <= 8'b01000010; //  332 :  66 - 0x42
      11'h14D: dout <= 8'b11011011; //  333 : 219 - 0xdb
      11'h14E: dout <= 8'b11011011; //  334 : 219 - 0xdb
      11'h14F: dout <= 8'b01000010; //  335 :  66 - 0x42
      11'h150: dout <= 8'b00100110; //  336 :  38 - 0x26
      11'h151: dout <= 8'b11011011; //  337 : 219 - 0xdb
      11'h152: dout <= 8'b01000010; //  338 :  66 - 0x42
      11'h153: dout <= 8'b11011011; //  339 : 219 - 0xdb
      11'h154: dout <= 8'b01000010; //  340 :  66 - 0x42
      11'h155: dout <= 8'b11011011; //  341 : 219 - 0xdb
      11'h156: dout <= 8'b01000010; //  342 :  66 - 0x42
      11'h157: dout <= 8'b11011011; //  343 : 219 - 0xdb
      11'h158: dout <= 8'b01000010; //  344 :  66 - 0x42
      11'h159: dout <= 8'b00100110; //  345 :  38 - 0x26
      11'h15A: dout <= 8'b01001010; //  346 :  74 - 0x4a
      11'h15B: dout <= 8'b00100100; //  347 :  36 - 0x24
      11'h15C: dout <= 8'b00100100; //  348 :  36 - 0x24
      11'h15D: dout <= 8'b00100100; //  349 :  36 - 0x24
      11'h15E: dout <= 8'b00100100; //  350 :  36 - 0x24
      11'h15F: dout <= 8'b00100100; //  351 :  36 - 0x24
      11'h160: dout <= 8'b00100100; //  352 :  36 - 0x24 -- line 0xb
      11'h161: dout <= 8'b00100100; //  353 :  36 - 0x24
      11'h162: dout <= 8'b00100100; //  354 :  36 - 0x24
      11'h163: dout <= 8'b00100100; //  355 :  36 - 0x24
      11'h164: dout <= 8'b00100100; //  356 :  36 - 0x24
      11'h165: dout <= 8'b01000110; //  357 :  70 - 0x46
      11'h166: dout <= 8'b11011011; //  358 : 219 - 0xdb
      11'h167: dout <= 8'b11011011; //  359 : 219 - 0xdb
      11'h168: dout <= 8'b11011011; //  360 : 219 - 0xdb
      11'h169: dout <= 8'b11011011; //  361 : 219 - 0xdb
      11'h16A: dout <= 8'b11011011; //  362 : 219 - 0xdb
      11'h16B: dout <= 8'b11011011; //  363 : 219 - 0xdb
      11'h16C: dout <= 8'b11011111; //  364 : 223 - 0xdf
      11'h16D: dout <= 8'b11011011; //  365 : 219 - 0xdb
      11'h16E: dout <= 8'b11011011; //  366 : 219 - 0xdb
      11'h16F: dout <= 8'b11011011; //  367 : 219 - 0xdb
      11'h170: dout <= 8'b00100110; //  368 :  38 - 0x26
      11'h171: dout <= 8'b11011011; //  369 : 219 - 0xdb
      11'h172: dout <= 8'b11011111; //  370 : 223 - 0xdf
      11'h173: dout <= 8'b11011011; //  371 : 219 - 0xdb
      11'h174: dout <= 8'b11011111; //  372 : 223 - 0xdf
      11'h175: dout <= 8'b11011011; //  373 : 219 - 0xdb
      11'h176: dout <= 8'b11011011; //  374 : 219 - 0xdb
      11'h177: dout <= 8'b11100100; //  375 : 228 - 0xe4
      11'h178: dout <= 8'b11100101; //  376 : 229 - 0xe5
      11'h179: dout <= 8'b00100110; //  377 :  38 - 0x26
      11'h17A: dout <= 8'b01001010; //  378 :  74 - 0x4a
      11'h17B: dout <= 8'b00100100; //  379 :  36 - 0x24
      11'h17C: dout <= 8'b00100100; //  380 :  36 - 0x24
      11'h17D: dout <= 8'b00100100; //  381 :  36 - 0x24
      11'h17E: dout <= 8'b00100100; //  382 :  36 - 0x24
      11'h17F: dout <= 8'b00100100; //  383 :  36 - 0x24
      11'h180: dout <= 8'b00100100; //  384 :  36 - 0x24 -- line 0xc
      11'h181: dout <= 8'b00100100; //  385 :  36 - 0x24
      11'h182: dout <= 8'b00100100; //  386 :  36 - 0x24
      11'h183: dout <= 8'b00100100; //  387 :  36 - 0x24
      11'h184: dout <= 8'b00100100; //  388 :  36 - 0x24
      11'h185: dout <= 8'b01000110; //  389 :  70 - 0x46
      11'h186: dout <= 8'b11011011; //  390 : 219 - 0xdb
      11'h187: dout <= 8'b11011011; //  391 : 219 - 0xdb
      11'h188: dout <= 8'b11011011; //  392 : 219 - 0xdb
      11'h189: dout <= 8'b11011110; //  393 : 222 - 0xde
      11'h18A: dout <= 8'b01000011; //  394 :  67 - 0x43
      11'h18B: dout <= 8'b11011011; //  395 : 219 - 0xdb
      11'h18C: dout <= 8'b11100000; //  396 : 224 - 0xe0
      11'h18D: dout <= 8'b11011011; //  397 : 219 - 0xdb
      11'h18E: dout <= 8'b11011011; //  398 : 219 - 0xdb
      11'h18F: dout <= 8'b11011011; //  399 : 219 - 0xdb
      11'h190: dout <= 8'b00100110; //  400 :  38 - 0x26
      11'h191: dout <= 8'b11011011; //  401 : 219 - 0xdb
      11'h192: dout <= 8'b11100011; //  402 : 227 - 0xe3
      11'h193: dout <= 8'b11011011; //  403 : 219 - 0xdb
      11'h194: dout <= 8'b11100000; //  404 : 224 - 0xe0
      11'h195: dout <= 8'b11011011; //  405 : 219 - 0xdb
      11'h196: dout <= 8'b11011011; //  406 : 219 - 0xdb
      11'h197: dout <= 8'b11100110; //  407 : 230 - 0xe6
      11'h198: dout <= 8'b11100011; //  408 : 227 - 0xe3
      11'h199: dout <= 8'b00100110; //  409 :  38 - 0x26
      11'h19A: dout <= 8'b01001010; //  410 :  74 - 0x4a
      11'h19B: dout <= 8'b00100100; //  411 :  36 - 0x24
      11'h19C: dout <= 8'b00100100; //  412 :  36 - 0x24
      11'h19D: dout <= 8'b00100100; //  413 :  36 - 0x24
      11'h19E: dout <= 8'b00100100; //  414 :  36 - 0x24
      11'h19F: dout <= 8'b00100100; //  415 :  36 - 0x24
      11'h1A0: dout <= 8'b00100100; //  416 :  36 - 0x24 -- line 0xd
      11'h1A1: dout <= 8'b00100100; //  417 :  36 - 0x24
      11'h1A2: dout <= 8'b00100100; //  418 :  36 - 0x24
      11'h1A3: dout <= 8'b00100100; //  419 :  36 - 0x24
      11'h1A4: dout <= 8'b00100100; //  420 :  36 - 0x24
      11'h1A5: dout <= 8'b01000110; //  421 :  70 - 0x46
      11'h1A6: dout <= 8'b11011011; //  422 : 219 - 0xdb
      11'h1A7: dout <= 8'b11011011; //  423 : 219 - 0xdb
      11'h1A8: dout <= 8'b11011011; //  424 : 219 - 0xdb
      11'h1A9: dout <= 8'b11011011; //  425 : 219 - 0xdb
      11'h1AA: dout <= 8'b01000010; //  426 :  66 - 0x42
      11'h1AB: dout <= 8'b11011011; //  427 : 219 - 0xdb
      11'h1AC: dout <= 8'b11011011; //  428 : 219 - 0xdb
      11'h1AD: dout <= 8'b11011011; //  429 : 219 - 0xdb
      11'h1AE: dout <= 8'b11010100; //  430 : 212 - 0xd4
      11'h1AF: dout <= 8'b11011001; //  431 : 217 - 0xd9
      11'h1B0: dout <= 8'b00100110; //  432 :  38 - 0x26
      11'h1B1: dout <= 8'b11011011; //  433 : 219 - 0xdb
      11'h1B2: dout <= 8'b11011001; //  434 : 217 - 0xd9
      11'h1B3: dout <= 8'b11011011; //  435 : 219 - 0xdb
      11'h1B4: dout <= 8'b11011011; //  436 : 219 - 0xdb
      11'h1B5: dout <= 8'b11010100; //  437 : 212 - 0xd4
      11'h1B6: dout <= 8'b11011001; //  438 : 217 - 0xd9
      11'h1B7: dout <= 8'b11010100; //  439 : 212 - 0xd4
      11'h1B8: dout <= 8'b11011001; //  440 : 217 - 0xd9
      11'h1B9: dout <= 8'b11100111; //  441 : 231 - 0xe7
      11'h1BA: dout <= 8'b01001010; //  442 :  74 - 0x4a
      11'h1BB: dout <= 8'b00100100; //  443 :  36 - 0x24
      11'h1BC: dout <= 8'b00100100; //  444 :  36 - 0x24
      11'h1BD: dout <= 8'b00100100; //  445 :  36 - 0x24
      11'h1BE: dout <= 8'b00100100; //  446 :  36 - 0x24
      11'h1BF: dout <= 8'b00100100; //  447 :  36 - 0x24
      11'h1C0: dout <= 8'b00100100; //  448 :  36 - 0x24 -- line 0xe
      11'h1C1: dout <= 8'b00100100; //  449 :  36 - 0x24
      11'h1C2: dout <= 8'b00100100; //  450 :  36 - 0x24
      11'h1C3: dout <= 8'b00100100; //  451 :  36 - 0x24
      11'h1C4: dout <= 8'b00100100; //  452 :  36 - 0x24
      11'h1C5: dout <= 8'b01011111; //  453 :  95 - 0x5f
      11'h1C6: dout <= 8'b10010101; //  454 : 149 - 0x95
      11'h1C7: dout <= 8'b10010101; //  455 : 149 - 0x95
      11'h1C8: dout <= 8'b10010101; //  456 : 149 - 0x95
      11'h1C9: dout <= 8'b10010101; //  457 : 149 - 0x95
      11'h1CA: dout <= 8'b10010101; //  458 : 149 - 0x95
      11'h1CB: dout <= 8'b10010101; //  459 : 149 - 0x95
      11'h1CC: dout <= 8'b10010101; //  460 : 149 - 0x95
      11'h1CD: dout <= 8'b10010101; //  461 : 149 - 0x95
      11'h1CE: dout <= 8'b10010111; //  462 : 151 - 0x97
      11'h1CF: dout <= 8'b10011000; //  463 : 152 - 0x98
      11'h1D0: dout <= 8'b01111000; //  464 : 120 - 0x78
      11'h1D1: dout <= 8'b10010101; //  465 : 149 - 0x95
      11'h1D2: dout <= 8'b10010110; //  466 : 150 - 0x96
      11'h1D3: dout <= 8'b10010101; //  467 : 149 - 0x95
      11'h1D4: dout <= 8'b10010101; //  468 : 149 - 0x95
      11'h1D5: dout <= 8'b10010111; //  469 : 151 - 0x97
      11'h1D6: dout <= 8'b10011000; //  470 : 152 - 0x98
      11'h1D7: dout <= 8'b10010111; //  471 : 151 - 0x97
      11'h1D8: dout <= 8'b10011000; //  472 : 152 - 0x98
      11'h1D9: dout <= 8'b10010101; //  473 : 149 - 0x95
      11'h1DA: dout <= 8'b01111010; //  474 : 122 - 0x7a
      11'h1DB: dout <= 8'b00100100; //  475 :  36 - 0x24
      11'h1DC: dout <= 8'b00100100; //  476 :  36 - 0x24
      11'h1DD: dout <= 8'b00100100; //  477 :  36 - 0x24
      11'h1DE: dout <= 8'b00100100; //  478 :  36 - 0x24
      11'h1DF: dout <= 8'b00100100; //  479 :  36 - 0x24
      11'h1E0: dout <= 8'b00100100; //  480 :  36 - 0x24 -- line 0xf
      11'h1E1: dout <= 8'b00100100; //  481 :  36 - 0x24
      11'h1E2: dout <= 8'b00100100; //  482 :  36 - 0x24
      11'h1E3: dout <= 8'b00100100; //  483 :  36 - 0x24
      11'h1E4: dout <= 8'b00100100; //  484 :  36 - 0x24
      11'h1E5: dout <= 8'b00100100; //  485 :  36 - 0x24
      11'h1E6: dout <= 8'b00100100; //  486 :  36 - 0x24
      11'h1E7: dout <= 8'b00100100; //  487 :  36 - 0x24
      11'h1E8: dout <= 8'b00100100; //  488 :  36 - 0x24
      11'h1E9: dout <= 8'b00100100; //  489 :  36 - 0x24
      11'h1EA: dout <= 8'b00100100; //  490 :  36 - 0x24
      11'h1EB: dout <= 8'b00100100; //  491 :  36 - 0x24
      11'h1EC: dout <= 8'b00100100; //  492 :  36 - 0x24
      11'h1ED: dout <= 8'b11001111; //  493 : 207 - 0xcf
      11'h1EE: dout <= 8'b00000001; //  494 :   1 - 0x1
      11'h1EF: dout <= 8'b00001001; //  495 :   9 - 0x9
      11'h1F0: dout <= 8'b00001000; //  496 :   8 - 0x8
      11'h1F1: dout <= 8'b00000101; //  497 :   5 - 0x5
      11'h1F2: dout <= 8'b00100100; //  498 :  36 - 0x24
      11'h1F3: dout <= 8'b00010111; //  499 :  23 - 0x17
      11'h1F4: dout <= 8'b00010010; //  500 :  18 - 0x12
      11'h1F5: dout <= 8'b00010111; //  501 :  23 - 0x17
      11'h1F6: dout <= 8'b00011101; //  502 :  29 - 0x1d
      11'h1F7: dout <= 8'b00001110; //  503 :  14 - 0xe
      11'h1F8: dout <= 8'b00010111; //  504 :  23 - 0x17
      11'h1F9: dout <= 8'b00001101; //  505 :  13 - 0xd
      11'h1FA: dout <= 8'b00011000; //  506 :  24 - 0x18
      11'h1FB: dout <= 8'b00100100; //  507 :  36 - 0x24
      11'h1FC: dout <= 8'b00100100; //  508 :  36 - 0x24
      11'h1FD: dout <= 8'b00100100; //  509 :  36 - 0x24
      11'h1FE: dout <= 8'b00100100; //  510 :  36 - 0x24
      11'h1FF: dout <= 8'b00100100; //  511 :  36 - 0x24
      11'h200: dout <= 8'b00100100; //  512 :  36 - 0x24 -- line 0x10
      11'h201: dout <= 8'b00100100; //  513 :  36 - 0x24
      11'h202: dout <= 8'b00100100; //  514 :  36 - 0x24
      11'h203: dout <= 8'b00100100; //  515 :  36 - 0x24
      11'h204: dout <= 8'b00100100; //  516 :  36 - 0x24
      11'h205: dout <= 8'b00100100; //  517 :  36 - 0x24
      11'h206: dout <= 8'b00100100; //  518 :  36 - 0x24
      11'h207: dout <= 8'b00100100; //  519 :  36 - 0x24
      11'h208: dout <= 8'b00100100; //  520 :  36 - 0x24
      11'h209: dout <= 8'b00100100; //  521 :  36 - 0x24
      11'h20A: dout <= 8'b00100100; //  522 :  36 - 0x24
      11'h20B: dout <= 8'b00100100; //  523 :  36 - 0x24
      11'h20C: dout <= 8'b00100100; //  524 :  36 - 0x24
      11'h20D: dout <= 8'b00100100; //  525 :  36 - 0x24
      11'h20E: dout <= 8'b00100100; //  526 :  36 - 0x24
      11'h20F: dout <= 8'b00100100; //  527 :  36 - 0x24
      11'h210: dout <= 8'b00100100; //  528 :  36 - 0x24
      11'h211: dout <= 8'b00100100; //  529 :  36 - 0x24
      11'h212: dout <= 8'b00100100; //  530 :  36 - 0x24
      11'h213: dout <= 8'b00100100; //  531 :  36 - 0x24
      11'h214: dout <= 8'b00100100; //  532 :  36 - 0x24
      11'h215: dout <= 8'b00100100; //  533 :  36 - 0x24
      11'h216: dout <= 8'b00100100; //  534 :  36 - 0x24
      11'h217: dout <= 8'b00100100; //  535 :  36 - 0x24
      11'h218: dout <= 8'b00100100; //  536 :  36 - 0x24
      11'h219: dout <= 8'b00100100; //  537 :  36 - 0x24
      11'h21A: dout <= 8'b00100100; //  538 :  36 - 0x24
      11'h21B: dout <= 8'b00100100; //  539 :  36 - 0x24
      11'h21C: dout <= 8'b00100100; //  540 :  36 - 0x24
      11'h21D: dout <= 8'b00100100; //  541 :  36 - 0x24
      11'h21E: dout <= 8'b00100100; //  542 :  36 - 0x24
      11'h21F: dout <= 8'b00100100; //  543 :  36 - 0x24
      11'h220: dout <= 8'b00100100; //  544 :  36 - 0x24 -- line 0x11
      11'h221: dout <= 8'b00100100; //  545 :  36 - 0x24
      11'h222: dout <= 8'b00100100; //  546 :  36 - 0x24
      11'h223: dout <= 8'b00100100; //  547 :  36 - 0x24
      11'h224: dout <= 8'b00100100; //  548 :  36 - 0x24
      11'h225: dout <= 8'b00100100; //  549 :  36 - 0x24
      11'h226: dout <= 8'b00100100; //  550 :  36 - 0x24
      11'h227: dout <= 8'b00100100; //  551 :  36 - 0x24
      11'h228: dout <= 8'b00100100; //  552 :  36 - 0x24
      11'h229: dout <= 8'b00100100; //  553 :  36 - 0x24
      11'h22A: dout <= 8'b00100100; //  554 :  36 - 0x24
      11'h22B: dout <= 8'b00100100; //  555 :  36 - 0x24
      11'h22C: dout <= 8'b00100100; //  556 :  36 - 0x24
      11'h22D: dout <= 8'b00100100; //  557 :  36 - 0x24
      11'h22E: dout <= 8'b00100100; //  558 :  36 - 0x24
      11'h22F: dout <= 8'b00100100; //  559 :  36 - 0x24
      11'h230: dout <= 8'b00100100; //  560 :  36 - 0x24
      11'h231: dout <= 8'b00100100; //  561 :  36 - 0x24
      11'h232: dout <= 8'b00100100; //  562 :  36 - 0x24
      11'h233: dout <= 8'b00100100; //  563 :  36 - 0x24
      11'h234: dout <= 8'b00100100; //  564 :  36 - 0x24
      11'h235: dout <= 8'b00100100; //  565 :  36 - 0x24
      11'h236: dout <= 8'b00100100; //  566 :  36 - 0x24
      11'h237: dout <= 8'b00100100; //  567 :  36 - 0x24
      11'h238: dout <= 8'b00100100; //  568 :  36 - 0x24
      11'h239: dout <= 8'b00100100; //  569 :  36 - 0x24
      11'h23A: dout <= 8'b00100100; //  570 :  36 - 0x24
      11'h23B: dout <= 8'b00100100; //  571 :  36 - 0x24
      11'h23C: dout <= 8'b00100100; //  572 :  36 - 0x24
      11'h23D: dout <= 8'b00100100; //  573 :  36 - 0x24
      11'h23E: dout <= 8'b00100100; //  574 :  36 - 0x24
      11'h23F: dout <= 8'b00100100; //  575 :  36 - 0x24
      11'h240: dout <= 8'b00100100; //  576 :  36 - 0x24 -- line 0x12
      11'h241: dout <= 8'b00100100; //  577 :  36 - 0x24
      11'h242: dout <= 8'b00100100; //  578 :  36 - 0x24
      11'h243: dout <= 8'b00100100; //  579 :  36 - 0x24
      11'h244: dout <= 8'b00100100; //  580 :  36 - 0x24
      11'h245: dout <= 8'b00100100; //  581 :  36 - 0x24
      11'h246: dout <= 8'b00100100; //  582 :  36 - 0x24
      11'h247: dout <= 8'b00100100; //  583 :  36 - 0x24
      11'h248: dout <= 8'b00100100; //  584 :  36 - 0x24
      11'h249: dout <= 8'b11001110; //  585 : 206 - 0xce
      11'h24A: dout <= 8'b00100100; //  586 :  36 - 0x24
      11'h24B: dout <= 8'b00000001; //  587 :   1 - 0x1
      11'h24C: dout <= 8'b00100100; //  588 :  36 - 0x24
      11'h24D: dout <= 8'b00011001; //  589 :  25 - 0x19
      11'h24E: dout <= 8'b00010101; //  590 :  21 - 0x15
      11'h24F: dout <= 8'b00001010; //  591 :  10 - 0xa
      11'h250: dout <= 8'b00100010; //  592 :  34 - 0x22
      11'h251: dout <= 8'b00001110; //  593 :  14 - 0xe
      11'h252: dout <= 8'b00011011; //  594 :  27 - 0x1b
      11'h253: dout <= 8'b00100100; //  595 :  36 - 0x24
      11'h254: dout <= 8'b00010000; //  596 :  16 - 0x10
      11'h255: dout <= 8'b00001010; //  597 :  10 - 0xa
      11'h256: dout <= 8'b00010110; //  598 :  22 - 0x16
      11'h257: dout <= 8'b00001110; //  599 :  14 - 0xe
      11'h258: dout <= 8'b00100100; //  600 :  36 - 0x24
      11'h259: dout <= 8'b00100100; //  601 :  36 - 0x24
      11'h25A: dout <= 8'b00100100; //  602 :  36 - 0x24
      11'h25B: dout <= 8'b00100100; //  603 :  36 - 0x24
      11'h25C: dout <= 8'b00100100; //  604 :  36 - 0x24
      11'h25D: dout <= 8'b00100100; //  605 :  36 - 0x24
      11'h25E: dout <= 8'b00100100; //  606 :  36 - 0x24
      11'h25F: dout <= 8'b00100100; //  607 :  36 - 0x24
      11'h260: dout <= 8'b00100100; //  608 :  36 - 0x24 -- line 0x13
      11'h261: dout <= 8'b00100100; //  609 :  36 - 0x24
      11'h262: dout <= 8'b00100100; //  610 :  36 - 0x24
      11'h263: dout <= 8'b00100100; //  611 :  36 - 0x24
      11'h264: dout <= 8'b00100100; //  612 :  36 - 0x24
      11'h265: dout <= 8'b00100100; //  613 :  36 - 0x24
      11'h266: dout <= 8'b00100100; //  614 :  36 - 0x24
      11'h267: dout <= 8'b00100100; //  615 :  36 - 0x24
      11'h268: dout <= 8'b00100100; //  616 :  36 - 0x24
      11'h269: dout <= 8'b00100100; //  617 :  36 - 0x24
      11'h26A: dout <= 8'b00100100; //  618 :  36 - 0x24
      11'h26B: dout <= 8'b00100100; //  619 :  36 - 0x24
      11'h26C: dout <= 8'b00100100; //  620 :  36 - 0x24
      11'h26D: dout <= 8'b00100100; //  621 :  36 - 0x24
      11'h26E: dout <= 8'b00100100; //  622 :  36 - 0x24
      11'h26F: dout <= 8'b00100100; //  623 :  36 - 0x24
      11'h270: dout <= 8'b00100100; //  624 :  36 - 0x24
      11'h271: dout <= 8'b00100100; //  625 :  36 - 0x24
      11'h272: dout <= 8'b00100100; //  626 :  36 - 0x24
      11'h273: dout <= 8'b00100100; //  627 :  36 - 0x24
      11'h274: dout <= 8'b00100100; //  628 :  36 - 0x24
      11'h275: dout <= 8'b00100100; //  629 :  36 - 0x24
      11'h276: dout <= 8'b00100100; //  630 :  36 - 0x24
      11'h277: dout <= 8'b00100100; //  631 :  36 - 0x24
      11'h278: dout <= 8'b00100100; //  632 :  36 - 0x24
      11'h279: dout <= 8'b00100100; //  633 :  36 - 0x24
      11'h27A: dout <= 8'b00100100; //  634 :  36 - 0x24
      11'h27B: dout <= 8'b00100100; //  635 :  36 - 0x24
      11'h27C: dout <= 8'b00100100; //  636 :  36 - 0x24
      11'h27D: dout <= 8'b00100100; //  637 :  36 - 0x24
      11'h27E: dout <= 8'b00100100; //  638 :  36 - 0x24
      11'h27F: dout <= 8'b00100100; //  639 :  36 - 0x24
      11'h280: dout <= 8'b00100100; //  640 :  36 - 0x24 -- line 0x14
      11'h281: dout <= 8'b00100100; //  641 :  36 - 0x24
      11'h282: dout <= 8'b00100100; //  642 :  36 - 0x24
      11'h283: dout <= 8'b00100100; //  643 :  36 - 0x24
      11'h284: dout <= 8'b00100100; //  644 :  36 - 0x24
      11'h285: dout <= 8'b00100100; //  645 :  36 - 0x24
      11'h286: dout <= 8'b00100100; //  646 :  36 - 0x24
      11'h287: dout <= 8'b00100100; //  647 :  36 - 0x24
      11'h288: dout <= 8'b00100100; //  648 :  36 - 0x24
      11'h289: dout <= 8'b00100100; //  649 :  36 - 0x24
      11'h28A: dout <= 8'b00100100; //  650 :  36 - 0x24
      11'h28B: dout <= 8'b00000010; //  651 :   2 - 0x2
      11'h28C: dout <= 8'b00100100; //  652 :  36 - 0x24
      11'h28D: dout <= 8'b00011001; //  653 :  25 - 0x19
      11'h28E: dout <= 8'b00010101; //  654 :  21 - 0x15
      11'h28F: dout <= 8'b00001010; //  655 :  10 - 0xa
      11'h290: dout <= 8'b00100010; //  656 :  34 - 0x22
      11'h291: dout <= 8'b00001110; //  657 :  14 - 0xe
      11'h292: dout <= 8'b00011011; //  658 :  27 - 0x1b
      11'h293: dout <= 8'b00100100; //  659 :  36 - 0x24
      11'h294: dout <= 8'b00010000; //  660 :  16 - 0x10
      11'h295: dout <= 8'b00001010; //  661 :  10 - 0xa
      11'h296: dout <= 8'b00010110; //  662 :  22 - 0x16
      11'h297: dout <= 8'b00001110; //  663 :  14 - 0xe
      11'h298: dout <= 8'b00100100; //  664 :  36 - 0x24
      11'h299: dout <= 8'b00100100; //  665 :  36 - 0x24
      11'h29A: dout <= 8'b00100100; //  666 :  36 - 0x24
      11'h29B: dout <= 8'b00100100; //  667 :  36 - 0x24
      11'h29C: dout <= 8'b00100100; //  668 :  36 - 0x24
      11'h29D: dout <= 8'b00100100; //  669 :  36 - 0x24
      11'h29E: dout <= 8'b00100100; //  670 :  36 - 0x24
      11'h29F: dout <= 8'b00100100; //  671 :  36 - 0x24
      11'h2A0: dout <= 8'b00100100; //  672 :  36 - 0x24 -- line 0x15
      11'h2A1: dout <= 8'b00100100; //  673 :  36 - 0x24
      11'h2A2: dout <= 8'b00100100; //  674 :  36 - 0x24
      11'h2A3: dout <= 8'b00100100; //  675 :  36 - 0x24
      11'h2A4: dout <= 8'b00110001; //  676 :  49 - 0x31
      11'h2A5: dout <= 8'b00110010; //  677 :  50 - 0x32
      11'h2A6: dout <= 8'b00100100; //  678 :  36 - 0x24
      11'h2A7: dout <= 8'b00100100; //  679 :  36 - 0x24
      11'h2A8: dout <= 8'b00100100; //  680 :  36 - 0x24
      11'h2A9: dout <= 8'b00100100; //  681 :  36 - 0x24
      11'h2AA: dout <= 8'b00100100; //  682 :  36 - 0x24
      11'h2AB: dout <= 8'b00100100; //  683 :  36 - 0x24
      11'h2AC: dout <= 8'b00100100; //  684 :  36 - 0x24
      11'h2AD: dout <= 8'b00100100; //  685 :  36 - 0x24
      11'h2AE: dout <= 8'b00100100; //  686 :  36 - 0x24
      11'h2AF: dout <= 8'b00100100; //  687 :  36 - 0x24
      11'h2B0: dout <= 8'b00100100; //  688 :  36 - 0x24
      11'h2B1: dout <= 8'b00100100; //  689 :  36 - 0x24
      11'h2B2: dout <= 8'b00100100; //  690 :  36 - 0x24
      11'h2B3: dout <= 8'b00100100; //  691 :  36 - 0x24
      11'h2B4: dout <= 8'b00100100; //  692 :  36 - 0x24
      11'h2B5: dout <= 8'b00100100; //  693 :  36 - 0x24
      11'h2B6: dout <= 8'b00100100; //  694 :  36 - 0x24
      11'h2B7: dout <= 8'b00100100; //  695 :  36 - 0x24
      11'h2B8: dout <= 8'b00100100; //  696 :  36 - 0x24
      11'h2B9: dout <= 8'b00100100; //  697 :  36 - 0x24
      11'h2BA: dout <= 8'b00100100; //  698 :  36 - 0x24
      11'h2BB: dout <= 8'b00100100; //  699 :  36 - 0x24
      11'h2BC: dout <= 8'b00100100; //  700 :  36 - 0x24
      11'h2BD: dout <= 8'b00100100; //  701 :  36 - 0x24
      11'h2BE: dout <= 8'b00100100; //  702 :  36 - 0x24
      11'h2BF: dout <= 8'b00100100; //  703 :  36 - 0x24
      11'h2C0: dout <= 8'b00100100; //  704 :  36 - 0x24 -- line 0x16
      11'h2C1: dout <= 8'b00100100; //  705 :  36 - 0x24
      11'h2C2: dout <= 8'b00100100; //  706 :  36 - 0x24
      11'h2C3: dout <= 8'b00110000; //  707 :  48 - 0x30
      11'h2C4: dout <= 8'b00100110; //  708 :  38 - 0x26
      11'h2C5: dout <= 8'b00110100; //  709 :  52 - 0x34
      11'h2C6: dout <= 8'b00110011; //  710 :  51 - 0x33
      11'h2C7: dout <= 8'b00100100; //  711 :  36 - 0x24
      11'h2C8: dout <= 8'b00100100; //  712 :  36 - 0x24
      11'h2C9: dout <= 8'b00100100; //  713 :  36 - 0x24
      11'h2CA: dout <= 8'b00100100; //  714 :  36 - 0x24
      11'h2CB: dout <= 8'b00100100; //  715 :  36 - 0x24
      11'h2CC: dout <= 8'b00100100; //  716 :  36 - 0x24
      11'h2CD: dout <= 8'b00100100; //  717 :  36 - 0x24
      11'h2CE: dout <= 8'b00100100; //  718 :  36 - 0x24
      11'h2CF: dout <= 8'b00100100; //  719 :  36 - 0x24
      11'h2D0: dout <= 8'b00100100; //  720 :  36 - 0x24
      11'h2D1: dout <= 8'b00100100; //  721 :  36 - 0x24
      11'h2D2: dout <= 8'b00100100; //  722 :  36 - 0x24
      11'h2D3: dout <= 8'b00100100; //  723 :  36 - 0x24
      11'h2D4: dout <= 8'b00100100; //  724 :  36 - 0x24
      11'h2D5: dout <= 8'b00100100; //  725 :  36 - 0x24
      11'h2D6: dout <= 8'b00100100; //  726 :  36 - 0x24
      11'h2D7: dout <= 8'b00100100; //  727 :  36 - 0x24
      11'h2D8: dout <= 8'b00100100; //  728 :  36 - 0x24
      11'h2D9: dout <= 8'b00100100; //  729 :  36 - 0x24
      11'h2DA: dout <= 8'b00100100; //  730 :  36 - 0x24
      11'h2DB: dout <= 8'b00100100; //  731 :  36 - 0x24
      11'h2DC: dout <= 8'b00100100; //  732 :  36 - 0x24
      11'h2DD: dout <= 8'b00100100; //  733 :  36 - 0x24
      11'h2DE: dout <= 8'b00100100; //  734 :  36 - 0x24
      11'h2DF: dout <= 8'b00100100; //  735 :  36 - 0x24
      11'h2E0: dout <= 8'b00100100; //  736 :  36 - 0x24 -- line 0x17
      11'h2E1: dout <= 8'b00100100; //  737 :  36 - 0x24
      11'h2E2: dout <= 8'b00110000; //  738 :  48 - 0x30
      11'h2E3: dout <= 8'b00100110; //  739 :  38 - 0x26
      11'h2E4: dout <= 8'b00100110; //  740 :  38 - 0x26
      11'h2E5: dout <= 8'b00100110; //  741 :  38 - 0x26
      11'h2E6: dout <= 8'b00100110; //  742 :  38 - 0x26
      11'h2E7: dout <= 8'b00110011; //  743 :  51 - 0x33
      11'h2E8: dout <= 8'b00100100; //  744 :  36 - 0x24
      11'h2E9: dout <= 8'b00100100; //  745 :  36 - 0x24
      11'h2EA: dout <= 8'b00100100; //  746 :  36 - 0x24
      11'h2EB: dout <= 8'b00100100; //  747 :  36 - 0x24
      11'h2EC: dout <= 8'b00011101; //  748 :  29 - 0x1d
      11'h2ED: dout <= 8'b00011000; //  749 :  24 - 0x18
      11'h2EE: dout <= 8'b00011001; //  750 :  25 - 0x19
      11'h2EF: dout <= 8'b00101000; //  751 :  40 - 0x28
      11'h2F0: dout <= 8'b00100100; //  752 :  36 - 0x24
      11'h2F1: dout <= 8'b00000000; //  753 :   0 - 0x0
      11'h2F2: dout <= 8'b00000000; //  754 :   0 - 0x0
      11'h2F3: dout <= 8'b00000000; //  755 :   0 - 0x0
      11'h2F4: dout <= 8'b00000000; //  756 :   0 - 0x0
      11'h2F5: dout <= 8'b00000000; //  757 :   0 - 0x0
      11'h2F6: dout <= 8'b00000000; //  758 :   0 - 0x0
      11'h2F7: dout <= 8'b00100100; //  759 :  36 - 0x24
      11'h2F8: dout <= 8'b00100100; //  760 :  36 - 0x24
      11'h2F9: dout <= 8'b00100100; //  761 :  36 - 0x24
      11'h2FA: dout <= 8'b00100100; //  762 :  36 - 0x24
      11'h2FB: dout <= 8'b00100100; //  763 :  36 - 0x24
      11'h2FC: dout <= 8'b00100100; //  764 :  36 - 0x24
      11'h2FD: dout <= 8'b00100100; //  765 :  36 - 0x24
      11'h2FE: dout <= 8'b00100100; //  766 :  36 - 0x24
      11'h2FF: dout <= 8'b00100100; //  767 :  36 - 0x24
      11'h300: dout <= 8'b00100100; //  768 :  36 - 0x24 -- line 0x18
      11'h301: dout <= 8'b00110000; //  769 :  48 - 0x30
      11'h302: dout <= 8'b00100110; //  770 :  38 - 0x26
      11'h303: dout <= 8'b00110100; //  771 :  52 - 0x34
      11'h304: dout <= 8'b00100110; //  772 :  38 - 0x26
      11'h305: dout <= 8'b00100110; //  773 :  38 - 0x26
      11'h306: dout <= 8'b00110100; //  774 :  52 - 0x34
      11'h307: dout <= 8'b00100110; //  775 :  38 - 0x26
      11'h308: dout <= 8'b00110011; //  776 :  51 - 0x33
      11'h309: dout <= 8'b00100100; //  777 :  36 - 0x24
      11'h30A: dout <= 8'b00100100; //  778 :  36 - 0x24
      11'h30B: dout <= 8'b00100100; //  779 :  36 - 0x24
      11'h30C: dout <= 8'b00100100; //  780 :  36 - 0x24
      11'h30D: dout <= 8'b00100100; //  781 :  36 - 0x24
      11'h30E: dout <= 8'b00100100; //  782 :  36 - 0x24
      11'h30F: dout <= 8'b00100100; //  783 :  36 - 0x24
      11'h310: dout <= 8'b00100100; //  784 :  36 - 0x24
      11'h311: dout <= 8'b00100100; //  785 :  36 - 0x24
      11'h312: dout <= 8'b00100100; //  786 :  36 - 0x24
      11'h313: dout <= 8'b00100100; //  787 :  36 - 0x24
      11'h314: dout <= 8'b00100100; //  788 :  36 - 0x24
      11'h315: dout <= 8'b00100100; //  789 :  36 - 0x24
      11'h316: dout <= 8'b00100100; //  790 :  36 - 0x24
      11'h317: dout <= 8'b00100100; //  791 :  36 - 0x24
      11'h318: dout <= 8'b00110110; //  792 :  54 - 0x36
      11'h319: dout <= 8'b00110111; //  793 :  55 - 0x37
      11'h31A: dout <= 8'b00110110; //  794 :  54 - 0x36
      11'h31B: dout <= 8'b00110111; //  795 :  55 - 0x37
      11'h31C: dout <= 8'b00110110; //  796 :  54 - 0x36
      11'h31D: dout <= 8'b00110111; //  797 :  55 - 0x37
      11'h31E: dout <= 8'b00100100; //  798 :  36 - 0x24
      11'h31F: dout <= 8'b00100100; //  799 :  36 - 0x24
      11'h320: dout <= 8'b00110000; //  800 :  48 - 0x30 -- line 0x19
      11'h321: dout <= 8'b00100110; //  801 :  38 - 0x26
      11'h322: dout <= 8'b00100110; //  802 :  38 - 0x26
      11'h323: dout <= 8'b00100110; //  803 :  38 - 0x26
      11'h324: dout <= 8'b00100110; //  804 :  38 - 0x26
      11'h325: dout <= 8'b00100110; //  805 :  38 - 0x26
      11'h326: dout <= 8'b00100110; //  806 :  38 - 0x26
      11'h327: dout <= 8'b00100110; //  807 :  38 - 0x26
      11'h328: dout <= 8'b00100110; //  808 :  38 - 0x26
      11'h329: dout <= 8'b00110011; //  809 :  51 - 0x33
      11'h32A: dout <= 8'b00100100; //  810 :  36 - 0x24
      11'h32B: dout <= 8'b00100100; //  811 :  36 - 0x24
      11'h32C: dout <= 8'b00100100; //  812 :  36 - 0x24
      11'h32D: dout <= 8'b00100100; //  813 :  36 - 0x24
      11'h32E: dout <= 8'b00100100; //  814 :  36 - 0x24
      11'h32F: dout <= 8'b00100100; //  815 :  36 - 0x24
      11'h330: dout <= 8'b00100100; //  816 :  36 - 0x24
      11'h331: dout <= 8'b00100100; //  817 :  36 - 0x24
      11'h332: dout <= 8'b00100100; //  818 :  36 - 0x24
      11'h333: dout <= 8'b00100100; //  819 :  36 - 0x24
      11'h334: dout <= 8'b00100100; //  820 :  36 - 0x24
      11'h335: dout <= 8'b00100100; //  821 :  36 - 0x24
      11'h336: dout <= 8'b00100100; //  822 :  36 - 0x24
      11'h337: dout <= 8'b00110101; //  823 :  53 - 0x35
      11'h338: dout <= 8'b00100101; //  824 :  37 - 0x25
      11'h339: dout <= 8'b00100101; //  825 :  37 - 0x25
      11'h33A: dout <= 8'b00100101; //  826 :  37 - 0x25
      11'h33B: dout <= 8'b00100101; //  827 :  37 - 0x25
      11'h33C: dout <= 8'b00100101; //  828 :  37 - 0x25
      11'h33D: dout <= 8'b00100101; //  829 :  37 - 0x25
      11'h33E: dout <= 8'b00111000; //  830 :  56 - 0x38
      11'h33F: dout <= 8'b00100100; //  831 :  36 - 0x24
      11'h340: dout <= 8'b10110100; //  832 : 180 - 0xb4 -- line 0x1a
      11'h341: dout <= 8'b10110101; //  833 : 181 - 0xb5
      11'h342: dout <= 8'b10110100; //  834 : 180 - 0xb4
      11'h343: dout <= 8'b10110101; //  835 : 181 - 0xb5
      11'h344: dout <= 8'b10110100; //  836 : 180 - 0xb4
      11'h345: dout <= 8'b10110101; //  837 : 181 - 0xb5
      11'h346: dout <= 8'b10110100; //  838 : 180 - 0xb4
      11'h347: dout <= 8'b10110101; //  839 : 181 - 0xb5
      11'h348: dout <= 8'b10110100; //  840 : 180 - 0xb4
      11'h349: dout <= 8'b10110101; //  841 : 181 - 0xb5
      11'h34A: dout <= 8'b10110100; //  842 : 180 - 0xb4
      11'h34B: dout <= 8'b10110101; //  843 : 181 - 0xb5
      11'h34C: dout <= 8'b10110100; //  844 : 180 - 0xb4
      11'h34D: dout <= 8'b10110101; //  845 : 181 - 0xb5
      11'h34E: dout <= 8'b10110100; //  846 : 180 - 0xb4
      11'h34F: dout <= 8'b10110101; //  847 : 181 - 0xb5
      11'h350: dout <= 8'b10110100; //  848 : 180 - 0xb4
      11'h351: dout <= 8'b10110101; //  849 : 181 - 0xb5
      11'h352: dout <= 8'b10110100; //  850 : 180 - 0xb4
      11'h353: dout <= 8'b10110101; //  851 : 181 - 0xb5
      11'h354: dout <= 8'b10110100; //  852 : 180 - 0xb4
      11'h355: dout <= 8'b10110101; //  853 : 181 - 0xb5
      11'h356: dout <= 8'b10110100; //  854 : 180 - 0xb4
      11'h357: dout <= 8'b10110101; //  855 : 181 - 0xb5
      11'h358: dout <= 8'b10110100; //  856 : 180 - 0xb4
      11'h359: dout <= 8'b10110101; //  857 : 181 - 0xb5
      11'h35A: dout <= 8'b10110100; //  858 : 180 - 0xb4
      11'h35B: dout <= 8'b10110101; //  859 : 181 - 0xb5
      11'h35C: dout <= 8'b10110100; //  860 : 180 - 0xb4
      11'h35D: dout <= 8'b10110101; //  861 : 181 - 0xb5
      11'h35E: dout <= 8'b10110100; //  862 : 180 - 0xb4
      11'h35F: dout <= 8'b10110101; //  863 : 181 - 0xb5
      11'h360: dout <= 8'b10110110; //  864 : 182 - 0xb6 -- line 0x1b
      11'h361: dout <= 8'b10110111; //  865 : 183 - 0xb7
      11'h362: dout <= 8'b10110110; //  866 : 182 - 0xb6
      11'h363: dout <= 8'b10110111; //  867 : 183 - 0xb7
      11'h364: dout <= 8'b10110110; //  868 : 182 - 0xb6
      11'h365: dout <= 8'b10110111; //  869 : 183 - 0xb7
      11'h366: dout <= 8'b10110110; //  870 : 182 - 0xb6
      11'h367: dout <= 8'b10110111; //  871 : 183 - 0xb7
      11'h368: dout <= 8'b10110110; //  872 : 182 - 0xb6
      11'h369: dout <= 8'b10110111; //  873 : 183 - 0xb7
      11'h36A: dout <= 8'b10110110; //  874 : 182 - 0xb6
      11'h36B: dout <= 8'b10110111; //  875 : 183 - 0xb7
      11'h36C: dout <= 8'b10110110; //  876 : 182 - 0xb6
      11'h36D: dout <= 8'b10110111; //  877 : 183 - 0xb7
      11'h36E: dout <= 8'b10110110; //  878 : 182 - 0xb6
      11'h36F: dout <= 8'b10110111; //  879 : 183 - 0xb7
      11'h370: dout <= 8'b10110110; //  880 : 182 - 0xb6
      11'h371: dout <= 8'b10110111; //  881 : 183 - 0xb7
      11'h372: dout <= 8'b10110110; //  882 : 182 - 0xb6
      11'h373: dout <= 8'b10110111; //  883 : 183 - 0xb7
      11'h374: dout <= 8'b10110110; //  884 : 182 - 0xb6
      11'h375: dout <= 8'b10110111; //  885 : 183 - 0xb7
      11'h376: dout <= 8'b10110110; //  886 : 182 - 0xb6
      11'h377: dout <= 8'b10110111; //  887 : 183 - 0xb7
      11'h378: dout <= 8'b10110110; //  888 : 182 - 0xb6
      11'h379: dout <= 8'b10110111; //  889 : 183 - 0xb7
      11'h37A: dout <= 8'b10110110; //  890 : 182 - 0xb6
      11'h37B: dout <= 8'b10110111; //  891 : 183 - 0xb7
      11'h37C: dout <= 8'b10110110; //  892 : 182 - 0xb6
      11'h37D: dout <= 8'b10110111; //  893 : 183 - 0xb7
      11'h37E: dout <= 8'b10110110; //  894 : 182 - 0xb6
      11'h37F: dout <= 8'b10110111; //  895 : 183 - 0xb7
      11'h380: dout <= 8'b10110100; //  896 : 180 - 0xb4 -- line 0x1c
      11'h381: dout <= 8'b10110101; //  897 : 181 - 0xb5
      11'h382: dout <= 8'b10110100; //  898 : 180 - 0xb4
      11'h383: dout <= 8'b10110101; //  899 : 181 - 0xb5
      11'h384: dout <= 8'b10110100; //  900 : 180 - 0xb4
      11'h385: dout <= 8'b10110101; //  901 : 181 - 0xb5
      11'h386: dout <= 8'b10110100; //  902 : 180 - 0xb4
      11'h387: dout <= 8'b10110101; //  903 : 181 - 0xb5
      11'h388: dout <= 8'b10110100; //  904 : 180 - 0xb4
      11'h389: dout <= 8'b10110101; //  905 : 181 - 0xb5
      11'h38A: dout <= 8'b10110100; //  906 : 180 - 0xb4
      11'h38B: dout <= 8'b10110101; //  907 : 181 - 0xb5
      11'h38C: dout <= 8'b10110100; //  908 : 180 - 0xb4
      11'h38D: dout <= 8'b10110101; //  909 : 181 - 0xb5
      11'h38E: dout <= 8'b10110100; //  910 : 180 - 0xb4
      11'h38F: dout <= 8'b10110101; //  911 : 181 - 0xb5
      11'h390: dout <= 8'b10110100; //  912 : 180 - 0xb4
      11'h391: dout <= 8'b10110101; //  913 : 181 - 0xb5
      11'h392: dout <= 8'b10110100; //  914 : 180 - 0xb4
      11'h393: dout <= 8'b10110101; //  915 : 181 - 0xb5
      11'h394: dout <= 8'b10110100; //  916 : 180 - 0xb4
      11'h395: dout <= 8'b10110101; //  917 : 181 - 0xb5
      11'h396: dout <= 8'b10110100; //  918 : 180 - 0xb4
      11'h397: dout <= 8'b10110101; //  919 : 181 - 0xb5
      11'h398: dout <= 8'b10110100; //  920 : 180 - 0xb4
      11'h399: dout <= 8'b10110101; //  921 : 181 - 0xb5
      11'h39A: dout <= 8'b10110100; //  922 : 180 - 0xb4
      11'h39B: dout <= 8'b10110101; //  923 : 181 - 0xb5
      11'h39C: dout <= 8'b10110100; //  924 : 180 - 0xb4
      11'h39D: dout <= 8'b10110101; //  925 : 181 - 0xb5
      11'h39E: dout <= 8'b10110100; //  926 : 180 - 0xb4
      11'h39F: dout <= 8'b10110101; //  927 : 181 - 0xb5
      11'h3A0: dout <= 8'b10110110; //  928 : 182 - 0xb6 -- line 0x1d
      11'h3A1: dout <= 8'b10110111; //  929 : 183 - 0xb7
      11'h3A2: dout <= 8'b10110110; //  930 : 182 - 0xb6
      11'h3A3: dout <= 8'b10110111; //  931 : 183 - 0xb7
      11'h3A4: dout <= 8'b10110110; //  932 : 182 - 0xb6
      11'h3A5: dout <= 8'b10110111; //  933 : 183 - 0xb7
      11'h3A6: dout <= 8'b10110110; //  934 : 182 - 0xb6
      11'h3A7: dout <= 8'b10110111; //  935 : 183 - 0xb7
      11'h3A8: dout <= 8'b10110110; //  936 : 182 - 0xb6
      11'h3A9: dout <= 8'b10110111; //  937 : 183 - 0xb7
      11'h3AA: dout <= 8'b10110110; //  938 : 182 - 0xb6
      11'h3AB: dout <= 8'b10110111; //  939 : 183 - 0xb7
      11'h3AC: dout <= 8'b10110110; //  940 : 182 - 0xb6
      11'h3AD: dout <= 8'b10110111; //  941 : 183 - 0xb7
      11'h3AE: dout <= 8'b10110110; //  942 : 182 - 0xb6
      11'h3AF: dout <= 8'b10110111; //  943 : 183 - 0xb7
      11'h3B0: dout <= 8'b10110110; //  944 : 182 - 0xb6
      11'h3B1: dout <= 8'b10110111; //  945 : 183 - 0xb7
      11'h3B2: dout <= 8'b10110110; //  946 : 182 - 0xb6
      11'h3B3: dout <= 8'b10110111; //  947 : 183 - 0xb7
      11'h3B4: dout <= 8'b10110110; //  948 : 182 - 0xb6
      11'h3B5: dout <= 8'b10110111; //  949 : 183 - 0xb7
      11'h3B6: dout <= 8'b10110110; //  950 : 182 - 0xb6
      11'h3B7: dout <= 8'b10110111; //  951 : 183 - 0xb7
      11'h3B8: dout <= 8'b10110110; //  952 : 182 - 0xb6
      11'h3B9: dout <= 8'b10110111; //  953 : 183 - 0xb7
      11'h3BA: dout <= 8'b10110110; //  954 : 182 - 0xb6
      11'h3BB: dout <= 8'b10110111; //  955 : 183 - 0xb7
      11'h3BC: dout <= 8'b10110110; //  956 : 182 - 0xb6
      11'h3BD: dout <= 8'b10110111; //  957 : 183 - 0xb7
      11'h3BE: dout <= 8'b10110110; //  958 : 182 - 0xb6
      11'h3BF: dout <= 8'b10110111; //  959 : 183 - 0xb7
        //-- Attribute Table 0----
      11'h3C0: dout <= 8'b10101010; //  960 : 170 - 0xaa
      11'h3C1: dout <= 8'b10101010; //  961 : 170 - 0xaa
      11'h3C2: dout <= 8'b11101010; //  962 : 234 - 0xea
      11'h3C3: dout <= 8'b10101010; //  963 : 170 - 0xaa
      11'h3C4: dout <= 8'b10101010; //  964 : 170 - 0xaa
      11'h3C5: dout <= 8'b10101010; //  965 : 170 - 0xaa
      11'h3C6: dout <= 8'b10101010; //  966 : 170 - 0xaa
      11'h3C7: dout <= 8'b10101010; //  967 : 170 - 0xaa
      11'h3C8: dout <= 8'b00000000; //  968 :   0 - 0x0
      11'h3C9: dout <= 8'b01010101; //  969 :  85 - 0x55
      11'h3CA: dout <= 8'b01010101; //  970 :  85 - 0x55
      11'h3CB: dout <= 8'b01010101; //  971 :  85 - 0x55
      11'h3CC: dout <= 8'b01010101; //  972 :  85 - 0x55
      11'h3CD: dout <= 8'b01010101; //  973 :  85 - 0x55
      11'h3CE: dout <= 8'b01010101; //  974 :  85 - 0x55
      11'h3CF: dout <= 8'b01010101; //  975 :  85 - 0x55
      11'h3D0: dout <= 8'b01010101; //  976 :  85 - 0x55
      11'h3D1: dout <= 8'b01010101; //  977 :  85 - 0x55
      11'h3D2: dout <= 8'b01010101; //  978 :  85 - 0x55
      11'h3D3: dout <= 8'b01010101; //  979 :  85 - 0x55
      11'h3D4: dout <= 8'b01010101; //  980 :  85 - 0x55
      11'h3D5: dout <= 8'b01010101; //  981 :  85 - 0x55
      11'h3D6: dout <= 8'b01010101; //  982 :  85 - 0x55
      11'h3D7: dout <= 8'b01010101; //  983 :  85 - 0x55
      11'h3D8: dout <= 8'b01010101; //  984 :  85 - 0x55
      11'h3D9: dout <= 8'b01010101; //  985 :  85 - 0x55
      11'h3DA: dout <= 8'b01010101; //  986 :  85 - 0x55
      11'h3DB: dout <= 8'b01010101; //  987 :  85 - 0x55
      11'h3DC: dout <= 8'b01010101; //  988 :  85 - 0x55
      11'h3DD: dout <= 8'b01010101; //  989 :  85 - 0x55
      11'h3DE: dout <= 8'b01010101; //  990 :  85 - 0x55
      11'h3DF: dout <= 8'b00000000; //  991 :   0 - 0x0
      11'h3E0: dout <= 8'b00000000; //  992 :   0 - 0x0
      11'h3E1: dout <= 8'b00000000; //  993 :   0 - 0x0
      11'h3E2: dout <= 8'b10011001; //  994 : 153 - 0x99
      11'h3E3: dout <= 8'b10101010; //  995 : 170 - 0xaa
      11'h3E4: dout <= 8'b10101010; //  996 : 170 - 0xaa
      11'h3E5: dout <= 8'b10101010; //  997 : 170 - 0xaa
      11'h3E6: dout <= 8'b00000000; //  998 :   0 - 0x0
      11'h3E7: dout <= 8'b00000000; //  999 :   0 - 0x0
      11'h3E8: dout <= 8'b00000000; // 1000 :   0 - 0x0
      11'h3E9: dout <= 8'b00000000; // 1001 :   0 - 0x0
      11'h3EA: dout <= 8'b10011001; // 1002 : 153 - 0x99
      11'h3EB: dout <= 8'b10101010; // 1003 : 170 - 0xaa
      11'h3EC: dout <= 8'b10101010; // 1004 : 170 - 0xaa
      11'h3ED: dout <= 8'b10101010; // 1005 : 170 - 0xaa
      11'h3EE: dout <= 8'b00000000; // 1006 :   0 - 0x0
      11'h3EF: dout <= 8'b00000000; // 1007 :   0 - 0x0
      11'h3F0: dout <= 8'b01010000; // 1008 :  80 - 0x50
      11'h3F1: dout <= 8'b01010000; // 1009 :  80 - 0x50
      11'h3F2: dout <= 8'b01010000; // 1010 :  80 - 0x50
      11'h3F3: dout <= 8'b01010000; // 1011 :  80 - 0x50
      11'h3F4: dout <= 8'b01010000; // 1012 :  80 - 0x50
      11'h3F5: dout <= 8'b01010000; // 1013 :  80 - 0x50
      11'h3F6: dout <= 8'b01010000; // 1014 :  80 - 0x50
      11'h3F7: dout <= 8'b01010000; // 1015 :  80 - 0x50
      11'h3F8: dout <= 8'b00000101; // 1016 :   5 - 0x5
      11'h3F9: dout <= 8'b00000101; // 1017 :   5 - 0x5
      11'h3FA: dout <= 8'b00000101; // 1018 :   5 - 0x5
      11'h3FB: dout <= 8'b00000101; // 1019 :   5 - 0x5
      11'h3FC: dout <= 8'b00000101; // 1020 :   5 - 0x5
      11'h3FD: dout <= 8'b00000101; // 1021 :   5 - 0x5
      11'h3FE: dout <= 8'b00000101; // 1022 :   5 - 0x5
      11'h3FF: dout <= 8'b00000101; // 1023 :   5 - 0x5
     //----- Name Table 1---------
      11'h400: dout <= 8'b00100100; // 1024 :  36 - 0x24 -- line 0x0
      11'h401: dout <= 8'b00100100; // 1025 :  36 - 0x24
      11'h402: dout <= 8'b00100100; // 1026 :  36 - 0x24
      11'h403: dout <= 8'b00100100; // 1027 :  36 - 0x24
      11'h404: dout <= 8'b00100100; // 1028 :  36 - 0x24
      11'h405: dout <= 8'b00100100; // 1029 :  36 - 0x24
      11'h406: dout <= 8'b00100100; // 1030 :  36 - 0x24
      11'h407: dout <= 8'b00100100; // 1031 :  36 - 0x24
      11'h408: dout <= 8'b00100100; // 1032 :  36 - 0x24
      11'h409: dout <= 8'b00100100; // 1033 :  36 - 0x24
      11'h40A: dout <= 8'b00100100; // 1034 :  36 - 0x24
      11'h40B: dout <= 8'b00100100; // 1035 :  36 - 0x24
      11'h40C: dout <= 8'b00100100; // 1036 :  36 - 0x24
      11'h40D: dout <= 8'b00100100; // 1037 :  36 - 0x24
      11'h40E: dout <= 8'b00100100; // 1038 :  36 - 0x24
      11'h40F: dout <= 8'b00100100; // 1039 :  36 - 0x24
      11'h410: dout <= 8'b00100100; // 1040 :  36 - 0x24
      11'h411: dout <= 8'b00100100; // 1041 :  36 - 0x24
      11'h412: dout <= 8'b00100100; // 1042 :  36 - 0x24
      11'h413: dout <= 8'b00100100; // 1043 :  36 - 0x24
      11'h414: dout <= 8'b00100100; // 1044 :  36 - 0x24
      11'h415: dout <= 8'b00100100; // 1045 :  36 - 0x24
      11'h416: dout <= 8'b00100100; // 1046 :  36 - 0x24
      11'h417: dout <= 8'b00100100; // 1047 :  36 - 0x24
      11'h418: dout <= 8'b00100100; // 1048 :  36 - 0x24
      11'h419: dout <= 8'b00100100; // 1049 :  36 - 0x24
      11'h41A: dout <= 8'b00100100; // 1050 :  36 - 0x24
      11'h41B: dout <= 8'b00100100; // 1051 :  36 - 0x24
      11'h41C: dout <= 8'b00100100; // 1052 :  36 - 0x24
      11'h41D: dout <= 8'b00100100; // 1053 :  36 - 0x24
      11'h41E: dout <= 8'b00100100; // 1054 :  36 - 0x24
      11'h41F: dout <= 8'b00100100; // 1055 :  36 - 0x24
      11'h420: dout <= 8'b00100100; // 1056 :  36 - 0x24 -- line 0x1
      11'h421: dout <= 8'b00100100; // 1057 :  36 - 0x24
      11'h422: dout <= 8'b00100100; // 1058 :  36 - 0x24
      11'h423: dout <= 8'b00100100; // 1059 :  36 - 0x24
      11'h424: dout <= 8'b00100100; // 1060 :  36 - 0x24
      11'h425: dout <= 8'b00100100; // 1061 :  36 - 0x24
      11'h426: dout <= 8'b00100100; // 1062 :  36 - 0x24
      11'h427: dout <= 8'b00100100; // 1063 :  36 - 0x24
      11'h428: dout <= 8'b00100100; // 1064 :  36 - 0x24
      11'h429: dout <= 8'b00100100; // 1065 :  36 - 0x24
      11'h42A: dout <= 8'b00100100; // 1066 :  36 - 0x24
      11'h42B: dout <= 8'b00100100; // 1067 :  36 - 0x24
      11'h42C: dout <= 8'b00100100; // 1068 :  36 - 0x24
      11'h42D: dout <= 8'b00100100; // 1069 :  36 - 0x24
      11'h42E: dout <= 8'b00100100; // 1070 :  36 - 0x24
      11'h42F: dout <= 8'b00100100; // 1071 :  36 - 0x24
      11'h430: dout <= 8'b00100100; // 1072 :  36 - 0x24
      11'h431: dout <= 8'b00100100; // 1073 :  36 - 0x24
      11'h432: dout <= 8'b00100100; // 1074 :  36 - 0x24
      11'h433: dout <= 8'b00100100; // 1075 :  36 - 0x24
      11'h434: dout <= 8'b00100100; // 1076 :  36 - 0x24
      11'h435: dout <= 8'b00100100; // 1077 :  36 - 0x24
      11'h436: dout <= 8'b00100100; // 1078 :  36 - 0x24
      11'h437: dout <= 8'b00100100; // 1079 :  36 - 0x24
      11'h438: dout <= 8'b00100100; // 1080 :  36 - 0x24
      11'h439: dout <= 8'b00100100; // 1081 :  36 - 0x24
      11'h43A: dout <= 8'b00100100; // 1082 :  36 - 0x24
      11'h43B: dout <= 8'b00100100; // 1083 :  36 - 0x24
      11'h43C: dout <= 8'b00100100; // 1084 :  36 - 0x24
      11'h43D: dout <= 8'b00100100; // 1085 :  36 - 0x24
      11'h43E: dout <= 8'b00100100; // 1086 :  36 - 0x24
      11'h43F: dout <= 8'b00100100; // 1087 :  36 - 0x24
      11'h440: dout <= 8'b00100100; // 1088 :  36 - 0x24 -- line 0x2
      11'h441: dout <= 8'b00100100; // 1089 :  36 - 0x24
      11'h442: dout <= 8'b00100100; // 1090 :  36 - 0x24
      11'h443: dout <= 8'b00100100; // 1091 :  36 - 0x24
      11'h444: dout <= 8'b00100100; // 1092 :  36 - 0x24
      11'h445: dout <= 8'b00100100; // 1093 :  36 - 0x24
      11'h446: dout <= 8'b00100100; // 1094 :  36 - 0x24
      11'h447: dout <= 8'b00100100; // 1095 :  36 - 0x24
      11'h448: dout <= 8'b00100100; // 1096 :  36 - 0x24
      11'h449: dout <= 8'b00100100; // 1097 :  36 - 0x24
      11'h44A: dout <= 8'b00100100; // 1098 :  36 - 0x24
      11'h44B: dout <= 8'b00100100; // 1099 :  36 - 0x24
      11'h44C: dout <= 8'b00100100; // 1100 :  36 - 0x24
      11'h44D: dout <= 8'b00100100; // 1101 :  36 - 0x24
      11'h44E: dout <= 8'b00100100; // 1102 :  36 - 0x24
      11'h44F: dout <= 8'b00100100; // 1103 :  36 - 0x24
      11'h450: dout <= 8'b00100100; // 1104 :  36 - 0x24
      11'h451: dout <= 8'b00100100; // 1105 :  36 - 0x24
      11'h452: dout <= 8'b00100100; // 1106 :  36 - 0x24
      11'h453: dout <= 8'b00100100; // 1107 :  36 - 0x24
      11'h454: dout <= 8'b00100100; // 1108 :  36 - 0x24
      11'h455: dout <= 8'b00100100; // 1109 :  36 - 0x24
      11'h456: dout <= 8'b00100100; // 1110 :  36 - 0x24
      11'h457: dout <= 8'b00100100; // 1111 :  36 - 0x24
      11'h458: dout <= 8'b00100100; // 1112 :  36 - 0x24
      11'h459: dout <= 8'b00100100; // 1113 :  36 - 0x24
      11'h45A: dout <= 8'b00100100; // 1114 :  36 - 0x24
      11'h45B: dout <= 8'b00100100; // 1115 :  36 - 0x24
      11'h45C: dout <= 8'b00100100; // 1116 :  36 - 0x24
      11'h45D: dout <= 8'b00100100; // 1117 :  36 - 0x24
      11'h45E: dout <= 8'b00100100; // 1118 :  36 - 0x24
      11'h45F: dout <= 8'b00100100; // 1119 :  36 - 0x24
      11'h460: dout <= 8'b00100100; // 1120 :  36 - 0x24 -- line 0x3
      11'h461: dout <= 8'b00100100; // 1121 :  36 - 0x24
      11'h462: dout <= 8'b00100100; // 1122 :  36 - 0x24
      11'h463: dout <= 8'b00100100; // 1123 :  36 - 0x24
      11'h464: dout <= 8'b00100100; // 1124 :  36 - 0x24
      11'h465: dout <= 8'b00100100; // 1125 :  36 - 0x24
      11'h466: dout <= 8'b00100100; // 1126 :  36 - 0x24
      11'h467: dout <= 8'b00100100; // 1127 :  36 - 0x24
      11'h468: dout <= 8'b00100100; // 1128 :  36 - 0x24
      11'h469: dout <= 8'b00100100; // 1129 :  36 - 0x24
      11'h46A: dout <= 8'b00100100; // 1130 :  36 - 0x24
      11'h46B: dout <= 8'b00100100; // 1131 :  36 - 0x24
      11'h46C: dout <= 8'b00100100; // 1132 :  36 - 0x24
      11'h46D: dout <= 8'b00100100; // 1133 :  36 - 0x24
      11'h46E: dout <= 8'b00100100; // 1134 :  36 - 0x24
      11'h46F: dout <= 8'b00100100; // 1135 :  36 - 0x24
      11'h470: dout <= 8'b00100100; // 1136 :  36 - 0x24
      11'h471: dout <= 8'b00100100; // 1137 :  36 - 0x24
      11'h472: dout <= 8'b00100100; // 1138 :  36 - 0x24
      11'h473: dout <= 8'b00100100; // 1139 :  36 - 0x24
      11'h474: dout <= 8'b00100100; // 1140 :  36 - 0x24
      11'h475: dout <= 8'b00100100; // 1141 :  36 - 0x24
      11'h476: dout <= 8'b00100100; // 1142 :  36 - 0x24
      11'h477: dout <= 8'b00100100; // 1143 :  36 - 0x24
      11'h478: dout <= 8'b00100100; // 1144 :  36 - 0x24
      11'h479: dout <= 8'b00100100; // 1145 :  36 - 0x24
      11'h47A: dout <= 8'b00100100; // 1146 :  36 - 0x24
      11'h47B: dout <= 8'b00100100; // 1147 :  36 - 0x24
      11'h47C: dout <= 8'b00100100; // 1148 :  36 - 0x24
      11'h47D: dout <= 8'b00100100; // 1149 :  36 - 0x24
      11'h47E: dout <= 8'b00100100; // 1150 :  36 - 0x24
      11'h47F: dout <= 8'b00100100; // 1151 :  36 - 0x24
      11'h480: dout <= 8'b00100100; // 1152 :  36 - 0x24 -- line 0x4
      11'h481: dout <= 8'b00100100; // 1153 :  36 - 0x24
      11'h482: dout <= 8'b00100100; // 1154 :  36 - 0x24
      11'h483: dout <= 8'b00100100; // 1155 :  36 - 0x24
      11'h484: dout <= 8'b00100100; // 1156 :  36 - 0x24
      11'h485: dout <= 8'b00100100; // 1157 :  36 - 0x24
      11'h486: dout <= 8'b00100100; // 1158 :  36 - 0x24
      11'h487: dout <= 8'b00100100; // 1159 :  36 - 0x24
      11'h488: dout <= 8'b00110110; // 1160 :  54 - 0x36
      11'h489: dout <= 8'b00110111; // 1161 :  55 - 0x37
      11'h48A: dout <= 8'b00100100; // 1162 :  36 - 0x24
      11'h48B: dout <= 8'b00100100; // 1163 :  36 - 0x24
      11'h48C: dout <= 8'b00100100; // 1164 :  36 - 0x24
      11'h48D: dout <= 8'b00100100; // 1165 :  36 - 0x24
      11'h48E: dout <= 8'b00100100; // 1166 :  36 - 0x24
      11'h48F: dout <= 8'b00100100; // 1167 :  36 - 0x24
      11'h490: dout <= 8'b00100100; // 1168 :  36 - 0x24
      11'h491: dout <= 8'b00100100; // 1169 :  36 - 0x24
      11'h492: dout <= 8'b00100100; // 1170 :  36 - 0x24
      11'h493: dout <= 8'b00100100; // 1171 :  36 - 0x24
      11'h494: dout <= 8'b00100100; // 1172 :  36 - 0x24
      11'h495: dout <= 8'b00100100; // 1173 :  36 - 0x24
      11'h496: dout <= 8'b00100100; // 1174 :  36 - 0x24
      11'h497: dout <= 8'b00100100; // 1175 :  36 - 0x24
      11'h498: dout <= 8'b00100100; // 1176 :  36 - 0x24
      11'h499: dout <= 8'b00100100; // 1177 :  36 - 0x24
      11'h49A: dout <= 8'b00100100; // 1178 :  36 - 0x24
      11'h49B: dout <= 8'b00100100; // 1179 :  36 - 0x24
      11'h49C: dout <= 8'b00100100; // 1180 :  36 - 0x24
      11'h49D: dout <= 8'b00100100; // 1181 :  36 - 0x24
      11'h49E: dout <= 8'b00100100; // 1182 :  36 - 0x24
      11'h49F: dout <= 8'b00100100; // 1183 :  36 - 0x24
      11'h4A0: dout <= 8'b00100100; // 1184 :  36 - 0x24 -- line 0x5
      11'h4A1: dout <= 8'b00100100; // 1185 :  36 - 0x24
      11'h4A2: dout <= 8'b00100100; // 1186 :  36 - 0x24
      11'h4A3: dout <= 8'b00100100; // 1187 :  36 - 0x24
      11'h4A4: dout <= 8'b00100100; // 1188 :  36 - 0x24
      11'h4A5: dout <= 8'b00100100; // 1189 :  36 - 0x24
      11'h4A6: dout <= 8'b00100100; // 1190 :  36 - 0x24
      11'h4A7: dout <= 8'b00110101; // 1191 :  53 - 0x35
      11'h4A8: dout <= 8'b00100101; // 1192 :  37 - 0x25
      11'h4A9: dout <= 8'b00100101; // 1193 :  37 - 0x25
      11'h4AA: dout <= 8'b00111000; // 1194 :  56 - 0x38
      11'h4AB: dout <= 8'b00100100; // 1195 :  36 - 0x24
      11'h4AC: dout <= 8'b00100100; // 1196 :  36 - 0x24
      11'h4AD: dout <= 8'b00100100; // 1197 :  36 - 0x24
      11'h4AE: dout <= 8'b00100100; // 1198 :  36 - 0x24
      11'h4AF: dout <= 8'b00100100; // 1199 :  36 - 0x24
      11'h4B0: dout <= 8'b00100100; // 1200 :  36 - 0x24
      11'h4B1: dout <= 8'b00100100; // 1201 :  36 - 0x24
      11'h4B2: dout <= 8'b00100100; // 1202 :  36 - 0x24
      11'h4B3: dout <= 8'b00100100; // 1203 :  36 - 0x24
      11'h4B4: dout <= 8'b00100100; // 1204 :  36 - 0x24
      11'h4B5: dout <= 8'b00100100; // 1205 :  36 - 0x24
      11'h4B6: dout <= 8'b00100100; // 1206 :  36 - 0x24
      11'h4B7: dout <= 8'b00100100; // 1207 :  36 - 0x24
      11'h4B8: dout <= 8'b00100100; // 1208 :  36 - 0x24
      11'h4B9: dout <= 8'b00100100; // 1209 :  36 - 0x24
      11'h4BA: dout <= 8'b00100100; // 1210 :  36 - 0x24
      11'h4BB: dout <= 8'b00100100; // 1211 :  36 - 0x24
      11'h4BC: dout <= 8'b00100100; // 1212 :  36 - 0x24
      11'h4BD: dout <= 8'b00100100; // 1213 :  36 - 0x24
      11'h4BE: dout <= 8'b00100100; // 1214 :  36 - 0x24
      11'h4BF: dout <= 8'b00100100; // 1215 :  36 - 0x24
      11'h4C0: dout <= 8'b00100100; // 1216 :  36 - 0x24 -- line 0x6
      11'h4C1: dout <= 8'b00100100; // 1217 :  36 - 0x24
      11'h4C2: dout <= 8'b00100100; // 1218 :  36 - 0x24
      11'h4C3: dout <= 8'b00100100; // 1219 :  36 - 0x24
      11'h4C4: dout <= 8'b00100100; // 1220 :  36 - 0x24
      11'h4C5: dout <= 8'b00100100; // 1221 :  36 - 0x24
      11'h4C6: dout <= 8'b00100100; // 1222 :  36 - 0x24
      11'h4C7: dout <= 8'b00111001; // 1223 :  57 - 0x39
      11'h4C8: dout <= 8'b00111010; // 1224 :  58 - 0x3a
      11'h4C9: dout <= 8'b00111011; // 1225 :  59 - 0x3b
      11'h4CA: dout <= 8'b00111100; // 1226 :  60 - 0x3c
      11'h4CB: dout <= 8'b00100100; // 1227 :  36 - 0x24
      11'h4CC: dout <= 8'b00100100; // 1228 :  36 - 0x24
      11'h4CD: dout <= 8'b00100100; // 1229 :  36 - 0x24
      11'h4CE: dout <= 8'b00100100; // 1230 :  36 - 0x24
      11'h4CF: dout <= 8'b00100100; // 1231 :  36 - 0x24
      11'h4D0: dout <= 8'b00100100; // 1232 :  36 - 0x24
      11'h4D1: dout <= 8'b00100100; // 1233 :  36 - 0x24
      11'h4D2: dout <= 8'b00100100; // 1234 :  36 - 0x24
      11'h4D3: dout <= 8'b00100100; // 1235 :  36 - 0x24
      11'h4D4: dout <= 8'b00100100; // 1236 :  36 - 0x24
      11'h4D5: dout <= 8'b00100100; // 1237 :  36 - 0x24
      11'h4D6: dout <= 8'b00100100; // 1238 :  36 - 0x24
      11'h4D7: dout <= 8'b00100100; // 1239 :  36 - 0x24
      11'h4D8: dout <= 8'b00100100; // 1240 :  36 - 0x24
      11'h4D9: dout <= 8'b00100100; // 1241 :  36 - 0x24
      11'h4DA: dout <= 8'b00100100; // 1242 :  36 - 0x24
      11'h4DB: dout <= 8'b00100100; // 1243 :  36 - 0x24
      11'h4DC: dout <= 8'b00100100; // 1244 :  36 - 0x24
      11'h4DD: dout <= 8'b00100100; // 1245 :  36 - 0x24
      11'h4DE: dout <= 8'b00100100; // 1246 :  36 - 0x24
      11'h4DF: dout <= 8'b00100100; // 1247 :  36 - 0x24
      11'h4E0: dout <= 8'b00100100; // 1248 :  36 - 0x24 -- line 0x7
      11'h4E1: dout <= 8'b00100100; // 1249 :  36 - 0x24
      11'h4E2: dout <= 8'b00100100; // 1250 :  36 - 0x24
      11'h4E3: dout <= 8'b00100100; // 1251 :  36 - 0x24
      11'h4E4: dout <= 8'b00100100; // 1252 :  36 - 0x24
      11'h4E5: dout <= 8'b00100100; // 1253 :  36 - 0x24
      11'h4E6: dout <= 8'b00100100; // 1254 :  36 - 0x24
      11'h4E7: dout <= 8'b00100100; // 1255 :  36 - 0x24
      11'h4E8: dout <= 8'b00100100; // 1256 :  36 - 0x24
      11'h4E9: dout <= 8'b00100100; // 1257 :  36 - 0x24
      11'h4EA: dout <= 8'b00100100; // 1258 :  36 - 0x24
      11'h4EB: dout <= 8'b00100100; // 1259 :  36 - 0x24
      11'h4EC: dout <= 8'b00100100; // 1260 :  36 - 0x24
      11'h4ED: dout <= 8'b00100100; // 1261 :  36 - 0x24
      11'h4EE: dout <= 8'b00100100; // 1262 :  36 - 0x24
      11'h4EF: dout <= 8'b00100100; // 1263 :  36 - 0x24
      11'h4F0: dout <= 8'b00100100; // 1264 :  36 - 0x24
      11'h4F1: dout <= 8'b00100100; // 1265 :  36 - 0x24
      11'h4F2: dout <= 8'b00100100; // 1266 :  36 - 0x24
      11'h4F3: dout <= 8'b00100100; // 1267 :  36 - 0x24
      11'h4F4: dout <= 8'b00100100; // 1268 :  36 - 0x24
      11'h4F5: dout <= 8'b00100100; // 1269 :  36 - 0x24
      11'h4F6: dout <= 8'b00100100; // 1270 :  36 - 0x24
      11'h4F7: dout <= 8'b00100100; // 1271 :  36 - 0x24
      11'h4F8: dout <= 8'b00100100; // 1272 :  36 - 0x24
      11'h4F9: dout <= 8'b00100100; // 1273 :  36 - 0x24
      11'h4FA: dout <= 8'b00100100; // 1274 :  36 - 0x24
      11'h4FB: dout <= 8'b00100100; // 1275 :  36 - 0x24
      11'h4FC: dout <= 8'b00100100; // 1276 :  36 - 0x24
      11'h4FD: dout <= 8'b00100100; // 1277 :  36 - 0x24
      11'h4FE: dout <= 8'b00100100; // 1278 :  36 - 0x24
      11'h4FF: dout <= 8'b00100100; // 1279 :  36 - 0x24
      11'h500: dout <= 8'b00100100; // 1280 :  36 - 0x24 -- line 0x8
      11'h501: dout <= 8'b00100100; // 1281 :  36 - 0x24
      11'h502: dout <= 8'b00100100; // 1282 :  36 - 0x24
      11'h503: dout <= 8'b00100100; // 1283 :  36 - 0x24
      11'h504: dout <= 8'b00100100; // 1284 :  36 - 0x24
      11'h505: dout <= 8'b00100100; // 1285 :  36 - 0x24
      11'h506: dout <= 8'b00100100; // 1286 :  36 - 0x24
      11'h507: dout <= 8'b00100100; // 1287 :  36 - 0x24
      11'h508: dout <= 8'b00100100; // 1288 :  36 - 0x24
      11'h509: dout <= 8'b00100100; // 1289 :  36 - 0x24
      11'h50A: dout <= 8'b00100100; // 1290 :  36 - 0x24
      11'h50B: dout <= 8'b00100100; // 1291 :  36 - 0x24
      11'h50C: dout <= 8'b00100100; // 1292 :  36 - 0x24
      11'h50D: dout <= 8'b00100100; // 1293 :  36 - 0x24
      11'h50E: dout <= 8'b00100100; // 1294 :  36 - 0x24
      11'h50F: dout <= 8'b00100100; // 1295 :  36 - 0x24
      11'h510: dout <= 8'b00100100; // 1296 :  36 - 0x24
      11'h511: dout <= 8'b00100100; // 1297 :  36 - 0x24
      11'h512: dout <= 8'b00100100; // 1298 :  36 - 0x24
      11'h513: dout <= 8'b00100100; // 1299 :  36 - 0x24
      11'h514: dout <= 8'b00100100; // 1300 :  36 - 0x24
      11'h515: dout <= 8'b00100100; // 1301 :  36 - 0x24
      11'h516: dout <= 8'b00100100; // 1302 :  36 - 0x24
      11'h517: dout <= 8'b00100100; // 1303 :  36 - 0x24
      11'h518: dout <= 8'b00100100; // 1304 :  36 - 0x24
      11'h519: dout <= 8'b00100100; // 1305 :  36 - 0x24
      11'h51A: dout <= 8'b00100100; // 1306 :  36 - 0x24
      11'h51B: dout <= 8'b00100100; // 1307 :  36 - 0x24
      11'h51C: dout <= 8'b00100100; // 1308 :  36 - 0x24
      11'h51D: dout <= 8'b00100100; // 1309 :  36 - 0x24
      11'h51E: dout <= 8'b00100100; // 1310 :  36 - 0x24
      11'h51F: dout <= 8'b00100100; // 1311 :  36 - 0x24
      11'h520: dout <= 8'b00100100; // 1312 :  36 - 0x24 -- line 0x9
      11'h521: dout <= 8'b00100100; // 1313 :  36 - 0x24
      11'h522: dout <= 8'b00100100; // 1314 :  36 - 0x24
      11'h523: dout <= 8'b00100100; // 1315 :  36 - 0x24
      11'h524: dout <= 8'b00100100; // 1316 :  36 - 0x24
      11'h525: dout <= 8'b00100100; // 1317 :  36 - 0x24
      11'h526: dout <= 8'b00100100; // 1318 :  36 - 0x24
      11'h527: dout <= 8'b00100100; // 1319 :  36 - 0x24
      11'h528: dout <= 8'b00100100; // 1320 :  36 - 0x24
      11'h529: dout <= 8'b00100100; // 1321 :  36 - 0x24
      11'h52A: dout <= 8'b00100100; // 1322 :  36 - 0x24
      11'h52B: dout <= 8'b00100100; // 1323 :  36 - 0x24
      11'h52C: dout <= 8'b00100100; // 1324 :  36 - 0x24
      11'h52D: dout <= 8'b00100100; // 1325 :  36 - 0x24
      11'h52E: dout <= 8'b00100100; // 1326 :  36 - 0x24
      11'h52F: dout <= 8'b00100100; // 1327 :  36 - 0x24
      11'h530: dout <= 8'b00100100; // 1328 :  36 - 0x24
      11'h531: dout <= 8'b00100100; // 1329 :  36 - 0x24
      11'h532: dout <= 8'b00100100; // 1330 :  36 - 0x24
      11'h533: dout <= 8'b00100100; // 1331 :  36 - 0x24
      11'h534: dout <= 8'b00100100; // 1332 :  36 - 0x24
      11'h535: dout <= 8'b00100100; // 1333 :  36 - 0x24
      11'h536: dout <= 8'b00100100; // 1334 :  36 - 0x24
      11'h537: dout <= 8'b00100100; // 1335 :  36 - 0x24
      11'h538: dout <= 8'b00100100; // 1336 :  36 - 0x24
      11'h539: dout <= 8'b00100100; // 1337 :  36 - 0x24
      11'h53A: dout <= 8'b00100100; // 1338 :  36 - 0x24
      11'h53B: dout <= 8'b00100100; // 1339 :  36 - 0x24
      11'h53C: dout <= 8'b00100100; // 1340 :  36 - 0x24
      11'h53D: dout <= 8'b00100100; // 1341 :  36 - 0x24
      11'h53E: dout <= 8'b00100100; // 1342 :  36 - 0x24
      11'h53F: dout <= 8'b00100100; // 1343 :  36 - 0x24
      11'h540: dout <= 8'b00100100; // 1344 :  36 - 0x24 -- line 0xa
      11'h541: dout <= 8'b00100100; // 1345 :  36 - 0x24
      11'h542: dout <= 8'b00100100; // 1346 :  36 - 0x24
      11'h543: dout <= 8'b00100100; // 1347 :  36 - 0x24
      11'h544: dout <= 8'b00100100; // 1348 :  36 - 0x24
      11'h545: dout <= 8'b00100100; // 1349 :  36 - 0x24
      11'h546: dout <= 8'b00100100; // 1350 :  36 - 0x24
      11'h547: dout <= 8'b00100100; // 1351 :  36 - 0x24
      11'h548: dout <= 8'b00100100; // 1352 :  36 - 0x24
      11'h549: dout <= 8'b00100100; // 1353 :  36 - 0x24
      11'h54A: dout <= 8'b00100100; // 1354 :  36 - 0x24
      11'h54B: dout <= 8'b00100100; // 1355 :  36 - 0x24
      11'h54C: dout <= 8'b01010011; // 1356 :  83 - 0x53
      11'h54D: dout <= 8'b01010100; // 1357 :  84 - 0x54
      11'h54E: dout <= 8'b00100100; // 1358 :  36 - 0x24
      11'h54F: dout <= 8'b00100100; // 1359 :  36 - 0x24
      11'h550: dout <= 8'b00100100; // 1360 :  36 - 0x24
      11'h551: dout <= 8'b00100100; // 1361 :  36 - 0x24
      11'h552: dout <= 8'b00100100; // 1362 :  36 - 0x24
      11'h553: dout <= 8'b00100100; // 1363 :  36 - 0x24
      11'h554: dout <= 8'b00100100; // 1364 :  36 - 0x24
      11'h555: dout <= 8'b00100100; // 1365 :  36 - 0x24
      11'h556: dout <= 8'b00100100; // 1366 :  36 - 0x24
      11'h557: dout <= 8'b00100100; // 1367 :  36 - 0x24
      11'h558: dout <= 8'b00100100; // 1368 :  36 - 0x24
      11'h559: dout <= 8'b00100100; // 1369 :  36 - 0x24
      11'h55A: dout <= 8'b00100100; // 1370 :  36 - 0x24
      11'h55B: dout <= 8'b00100100; // 1371 :  36 - 0x24
      11'h55C: dout <= 8'b00100100; // 1372 :  36 - 0x24
      11'h55D: dout <= 8'b00100100; // 1373 :  36 - 0x24
      11'h55E: dout <= 8'b00100100; // 1374 :  36 - 0x24
      11'h55F: dout <= 8'b00100100; // 1375 :  36 - 0x24
      11'h560: dout <= 8'b00100100; // 1376 :  36 - 0x24 -- line 0xb
      11'h561: dout <= 8'b00100100; // 1377 :  36 - 0x24
      11'h562: dout <= 8'b00100100; // 1378 :  36 - 0x24
      11'h563: dout <= 8'b00100100; // 1379 :  36 - 0x24
      11'h564: dout <= 8'b00100100; // 1380 :  36 - 0x24
      11'h565: dout <= 8'b00100100; // 1381 :  36 - 0x24
      11'h566: dout <= 8'b00100100; // 1382 :  36 - 0x24
      11'h567: dout <= 8'b00100100; // 1383 :  36 - 0x24
      11'h568: dout <= 8'b00100100; // 1384 :  36 - 0x24
      11'h569: dout <= 8'b00100100; // 1385 :  36 - 0x24
      11'h56A: dout <= 8'b00100100; // 1386 :  36 - 0x24
      11'h56B: dout <= 8'b00100100; // 1387 :  36 - 0x24
      11'h56C: dout <= 8'b01010101; // 1388 :  85 - 0x55
      11'h56D: dout <= 8'b01010110; // 1389 :  86 - 0x56
      11'h56E: dout <= 8'b00100100; // 1390 :  36 - 0x24
      11'h56F: dout <= 8'b00100100; // 1391 :  36 - 0x24
      11'h570: dout <= 8'b00100100; // 1392 :  36 - 0x24
      11'h571: dout <= 8'b00100100; // 1393 :  36 - 0x24
      11'h572: dout <= 8'b00100100; // 1394 :  36 - 0x24
      11'h573: dout <= 8'b00100100; // 1395 :  36 - 0x24
      11'h574: dout <= 8'b00100100; // 1396 :  36 - 0x24
      11'h575: dout <= 8'b00100100; // 1397 :  36 - 0x24
      11'h576: dout <= 8'b00100100; // 1398 :  36 - 0x24
      11'h577: dout <= 8'b00100100; // 1399 :  36 - 0x24
      11'h578: dout <= 8'b00100100; // 1400 :  36 - 0x24
      11'h579: dout <= 8'b00100100; // 1401 :  36 - 0x24
      11'h57A: dout <= 8'b00100100; // 1402 :  36 - 0x24
      11'h57B: dout <= 8'b00100100; // 1403 :  36 - 0x24
      11'h57C: dout <= 8'b00100100; // 1404 :  36 - 0x24
      11'h57D: dout <= 8'b00100100; // 1405 :  36 - 0x24
      11'h57E: dout <= 8'b00100100; // 1406 :  36 - 0x24
      11'h57F: dout <= 8'b00100100; // 1407 :  36 - 0x24
      11'h580: dout <= 8'b00100100; // 1408 :  36 - 0x24 -- line 0xc
      11'h581: dout <= 8'b00100100; // 1409 :  36 - 0x24
      11'h582: dout <= 8'b00100100; // 1410 :  36 - 0x24
      11'h583: dout <= 8'b00100100; // 1411 :  36 - 0x24
      11'h584: dout <= 8'b00100100; // 1412 :  36 - 0x24
      11'h585: dout <= 8'b00100100; // 1413 :  36 - 0x24
      11'h586: dout <= 8'b00100100; // 1414 :  36 - 0x24
      11'h587: dout <= 8'b00100100; // 1415 :  36 - 0x24
      11'h588: dout <= 8'b00100100; // 1416 :  36 - 0x24
      11'h589: dout <= 8'b00100100; // 1417 :  36 - 0x24
      11'h58A: dout <= 8'b00100100; // 1418 :  36 - 0x24
      11'h58B: dout <= 8'b00100100; // 1419 :  36 - 0x24
      11'h58C: dout <= 8'b00100100; // 1420 :  36 - 0x24
      11'h58D: dout <= 8'b00100100; // 1421 :  36 - 0x24
      11'h58E: dout <= 8'b00100100; // 1422 :  36 - 0x24
      11'h58F: dout <= 8'b00100100; // 1423 :  36 - 0x24
      11'h590: dout <= 8'b00100100; // 1424 :  36 - 0x24
      11'h591: dout <= 8'b00100100; // 1425 :  36 - 0x24
      11'h592: dout <= 8'b00100100; // 1426 :  36 - 0x24
      11'h593: dout <= 8'b00100100; // 1427 :  36 - 0x24
      11'h594: dout <= 8'b00100100; // 1428 :  36 - 0x24
      11'h595: dout <= 8'b00100100; // 1429 :  36 - 0x24
      11'h596: dout <= 8'b00100100; // 1430 :  36 - 0x24
      11'h597: dout <= 8'b00100100; // 1431 :  36 - 0x24
      11'h598: dout <= 8'b00100100; // 1432 :  36 - 0x24
      11'h599: dout <= 8'b00100100; // 1433 :  36 - 0x24
      11'h59A: dout <= 8'b00100100; // 1434 :  36 - 0x24
      11'h59B: dout <= 8'b00100100; // 1435 :  36 - 0x24
      11'h59C: dout <= 8'b00100100; // 1436 :  36 - 0x24
      11'h59D: dout <= 8'b00100100; // 1437 :  36 - 0x24
      11'h59E: dout <= 8'b00100100; // 1438 :  36 - 0x24
      11'h59F: dout <= 8'b00100100; // 1439 :  36 - 0x24
      11'h5A0: dout <= 8'b00100100; // 1440 :  36 - 0x24 -- line 0xd
      11'h5A1: dout <= 8'b00100100; // 1441 :  36 - 0x24
      11'h5A2: dout <= 8'b00100100; // 1442 :  36 - 0x24
      11'h5A3: dout <= 8'b00100100; // 1443 :  36 - 0x24
      11'h5A4: dout <= 8'b00100100; // 1444 :  36 - 0x24
      11'h5A5: dout <= 8'b00100100; // 1445 :  36 - 0x24
      11'h5A6: dout <= 8'b00100100; // 1446 :  36 - 0x24
      11'h5A7: dout <= 8'b00100100; // 1447 :  36 - 0x24
      11'h5A8: dout <= 8'b00100100; // 1448 :  36 - 0x24
      11'h5A9: dout <= 8'b00100100; // 1449 :  36 - 0x24
      11'h5AA: dout <= 8'b00100100; // 1450 :  36 - 0x24
      11'h5AB: dout <= 8'b00100100; // 1451 :  36 - 0x24
      11'h5AC: dout <= 8'b00100100; // 1452 :  36 - 0x24
      11'h5AD: dout <= 8'b00100100; // 1453 :  36 - 0x24
      11'h5AE: dout <= 8'b00100100; // 1454 :  36 - 0x24
      11'h5AF: dout <= 8'b00100100; // 1455 :  36 - 0x24
      11'h5B0: dout <= 8'b00100100; // 1456 :  36 - 0x24
      11'h5B1: dout <= 8'b00100100; // 1457 :  36 - 0x24
      11'h5B2: dout <= 8'b00100100; // 1458 :  36 - 0x24
      11'h5B3: dout <= 8'b00100100; // 1459 :  36 - 0x24
      11'h5B4: dout <= 8'b00100100; // 1460 :  36 - 0x24
      11'h5B5: dout <= 8'b00100100; // 1461 :  36 - 0x24
      11'h5B6: dout <= 8'b00100100; // 1462 :  36 - 0x24
      11'h5B7: dout <= 8'b00100100; // 1463 :  36 - 0x24
      11'h5B8: dout <= 8'b00100100; // 1464 :  36 - 0x24
      11'h5B9: dout <= 8'b00100100; // 1465 :  36 - 0x24
      11'h5BA: dout <= 8'b00100100; // 1466 :  36 - 0x24
      11'h5BB: dout <= 8'b00100100; // 1467 :  36 - 0x24
      11'h5BC: dout <= 8'b00100100; // 1468 :  36 - 0x24
      11'h5BD: dout <= 8'b00100100; // 1469 :  36 - 0x24
      11'h5BE: dout <= 8'b00100100; // 1470 :  36 - 0x24
      11'h5BF: dout <= 8'b00100100; // 1471 :  36 - 0x24
      11'h5C0: dout <= 8'b00100100; // 1472 :  36 - 0x24 -- line 0xe
      11'h5C1: dout <= 8'b00100100; // 1473 :  36 - 0x24
      11'h5C2: dout <= 8'b00100100; // 1474 :  36 - 0x24
      11'h5C3: dout <= 8'b00100100; // 1475 :  36 - 0x24
      11'h5C4: dout <= 8'b00100100; // 1476 :  36 - 0x24
      11'h5C5: dout <= 8'b00100100; // 1477 :  36 - 0x24
      11'h5C6: dout <= 8'b00100100; // 1478 :  36 - 0x24
      11'h5C7: dout <= 8'b00100100; // 1479 :  36 - 0x24
      11'h5C8: dout <= 8'b00100100; // 1480 :  36 - 0x24
      11'h5C9: dout <= 8'b00100100; // 1481 :  36 - 0x24
      11'h5CA: dout <= 8'b00100100; // 1482 :  36 - 0x24
      11'h5CB: dout <= 8'b00100100; // 1483 :  36 - 0x24
      11'h5CC: dout <= 8'b00100100; // 1484 :  36 - 0x24
      11'h5CD: dout <= 8'b00100100; // 1485 :  36 - 0x24
      11'h5CE: dout <= 8'b00100100; // 1486 :  36 - 0x24
      11'h5CF: dout <= 8'b00100100; // 1487 :  36 - 0x24
      11'h5D0: dout <= 8'b00100100; // 1488 :  36 - 0x24
      11'h5D1: dout <= 8'b00100100; // 1489 :  36 - 0x24
      11'h5D2: dout <= 8'b00100100; // 1490 :  36 - 0x24
      11'h5D3: dout <= 8'b00100100; // 1491 :  36 - 0x24
      11'h5D4: dout <= 8'b00100100; // 1492 :  36 - 0x24
      11'h5D5: dout <= 8'b00100100; // 1493 :  36 - 0x24
      11'h5D6: dout <= 8'b00100100; // 1494 :  36 - 0x24
      11'h5D7: dout <= 8'b00100100; // 1495 :  36 - 0x24
      11'h5D8: dout <= 8'b00100100; // 1496 :  36 - 0x24
      11'h5D9: dout <= 8'b00100100; // 1497 :  36 - 0x24
      11'h5DA: dout <= 8'b00100100; // 1498 :  36 - 0x24
      11'h5DB: dout <= 8'b00100100; // 1499 :  36 - 0x24
      11'h5DC: dout <= 8'b00100100; // 1500 :  36 - 0x24
      11'h5DD: dout <= 8'b00100100; // 1501 :  36 - 0x24
      11'h5DE: dout <= 8'b00100100; // 1502 :  36 - 0x24
      11'h5DF: dout <= 8'b00100100; // 1503 :  36 - 0x24
      11'h5E0: dout <= 8'b00100100; // 1504 :  36 - 0x24 -- line 0xf
      11'h5E1: dout <= 8'b00100100; // 1505 :  36 - 0x24
      11'h5E2: dout <= 8'b00100100; // 1506 :  36 - 0x24
      11'h5E3: dout <= 8'b00100100; // 1507 :  36 - 0x24
      11'h5E4: dout <= 8'b00100100; // 1508 :  36 - 0x24
      11'h5E5: dout <= 8'b00100100; // 1509 :  36 - 0x24
      11'h5E6: dout <= 8'b00100100; // 1510 :  36 - 0x24
      11'h5E7: dout <= 8'b00100100; // 1511 :  36 - 0x24
      11'h5E8: dout <= 8'b00100100; // 1512 :  36 - 0x24
      11'h5E9: dout <= 8'b00100100; // 1513 :  36 - 0x24
      11'h5EA: dout <= 8'b00100100; // 1514 :  36 - 0x24
      11'h5EB: dout <= 8'b00100100; // 1515 :  36 - 0x24
      11'h5EC: dout <= 8'b00100100; // 1516 :  36 - 0x24
      11'h5ED: dout <= 8'b00100100; // 1517 :  36 - 0x24
      11'h5EE: dout <= 8'b00100100; // 1518 :  36 - 0x24
      11'h5EF: dout <= 8'b00100100; // 1519 :  36 - 0x24
      11'h5F0: dout <= 8'b00100100; // 1520 :  36 - 0x24
      11'h5F1: dout <= 8'b00100100; // 1521 :  36 - 0x24
      11'h5F2: dout <= 8'b00100100; // 1522 :  36 - 0x24
      11'h5F3: dout <= 8'b00100100; // 1523 :  36 - 0x24
      11'h5F4: dout <= 8'b00100100; // 1524 :  36 - 0x24
      11'h5F5: dout <= 8'b00100100; // 1525 :  36 - 0x24
      11'h5F6: dout <= 8'b00100100; // 1526 :  36 - 0x24
      11'h5F7: dout <= 8'b00100100; // 1527 :  36 - 0x24
      11'h5F8: dout <= 8'b00100100; // 1528 :  36 - 0x24
      11'h5F9: dout <= 8'b00100100; // 1529 :  36 - 0x24
      11'h5FA: dout <= 8'b00100100; // 1530 :  36 - 0x24
      11'h5FB: dout <= 8'b00100100; // 1531 :  36 - 0x24
      11'h5FC: dout <= 8'b00100100; // 1532 :  36 - 0x24
      11'h5FD: dout <= 8'b00100100; // 1533 :  36 - 0x24
      11'h5FE: dout <= 8'b00100100; // 1534 :  36 - 0x24
      11'h5FF: dout <= 8'b00100100; // 1535 :  36 - 0x24
      11'h600: dout <= 8'b00100100; // 1536 :  36 - 0x24 -- line 0x10
      11'h601: dout <= 8'b00100100; // 1537 :  36 - 0x24
      11'h602: dout <= 8'b00100100; // 1538 :  36 - 0x24
      11'h603: dout <= 8'b00100100; // 1539 :  36 - 0x24
      11'h604: dout <= 8'b00100100; // 1540 :  36 - 0x24
      11'h605: dout <= 8'b00100100; // 1541 :  36 - 0x24
      11'h606: dout <= 8'b00100100; // 1542 :  36 - 0x24
      11'h607: dout <= 8'b00100100; // 1543 :  36 - 0x24
      11'h608: dout <= 8'b00100100; // 1544 :  36 - 0x24
      11'h609: dout <= 8'b00100100; // 1545 :  36 - 0x24
      11'h60A: dout <= 8'b00100100; // 1546 :  36 - 0x24
      11'h60B: dout <= 8'b00100100; // 1547 :  36 - 0x24
      11'h60C: dout <= 8'b00100100; // 1548 :  36 - 0x24
      11'h60D: dout <= 8'b00100100; // 1549 :  36 - 0x24
      11'h60E: dout <= 8'b00100100; // 1550 :  36 - 0x24
      11'h60F: dout <= 8'b00100100; // 1551 :  36 - 0x24
      11'h610: dout <= 8'b00100100; // 1552 :  36 - 0x24
      11'h611: dout <= 8'b00100100; // 1553 :  36 - 0x24
      11'h612: dout <= 8'b00100100; // 1554 :  36 - 0x24
      11'h613: dout <= 8'b00100100; // 1555 :  36 - 0x24
      11'h614: dout <= 8'b00100100; // 1556 :  36 - 0x24
      11'h615: dout <= 8'b00100100; // 1557 :  36 - 0x24
      11'h616: dout <= 8'b00100100; // 1558 :  36 - 0x24
      11'h617: dout <= 8'b00100100; // 1559 :  36 - 0x24
      11'h618: dout <= 8'b00100100; // 1560 :  36 - 0x24
      11'h619: dout <= 8'b00100100; // 1561 :  36 - 0x24
      11'h61A: dout <= 8'b00100100; // 1562 :  36 - 0x24
      11'h61B: dout <= 8'b00100100; // 1563 :  36 - 0x24
      11'h61C: dout <= 8'b00100100; // 1564 :  36 - 0x24
      11'h61D: dout <= 8'b00100100; // 1565 :  36 - 0x24
      11'h61E: dout <= 8'b00100100; // 1566 :  36 - 0x24
      11'h61F: dout <= 8'b00100100; // 1567 :  36 - 0x24
      11'h620: dout <= 8'b00100100; // 1568 :  36 - 0x24 -- line 0x11
      11'h621: dout <= 8'b00100100; // 1569 :  36 - 0x24
      11'h622: dout <= 8'b00100100; // 1570 :  36 - 0x24
      11'h623: dout <= 8'b00100100; // 1571 :  36 - 0x24
      11'h624: dout <= 8'b00100100; // 1572 :  36 - 0x24
      11'h625: dout <= 8'b00100100; // 1573 :  36 - 0x24
      11'h626: dout <= 8'b00100100; // 1574 :  36 - 0x24
      11'h627: dout <= 8'b00100100; // 1575 :  36 - 0x24
      11'h628: dout <= 8'b00100100; // 1576 :  36 - 0x24
      11'h629: dout <= 8'b00100100; // 1577 :  36 - 0x24
      11'h62A: dout <= 8'b00100100; // 1578 :  36 - 0x24
      11'h62B: dout <= 8'b00100100; // 1579 :  36 - 0x24
      11'h62C: dout <= 8'b00100100; // 1580 :  36 - 0x24
      11'h62D: dout <= 8'b00100100; // 1581 :  36 - 0x24
      11'h62E: dout <= 8'b00100100; // 1582 :  36 - 0x24
      11'h62F: dout <= 8'b00100100; // 1583 :  36 - 0x24
      11'h630: dout <= 8'b00100100; // 1584 :  36 - 0x24
      11'h631: dout <= 8'b00100100; // 1585 :  36 - 0x24
      11'h632: dout <= 8'b00100100; // 1586 :  36 - 0x24
      11'h633: dout <= 8'b00100100; // 1587 :  36 - 0x24
      11'h634: dout <= 8'b00100100; // 1588 :  36 - 0x24
      11'h635: dout <= 8'b00100100; // 1589 :  36 - 0x24
      11'h636: dout <= 8'b00100100; // 1590 :  36 - 0x24
      11'h637: dout <= 8'b00100100; // 1591 :  36 - 0x24
      11'h638: dout <= 8'b00100100; // 1592 :  36 - 0x24
      11'h639: dout <= 8'b00100100; // 1593 :  36 - 0x24
      11'h63A: dout <= 8'b00100100; // 1594 :  36 - 0x24
      11'h63B: dout <= 8'b00100100; // 1595 :  36 - 0x24
      11'h63C: dout <= 8'b00100100; // 1596 :  36 - 0x24
      11'h63D: dout <= 8'b00100100; // 1597 :  36 - 0x24
      11'h63E: dout <= 8'b00100100; // 1598 :  36 - 0x24
      11'h63F: dout <= 8'b00100100; // 1599 :  36 - 0x24
      11'h640: dout <= 8'b01010011; // 1600 :  83 - 0x53 -- line 0x12
      11'h641: dout <= 8'b01010100; // 1601 :  84 - 0x54
      11'h642: dout <= 8'b00100100; // 1602 :  36 - 0x24
      11'h643: dout <= 8'b00100100; // 1603 :  36 - 0x24
      11'h644: dout <= 8'b00100100; // 1604 :  36 - 0x24
      11'h645: dout <= 8'b00100100; // 1605 :  36 - 0x24
      11'h646: dout <= 8'b00100100; // 1606 :  36 - 0x24
      11'h647: dout <= 8'b00100100; // 1607 :  36 - 0x24
      11'h648: dout <= 8'b01000101; // 1608 :  69 - 0x45
      11'h649: dout <= 8'b01000101; // 1609 :  69 - 0x45
      11'h64A: dout <= 8'b01010011; // 1610 :  83 - 0x53
      11'h64B: dout <= 8'b01010100; // 1611 :  84 - 0x54
      11'h64C: dout <= 8'b01000101; // 1612 :  69 - 0x45
      11'h64D: dout <= 8'b01000101; // 1613 :  69 - 0x45
      11'h64E: dout <= 8'b01010011; // 1614 :  83 - 0x53
      11'h64F: dout <= 8'b01010100; // 1615 :  84 - 0x54
      11'h650: dout <= 8'b00100100; // 1616 :  36 - 0x24
      11'h651: dout <= 8'b00100100; // 1617 :  36 - 0x24
      11'h652: dout <= 8'b00100100; // 1618 :  36 - 0x24
      11'h653: dout <= 8'b00100100; // 1619 :  36 - 0x24
      11'h654: dout <= 8'b00100100; // 1620 :  36 - 0x24
      11'h655: dout <= 8'b00100100; // 1621 :  36 - 0x24
      11'h656: dout <= 8'b00100100; // 1622 :  36 - 0x24
      11'h657: dout <= 8'b00100100; // 1623 :  36 - 0x24
      11'h658: dout <= 8'b00100100; // 1624 :  36 - 0x24
      11'h659: dout <= 8'b00100100; // 1625 :  36 - 0x24
      11'h65A: dout <= 8'b00100100; // 1626 :  36 - 0x24
      11'h65B: dout <= 8'b00100100; // 1627 :  36 - 0x24
      11'h65C: dout <= 8'b00100100; // 1628 :  36 - 0x24
      11'h65D: dout <= 8'b00100100; // 1629 :  36 - 0x24
      11'h65E: dout <= 8'b00100100; // 1630 :  36 - 0x24
      11'h65F: dout <= 8'b00100100; // 1631 :  36 - 0x24
      11'h660: dout <= 8'b01010101; // 1632 :  85 - 0x55 -- line 0x13
      11'h661: dout <= 8'b01010110; // 1633 :  86 - 0x56
      11'h662: dout <= 8'b00100100; // 1634 :  36 - 0x24
      11'h663: dout <= 8'b00100100; // 1635 :  36 - 0x24
      11'h664: dout <= 8'b00100100; // 1636 :  36 - 0x24
      11'h665: dout <= 8'b00100100; // 1637 :  36 - 0x24
      11'h666: dout <= 8'b00100100; // 1638 :  36 - 0x24
      11'h667: dout <= 8'b00100100; // 1639 :  36 - 0x24
      11'h668: dout <= 8'b01000111; // 1640 :  71 - 0x47
      11'h669: dout <= 8'b01000111; // 1641 :  71 - 0x47
      11'h66A: dout <= 8'b01010101; // 1642 :  85 - 0x55
      11'h66B: dout <= 8'b01010110; // 1643 :  86 - 0x56
      11'h66C: dout <= 8'b01000111; // 1644 :  71 - 0x47
      11'h66D: dout <= 8'b01000111; // 1645 :  71 - 0x47
      11'h66E: dout <= 8'b01010101; // 1646 :  85 - 0x55
      11'h66F: dout <= 8'b01010110; // 1647 :  86 - 0x56
      11'h670: dout <= 8'b00100100; // 1648 :  36 - 0x24
      11'h671: dout <= 8'b00100100; // 1649 :  36 - 0x24
      11'h672: dout <= 8'b00100100; // 1650 :  36 - 0x24
      11'h673: dout <= 8'b00100100; // 1651 :  36 - 0x24
      11'h674: dout <= 8'b00100100; // 1652 :  36 - 0x24
      11'h675: dout <= 8'b00100100; // 1653 :  36 - 0x24
      11'h676: dout <= 8'b00100100; // 1654 :  36 - 0x24
      11'h677: dout <= 8'b00100100; // 1655 :  36 - 0x24
      11'h678: dout <= 8'b00100100; // 1656 :  36 - 0x24
      11'h679: dout <= 8'b00100100; // 1657 :  36 - 0x24
      11'h67A: dout <= 8'b00100100; // 1658 :  36 - 0x24
      11'h67B: dout <= 8'b00100100; // 1659 :  36 - 0x24
      11'h67C: dout <= 8'b00100100; // 1660 :  36 - 0x24
      11'h67D: dout <= 8'b00100100; // 1661 :  36 - 0x24
      11'h67E: dout <= 8'b00100100; // 1662 :  36 - 0x24
      11'h67F: dout <= 8'b00100100; // 1663 :  36 - 0x24
      11'h680: dout <= 8'b00100100; // 1664 :  36 - 0x24 -- line 0x14
      11'h681: dout <= 8'b00100100; // 1665 :  36 - 0x24
      11'h682: dout <= 8'b00100100; // 1666 :  36 - 0x24
      11'h683: dout <= 8'b00100100; // 1667 :  36 - 0x24
      11'h684: dout <= 8'b00100100; // 1668 :  36 - 0x24
      11'h685: dout <= 8'b00100100; // 1669 :  36 - 0x24
      11'h686: dout <= 8'b00100100; // 1670 :  36 - 0x24
      11'h687: dout <= 8'b00100100; // 1671 :  36 - 0x24
      11'h688: dout <= 8'b00100100; // 1672 :  36 - 0x24
      11'h689: dout <= 8'b00100100; // 1673 :  36 - 0x24
      11'h68A: dout <= 8'b00100100; // 1674 :  36 - 0x24
      11'h68B: dout <= 8'b00100100; // 1675 :  36 - 0x24
      11'h68C: dout <= 8'b00100100; // 1676 :  36 - 0x24
      11'h68D: dout <= 8'b00100100; // 1677 :  36 - 0x24
      11'h68E: dout <= 8'b00100100; // 1678 :  36 - 0x24
      11'h68F: dout <= 8'b00100100; // 1679 :  36 - 0x24
      11'h690: dout <= 8'b00100100; // 1680 :  36 - 0x24
      11'h691: dout <= 8'b00100100; // 1681 :  36 - 0x24
      11'h692: dout <= 8'b00100100; // 1682 :  36 - 0x24
      11'h693: dout <= 8'b00100100; // 1683 :  36 - 0x24
      11'h694: dout <= 8'b00100100; // 1684 :  36 - 0x24
      11'h695: dout <= 8'b00100100; // 1685 :  36 - 0x24
      11'h696: dout <= 8'b00100100; // 1686 :  36 - 0x24
      11'h697: dout <= 8'b00100100; // 1687 :  36 - 0x24
      11'h698: dout <= 8'b00100100; // 1688 :  36 - 0x24
      11'h699: dout <= 8'b00100100; // 1689 :  36 - 0x24
      11'h69A: dout <= 8'b00100100; // 1690 :  36 - 0x24
      11'h69B: dout <= 8'b00100100; // 1691 :  36 - 0x24
      11'h69C: dout <= 8'b00100100; // 1692 :  36 - 0x24
      11'h69D: dout <= 8'b00100100; // 1693 :  36 - 0x24
      11'h69E: dout <= 8'b00100100; // 1694 :  36 - 0x24
      11'h69F: dout <= 8'b00100100; // 1695 :  36 - 0x24
      11'h6A0: dout <= 8'b00100100; // 1696 :  36 - 0x24 -- line 0x15
      11'h6A1: dout <= 8'b00100100; // 1697 :  36 - 0x24
      11'h6A2: dout <= 8'b00100100; // 1698 :  36 - 0x24
      11'h6A3: dout <= 8'b00100100; // 1699 :  36 - 0x24
      11'h6A4: dout <= 8'b00100100; // 1700 :  36 - 0x24
      11'h6A5: dout <= 8'b00100100; // 1701 :  36 - 0x24
      11'h6A6: dout <= 8'b00100100; // 1702 :  36 - 0x24
      11'h6A7: dout <= 8'b00100100; // 1703 :  36 - 0x24
      11'h6A8: dout <= 8'b00100100; // 1704 :  36 - 0x24
      11'h6A9: dout <= 8'b00100100; // 1705 :  36 - 0x24
      11'h6AA: dout <= 8'b00100100; // 1706 :  36 - 0x24
      11'h6AB: dout <= 8'b00100100; // 1707 :  36 - 0x24
      11'h6AC: dout <= 8'b00100100; // 1708 :  36 - 0x24
      11'h6AD: dout <= 8'b00100100; // 1709 :  36 - 0x24
      11'h6AE: dout <= 8'b00100100; // 1710 :  36 - 0x24
      11'h6AF: dout <= 8'b00100100; // 1711 :  36 - 0x24
      11'h6B0: dout <= 8'b00100100; // 1712 :  36 - 0x24
      11'h6B1: dout <= 8'b00100100; // 1713 :  36 - 0x24
      11'h6B2: dout <= 8'b00100100; // 1714 :  36 - 0x24
      11'h6B3: dout <= 8'b00100100; // 1715 :  36 - 0x24
      11'h6B4: dout <= 8'b00100100; // 1716 :  36 - 0x24
      11'h6B5: dout <= 8'b00100100; // 1717 :  36 - 0x24
      11'h6B6: dout <= 8'b00100100; // 1718 :  36 - 0x24
      11'h6B7: dout <= 8'b00100100; // 1719 :  36 - 0x24
      11'h6B8: dout <= 8'b00100100; // 1720 :  36 - 0x24
      11'h6B9: dout <= 8'b00100100; // 1721 :  36 - 0x24
      11'h6BA: dout <= 8'b00100100; // 1722 :  36 - 0x24
      11'h6BB: dout <= 8'b00100100; // 1723 :  36 - 0x24
      11'h6BC: dout <= 8'b00100100; // 1724 :  36 - 0x24
      11'h6BD: dout <= 8'b00100100; // 1725 :  36 - 0x24
      11'h6BE: dout <= 8'b00100100; // 1726 :  36 - 0x24
      11'h6BF: dout <= 8'b00100100; // 1727 :  36 - 0x24
      11'h6C0: dout <= 8'b00100100; // 1728 :  36 - 0x24 -- line 0x16
      11'h6C1: dout <= 8'b00100100; // 1729 :  36 - 0x24
      11'h6C2: dout <= 8'b00100100; // 1730 :  36 - 0x24
      11'h6C3: dout <= 8'b00100100; // 1731 :  36 - 0x24
      11'h6C4: dout <= 8'b00100100; // 1732 :  36 - 0x24
      11'h6C5: dout <= 8'b00100100; // 1733 :  36 - 0x24
      11'h6C6: dout <= 8'b00100100; // 1734 :  36 - 0x24
      11'h6C7: dout <= 8'b00100100; // 1735 :  36 - 0x24
      11'h6C8: dout <= 8'b00100100; // 1736 :  36 - 0x24
      11'h6C9: dout <= 8'b00100100; // 1737 :  36 - 0x24
      11'h6CA: dout <= 8'b00100100; // 1738 :  36 - 0x24
      11'h6CB: dout <= 8'b00100100; // 1739 :  36 - 0x24
      11'h6CC: dout <= 8'b00100100; // 1740 :  36 - 0x24
      11'h6CD: dout <= 8'b00100100; // 1741 :  36 - 0x24
      11'h6CE: dout <= 8'b00100100; // 1742 :  36 - 0x24
      11'h6CF: dout <= 8'b00100100; // 1743 :  36 - 0x24
      11'h6D0: dout <= 8'b00100100; // 1744 :  36 - 0x24
      11'h6D1: dout <= 8'b00100100; // 1745 :  36 - 0x24
      11'h6D2: dout <= 8'b00100100; // 1746 :  36 - 0x24
      11'h6D3: dout <= 8'b00100100; // 1747 :  36 - 0x24
      11'h6D4: dout <= 8'b00100100; // 1748 :  36 - 0x24
      11'h6D5: dout <= 8'b00100100; // 1749 :  36 - 0x24
      11'h6D6: dout <= 8'b00100100; // 1750 :  36 - 0x24
      11'h6D7: dout <= 8'b00100100; // 1751 :  36 - 0x24
      11'h6D8: dout <= 8'b00100100; // 1752 :  36 - 0x24
      11'h6D9: dout <= 8'b00100100; // 1753 :  36 - 0x24
      11'h6DA: dout <= 8'b00100100; // 1754 :  36 - 0x24
      11'h6DB: dout <= 8'b00100100; // 1755 :  36 - 0x24
      11'h6DC: dout <= 8'b00100100; // 1756 :  36 - 0x24
      11'h6DD: dout <= 8'b00100100; // 1757 :  36 - 0x24
      11'h6DE: dout <= 8'b00100100; // 1758 :  36 - 0x24
      11'h6DF: dout <= 8'b00100100; // 1759 :  36 - 0x24
      11'h6E0: dout <= 8'b00100100; // 1760 :  36 - 0x24 -- line 0x17
      11'h6E1: dout <= 8'b00100100; // 1761 :  36 - 0x24
      11'h6E2: dout <= 8'b00110001; // 1762 :  49 - 0x31
      11'h6E3: dout <= 8'b00110010; // 1763 :  50 - 0x32
      11'h6E4: dout <= 8'b00100100; // 1764 :  36 - 0x24
      11'h6E5: dout <= 8'b00100100; // 1765 :  36 - 0x24
      11'h6E6: dout <= 8'b00100100; // 1766 :  36 - 0x24
      11'h6E7: dout <= 8'b00100100; // 1767 :  36 - 0x24
      11'h6E8: dout <= 8'b00100100; // 1768 :  36 - 0x24
      11'h6E9: dout <= 8'b00100100; // 1769 :  36 - 0x24
      11'h6EA: dout <= 8'b00100100; // 1770 :  36 - 0x24
      11'h6EB: dout <= 8'b00100100; // 1771 :  36 - 0x24
      11'h6EC: dout <= 8'b00100100; // 1772 :  36 - 0x24
      11'h6ED: dout <= 8'b00100100; // 1773 :  36 - 0x24
      11'h6EE: dout <= 8'b00100100; // 1774 :  36 - 0x24
      11'h6EF: dout <= 8'b00100100; // 1775 :  36 - 0x24
      11'h6F0: dout <= 8'b00100100; // 1776 :  36 - 0x24
      11'h6F1: dout <= 8'b00100100; // 1777 :  36 - 0x24
      11'h6F2: dout <= 8'b00100100; // 1778 :  36 - 0x24
      11'h6F3: dout <= 8'b00100100; // 1779 :  36 - 0x24
      11'h6F4: dout <= 8'b00100100; // 1780 :  36 - 0x24
      11'h6F5: dout <= 8'b00100100; // 1781 :  36 - 0x24
      11'h6F6: dout <= 8'b00100100; // 1782 :  36 - 0x24
      11'h6F7: dout <= 8'b00100100; // 1783 :  36 - 0x24
      11'h6F8: dout <= 8'b00100100; // 1784 :  36 - 0x24
      11'h6F9: dout <= 8'b00100100; // 1785 :  36 - 0x24
      11'h6FA: dout <= 8'b00100100; // 1786 :  36 - 0x24
      11'h6FB: dout <= 8'b00100100; // 1787 :  36 - 0x24
      11'h6FC: dout <= 8'b00100100; // 1788 :  36 - 0x24
      11'h6FD: dout <= 8'b00100100; // 1789 :  36 - 0x24
      11'h6FE: dout <= 8'b00100100; // 1790 :  36 - 0x24
      11'h6FF: dout <= 8'b00100100; // 1791 :  36 - 0x24
      11'h700: dout <= 8'b00100100; // 1792 :  36 - 0x24 -- line 0x18
      11'h701: dout <= 8'b00110000; // 1793 :  48 - 0x30
      11'h702: dout <= 8'b00100110; // 1794 :  38 - 0x26
      11'h703: dout <= 8'b00110100; // 1795 :  52 - 0x34
      11'h704: dout <= 8'b00110011; // 1796 :  51 - 0x33
      11'h705: dout <= 8'b00100100; // 1797 :  36 - 0x24
      11'h706: dout <= 8'b00100100; // 1798 :  36 - 0x24
      11'h707: dout <= 8'b00100100; // 1799 :  36 - 0x24
      11'h708: dout <= 8'b00100100; // 1800 :  36 - 0x24
      11'h709: dout <= 8'b00100100; // 1801 :  36 - 0x24
      11'h70A: dout <= 8'b00100100; // 1802 :  36 - 0x24
      11'h70B: dout <= 8'b00100100; // 1803 :  36 - 0x24
      11'h70C: dout <= 8'b00100100; // 1804 :  36 - 0x24
      11'h70D: dout <= 8'b00100100; // 1805 :  36 - 0x24
      11'h70E: dout <= 8'b00100100; // 1806 :  36 - 0x24
      11'h70F: dout <= 8'b00100100; // 1807 :  36 - 0x24
      11'h710: dout <= 8'b00100100; // 1808 :  36 - 0x24
      11'h711: dout <= 8'b00100100; // 1809 :  36 - 0x24
      11'h712: dout <= 8'b00100100; // 1810 :  36 - 0x24
      11'h713: dout <= 8'b00100100; // 1811 :  36 - 0x24
      11'h714: dout <= 8'b00100100; // 1812 :  36 - 0x24
      11'h715: dout <= 8'b00100100; // 1813 :  36 - 0x24
      11'h716: dout <= 8'b00100100; // 1814 :  36 - 0x24
      11'h717: dout <= 8'b00100100; // 1815 :  36 - 0x24
      11'h718: dout <= 8'b00100100; // 1816 :  36 - 0x24
      11'h719: dout <= 8'b00100100; // 1817 :  36 - 0x24
      11'h71A: dout <= 8'b00100100; // 1818 :  36 - 0x24
      11'h71B: dout <= 8'b00100100; // 1819 :  36 - 0x24
      11'h71C: dout <= 8'b00100100; // 1820 :  36 - 0x24
      11'h71D: dout <= 8'b00100100; // 1821 :  36 - 0x24
      11'h71E: dout <= 8'b00100100; // 1822 :  36 - 0x24
      11'h71F: dout <= 8'b00100100; // 1823 :  36 - 0x24
      11'h720: dout <= 8'b00110000; // 1824 :  48 - 0x30 -- line 0x19
      11'h721: dout <= 8'b00100110; // 1825 :  38 - 0x26
      11'h722: dout <= 8'b00100110; // 1826 :  38 - 0x26
      11'h723: dout <= 8'b00100110; // 1827 :  38 - 0x26
      11'h724: dout <= 8'b00100110; // 1828 :  38 - 0x26
      11'h725: dout <= 8'b00110011; // 1829 :  51 - 0x33
      11'h726: dout <= 8'b00100100; // 1830 :  36 - 0x24
      11'h727: dout <= 8'b00100100; // 1831 :  36 - 0x24
      11'h728: dout <= 8'b00100100; // 1832 :  36 - 0x24
      11'h729: dout <= 8'b00100100; // 1833 :  36 - 0x24
      11'h72A: dout <= 8'b00100100; // 1834 :  36 - 0x24
      11'h72B: dout <= 8'b00100100; // 1835 :  36 - 0x24
      11'h72C: dout <= 8'b00100100; // 1836 :  36 - 0x24
      11'h72D: dout <= 8'b00100100; // 1837 :  36 - 0x24
      11'h72E: dout <= 8'b00100100; // 1838 :  36 - 0x24
      11'h72F: dout <= 8'b00110101; // 1839 :  53 - 0x35
      11'h730: dout <= 8'b00100100; // 1840 :  36 - 0x24
      11'h731: dout <= 8'b00100100; // 1841 :  36 - 0x24
      11'h732: dout <= 8'b00100100; // 1842 :  36 - 0x24
      11'h733: dout <= 8'b00100100; // 1843 :  36 - 0x24
      11'h734: dout <= 8'b00100100; // 1844 :  36 - 0x24
      11'h735: dout <= 8'b00100100; // 1845 :  36 - 0x24
      11'h736: dout <= 8'b00100100; // 1846 :  36 - 0x24
      11'h737: dout <= 8'b00100100; // 1847 :  36 - 0x24
      11'h738: dout <= 8'b00100100; // 1848 :  36 - 0x24
      11'h739: dout <= 8'b00100100; // 1849 :  36 - 0x24
      11'h73A: dout <= 8'b00100100; // 1850 :  36 - 0x24
      11'h73B: dout <= 8'b00100100; // 1851 :  36 - 0x24
      11'h73C: dout <= 8'b00100100; // 1852 :  36 - 0x24
      11'h73D: dout <= 8'b00100100; // 1853 :  36 - 0x24
      11'h73E: dout <= 8'b00100100; // 1854 :  36 - 0x24
      11'h73F: dout <= 8'b00100100; // 1855 :  36 - 0x24
      11'h740: dout <= 8'b10110100; // 1856 : 180 - 0xb4 -- line 0x1a
      11'h741: dout <= 8'b10110101; // 1857 : 181 - 0xb5
      11'h742: dout <= 8'b10110100; // 1858 : 180 - 0xb4
      11'h743: dout <= 8'b10110101; // 1859 : 181 - 0xb5
      11'h744: dout <= 8'b10110100; // 1860 : 180 - 0xb4
      11'h745: dout <= 8'b10110101; // 1861 : 181 - 0xb5
      11'h746: dout <= 8'b10110100; // 1862 : 180 - 0xb4
      11'h747: dout <= 8'b10110101; // 1863 : 181 - 0xb5
      11'h748: dout <= 8'b10110100; // 1864 : 180 - 0xb4
      11'h749: dout <= 8'b10110101; // 1865 : 181 - 0xb5
      11'h74A: dout <= 8'b10110100; // 1866 : 180 - 0xb4
      11'h74B: dout <= 8'b10110101; // 1867 : 181 - 0xb5
      11'h74C: dout <= 8'b10110100; // 1868 : 180 - 0xb4
      11'h74D: dout <= 8'b10110101; // 1869 : 181 - 0xb5
      11'h74E: dout <= 8'b10110100; // 1870 : 180 - 0xb4
      11'h74F: dout <= 8'b10110101; // 1871 : 181 - 0xb5
      11'h750: dout <= 8'b00100100; // 1872 :  36 - 0x24
      11'h751: dout <= 8'b00100100; // 1873 :  36 - 0x24
      11'h752: dout <= 8'b00100100; // 1874 :  36 - 0x24
      11'h753: dout <= 8'b00100100; // 1875 :  36 - 0x24
      11'h754: dout <= 8'b00100100; // 1876 :  36 - 0x24
      11'h755: dout <= 8'b00100100; // 1877 :  36 - 0x24
      11'h756: dout <= 8'b00100100; // 1878 :  36 - 0x24
      11'h757: dout <= 8'b00100100; // 1879 :  36 - 0x24
      11'h758: dout <= 8'b00100100; // 1880 :  36 - 0x24
      11'h759: dout <= 8'b00100100; // 1881 :  36 - 0x24
      11'h75A: dout <= 8'b00100100; // 1882 :  36 - 0x24
      11'h75B: dout <= 8'b00100100; // 1883 :  36 - 0x24
      11'h75C: dout <= 8'b00100100; // 1884 :  36 - 0x24
      11'h75D: dout <= 8'b00100100; // 1885 :  36 - 0x24
      11'h75E: dout <= 8'b00100100; // 1886 :  36 - 0x24
      11'h75F: dout <= 8'b00100100; // 1887 :  36 - 0x24
      11'h760: dout <= 8'b10110110; // 1888 : 182 - 0xb6 -- line 0x1b
      11'h761: dout <= 8'b10110111; // 1889 : 183 - 0xb7
      11'h762: dout <= 8'b10110110; // 1890 : 182 - 0xb6
      11'h763: dout <= 8'b10110111; // 1891 : 183 - 0xb7
      11'h764: dout <= 8'b10110110; // 1892 : 182 - 0xb6
      11'h765: dout <= 8'b10110111; // 1893 : 183 - 0xb7
      11'h766: dout <= 8'b10110110; // 1894 : 182 - 0xb6
      11'h767: dout <= 8'b10110111; // 1895 : 183 - 0xb7
      11'h768: dout <= 8'b10110110; // 1896 : 182 - 0xb6
      11'h769: dout <= 8'b10110111; // 1897 : 183 - 0xb7
      11'h76A: dout <= 8'b10110110; // 1898 : 182 - 0xb6
      11'h76B: dout <= 8'b10110111; // 1899 : 183 - 0xb7
      11'h76C: dout <= 8'b10110110; // 1900 : 182 - 0xb6
      11'h76D: dout <= 8'b10110111; // 1901 : 183 - 0xb7
      11'h76E: dout <= 8'b10110110; // 1902 : 182 - 0xb6
      11'h76F: dout <= 8'b10110111; // 1903 : 183 - 0xb7
      11'h770: dout <= 8'b00100100; // 1904 :  36 - 0x24
      11'h771: dout <= 8'b00100100; // 1905 :  36 - 0x24
      11'h772: dout <= 8'b00100100; // 1906 :  36 - 0x24
      11'h773: dout <= 8'b00100100; // 1907 :  36 - 0x24
      11'h774: dout <= 8'b00100100; // 1908 :  36 - 0x24
      11'h775: dout <= 8'b00100100; // 1909 :  36 - 0x24
      11'h776: dout <= 8'b00100100; // 1910 :  36 - 0x24
      11'h777: dout <= 8'b00100100; // 1911 :  36 - 0x24
      11'h778: dout <= 8'b00100100; // 1912 :  36 - 0x24
      11'h779: dout <= 8'b00100100; // 1913 :  36 - 0x24
      11'h77A: dout <= 8'b00100100; // 1914 :  36 - 0x24
      11'h77B: dout <= 8'b00100100; // 1915 :  36 - 0x24
      11'h77C: dout <= 8'b00100100; // 1916 :  36 - 0x24
      11'h77D: dout <= 8'b00100100; // 1917 :  36 - 0x24
      11'h77E: dout <= 8'b00100100; // 1918 :  36 - 0x24
      11'h77F: dout <= 8'b00100100; // 1919 :  36 - 0x24
      11'h780: dout <= 8'b10110100; // 1920 : 180 - 0xb4 -- line 0x1c
      11'h781: dout <= 8'b10110101; // 1921 : 181 - 0xb5
      11'h782: dout <= 8'b10110100; // 1922 : 180 - 0xb4
      11'h783: dout <= 8'b10110101; // 1923 : 181 - 0xb5
      11'h784: dout <= 8'b10110100; // 1924 : 180 - 0xb4
      11'h785: dout <= 8'b10110101; // 1925 : 181 - 0xb5
      11'h786: dout <= 8'b10110100; // 1926 : 180 - 0xb4
      11'h787: dout <= 8'b10110101; // 1927 : 181 - 0xb5
      11'h788: dout <= 8'b10110100; // 1928 : 180 - 0xb4
      11'h789: dout <= 8'b10110101; // 1929 : 181 - 0xb5
      11'h78A: dout <= 8'b10110100; // 1930 : 180 - 0xb4
      11'h78B: dout <= 8'b10110101; // 1931 : 181 - 0xb5
      11'h78C: dout <= 8'b10110100; // 1932 : 180 - 0xb4
      11'h78D: dout <= 8'b10110101; // 1933 : 181 - 0xb5
      11'h78E: dout <= 8'b10110100; // 1934 : 180 - 0xb4
      11'h78F: dout <= 8'b10110101; // 1935 : 181 - 0xb5
      11'h790: dout <= 8'b00100100; // 1936 :  36 - 0x24
      11'h791: dout <= 8'b00100100; // 1937 :  36 - 0x24
      11'h792: dout <= 8'b00100100; // 1938 :  36 - 0x24
      11'h793: dout <= 8'b00100100; // 1939 :  36 - 0x24
      11'h794: dout <= 8'b00100100; // 1940 :  36 - 0x24
      11'h795: dout <= 8'b00100100; // 1941 :  36 - 0x24
      11'h796: dout <= 8'b00100100; // 1942 :  36 - 0x24
      11'h797: dout <= 8'b00100100; // 1943 :  36 - 0x24
      11'h798: dout <= 8'b00100100; // 1944 :  36 - 0x24
      11'h799: dout <= 8'b00100100; // 1945 :  36 - 0x24
      11'h79A: dout <= 8'b00100100; // 1946 :  36 - 0x24
      11'h79B: dout <= 8'b00100100; // 1947 :  36 - 0x24
      11'h79C: dout <= 8'b00100100; // 1948 :  36 - 0x24
      11'h79D: dout <= 8'b00100100; // 1949 :  36 - 0x24
      11'h79E: dout <= 8'b00100100; // 1950 :  36 - 0x24
      11'h79F: dout <= 8'b00100100; // 1951 :  36 - 0x24
      11'h7A0: dout <= 8'b10110110; // 1952 : 182 - 0xb6 -- line 0x1d
      11'h7A1: dout <= 8'b10110111; // 1953 : 183 - 0xb7
      11'h7A2: dout <= 8'b10110110; // 1954 : 182 - 0xb6
      11'h7A3: dout <= 8'b10110111; // 1955 : 183 - 0xb7
      11'h7A4: dout <= 8'b10110110; // 1956 : 182 - 0xb6
      11'h7A5: dout <= 8'b10110111; // 1957 : 183 - 0xb7
      11'h7A6: dout <= 8'b10110110; // 1958 : 182 - 0xb6
      11'h7A7: dout <= 8'b10110111; // 1959 : 183 - 0xb7
      11'h7A8: dout <= 8'b10110110; // 1960 : 182 - 0xb6
      11'h7A9: dout <= 8'b10110111; // 1961 : 183 - 0xb7
      11'h7AA: dout <= 8'b10110110; // 1962 : 182 - 0xb6
      11'h7AB: dout <= 8'b10110111; // 1963 : 183 - 0xb7
      11'h7AC: dout <= 8'b10110110; // 1964 : 182 - 0xb6
      11'h7AD: dout <= 8'b10110111; // 1965 : 183 - 0xb7
      11'h7AE: dout <= 8'b10110110; // 1966 : 182 - 0xb6
      11'h7AF: dout <= 8'b10110111; // 1967 : 183 - 0xb7
      11'h7B0: dout <= 8'b00100100; // 1968 :  36 - 0x24
      11'h7B1: dout <= 8'b00100100; // 1969 :  36 - 0x24
      11'h7B2: dout <= 8'b00100100; // 1970 :  36 - 0x24
      11'h7B3: dout <= 8'b00100100; // 1971 :  36 - 0x24
      11'h7B4: dout <= 8'b00100100; // 1972 :  36 - 0x24
      11'h7B5: dout <= 8'b00100100; // 1973 :  36 - 0x24
      11'h7B6: dout <= 8'b00100100; // 1974 :  36 - 0x24
      11'h7B7: dout <= 8'b00100100; // 1975 :  36 - 0x24
      11'h7B8: dout <= 8'b00100100; // 1976 :  36 - 0x24
      11'h7B9: dout <= 8'b00100100; // 1977 :  36 - 0x24
      11'h7BA: dout <= 8'b00100100; // 1978 :  36 - 0x24
      11'h7BB: dout <= 8'b00100100; // 1979 :  36 - 0x24
      11'h7BC: dout <= 8'b00100100; // 1980 :  36 - 0x24
      11'h7BD: dout <= 8'b00100100; // 1981 :  36 - 0x24
      11'h7BE: dout <= 8'b00100100; // 1982 :  36 - 0x24
      11'h7BF: dout <= 8'b00100100; // 1983 :  36 - 0x24
        //-- Attribute Table 1----
      11'h7C0: dout <= 8'b00000000; // 1984 :   0 - 0x0
      11'h7C1: dout <= 8'b00000000; // 1985 :   0 - 0x0
      11'h7C2: dout <= 8'b00000000; // 1986 :   0 - 0x0
      11'h7C3: dout <= 8'b00000000; // 1987 :   0 - 0x0
      11'h7C4: dout <= 8'b00000000; // 1988 :   0 - 0x0
      11'h7C5: dout <= 8'b00000000; // 1989 :   0 - 0x0
      11'h7C6: dout <= 8'b00000000; // 1990 :   0 - 0x0
      11'h7C7: dout <= 8'b00000000; // 1991 :   0 - 0x0
      11'h7C8: dout <= 8'b00000000; // 1992 :   0 - 0x0
      11'h7C9: dout <= 8'b10001000; // 1993 : 136 - 0x88
      11'h7CA: dout <= 8'b10101010; // 1994 : 170 - 0xaa
      11'h7CB: dout <= 8'b00000000; // 1995 :   0 - 0x0
      11'h7CC: dout <= 8'b00000000; // 1996 :   0 - 0x0
      11'h7CD: dout <= 8'b00000000; // 1997 :   0 - 0x0
      11'h7CE: dout <= 8'b00000000; // 1998 :   0 - 0x0
      11'h7CF: dout <= 8'b00000000; // 1999 :   0 - 0x0
      11'h7D0: dout <= 8'b00000000; // 2000 :   0 - 0x0
      11'h7D1: dout <= 8'b00000000; // 2001 :   0 - 0x0
      11'h7D2: dout <= 8'b00000000; // 2002 :   0 - 0x0
      11'h7D3: dout <= 8'b00110000; // 2003 :  48 - 0x30
      11'h7D4: dout <= 8'b00000000; // 2004 :   0 - 0x0
      11'h7D5: dout <= 8'b00000000; // 2005 :   0 - 0x0
      11'h7D6: dout <= 8'b00000000; // 2006 :   0 - 0x0
      11'h7D7: dout <= 8'b00000000; // 2007 :   0 - 0x0
      11'h7D8: dout <= 8'b00000000; // 2008 :   0 - 0x0
      11'h7D9: dout <= 8'b00000000; // 2009 :   0 - 0x0
      11'h7DA: dout <= 8'b00000000; // 2010 :   0 - 0x0
      11'h7DB: dout <= 8'b00000000; // 2011 :   0 - 0x0
      11'h7DC: dout <= 8'b00000000; // 2012 :   0 - 0x0
      11'h7DD: dout <= 8'b00000000; // 2013 :   0 - 0x0
      11'h7DE: dout <= 8'b00000000; // 2014 :   0 - 0x0
      11'h7DF: dout <= 8'b00000000; // 2015 :   0 - 0x0
      11'h7E0: dout <= 8'b00110000; // 2016 :  48 - 0x30
      11'h7E1: dout <= 8'b00000000; // 2017 :   0 - 0x0
      11'h7E2: dout <= 8'b11010000; // 2018 : 208 - 0xd0
      11'h7E3: dout <= 8'b11010000; // 2019 : 208 - 0xd0
      11'h7E4: dout <= 8'b00000000; // 2020 :   0 - 0x0
      11'h7E5: dout <= 8'b00000000; // 2021 :   0 - 0x0
      11'h7E6: dout <= 8'b00000000; // 2022 :   0 - 0x0
      11'h7E7: dout <= 8'b00000000; // 2023 :   0 - 0x0
      11'h7E8: dout <= 8'b00000000; // 2024 :   0 - 0x0
      11'h7E9: dout <= 8'b00000000; // 2025 :   0 - 0x0
      11'h7EA: dout <= 8'b00000000; // 2026 :   0 - 0x0
      11'h7EB: dout <= 8'b00000000; // 2027 :   0 - 0x0
      11'h7EC: dout <= 8'b00000000; // 2028 :   0 - 0x0
      11'h7ED: dout <= 8'b00000000; // 2029 :   0 - 0x0
      11'h7EE: dout <= 8'b00000000; // 2030 :   0 - 0x0
      11'h7EF: dout <= 8'b00000000; // 2031 :   0 - 0x0
      11'h7F0: dout <= 8'b01010000; // 2032 :  80 - 0x50
      11'h7F1: dout <= 8'b01010000; // 2033 :  80 - 0x50
      11'h7F2: dout <= 8'b01010000; // 2034 :  80 - 0x50
      11'h7F3: dout <= 8'b01010000; // 2035 :  80 - 0x50
      11'h7F4: dout <= 8'b00000000; // 2036 :   0 - 0x0
      11'h7F5: dout <= 8'b00000000; // 2037 :   0 - 0x0
      11'h7F6: dout <= 8'b00000000; // 2038 :   0 - 0x0
      11'h7F7: dout <= 8'b00000000; // 2039 :   0 - 0x0
      11'h7F8: dout <= 8'b00000101; // 2040 :   5 - 0x5
      11'h7F9: dout <= 8'b00000101; // 2041 :   5 - 0x5
      11'h7FA: dout <= 8'b00000101; // 2042 :   5 - 0x5
      11'h7FB: dout <= 8'b00000101; // 2043 :   5 - 0x5
      11'h7FC: dout <= 8'b00000000; // 2044 :   0 - 0x0
      11'h7FD: dout <= 8'b00000000; // 2045 :   0 - 0x0
      11'h7FE: dout <= 8'b00000000; // 2046 :   0 - 0x0
      11'h7FF: dout <= 8'b00000000; // 2047 :   0 - 0x0
    endcase
  end

endmodule
