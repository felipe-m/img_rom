---   Background Pattern table BOTH COLOR PLANES
-- https://wiki.nesdev.com/w/index.php/PPU_pattern_tables
--- Autcmatically generated VHDL ROM from a NES memory file----


---  Original memory dump file name: nova_ptable.dmp --
------ Felipe Machado -----------------------------------
------ Area de Tecnologia Electronica -----------
------ Universidad Rey Juan Carlos ----------------------
------ https://github.com/felipe-m ----------------------
---------------------------------------------------------
----- Memory without clock -----

----- Ports ---------------------------------------------
-- Inputs   ---------------------------------------------
--   -- clk  :  clock signal
--    addr :  memory address
-- Salidas  ---------------------------------------------
--    dout :  memory data out  (no clock: in the same clock cycle)


library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;


entity ROM_PTABLE_NOVA_BG is
  port (
    --clk  : in  std_logic;   -- clock
    addr : in  std_logic_vector(12-1 downto 0);  --4096 memory positions
    dout : out std_logic_vector(8-1 downto 0) -- memory data width
  );
end ROM_PTABLE_NOVA_BG;

architecture BEHAVIORAL of ROM_PTABLE_NOVA_BG is
  signal addr_int  : natural range 0 to 2**12-1;
  type memostruct is array (natural range<>) of std_logic_vector(8-1 downto 0);
  constant table_mem : memostruct := (
                --    address   :    value 
                --  dec -  hex  :  dec - hex
          -- Background pattern Table both color planes
    "11111111", --    0 -  0x0  :  255 - 0xff -- Background 0x0
    "11111111", --    1 -  0x1  :  255 - 0xff
    "11000000", --    2 -  0x2  :  192 - 0xc0
    "11000000", --    3 -  0x3  :  192 - 0xc0
    "11000000", --    4 -  0x4  :  192 - 0xc0
    "11000000", --    5 -  0x5  :  192 - 0xc0
    "11010101", --    6 -  0x6  :  213 - 0xd5
    "11111111", --    7 -  0x7  :  255 - 0xff
    "00000000", --    8 -  0x8  :    0 - 0x0 -- plane 1
    "01111111", --    9 -  0x9  :  127 - 0x7f
    "01111111", --   10 -  0xa  :  127 - 0x7f
    "01111111", --   11 -  0xb  :  127 - 0x7f
    "01111111", --   12 -  0xc  :  127 - 0x7f
    "01111111", --   13 -  0xd  :  127 - 0x7f
    "01101010", --   14 -  0xe  :  106 - 0x6a
    "00000000", --   15 -  0xf  :    0 - 0x0
    "11111111", --   16 - 0x10  :  255 - 0xff -- Background 0x1
    "11111111", --   17 - 0x11  :  255 - 0xff
    "11001110", --   18 - 0x12  :  206 - 0xce
    "11000110", --   19 - 0x13  :  198 - 0xc6
    "11001110", --   20 - 0x14  :  206 - 0xce
    "11000110", --   21 - 0x15  :  198 - 0xc6
    "11101110", --   22 - 0x16  :  238 - 0xee
    "11111111", --   23 - 0x17  :  255 - 0xff
    "00000000", --   24 - 0x18  :    0 - 0x0 -- plane 1
    "01111011", --   25 - 0x19  :  123 - 0x7b
    "01110011", --   26 - 0x1a  :  115 - 0x73
    "01111011", --   27 - 0x1b  :  123 - 0x7b
    "01110011", --   28 - 0x1c  :  115 - 0x73
    "01111011", --   29 - 0x1d  :  123 - 0x7b
    "01010011", --   30 - 0x1e  :   83 - 0x53
    "00000000", --   31 - 0x1f  :    0 - 0x0
    "11111111", --   32 - 0x20  :  255 - 0xff -- Background 0x2
    "11111111", --   33 - 0x21  :  255 - 0xff
    "01110001", --   34 - 0x22  :  113 - 0x71
    "00110011", --   35 - 0x23  :   51 - 0x33
    "01110001", --   36 - 0x24  :  113 - 0x71
    "00110011", --   37 - 0x25  :   51 - 0x33
    "01110101", --   38 - 0x26  :  117 - 0x75
    "11111111", --   39 - 0x27  :  255 - 0xff
    "00000000", --   40 - 0x28  :    0 - 0x0 -- plane 1
    "11011110", --   41 - 0x29  :  222 - 0xde
    "10011110", --   42 - 0x2a  :  158 - 0x9e
    "11011100", --   43 - 0x2b  :  220 - 0xdc
    "10011110", --   44 - 0x2c  :  158 - 0x9e
    "11011100", --   45 - 0x2d  :  220 - 0xdc
    "10011010", --   46 - 0x2e  :  154 - 0x9a
    "00000000", --   47 - 0x2f  :    0 - 0x0
    "11111111", --   48 - 0x30  :  255 - 0xff -- Background 0x3
    "11111111", --   49 - 0x31  :  255 - 0xff
    "00000011", --   50 - 0x32  :    3 - 0x3
    "00000001", --   51 - 0x33  :    1 - 0x1
    "00000011", --   52 - 0x34  :    3 - 0x3
    "00000001", --   53 - 0x35  :    1 - 0x1
    "10101011", --   54 - 0x36  :  171 - 0xab
    "11111111", --   55 - 0x37  :  255 - 0xff
    "00000000", --   56 - 0x38  :    0 - 0x0 -- plane 1
    "11111110", --   57 - 0x39  :  254 - 0xfe
    "11111100", --   58 - 0x3a  :  252 - 0xfc
    "11111110", --   59 - 0x3b  :  254 - 0xfe
    "11111100", --   60 - 0x3c  :  252 - 0xfc
    "11111110", --   61 - 0x3d  :  254 - 0xfe
    "01010100", --   62 - 0x3e  :   84 - 0x54
    "00000000", --   63 - 0x3f  :    0 - 0x0
    "11111111", --   64 - 0x40  :  255 - 0xff -- Background 0x4
    "11111111", --   65 - 0x41  :  255 - 0xff
    "11100000", --   66 - 0x42  :  224 - 0xe0
    "11000110", --   67 - 0x43  :  198 - 0xc6
    "11000110", --   68 - 0x44  :  198 - 0xc6
    "11110110", --   69 - 0x45  :  246 - 0xf6
    "11110000", --   70 - 0x46  :  240 - 0xf0
    "11110001", --   71 - 0x47  :  241 - 0xf1
    "00000000", --   72 - 0x48  :    0 - 0x0 -- plane 1
    "01111111", --   73 - 0x49  :  127 - 0x7f
    "01011111", --   74 - 0x4a  :   95 - 0x5f
    "01111001", --   75 - 0x4b  :  121 - 0x79
    "01111001", --   76 - 0x4c  :  121 - 0x79
    "01001001", --   77 - 0x4d  :   73 - 0x49
    "01001111", --   78 - 0x4e  :   79 - 0x4f
    "01001110", --   79 - 0x4f  :   78 - 0x4e
    "11000111", --   80 - 0x50  :  199 - 0xc7 -- Background 0x5
    "11001111", --   81 - 0x51  :  207 - 0xcf
    "11011111", --   82 - 0x52  :  223 - 0xdf
    "11011111", --   83 - 0x53  :  223 - 0xdf
    "11001110", --   84 - 0x54  :  206 - 0xce
    "11100000", --   85 - 0x55  :  224 - 0xe0
    "11111111", --   86 - 0x56  :  255 - 0xff
    "11111111", --   87 - 0x57  :  255 - 0xff
    "01111000", --   88 - 0x58  :  120 - 0x78 -- plane 1
    "01110000", --   89 - 0x59  :  112 - 0x70
    "01100000", --   90 - 0x5a  :   96 - 0x60
    "01100000", --   91 - 0x5b  :   96 - 0x60
    "01110001", --   92 - 0x5c  :  113 - 0x71
    "01011111", --   93 - 0x5d  :   95 - 0x5f
    "01111111", --   94 - 0x5e  :  127 - 0x7f
    "00000000", --   95 - 0x5f  :    0 - 0x0
    "11111111", --   96 - 0x60  :  255 - 0xff -- Background 0x6
    "11111111", --   97 - 0x61  :  255 - 0xff
    "00000111", --   98 - 0x62  :    7 - 0x7
    "01100011", --   99 - 0x63  :   99 - 0x63
    "01100011", --  100 - 0x64  :   99 - 0x63
    "01101111", --  101 - 0x65  :  111 - 0x6f
    "00001111", --  102 - 0x66  :   15 - 0xf
    "10001111", --  103 - 0x67  :  143 - 0x8f
    "00000000", --  104 - 0x68  :    0 - 0x0 -- plane 1
    "11111110", --  105 - 0x69  :  254 - 0xfe
    "11111010", --  106 - 0x6a  :  250 - 0xfa
    "10011110", --  107 - 0x6b  :  158 - 0x9e
    "10011110", --  108 - 0x6c  :  158 - 0x9e
    "10010010", --  109 - 0x6d  :  146 - 0x92
    "11110010", --  110 - 0x6e  :  242 - 0xf2
    "01110010", --  111 - 0x6f  :  114 - 0x72
    "11100011", --  112 - 0x70  :  227 - 0xe3 -- Background 0x7
    "11110011", --  113 - 0x71  :  243 - 0xf3
    "11111011", --  114 - 0x72  :  251 - 0xfb
    "11111011", --  115 - 0x73  :  251 - 0xfb
    "01110011", --  116 - 0x74  :  115 - 0x73
    "00000111", --  117 - 0x75  :    7 - 0x7
    "11111111", --  118 - 0x76  :  255 - 0xff
    "11111111", --  119 - 0x77  :  255 - 0xff
    "00011110", --  120 - 0x78  :   30 - 0x1e -- plane 1
    "00001110", --  121 - 0x79  :   14 - 0xe
    "00000110", --  122 - 0x7a  :    6 - 0x6
    "00000110", --  123 - 0x7b  :    6 - 0x6
    "10001110", --  124 - 0x7c  :  142 - 0x8e
    "11111010", --  125 - 0x7d  :  250 - 0xfa
    "11111110", --  126 - 0x7e  :  254 - 0xfe
    "00000000", --  127 - 0x7f  :    0 - 0x0
    "11111111", --  128 - 0x80  :  255 - 0xff -- Background 0x8
    "11010101", --  129 - 0x81  :  213 - 0xd5
    "10101010", --  130 - 0x82  :  170 - 0xaa
    "11010101", --  131 - 0x83  :  213 - 0xd5
    "10101010", --  132 - 0x84  :  170 - 0xaa
    "11010101", --  133 - 0x85  :  213 - 0xd5
    "10101010", --  134 - 0x86  :  170 - 0xaa
    "11010101", --  135 - 0x87  :  213 - 0xd5
    "00000000", --  136 - 0x88  :    0 - 0x0 -- plane 1
    "01111111", --  137 - 0x89  :  127 - 0x7f
    "01011111", --  138 - 0x8a  :   95 - 0x5f
    "01111111", --  139 - 0x8b  :  127 - 0x7f
    "01111111", --  140 - 0x8c  :  127 - 0x7f
    "01111111", --  141 - 0x8d  :  127 - 0x7f
    "01111111", --  142 - 0x8e  :  127 - 0x7f
    "01111111", --  143 - 0x8f  :  127 - 0x7f
    "10101010", --  144 - 0x90  :  170 - 0xaa -- Background 0x9
    "11010101", --  145 - 0x91  :  213 - 0xd5
    "10101010", --  146 - 0x92  :  170 - 0xaa
    "11010101", --  147 - 0x93  :  213 - 0xd5
    "10101010", --  148 - 0x94  :  170 - 0xaa
    "11110101", --  149 - 0x95  :  245 - 0xf5
    "10101010", --  150 - 0x96  :  170 - 0xaa
    "11111111", --  151 - 0x97  :  255 - 0xff
    "01111111", --  152 - 0x98  :  127 - 0x7f -- plane 1
    "01111111", --  153 - 0x99  :  127 - 0x7f
    "01111111", --  154 - 0x9a  :  127 - 0x7f
    "01111111", --  155 - 0x9b  :  127 - 0x7f
    "01111111", --  156 - 0x9c  :  127 - 0x7f
    "01011111", --  157 - 0x9d  :   95 - 0x5f
    "01111111", --  158 - 0x9e  :  127 - 0x7f
    "00000000", --  159 - 0x9f  :    0 - 0x0
    "11111111", --  160 - 0xa0  :  255 - 0xff -- Background 0xa
    "01010101", --  161 - 0xa1  :   85 - 0x55
    "10101111", --  162 - 0xa2  :  175 - 0xaf
    "01010101", --  163 - 0xa3  :   85 - 0x55
    "10101011", --  164 - 0xa4  :  171 - 0xab
    "01010101", --  165 - 0xa5  :   85 - 0x55
    "10101011", --  166 - 0xa6  :  171 - 0xab
    "01010101", --  167 - 0xa7  :   85 - 0x55
    "00000000", --  168 - 0xa8  :    0 - 0x0 -- plane 1
    "11111110", --  169 - 0xa9  :  254 - 0xfe
    "11111010", --  170 - 0xaa  :  250 - 0xfa
    "11111110", --  171 - 0xab  :  254 - 0xfe
    "11111110", --  172 - 0xac  :  254 - 0xfe
    "11111110", --  173 - 0xad  :  254 - 0xfe
    "11111110", --  174 - 0xae  :  254 - 0xfe
    "11111110", --  175 - 0xaf  :  254 - 0xfe
    "10101011", --  176 - 0xb0  :  171 - 0xab -- Background 0xb
    "01010101", --  177 - 0xb1  :   85 - 0x55
    "10101011", --  178 - 0xb2  :  171 - 0xab
    "01010101", --  179 - 0xb3  :   85 - 0x55
    "10101011", --  180 - 0xb4  :  171 - 0xab
    "01010101", --  181 - 0xb5  :   85 - 0x55
    "10101011", --  182 - 0xb6  :  171 - 0xab
    "11111111", --  183 - 0xb7  :  255 - 0xff
    "11111110", --  184 - 0xb8  :  254 - 0xfe -- plane 1
    "11111110", --  185 - 0xb9  :  254 - 0xfe
    "11111110", --  186 - 0xba  :  254 - 0xfe
    "11111110", --  187 - 0xbb  :  254 - 0xfe
    "11111110", --  188 - 0xbc  :  254 - 0xfe
    "11111010", --  189 - 0xbd  :  250 - 0xfa
    "11111110", --  190 - 0xbe  :  254 - 0xfe
    "00000000", --  191 - 0xbf  :    0 - 0x0
    "11111111", --  192 - 0xc0  :  255 - 0xff -- Background 0xc
    "11010101", --  193 - 0xc1  :  213 - 0xd5
    "10100000", --  194 - 0xc2  :  160 - 0xa0
    "11010000", --  195 - 0xc3  :  208 - 0xd0
    "10001111", --  196 - 0xc4  :  143 - 0x8f
    "11001000", --  197 - 0xc5  :  200 - 0xc8
    "10001000", --  198 - 0xc6  :  136 - 0x88
    "11001000", --  199 - 0xc7  :  200 - 0xc8
    "00000000", --  200 - 0xc8  :    0 - 0x0 -- plane 1
    "00111111", --  201 - 0xc9  :   63 - 0x3f
    "01011111", --  202 - 0xca  :   95 - 0x5f
    "01101111", --  203 - 0xcb  :  111 - 0x6f
    "01110000", --  204 - 0xcc  :  112 - 0x70
    "01110111", --  205 - 0xcd  :  119 - 0x77
    "01110111", --  206 - 0xce  :  119 - 0x77
    "01110111", --  207 - 0xcf  :  119 - 0x77
    "10001000", --  208 - 0xd0  :  136 - 0x88 -- Background 0xd
    "11001000", --  209 - 0xd1  :  200 - 0xc8
    "10001000", --  210 - 0xd2  :  136 - 0x88
    "11001111", --  211 - 0xd3  :  207 - 0xcf
    "10010000", --  212 - 0xd4  :  144 - 0x90
    "11100000", --  213 - 0xd5  :  224 - 0xe0
    "11101010", --  214 - 0xd6  :  234 - 0xea
    "11111111", --  215 - 0xd7  :  255 - 0xff
    "01110111", --  216 - 0xd8  :  119 - 0x77 -- plane 1
    "01110111", --  217 - 0xd9  :  119 - 0x77
    "01110111", --  218 - 0xda  :  119 - 0x77
    "01110000", --  219 - 0xdb  :  112 - 0x70
    "01101111", --  220 - 0xdc  :  111 - 0x6f
    "01011111", --  221 - 0xdd  :   95 - 0x5f
    "00010101", --  222 - 0xde  :   21 - 0x15
    "00000000", --  223 - 0xdf  :    0 - 0x0
    "11111111", --  224 - 0xe0  :  255 - 0xff -- Background 0xe
    "01011011", --  225 - 0xe1  :   91 - 0x5b
    "00000111", --  226 - 0xe2  :    7 - 0x7
    "00001001", --  227 - 0xe3  :    9 - 0x9
    "11110011", --  228 - 0xe4  :  243 - 0xf3
    "00010001", --  229 - 0xe5  :   17 - 0x11
    "00010011", --  230 - 0xe6  :   19 - 0x13
    "00010001", --  231 - 0xe7  :   17 - 0x11
    "00000000", --  232 - 0xe8  :    0 - 0x0 -- plane 1
    "11111100", --  233 - 0xe9  :  252 - 0xfc
    "11111000", --  234 - 0xea  :  248 - 0xf8
    "11110110", --  235 - 0xeb  :  246 - 0xf6
    "00001100", --  236 - 0xec  :   12 - 0xc
    "11101110", --  237 - 0xed  :  238 - 0xee
    "11101100", --  238 - 0xee  :  236 - 0xec
    "11101110", --  239 - 0xef  :  238 - 0xee
    "00010011", --  240 - 0xf0  :   19 - 0x13 -- Background 0xf
    "00010001", --  241 - 0xf1  :   17 - 0x11
    "00010011", --  242 - 0xf2  :   19 - 0x13
    "11110001", --  243 - 0xf3  :  241 - 0xf1
    "00001011", --  244 - 0xf4  :   11 - 0xb
    "00000101", --  245 - 0xf5  :    5 - 0x5
    "10101011", --  246 - 0xf6  :  171 - 0xab
    "11111111", --  247 - 0xf7  :  255 - 0xff
    "11101100", --  248 - 0xf8  :  236 - 0xec -- plane 1
    "11101110", --  249 - 0xf9  :  238 - 0xee
    "11101100", --  250 - 0xfa  :  236 - 0xec
    "00001110", --  251 - 0xfb  :   14 - 0xe
    "11110100", --  252 - 0xfc  :  244 - 0xf4
    "11111010", --  253 - 0xfd  :  250 - 0xfa
    "01010100", --  254 - 0xfe  :   84 - 0x54
    "00000000", --  255 - 0xff  :    0 - 0x0
    "11010000", --  256 - 0x100  :  208 - 0xd0 -- Background 0x10
    "10010000", --  257 - 0x101  :  144 - 0x90
    "11011111", --  258 - 0x102  :  223 - 0xdf
    "10011010", --  259 - 0x103  :  154 - 0x9a
    "11010101", --  260 - 0x104  :  213 - 0xd5
    "10011111", --  261 - 0x105  :  159 - 0x9f
    "11010000", --  262 - 0x106  :  208 - 0xd0
    "10010000", --  263 - 0x107  :  144 - 0x90
    "01100000", --  264 - 0x108  :   96 - 0x60 -- plane 1
    "01100000", --  265 - 0x109  :   96 - 0x60
    "01100000", --  266 - 0x10a  :   96 - 0x60
    "01101111", --  267 - 0x10b  :  111 - 0x6f
    "01101010", --  268 - 0x10c  :  106 - 0x6a
    "01100000", --  269 - 0x10d  :   96 - 0x60
    "01100000", --  270 - 0x10e  :   96 - 0x60
    "01100000", --  271 - 0x10f  :   96 - 0x60
    "00001001", --  272 - 0x110  :    9 - 0x9 -- Background 0x11
    "00001011", --  273 - 0x111  :   11 - 0xb
    "11111001", --  274 - 0x112  :  249 - 0xf9
    "10101011", --  275 - 0x113  :  171 - 0xab
    "01011001", --  276 - 0x114  :   89 - 0x59
    "11111011", --  277 - 0x115  :  251 - 0xfb
    "00001001", --  278 - 0x116  :    9 - 0x9
    "00001011", --  279 - 0x117  :   11 - 0xb
    "00000110", --  280 - 0x118  :    6 - 0x6 -- plane 1
    "00000100", --  281 - 0x119  :    4 - 0x4
    "00000110", --  282 - 0x11a  :    6 - 0x6
    "11110100", --  283 - 0x11b  :  244 - 0xf4
    "10100110", --  284 - 0x11c  :  166 - 0xa6
    "00000100", --  285 - 0x11d  :    4 - 0x4
    "00000110", --  286 - 0x11e  :    6 - 0x6
    "00000100", --  287 - 0x11f  :    4 - 0x4
    "00011000", --  288 - 0x120  :   24 - 0x18 -- Background 0x12
    "00010100", --  289 - 0x121  :   20 - 0x14
    "00010100", --  290 - 0x122  :   20 - 0x14
    "00111010", --  291 - 0x123  :   58 - 0x3a
    "00111010", --  292 - 0x124  :   58 - 0x3a
    "01111010", --  293 - 0x125  :  122 - 0x7a
    "01111010", --  294 - 0x126  :  122 - 0x7a
    "01111010", --  295 - 0x127  :  122 - 0x7a
    "00000000", --  296 - 0x128  :    0 - 0x0 -- plane 1
    "00001000", --  297 - 0x129  :    8 - 0x8
    "00001000", --  298 - 0x12a  :    8 - 0x8
    "00011100", --  299 - 0x12b  :   28 - 0x1c
    "00011100", --  300 - 0x12c  :   28 - 0x1c
    "00111100", --  301 - 0x12d  :   60 - 0x3c
    "00111100", --  302 - 0x12e  :   60 - 0x3c
    "00111100", --  303 - 0x12f  :   60 - 0x3c
    "11111011", --  304 - 0x130  :  251 - 0xfb -- Background 0x13
    "11111101", --  305 - 0x131  :  253 - 0xfd
    "11111101", --  306 - 0x132  :  253 - 0xfd
    "11111101", --  307 - 0x133  :  253 - 0xfd
    "11111101", --  308 - 0x134  :  253 - 0xfd
    "11111101", --  309 - 0x135  :  253 - 0xfd
    "10000001", --  310 - 0x136  :  129 - 0x81
    "11111111", --  311 - 0x137  :  255 - 0xff
    "00111100", --  312 - 0x138  :   60 - 0x3c -- plane 1
    "01111110", --  313 - 0x139  :  126 - 0x7e
    "01111110", --  314 - 0x13a  :  126 - 0x7e
    "01111110", --  315 - 0x13b  :  126 - 0x7e
    "01111110", --  316 - 0x13c  :  126 - 0x7e
    "01111110", --  317 - 0x13d  :  126 - 0x7e
    "01111110", --  318 - 0x13e  :  126 - 0x7e
    "00000000", --  319 - 0x13f  :    0 - 0x0
    "00000000", --  320 - 0x140  :    0 - 0x0 -- Background 0x14
    "00000111", --  321 - 0x141  :    7 - 0x7
    "00000010", --  322 - 0x142  :    2 - 0x2
    "00000100", --  323 - 0x143  :    4 - 0x4
    "00000011", --  324 - 0x144  :    3 - 0x3
    "00000011", --  325 - 0x145  :    3 - 0x3
    "00001101", --  326 - 0x146  :   13 - 0xd
    "00010111", --  327 - 0x147  :   23 - 0x17
    "00000000", --  328 - 0x148  :    0 - 0x0 -- plane 1
    "00000000", --  329 - 0x149  :    0 - 0x0
    "00000101", --  330 - 0x14a  :    5 - 0x5
    "00000011", --  331 - 0x14b  :    3 - 0x3
    "00000000", --  332 - 0x14c  :    0 - 0x0
    "00000000", --  333 - 0x14d  :    0 - 0x0
    "00000010", --  334 - 0x14e  :    2 - 0x2
    "00001111", --  335 - 0x14f  :   15 - 0xf
    "00101111", --  336 - 0x150  :   47 - 0x2f -- Background 0x15
    "01001111", --  337 - 0x151  :   79 - 0x4f
    "01001111", --  338 - 0x152  :   79 - 0x4f
    "01001111", --  339 - 0x153  :   79 - 0x4f
    "01001111", --  340 - 0x154  :   79 - 0x4f
    "00100111", --  341 - 0x155  :   39 - 0x27
    "00010000", --  342 - 0x156  :   16 - 0x10
    "00001111", --  343 - 0x157  :   15 - 0xf
    "00011100", --  344 - 0x158  :   28 - 0x1c -- plane 1
    "00111010", --  345 - 0x159  :   58 - 0x3a
    "00111100", --  346 - 0x15a  :   60 - 0x3c
    "00111111", --  347 - 0x15b  :   63 - 0x3f
    "00111000", --  348 - 0x15c  :   56 - 0x38
    "00011110", --  349 - 0x15d  :   30 - 0x1e
    "00001111", --  350 - 0x15e  :   15 - 0xf
    "00000000", --  351 - 0x15f  :    0 - 0x0
    "00000000", --  352 - 0x160  :    0 - 0x0 -- Background 0x16
    "11100000", --  353 - 0x161  :  224 - 0xe0
    "10100000", --  354 - 0x162  :  160 - 0xa0
    "00100000", --  355 - 0x163  :   32 - 0x20
    "11000000", --  356 - 0x164  :  192 - 0xc0
    "01000000", --  357 - 0x165  :   64 - 0x40
    "00110000", --  358 - 0x166  :   48 - 0x30
    "11101000", --  359 - 0x167  :  232 - 0xe8
    "00000000", --  360 - 0x168  :    0 - 0x0 -- plane 1
    "00000000", --  361 - 0x169  :    0 - 0x0
    "01000000", --  362 - 0x16a  :   64 - 0x40
    "11000000", --  363 - 0x16b  :  192 - 0xc0
    "00000000", --  364 - 0x16c  :    0 - 0x0
    "10000000", --  365 - 0x16d  :  128 - 0x80
    "11000000", --  366 - 0x16e  :  192 - 0xc0
    "01110000", --  367 - 0x16f  :  112 - 0x70
    "11110100", --  368 - 0x170  :  244 - 0xf4 -- Background 0x17
    "11110010", --  369 - 0x171  :  242 - 0xf2
    "11110010", --  370 - 0x172  :  242 - 0xf2
    "11110010", --  371 - 0x173  :  242 - 0xf2
    "11110010", --  372 - 0x174  :  242 - 0xf2
    "11100100", --  373 - 0x175  :  228 - 0xe4
    "00001000", --  374 - 0x176  :    8 - 0x8
    "11110000", --  375 - 0x177  :  240 - 0xf0
    "00011000", --  376 - 0x178  :   24 - 0x18 -- plane 1
    "11111100", --  377 - 0x179  :  252 - 0xfc
    "00111100", --  378 - 0x17a  :   60 - 0x3c
    "01011100", --  379 - 0x17b  :   92 - 0x5c
    "00111100", --  380 - 0x17c  :   60 - 0x3c
    "11111000", --  381 - 0x17d  :  248 - 0xf8
    "11110000", --  382 - 0x17e  :  240 - 0xf0
    "00000000", --  383 - 0x17f  :    0 - 0x0
    "00111111", --  384 - 0x180  :   63 - 0x3f -- Background 0x18
    "01000000", --  385 - 0x181  :   64 - 0x40
    "01000000", --  386 - 0x182  :   64 - 0x40
    "10000000", --  387 - 0x183  :  128 - 0x80
    "10000000", --  388 - 0x184  :  128 - 0x80
    "01111111", --  389 - 0x185  :  127 - 0x7f
    "00000001", --  390 - 0x186  :    1 - 0x1
    "01111111", --  391 - 0x187  :  127 - 0x7f
    "00000000", --  392 - 0x188  :    0 - 0x0 -- plane 1
    "00111111", --  393 - 0x189  :   63 - 0x3f
    "00111111", --  394 - 0x18a  :   63 - 0x3f
    "01111111", --  395 - 0x18b  :  127 - 0x7f
    "01111111", --  396 - 0x18c  :  127 - 0x7f
    "00000000", --  397 - 0x18d  :    0 - 0x0
    "00000000", --  398 - 0x18e  :    0 - 0x0
    "00000000", --  399 - 0x18f  :    0 - 0x0
    "11111100", --  400 - 0x190  :  252 - 0xfc -- Background 0x19
    "00000010", --  401 - 0x191  :    2 - 0x2
    "00000010", --  402 - 0x192  :    2 - 0x2
    "00000001", --  403 - 0x193  :    1 - 0x1
    "00000001", --  404 - 0x194  :    1 - 0x1
    "11111110", --  405 - 0x195  :  254 - 0xfe
    "10000000", --  406 - 0x196  :  128 - 0x80
    "11111110", --  407 - 0x197  :  254 - 0xfe
    "00000000", --  408 - 0x198  :    0 - 0x0 -- plane 1
    "11111100", --  409 - 0x199  :  252 - 0xfc
    "11111100", --  410 - 0x19a  :  252 - 0xfc
    "11111110", --  411 - 0x19b  :  254 - 0xfe
    "11111110", --  412 - 0x19c  :  254 - 0xfe
    "00000000", --  413 - 0x19d  :    0 - 0x0
    "00000000", --  414 - 0x19e  :    0 - 0x0
    "00000000", --  415 - 0x19f  :    0 - 0x0
    "00000000", --  416 - 0x1a0  :    0 - 0x0 -- Background 0x1a
    "00000000", --  417 - 0x1a1  :    0 - 0x0
    "00111111", --  418 - 0x1a2  :   63 - 0x3f
    "01000000", --  419 - 0x1a3  :   64 - 0x40
    "01000000", --  420 - 0x1a4  :   64 - 0x40
    "10000000", --  421 - 0x1a5  :  128 - 0x80
    "10000000", --  422 - 0x1a6  :  128 - 0x80
    "01111111", --  423 - 0x1a7  :  127 - 0x7f
    "00000000", --  424 - 0x1a8  :    0 - 0x0 -- plane 1
    "00000000", --  425 - 0x1a9  :    0 - 0x0
    "00000000", --  426 - 0x1aa  :    0 - 0x0
    "00111111", --  427 - 0x1ab  :   63 - 0x3f
    "00111111", --  428 - 0x1ac  :   63 - 0x3f
    "01111111", --  429 - 0x1ad  :  127 - 0x7f
    "01111111", --  430 - 0x1ae  :  127 - 0x7f
    "00000000", --  431 - 0x1af  :    0 - 0x0
    "00000000", --  432 - 0x1b0  :    0 - 0x0 -- Background 0x1b
    "00000000", --  433 - 0x1b1  :    0 - 0x0
    "11111100", --  434 - 0x1b2  :  252 - 0xfc
    "00000010", --  435 - 0x1b3  :    2 - 0x2
    "00000010", --  436 - 0x1b4  :    2 - 0x2
    "00000001", --  437 - 0x1b5  :    1 - 0x1
    "00000001", --  438 - 0x1b6  :    1 - 0x1
    "11111110", --  439 - 0x1b7  :  254 - 0xfe
    "00000000", --  440 - 0x1b8  :    0 - 0x0 -- plane 1
    "00000000", --  441 - 0x1b9  :    0 - 0x0
    "00000000", --  442 - 0x1ba  :    0 - 0x0
    "11111100", --  443 - 0x1bb  :  252 - 0xfc
    "11111100", --  444 - 0x1bc  :  252 - 0xfc
    "11111110", --  445 - 0x1bd  :  254 - 0xfe
    "11111110", --  446 - 0x1be  :  254 - 0xfe
    "00000000", --  447 - 0x1bf  :    0 - 0x0
    "01111111", --  448 - 0x1c0  :  127 - 0x7f -- Background 0x1c
    "10000000", --  449 - 0x1c1  :  128 - 0x80
    "10000000", --  450 - 0x1c2  :  128 - 0x80
    "10000000", --  451 - 0x1c3  :  128 - 0x80
    "10011011", --  452 - 0x1c4  :  155 - 0x9b
    "10100100", --  453 - 0x1c5  :  164 - 0xa4
    "10100110", --  454 - 0x1c6  :  166 - 0xa6
    "10000000", --  455 - 0x1c7  :  128 - 0x80
    "00000000", --  456 - 0x1c8  :    0 - 0x0 -- plane 1
    "01111111", --  457 - 0x1c9  :  127 - 0x7f
    "01111111", --  458 - 0x1ca  :  127 - 0x7f
    "01111111", --  459 - 0x1cb  :  127 - 0x7f
    "01100100", --  460 - 0x1cc  :  100 - 0x64
    "01011011", --  461 - 0x1cd  :   91 - 0x5b
    "01011001", --  462 - 0x1ce  :   89 - 0x59
    "01111111", --  463 - 0x1cf  :  127 - 0x7f
    "10000000", --  464 - 0x1d0  :  128 - 0x80 -- Background 0x1d
    "01111111", --  465 - 0x1d1  :  127 - 0x7f
    "00000010", --  466 - 0x1d2  :    2 - 0x2
    "00000010", --  467 - 0x1d3  :    2 - 0x2
    "00000010", --  468 - 0x1d4  :    2 - 0x2
    "00000010", --  469 - 0x1d5  :    2 - 0x2
    "00000010", --  470 - 0x1d6  :    2 - 0x2
    "00001111", --  471 - 0x1d7  :   15 - 0xf
    "01111111", --  472 - 0x1d8  :  127 - 0x7f -- plane 1
    "00000000", --  473 - 0x1d9  :    0 - 0x0
    "00000001", --  474 - 0x1da  :    1 - 0x1
    "00000001", --  475 - 0x1db  :    1 - 0x1
    "00000001", --  476 - 0x1dc  :    1 - 0x1
    "00000001", --  477 - 0x1dd  :    1 - 0x1
    "00000001", --  478 - 0x1de  :    1 - 0x1
    "00000000", --  479 - 0x1df  :    0 - 0x0
    "11111110", --  480 - 0x1e0  :  254 - 0xfe -- Background 0x1e
    "00000001", --  481 - 0x1e1  :    1 - 0x1
    "00000001", --  482 - 0x1e2  :    1 - 0x1
    "00000001", --  483 - 0x1e3  :    1 - 0x1
    "01000001", --  484 - 0x1e4  :   65 - 0x41
    "11110101", --  485 - 0x1e5  :  245 - 0xf5
    "00011101", --  486 - 0x1e6  :   29 - 0x1d
    "00000001", --  487 - 0x1e7  :    1 - 0x1
    "00000000", --  488 - 0x1e8  :    0 - 0x0 -- plane 1
    "11111110", --  489 - 0x1e9  :  254 - 0xfe
    "11111110", --  490 - 0x1ea  :  254 - 0xfe
    "11111110", --  491 - 0x1eb  :  254 - 0xfe
    "10111110", --  492 - 0x1ec  :  190 - 0xbe
    "00001010", --  493 - 0x1ed  :   10 - 0xa
    "11100010", --  494 - 0x1ee  :  226 - 0xe2
    "11111110", --  495 - 0x1ef  :  254 - 0xfe
    "00000001", --  496 - 0x1f0  :    1 - 0x1 -- Background 0x1f
    "11111110", --  497 - 0x1f1  :  254 - 0xfe
    "01000000", --  498 - 0x1f2  :   64 - 0x40
    "01000000", --  499 - 0x1f3  :   64 - 0x40
    "01000000", --  500 - 0x1f4  :   64 - 0x40
    "01000000", --  501 - 0x1f5  :   64 - 0x40
    "01000000", --  502 - 0x1f6  :   64 - 0x40
    "11110000", --  503 - 0x1f7  :  240 - 0xf0
    "11111110", --  504 - 0x1f8  :  254 - 0xfe -- plane 1
    "00000000", --  505 - 0x1f9  :    0 - 0x0
    "10000000", --  506 - 0x1fa  :  128 - 0x80
    "10000000", --  507 - 0x1fb  :  128 - 0x80
    "10000000", --  508 - 0x1fc  :  128 - 0x80
    "10000000", --  509 - 0x1fd  :  128 - 0x80
    "10000000", --  510 - 0x1fe  :  128 - 0x80
    "00000000", --  511 - 0x1ff  :    0 - 0x0
    "00000111", --  512 - 0x200  :    7 - 0x7 -- Background 0x20
    "00011111", --  513 - 0x201  :   31 - 0x1f
    "00111111", --  514 - 0x202  :   63 - 0x3f
    "01111111", --  515 - 0x203  :  127 - 0x7f
    "01111111", --  516 - 0x204  :  127 - 0x7f
    "11111111", --  517 - 0x205  :  255 - 0xff
    "11111111", --  518 - 0x206  :  255 - 0xff
    "11111111", --  519 - 0x207  :  255 - 0xff
    "00000000", --  520 - 0x208  :    0 - 0x0 -- plane 1
    "00000000", --  521 - 0x209  :    0 - 0x0
    "00000000", --  522 - 0x20a  :    0 - 0x0
    "00000000", --  523 - 0x20b  :    0 - 0x0
    "00000000", --  524 - 0x20c  :    0 - 0x0
    "00000000", --  525 - 0x20d  :    0 - 0x0
    "00000000", --  526 - 0x20e  :    0 - 0x0
    "00000000", --  527 - 0x20f  :    0 - 0x0
    "11100000", --  528 - 0x210  :  224 - 0xe0 -- Background 0x21
    "11111000", --  529 - 0x211  :  248 - 0xf8
    "11111100", --  530 - 0x212  :  252 - 0xfc
    "11111110", --  531 - 0x213  :  254 - 0xfe
    "11111110", --  532 - 0x214  :  254 - 0xfe
    "11111111", --  533 - 0x215  :  255 - 0xff
    "11111111", --  534 - 0x216  :  255 - 0xff
    "11111111", --  535 - 0x217  :  255 - 0xff
    "00000000", --  536 - 0x218  :    0 - 0x0 -- plane 1
    "00000000", --  537 - 0x219  :    0 - 0x0
    "00000000", --  538 - 0x21a  :    0 - 0x0
    "00000000", --  539 - 0x21b  :    0 - 0x0
    "00000000", --  540 - 0x21c  :    0 - 0x0
    "00000000", --  541 - 0x21d  :    0 - 0x0
    "00000000", --  542 - 0x21e  :    0 - 0x0
    "00000000", --  543 - 0x21f  :    0 - 0x0
    "00000111", --  544 - 0x220  :    7 - 0x7 -- Background 0x22
    "00011111", --  545 - 0x221  :   31 - 0x1f
    "00111111", --  546 - 0x222  :   63 - 0x3f
    "01111111", --  547 - 0x223  :  127 - 0x7f
    "01111111", --  548 - 0x224  :  127 - 0x7f
    "11111111", --  549 - 0x225  :  255 - 0xff
    "11111111", --  550 - 0x226  :  255 - 0xff
    "11111111", --  551 - 0x227  :  255 - 0xff
    "00000000", --  552 - 0x228  :    0 - 0x0 -- plane 1
    "00000000", --  553 - 0x229  :    0 - 0x0
    "00011000", --  554 - 0x22a  :   24 - 0x18
    "00010000", --  555 - 0x22b  :   16 - 0x10
    "00011010", --  556 - 0x22c  :   26 - 0x1a
    "00010001", --  557 - 0x22d  :   17 - 0x11
    "00011010", --  558 - 0x22e  :   26 - 0x1a
    "00000000", --  559 - 0x22f  :    0 - 0x0
    "11100000", --  560 - 0x230  :  224 - 0xe0 -- Background 0x23
    "11111000", --  561 - 0x231  :  248 - 0xf8
    "11111100", --  562 - 0x232  :  252 - 0xfc
    "11111110", --  563 - 0x233  :  254 - 0xfe
    "11111110", --  564 - 0x234  :  254 - 0xfe
    "11111111", --  565 - 0x235  :  255 - 0xff
    "11111111", --  566 - 0x236  :  255 - 0xff
    "11111111", --  567 - 0x237  :  255 - 0xff
    "00000000", --  568 - 0x238  :    0 - 0x0 -- plane 1
    "00000000", --  569 - 0x239  :    0 - 0x0
    "00000000", --  570 - 0x23a  :    0 - 0x0
    "00101000", --  571 - 0x23b  :   40 - 0x28
    "10001100", --  572 - 0x23c  :  140 - 0x8c
    "00101000", --  573 - 0x23d  :   40 - 0x28
    "10101100", --  574 - 0x23e  :  172 - 0xac
    "00000000", --  575 - 0x23f  :    0 - 0x0
    "00000000", --  576 - 0x240  :    0 - 0x0 -- Background 0x24
    "00000000", --  577 - 0x241  :    0 - 0x0
    "00000000", --  578 - 0x242  :    0 - 0x0
    "00000000", --  579 - 0x243  :    0 - 0x0
    "00000000", --  580 - 0x244  :    0 - 0x0
    "00000000", --  581 - 0x245  :    0 - 0x0
    "00000000", --  582 - 0x246  :    0 - 0x0
    "00000000", --  583 - 0x247  :    0 - 0x0
    "00000000", --  584 - 0x248  :    0 - 0x0 -- plane 1
    "00000000", --  585 - 0x249  :    0 - 0x0
    "00000000", --  586 - 0x24a  :    0 - 0x0
    "00000000", --  587 - 0x24b  :    0 - 0x0
    "00000000", --  588 - 0x24c  :    0 - 0x0
    "00000000", --  589 - 0x24d  :    0 - 0x0
    "00000000", --  590 - 0x24e  :    0 - 0x0
    "00000000", --  591 - 0x24f  :    0 - 0x0
    "00101111", --  592 - 0x250  :   47 - 0x2f -- Background 0x25
    "01001111", --  593 - 0x251  :   79 - 0x4f
    "01001111", --  594 - 0x252  :   79 - 0x4f
    "01001111", --  595 - 0x253  :   79 - 0x4f
    "01001111", --  596 - 0x254  :   79 - 0x4f
    "00100111", --  597 - 0x255  :   39 - 0x27
    "00010000", --  598 - 0x256  :   16 - 0x10
    "00001111", --  599 - 0x257  :   15 - 0xf
    "00011100", --  600 - 0x258  :   28 - 0x1c -- plane 1
    "00111001", --  601 - 0x259  :   57 - 0x39
    "00111111", --  602 - 0x25a  :   63 - 0x3f
    "00111110", --  603 - 0x25b  :   62 - 0x3e
    "00111111", --  604 - 0x25c  :   63 - 0x3f
    "00011110", --  605 - 0x25d  :   30 - 0x1e
    "00001111", --  606 - 0x25e  :   15 - 0xf
    "00000000", --  607 - 0x25f  :    0 - 0x0
    "00000000", --  608 - 0x260  :    0 - 0x0 -- Background 0x26
    "11100000", --  609 - 0x261  :  224 - 0xe0
    "10100000", --  610 - 0x262  :  160 - 0xa0
    "00100000", --  611 - 0x263  :   32 - 0x20
    "11000000", --  612 - 0x264  :  192 - 0xc0
    "01000000", --  613 - 0x265  :   64 - 0x40
    "00110000", --  614 - 0x266  :   48 - 0x30
    "11101000", --  615 - 0x267  :  232 - 0xe8
    "00000000", --  616 - 0x268  :    0 - 0x0 -- plane 1
    "00000000", --  617 - 0x269  :    0 - 0x0
    "01000000", --  618 - 0x26a  :   64 - 0x40
    "11000000", --  619 - 0x26b  :  192 - 0xc0
    "00000000", --  620 - 0x26c  :    0 - 0x0
    "10000000", --  621 - 0x26d  :  128 - 0x80
    "11000000", --  622 - 0x26e  :  192 - 0xc0
    "11110000", --  623 - 0x26f  :  240 - 0xf0
    "11110100", --  624 - 0x270  :  244 - 0xf4 -- Background 0x27
    "11110010", --  625 - 0x271  :  242 - 0xf2
    "11110010", --  626 - 0x272  :  242 - 0xf2
    "11110010", --  627 - 0x273  :  242 - 0xf2
    "11110010", --  628 - 0x274  :  242 - 0xf2
    "11100100", --  629 - 0x275  :  228 - 0xe4
    "00001000", --  630 - 0x276  :    8 - 0x8
    "11110000", --  631 - 0x277  :  240 - 0xf0
    "00111000", --  632 - 0x278  :   56 - 0x38 -- plane 1
    "10011100", --  633 - 0x279  :  156 - 0x9c
    "10011100", --  634 - 0x27a  :  156 - 0x9c
    "00111100", --  635 - 0x27b  :   60 - 0x3c
    "11111100", --  636 - 0x27c  :  252 - 0xfc
    "01111000", --  637 - 0x27d  :  120 - 0x78
    "11110000", --  638 - 0x27e  :  240 - 0xf0
    "00000000", --  639 - 0x27f  :    0 - 0x0
    "11111111", --  640 - 0x280  :  255 - 0xff -- Background 0x28
    "11010101", --  641 - 0x281  :  213 - 0xd5
    "10100011", --  642 - 0x282  :  163 - 0xa3
    "11010111", --  643 - 0x283  :  215 - 0xd7
    "10001111", --  644 - 0x284  :  143 - 0x8f
    "11001111", --  645 - 0x285  :  207 - 0xcf
    "10001011", --  646 - 0x286  :  139 - 0x8b
    "11001011", --  647 - 0x287  :  203 - 0xcb
    "00000000", --  648 - 0x288  :    0 - 0x0 -- plane 1
    "00111110", --  649 - 0x289  :   62 - 0x3e
    "01011101", --  650 - 0x28a  :   93 - 0x5d
    "01101011", --  651 - 0x28b  :  107 - 0x6b
    "01110101", --  652 - 0x28c  :  117 - 0x75
    "01110001", --  653 - 0x28d  :  113 - 0x71
    "01110101", --  654 - 0x28e  :  117 - 0x75
    "01110100", --  655 - 0x28f  :  116 - 0x74
    "10001111", --  656 - 0x290  :  143 - 0x8f -- Background 0x29
    "11001111", --  657 - 0x291  :  207 - 0xcf
    "10001111", --  658 - 0x292  :  143 - 0x8f
    "11001111", --  659 - 0x293  :  207 - 0xcf
    "10010000", --  660 - 0x294  :  144 - 0x90
    "11100000", --  661 - 0x295  :  224 - 0xe0
    "11101010", --  662 - 0x296  :  234 - 0xea
    "11111111", --  663 - 0x297  :  255 - 0xff
    "01110000", --  664 - 0x298  :  112 - 0x70 -- plane 1
    "01110111", --  665 - 0x299  :  119 - 0x77
    "01110111", --  666 - 0x29a  :  119 - 0x77
    "01110000", --  667 - 0x29b  :  112 - 0x70
    "01101111", --  668 - 0x29c  :  111 - 0x6f
    "01011111", --  669 - 0x29d  :   95 - 0x5f
    "00010101", --  670 - 0x29e  :   21 - 0x15
    "00000000", --  671 - 0x29f  :    0 - 0x0
    "11111111", --  672 - 0x2a0  :  255 - 0xff -- Background 0x2a
    "11011011", --  673 - 0x2a1  :  219 - 0xdb
    "11000111", --  674 - 0x2a2  :  199 - 0xc7
    "11101001", --  675 - 0x2a3  :  233 - 0xe9
    "11110011", --  676 - 0x2a4  :  243 - 0xf3
    "11110001", --  677 - 0x2a5  :  241 - 0xf1
    "11010011", --  678 - 0x2a6  :  211 - 0xd3
    "11010001", --  679 - 0x2a7  :  209 - 0xd1
    "00000000", --  680 - 0x2a8  :    0 - 0x0 -- plane 1
    "01111100", --  681 - 0x2a9  :  124 - 0x7c
    "10111000", --  682 - 0x2aa  :  184 - 0xb8
    "11010110", --  683 - 0x2ab  :  214 - 0xd6
    "10101100", --  684 - 0x2ac  :  172 - 0xac
    "10001110", --  685 - 0x2ad  :  142 - 0x8e
    "10101100", --  686 - 0x2ae  :  172 - 0xac
    "00101110", --  687 - 0x2af  :   46 - 0x2e
    "11110011", --  688 - 0x2b0  :  243 - 0xf3 -- Background 0x2b
    "11110001", --  689 - 0x2b1  :  241 - 0xf1
    "11110011", --  690 - 0x2b2  :  243 - 0xf3
    "11110001", --  691 - 0x2b3  :  241 - 0xf1
    "00001011", --  692 - 0x2b4  :   11 - 0xb
    "00000101", --  693 - 0x2b5  :    5 - 0x5
    "10101011", --  694 - 0x2b6  :  171 - 0xab
    "11111111", --  695 - 0x2b7  :  255 - 0xff
    "00001100", --  696 - 0x2b8  :   12 - 0xc -- plane 1
    "11101110", --  697 - 0x2b9  :  238 - 0xee
    "11101100", --  698 - 0x2ba  :  236 - 0xec
    "00001110", --  699 - 0x2bb  :   14 - 0xe
    "11110100", --  700 - 0x2bc  :  244 - 0xf4
    "11111010", --  701 - 0x2bd  :  250 - 0xfa
    "01010100", --  702 - 0x2be  :   84 - 0x54
    "00000000", --  703 - 0x2bf  :    0 - 0x0
    "00000000", --  704 - 0x2c0  :    0 - 0x0 -- Background 0x2c
    "00000000", --  705 - 0x2c1  :    0 - 0x0
    "00000000", --  706 - 0x2c2  :    0 - 0x0
    "00000000", --  707 - 0x2c3  :    0 - 0x0
    "00000000", --  708 - 0x2c4  :    0 - 0x0
    "00000000", --  709 - 0x2c5  :    0 - 0x0
    "00000000", --  710 - 0x2c6  :    0 - 0x0
    "00000000", --  711 - 0x2c7  :    0 - 0x0
    "00000000", --  712 - 0x2c8  :    0 - 0x0 -- plane 1
    "00000000", --  713 - 0x2c9  :    0 - 0x0
    "00000000", --  714 - 0x2ca  :    0 - 0x0
    "00000000", --  715 - 0x2cb  :    0 - 0x0
    "00000000", --  716 - 0x2cc  :    0 - 0x0
    "00000000", --  717 - 0x2cd  :    0 - 0x0
    "00000000", --  718 - 0x2ce  :    0 - 0x0
    "00000000", --  719 - 0x2cf  :    0 - 0x0
    "00101111", --  720 - 0x2d0  :   47 - 0x2f -- Background 0x2d
    "01001111", --  721 - 0x2d1  :   79 - 0x4f
    "01001111", --  722 - 0x2d2  :   79 - 0x4f
    "01001111", --  723 - 0x2d3  :   79 - 0x4f
    "01001111", --  724 - 0x2d4  :   79 - 0x4f
    "00100111", --  725 - 0x2d5  :   39 - 0x27
    "00010000", --  726 - 0x2d6  :   16 - 0x10
    "00001111", --  727 - 0x2d7  :   15 - 0xf
    "00011110", --  728 - 0x2d8  :   30 - 0x1e -- plane 1
    "00111110", --  729 - 0x2d9  :   62 - 0x3e
    "00111110", --  730 - 0x2da  :   62 - 0x3e
    "00111110", --  731 - 0x2db  :   62 - 0x3e
    "00111111", --  732 - 0x2dc  :   63 - 0x3f
    "00011110", --  733 - 0x2dd  :   30 - 0x1e
    "00001111", --  734 - 0x2de  :   15 - 0xf
    "00000000", --  735 - 0x2df  :    0 - 0x0
    "00000000", --  736 - 0x2e0  :    0 - 0x0 -- Background 0x2e
    "00000000", --  737 - 0x2e1  :    0 - 0x0
    "00000000", --  738 - 0x2e2  :    0 - 0x0
    "00000000", --  739 - 0x2e3  :    0 - 0x0
    "00000000", --  740 - 0x2e4  :    0 - 0x0
    "00000000", --  741 - 0x2e5  :    0 - 0x0
    "00000000", --  742 - 0x2e6  :    0 - 0x0
    "00000000", --  743 - 0x2e7  :    0 - 0x0
    "00000000", --  744 - 0x2e8  :    0 - 0x0 -- plane 1
    "00000000", --  745 - 0x2e9  :    0 - 0x0
    "00000000", --  746 - 0x2ea  :    0 - 0x0
    "00000000", --  747 - 0x2eb  :    0 - 0x0
    "00000000", --  748 - 0x2ec  :    0 - 0x0
    "00000000", --  749 - 0x2ed  :    0 - 0x0
    "00000000", --  750 - 0x2ee  :    0 - 0x0
    "00000000", --  751 - 0x2ef  :    0 - 0x0
    "11110100", --  752 - 0x2f0  :  244 - 0xf4 -- Background 0x2f
    "11110010", --  753 - 0x2f1  :  242 - 0xf2
    "11110010", --  754 - 0x2f2  :  242 - 0xf2
    "11110010", --  755 - 0x2f3  :  242 - 0xf2
    "11110010", --  756 - 0x2f4  :  242 - 0xf2
    "11100100", --  757 - 0x2f5  :  228 - 0xe4
    "00001000", --  758 - 0x2f6  :    8 - 0x8
    "11110000", --  759 - 0x2f7  :  240 - 0xf0
    "01111000", --  760 - 0x2f8  :  120 - 0x78 -- plane 1
    "01111100", --  761 - 0x2f9  :  124 - 0x7c
    "01111100", --  762 - 0x2fa  :  124 - 0x7c
    "01111100", --  763 - 0x2fb  :  124 - 0x7c
    "11111100", --  764 - 0x2fc  :  252 - 0xfc
    "01111000", --  765 - 0x2fd  :  120 - 0x78
    "11110000", --  766 - 0x2fe  :  240 - 0xf0
    "00000000", --  767 - 0x2ff  :    0 - 0x0
    "00011000", --  768 - 0x300  :   24 - 0x18 -- Background 0x30
    "00100100", --  769 - 0x301  :   36 - 0x24
    "01000010", --  770 - 0x302  :   66 - 0x42
    "10100101", --  771 - 0x303  :  165 - 0xa5
    "11100111", --  772 - 0x304  :  231 - 0xe7
    "00100100", --  773 - 0x305  :   36 - 0x24
    "00100100", --  774 - 0x306  :   36 - 0x24
    "00111100", --  775 - 0x307  :   60 - 0x3c
    "00000000", --  776 - 0x308  :    0 - 0x0 -- plane 1
    "00011000", --  777 - 0x309  :   24 - 0x18
    "00111100", --  778 - 0x30a  :   60 - 0x3c
    "01011010", --  779 - 0x30b  :   90 - 0x5a
    "00011000", --  780 - 0x30c  :   24 - 0x18
    "00011000", --  781 - 0x30d  :   24 - 0x18
    "00011000", --  782 - 0x30e  :   24 - 0x18
    "00000000", --  783 - 0x30f  :    0 - 0x0
    "00111100", --  784 - 0x310  :   60 - 0x3c -- Background 0x31
    "00100100", --  785 - 0x311  :   36 - 0x24
    "00100100", --  786 - 0x312  :   36 - 0x24
    "01100110", --  787 - 0x313  :  102 - 0x66
    "10100101", --  788 - 0x314  :  165 - 0xa5
    "01000010", --  789 - 0x315  :   66 - 0x42
    "00100100", --  790 - 0x316  :   36 - 0x24
    "00011000", --  791 - 0x317  :   24 - 0x18
    "00000000", --  792 - 0x318  :    0 - 0x0 -- plane 1
    "00011000", --  793 - 0x319  :   24 - 0x18
    "00011000", --  794 - 0x31a  :   24 - 0x18
    "00011000", --  795 - 0x31b  :   24 - 0x18
    "01011010", --  796 - 0x31c  :   90 - 0x5a
    "00111100", --  797 - 0x31d  :   60 - 0x3c
    "00011000", --  798 - 0x31e  :   24 - 0x18
    "00000000", --  799 - 0x31f  :    0 - 0x0
    "00000010", --  800 - 0x320  :    2 - 0x2 -- Background 0x32
    "00000010", --  801 - 0x321  :    2 - 0x2
    "00000011", --  802 - 0x322  :    3 - 0x3
    "00000010", --  803 - 0x323  :    2 - 0x2
    "00000010", --  804 - 0x324  :    2 - 0x2
    "00000010", --  805 - 0x325  :    2 - 0x2
    "00000011", --  806 - 0x326  :    3 - 0x3
    "00000010", --  807 - 0x327  :    2 - 0x2
    "00000001", --  808 - 0x328  :    1 - 0x1 -- plane 1
    "00000001", --  809 - 0x329  :    1 - 0x1
    "00000000", --  810 - 0x32a  :    0 - 0x0
    "00000001", --  811 - 0x32b  :    1 - 0x1
    "00000001", --  812 - 0x32c  :    1 - 0x1
    "00000001", --  813 - 0x32d  :    1 - 0x1
    "00000000", --  814 - 0x32e  :    0 - 0x0
    "00000001", --  815 - 0x32f  :    1 - 0x1
    "01000000", --  816 - 0x330  :   64 - 0x40 -- Background 0x33
    "11000000", --  817 - 0x331  :  192 - 0xc0
    "01000000", --  818 - 0x332  :   64 - 0x40
    "01000000", --  819 - 0x333  :   64 - 0x40
    "01000000", --  820 - 0x334  :   64 - 0x40
    "11000000", --  821 - 0x335  :  192 - 0xc0
    "01000000", --  822 - 0x336  :   64 - 0x40
    "01000000", --  823 - 0x337  :   64 - 0x40
    "10000000", --  824 - 0x338  :  128 - 0x80 -- plane 1
    "00000000", --  825 - 0x339  :    0 - 0x0
    "10000000", --  826 - 0x33a  :  128 - 0x80
    "10000000", --  827 - 0x33b  :  128 - 0x80
    "10000000", --  828 - 0x33c  :  128 - 0x80
    "00000000", --  829 - 0x33d  :    0 - 0x0
    "10000000", --  830 - 0x33e  :  128 - 0x80
    "10000000", --  831 - 0x33f  :  128 - 0x80
    "00000000", --  832 - 0x340  :    0 - 0x0 -- Background 0x34
    "00011000", --  833 - 0x341  :   24 - 0x18
    "00111100", --  834 - 0x342  :   60 - 0x3c
    "01100010", --  835 - 0x343  :   98 - 0x62
    "01100001", --  836 - 0x344  :   97 - 0x61
    "11000000", --  837 - 0x345  :  192 - 0xc0
    "11000000", --  838 - 0x346  :  192 - 0xc0
    "11000000", --  839 - 0x347  :  192 - 0xc0
    "00000000", --  840 - 0x348  :    0 - 0x0 -- plane 1
    "00000000", --  841 - 0x349  :    0 - 0x0
    "00011000", --  842 - 0x34a  :   24 - 0x18
    "00111100", --  843 - 0x34b  :   60 - 0x3c
    "00111110", --  844 - 0x34c  :   62 - 0x3e
    "01111111", --  845 - 0x34d  :  127 - 0x7f
    "01111111", --  846 - 0x34e  :  127 - 0x7f
    "01111111", --  847 - 0x34f  :  127 - 0x7f
    "01100000", --  848 - 0x350  :   96 - 0x60 -- Background 0x35
    "01100000", --  849 - 0x351  :   96 - 0x60
    "00110000", --  850 - 0x352  :   48 - 0x30
    "00011000", --  851 - 0x353  :   24 - 0x18
    "00001100", --  852 - 0x354  :   12 - 0xc
    "00000110", --  853 - 0x355  :    6 - 0x6
    "00000010", --  854 - 0x356  :    2 - 0x2
    "00000001", --  855 - 0x357  :    1 - 0x1
    "00111111", --  856 - 0x358  :   63 - 0x3f -- plane 1
    "00111111", --  857 - 0x359  :   63 - 0x3f
    "00011111", --  858 - 0x35a  :   31 - 0x1f
    "00001111", --  859 - 0x35b  :   15 - 0xf
    "00000111", --  860 - 0x35c  :    7 - 0x7
    "00000011", --  861 - 0x35d  :    3 - 0x3
    "00000001", --  862 - 0x35e  :    1 - 0x1
    "00000000", --  863 - 0x35f  :    0 - 0x0
    "00000000", --  864 - 0x360  :    0 - 0x0 -- Background 0x36
    "00011000", --  865 - 0x361  :   24 - 0x18
    "00100100", --  866 - 0x362  :   36 - 0x24
    "01000010", --  867 - 0x363  :   66 - 0x42
    "10000010", --  868 - 0x364  :  130 - 0x82
    "00000001", --  869 - 0x365  :    1 - 0x1
    "00000001", --  870 - 0x366  :    1 - 0x1
    "00000001", --  871 - 0x367  :    1 - 0x1
    "00000000", --  872 - 0x368  :    0 - 0x0 -- plane 1
    "00000000", --  873 - 0x369  :    0 - 0x0
    "00011000", --  874 - 0x36a  :   24 - 0x18
    "00111100", --  875 - 0x36b  :   60 - 0x3c
    "01111100", --  876 - 0x36c  :  124 - 0x7c
    "11111110", --  877 - 0x36d  :  254 - 0xfe
    "11111110", --  878 - 0x36e  :  254 - 0xfe
    "11111110", --  879 - 0x36f  :  254 - 0xfe
    "00000010", --  880 - 0x370  :    2 - 0x2 -- Background 0x37
    "00000010", --  881 - 0x371  :    2 - 0x2
    "00000100", --  882 - 0x372  :    4 - 0x4
    "00001000", --  883 - 0x373  :    8 - 0x8
    "00010000", --  884 - 0x374  :   16 - 0x10
    "00100000", --  885 - 0x375  :   32 - 0x20
    "01000000", --  886 - 0x376  :   64 - 0x40
    "10000000", --  887 - 0x377  :  128 - 0x80
    "11111100", --  888 - 0x378  :  252 - 0xfc -- plane 1
    "11111100", --  889 - 0x379  :  252 - 0xfc
    "11111000", --  890 - 0x37a  :  248 - 0xf8
    "11110000", --  891 - 0x37b  :  240 - 0xf0
    "11100000", --  892 - 0x37c  :  224 - 0xe0
    "11000000", --  893 - 0x37d  :  192 - 0xc0
    "10000000", --  894 - 0x37e  :  128 - 0x80
    "00000000", --  895 - 0x37f  :    0 - 0x0
    "00000000", --  896 - 0x380  :    0 - 0x0 -- Background 0x38
    "00000110", --  897 - 0x381  :    6 - 0x6
    "00001101", --  898 - 0x382  :   13 - 0xd
    "00001100", --  899 - 0x383  :   12 - 0xc
    "00001100", --  900 - 0x384  :   12 - 0xc
    "00000110", --  901 - 0x385  :    6 - 0x6
    "00000010", --  902 - 0x386  :    2 - 0x2
    "00000001", --  903 - 0x387  :    1 - 0x1
    "00000000", --  904 - 0x388  :    0 - 0x0 -- plane 1
    "00000000", --  905 - 0x389  :    0 - 0x0
    "00000110", --  906 - 0x38a  :    6 - 0x6
    "00000111", --  907 - 0x38b  :    7 - 0x7
    "00000111", --  908 - 0x38c  :    7 - 0x7
    "00000011", --  909 - 0x38d  :    3 - 0x3
    "00000001", --  910 - 0x38e  :    1 - 0x1
    "00000000", --  911 - 0x38f  :    0 - 0x0
    "11111111", --  912 - 0x390  :  255 - 0xff -- Background 0x39
    "00000000", --  913 - 0x391  :    0 - 0x0
    "00000000", --  914 - 0x392  :    0 - 0x0
    "00000000", --  915 - 0x393  :    0 - 0x0
    "00000000", --  916 - 0x394  :    0 - 0x0
    "00000000", --  917 - 0x395  :    0 - 0x0
    "00000000", --  918 - 0x396  :    0 - 0x0
    "00000000", --  919 - 0x397  :    0 - 0x0
    "00000000", --  920 - 0x398  :    0 - 0x0 -- plane 1
    "00000000", --  921 - 0x399  :    0 - 0x0
    "00000000", --  922 - 0x39a  :    0 - 0x0
    "00000000", --  923 - 0x39b  :    0 - 0x0
    "00000000", --  924 - 0x39c  :    0 - 0x0
    "00000000", --  925 - 0x39d  :    0 - 0x0
    "00000000", --  926 - 0x39e  :    0 - 0x0
    "00000000", --  927 - 0x39f  :    0 - 0x0
    "00000000", --  928 - 0x3a0  :    0 - 0x0 -- Background 0x3a
    "01100000", --  929 - 0x3a1  :   96 - 0x60
    "10010000", --  930 - 0x3a2  :  144 - 0x90
    "00010000", --  931 - 0x3a3  :   16 - 0x10
    "00010000", --  932 - 0x3a4  :   16 - 0x10
    "00100000", --  933 - 0x3a5  :   32 - 0x20
    "01000000", --  934 - 0x3a6  :   64 - 0x40
    "10000000", --  935 - 0x3a7  :  128 - 0x80
    "00000000", --  936 - 0x3a8  :    0 - 0x0 -- plane 1
    "00000000", --  937 - 0x3a9  :    0 - 0x0
    "01100000", --  938 - 0x3aa  :   96 - 0x60
    "11100000", --  939 - 0x3ab  :  224 - 0xe0
    "11100000", --  940 - 0x3ac  :  224 - 0xe0
    "11000000", --  941 - 0x3ad  :  192 - 0xc0
    "10000000", --  942 - 0x3ae  :  128 - 0x80
    "00000000", --  943 - 0x3af  :    0 - 0x0
    "00000000", --  944 - 0x3b0  :    0 - 0x0 -- Background 0x3b
    "01010100", --  945 - 0x3b1  :   84 - 0x54
    "00000010", --  946 - 0x3b2  :    2 - 0x2
    "01000000", --  947 - 0x3b3  :   64 - 0x40
    "00000010", --  948 - 0x3b4  :    2 - 0x2
    "01000000", --  949 - 0x3b5  :   64 - 0x40
    "00101010", --  950 - 0x3b6  :   42 - 0x2a
    "00000000", --  951 - 0x3b7  :    0 - 0x0
    "00000000", --  952 - 0x3b8  :    0 - 0x0 -- plane 1
    "00101010", --  953 - 0x3b9  :   42 - 0x2a
    "01000000", --  954 - 0x3ba  :   64 - 0x40
    "00000010", --  955 - 0x3bb  :    2 - 0x2
    "01000000", --  956 - 0x3bc  :   64 - 0x40
    "00000010", --  957 - 0x3bd  :    2 - 0x2
    "01010100", --  958 - 0x3be  :   84 - 0x54
    "00000000", --  959 - 0x3bf  :    0 - 0x0
    "11111111", --  960 - 0x3c0  :  255 - 0xff -- Background 0x3c
    "11111111", --  961 - 0x3c1  :  255 - 0xff
    "11111111", --  962 - 0x3c2  :  255 - 0xff
    "11111111", --  963 - 0x3c3  :  255 - 0xff
    "11111111", --  964 - 0x3c4  :  255 - 0xff
    "11111111", --  965 - 0x3c5  :  255 - 0xff
    "11111111", --  966 - 0x3c6  :  255 - 0xff
    "11111111", --  967 - 0x3c7  :  255 - 0xff
    "00000000", --  968 - 0x3c8  :    0 - 0x0 -- plane 1
    "00000000", --  969 - 0x3c9  :    0 - 0x0
    "00000000", --  970 - 0x3ca  :    0 - 0x0
    "00000000", --  971 - 0x3cb  :    0 - 0x0
    "00000000", --  972 - 0x3cc  :    0 - 0x0
    "00000000", --  973 - 0x3cd  :    0 - 0x0
    "00000000", --  974 - 0x3ce  :    0 - 0x0
    "00000000", --  975 - 0x3cf  :    0 - 0x0
    "00000000", --  976 - 0x3d0  :    0 - 0x0 -- Background 0x3d
    "00000000", --  977 - 0x3d1  :    0 - 0x0
    "00000000", --  978 - 0x3d2  :    0 - 0x0
    "00000000", --  979 - 0x3d3  :    0 - 0x0
    "00000000", --  980 - 0x3d4  :    0 - 0x0
    "00000000", --  981 - 0x3d5  :    0 - 0x0
    "00000000", --  982 - 0x3d6  :    0 - 0x0
    "00000000", --  983 - 0x3d7  :    0 - 0x0
    "11111111", --  984 - 0x3d8  :  255 - 0xff -- plane 1
    "11111111", --  985 - 0x3d9  :  255 - 0xff
    "11111111", --  986 - 0x3da  :  255 - 0xff
    "11111111", --  987 - 0x3db  :  255 - 0xff
    "11111111", --  988 - 0x3dc  :  255 - 0xff
    "11111111", --  989 - 0x3dd  :  255 - 0xff
    "11111111", --  990 - 0x3de  :  255 - 0xff
    "11111111", --  991 - 0x3df  :  255 - 0xff
    "11111111", --  992 - 0x3e0  :  255 - 0xff -- Background 0x3e
    "11111111", --  993 - 0x3e1  :  255 - 0xff
    "11111111", --  994 - 0x3e2  :  255 - 0xff
    "11111111", --  995 - 0x3e3  :  255 - 0xff
    "11111111", --  996 - 0x3e4  :  255 - 0xff
    "11111111", --  997 - 0x3e5  :  255 - 0xff
    "11111111", --  998 - 0x3e6  :  255 - 0xff
    "11111111", --  999 - 0x3e7  :  255 - 0xff
    "11111111", -- 1000 - 0x3e8  :  255 - 0xff -- plane 1
    "11111111", -- 1001 - 0x3e9  :  255 - 0xff
    "11111111", -- 1002 - 0x3ea  :  255 - 0xff
    "11111111", -- 1003 - 0x3eb  :  255 - 0xff
    "11111111", -- 1004 - 0x3ec  :  255 - 0xff
    "11111111", -- 1005 - 0x3ed  :  255 - 0xff
    "11111111", -- 1006 - 0x3ee  :  255 - 0xff
    "11111111", -- 1007 - 0x3ef  :  255 - 0xff
    "00000000", -- 1008 - 0x3f0  :    0 - 0x0 -- Background 0x3f
    "00000000", -- 1009 - 0x3f1  :    0 - 0x0
    "00000000", -- 1010 - 0x3f2  :    0 - 0x0
    "00000000", -- 1011 - 0x3f3  :    0 - 0x0
    "00000000", -- 1012 - 0x3f4  :    0 - 0x0
    "00000000", -- 1013 - 0x3f5  :    0 - 0x0
    "00000000", -- 1014 - 0x3f6  :    0 - 0x0
    "00000000", -- 1015 - 0x3f7  :    0 - 0x0
    "00000000", -- 1016 - 0x3f8  :    0 - 0x0 -- plane 1
    "00000000", -- 1017 - 0x3f9  :    0 - 0x0
    "00000000", -- 1018 - 0x3fa  :    0 - 0x0
    "00000000", -- 1019 - 0x3fb  :    0 - 0x0
    "00000000", -- 1020 - 0x3fc  :    0 - 0x0
    "00000000", -- 1021 - 0x3fd  :    0 - 0x0
    "00000000", -- 1022 - 0x3fe  :    0 - 0x0
    "00000000", -- 1023 - 0x3ff  :    0 - 0x0
    "00111100", -- 1024 - 0x400  :   60 - 0x3c -- Background 0x40
    "01000010", -- 1025 - 0x401  :   66 - 0x42
    "10011001", -- 1026 - 0x402  :  153 - 0x99
    "10100101", -- 1027 - 0x403  :  165 - 0xa5
    "10100101", -- 1028 - 0x404  :  165 - 0xa5
    "10011010", -- 1029 - 0x405  :  154 - 0x9a
    "01000000", -- 1030 - 0x406  :   64 - 0x40
    "00111100", -- 1031 - 0x407  :   60 - 0x3c
    "00000000", -- 1032 - 0x408  :    0 - 0x0 -- plane 1
    "00000000", -- 1033 - 0x409  :    0 - 0x0
    "00000000", -- 1034 - 0x40a  :    0 - 0x0
    "00000000", -- 1035 - 0x40b  :    0 - 0x0
    "00000000", -- 1036 - 0x40c  :    0 - 0x0
    "00000000", -- 1037 - 0x40d  :    0 - 0x0
    "00000000", -- 1038 - 0x40e  :    0 - 0x0
    "00000000", -- 1039 - 0x40f  :    0 - 0x0
    "00001100", -- 1040 - 0x410  :   12 - 0xc -- Background 0x41
    "00010010", -- 1041 - 0x411  :   18 - 0x12
    "00100010", -- 1042 - 0x412  :   34 - 0x22
    "00100010", -- 1043 - 0x413  :   34 - 0x22
    "01111110", -- 1044 - 0x414  :  126 - 0x7e
    "00100010", -- 1045 - 0x415  :   34 - 0x22
    "00100100", -- 1046 - 0x416  :   36 - 0x24
    "00000000", -- 1047 - 0x417  :    0 - 0x0
    "00000000", -- 1048 - 0x418  :    0 - 0x0 -- plane 1
    "00000000", -- 1049 - 0x419  :    0 - 0x0
    "00000000", -- 1050 - 0x41a  :    0 - 0x0
    "00000000", -- 1051 - 0x41b  :    0 - 0x0
    "00000000", -- 1052 - 0x41c  :    0 - 0x0
    "00000000", -- 1053 - 0x41d  :    0 - 0x0
    "00000000", -- 1054 - 0x41e  :    0 - 0x0
    "00000000", -- 1055 - 0x41f  :    0 - 0x0
    "00111100", -- 1056 - 0x420  :   60 - 0x3c -- Background 0x42
    "01000010", -- 1057 - 0x421  :   66 - 0x42
    "01010010", -- 1058 - 0x422  :   82 - 0x52
    "00011100", -- 1059 - 0x423  :   28 - 0x1c
    "00010010", -- 1060 - 0x424  :   18 - 0x12
    "00110010", -- 1061 - 0x425  :   50 - 0x32
    "00011100", -- 1062 - 0x426  :   28 - 0x1c
    "00000000", -- 1063 - 0x427  :    0 - 0x0
    "00000000", -- 1064 - 0x428  :    0 - 0x0 -- plane 1
    "00000000", -- 1065 - 0x429  :    0 - 0x0
    "00000000", -- 1066 - 0x42a  :    0 - 0x0
    "00000000", -- 1067 - 0x42b  :    0 - 0x0
    "00000000", -- 1068 - 0x42c  :    0 - 0x0
    "00000000", -- 1069 - 0x42d  :    0 - 0x0
    "00000000", -- 1070 - 0x42e  :    0 - 0x0
    "00000000", -- 1071 - 0x42f  :    0 - 0x0
    "00011000", -- 1072 - 0x430  :   24 - 0x18 -- Background 0x43
    "00100100", -- 1073 - 0x431  :   36 - 0x24
    "01010100", -- 1074 - 0x432  :   84 - 0x54
    "01001000", -- 1075 - 0x433  :   72 - 0x48
    "01000010", -- 1076 - 0x434  :   66 - 0x42
    "00100100", -- 1077 - 0x435  :   36 - 0x24
    "00011000", -- 1078 - 0x436  :   24 - 0x18
    "00000000", -- 1079 - 0x437  :    0 - 0x0
    "00000000", -- 1080 - 0x438  :    0 - 0x0 -- plane 1
    "00000000", -- 1081 - 0x439  :    0 - 0x0
    "00000000", -- 1082 - 0x43a  :    0 - 0x0
    "00000000", -- 1083 - 0x43b  :    0 - 0x0
    "00000000", -- 1084 - 0x43c  :    0 - 0x0
    "00000000", -- 1085 - 0x43d  :    0 - 0x0
    "00000000", -- 1086 - 0x43e  :    0 - 0x0
    "00000000", -- 1087 - 0x43f  :    0 - 0x0
    "01011000", -- 1088 - 0x440  :   88 - 0x58 -- Background 0x44
    "11100100", -- 1089 - 0x441  :  228 - 0xe4
    "01000010", -- 1090 - 0x442  :   66 - 0x42
    "01000010", -- 1091 - 0x443  :   66 - 0x42
    "00100010", -- 1092 - 0x444  :   34 - 0x22
    "01100100", -- 1093 - 0x445  :  100 - 0x64
    "00111000", -- 1094 - 0x446  :   56 - 0x38
    "00000000", -- 1095 - 0x447  :    0 - 0x0
    "00000000", -- 1096 - 0x448  :    0 - 0x0 -- plane 1
    "00000000", -- 1097 - 0x449  :    0 - 0x0
    "00000000", -- 1098 - 0x44a  :    0 - 0x0
    "00000000", -- 1099 - 0x44b  :    0 - 0x0
    "00000000", -- 1100 - 0x44c  :    0 - 0x0
    "00000000", -- 1101 - 0x44d  :    0 - 0x0
    "00000000", -- 1102 - 0x44e  :    0 - 0x0
    "00000000", -- 1103 - 0x44f  :    0 - 0x0
    "00011100", -- 1104 - 0x450  :   28 - 0x1c -- Background 0x45
    "00100000", -- 1105 - 0x451  :   32 - 0x20
    "00100000", -- 1106 - 0x452  :   32 - 0x20
    "00101100", -- 1107 - 0x453  :   44 - 0x2c
    "01110000", -- 1108 - 0x454  :  112 - 0x70
    "00100010", -- 1109 - 0x455  :   34 - 0x22
    "00011100", -- 1110 - 0x456  :   28 - 0x1c
    "00000000", -- 1111 - 0x457  :    0 - 0x0
    "00000000", -- 1112 - 0x458  :    0 - 0x0 -- plane 1
    "00000000", -- 1113 - 0x459  :    0 - 0x0
    "00000000", -- 1114 - 0x45a  :    0 - 0x0
    "00000000", -- 1115 - 0x45b  :    0 - 0x0
    "00000000", -- 1116 - 0x45c  :    0 - 0x0
    "00000000", -- 1117 - 0x45d  :    0 - 0x0
    "00000000", -- 1118 - 0x45e  :    0 - 0x0
    "00000000", -- 1119 - 0x45f  :    0 - 0x0
    "00011100", -- 1120 - 0x460  :   28 - 0x1c -- Background 0x46
    "00100000", -- 1121 - 0x461  :   32 - 0x20
    "00100000", -- 1122 - 0x462  :   32 - 0x20
    "00101100", -- 1123 - 0x463  :   44 - 0x2c
    "01110000", -- 1124 - 0x464  :  112 - 0x70
    "00010000", -- 1125 - 0x465  :   16 - 0x10
    "00010000", -- 1126 - 0x466  :   16 - 0x10
    "00000000", -- 1127 - 0x467  :    0 - 0x0
    "00000000", -- 1128 - 0x468  :    0 - 0x0 -- plane 1
    "00000000", -- 1129 - 0x469  :    0 - 0x0
    "00000000", -- 1130 - 0x46a  :    0 - 0x0
    "00000000", -- 1131 - 0x46b  :    0 - 0x0
    "00000000", -- 1132 - 0x46c  :    0 - 0x0
    "00000000", -- 1133 - 0x46d  :    0 - 0x0
    "00000000", -- 1134 - 0x46e  :    0 - 0x0
    "00000000", -- 1135 - 0x46f  :    0 - 0x0
    "00011000", -- 1136 - 0x470  :   24 - 0x18 -- Background 0x47
    "00100100", -- 1137 - 0x471  :   36 - 0x24
    "01000000", -- 1138 - 0x472  :   64 - 0x40
    "01001110", -- 1139 - 0x473  :   78 - 0x4e
    "01000010", -- 1140 - 0x474  :   66 - 0x42
    "00100100", -- 1141 - 0x475  :   36 - 0x24
    "00011000", -- 1142 - 0x476  :   24 - 0x18
    "00000000", -- 1143 - 0x477  :    0 - 0x0
    "00000000", -- 1144 - 0x478  :    0 - 0x0 -- plane 1
    "00000000", -- 1145 - 0x479  :    0 - 0x0
    "00000000", -- 1146 - 0x47a  :    0 - 0x0
    "00000000", -- 1147 - 0x47b  :    0 - 0x0
    "00000000", -- 1148 - 0x47c  :    0 - 0x0
    "00000000", -- 1149 - 0x47d  :    0 - 0x0
    "00000000", -- 1150 - 0x47e  :    0 - 0x0
    "00000000", -- 1151 - 0x47f  :    0 - 0x0
    "00100000", -- 1152 - 0x480  :   32 - 0x20 -- Background 0x48
    "01000100", -- 1153 - 0x481  :   68 - 0x44
    "01000100", -- 1154 - 0x482  :   68 - 0x44
    "01000100", -- 1155 - 0x483  :   68 - 0x44
    "11111100", -- 1156 - 0x484  :  252 - 0xfc
    "01000100", -- 1157 - 0x485  :   68 - 0x44
    "01001000", -- 1158 - 0x486  :   72 - 0x48
    "00000000", -- 1159 - 0x487  :    0 - 0x0
    "00000000", -- 1160 - 0x488  :    0 - 0x0 -- plane 1
    "00000000", -- 1161 - 0x489  :    0 - 0x0
    "00000000", -- 1162 - 0x48a  :    0 - 0x0
    "00000000", -- 1163 - 0x48b  :    0 - 0x0
    "00000000", -- 1164 - 0x48c  :    0 - 0x0
    "00000000", -- 1165 - 0x48d  :    0 - 0x0
    "00000000", -- 1166 - 0x48e  :    0 - 0x0
    "00000000", -- 1167 - 0x48f  :    0 - 0x0
    "00010000", -- 1168 - 0x490  :   16 - 0x10 -- Background 0x49
    "00010000", -- 1169 - 0x491  :   16 - 0x10
    "00010000", -- 1170 - 0x492  :   16 - 0x10
    "00010000", -- 1171 - 0x493  :   16 - 0x10
    "00010000", -- 1172 - 0x494  :   16 - 0x10
    "00001000", -- 1173 - 0x495  :    8 - 0x8
    "00001000", -- 1174 - 0x496  :    8 - 0x8
    "00000000", -- 1175 - 0x497  :    0 - 0x0
    "00000000", -- 1176 - 0x498  :    0 - 0x0 -- plane 1
    "00000000", -- 1177 - 0x499  :    0 - 0x0
    "00000000", -- 1178 - 0x49a  :    0 - 0x0
    "00000000", -- 1179 - 0x49b  :    0 - 0x0
    "00000000", -- 1180 - 0x49c  :    0 - 0x0
    "00000000", -- 1181 - 0x49d  :    0 - 0x0
    "00000000", -- 1182 - 0x49e  :    0 - 0x0
    "00000000", -- 1183 - 0x49f  :    0 - 0x0
    "00001000", -- 1184 - 0x4a0  :    8 - 0x8 -- Background 0x4a
    "00001000", -- 1185 - 0x4a1  :    8 - 0x8
    "00000100", -- 1186 - 0x4a2  :    4 - 0x4
    "00000100", -- 1187 - 0x4a3  :    4 - 0x4
    "01000100", -- 1188 - 0x4a4  :   68 - 0x44
    "01001000", -- 1189 - 0x4a5  :   72 - 0x48
    "00110000", -- 1190 - 0x4a6  :   48 - 0x30
    "00000000", -- 1191 - 0x4a7  :    0 - 0x0
    "00000000", -- 1192 - 0x4a8  :    0 - 0x0 -- plane 1
    "00000000", -- 1193 - 0x4a9  :    0 - 0x0
    "00000000", -- 1194 - 0x4aa  :    0 - 0x0
    "00000000", -- 1195 - 0x4ab  :    0 - 0x0
    "00000000", -- 1196 - 0x4ac  :    0 - 0x0
    "00000000", -- 1197 - 0x4ad  :    0 - 0x0
    "00000000", -- 1198 - 0x4ae  :    0 - 0x0
    "00000000", -- 1199 - 0x4af  :    0 - 0x0
    "01000100", -- 1200 - 0x4b0  :   68 - 0x44 -- Background 0x4b
    "01000100", -- 1201 - 0x4b1  :   68 - 0x44
    "01001000", -- 1202 - 0x4b2  :   72 - 0x48
    "01110000", -- 1203 - 0x4b3  :  112 - 0x70
    "01001000", -- 1204 - 0x4b4  :   72 - 0x48
    "00100100", -- 1205 - 0x4b5  :   36 - 0x24
    "00100010", -- 1206 - 0x4b6  :   34 - 0x22
    "00000000", -- 1207 - 0x4b7  :    0 - 0x0
    "00000000", -- 1208 - 0x4b8  :    0 - 0x0 -- plane 1
    "00000000", -- 1209 - 0x4b9  :    0 - 0x0
    "00000000", -- 1210 - 0x4ba  :    0 - 0x0
    "00000000", -- 1211 - 0x4bb  :    0 - 0x0
    "00000000", -- 1212 - 0x4bc  :    0 - 0x0
    "00000000", -- 1213 - 0x4bd  :    0 - 0x0
    "00000000", -- 1214 - 0x4be  :    0 - 0x0
    "00000000", -- 1215 - 0x4bf  :    0 - 0x0
    "00010000", -- 1216 - 0x4c0  :   16 - 0x10 -- Background 0x4c
    "00100000", -- 1217 - 0x4c1  :   32 - 0x20
    "00100000", -- 1218 - 0x4c2  :   32 - 0x20
    "00100000", -- 1219 - 0x4c3  :   32 - 0x20
    "01000000", -- 1220 - 0x4c4  :   64 - 0x40
    "01000000", -- 1221 - 0x4c5  :   64 - 0x40
    "01000110", -- 1222 - 0x4c6  :   70 - 0x46
    "00111000", -- 1223 - 0x4c7  :   56 - 0x38
    "00000000", -- 1224 - 0x4c8  :    0 - 0x0 -- plane 1
    "00000000", -- 1225 - 0x4c9  :    0 - 0x0
    "00000000", -- 1226 - 0x4ca  :    0 - 0x0
    "00000000", -- 1227 - 0x4cb  :    0 - 0x0
    "00000000", -- 1228 - 0x4cc  :    0 - 0x0
    "00000000", -- 1229 - 0x4cd  :    0 - 0x0
    "00000000", -- 1230 - 0x4ce  :    0 - 0x0
    "00000000", -- 1231 - 0x4cf  :    0 - 0x0
    "00100100", -- 1232 - 0x4d0  :   36 - 0x24 -- Background 0x4d
    "01011010", -- 1233 - 0x4d1  :   90 - 0x5a
    "01011010", -- 1234 - 0x4d2  :   90 - 0x5a
    "01011010", -- 1235 - 0x4d3  :   90 - 0x5a
    "01000010", -- 1236 - 0x4d4  :   66 - 0x42
    "01000010", -- 1237 - 0x4d5  :   66 - 0x42
    "00100010", -- 1238 - 0x4d6  :   34 - 0x22
    "00000000", -- 1239 - 0x4d7  :    0 - 0x0
    "00000000", -- 1240 - 0x4d8  :    0 - 0x0 -- plane 1
    "00000000", -- 1241 - 0x4d9  :    0 - 0x0
    "00000000", -- 1242 - 0x4da  :    0 - 0x0
    "00000000", -- 1243 - 0x4db  :    0 - 0x0
    "00000000", -- 1244 - 0x4dc  :    0 - 0x0
    "00000000", -- 1245 - 0x4dd  :    0 - 0x0
    "00000000", -- 1246 - 0x4de  :    0 - 0x0
    "00000000", -- 1247 - 0x4df  :    0 - 0x0
    "00100100", -- 1248 - 0x4e0  :   36 - 0x24 -- Background 0x4e
    "01010010", -- 1249 - 0x4e1  :   82 - 0x52
    "01010010", -- 1250 - 0x4e2  :   82 - 0x52
    "01010010", -- 1251 - 0x4e3  :   82 - 0x52
    "01010010", -- 1252 - 0x4e4  :   82 - 0x52
    "01010010", -- 1253 - 0x4e5  :   82 - 0x52
    "01001100", -- 1254 - 0x4e6  :   76 - 0x4c
    "00000000", -- 1255 - 0x4e7  :    0 - 0x0
    "00000000", -- 1256 - 0x4e8  :    0 - 0x0 -- plane 1
    "00000000", -- 1257 - 0x4e9  :    0 - 0x0
    "00000000", -- 1258 - 0x4ea  :    0 - 0x0
    "00000000", -- 1259 - 0x4eb  :    0 - 0x0
    "00000000", -- 1260 - 0x4ec  :    0 - 0x0
    "00000000", -- 1261 - 0x4ed  :    0 - 0x0
    "00000000", -- 1262 - 0x4ee  :    0 - 0x0
    "00000000", -- 1263 - 0x4ef  :    0 - 0x0
    "00111000", -- 1264 - 0x4f0  :   56 - 0x38 -- Background 0x4f
    "01000100", -- 1265 - 0x4f1  :   68 - 0x44
    "10000010", -- 1266 - 0x4f2  :  130 - 0x82
    "10000010", -- 1267 - 0x4f3  :  130 - 0x82
    "10000010", -- 1268 - 0x4f4  :  130 - 0x82
    "01000100", -- 1269 - 0x4f5  :   68 - 0x44
    "00111000", -- 1270 - 0x4f6  :   56 - 0x38
    "00000000", -- 1271 - 0x4f7  :    0 - 0x0
    "00000000", -- 1272 - 0x4f8  :    0 - 0x0 -- plane 1
    "00000000", -- 1273 - 0x4f9  :    0 - 0x0
    "00000000", -- 1274 - 0x4fa  :    0 - 0x0
    "00000000", -- 1275 - 0x4fb  :    0 - 0x0
    "00000000", -- 1276 - 0x4fc  :    0 - 0x0
    "00000000", -- 1277 - 0x4fd  :    0 - 0x0
    "00000000", -- 1278 - 0x4fe  :    0 - 0x0
    "00000000", -- 1279 - 0x4ff  :    0 - 0x0
    "01111111", -- 1280 - 0x500  :  127 - 0x7f -- Background 0x50
    "11000000", -- 1281 - 0x501  :  192 - 0xc0
    "10000000", -- 1282 - 0x502  :  128 - 0x80
    "10000000", -- 1283 - 0x503  :  128 - 0x80
    "10000000", -- 1284 - 0x504  :  128 - 0x80
    "11000011", -- 1285 - 0x505  :  195 - 0xc3
    "11111111", -- 1286 - 0x506  :  255 - 0xff
    "11111111", -- 1287 - 0x507  :  255 - 0xff
    "00000000", -- 1288 - 0x508  :    0 - 0x0 -- plane 1
    "00111111", -- 1289 - 0x509  :   63 - 0x3f
    "01111111", -- 1290 - 0x50a  :  127 - 0x7f
    "01111111", -- 1291 - 0x50b  :  127 - 0x7f
    "01111111", -- 1292 - 0x50c  :  127 - 0x7f
    "00111100", -- 1293 - 0x50d  :   60 - 0x3c
    "00000000", -- 1294 - 0x50e  :    0 - 0x0
    "01000000", -- 1295 - 0x50f  :   64 - 0x40
    "11111110", -- 1296 - 0x510  :  254 - 0xfe -- Background 0x51
    "00000011", -- 1297 - 0x511  :    3 - 0x3
    "00000001", -- 1298 - 0x512  :    1 - 0x1
    "00000001", -- 1299 - 0x513  :    1 - 0x1
    "00000001", -- 1300 - 0x514  :    1 - 0x1
    "11000011", -- 1301 - 0x515  :  195 - 0xc3
    "11111111", -- 1302 - 0x516  :  255 - 0xff
    "11111111", -- 1303 - 0x517  :  255 - 0xff
    "00000000", -- 1304 - 0x518  :    0 - 0x0 -- plane 1
    "11111100", -- 1305 - 0x519  :  252 - 0xfc
    "11111110", -- 1306 - 0x51a  :  254 - 0xfe
    "11111110", -- 1307 - 0x51b  :  254 - 0xfe
    "11111110", -- 1308 - 0x51c  :  254 - 0xfe
    "00111100", -- 1309 - 0x51d  :   60 - 0x3c
    "00000000", -- 1310 - 0x51e  :    0 - 0x0
    "00000010", -- 1311 - 0x51f  :    2 - 0x2
    "00000000", -- 1312 - 0x520  :    0 - 0x0 -- Background 0x52
    "00000111", -- 1313 - 0x521  :    7 - 0x7
    "00001100", -- 1314 - 0x522  :   12 - 0xc
    "00011000", -- 1315 - 0x523  :   24 - 0x18
    "00110000", -- 1316 - 0x524  :   48 - 0x30
    "01100000", -- 1317 - 0x525  :   96 - 0x60
    "01000000", -- 1318 - 0x526  :   64 - 0x40
    "01001111", -- 1319 - 0x527  :   79 - 0x4f
    "00000000", -- 1320 - 0x528  :    0 - 0x0 -- plane 1
    "00000000", -- 1321 - 0x529  :    0 - 0x0
    "00000011", -- 1322 - 0x52a  :    3 - 0x3
    "00000111", -- 1323 - 0x52b  :    7 - 0x7
    "00001111", -- 1324 - 0x52c  :   15 - 0xf
    "00011111", -- 1325 - 0x52d  :   31 - 0x1f
    "00111111", -- 1326 - 0x52e  :   63 - 0x3f
    "00110000", -- 1327 - 0x52f  :   48 - 0x30
    "00000000", -- 1328 - 0x530  :    0 - 0x0 -- Background 0x53
    "11110000", -- 1329 - 0x531  :  240 - 0xf0
    "01010000", -- 1330 - 0x532  :   80 - 0x50
    "01001000", -- 1331 - 0x533  :   72 - 0x48
    "01001100", -- 1332 - 0x534  :   76 - 0x4c
    "01000100", -- 1333 - 0x535  :   68 - 0x44
    "10000010", -- 1334 - 0x536  :  130 - 0x82
    "10000011", -- 1335 - 0x537  :  131 - 0x83
    "00000000", -- 1336 - 0x538  :    0 - 0x0 -- plane 1
    "00000000", -- 1337 - 0x539  :    0 - 0x0
    "10100000", -- 1338 - 0x53a  :  160 - 0xa0
    "10110000", -- 1339 - 0x53b  :  176 - 0xb0
    "10110000", -- 1340 - 0x53c  :  176 - 0xb0
    "10111000", -- 1341 - 0x53d  :  184 - 0xb8
    "01111100", -- 1342 - 0x53e  :  124 - 0x7c
    "01111100", -- 1343 - 0x53f  :  124 - 0x7c
    "01111111", -- 1344 - 0x540  :  127 - 0x7f -- Background 0x54
    "11011110", -- 1345 - 0x541  :  222 - 0xde
    "10001110", -- 1346 - 0x542  :  142 - 0x8e
    "11000101", -- 1347 - 0x543  :  197 - 0xc5
    "10010010", -- 1348 - 0x544  :  146 - 0x92
    "11000111", -- 1349 - 0x545  :  199 - 0xc7
    "11100010", -- 1350 - 0x546  :  226 - 0xe2
    "11010000", -- 1351 - 0x547  :  208 - 0xd0
    "00000000", -- 1352 - 0x548  :    0 - 0x0 -- plane 1
    "00100001", -- 1353 - 0x549  :   33 - 0x21
    "01110001", -- 1354 - 0x54a  :  113 - 0x71
    "00111010", -- 1355 - 0x54b  :   58 - 0x3a
    "01101101", -- 1356 - 0x54c  :  109 - 0x6d
    "00111000", -- 1357 - 0x54d  :   56 - 0x38
    "00011101", -- 1358 - 0x54e  :   29 - 0x1d
    "00101111", -- 1359 - 0x54f  :   47 - 0x2f
    "11111111", -- 1360 - 0x550  :  255 - 0xff -- Background 0x55
    "11011110", -- 1361 - 0x551  :  222 - 0xde
    "10001110", -- 1362 - 0x552  :  142 - 0x8e
    "11000101", -- 1363 - 0x553  :  197 - 0xc5
    "10010010", -- 1364 - 0x554  :  146 - 0x92
    "01000111", -- 1365 - 0x555  :   71 - 0x47
    "11100010", -- 1366 - 0x556  :  226 - 0xe2
    "01010000", -- 1367 - 0x557  :   80 - 0x50
    "00000000", -- 1368 - 0x558  :    0 - 0x0 -- plane 1
    "00100001", -- 1369 - 0x559  :   33 - 0x21
    "01110001", -- 1370 - 0x55a  :  113 - 0x71
    "00111010", -- 1371 - 0x55b  :   58 - 0x3a
    "01101101", -- 1372 - 0x55c  :  109 - 0x6d
    "10111000", -- 1373 - 0x55d  :  184 - 0xb8
    "00011101", -- 1374 - 0x55e  :   29 - 0x1d
    "10101111", -- 1375 - 0x55f  :  175 - 0xaf
    "11111110", -- 1376 - 0x560  :  254 - 0xfe -- Background 0x56
    "11011111", -- 1377 - 0x561  :  223 - 0xdf
    "10001111", -- 1378 - 0x562  :  143 - 0x8f
    "11000101", -- 1379 - 0x563  :  197 - 0xc5
    "10010011", -- 1380 - 0x564  :  147 - 0x93
    "01000111", -- 1381 - 0x565  :   71 - 0x47
    "11100011", -- 1382 - 0x566  :  227 - 0xe3
    "01010001", -- 1383 - 0x567  :   81 - 0x51
    "00000000", -- 1384 - 0x568  :    0 - 0x0 -- plane 1
    "00100000", -- 1385 - 0x569  :   32 - 0x20
    "01110000", -- 1386 - 0x56a  :  112 - 0x70
    "00111010", -- 1387 - 0x56b  :   58 - 0x3a
    "01101100", -- 1388 - 0x56c  :  108 - 0x6c
    "10111000", -- 1389 - 0x56d  :  184 - 0xb8
    "00011100", -- 1390 - 0x56e  :   28 - 0x1c
    "10101110", -- 1391 - 0x56f  :  174 - 0xae
    "01111111", -- 1392 - 0x570  :  127 - 0x7f -- Background 0x57
    "10000000", -- 1393 - 0x571  :  128 - 0x80
    "10110011", -- 1394 - 0x572  :  179 - 0xb3
    "01001100", -- 1395 - 0x573  :   76 - 0x4c
    "00111111", -- 1396 - 0x574  :   63 - 0x3f
    "00000011", -- 1397 - 0x575  :    3 - 0x3
    "00000000", -- 1398 - 0x576  :    0 - 0x0
    "00000000", -- 1399 - 0x577  :    0 - 0x0
    "00000000", -- 1400 - 0x578  :    0 - 0x0 -- plane 1
    "01111111", -- 1401 - 0x579  :  127 - 0x7f
    "01001100", -- 1402 - 0x57a  :   76 - 0x4c
    "00110011", -- 1403 - 0x57b  :   51 - 0x33
    "00000000", -- 1404 - 0x57c  :    0 - 0x0
    "00000000", -- 1405 - 0x57d  :    0 - 0x0
    "00000000", -- 1406 - 0x57e  :    0 - 0x0
    "00000000", -- 1407 - 0x57f  :    0 - 0x0
    "11111111", -- 1408 - 0x580  :  255 - 0xff -- Background 0x58
    "00000000", -- 1409 - 0x581  :    0 - 0x0
    "00110011", -- 1410 - 0x582  :   51 - 0x33
    "11001100", -- 1411 - 0x583  :  204 - 0xcc
    "00110011", -- 1412 - 0x584  :   51 - 0x33
    "11111111", -- 1413 - 0x585  :  255 - 0xff
    "00000000", -- 1414 - 0x586  :    0 - 0x0
    "00000000", -- 1415 - 0x587  :    0 - 0x0
    "00000000", -- 1416 - 0x588  :    0 - 0x0 -- plane 1
    "11111111", -- 1417 - 0x589  :  255 - 0xff
    "11001100", -- 1418 - 0x58a  :  204 - 0xcc
    "00110011", -- 1419 - 0x58b  :   51 - 0x33
    "11001100", -- 1420 - 0x58c  :  204 - 0xcc
    "00000000", -- 1421 - 0x58d  :    0 - 0x0
    "00000000", -- 1422 - 0x58e  :    0 - 0x0
    "00000000", -- 1423 - 0x58f  :    0 - 0x0
    "11111110", -- 1424 - 0x590  :  254 - 0xfe -- Background 0x59
    "00000001", -- 1425 - 0x591  :    1 - 0x1
    "00110011", -- 1426 - 0x592  :   51 - 0x33
    "11001110", -- 1427 - 0x593  :  206 - 0xce
    "00111100", -- 1428 - 0x594  :   60 - 0x3c
    "11000000", -- 1429 - 0x595  :  192 - 0xc0
    "00000000", -- 1430 - 0x596  :    0 - 0x0
    "00000000", -- 1431 - 0x597  :    0 - 0x0
    "00000000", -- 1432 - 0x598  :    0 - 0x0 -- plane 1
    "11111110", -- 1433 - 0x599  :  254 - 0xfe
    "11001100", -- 1434 - 0x59a  :  204 - 0xcc
    "00110000", -- 1435 - 0x59b  :   48 - 0x30
    "11000000", -- 1436 - 0x59c  :  192 - 0xc0
    "00000000", -- 1437 - 0x59d  :    0 - 0x0
    "00000000", -- 1438 - 0x59e  :    0 - 0x0
    "00000000", -- 1439 - 0x59f  :    0 - 0x0
    "00000000", -- 1440 - 0x5a0  :    0 - 0x0 -- Background 0x5a
    "00000000", -- 1441 - 0x5a1  :    0 - 0x0
    "00000000", -- 1442 - 0x5a2  :    0 - 0x0
    "00000000", -- 1443 - 0x5a3  :    0 - 0x0
    "00000000", -- 1444 - 0x5a4  :    0 - 0x0
    "00000000", -- 1445 - 0x5a5  :    0 - 0x0
    "00000000", -- 1446 - 0x5a6  :    0 - 0x0
    "00000000", -- 1447 - 0x5a7  :    0 - 0x0
    "00000000", -- 1448 - 0x5a8  :    0 - 0x0 -- plane 1
    "00000000", -- 1449 - 0x5a9  :    0 - 0x0
    "00000000", -- 1450 - 0x5aa  :    0 - 0x0
    "00000000", -- 1451 - 0x5ab  :    0 - 0x0
    "00000000", -- 1452 - 0x5ac  :    0 - 0x0
    "00000000", -- 1453 - 0x5ad  :    0 - 0x0
    "00000000", -- 1454 - 0x5ae  :    0 - 0x0
    "00000000", -- 1455 - 0x5af  :    0 - 0x0
    "00000000", -- 1456 - 0x5b0  :    0 - 0x0 -- Background 0x5b
    "00000000", -- 1457 - 0x5b1  :    0 - 0x0
    "00000000", -- 1458 - 0x5b2  :    0 - 0x0
    "00000001", -- 1459 - 0x5b3  :    1 - 0x1
    "00000011", -- 1460 - 0x5b4  :    3 - 0x3
    "00000011", -- 1461 - 0x5b5  :    3 - 0x3
    "00000111", -- 1462 - 0x5b6  :    7 - 0x7
    "00111111", -- 1463 - 0x5b7  :   63 - 0x3f
    "00000000", -- 1464 - 0x5b8  :    0 - 0x0 -- plane 1
    "00000000", -- 1465 - 0x5b9  :    0 - 0x0
    "00000000", -- 1466 - 0x5ba  :    0 - 0x0
    "00000000", -- 1467 - 0x5bb  :    0 - 0x0
    "00000001", -- 1468 - 0x5bc  :    1 - 0x1
    "00000001", -- 1469 - 0x5bd  :    1 - 0x1
    "00000011", -- 1470 - 0x5be  :    3 - 0x3
    "00000011", -- 1471 - 0x5bf  :    3 - 0x3
    "00000000", -- 1472 - 0x5c0  :    0 - 0x0 -- Background 0x5c
    "00000001", -- 1473 - 0x5c1  :    1 - 0x1
    "01111111", -- 1474 - 0x5c2  :  127 - 0x7f
    "11111111", -- 1475 - 0x5c3  :  255 - 0xff
    "11111111", -- 1476 - 0x5c4  :  255 - 0xff
    "11111111", -- 1477 - 0x5c5  :  255 - 0xff
    "11111111", -- 1478 - 0x5c6  :  255 - 0xff
    "11111111", -- 1479 - 0x5c7  :  255 - 0xff
    "00000000", -- 1480 - 0x5c8  :    0 - 0x0 -- plane 1
    "00000000", -- 1481 - 0x5c9  :    0 - 0x0
    "00000001", -- 1482 - 0x5ca  :    1 - 0x1
    "01111110", -- 1483 - 0x5cb  :  126 - 0x7e
    "11111111", -- 1484 - 0x5cc  :  255 - 0xff
    "11111111", -- 1485 - 0x5cd  :  255 - 0xff
    "11111111", -- 1486 - 0x5ce  :  255 - 0xff
    "11111111", -- 1487 - 0x5cf  :  255 - 0xff
    "11111111", -- 1488 - 0x5d0  :  255 - 0xff -- Background 0x5d
    "11111111", -- 1489 - 0x5d1  :  255 - 0xff
    "11111111", -- 1490 - 0x5d2  :  255 - 0xff
    "11111111", -- 1491 - 0x5d3  :  255 - 0xff
    "11111111", -- 1492 - 0x5d4  :  255 - 0xff
    "11111111", -- 1493 - 0x5d5  :  255 - 0xff
    "11111111", -- 1494 - 0x5d6  :  255 - 0xff
    "11111111", -- 1495 - 0x5d7  :  255 - 0xff
    "00000000", -- 1496 - 0x5d8  :    0 - 0x0 -- plane 1
    "11111111", -- 1497 - 0x5d9  :  255 - 0xff
    "11111111", -- 1498 - 0x5da  :  255 - 0xff
    "11111111", -- 1499 - 0x5db  :  255 - 0xff
    "01111111", -- 1500 - 0x5dc  :  127 - 0x7f
    "11111111", -- 1501 - 0x5dd  :  255 - 0xff
    "11111111", -- 1502 - 0x5de  :  255 - 0xff
    "11111111", -- 1503 - 0x5df  :  255 - 0xff
    "00000000", -- 1504 - 0x5e0  :    0 - 0x0 -- Background 0x5e
    "10000000", -- 1505 - 0x5e1  :  128 - 0x80
    "11111110", -- 1506 - 0x5e2  :  254 - 0xfe
    "11111111", -- 1507 - 0x5e3  :  255 - 0xff
    "11111111", -- 1508 - 0x5e4  :  255 - 0xff
    "11111111", -- 1509 - 0x5e5  :  255 - 0xff
    "11111111", -- 1510 - 0x5e6  :  255 - 0xff
    "11111111", -- 1511 - 0x5e7  :  255 - 0xff
    "00000000", -- 1512 - 0x5e8  :    0 - 0x0 -- plane 1
    "00000000", -- 1513 - 0x5e9  :    0 - 0x0
    "10000000", -- 1514 - 0x5ea  :  128 - 0x80
    "01111110", -- 1515 - 0x5eb  :  126 - 0x7e
    "10111111", -- 1516 - 0x5ec  :  191 - 0xbf
    "11111111", -- 1517 - 0x5ed  :  255 - 0xff
    "11111111", -- 1518 - 0x5ee  :  255 - 0xff
    "11111111", -- 1519 - 0x5ef  :  255 - 0xff
    "00000000", -- 1520 - 0x5f0  :    0 - 0x0 -- Background 0x5f
    "00000000", -- 1521 - 0x5f1  :    0 - 0x0
    "00000000", -- 1522 - 0x5f2  :    0 - 0x0
    "10000000", -- 1523 - 0x5f3  :  128 - 0x80
    "11000000", -- 1524 - 0x5f4  :  192 - 0xc0
    "11000000", -- 1525 - 0x5f5  :  192 - 0xc0
    "11100000", -- 1526 - 0x5f6  :  224 - 0xe0
    "11111000", -- 1527 - 0x5f7  :  248 - 0xf8
    "00000000", -- 1528 - 0x5f8  :    0 - 0x0 -- plane 1
    "00000000", -- 1529 - 0x5f9  :    0 - 0x0
    "00000000", -- 1530 - 0x5fa  :    0 - 0x0
    "00000000", -- 1531 - 0x5fb  :    0 - 0x0
    "10000000", -- 1532 - 0x5fc  :  128 - 0x80
    "10000000", -- 1533 - 0x5fd  :  128 - 0x80
    "11000000", -- 1534 - 0x5fe  :  192 - 0xc0
    "11000000", -- 1535 - 0x5ff  :  192 - 0xc0
    "11111111", -- 1536 - 0x600  :  255 - 0xff -- Background 0x60
    "11111111", -- 1537 - 0x601  :  255 - 0xff
    "11111111", -- 1538 - 0x602  :  255 - 0xff
    "11111111", -- 1539 - 0x603  :  255 - 0xff
    "11111111", -- 1540 - 0x604  :  255 - 0xff
    "11111111", -- 1541 - 0x605  :  255 - 0xff
    "11111111", -- 1542 - 0x606  :  255 - 0xff
    "11111111", -- 1543 - 0x607  :  255 - 0xff
    "01111111", -- 1544 - 0x608  :  127 - 0x7f -- plane 1
    "01111111", -- 1545 - 0x609  :  127 - 0x7f
    "01111101", -- 1546 - 0x60a  :  125 - 0x7d
    "01111111", -- 1547 - 0x60b  :  127 - 0x7f
    "00111111", -- 1548 - 0x60c  :   63 - 0x3f
    "01111111", -- 1549 - 0x60d  :  127 - 0x7f
    "01111111", -- 1550 - 0x60e  :  127 - 0x7f
    "01110111", -- 1551 - 0x60f  :  119 - 0x77
    "11111111", -- 1552 - 0x610  :  255 - 0xff -- Background 0x61
    "11111111", -- 1553 - 0x611  :  255 - 0xff
    "11111111", -- 1554 - 0x612  :  255 - 0xff
    "11111111", -- 1555 - 0x613  :  255 - 0xff
    "11111111", -- 1556 - 0x614  :  255 - 0xff
    "11111111", -- 1557 - 0x615  :  255 - 0xff
    "11111111", -- 1558 - 0x616  :  255 - 0xff
    "11111111", -- 1559 - 0x617  :  255 - 0xff
    "11111110", -- 1560 - 0x618  :  254 - 0xfe -- plane 1
    "11111110", -- 1561 - 0x619  :  254 - 0xfe
    "11111100", -- 1562 - 0x61a  :  252 - 0xfc
    "11111110", -- 1563 - 0x61b  :  254 - 0xfe
    "10111110", -- 1564 - 0x61c  :  190 - 0xbe
    "11111110", -- 1565 - 0x61d  :  254 - 0xfe
    "11111110", -- 1566 - 0x61e  :  254 - 0xfe
    "11110110", -- 1567 - 0x61f  :  246 - 0xf6
    "01111000", -- 1568 - 0x620  :  120 - 0x78 -- Background 0x62
    "01100000", -- 1569 - 0x621  :   96 - 0x60
    "01000000", -- 1570 - 0x622  :   64 - 0x40
    "01000000", -- 1571 - 0x623  :   64 - 0x40
    "01000000", -- 1572 - 0x624  :   64 - 0x40
    "01100000", -- 1573 - 0x625  :   96 - 0x60
    "00110000", -- 1574 - 0x626  :   48 - 0x30
    "00011111", -- 1575 - 0x627  :   31 - 0x1f
    "00000111", -- 1576 - 0x628  :    7 - 0x7 -- plane 1
    "00011111", -- 1577 - 0x629  :   31 - 0x1f
    "00111111", -- 1578 - 0x62a  :   63 - 0x3f
    "00111111", -- 1579 - 0x62b  :   63 - 0x3f
    "00111111", -- 1580 - 0x62c  :   63 - 0x3f
    "00011111", -- 1581 - 0x62d  :   31 - 0x1f
    "00001111", -- 1582 - 0x62e  :   15 - 0xf
    "00000000", -- 1583 - 0x62f  :    0 - 0x0
    "10000001", -- 1584 - 0x630  :  129 - 0x81 -- Background 0x63
    "10000011", -- 1585 - 0x631  :  131 - 0x83
    "11000001", -- 1586 - 0x632  :  193 - 0xc1
    "01000011", -- 1587 - 0x633  :   67 - 0x43
    "01000001", -- 1588 - 0x634  :   65 - 0x41
    "01100011", -- 1589 - 0x635  :   99 - 0x63
    "00100110", -- 1590 - 0x636  :   38 - 0x26
    "11111000", -- 1591 - 0x637  :  248 - 0xf8
    "01111110", -- 1592 - 0x638  :  126 - 0x7e -- plane 1
    "01111100", -- 1593 - 0x639  :  124 - 0x7c
    "00111110", -- 1594 - 0x63a  :   62 - 0x3e
    "10111100", -- 1595 - 0x63b  :  188 - 0xbc
    "10111110", -- 1596 - 0x63c  :  190 - 0xbe
    "10011100", -- 1597 - 0x63d  :  156 - 0x9c
    "11011000", -- 1598 - 0x63e  :  216 - 0xd8
    "00000000", -- 1599 - 0x63f  :    0 - 0x0
    "10111001", -- 1600 - 0x640  :  185 - 0xb9 -- Background 0x64
    "10010100", -- 1601 - 0x641  :  148 - 0x94
    "10001110", -- 1602 - 0x642  :  142 - 0x8e
    "11000101", -- 1603 - 0x643  :  197 - 0xc5
    "10010010", -- 1604 - 0x644  :  146 - 0x92
    "11000111", -- 1605 - 0x645  :  199 - 0xc7
    "11100010", -- 1606 - 0x646  :  226 - 0xe2
    "11010000", -- 1607 - 0x647  :  208 - 0xd0
    "01000110", -- 1608 - 0x648  :   70 - 0x46 -- plane 1
    "01101011", -- 1609 - 0x649  :  107 - 0x6b
    "01110001", -- 1610 - 0x64a  :  113 - 0x71
    "00111010", -- 1611 - 0x64b  :   58 - 0x3a
    "01101101", -- 1612 - 0x64c  :  109 - 0x6d
    "00111000", -- 1613 - 0x64d  :   56 - 0x38
    "00011101", -- 1614 - 0x64e  :   29 - 0x1d
    "00101111", -- 1615 - 0x64f  :   47 - 0x2f
    "10111001", -- 1616 - 0x650  :  185 - 0xb9 -- Background 0x65
    "00010100", -- 1617 - 0x651  :   20 - 0x14
    "10001110", -- 1618 - 0x652  :  142 - 0x8e
    "11000101", -- 1619 - 0x653  :  197 - 0xc5
    "10010010", -- 1620 - 0x654  :  146 - 0x92
    "01000111", -- 1621 - 0x655  :   71 - 0x47
    "11100010", -- 1622 - 0x656  :  226 - 0xe2
    "01010000", -- 1623 - 0x657  :   80 - 0x50
    "01000110", -- 1624 - 0x658  :   70 - 0x46 -- plane 1
    "11101011", -- 1625 - 0x659  :  235 - 0xeb
    "01110001", -- 1626 - 0x65a  :  113 - 0x71
    "00111010", -- 1627 - 0x65b  :   58 - 0x3a
    "01101101", -- 1628 - 0x65c  :  109 - 0x6d
    "10111000", -- 1629 - 0x65d  :  184 - 0xb8
    "00011101", -- 1630 - 0x65e  :   29 - 0x1d
    "10101111", -- 1631 - 0x65f  :  175 - 0xaf
    "10111001", -- 1632 - 0x660  :  185 - 0xb9 -- Background 0x66
    "00010101", -- 1633 - 0x661  :   21 - 0x15
    "10001111", -- 1634 - 0x662  :  143 - 0x8f
    "11000101", -- 1635 - 0x663  :  197 - 0xc5
    "10010011", -- 1636 - 0x664  :  147 - 0x93
    "01000111", -- 1637 - 0x665  :   71 - 0x47
    "11100011", -- 1638 - 0x666  :  227 - 0xe3
    "01010001", -- 1639 - 0x667  :   81 - 0x51
    "01000110", -- 1640 - 0x668  :   70 - 0x46 -- plane 1
    "11101010", -- 1641 - 0x669  :  234 - 0xea
    "01110000", -- 1642 - 0x66a  :  112 - 0x70
    "00111010", -- 1643 - 0x66b  :   58 - 0x3a
    "01101100", -- 1644 - 0x66c  :  108 - 0x6c
    "10111000", -- 1645 - 0x66d  :  184 - 0xb8
    "00011100", -- 1646 - 0x66e  :   28 - 0x1c
    "10101110", -- 1647 - 0x66f  :  174 - 0xae
    "01111111", -- 1648 - 0x670  :  127 - 0x7f -- Background 0x67
    "10000000", -- 1649 - 0x671  :  128 - 0x80
    "11001100", -- 1650 - 0x672  :  204 - 0xcc
    "01111111", -- 1651 - 0x673  :  127 - 0x7f
    "00111111", -- 1652 - 0x674  :   63 - 0x3f
    "00000011", -- 1653 - 0x675  :    3 - 0x3
    "00000000", -- 1654 - 0x676  :    0 - 0x0
    "00000000", -- 1655 - 0x677  :    0 - 0x0
    "00000000", -- 1656 - 0x678  :    0 - 0x0 -- plane 1
    "01111111", -- 1657 - 0x679  :  127 - 0x7f
    "01111111", -- 1658 - 0x67a  :  127 - 0x7f
    "00110011", -- 1659 - 0x67b  :   51 - 0x33
    "00000000", -- 1660 - 0x67c  :    0 - 0x0
    "00000000", -- 1661 - 0x67d  :    0 - 0x0
    "00000000", -- 1662 - 0x67e  :    0 - 0x0
    "00000000", -- 1663 - 0x67f  :    0 - 0x0
    "11111111", -- 1664 - 0x680  :  255 - 0xff -- Background 0x68
    "00000000", -- 1665 - 0x681  :    0 - 0x0
    "11001100", -- 1666 - 0x682  :  204 - 0xcc
    "00110011", -- 1667 - 0x683  :   51 - 0x33
    "11111111", -- 1668 - 0x684  :  255 - 0xff
    "11111111", -- 1669 - 0x685  :  255 - 0xff
    "00000000", -- 1670 - 0x686  :    0 - 0x0
    "00000000", -- 1671 - 0x687  :    0 - 0x0
    "00000000", -- 1672 - 0x688  :    0 - 0x0 -- plane 1
    "11111111", -- 1673 - 0x689  :  255 - 0xff
    "11111111", -- 1674 - 0x68a  :  255 - 0xff
    "11111111", -- 1675 - 0x68b  :  255 - 0xff
    "11001100", -- 1676 - 0x68c  :  204 - 0xcc
    "00000000", -- 1677 - 0x68d  :    0 - 0x0
    "00000000", -- 1678 - 0x68e  :    0 - 0x0
    "00000000", -- 1679 - 0x68f  :    0 - 0x0
    "11111110", -- 1680 - 0x690  :  254 - 0xfe -- Background 0x69
    "00000001", -- 1681 - 0x691  :    1 - 0x1
    "11001101", -- 1682 - 0x692  :  205 - 0xcd
    "00111110", -- 1683 - 0x693  :   62 - 0x3e
    "11111100", -- 1684 - 0x694  :  252 - 0xfc
    "11000000", -- 1685 - 0x695  :  192 - 0xc0
    "00000000", -- 1686 - 0x696  :    0 - 0x0
    "00000000", -- 1687 - 0x697  :    0 - 0x0
    "00000000", -- 1688 - 0x698  :    0 - 0x0 -- plane 1
    "11111110", -- 1689 - 0x699  :  254 - 0xfe
    "11111110", -- 1690 - 0x69a  :  254 - 0xfe
    "11110000", -- 1691 - 0x69b  :  240 - 0xf0
    "11000000", -- 1692 - 0x69c  :  192 - 0xc0
    "00000000", -- 1693 - 0x69d  :    0 - 0x0
    "00000000", -- 1694 - 0x69e  :    0 - 0x0
    "00000000", -- 1695 - 0x69f  :    0 - 0x0
    "00000000", -- 1696 - 0x6a0  :    0 - 0x0 -- Background 0x6a
    "00000000", -- 1697 - 0x6a1  :    0 - 0x0
    "00000000", -- 1698 - 0x6a2  :    0 - 0x0
    "00000000", -- 1699 - 0x6a3  :    0 - 0x0
    "00000000", -- 1700 - 0x6a4  :    0 - 0x0
    "00000000", -- 1701 - 0x6a5  :    0 - 0x0
    "00000000", -- 1702 - 0x6a6  :    0 - 0x0
    "00000000", -- 1703 - 0x6a7  :    0 - 0x0
    "00000000", -- 1704 - 0x6a8  :    0 - 0x0 -- plane 1
    "00000000", -- 1705 - 0x6a9  :    0 - 0x0
    "00000000", -- 1706 - 0x6aa  :    0 - 0x0
    "00000000", -- 1707 - 0x6ab  :    0 - 0x0
    "00000000", -- 1708 - 0x6ac  :    0 - 0x0
    "00000000", -- 1709 - 0x6ad  :    0 - 0x0
    "00000000", -- 1710 - 0x6ae  :    0 - 0x0
    "00000000", -- 1711 - 0x6af  :    0 - 0x0
    "01111111", -- 1712 - 0x6b0  :  127 - 0x7f -- Background 0x6b
    "11111111", -- 1713 - 0x6b1  :  255 - 0xff
    "11111111", -- 1714 - 0x6b2  :  255 - 0xff
    "11111111", -- 1715 - 0x6b3  :  255 - 0xff
    "01111111", -- 1716 - 0x6b4  :  127 - 0x7f
    "00110000", -- 1717 - 0x6b5  :   48 - 0x30
    "00001111", -- 1718 - 0x6b6  :   15 - 0xf
    "00000000", -- 1719 - 0x6b7  :    0 - 0x0
    "00111101", -- 1720 - 0x6b8  :   61 - 0x3d -- plane 1
    "01111111", -- 1721 - 0x6b9  :  127 - 0x7f
    "01111111", -- 1722 - 0x6ba  :  127 - 0x7f
    "01111111", -- 1723 - 0x6bb  :  127 - 0x7f
    "00111111", -- 1724 - 0x6bc  :   63 - 0x3f
    "00001111", -- 1725 - 0x6bd  :   15 - 0xf
    "00000000", -- 1726 - 0x6be  :    0 - 0x0
    "00000000", -- 1727 - 0x6bf  :    0 - 0x0
    "11111111", -- 1728 - 0x6c0  :  255 - 0xff -- Background 0x6c
    "11111111", -- 1729 - 0x6c1  :  255 - 0xff
    "11111111", -- 1730 - 0x6c2  :  255 - 0xff
    "11111111", -- 1731 - 0x6c3  :  255 - 0xff
    "11111111", -- 1732 - 0x6c4  :  255 - 0xff
    "11111110", -- 1733 - 0x6c5  :  254 - 0xfe
    "00000001", -- 1734 - 0x6c6  :    1 - 0x1
    "11111110", -- 1735 - 0x6c7  :  254 - 0xfe
    "11111111", -- 1736 - 0x6c8  :  255 - 0xff -- plane 1
    "11111111", -- 1737 - 0x6c9  :  255 - 0xff
    "11111111", -- 1738 - 0x6ca  :  255 - 0xff
    "11111111", -- 1739 - 0x6cb  :  255 - 0xff
    "11111111", -- 1740 - 0x6cc  :  255 - 0xff
    "11111111", -- 1741 - 0x6cd  :  255 - 0xff
    "11111110", -- 1742 - 0x6ce  :  254 - 0xfe
    "00000000", -- 1743 - 0x6cf  :    0 - 0x0
    "00000000", -- 1744 - 0x6d0  :    0 - 0x0 -- Background 0x6d
    "00000000", -- 1745 - 0x6d1  :    0 - 0x0
    "00000000", -- 1746 - 0x6d2  :    0 - 0x0
    "00000000", -- 1747 - 0x6d3  :    0 - 0x0
    "00000000", -- 1748 - 0x6d4  :    0 - 0x0
    "00000000", -- 1749 - 0x6d5  :    0 - 0x0
    "00000000", -- 1750 - 0x6d6  :    0 - 0x0
    "00000000", -- 1751 - 0x6d7  :    0 - 0x0
    "00000000", -- 1752 - 0x6d8  :    0 - 0x0 -- plane 1
    "00000000", -- 1753 - 0x6d9  :    0 - 0x0
    "00000000", -- 1754 - 0x6da  :    0 - 0x0
    "00000000", -- 1755 - 0x6db  :    0 - 0x0
    "00000000", -- 1756 - 0x6dc  :    0 - 0x0
    "00000000", -- 1757 - 0x6dd  :    0 - 0x0
    "00000000", -- 1758 - 0x6de  :    0 - 0x0
    "00000000", -- 1759 - 0x6df  :    0 - 0x0
    "00000000", -- 1760 - 0x6e0  :    0 - 0x0 -- Background 0x6e
    "00000000", -- 1761 - 0x6e1  :    0 - 0x0
    "00000000", -- 1762 - 0x6e2  :    0 - 0x0
    "00000000", -- 1763 - 0x6e3  :    0 - 0x0
    "00000000", -- 1764 - 0x6e4  :    0 - 0x0
    "00000000", -- 1765 - 0x6e5  :    0 - 0x0
    "00000000", -- 1766 - 0x6e6  :    0 - 0x0
    "00000000", -- 1767 - 0x6e7  :    0 - 0x0
    "00000000", -- 1768 - 0x6e8  :    0 - 0x0 -- plane 1
    "00000000", -- 1769 - 0x6e9  :    0 - 0x0
    "00000000", -- 1770 - 0x6ea  :    0 - 0x0
    "00000000", -- 1771 - 0x6eb  :    0 - 0x0
    "00000000", -- 1772 - 0x6ec  :    0 - 0x0
    "00000000", -- 1773 - 0x6ed  :    0 - 0x0
    "00000000", -- 1774 - 0x6ee  :    0 - 0x0
    "00000000", -- 1775 - 0x6ef  :    0 - 0x0
    "11111100", -- 1776 - 0x6f0  :  252 - 0xfc -- Background 0x6f
    "11111110", -- 1777 - 0x6f1  :  254 - 0xfe
    "11111111", -- 1778 - 0x6f2  :  255 - 0xff
    "11111111", -- 1779 - 0x6f3  :  255 - 0xff
    "11110010", -- 1780 - 0x6f4  :  242 - 0xf2
    "00001100", -- 1781 - 0x6f5  :   12 - 0xc
    "11110000", -- 1782 - 0x6f6  :  240 - 0xf0
    "00000000", -- 1783 - 0x6f7  :    0 - 0x0
    "10111000", -- 1784 - 0x6f8  :  184 - 0xb8 -- plane 1
    "11111100", -- 1785 - 0x6f9  :  252 - 0xfc
    "11111110", -- 1786 - 0x6fa  :  254 - 0xfe
    "11111110", -- 1787 - 0x6fb  :  254 - 0xfe
    "11111100", -- 1788 - 0x6fc  :  252 - 0xfc
    "11110000", -- 1789 - 0x6fd  :  240 - 0xf0
    "00000000", -- 1790 - 0x6fe  :    0 - 0x0
    "00000000", -- 1791 - 0x6ff  :    0 - 0x0
    "01111111", -- 1792 - 0x700  :  127 - 0x7f -- Background 0x70
    "11000000", -- 1793 - 0x701  :  192 - 0xc0
    "10000000", -- 1794 - 0x702  :  128 - 0x80
    "10000000", -- 1795 - 0x703  :  128 - 0x80
    "11100011", -- 1796 - 0x704  :  227 - 0xe3
    "11111111", -- 1797 - 0x705  :  255 - 0xff
    "11111111", -- 1798 - 0x706  :  255 - 0xff
    "11111111", -- 1799 - 0x707  :  255 - 0xff
    "00000000", -- 1800 - 0x708  :    0 - 0x0 -- plane 1
    "00111111", -- 1801 - 0x709  :   63 - 0x3f
    "01111111", -- 1802 - 0x70a  :  127 - 0x7f
    "01111111", -- 1803 - 0x70b  :  127 - 0x7f
    "00011100", -- 1804 - 0x70c  :   28 - 0x1c
    "00000000", -- 1805 - 0x70d  :    0 - 0x0
    "00000000", -- 1806 - 0x70e  :    0 - 0x0
    "00000000", -- 1807 - 0x70f  :    0 - 0x0
    "11111111", -- 1808 - 0x710  :  255 - 0xff -- Background 0x71
    "00000000", -- 1809 - 0x711  :    0 - 0x0
    "00000000", -- 1810 - 0x712  :    0 - 0x0
    "00000000", -- 1811 - 0x713  :    0 - 0x0
    "00000000", -- 1812 - 0x714  :    0 - 0x0
    "11000011", -- 1813 - 0x715  :  195 - 0xc3
    "11111111", -- 1814 - 0x716  :  255 - 0xff
    "11111111", -- 1815 - 0x717  :  255 - 0xff
    "00000000", -- 1816 - 0x718  :    0 - 0x0 -- plane 1
    "11111111", -- 1817 - 0x719  :  255 - 0xff
    "11111111", -- 1818 - 0x71a  :  255 - 0xff
    "11111111", -- 1819 - 0x71b  :  255 - 0xff
    "11111111", -- 1820 - 0x71c  :  255 - 0xff
    "00111100", -- 1821 - 0x71d  :   60 - 0x3c
    "00000000", -- 1822 - 0x71e  :    0 - 0x0
    "00000000", -- 1823 - 0x71f  :    0 - 0x0
    "11111110", -- 1824 - 0x720  :  254 - 0xfe -- Background 0x72
    "00000011", -- 1825 - 0x721  :    3 - 0x3
    "00000001", -- 1826 - 0x722  :    1 - 0x1
    "00000001", -- 1827 - 0x723  :    1 - 0x1
    "11000111", -- 1828 - 0x724  :  199 - 0xc7
    "11111111", -- 1829 - 0x725  :  255 - 0xff
    "11111111", -- 1830 - 0x726  :  255 - 0xff
    "11111111", -- 1831 - 0x727  :  255 - 0xff
    "00000000", -- 1832 - 0x728  :    0 - 0x0 -- plane 1
    "11111100", -- 1833 - 0x729  :  252 - 0xfc
    "11111110", -- 1834 - 0x72a  :  254 - 0xfe
    "11111110", -- 1835 - 0x72b  :  254 - 0xfe
    "00111000", -- 1836 - 0x72c  :   56 - 0x38
    "00000000", -- 1837 - 0x72d  :    0 - 0x0
    "00000000", -- 1838 - 0x72e  :    0 - 0x0
    "00000000", -- 1839 - 0x72f  :    0 - 0x0
    "11111111", -- 1840 - 0x730  :  255 - 0xff -- Background 0x73
    "11111111", -- 1841 - 0x731  :  255 - 0xff
    "11111111", -- 1842 - 0x732  :  255 - 0xff
    "11111111", -- 1843 - 0x733  :  255 - 0xff
    "11111111", -- 1844 - 0x734  :  255 - 0xff
    "11111111", -- 1845 - 0x735  :  255 - 0xff
    "11111111", -- 1846 - 0x736  :  255 - 0xff
    "11111111", -- 1847 - 0x737  :  255 - 0xff
    "11111111", -- 1848 - 0x738  :  255 - 0xff -- plane 1
    "11111111", -- 1849 - 0x739  :  255 - 0xff
    "11111101", -- 1850 - 0x73a  :  253 - 0xfd
    "11111111", -- 1851 - 0x73b  :  255 - 0xff
    "10111111", -- 1852 - 0x73c  :  191 - 0xbf
    "11111111", -- 1853 - 0x73d  :  255 - 0xff
    "11111111", -- 1854 - 0x73e  :  255 - 0xff
    "11110111", -- 1855 - 0x73f  :  247 - 0xf7
    "10111001", -- 1856 - 0x740  :  185 - 0xb9 -- Background 0x74
    "10010100", -- 1857 - 0x741  :  148 - 0x94
    "10001110", -- 1858 - 0x742  :  142 - 0x8e
    "11000101", -- 1859 - 0x743  :  197 - 0xc5
    "10010010", -- 1860 - 0x744  :  146 - 0x92
    "11000111", -- 1861 - 0x745  :  199 - 0xc7
    "11100010", -- 1862 - 0x746  :  226 - 0xe2
    "01111111", -- 1863 - 0x747  :  127 - 0x7f
    "01000110", -- 1864 - 0x748  :   70 - 0x46 -- plane 1
    "01101011", -- 1865 - 0x749  :  107 - 0x6b
    "01110001", -- 1866 - 0x74a  :  113 - 0x71
    "00111010", -- 1867 - 0x74b  :   58 - 0x3a
    "01101101", -- 1868 - 0x74c  :  109 - 0x6d
    "00111000", -- 1869 - 0x74d  :   56 - 0x38
    "00011101", -- 1870 - 0x74e  :   29 - 0x1d
    "00000000", -- 1871 - 0x74f  :    0 - 0x0
    "10111001", -- 1872 - 0x750  :  185 - 0xb9 -- Background 0x75
    "00010100", -- 1873 - 0x751  :   20 - 0x14
    "10001110", -- 1874 - 0x752  :  142 - 0x8e
    "11000101", -- 1875 - 0x753  :  197 - 0xc5
    "10010010", -- 1876 - 0x754  :  146 - 0x92
    "01000111", -- 1877 - 0x755  :   71 - 0x47
    "11100010", -- 1878 - 0x756  :  226 - 0xe2
    "11111111", -- 1879 - 0x757  :  255 - 0xff
    "01000110", -- 1880 - 0x758  :   70 - 0x46 -- plane 1
    "11101011", -- 1881 - 0x759  :  235 - 0xeb
    "01110001", -- 1882 - 0x75a  :  113 - 0x71
    "00111010", -- 1883 - 0x75b  :   58 - 0x3a
    "01101101", -- 1884 - 0x75c  :  109 - 0x6d
    "10111000", -- 1885 - 0x75d  :  184 - 0xb8
    "00011101", -- 1886 - 0x75e  :   29 - 0x1d
    "00000000", -- 1887 - 0x75f  :    0 - 0x0
    "10111001", -- 1888 - 0x760  :  185 - 0xb9 -- Background 0x76
    "00010101", -- 1889 - 0x761  :   21 - 0x15
    "10001111", -- 1890 - 0x762  :  143 - 0x8f
    "11000101", -- 1891 - 0x763  :  197 - 0xc5
    "10010011", -- 1892 - 0x764  :  147 - 0x93
    "01000111", -- 1893 - 0x765  :   71 - 0x47
    "11100011", -- 1894 - 0x766  :  227 - 0xe3
    "11111110", -- 1895 - 0x767  :  254 - 0xfe
    "01000110", -- 1896 - 0x768  :   70 - 0x46 -- plane 1
    "11101010", -- 1897 - 0x769  :  234 - 0xea
    "01110000", -- 1898 - 0x76a  :  112 - 0x70
    "00111010", -- 1899 - 0x76b  :   58 - 0x3a
    "01101100", -- 1900 - 0x76c  :  108 - 0x6c
    "10111000", -- 1901 - 0x76d  :  184 - 0xb8
    "00011100", -- 1902 - 0x76e  :   28 - 0x1c
    "00000000", -- 1903 - 0x76f  :    0 - 0x0
    "11111111", -- 1904 - 0x770  :  255 - 0xff -- Background 0x77
    "11111111", -- 1905 - 0x771  :  255 - 0xff
    "11111111", -- 1906 - 0x772  :  255 - 0xff
    "11111111", -- 1907 - 0x773  :  255 - 0xff
    "11111111", -- 1908 - 0x774  :  255 - 0xff
    "11111111", -- 1909 - 0x775  :  255 - 0xff
    "11111111", -- 1910 - 0x776  :  255 - 0xff
    "11111111", -- 1911 - 0x777  :  255 - 0xff
    "10000001", -- 1912 - 0x778  :  129 - 0x81 -- plane 1
    "11111111", -- 1913 - 0x779  :  255 - 0xff
    "11111101", -- 1914 - 0x77a  :  253 - 0xfd
    "11111111", -- 1915 - 0x77b  :  255 - 0xff
    "10111111", -- 1916 - 0x77c  :  191 - 0xbf
    "11111111", -- 1917 - 0x77d  :  255 - 0xff
    "11111111", -- 1918 - 0x77e  :  255 - 0xff
    "11110111", -- 1919 - 0x77f  :  247 - 0xf7
    "00000000", -- 1920 - 0x780  :    0 - 0x0 -- Background 0x78
    "00000000", -- 1921 - 0x781  :    0 - 0x0
    "00000000", -- 1922 - 0x782  :    0 - 0x0
    "00000000", -- 1923 - 0x783  :    0 - 0x0
    "00000000", -- 1924 - 0x784  :    0 - 0x0
    "00000000", -- 1925 - 0x785  :    0 - 0x0
    "00000000", -- 1926 - 0x786  :    0 - 0x0
    "00000000", -- 1927 - 0x787  :    0 - 0x0
    "00000000", -- 1928 - 0x788  :    0 - 0x0 -- plane 1
    "00000000", -- 1929 - 0x789  :    0 - 0x0
    "00000000", -- 1930 - 0x78a  :    0 - 0x0
    "00000000", -- 1931 - 0x78b  :    0 - 0x0
    "00000000", -- 1932 - 0x78c  :    0 - 0x0
    "00000000", -- 1933 - 0x78d  :    0 - 0x0
    "00000000", -- 1934 - 0x78e  :    0 - 0x0
    "00000000", -- 1935 - 0x78f  :    0 - 0x0
    "00000000", -- 1936 - 0x790  :    0 - 0x0 -- Background 0x79
    "00000000", -- 1937 - 0x791  :    0 - 0x0
    "00000000", -- 1938 - 0x792  :    0 - 0x0
    "00000000", -- 1939 - 0x793  :    0 - 0x0
    "00000000", -- 1940 - 0x794  :    0 - 0x0
    "00000000", -- 1941 - 0x795  :    0 - 0x0
    "00000000", -- 1942 - 0x796  :    0 - 0x0
    "00000000", -- 1943 - 0x797  :    0 - 0x0
    "00000000", -- 1944 - 0x798  :    0 - 0x0 -- plane 1
    "00000000", -- 1945 - 0x799  :    0 - 0x0
    "00000000", -- 1946 - 0x79a  :    0 - 0x0
    "00000000", -- 1947 - 0x79b  :    0 - 0x0
    "00000000", -- 1948 - 0x79c  :    0 - 0x0
    "00000000", -- 1949 - 0x79d  :    0 - 0x0
    "00000000", -- 1950 - 0x79e  :    0 - 0x0
    "00000000", -- 1951 - 0x79f  :    0 - 0x0
    "00000000", -- 1952 - 0x7a0  :    0 - 0x0 -- Background 0x7a
    "00000000", -- 1953 - 0x7a1  :    0 - 0x0
    "00000000", -- 1954 - 0x7a2  :    0 - 0x0
    "00000000", -- 1955 - 0x7a3  :    0 - 0x0
    "00000000", -- 1956 - 0x7a4  :    0 - 0x0
    "00000000", -- 1957 - 0x7a5  :    0 - 0x0
    "00000000", -- 1958 - 0x7a6  :    0 - 0x0
    "00000000", -- 1959 - 0x7a7  :    0 - 0x0
    "00000000", -- 1960 - 0x7a8  :    0 - 0x0 -- plane 1
    "00000000", -- 1961 - 0x7a9  :    0 - 0x0
    "00000000", -- 1962 - 0x7aa  :    0 - 0x0
    "00000000", -- 1963 - 0x7ab  :    0 - 0x0
    "00000000", -- 1964 - 0x7ac  :    0 - 0x0
    "00000000", -- 1965 - 0x7ad  :    0 - 0x0
    "00000000", -- 1966 - 0x7ae  :    0 - 0x0
    "00000000", -- 1967 - 0x7af  :    0 - 0x0
    "00000000", -- 1968 - 0x7b0  :    0 - 0x0 -- Background 0x7b
    "00000000", -- 1969 - 0x7b1  :    0 - 0x0
    "00000000", -- 1970 - 0x7b2  :    0 - 0x0
    "00000000", -- 1971 - 0x7b3  :    0 - 0x0
    "00000000", -- 1972 - 0x7b4  :    0 - 0x0
    "00000000", -- 1973 - 0x7b5  :    0 - 0x0
    "00000000", -- 1974 - 0x7b6  :    0 - 0x0
    "00000000", -- 1975 - 0x7b7  :    0 - 0x0
    "00000000", -- 1976 - 0x7b8  :    0 - 0x0 -- plane 1
    "00000000", -- 1977 - 0x7b9  :    0 - 0x0
    "00000000", -- 1978 - 0x7ba  :    0 - 0x0
    "00000000", -- 1979 - 0x7bb  :    0 - 0x0
    "00000000", -- 1980 - 0x7bc  :    0 - 0x0
    "00000000", -- 1981 - 0x7bd  :    0 - 0x0
    "00000000", -- 1982 - 0x7be  :    0 - 0x0
    "00000000", -- 1983 - 0x7bf  :    0 - 0x0
    "00100010", -- 1984 - 0x7c0  :   34 - 0x22 -- Background 0x7c
    "01010101", -- 1985 - 0x7c1  :   85 - 0x55
    "10101010", -- 1986 - 0x7c2  :  170 - 0xaa
    "00000101", -- 1987 - 0x7c3  :    5 - 0x5
    "00000100", -- 1988 - 0x7c4  :    4 - 0x4
    "00001010", -- 1989 - 0x7c5  :   10 - 0xa
    "01010000", -- 1990 - 0x7c6  :   80 - 0x50
    "00000010", -- 1991 - 0x7c7  :    2 - 0x2
    "00000000", -- 1992 - 0x7c8  :    0 - 0x0 -- plane 1
    "00100010", -- 1993 - 0x7c9  :   34 - 0x22
    "01110111", -- 1994 - 0x7ca  :  119 - 0x77
    "11111111", -- 1995 - 0x7cb  :  255 - 0xff
    "11111011", -- 1996 - 0x7cc  :  251 - 0xfb
    "11110101", -- 1997 - 0x7cd  :  245 - 0xf5
    "11101111", -- 1998 - 0x7ce  :  239 - 0xef
    "11111111", -- 1999 - 0x7cf  :  255 - 0xff
    "01110011", -- 2000 - 0x7d0  :  115 - 0x73 -- Background 0x7d
    "11111111", -- 2001 - 0x7d1  :  255 - 0xff
    "11111111", -- 2002 - 0x7d2  :  255 - 0xff
    "10111101", -- 2003 - 0x7d3  :  189 - 0xbd
    "01101110", -- 2004 - 0x7d4  :  110 - 0x6e
    "00001010", -- 2005 - 0x7d5  :   10 - 0xa
    "01010000", -- 2006 - 0x7d6  :   80 - 0x50
    "00000010", -- 2007 - 0x7d7  :    2 - 0x2
    "00000000", -- 2008 - 0x7d8  :    0 - 0x0 -- plane 1
    "01110011", -- 2009 - 0x7d9  :  115 - 0x73
    "11111111", -- 2010 - 0x7da  :  255 - 0xff
    "11111111", -- 2011 - 0x7db  :  255 - 0xff
    "11111011", -- 2012 - 0x7dc  :  251 - 0xfb
    "11111101", -- 2013 - 0x7dd  :  253 - 0xfd
    "11101111", -- 2014 - 0x7de  :  239 - 0xef
    "11111111", -- 2015 - 0x7df  :  255 - 0xff
    "00100000", -- 2016 - 0x7e0  :   32 - 0x20 -- Background 0x7e
    "01010000", -- 2017 - 0x7e1  :   80 - 0x50
    "10000100", -- 2018 - 0x7e2  :  132 - 0x84
    "00000000", -- 2019 - 0x7e3  :    0 - 0x0
    "00100100", -- 2020 - 0x7e4  :   36 - 0x24
    "01011010", -- 2021 - 0x7e5  :   90 - 0x5a
    "00010000", -- 2022 - 0x7e6  :   16 - 0x10
    "00000000", -- 2023 - 0x7e7  :    0 - 0x0
    "11011111", -- 2024 - 0x7e8  :  223 - 0xdf -- plane 1
    "10101111", -- 2025 - 0x7e9  :  175 - 0xaf
    "01111111", -- 2026 - 0x7ea  :  127 - 0x7f
    "11111111", -- 2027 - 0x7eb  :  255 - 0xff
    "11111011", -- 2028 - 0x7ec  :  251 - 0xfb
    "11110101", -- 2029 - 0x7ed  :  245 - 0xf5
    "11101111", -- 2030 - 0x7ee  :  239 - 0xef
    "11111111", -- 2031 - 0x7ef  :  255 - 0xff
    "11111111", -- 2032 - 0x7f0  :  255 - 0xff -- Background 0x7f
    "01010000", -- 2033 - 0x7f1  :   80 - 0x50
    "10000100", -- 2034 - 0x7f2  :  132 - 0x84
    "00000000", -- 2035 - 0x7f3  :    0 - 0x0
    "00100100", -- 2036 - 0x7f4  :   36 - 0x24
    "01011010", -- 2037 - 0x7f5  :   90 - 0x5a
    "00010000", -- 2038 - 0x7f6  :   16 - 0x10
    "00000000", -- 2039 - 0x7f7  :    0 - 0x0
    "00000000", -- 2040 - 0x7f8  :    0 - 0x0 -- plane 1
    "10101111", -- 2041 - 0x7f9  :  175 - 0xaf
    "01111111", -- 2042 - 0x7fa  :  127 - 0x7f
    "11111111", -- 2043 - 0x7fb  :  255 - 0xff
    "11111011", -- 2044 - 0x7fc  :  251 - 0xfb
    "11110101", -- 2045 - 0x7fd  :  245 - 0xf5
    "11101111", -- 2046 - 0x7fe  :  239 - 0xef
    "11111111", -- 2047 - 0x7ff  :  255 - 0xff
    "11111111", -- 2048 - 0x800  :  255 - 0xff -- Background 0x80
    "10000000", -- 2049 - 0x801  :  128 - 0x80
    "11001111", -- 2050 - 0x802  :  207 - 0xcf
    "01001000", -- 2051 - 0x803  :   72 - 0x48
    "11001111", -- 2052 - 0x804  :  207 - 0xcf
    "10000000", -- 2053 - 0x805  :  128 - 0x80
    "11001111", -- 2054 - 0x806  :  207 - 0xcf
    "01001000", -- 2055 - 0x807  :   72 - 0x48
    "00000000", -- 2056 - 0x808  :    0 - 0x0 -- plane 1
    "01111111", -- 2057 - 0x809  :  127 - 0x7f
    "00110000", -- 2058 - 0x80a  :   48 - 0x30
    "00110000", -- 2059 - 0x80b  :   48 - 0x30
    "00110000", -- 2060 - 0x80c  :   48 - 0x30
    "01111111", -- 2061 - 0x80d  :  127 - 0x7f
    "00110000", -- 2062 - 0x80e  :   48 - 0x30
    "00110000", -- 2063 - 0x80f  :   48 - 0x30
    "11111111", -- 2064 - 0x810  :  255 - 0xff -- Background 0x81
    "10000000", -- 2065 - 0x811  :  128 - 0x80
    "11111111", -- 2066 - 0x812  :  255 - 0xff
    "10000000", -- 2067 - 0x813  :  128 - 0x80
    "10000000", -- 2068 - 0x814  :  128 - 0x80
    "11011111", -- 2069 - 0x815  :  223 - 0xdf
    "10110000", -- 2070 - 0x816  :  176 - 0xb0
    "11000000", -- 2071 - 0x817  :  192 - 0xc0
    "00000000", -- 2072 - 0x818  :    0 - 0x0 -- plane 1
    "01111111", -- 2073 - 0x819  :  127 - 0x7f
    "00000000", -- 2074 - 0x81a  :    0 - 0x0
    "01111111", -- 2075 - 0x81b  :  127 - 0x7f
    "01111111", -- 2076 - 0x81c  :  127 - 0x7f
    "00100000", -- 2077 - 0x81d  :   32 - 0x20
    "01000000", -- 2078 - 0x81e  :   64 - 0x40
    "00000000", -- 2079 - 0x81f  :    0 - 0x0
    "11111111", -- 2080 - 0x820  :  255 - 0xff -- Background 0x82
    "00000001", -- 2081 - 0x821  :    1 - 0x1
    "11110011", -- 2082 - 0x822  :  243 - 0xf3
    "00010010", -- 2083 - 0x823  :   18 - 0x12
    "11110011", -- 2084 - 0x824  :  243 - 0xf3
    "00000001", -- 2085 - 0x825  :    1 - 0x1
    "11110011", -- 2086 - 0x826  :  243 - 0xf3
    "00010010", -- 2087 - 0x827  :   18 - 0x12
    "00000000", -- 2088 - 0x828  :    0 - 0x0 -- plane 1
    "11111110", -- 2089 - 0x829  :  254 - 0xfe
    "00001100", -- 2090 - 0x82a  :   12 - 0xc
    "00001100", -- 2091 - 0x82b  :   12 - 0xc
    "00001100", -- 2092 - 0x82c  :   12 - 0xc
    "11111110", -- 2093 - 0x82d  :  254 - 0xfe
    "00001100", -- 2094 - 0x82e  :   12 - 0xc
    "00001100", -- 2095 - 0x82f  :   12 - 0xc
    "11111111", -- 2096 - 0x830  :  255 - 0xff -- Background 0x83
    "00000000", -- 2097 - 0x831  :    0 - 0x0
    "11111111", -- 2098 - 0x832  :  255 - 0xff
    "00000000", -- 2099 - 0x833  :    0 - 0x0
    "00000000", -- 2100 - 0x834  :    0 - 0x0
    "11111111", -- 2101 - 0x835  :  255 - 0xff
    "00000000", -- 2102 - 0x836  :    0 - 0x0
    "00000000", -- 2103 - 0x837  :    0 - 0x0
    "00000000", -- 2104 - 0x838  :    0 - 0x0 -- plane 1
    "11111111", -- 2105 - 0x839  :  255 - 0xff
    "00000000", -- 2106 - 0x83a  :    0 - 0x0
    "11111111", -- 2107 - 0x83b  :  255 - 0xff
    "11111111", -- 2108 - 0x83c  :  255 - 0xff
    "00000000", -- 2109 - 0x83d  :    0 - 0x0
    "00000000", -- 2110 - 0x83e  :    0 - 0x0
    "00000000", -- 2111 - 0x83f  :    0 - 0x0
    "11111111", -- 2112 - 0x840  :  255 - 0xff -- Background 0x84
    "10000010", -- 2113 - 0x841  :  130 - 0x82
    "00010000", -- 2114 - 0x842  :   16 - 0x10
    "00000000", -- 2115 - 0x843  :    0 - 0x0
    "00000000", -- 2116 - 0x844  :    0 - 0x0
    "00010000", -- 2117 - 0x845  :   16 - 0x10
    "01000100", -- 2118 - 0x846  :   68 - 0x44
    "11111111", -- 2119 - 0x847  :  255 - 0xff
    "00000000", -- 2120 - 0x848  :    0 - 0x0 -- plane 1
    "11111111", -- 2121 - 0x849  :  255 - 0xff
    "11111111", -- 2122 - 0x84a  :  255 - 0xff
    "11111111", -- 2123 - 0x84b  :  255 - 0xff
    "11111111", -- 2124 - 0x84c  :  255 - 0xff
    "11101111", -- 2125 - 0x84d  :  239 - 0xef
    "10111011", -- 2126 - 0x84e  :  187 - 0xbb
    "00000000", -- 2127 - 0x84f  :    0 - 0x0
    "11111111", -- 2128 - 0x850  :  255 - 0xff -- Background 0x85
    "00000001", -- 2129 - 0x851  :    1 - 0x1
    "11111111", -- 2130 - 0x852  :  255 - 0xff
    "00000001", -- 2131 - 0x853  :    1 - 0x1
    "00000001", -- 2132 - 0x854  :    1 - 0x1
    "11110011", -- 2133 - 0x855  :  243 - 0xf3
    "00001101", -- 2134 - 0x856  :   13 - 0xd
    "00000011", -- 2135 - 0x857  :    3 - 0x3
    "00000000", -- 2136 - 0x858  :    0 - 0x0 -- plane 1
    "11111110", -- 2137 - 0x859  :  254 - 0xfe
    "00000000", -- 2138 - 0x85a  :    0 - 0x0
    "11111110", -- 2139 - 0x85b  :  254 - 0xfe
    "11111110", -- 2140 - 0x85c  :  254 - 0xfe
    "00001100", -- 2141 - 0x85d  :   12 - 0xc
    "00000010", -- 2142 - 0x85e  :    2 - 0x2
    "00000000", -- 2143 - 0x85f  :    0 - 0x0
    "00000000", -- 2144 - 0x860  :    0 - 0x0 -- Background 0x86
    "00000000", -- 2145 - 0x861  :    0 - 0x0
    "00000000", -- 2146 - 0x862  :    0 - 0x0
    "00000000", -- 2147 - 0x863  :    0 - 0x0
    "00000000", -- 2148 - 0x864  :    0 - 0x0
    "00000000", -- 2149 - 0x865  :    0 - 0x0
    "00000000", -- 2150 - 0x866  :    0 - 0x0
    "00000000", -- 2151 - 0x867  :    0 - 0x0
    "00000000", -- 2152 - 0x868  :    0 - 0x0 -- plane 1
    "00000000", -- 2153 - 0x869  :    0 - 0x0
    "00000000", -- 2154 - 0x86a  :    0 - 0x0
    "00000000", -- 2155 - 0x86b  :    0 - 0x0
    "00000000", -- 2156 - 0x86c  :    0 - 0x0
    "00000000", -- 2157 - 0x86d  :    0 - 0x0
    "00000000", -- 2158 - 0x86e  :    0 - 0x0
    "00000000", -- 2159 - 0x86f  :    0 - 0x0
    "00000000", -- 2160 - 0x870  :    0 - 0x0 -- Background 0x87
    "00000000", -- 2161 - 0x871  :    0 - 0x0
    "00000000", -- 2162 - 0x872  :    0 - 0x0
    "00000000", -- 2163 - 0x873  :    0 - 0x0
    "00000000", -- 2164 - 0x874  :    0 - 0x0
    "00000000", -- 2165 - 0x875  :    0 - 0x0
    "00000000", -- 2166 - 0x876  :    0 - 0x0
    "00000000", -- 2167 - 0x877  :    0 - 0x0
    "00000000", -- 2168 - 0x878  :    0 - 0x0 -- plane 1
    "00000000", -- 2169 - 0x879  :    0 - 0x0
    "00000000", -- 2170 - 0x87a  :    0 - 0x0
    "00000000", -- 2171 - 0x87b  :    0 - 0x0
    "00000000", -- 2172 - 0x87c  :    0 - 0x0
    "00000000", -- 2173 - 0x87d  :    0 - 0x0
    "00000000", -- 2174 - 0x87e  :    0 - 0x0
    "00000000", -- 2175 - 0x87f  :    0 - 0x0
    "00000111", -- 2176 - 0x880  :    7 - 0x7 -- Background 0x88
    "00011110", -- 2177 - 0x881  :   30 - 0x1e
    "00101111", -- 2178 - 0x882  :   47 - 0x2f
    "01010011", -- 2179 - 0x883  :   83 - 0x53
    "01101110", -- 2180 - 0x884  :  110 - 0x6e
    "11011011", -- 2181 - 0x885  :  219 - 0xdb
    "11111010", -- 2182 - 0x886  :  250 - 0xfa
    "11010101", -- 2183 - 0x887  :  213 - 0xd5
    "00000000", -- 2184 - 0x888  :    0 - 0x0 -- plane 1
    "00000111", -- 2185 - 0x889  :    7 - 0x7
    "00011111", -- 2186 - 0x88a  :   31 - 0x1f
    "00111100", -- 2187 - 0x88b  :   60 - 0x3c
    "00110001", -- 2188 - 0x88c  :   49 - 0x31
    "01110100", -- 2189 - 0x88d  :  116 - 0x74
    "01100101", -- 2190 - 0x88e  :  101 - 0x65
    "01101010", -- 2191 - 0x88f  :  106 - 0x6a
    "10111011", -- 2192 - 0x890  :  187 - 0xbb -- Background 0x89
    "11110010", -- 2193 - 0x891  :  242 - 0xf2
    "11011101", -- 2194 - 0x892  :  221 - 0xdd
    "01001111", -- 2195 - 0x893  :   79 - 0x4f
    "01111011", -- 2196 - 0x894  :  123 - 0x7b
    "00110010", -- 2197 - 0x895  :   50 - 0x32
    "00011111", -- 2198 - 0x896  :   31 - 0x1f
    "00000111", -- 2199 - 0x897  :    7 - 0x7
    "01100100", -- 2200 - 0x898  :  100 - 0x64 -- plane 1
    "01101101", -- 2201 - 0x899  :  109 - 0x6d
    "01110010", -- 2202 - 0x89a  :  114 - 0x72
    "00110000", -- 2203 - 0x89b  :   48 - 0x30
    "00111100", -- 2204 - 0x89c  :   60 - 0x3c
    "00011111", -- 2205 - 0x89d  :   31 - 0x1f
    "00000111", -- 2206 - 0x89e  :    7 - 0x7
    "00000000", -- 2207 - 0x89f  :    0 - 0x0
    "11100000", -- 2208 - 0x8a0  :  224 - 0xe0 -- Background 0x8a
    "11011000", -- 2209 - 0x8a1  :  216 - 0xd8
    "01010100", -- 2210 - 0x8a2  :   84 - 0x54
    "11101010", -- 2211 - 0x8a3  :  234 - 0xea
    "10111010", -- 2212 - 0x8a4  :  186 - 0xba
    "10010011", -- 2213 - 0x8a5  :  147 - 0x93
    "11011111", -- 2214 - 0x8a6  :  223 - 0xdf
    "10111101", -- 2215 - 0x8a7  :  189 - 0xbd
    "00000000", -- 2216 - 0x8a8  :    0 - 0x0 -- plane 1
    "11100000", -- 2217 - 0x8a9  :  224 - 0xe0
    "11111000", -- 2218 - 0x8aa  :  248 - 0xf8
    "00111100", -- 2219 - 0x8ab  :   60 - 0x3c
    "01001100", -- 2220 - 0x8ac  :   76 - 0x4c
    "01101110", -- 2221 - 0x8ad  :  110 - 0x6e
    "00100110", -- 2222 - 0x8ae  :   38 - 0x26
    "01000110", -- 2223 - 0x8af  :   70 - 0x46
    "01101011", -- 2224 - 0x8b0  :  107 - 0x6b -- Background 0x8b
    "10011111", -- 2225 - 0x8b1  :  159 - 0x9f
    "01011101", -- 2226 - 0x8b2  :   93 - 0x5d
    "10110110", -- 2227 - 0x8b3  :  182 - 0xb6
    "11101010", -- 2228 - 0x8b4  :  234 - 0xea
    "11001100", -- 2229 - 0x8b5  :  204 - 0xcc
    "01111000", -- 2230 - 0x8b6  :  120 - 0x78
    "11100000", -- 2231 - 0x8b7  :  224 - 0xe0
    "10010110", -- 2232 - 0x8b8  :  150 - 0x96 -- plane 1
    "01100110", -- 2233 - 0x8b9  :  102 - 0x66
    "10101110", -- 2234 - 0x8ba  :  174 - 0xae
    "01001100", -- 2235 - 0x8bb  :   76 - 0x4c
    "00111100", -- 2236 - 0x8bc  :   60 - 0x3c
    "11111000", -- 2237 - 0x8bd  :  248 - 0xf8
    "11100000", -- 2238 - 0x8be  :  224 - 0xe0
    "00000000", -- 2239 - 0x8bf  :    0 - 0x0
    "00000111", -- 2240 - 0x8c0  :    7 - 0x7 -- Background 0x8c
    "00011000", -- 2241 - 0x8c1  :   24 - 0x18
    "00100011", -- 2242 - 0x8c2  :   35 - 0x23
    "01001100", -- 2243 - 0x8c3  :   76 - 0x4c
    "01110000", -- 2244 - 0x8c4  :  112 - 0x70
    "10100001", -- 2245 - 0x8c5  :  161 - 0xa1
    "10100110", -- 2246 - 0x8c6  :  166 - 0xa6
    "10101000", -- 2247 - 0x8c7  :  168 - 0xa8
    "00000000", -- 2248 - 0x8c8  :    0 - 0x0 -- plane 1
    "00000111", -- 2249 - 0x8c9  :    7 - 0x7
    "00011111", -- 2250 - 0x8ca  :   31 - 0x1f
    "00111111", -- 2251 - 0x8cb  :   63 - 0x3f
    "00111111", -- 2252 - 0x8cc  :   63 - 0x3f
    "01111111", -- 2253 - 0x8cd  :  127 - 0x7f
    "01111111", -- 2254 - 0x8ce  :  127 - 0x7f
    "01111111", -- 2255 - 0x8cf  :  127 - 0x7f
    "10100101", -- 2256 - 0x8d0  :  165 - 0xa5 -- Background 0x8d
    "10100010", -- 2257 - 0x8d1  :  162 - 0xa2
    "10010000", -- 2258 - 0x8d2  :  144 - 0x90
    "01001000", -- 2259 - 0x8d3  :   72 - 0x48
    "01000111", -- 2260 - 0x8d4  :   71 - 0x47
    "00100000", -- 2261 - 0x8d5  :   32 - 0x20
    "00011001", -- 2262 - 0x8d6  :   25 - 0x19
    "00000111", -- 2263 - 0x8d7  :    7 - 0x7
    "01111111", -- 2264 - 0x8d8  :  127 - 0x7f -- plane 1
    "01111111", -- 2265 - 0x8d9  :  127 - 0x7f
    "01111111", -- 2266 - 0x8da  :  127 - 0x7f
    "00111111", -- 2267 - 0x8db  :   63 - 0x3f
    "00111111", -- 2268 - 0x8dc  :   63 - 0x3f
    "00011111", -- 2269 - 0x8dd  :   31 - 0x1f
    "00000111", -- 2270 - 0x8de  :    7 - 0x7
    "00000000", -- 2271 - 0x8df  :    0 - 0x0
    "11100000", -- 2272 - 0x8e0  :  224 - 0xe0 -- Background 0x8e
    "00011000", -- 2273 - 0x8e1  :   24 - 0x18
    "00000100", -- 2274 - 0x8e2  :    4 - 0x4
    "11000010", -- 2275 - 0x8e3  :  194 - 0xc2
    "00110010", -- 2276 - 0x8e4  :   50 - 0x32
    "00001001", -- 2277 - 0x8e5  :    9 - 0x9
    "11000101", -- 2278 - 0x8e6  :  197 - 0xc5
    "00100101", -- 2279 - 0x8e7  :   37 - 0x25
    "00000000", -- 2280 - 0x8e8  :    0 - 0x0 -- plane 1
    "11100000", -- 2281 - 0x8e9  :  224 - 0xe0
    "11111000", -- 2282 - 0x8ea  :  248 - 0xf8
    "11111100", -- 2283 - 0x8eb  :  252 - 0xfc
    "11111100", -- 2284 - 0x8ec  :  252 - 0xfc
    "11111110", -- 2285 - 0x8ed  :  254 - 0xfe
    "11111110", -- 2286 - 0x8ee  :  254 - 0xfe
    "11111110", -- 2287 - 0x8ef  :  254 - 0xfe
    "10100101", -- 2288 - 0x8f0  :  165 - 0xa5 -- Background 0x8f
    "01100101", -- 2289 - 0x8f1  :  101 - 0x65
    "01000101", -- 2290 - 0x8f2  :   69 - 0x45
    "10001010", -- 2291 - 0x8f3  :  138 - 0x8a
    "10010010", -- 2292 - 0x8f4  :  146 - 0x92
    "00100100", -- 2293 - 0x8f5  :   36 - 0x24
    "11011000", -- 2294 - 0x8f6  :  216 - 0xd8
    "11100000", -- 2295 - 0x8f7  :  224 - 0xe0
    "11111110", -- 2296 - 0x8f8  :  254 - 0xfe -- plane 1
    "11111110", -- 2297 - 0x8f9  :  254 - 0xfe
    "11111110", -- 2298 - 0x8fa  :  254 - 0xfe
    "11111100", -- 2299 - 0x8fb  :  252 - 0xfc
    "11111100", -- 2300 - 0x8fc  :  252 - 0xfc
    "11111000", -- 2301 - 0x8fd  :  248 - 0xf8
    "11100000", -- 2302 - 0x8fe  :  224 - 0xe0
    "00000000", -- 2303 - 0x8ff  :    0 - 0x0
    "00000000", -- 2304 - 0x900  :    0 - 0x0 -- Background 0x90
    "00000000", -- 2305 - 0x901  :    0 - 0x0
    "00100000", -- 2306 - 0x902  :   32 - 0x20
    "00110000", -- 2307 - 0x903  :   48 - 0x30
    "00101100", -- 2308 - 0x904  :   44 - 0x2c
    "00100010", -- 2309 - 0x905  :   34 - 0x22
    "00010001", -- 2310 - 0x906  :   17 - 0x11
    "00001000", -- 2311 - 0x907  :    8 - 0x8
    "00000000", -- 2312 - 0x908  :    0 - 0x0 -- plane 1
    "00000000", -- 2313 - 0x909  :    0 - 0x0
    "00000000", -- 2314 - 0x90a  :    0 - 0x0
    "00000000", -- 2315 - 0x90b  :    0 - 0x0
    "00010000", -- 2316 - 0x90c  :   16 - 0x10
    "00011100", -- 2317 - 0x90d  :   28 - 0x1c
    "00001110", -- 2318 - 0x90e  :   14 - 0xe
    "00000111", -- 2319 - 0x90f  :    7 - 0x7
    "00000100", -- 2320 - 0x910  :    4 - 0x4 -- Background 0x91
    "11110010", -- 2321 - 0x911  :  242 - 0xf2
    "11001111", -- 2322 - 0x912  :  207 - 0xcf
    "00110000", -- 2323 - 0x913  :   48 - 0x30
    "00001100", -- 2324 - 0x914  :   12 - 0xc
    "11111111", -- 2325 - 0x915  :  255 - 0xff
    "10000000", -- 2326 - 0x916  :  128 - 0x80
    "11111111", -- 2327 - 0x917  :  255 - 0xff
    "00000011", -- 2328 - 0x918  :    3 - 0x3 -- plane 1
    "00000001", -- 2329 - 0x919  :    1 - 0x1
    "00110000", -- 2330 - 0x91a  :   48 - 0x30
    "00001111", -- 2331 - 0x91b  :   15 - 0xf
    "00000011", -- 2332 - 0x91c  :    3 - 0x3
    "00000000", -- 2333 - 0x91d  :    0 - 0x0
    "01111111", -- 2334 - 0x91e  :  127 - 0x7f
    "00000000", -- 2335 - 0x91f  :    0 - 0x0
    "01000010", -- 2336 - 0x920  :   66 - 0x42 -- Background 0x92
    "10100101", -- 2337 - 0x921  :  165 - 0xa5
    "10100101", -- 2338 - 0x922  :  165 - 0xa5
    "10011001", -- 2339 - 0x923  :  153 - 0x99
    "10011001", -- 2340 - 0x924  :  153 - 0x99
    "10011001", -- 2341 - 0x925  :  153 - 0x99
    "00000001", -- 2342 - 0x926  :    1 - 0x1
    "00000000", -- 2343 - 0x927  :    0 - 0x0
    "00000000", -- 2344 - 0x928  :    0 - 0x0 -- plane 1
    "01000010", -- 2345 - 0x929  :   66 - 0x42
    "01000010", -- 2346 - 0x92a  :   66 - 0x42
    "01100110", -- 2347 - 0x92b  :  102 - 0x66
    "01100110", -- 2348 - 0x92c  :  102 - 0x66
    "01100110", -- 2349 - 0x92d  :  102 - 0x66
    "11111110", -- 2350 - 0x92e  :  254 - 0xfe
    "11111111", -- 2351 - 0x92f  :  255 - 0xff
    "11111111", -- 2352 - 0x930  :  255 - 0xff -- Background 0x93
    "11111111", -- 2353 - 0x931  :  255 - 0xff
    "11111111", -- 2354 - 0x932  :  255 - 0xff
    "10000001", -- 2355 - 0x933  :  129 - 0x81
    "11111111", -- 2356 - 0x934  :  255 - 0xff
    "11111111", -- 2357 - 0x935  :  255 - 0xff
    "11111111", -- 2358 - 0x936  :  255 - 0xff
    "10000001", -- 2359 - 0x937  :  129 - 0x81
    "01111110", -- 2360 - 0x938  :  126 - 0x7e -- plane 1
    "01111110", -- 2361 - 0x939  :  126 - 0x7e
    "01111110", -- 2362 - 0x93a  :  126 - 0x7e
    "01111110", -- 2363 - 0x93b  :  126 - 0x7e
    "01111110", -- 2364 - 0x93c  :  126 - 0x7e
    "01111110", -- 2365 - 0x93d  :  126 - 0x7e
    "01111110", -- 2366 - 0x93e  :  126 - 0x7e
    "01111110", -- 2367 - 0x93f  :  126 - 0x7e
    "00000000", -- 2368 - 0x940  :    0 - 0x0 -- Background 0x94
    "00000000", -- 2369 - 0x941  :    0 - 0x0
    "00000100", -- 2370 - 0x942  :    4 - 0x4
    "00001100", -- 2371 - 0x943  :   12 - 0xc
    "00110100", -- 2372 - 0x944  :   52 - 0x34
    "01000100", -- 2373 - 0x945  :   68 - 0x44
    "10001000", -- 2374 - 0x946  :  136 - 0x88
    "00010000", -- 2375 - 0x947  :   16 - 0x10
    "00000000", -- 2376 - 0x948  :    0 - 0x0 -- plane 1
    "00000000", -- 2377 - 0x949  :    0 - 0x0
    "00000000", -- 2378 - 0x94a  :    0 - 0x0
    "00000000", -- 2379 - 0x94b  :    0 - 0x0
    "00001000", -- 2380 - 0x94c  :    8 - 0x8
    "00111000", -- 2381 - 0x94d  :   56 - 0x38
    "01110000", -- 2382 - 0x94e  :  112 - 0x70
    "11100000", -- 2383 - 0x94f  :  224 - 0xe0
    "00100000", -- 2384 - 0x950  :   32 - 0x20 -- Background 0x95
    "01001111", -- 2385 - 0x951  :   79 - 0x4f
    "11110011", -- 2386 - 0x952  :  243 - 0xf3
    "00001100", -- 2387 - 0x953  :   12 - 0xc
    "00110000", -- 2388 - 0x954  :   48 - 0x30
    "11111111", -- 2389 - 0x955  :  255 - 0xff
    "00000001", -- 2390 - 0x956  :    1 - 0x1
    "11111111", -- 2391 - 0x957  :  255 - 0xff
    "11000000", -- 2392 - 0x958  :  192 - 0xc0 -- plane 1
    "10000000", -- 2393 - 0x959  :  128 - 0x80
    "00001100", -- 2394 - 0x95a  :   12 - 0xc
    "11110000", -- 2395 - 0x95b  :  240 - 0xf0
    "11000000", -- 2396 - 0x95c  :  192 - 0xc0
    "00000000", -- 2397 - 0x95d  :    0 - 0x0
    "11111110", -- 2398 - 0x95e  :  254 - 0xfe
    "00000000", -- 2399 - 0x95f  :    0 - 0x0
    "01111111", -- 2400 - 0x960  :  127 - 0x7f -- Background 0x96
    "11111111", -- 2401 - 0x961  :  255 - 0xff
    "11111111", -- 2402 - 0x962  :  255 - 0xff
    "11111111", -- 2403 - 0x963  :  255 - 0xff
    "11111011", -- 2404 - 0x964  :  251 - 0xfb
    "11111111", -- 2405 - 0x965  :  255 - 0xff
    "11111111", -- 2406 - 0x966  :  255 - 0xff
    "11111111", -- 2407 - 0x967  :  255 - 0xff
    "00000000", -- 2408 - 0x968  :    0 - 0x0 -- plane 1
    "00111111", -- 2409 - 0x969  :   63 - 0x3f
    "01111111", -- 2410 - 0x96a  :  127 - 0x7f
    "01111111", -- 2411 - 0x96b  :  127 - 0x7f
    "01111111", -- 2412 - 0x96c  :  127 - 0x7f
    "01111111", -- 2413 - 0x96d  :  127 - 0x7f
    "01111111", -- 2414 - 0x96e  :  127 - 0x7f
    "01111111", -- 2415 - 0x96f  :  127 - 0x7f
    "11111111", -- 2416 - 0x970  :  255 - 0xff -- Background 0x97
    "11111111", -- 2417 - 0x971  :  255 - 0xff
    "11111111", -- 2418 - 0x972  :  255 - 0xff
    "11111111", -- 2419 - 0x973  :  255 - 0xff
    "11111111", -- 2420 - 0x974  :  255 - 0xff
    "11111111", -- 2421 - 0x975  :  255 - 0xff
    "11111110", -- 2422 - 0x976  :  254 - 0xfe
    "11111111", -- 2423 - 0x977  :  255 - 0xff
    "01111111", -- 2424 - 0x978  :  127 - 0x7f -- plane 1
    "01111111", -- 2425 - 0x979  :  127 - 0x7f
    "00111111", -- 2426 - 0x97a  :   63 - 0x3f
    "01111111", -- 2427 - 0x97b  :  127 - 0x7f
    "01111111", -- 2428 - 0x97c  :  127 - 0x7f
    "01111111", -- 2429 - 0x97d  :  127 - 0x7f
    "01111111", -- 2430 - 0x97e  :  127 - 0x7f
    "01111111", -- 2431 - 0x97f  :  127 - 0x7f
    "11111111", -- 2432 - 0x980  :  255 - 0xff -- Background 0x98
    "10111111", -- 2433 - 0x981  :  191 - 0xbf
    "11111111", -- 2434 - 0x982  :  255 - 0xff
    "11111111", -- 2435 - 0x983  :  255 - 0xff
    "11111011", -- 2436 - 0x984  :  251 - 0xfb
    "11111111", -- 2437 - 0x985  :  255 - 0xff
    "11111111", -- 2438 - 0x986  :  255 - 0xff
    "11111111", -- 2439 - 0x987  :  255 - 0xff
    "00000000", -- 2440 - 0x988  :    0 - 0x0 -- plane 1
    "11011111", -- 2441 - 0x989  :  223 - 0xdf
    "11111111", -- 2442 - 0x98a  :  255 - 0xff
    "11111111", -- 2443 - 0x98b  :  255 - 0xff
    "11111111", -- 2444 - 0x98c  :  255 - 0xff
    "11111111", -- 2445 - 0x98d  :  255 - 0xff
    "11111111", -- 2446 - 0x98e  :  255 - 0xff
    "11111111", -- 2447 - 0x98f  :  255 - 0xff
    "11111111", -- 2448 - 0x990  :  255 - 0xff -- Background 0x99
    "11111111", -- 2449 - 0x991  :  255 - 0xff
    "11111111", -- 2450 - 0x992  :  255 - 0xff
    "11111111", -- 2451 - 0x993  :  255 - 0xff
    "11111111", -- 2452 - 0x994  :  255 - 0xff
    "11111111", -- 2453 - 0x995  :  255 - 0xff
    "11111110", -- 2454 - 0x996  :  254 - 0xfe
    "11111111", -- 2455 - 0x997  :  255 - 0xff
    "11111111", -- 2456 - 0x998  :  255 - 0xff -- plane 1
    "11111111", -- 2457 - 0x999  :  255 - 0xff
    "10111111", -- 2458 - 0x99a  :  191 - 0xbf
    "11111111", -- 2459 - 0x99b  :  255 - 0xff
    "11111111", -- 2460 - 0x99c  :  255 - 0xff
    "11111111", -- 2461 - 0x99d  :  255 - 0xff
    "11111111", -- 2462 - 0x99e  :  255 - 0xff
    "11111111", -- 2463 - 0x99f  :  255 - 0xff
    "11111110", -- 2464 - 0x9a0  :  254 - 0xfe -- Background 0x9a
    "11111111", -- 2465 - 0x9a1  :  255 - 0xff
    "11111111", -- 2466 - 0x9a2  :  255 - 0xff
    "11111111", -- 2467 - 0x9a3  :  255 - 0xff
    "11111011", -- 2468 - 0x9a4  :  251 - 0xfb
    "11111111", -- 2469 - 0x9a5  :  255 - 0xff
    "11111111", -- 2470 - 0x9a6  :  255 - 0xff
    "11111111", -- 2471 - 0x9a7  :  255 - 0xff
    "00000000", -- 2472 - 0x9a8  :    0 - 0x0 -- plane 1
    "10111100", -- 2473 - 0x9a9  :  188 - 0xbc
    "11111110", -- 2474 - 0x9aa  :  254 - 0xfe
    "11111110", -- 2475 - 0x9ab  :  254 - 0xfe
    "11111110", -- 2476 - 0x9ac  :  254 - 0xfe
    "11111110", -- 2477 - 0x9ad  :  254 - 0xfe
    "11111110", -- 2478 - 0x9ae  :  254 - 0xfe
    "11111110", -- 2479 - 0x9af  :  254 - 0xfe
    "11111111", -- 2480 - 0x9b0  :  255 - 0xff -- Background 0x9b
    "11111111", -- 2481 - 0x9b1  :  255 - 0xff
    "11111111", -- 2482 - 0x9b2  :  255 - 0xff
    "11111111", -- 2483 - 0x9b3  :  255 - 0xff
    "11111111", -- 2484 - 0x9b4  :  255 - 0xff
    "11111111", -- 2485 - 0x9b5  :  255 - 0xff
    "11111111", -- 2486 - 0x9b6  :  255 - 0xff
    "11111111", -- 2487 - 0x9b7  :  255 - 0xff
    "11111110", -- 2488 - 0x9b8  :  254 - 0xfe -- plane 1
    "11111110", -- 2489 - 0x9b9  :  254 - 0xfe
    "10111110", -- 2490 - 0x9ba  :  190 - 0xbe
    "11111110", -- 2491 - 0x9bb  :  254 - 0xfe
    "11111110", -- 2492 - 0x9bc  :  254 - 0xfe
    "11111110", -- 2493 - 0x9bd  :  254 - 0xfe
    "11111110", -- 2494 - 0x9be  :  254 - 0xfe
    "11111110", -- 2495 - 0x9bf  :  254 - 0xfe
    "11111111", -- 2496 - 0x9c0  :  255 - 0xff -- Background 0x9c
    "11111111", -- 2497 - 0x9c1  :  255 - 0xff
    "10100000", -- 2498 - 0x9c2  :  160 - 0xa0
    "10010000", -- 2499 - 0x9c3  :  144 - 0x90
    "10001000", -- 2500 - 0x9c4  :  136 - 0x88
    "10000100", -- 2501 - 0x9c5  :  132 - 0x84
    "01101010", -- 2502 - 0x9c6  :  106 - 0x6a
    "00111111", -- 2503 - 0x9c7  :   63 - 0x3f
    "00000000", -- 2504 - 0x9c8  :    0 - 0x0 -- plane 1
    "00111111", -- 2505 - 0x9c9  :   63 - 0x3f
    "01011111", -- 2506 - 0x9ca  :   95 - 0x5f
    "01101111", -- 2507 - 0x9cb  :  111 - 0x6f
    "01110111", -- 2508 - 0x9cc  :  119 - 0x77
    "01111011", -- 2509 - 0x9cd  :  123 - 0x7b
    "00010101", -- 2510 - 0x9ce  :   21 - 0x15
    "00000000", -- 2511 - 0x9cf  :    0 - 0x0
    "11111111", -- 2512 - 0x9d0  :  255 - 0xff -- Background 0x9d
    "11111111", -- 2513 - 0x9d1  :  255 - 0xff
    "00100001", -- 2514 - 0x9d2  :   33 - 0x21
    "00010001", -- 2515 - 0x9d3  :   17 - 0x11
    "00001001", -- 2516 - 0x9d4  :    9 - 0x9
    "00000101", -- 2517 - 0x9d5  :    5 - 0x5
    "10101010", -- 2518 - 0x9d6  :  170 - 0xaa
    "11111100", -- 2519 - 0x9d7  :  252 - 0xfc
    "00000000", -- 2520 - 0x9d8  :    0 - 0x0 -- plane 1
    "10111110", -- 2521 - 0x9d9  :  190 - 0xbe
    "11011110", -- 2522 - 0x9da  :  222 - 0xde
    "11101110", -- 2523 - 0x9db  :  238 - 0xee
    "11110110", -- 2524 - 0x9dc  :  246 - 0xf6
    "11111010", -- 2525 - 0x9dd  :  250 - 0xfa
    "01010100", -- 2526 - 0x9de  :   84 - 0x54
    "00000000", -- 2527 - 0x9df  :    0 - 0x0
    "11111111", -- 2528 - 0x9e0  :  255 - 0xff -- Background 0x9e
    "11111111", -- 2529 - 0x9e1  :  255 - 0xff
    "00100000", -- 2530 - 0x9e2  :   32 - 0x20
    "00010000", -- 2531 - 0x9e3  :   16 - 0x10
    "00001000", -- 2532 - 0x9e4  :    8 - 0x8
    "00000100", -- 2533 - 0x9e5  :    4 - 0x4
    "10101010", -- 2534 - 0x9e6  :  170 - 0xaa
    "11111111", -- 2535 - 0x9e7  :  255 - 0xff
    "00000000", -- 2536 - 0x9e8  :    0 - 0x0 -- plane 1
    "10111111", -- 2537 - 0x9e9  :  191 - 0xbf
    "11011111", -- 2538 - 0x9ea  :  223 - 0xdf
    "11101111", -- 2539 - 0x9eb  :  239 - 0xef
    "11110111", -- 2540 - 0x9ec  :  247 - 0xf7
    "11111011", -- 2541 - 0x9ed  :  251 - 0xfb
    "01010101", -- 2542 - 0x9ee  :   85 - 0x55
    "00000000", -- 2543 - 0x9ef  :    0 - 0x0
    "00000000", -- 2544 - 0x9f0  :    0 - 0x0 -- Background 0x9f
    "00000000", -- 2545 - 0x9f1  :    0 - 0x0
    "00000000", -- 2546 - 0x9f2  :    0 - 0x0
    "00000000", -- 2547 - 0x9f3  :    0 - 0x0
    "00000000", -- 2548 - 0x9f4  :    0 - 0x0
    "00000000", -- 2549 - 0x9f5  :    0 - 0x0
    "00000000", -- 2550 - 0x9f6  :    0 - 0x0
    "00000000", -- 2551 - 0x9f7  :    0 - 0x0
    "00000000", -- 2552 - 0x9f8  :    0 - 0x0 -- plane 1
    "00000000", -- 2553 - 0x9f9  :    0 - 0x0
    "00000000", -- 2554 - 0x9fa  :    0 - 0x0
    "00000000", -- 2555 - 0x9fb  :    0 - 0x0
    "00000000", -- 2556 - 0x9fc  :    0 - 0x0
    "00000000", -- 2557 - 0x9fd  :    0 - 0x0
    "00000000", -- 2558 - 0x9fe  :    0 - 0x0
    "00000000", -- 2559 - 0x9ff  :    0 - 0x0
    "11111111", -- 2560 - 0xa00  :  255 - 0xff -- Background 0xa0
    "11010101", -- 2561 - 0xa01  :  213 - 0xd5
    "11111111", -- 2562 - 0xa02  :  255 - 0xff
    "00000010", -- 2563 - 0xa03  :    2 - 0x2
    "00000010", -- 2564 - 0xa04  :    2 - 0x2
    "00000010", -- 2565 - 0xa05  :    2 - 0x2
    "00000010", -- 2566 - 0xa06  :    2 - 0x2
    "00000010", -- 2567 - 0xa07  :    2 - 0x2
    "00000000", -- 2568 - 0xa08  :    0 - 0x0 -- plane 1
    "01111111", -- 2569 - 0xa09  :  127 - 0x7f
    "00000000", -- 2570 - 0xa0a  :    0 - 0x0
    "00000001", -- 2571 - 0xa0b  :    1 - 0x1
    "00000001", -- 2572 - 0xa0c  :    1 - 0x1
    "00000001", -- 2573 - 0xa0d  :    1 - 0x1
    "00000001", -- 2574 - 0xa0e  :    1 - 0x1
    "00000001", -- 2575 - 0xa0f  :    1 - 0x1
    "00000010", -- 2576 - 0xa10  :    2 - 0x2 -- Background 0xa1
    "00000010", -- 2577 - 0xa11  :    2 - 0x2
    "00000010", -- 2578 - 0xa12  :    2 - 0x2
    "00000010", -- 2579 - 0xa13  :    2 - 0x2
    "00000010", -- 2580 - 0xa14  :    2 - 0x2
    "00000010", -- 2581 - 0xa15  :    2 - 0x2
    "00000010", -- 2582 - 0xa16  :    2 - 0x2
    "00000010", -- 2583 - 0xa17  :    2 - 0x2
    "00000001", -- 2584 - 0xa18  :    1 - 0x1 -- plane 1
    "00000001", -- 2585 - 0xa19  :    1 - 0x1
    "00000001", -- 2586 - 0xa1a  :    1 - 0x1
    "00000001", -- 2587 - 0xa1b  :    1 - 0x1
    "00000001", -- 2588 - 0xa1c  :    1 - 0x1
    "00000001", -- 2589 - 0xa1d  :    1 - 0x1
    "00000001", -- 2590 - 0xa1e  :    1 - 0x1
    "00000001", -- 2591 - 0xa1f  :    1 - 0x1
    "11111111", -- 2592 - 0xa20  :  255 - 0xff -- Background 0xa2
    "01010101", -- 2593 - 0xa21  :   85 - 0x55
    "11111111", -- 2594 - 0xa22  :  255 - 0xff
    "01000000", -- 2595 - 0xa23  :   64 - 0x40
    "01000000", -- 2596 - 0xa24  :   64 - 0x40
    "01000000", -- 2597 - 0xa25  :   64 - 0x40
    "01000000", -- 2598 - 0xa26  :   64 - 0x40
    "01000000", -- 2599 - 0xa27  :   64 - 0x40
    "00000000", -- 2600 - 0xa28  :    0 - 0x0 -- plane 1
    "11111110", -- 2601 - 0xa29  :  254 - 0xfe
    "00000000", -- 2602 - 0xa2a  :    0 - 0x0
    "10000000", -- 2603 - 0xa2b  :  128 - 0x80
    "10000000", -- 2604 - 0xa2c  :  128 - 0x80
    "10000000", -- 2605 - 0xa2d  :  128 - 0x80
    "10000000", -- 2606 - 0xa2e  :  128 - 0x80
    "10000000", -- 2607 - 0xa2f  :  128 - 0x80
    "01000000", -- 2608 - 0xa30  :   64 - 0x40 -- Background 0xa3
    "01000000", -- 2609 - 0xa31  :   64 - 0x40
    "01000000", -- 2610 - 0xa32  :   64 - 0x40
    "01000000", -- 2611 - 0xa33  :   64 - 0x40
    "01000000", -- 2612 - 0xa34  :   64 - 0x40
    "01000000", -- 2613 - 0xa35  :   64 - 0x40
    "01000000", -- 2614 - 0xa36  :   64 - 0x40
    "01000000", -- 2615 - 0xa37  :   64 - 0x40
    "10000000", -- 2616 - 0xa38  :  128 - 0x80 -- plane 1
    "10000000", -- 2617 - 0xa39  :  128 - 0x80
    "10000000", -- 2618 - 0xa3a  :  128 - 0x80
    "10000000", -- 2619 - 0xa3b  :  128 - 0x80
    "10000000", -- 2620 - 0xa3c  :  128 - 0x80
    "10000000", -- 2621 - 0xa3d  :  128 - 0x80
    "10000000", -- 2622 - 0xa3e  :  128 - 0x80
    "10000000", -- 2623 - 0xa3f  :  128 - 0x80
    "00110001", -- 2624 - 0xa40  :   49 - 0x31 -- Background 0xa4
    "01001000", -- 2625 - 0xa41  :   72 - 0x48
    "01000101", -- 2626 - 0xa42  :   69 - 0x45
    "10000101", -- 2627 - 0xa43  :  133 - 0x85
    "10000011", -- 2628 - 0xa44  :  131 - 0x83
    "10000010", -- 2629 - 0xa45  :  130 - 0x82
    "01100010", -- 2630 - 0xa46  :   98 - 0x62
    "00010010", -- 2631 - 0xa47  :   18 - 0x12
    "00000000", -- 2632 - 0xa48  :    0 - 0x0 -- plane 1
    "00110000", -- 2633 - 0xa49  :   48 - 0x30
    "00111000", -- 2634 - 0xa4a  :   56 - 0x38
    "01111000", -- 2635 - 0xa4b  :  120 - 0x78
    "01111100", -- 2636 - 0xa4c  :  124 - 0x7c
    "01111101", -- 2637 - 0xa4d  :  125 - 0x7d
    "00011101", -- 2638 - 0xa4e  :   29 - 0x1d
    "00001101", -- 2639 - 0xa4f  :   13 - 0xd
    "00110010", -- 2640 - 0xa50  :   50 - 0x32 -- Background 0xa5
    "00100010", -- 2641 - 0xa51  :   34 - 0x22
    "01000010", -- 2642 - 0xa52  :   66 - 0x42
    "01000000", -- 2643 - 0xa53  :   64 - 0x40
    "01000000", -- 2644 - 0xa54  :   64 - 0x40
    "00100000", -- 2645 - 0xa55  :   32 - 0x20
    "00011110", -- 2646 - 0xa56  :   30 - 0x1e
    "00000111", -- 2647 - 0xa57  :    7 - 0x7
    "00001101", -- 2648 - 0xa58  :   13 - 0xd -- plane 1
    "00011101", -- 2649 - 0xa59  :   29 - 0x1d
    "00111101", -- 2650 - 0xa5a  :   61 - 0x3d
    "00111111", -- 2651 - 0xa5b  :   63 - 0x3f
    "00111111", -- 2652 - 0xa5c  :   63 - 0x3f
    "00011111", -- 2653 - 0xa5d  :   31 - 0x1f
    "00000001", -- 2654 - 0xa5e  :    1 - 0x1
    "00000000", -- 2655 - 0xa5f  :    0 - 0x0
    "10000000", -- 2656 - 0xa60  :  128 - 0x80 -- Background 0xa6
    "11100000", -- 2657 - 0xa61  :  224 - 0xe0
    "00111000", -- 2658 - 0xa62  :   56 - 0x38
    "00100100", -- 2659 - 0xa63  :   36 - 0x24
    "00000100", -- 2660 - 0xa64  :    4 - 0x4
    "00001000", -- 2661 - 0xa65  :    8 - 0x8
    "00110000", -- 2662 - 0xa66  :   48 - 0x30
    "00100000", -- 2663 - 0xa67  :   32 - 0x20
    "00000000", -- 2664 - 0xa68  :    0 - 0x0 -- plane 1
    "00000000", -- 2665 - 0xa69  :    0 - 0x0
    "11100000", -- 2666 - 0xa6a  :  224 - 0xe0
    "11111000", -- 2667 - 0xa6b  :  248 - 0xf8
    "11111000", -- 2668 - 0xa6c  :  248 - 0xf8
    "11110000", -- 2669 - 0xa6d  :  240 - 0xf0
    "11000000", -- 2670 - 0xa6e  :  192 - 0xc0
    "11000000", -- 2671 - 0xa6f  :  192 - 0xc0
    "00110000", -- 2672 - 0xa70  :   48 - 0x30 -- Background 0xa7
    "00001000", -- 2673 - 0xa71  :    8 - 0x8
    "00001000", -- 2674 - 0xa72  :    8 - 0x8
    "00110000", -- 2675 - 0xa73  :   48 - 0x30
    "00100000", -- 2676 - 0xa74  :   32 - 0x20
    "00100000", -- 2677 - 0xa75  :   32 - 0x20
    "00110000", -- 2678 - 0xa76  :   48 - 0x30
    "11110000", -- 2679 - 0xa77  :  240 - 0xf0
    "11000000", -- 2680 - 0xa78  :  192 - 0xc0 -- plane 1
    "11110000", -- 2681 - 0xa79  :  240 - 0xf0
    "11110000", -- 2682 - 0xa7a  :  240 - 0xf0
    "11000000", -- 2683 - 0xa7b  :  192 - 0xc0
    "11000000", -- 2684 - 0xa7c  :  192 - 0xc0
    "11000000", -- 2685 - 0xa7d  :  192 - 0xc0
    "11000000", -- 2686 - 0xa7e  :  192 - 0xc0
    "00000000", -- 2687 - 0xa7f  :    0 - 0x0
    "11111111", -- 2688 - 0xa80  :  255 - 0xff -- Background 0xa8
    "11010010", -- 2689 - 0xa81  :  210 - 0xd2
    "11110100", -- 2690 - 0xa82  :  244 - 0xf4
    "11011000", -- 2691 - 0xa83  :  216 - 0xd8
    "11111000", -- 2692 - 0xa84  :  248 - 0xf8
    "11010100", -- 2693 - 0xa85  :  212 - 0xd4
    "11110010", -- 2694 - 0xa86  :  242 - 0xf2
    "11010001", -- 2695 - 0xa87  :  209 - 0xd1
    "00000000", -- 2696 - 0xa88  :    0 - 0x0 -- plane 1
    "01100000", -- 2697 - 0xa89  :   96 - 0x60
    "01100000", -- 2698 - 0xa8a  :   96 - 0x60
    "01100000", -- 2699 - 0xa8b  :   96 - 0x60
    "01100000", -- 2700 - 0xa8c  :   96 - 0x60
    "01100000", -- 2701 - 0xa8d  :   96 - 0x60
    "01100000", -- 2702 - 0xa8e  :   96 - 0x60
    "01100000", -- 2703 - 0xa8f  :   96 - 0x60
    "11110001", -- 2704 - 0xa90  :  241 - 0xf1 -- Background 0xa9
    "11010010", -- 2705 - 0xa91  :  210 - 0xd2
    "11110100", -- 2706 - 0xa92  :  244 - 0xf4
    "11011000", -- 2707 - 0xa93  :  216 - 0xd8
    "11111000", -- 2708 - 0xa94  :  248 - 0xf8
    "11010100", -- 2709 - 0xa95  :  212 - 0xd4
    "11110010", -- 2710 - 0xa96  :  242 - 0xf2
    "11111111", -- 2711 - 0xa97  :  255 - 0xff
    "01100000", -- 2712 - 0xa98  :   96 - 0x60 -- plane 1
    "01100000", -- 2713 - 0xa99  :   96 - 0x60
    "01100000", -- 2714 - 0xa9a  :   96 - 0x60
    "01100000", -- 2715 - 0xa9b  :   96 - 0x60
    "01100000", -- 2716 - 0xa9c  :   96 - 0x60
    "01100000", -- 2717 - 0xa9d  :   96 - 0x60
    "01100000", -- 2718 - 0xa9e  :   96 - 0x60
    "00000000", -- 2719 - 0xa9f  :    0 - 0x0
    "11111111", -- 2720 - 0xaa0  :  255 - 0xff -- Background 0xaa
    "01000010", -- 2721 - 0xaa1  :   66 - 0x42
    "00100100", -- 2722 - 0xaa2  :   36 - 0x24
    "00011000", -- 2723 - 0xaa3  :   24 - 0x18
    "00011000", -- 2724 - 0xaa4  :   24 - 0x18
    "00100100", -- 2725 - 0xaa5  :   36 - 0x24
    "01000010", -- 2726 - 0xaa6  :   66 - 0x42
    "10000001", -- 2727 - 0xaa7  :  129 - 0x81
    "00000000", -- 2728 - 0xaa8  :    0 - 0x0 -- plane 1
    "00000000", -- 2729 - 0xaa9  :    0 - 0x0
    "00000000", -- 2730 - 0xaaa  :    0 - 0x0
    "00000000", -- 2731 - 0xaab  :    0 - 0x0
    "00000000", -- 2732 - 0xaac  :    0 - 0x0
    "00000000", -- 2733 - 0xaad  :    0 - 0x0
    "00000000", -- 2734 - 0xaae  :    0 - 0x0
    "00000000", -- 2735 - 0xaaf  :    0 - 0x0
    "10000001", -- 2736 - 0xab0  :  129 - 0x81 -- Background 0xab
    "01000010", -- 2737 - 0xab1  :   66 - 0x42
    "00100100", -- 2738 - 0xab2  :   36 - 0x24
    "00011000", -- 2739 - 0xab3  :   24 - 0x18
    "00011000", -- 2740 - 0xab4  :   24 - 0x18
    "00100100", -- 2741 - 0xab5  :   36 - 0x24
    "01000010", -- 2742 - 0xab6  :   66 - 0x42
    "11111111", -- 2743 - 0xab7  :  255 - 0xff
    "00000000", -- 2744 - 0xab8  :    0 - 0x0 -- plane 1
    "00000000", -- 2745 - 0xab9  :    0 - 0x0
    "00000000", -- 2746 - 0xaba  :    0 - 0x0
    "00000000", -- 2747 - 0xabb  :    0 - 0x0
    "00000000", -- 2748 - 0xabc  :    0 - 0x0
    "00000000", -- 2749 - 0xabd  :    0 - 0x0
    "00000000", -- 2750 - 0xabe  :    0 - 0x0
    "00000000", -- 2751 - 0xabf  :    0 - 0x0
    "11111111", -- 2752 - 0xac0  :  255 - 0xff -- Background 0xac
    "01001101", -- 2753 - 0xac1  :   77 - 0x4d
    "00101111", -- 2754 - 0xac2  :   47 - 0x2f
    "00011101", -- 2755 - 0xac3  :   29 - 0x1d
    "00011111", -- 2756 - 0xac4  :   31 - 0x1f
    "00101101", -- 2757 - 0xac5  :   45 - 0x2d
    "01001111", -- 2758 - 0xac6  :   79 - 0x4f
    "10001101", -- 2759 - 0xac7  :  141 - 0x8d
    "00000000", -- 2760 - 0xac8  :    0 - 0x0 -- plane 1
    "00000110", -- 2761 - 0xac9  :    6 - 0x6
    "00000110", -- 2762 - 0xaca  :    6 - 0x6
    "00000110", -- 2763 - 0xacb  :    6 - 0x6
    "00000110", -- 2764 - 0xacc  :    6 - 0x6
    "00000110", -- 2765 - 0xacd  :    6 - 0x6
    "00000110", -- 2766 - 0xace  :    6 - 0x6
    "00000110", -- 2767 - 0xacf  :    6 - 0x6
    "10001111", -- 2768 - 0xad0  :  143 - 0x8f -- Background 0xad
    "01001101", -- 2769 - 0xad1  :   77 - 0x4d
    "00101111", -- 2770 - 0xad2  :   47 - 0x2f
    "00011101", -- 2771 - 0xad3  :   29 - 0x1d
    "00011111", -- 2772 - 0xad4  :   31 - 0x1f
    "00101101", -- 2773 - 0xad5  :   45 - 0x2d
    "01001111", -- 2774 - 0xad6  :   79 - 0x4f
    "11111111", -- 2775 - 0xad7  :  255 - 0xff
    "00000110", -- 2776 - 0xad8  :    6 - 0x6 -- plane 1
    "00000110", -- 2777 - 0xad9  :    6 - 0x6
    "00000110", -- 2778 - 0xada  :    6 - 0x6
    "00000110", -- 2779 - 0xadb  :    6 - 0x6
    "00000110", -- 2780 - 0xadc  :    6 - 0x6
    "00000110", -- 2781 - 0xadd  :    6 - 0x6
    "00000110", -- 2782 - 0xade  :    6 - 0x6
    "00000000", -- 2783 - 0xadf  :    0 - 0x0
    "00000001", -- 2784 - 0xae0  :    1 - 0x1 -- Background 0xae
    "00000011", -- 2785 - 0xae1  :    3 - 0x3
    "00000110", -- 2786 - 0xae2  :    6 - 0x6
    "00000111", -- 2787 - 0xae3  :    7 - 0x7
    "00000111", -- 2788 - 0xae4  :    7 - 0x7
    "00000111", -- 2789 - 0xae5  :    7 - 0x7
    "00000110", -- 2790 - 0xae6  :    6 - 0x6
    "00000111", -- 2791 - 0xae7  :    7 - 0x7
    "00000000", -- 2792 - 0xae8  :    0 - 0x0 -- plane 1
    "00000001", -- 2793 - 0xae9  :    1 - 0x1
    "00000011", -- 2794 - 0xaea  :    3 - 0x3
    "00000010", -- 2795 - 0xaeb  :    2 - 0x2
    "00000010", -- 2796 - 0xaec  :    2 - 0x2
    "00000000", -- 2797 - 0xaed  :    0 - 0x0
    "00000011", -- 2798 - 0xaee  :    3 - 0x3
    "00000010", -- 2799 - 0xaef  :    2 - 0x2
    "00000110", -- 2800 - 0xaf0  :    6 - 0x6 -- Background 0xaf
    "00000110", -- 2801 - 0xaf1  :    6 - 0x6
    "00001110", -- 2802 - 0xaf2  :   14 - 0xe
    "00001111", -- 2803 - 0xaf3  :   15 - 0xf
    "00001110", -- 2804 - 0xaf4  :   14 - 0xe
    "00011010", -- 2805 - 0xaf5  :   26 - 0x1a
    "00011011", -- 2806 - 0xaf6  :   27 - 0x1b
    "00001111", -- 2807 - 0xaf7  :   15 - 0xf
    "00000001", -- 2808 - 0xaf8  :    1 - 0x1 -- plane 1
    "00000011", -- 2809 - 0xaf9  :    3 - 0x3
    "00000101", -- 2810 - 0xafa  :    5 - 0x5
    "00000100", -- 2811 - 0xafb  :    4 - 0x4
    "00000101", -- 2812 - 0xafc  :    5 - 0x5
    "00001101", -- 2813 - 0xafd  :   13 - 0xd
    "00001100", -- 2814 - 0xafe  :   12 - 0xc
    "00000001", -- 2815 - 0xaff  :    1 - 0x1
    "00000000", -- 2816 - 0xb00  :    0 - 0x0 -- Background 0xb0
    "11000000", -- 2817 - 0xb01  :  192 - 0xc0
    "11110000", -- 2818 - 0xb02  :  240 - 0xf0
    "10001000", -- 2819 - 0xb03  :  136 - 0x88
    "00010100", -- 2820 - 0xb04  :   20 - 0x14
    "01101000", -- 2821 - 0xb05  :  104 - 0x68
    "10101000", -- 2822 - 0xb06  :  168 - 0xa8
    "00101100", -- 2823 - 0xb07  :   44 - 0x2c
    "00000000", -- 2824 - 0xb08  :    0 - 0x0 -- plane 1
    "00000000", -- 2825 - 0xb09  :    0 - 0x0
    "01000000", -- 2826 - 0xb0a  :   64 - 0x40
    "11110000", -- 2827 - 0xb0b  :  240 - 0xf0
    "11101000", -- 2828 - 0xb0c  :  232 - 0xe8
    "10010000", -- 2829 - 0xb0d  :  144 - 0x90
    "01010000", -- 2830 - 0xb0e  :   80 - 0x50
    "11010000", -- 2831 - 0xb0f  :  208 - 0xd0
    "00000100", -- 2832 - 0xb10  :    4 - 0x4 -- Background 0xb1
    "00111000", -- 2833 - 0xb11  :   56 - 0x38
    "00010000", -- 2834 - 0xb12  :   16 - 0x10
    "10100000", -- 2835 - 0xb13  :  160 - 0xa0
    "01100000", -- 2836 - 0xb14  :   96 - 0x60
    "00100000", -- 2837 - 0xb15  :   32 - 0x20
    "00010000", -- 2838 - 0xb16  :   16 - 0x10
    "10001000", -- 2839 - 0xb17  :  136 - 0x88
    "11111000", -- 2840 - 0xb18  :  248 - 0xf8 -- plane 1
    "11000000", -- 2841 - 0xb19  :  192 - 0xc0
    "11100000", -- 2842 - 0xb1a  :  224 - 0xe0
    "01000000", -- 2843 - 0xb1b  :   64 - 0x40
    "10000000", -- 2844 - 0xb1c  :  128 - 0x80
    "11000000", -- 2845 - 0xb1d  :  192 - 0xc0
    "11100000", -- 2846 - 0xb1e  :  224 - 0xe0
    "01110000", -- 2847 - 0xb1f  :  112 - 0x70
    "00001111", -- 2848 - 0xb20  :   15 - 0xf -- Background 0xb2
    "00011011", -- 2849 - 0xb21  :   27 - 0x1b
    "00011011", -- 2850 - 0xb22  :   27 - 0x1b
    "00001110", -- 2851 - 0xb23  :   14 - 0xe
    "00000110", -- 2852 - 0xb24  :    6 - 0x6
    "00001100", -- 2853 - 0xb25  :   12 - 0xc
    "00001100", -- 2854 - 0xb26  :   12 - 0xc
    "00111111", -- 2855 - 0xb27  :   63 - 0x3f
    "00000001", -- 2856 - 0xb28  :    1 - 0x1 -- plane 1
    "00001101", -- 2857 - 0xb29  :   13 - 0xd
    "00001101", -- 2858 - 0xb2a  :   13 - 0xd
    "00000011", -- 2859 - 0xb2b  :    3 - 0x3
    "00000011", -- 2860 - 0xb2c  :    3 - 0x3
    "00000111", -- 2861 - 0xb2d  :    7 - 0x7
    "00000111", -- 2862 - 0xb2e  :    7 - 0x7
    "00000000", -- 2863 - 0xb2f  :    0 - 0x0
    "01111111", -- 2864 - 0xb30  :  127 - 0x7f -- Background 0xb3
    "01100000", -- 2865 - 0xb31  :   96 - 0x60
    "01100000", -- 2866 - 0xb32  :   96 - 0x60
    "01100000", -- 2867 - 0xb33  :   96 - 0x60
    "01100000", -- 2868 - 0xb34  :   96 - 0x60
    "01100000", -- 2869 - 0xb35  :   96 - 0x60
    "01101010", -- 2870 - 0xb36  :  106 - 0x6a
    "01111111", -- 2871 - 0xb37  :  127 - 0x7f
    "00111111", -- 2872 - 0xb38  :   63 - 0x3f -- plane 1
    "00111111", -- 2873 - 0xb39  :   63 - 0x3f
    "00111111", -- 2874 - 0xb3a  :   63 - 0x3f
    "00111111", -- 2875 - 0xb3b  :   63 - 0x3f
    "00111111", -- 2876 - 0xb3c  :   63 - 0x3f
    "00111111", -- 2877 - 0xb3d  :   63 - 0x3f
    "00110101", -- 2878 - 0xb3e  :   53 - 0x35
    "00000000", -- 2879 - 0xb3f  :    0 - 0x0
    "01001000", -- 2880 - 0xb40  :   72 - 0x48 -- Background 0xb4
    "00110000", -- 2881 - 0xb41  :   48 - 0x30
    "00010000", -- 2882 - 0xb42  :   16 - 0x10
    "00010000", -- 2883 - 0xb43  :   16 - 0x10
    "00001000", -- 2884 - 0xb44  :    8 - 0x8
    "00001000", -- 2885 - 0xb45  :    8 - 0x8
    "00001000", -- 2886 - 0xb46  :    8 - 0x8
    "11111100", -- 2887 - 0xb47  :  252 - 0xfc
    "10110000", -- 2888 - 0xb48  :  176 - 0xb0 -- plane 1
    "11000000", -- 2889 - 0xb49  :  192 - 0xc0
    "11100000", -- 2890 - 0xb4a  :  224 - 0xe0
    "11100000", -- 2891 - 0xb4b  :  224 - 0xe0
    "11110000", -- 2892 - 0xb4c  :  240 - 0xf0
    "11110000", -- 2893 - 0xb4d  :  240 - 0xf0
    "11110000", -- 2894 - 0xb4e  :  240 - 0xf0
    "00000000", -- 2895 - 0xb4f  :    0 - 0x0
    "11111110", -- 2896 - 0xb50  :  254 - 0xfe -- Background 0xb5
    "00000110", -- 2897 - 0xb51  :    6 - 0x6
    "00000010", -- 2898 - 0xb52  :    2 - 0x2
    "00000110", -- 2899 - 0xb53  :    6 - 0x6
    "00000010", -- 2900 - 0xb54  :    2 - 0x2
    "00000110", -- 2901 - 0xb55  :    6 - 0x6
    "10101010", -- 2902 - 0xb56  :  170 - 0xaa
    "11111110", -- 2903 - 0xb57  :  254 - 0xfe
    "11111100", -- 2904 - 0xb58  :  252 - 0xfc -- plane 1
    "11111000", -- 2905 - 0xb59  :  248 - 0xf8
    "11111100", -- 2906 - 0xb5a  :  252 - 0xfc
    "11111000", -- 2907 - 0xb5b  :  248 - 0xf8
    "11111100", -- 2908 - 0xb5c  :  252 - 0xfc
    "11111000", -- 2909 - 0xb5d  :  248 - 0xf8
    "01010100", -- 2910 - 0xb5e  :   84 - 0x54
    "00000000", -- 2911 - 0xb5f  :    0 - 0x0
    "11111111", -- 2912 - 0xb60  :  255 - 0xff -- Background 0xb6
    "10000000", -- 2913 - 0xb61  :  128 - 0x80
    "10000000", -- 2914 - 0xb62  :  128 - 0x80
    "10000000", -- 2915 - 0xb63  :  128 - 0x80
    "10000000", -- 2916 - 0xb64  :  128 - 0x80
    "10000000", -- 2917 - 0xb65  :  128 - 0x80
    "10010101", -- 2918 - 0xb66  :  149 - 0x95
    "11111111", -- 2919 - 0xb67  :  255 - 0xff
    "00000000", -- 2920 - 0xb68  :    0 - 0x0 -- plane 1
    "01111111", -- 2921 - 0xb69  :  127 - 0x7f
    "01111111", -- 2922 - 0xb6a  :  127 - 0x7f
    "01111111", -- 2923 - 0xb6b  :  127 - 0x7f
    "01111111", -- 2924 - 0xb6c  :  127 - 0x7f
    "01111111", -- 2925 - 0xb6d  :  127 - 0x7f
    "01101010", -- 2926 - 0xb6e  :  106 - 0x6a
    "00000000", -- 2927 - 0xb6f  :    0 - 0x0
    "11111111", -- 2928 - 0xb70  :  255 - 0xff -- Background 0xb7
    "10000100", -- 2929 - 0xb71  :  132 - 0x84
    "10001100", -- 2930 - 0xb72  :  140 - 0x8c
    "10000100", -- 2931 - 0xb73  :  132 - 0x84
    "10001100", -- 2932 - 0xb74  :  140 - 0x8c
    "10000100", -- 2933 - 0xb75  :  132 - 0x84
    "10101100", -- 2934 - 0xb76  :  172 - 0xac
    "11111111", -- 2935 - 0xb77  :  255 - 0xff
    "00000000", -- 2936 - 0xb78  :    0 - 0x0 -- plane 1
    "01111011", -- 2937 - 0xb79  :  123 - 0x7b
    "01110011", -- 2938 - 0xb7a  :  115 - 0x73
    "01111011", -- 2939 - 0xb7b  :  123 - 0x7b
    "01110011", -- 2940 - 0xb7c  :  115 - 0x73
    "01111011", -- 2941 - 0xb7d  :  123 - 0x7b
    "01010011", -- 2942 - 0xb7e  :   83 - 0x53
    "00000000", -- 2943 - 0xb7f  :    0 - 0x0
    "11111111", -- 2944 - 0xb80  :  255 - 0xff -- Background 0xb8
    "00100001", -- 2945 - 0xb81  :   33 - 0x21
    "01100001", -- 2946 - 0xb82  :   97 - 0x61
    "00100011", -- 2947 - 0xb83  :   35 - 0x23
    "01100001", -- 2948 - 0xb84  :   97 - 0x61
    "00100011", -- 2949 - 0xb85  :   35 - 0x23
    "01100101", -- 2950 - 0xb86  :  101 - 0x65
    "11111111", -- 2951 - 0xb87  :  255 - 0xff
    "00000000", -- 2952 - 0xb88  :    0 - 0x0 -- plane 1
    "11011110", -- 2953 - 0xb89  :  222 - 0xde
    "10011110", -- 2954 - 0xb8a  :  158 - 0x9e
    "11011100", -- 2955 - 0xb8b  :  220 - 0xdc
    "10011110", -- 2956 - 0xb8c  :  158 - 0x9e
    "11011100", -- 2957 - 0xb8d  :  220 - 0xdc
    "10011010", -- 2958 - 0xb8e  :  154 - 0x9a
    "00000000", -- 2959 - 0xb8f  :    0 - 0x0
    "11111111", -- 2960 - 0xb90  :  255 - 0xff -- Background 0xb9
    "00000001", -- 2961 - 0xb91  :    1 - 0x1
    "00000011", -- 2962 - 0xb92  :    3 - 0x3
    "00000001", -- 2963 - 0xb93  :    1 - 0x1
    "00000011", -- 2964 - 0xb94  :    3 - 0x3
    "00000001", -- 2965 - 0xb95  :    1 - 0x1
    "10101011", -- 2966 - 0xb96  :  171 - 0xab
    "11111111", -- 2967 - 0xb97  :  255 - 0xff
    "00000000", -- 2968 - 0xb98  :    0 - 0x0 -- plane 1
    "11111110", -- 2969 - 0xb99  :  254 - 0xfe
    "11111100", -- 2970 - 0xb9a  :  252 - 0xfc
    "11111110", -- 2971 - 0xb9b  :  254 - 0xfe
    "11111100", -- 2972 - 0xb9c  :  252 - 0xfc
    "11111110", -- 2973 - 0xb9d  :  254 - 0xfe
    "01010100", -- 2974 - 0xb9e  :   84 - 0x54
    "00000000", -- 2975 - 0xb9f  :    0 - 0x0
    "11111111", -- 2976 - 0xba0  :  255 - 0xff -- Background 0xba
    "11010101", -- 2977 - 0xba1  :  213 - 0xd5
    "10101010", -- 2978 - 0xba2  :  170 - 0xaa
    "11111111", -- 2979 - 0xba3  :  255 - 0xff
    "10000000", -- 2980 - 0xba4  :  128 - 0x80
    "10000000", -- 2981 - 0xba5  :  128 - 0x80
    "10010101", -- 2982 - 0xba6  :  149 - 0x95
    "11111111", -- 2983 - 0xba7  :  255 - 0xff
    "00000000", -- 2984 - 0xba8  :    0 - 0x0 -- plane 1
    "01111111", -- 2985 - 0xba9  :  127 - 0x7f
    "01111111", -- 2986 - 0xbaa  :  127 - 0x7f
    "00000000", -- 2987 - 0xbab  :    0 - 0x0
    "01111111", -- 2988 - 0xbac  :  127 - 0x7f
    "01111111", -- 2989 - 0xbad  :  127 - 0x7f
    "01101010", -- 2990 - 0xbae  :  106 - 0x6a
    "00000000", -- 2991 - 0xbaf  :    0 - 0x0
    "00000000", -- 2992 - 0xbb0  :    0 - 0x0 -- Background 0xbb
    "00000000", -- 2993 - 0xbb1  :    0 - 0x0
    "00000000", -- 2994 - 0xbb2  :    0 - 0x0
    "00000000", -- 2995 - 0xbb3  :    0 - 0x0
    "00000000", -- 2996 - 0xbb4  :    0 - 0x0
    "00000000", -- 2997 - 0xbb5  :    0 - 0x0
    "00000000", -- 2998 - 0xbb6  :    0 - 0x0
    "00000000", -- 2999 - 0xbb7  :    0 - 0x0
    "00000000", -- 3000 - 0xbb8  :    0 - 0x0 -- plane 1
    "00000000", -- 3001 - 0xbb9  :    0 - 0x0
    "00000000", -- 3002 - 0xbba  :    0 - 0x0
    "00000000", -- 3003 - 0xbbb  :    0 - 0x0
    "00000000", -- 3004 - 0xbbc  :    0 - 0x0
    "00000000", -- 3005 - 0xbbd  :    0 - 0x0
    "00000000", -- 3006 - 0xbbe  :    0 - 0x0
    "00000000", -- 3007 - 0xbbf  :    0 - 0x0
    "11111111", -- 3008 - 0xbc0  :  255 - 0xff -- Background 0xbc
    "01010101", -- 3009 - 0xbc1  :   85 - 0x55
    "10101011", -- 3010 - 0xbc2  :  171 - 0xab
    "11111111", -- 3011 - 0xbc3  :  255 - 0xff
    "01100001", -- 3012 - 0xbc4  :   97 - 0x61
    "00100011", -- 3013 - 0xbc5  :   35 - 0x23
    "01100101", -- 3014 - 0xbc6  :  101 - 0x65
    "11111111", -- 3015 - 0xbc7  :  255 - 0xff
    "00000000", -- 3016 - 0xbc8  :    0 - 0x0 -- plane 1
    "11111110", -- 3017 - 0xbc9  :  254 - 0xfe
    "11111110", -- 3018 - 0xbca  :  254 - 0xfe
    "00000000", -- 3019 - 0xbcb  :    0 - 0x0
    "10011110", -- 3020 - 0xbcc  :  158 - 0x9e
    "11011100", -- 3021 - 0xbcd  :  220 - 0xdc
    "10011010", -- 3022 - 0xbce  :  154 - 0x9a
    "00000000", -- 3023 - 0xbcf  :    0 - 0x0
    "00000000", -- 3024 - 0xbd0  :    0 - 0x0 -- Background 0xbd
    "00000000", -- 3025 - 0xbd1  :    0 - 0x0
    "00000000", -- 3026 - 0xbd2  :    0 - 0x0
    "00000000", -- 3027 - 0xbd3  :    0 - 0x0
    "00000000", -- 3028 - 0xbd4  :    0 - 0x0
    "00000000", -- 3029 - 0xbd5  :    0 - 0x0
    "00000000", -- 3030 - 0xbd6  :    0 - 0x0
    "00000000", -- 3031 - 0xbd7  :    0 - 0x0
    "00000000", -- 3032 - 0xbd8  :    0 - 0x0 -- plane 1
    "00000000", -- 3033 - 0xbd9  :    0 - 0x0
    "00000000", -- 3034 - 0xbda  :    0 - 0x0
    "00000000", -- 3035 - 0xbdb  :    0 - 0x0
    "00000000", -- 3036 - 0xbdc  :    0 - 0x0
    "00000000", -- 3037 - 0xbdd  :    0 - 0x0
    "00000000", -- 3038 - 0xbde  :    0 - 0x0
    "00000000", -- 3039 - 0xbdf  :    0 - 0x0
    "00000000", -- 3040 - 0xbe0  :    0 - 0x0 -- Background 0xbe
    "00000000", -- 3041 - 0xbe1  :    0 - 0x0
    "00000000", -- 3042 - 0xbe2  :    0 - 0x0
    "00000000", -- 3043 - 0xbe3  :    0 - 0x0
    "00000000", -- 3044 - 0xbe4  :    0 - 0x0
    "00000000", -- 3045 - 0xbe5  :    0 - 0x0
    "00000000", -- 3046 - 0xbe6  :    0 - 0x0
    "00000000", -- 3047 - 0xbe7  :    0 - 0x0
    "00000000", -- 3048 - 0xbe8  :    0 - 0x0 -- plane 1
    "00000000", -- 3049 - 0xbe9  :    0 - 0x0
    "00000000", -- 3050 - 0xbea  :    0 - 0x0
    "00000000", -- 3051 - 0xbeb  :    0 - 0x0
    "00000000", -- 3052 - 0xbec  :    0 - 0x0
    "00000000", -- 3053 - 0xbed  :    0 - 0x0
    "00000000", -- 3054 - 0xbee  :    0 - 0x0
    "00000000", -- 3055 - 0xbef  :    0 - 0x0
    "00000000", -- 3056 - 0xbf0  :    0 - 0x0 -- Background 0xbf
    "00000000", -- 3057 - 0xbf1  :    0 - 0x0
    "00000000", -- 3058 - 0xbf2  :    0 - 0x0
    "00000000", -- 3059 - 0xbf3  :    0 - 0x0
    "00000000", -- 3060 - 0xbf4  :    0 - 0x0
    "00000000", -- 3061 - 0xbf5  :    0 - 0x0
    "00000000", -- 3062 - 0xbf6  :    0 - 0x0
    "00000000", -- 3063 - 0xbf7  :    0 - 0x0
    "00000000", -- 3064 - 0xbf8  :    0 - 0x0 -- plane 1
    "00000000", -- 3065 - 0xbf9  :    0 - 0x0
    "00000000", -- 3066 - 0xbfa  :    0 - 0x0
    "00000000", -- 3067 - 0xbfb  :    0 - 0x0
    "00000000", -- 3068 - 0xbfc  :    0 - 0x0
    "00000000", -- 3069 - 0xbfd  :    0 - 0x0
    "00000000", -- 3070 - 0xbfe  :    0 - 0x0
    "00000000", -- 3071 - 0xbff  :    0 - 0x0
    "00000000", -- 3072 - 0xc00  :    0 - 0x0 -- Background 0xc0
    "00000000", -- 3073 - 0xc01  :    0 - 0x0
    "00000000", -- 3074 - 0xc02  :    0 - 0x0
    "00000000", -- 3075 - 0xc03  :    0 - 0x0
    "00000000", -- 3076 - 0xc04  :    0 - 0x0
    "00000000", -- 3077 - 0xc05  :    0 - 0x0
    "00000000", -- 3078 - 0xc06  :    0 - 0x0
    "00000000", -- 3079 - 0xc07  :    0 - 0x0
    "00000000", -- 3080 - 0xc08  :    0 - 0x0 -- plane 1
    "00000000", -- 3081 - 0xc09  :    0 - 0x0
    "00000000", -- 3082 - 0xc0a  :    0 - 0x0
    "00000000", -- 3083 - 0xc0b  :    0 - 0x0
    "00000000", -- 3084 - 0xc0c  :    0 - 0x0
    "00000000", -- 3085 - 0xc0d  :    0 - 0x0
    "00000000", -- 3086 - 0xc0e  :    0 - 0x0
    "00000000", -- 3087 - 0xc0f  :    0 - 0x0
    "00000000", -- 3088 - 0xc10  :    0 - 0x0 -- Background 0xc1
    "00000000", -- 3089 - 0xc11  :    0 - 0x0
    "00000000", -- 3090 - 0xc12  :    0 - 0x0
    "00000000", -- 3091 - 0xc13  :    0 - 0x0
    "00000000", -- 3092 - 0xc14  :    0 - 0x0
    "00000000", -- 3093 - 0xc15  :    0 - 0x0
    "00000000", -- 3094 - 0xc16  :    0 - 0x0
    "00000000", -- 3095 - 0xc17  :    0 - 0x0
    "00000000", -- 3096 - 0xc18  :    0 - 0x0 -- plane 1
    "00000000", -- 3097 - 0xc19  :    0 - 0x0
    "00000000", -- 3098 - 0xc1a  :    0 - 0x0
    "00000000", -- 3099 - 0xc1b  :    0 - 0x0
    "00000000", -- 3100 - 0xc1c  :    0 - 0x0
    "00000000", -- 3101 - 0xc1d  :    0 - 0x0
    "00000000", -- 3102 - 0xc1e  :    0 - 0x0
    "00000000", -- 3103 - 0xc1f  :    0 - 0x0
    "00000000", -- 3104 - 0xc20  :    0 - 0x0 -- Background 0xc2
    "00000000", -- 3105 - 0xc21  :    0 - 0x0
    "00000000", -- 3106 - 0xc22  :    0 - 0x0
    "00000000", -- 3107 - 0xc23  :    0 - 0x0
    "00000000", -- 3108 - 0xc24  :    0 - 0x0
    "00000000", -- 3109 - 0xc25  :    0 - 0x0
    "00000000", -- 3110 - 0xc26  :    0 - 0x0
    "00000000", -- 3111 - 0xc27  :    0 - 0x0
    "00000000", -- 3112 - 0xc28  :    0 - 0x0 -- plane 1
    "00000000", -- 3113 - 0xc29  :    0 - 0x0
    "00000000", -- 3114 - 0xc2a  :    0 - 0x0
    "00000000", -- 3115 - 0xc2b  :    0 - 0x0
    "00000000", -- 3116 - 0xc2c  :    0 - 0x0
    "00000000", -- 3117 - 0xc2d  :    0 - 0x0
    "00000000", -- 3118 - 0xc2e  :    0 - 0x0
    "00000000", -- 3119 - 0xc2f  :    0 - 0x0
    "00000000", -- 3120 - 0xc30  :    0 - 0x0 -- Background 0xc3
    "00000000", -- 3121 - 0xc31  :    0 - 0x0
    "00000000", -- 3122 - 0xc32  :    0 - 0x0
    "00000000", -- 3123 - 0xc33  :    0 - 0x0
    "00000000", -- 3124 - 0xc34  :    0 - 0x0
    "00000000", -- 3125 - 0xc35  :    0 - 0x0
    "00000000", -- 3126 - 0xc36  :    0 - 0x0
    "00000000", -- 3127 - 0xc37  :    0 - 0x0
    "00000000", -- 3128 - 0xc38  :    0 - 0x0 -- plane 1
    "00000000", -- 3129 - 0xc39  :    0 - 0x0
    "00000000", -- 3130 - 0xc3a  :    0 - 0x0
    "00000000", -- 3131 - 0xc3b  :    0 - 0x0
    "00000000", -- 3132 - 0xc3c  :    0 - 0x0
    "00000000", -- 3133 - 0xc3d  :    0 - 0x0
    "00000000", -- 3134 - 0xc3e  :    0 - 0x0
    "00000000", -- 3135 - 0xc3f  :    0 - 0x0
    "00000000", -- 3136 - 0xc40  :    0 - 0x0 -- Background 0xc4
    "00000000", -- 3137 - 0xc41  :    0 - 0x0
    "00000000", -- 3138 - 0xc42  :    0 - 0x0
    "00000000", -- 3139 - 0xc43  :    0 - 0x0
    "00000000", -- 3140 - 0xc44  :    0 - 0x0
    "00000000", -- 3141 - 0xc45  :    0 - 0x0
    "00000000", -- 3142 - 0xc46  :    0 - 0x0
    "00000000", -- 3143 - 0xc47  :    0 - 0x0
    "00000000", -- 3144 - 0xc48  :    0 - 0x0 -- plane 1
    "00000000", -- 3145 - 0xc49  :    0 - 0x0
    "00000000", -- 3146 - 0xc4a  :    0 - 0x0
    "00000000", -- 3147 - 0xc4b  :    0 - 0x0
    "00000000", -- 3148 - 0xc4c  :    0 - 0x0
    "00000000", -- 3149 - 0xc4d  :    0 - 0x0
    "00000000", -- 3150 - 0xc4e  :    0 - 0x0
    "00000000", -- 3151 - 0xc4f  :    0 - 0x0
    "00000000", -- 3152 - 0xc50  :    0 - 0x0 -- Background 0xc5
    "00000000", -- 3153 - 0xc51  :    0 - 0x0
    "00000001", -- 3154 - 0xc52  :    1 - 0x1
    "00000110", -- 3155 - 0xc53  :    6 - 0x6
    "00001010", -- 3156 - 0xc54  :   10 - 0xa
    "00010100", -- 3157 - 0xc55  :   20 - 0x14
    "00010000", -- 3158 - 0xc56  :   16 - 0x10
    "00101000", -- 3159 - 0xc57  :   40 - 0x28
    "00000000", -- 3160 - 0xc58  :    0 - 0x0 -- plane 1
    "00000000", -- 3161 - 0xc59  :    0 - 0x0
    "00000000", -- 3162 - 0xc5a  :    0 - 0x0
    "00000001", -- 3163 - 0xc5b  :    1 - 0x1
    "00000111", -- 3164 - 0xc5c  :    7 - 0x7
    "00001111", -- 3165 - 0xc5d  :   15 - 0xf
    "00001111", -- 3166 - 0xc5e  :   15 - 0xf
    "00011111", -- 3167 - 0xc5f  :   31 - 0x1f
    "00011111", -- 3168 - 0xc60  :   31 - 0x1f -- Background 0xc6
    "01100000", -- 3169 - 0xc61  :   96 - 0x60
    "10100000", -- 3170 - 0xc62  :  160 - 0xa0
    "01000000", -- 3171 - 0xc63  :   64 - 0x40
    "00000000", -- 3172 - 0xc64  :    0 - 0x0
    "00000000", -- 3173 - 0xc65  :    0 - 0x0
    "00000000", -- 3174 - 0xc66  :    0 - 0x0
    "00000000", -- 3175 - 0xc67  :    0 - 0x0
    "00000000", -- 3176 - 0xc68  :    0 - 0x0 -- plane 1
    "00011111", -- 3177 - 0xc69  :   31 - 0x1f
    "01111111", -- 3178 - 0xc6a  :  127 - 0x7f
    "11111111", -- 3179 - 0xc6b  :  255 - 0xff
    "11111111", -- 3180 - 0xc6c  :  255 - 0xff
    "11111111", -- 3181 - 0xc6d  :  255 - 0xff
    "11111111", -- 3182 - 0xc6e  :  255 - 0xff
    "11111111", -- 3183 - 0xc6f  :  255 - 0xff
    "00110000", -- 3184 - 0xc70  :   48 - 0x30 -- Background 0xc7
    "01000000", -- 3185 - 0xc71  :   64 - 0x40
    "01100000", -- 3186 - 0xc72  :   96 - 0x60
    "11000000", -- 3187 - 0xc73  :  192 - 0xc0
    "10000000", -- 3188 - 0xc74  :  128 - 0x80
    "10100000", -- 3189 - 0xc75  :  160 - 0xa0
    "11000000", -- 3190 - 0xc76  :  192 - 0xc0
    "10000000", -- 3191 - 0xc77  :  128 - 0x80
    "00011111", -- 3192 - 0xc78  :   31 - 0x1f -- plane 1
    "00111111", -- 3193 - 0xc79  :   63 - 0x3f
    "00111111", -- 3194 - 0xc7a  :   63 - 0x3f
    "01111111", -- 3195 - 0xc7b  :  127 - 0x7f
    "01111111", -- 3196 - 0xc7c  :  127 - 0x7f
    "01111111", -- 3197 - 0xc7d  :  127 - 0x7f
    "01111111", -- 3198 - 0xc7e  :  127 - 0x7f
    "01111111", -- 3199 - 0xc7f  :  127 - 0x7f
    "11111111", -- 3200 - 0xc80  :  255 - 0xff -- Background 0xc8
    "00000000", -- 3201 - 0xc81  :    0 - 0x0
    "00000000", -- 3202 - 0xc82  :    0 - 0x0
    "00000000", -- 3203 - 0xc83  :    0 - 0x0
    "00000000", -- 3204 - 0xc84  :    0 - 0x0
    "00000000", -- 3205 - 0xc85  :    0 - 0x0
    "00000000", -- 3206 - 0xc86  :    0 - 0x0
    "00000000", -- 3207 - 0xc87  :    0 - 0x0
    "00000000", -- 3208 - 0xc88  :    0 - 0x0 -- plane 1
    "11111111", -- 3209 - 0xc89  :  255 - 0xff
    "11111111", -- 3210 - 0xc8a  :  255 - 0xff
    "11111111", -- 3211 - 0xc8b  :  255 - 0xff
    "11111111", -- 3212 - 0xc8c  :  255 - 0xff
    "11111111", -- 3213 - 0xc8d  :  255 - 0xff
    "11111111", -- 3214 - 0xc8e  :  255 - 0xff
    "11111111", -- 3215 - 0xc8f  :  255 - 0xff
    "00010100", -- 3216 - 0xc90  :   20 - 0x14 -- Background 0xc9
    "00101010", -- 3217 - 0xc91  :   42 - 0x2a
    "00010110", -- 3218 - 0xc92  :   22 - 0x16
    "00101011", -- 3219 - 0xc93  :   43 - 0x2b
    "00010101", -- 3220 - 0xc94  :   21 - 0x15
    "00101011", -- 3221 - 0xc95  :   43 - 0x2b
    "00010101", -- 3222 - 0xc96  :   21 - 0x15
    "00101011", -- 3223 - 0xc97  :   43 - 0x2b
    "11101000", -- 3224 - 0xc98  :  232 - 0xe8 -- plane 1
    "11010100", -- 3225 - 0xc99  :  212 - 0xd4
    "11101000", -- 3226 - 0xc9a  :  232 - 0xe8
    "11010100", -- 3227 - 0xc9b  :  212 - 0xd4
    "11101010", -- 3228 - 0xc9c  :  234 - 0xea
    "11010100", -- 3229 - 0xc9d  :  212 - 0xd4
    "11101010", -- 3230 - 0xc9e  :  234 - 0xea
    "11010100", -- 3231 - 0xc9f  :  212 - 0xd4
    "00000000", -- 3232 - 0xca0  :    0 - 0x0 -- Background 0xca
    "00000100", -- 3233 - 0xca1  :    4 - 0x4
    "00000100", -- 3234 - 0xca2  :    4 - 0x4
    "00000101", -- 3235 - 0xca3  :    5 - 0x5
    "00010101", -- 3236 - 0xca4  :   21 - 0x15
    "00010101", -- 3237 - 0xca5  :   21 - 0x15
    "01010101", -- 3238 - 0xca6  :   85 - 0x55
    "01010101", -- 3239 - 0xca7  :   85 - 0x55
    "00000000", -- 3240 - 0xca8  :    0 - 0x0 -- plane 1
    "00000000", -- 3241 - 0xca9  :    0 - 0x0
    "00000000", -- 3242 - 0xcaa  :    0 - 0x0
    "00000000", -- 3243 - 0xcab  :    0 - 0x0
    "00000000", -- 3244 - 0xcac  :    0 - 0x0
    "00000000", -- 3245 - 0xcad  :    0 - 0x0
    "00000000", -- 3246 - 0xcae  :    0 - 0x0
    "00000000", -- 3247 - 0xcaf  :    0 - 0x0
    "00000000", -- 3248 - 0xcb0  :    0 - 0x0 -- Background 0xcb
    "00000000", -- 3249 - 0xcb1  :    0 - 0x0
    "00010000", -- 3250 - 0xcb2  :   16 - 0x10
    "00010000", -- 3251 - 0xcb3  :   16 - 0x10
    "01010001", -- 3252 - 0xcb4  :   81 - 0x51
    "01010101", -- 3253 - 0xcb5  :   85 - 0x55
    "01010101", -- 3254 - 0xcb6  :   85 - 0x55
    "01010101", -- 3255 - 0xcb7  :   85 - 0x55
    "00000000", -- 3256 - 0xcb8  :    0 - 0x0 -- plane 1
    "00000000", -- 3257 - 0xcb9  :    0 - 0x0
    "00000000", -- 3258 - 0xcba  :    0 - 0x0
    "00000000", -- 3259 - 0xcbb  :    0 - 0x0
    "00000000", -- 3260 - 0xcbc  :    0 - 0x0
    "00000000", -- 3261 - 0xcbd  :    0 - 0x0
    "00000000", -- 3262 - 0xcbe  :    0 - 0x0
    "00000000", -- 3263 - 0xcbf  :    0 - 0x0
    "00000000", -- 3264 - 0xcc0  :    0 - 0x0 -- Background 0xcc
    "00000000", -- 3265 - 0xcc1  :    0 - 0x0
    "00000000", -- 3266 - 0xcc2  :    0 - 0x0
    "00000101", -- 3267 - 0xcc3  :    5 - 0x5
    "00001111", -- 3268 - 0xcc4  :   15 - 0xf
    "00000111", -- 3269 - 0xcc5  :    7 - 0x7
    "00000011", -- 3270 - 0xcc6  :    3 - 0x3
    "00000001", -- 3271 - 0xcc7  :    1 - 0x1
    "00000000", -- 3272 - 0xcc8  :    0 - 0x0 -- plane 1
    "00000000", -- 3273 - 0xcc9  :    0 - 0x0
    "00000000", -- 3274 - 0xcca  :    0 - 0x0
    "00000000", -- 3275 - 0xccb  :    0 - 0x0
    "00000101", -- 3276 - 0xccc  :    5 - 0x5
    "00000010", -- 3277 - 0xccd  :    2 - 0x2
    "00000001", -- 3278 - 0xcce  :    1 - 0x1
    "00000000", -- 3279 - 0xccf  :    0 - 0x0
    "00000000", -- 3280 - 0xcd0  :    0 - 0x0 -- Background 0xcd
    "00000000", -- 3281 - 0xcd1  :    0 - 0x0
    "10000000", -- 3282 - 0xcd2  :  128 - 0x80
    "11010000", -- 3283 - 0xcd3  :  208 - 0xd0
    "11111000", -- 3284 - 0xcd4  :  248 - 0xf8
    "11110000", -- 3285 - 0xcd5  :  240 - 0xf0
    "11100000", -- 3286 - 0xcd6  :  224 - 0xe0
    "11000000", -- 3287 - 0xcd7  :  192 - 0xc0
    "00000000", -- 3288 - 0xcd8  :    0 - 0x0 -- plane 1
    "00000000", -- 3289 - 0xcd9  :    0 - 0x0
    "00000000", -- 3290 - 0xcda  :    0 - 0x0
    "10000000", -- 3291 - 0xcdb  :  128 - 0x80
    "01010000", -- 3292 - 0xcdc  :   80 - 0x50
    "10100000", -- 3293 - 0xcdd  :  160 - 0xa0
    "01000000", -- 3294 - 0xcde  :   64 - 0x40
    "10000000", -- 3295 - 0xcdf  :  128 - 0x80
    "00000000", -- 3296 - 0xce0  :    0 - 0x0 -- Background 0xce
    "00000000", -- 3297 - 0xce1  :    0 - 0x0
    "00000000", -- 3298 - 0xce2  :    0 - 0x0
    "01111000", -- 3299 - 0xce3  :  120 - 0x78
    "11001111", -- 3300 - 0xce4  :  207 - 0xcf
    "10000000", -- 3301 - 0xce5  :  128 - 0x80
    "11001111", -- 3302 - 0xce6  :  207 - 0xcf
    "01001000", -- 3303 - 0xce7  :   72 - 0x48
    "00000000", -- 3304 - 0xce8  :    0 - 0x0 -- plane 1
    "00000000", -- 3305 - 0xce9  :    0 - 0x0
    "00000000", -- 3306 - 0xcea  :    0 - 0x0
    "00000000", -- 3307 - 0xceb  :    0 - 0x0
    "00110000", -- 3308 - 0xcec  :   48 - 0x30
    "01111111", -- 3309 - 0xced  :  127 - 0x7f
    "00110000", -- 3310 - 0xcee  :   48 - 0x30
    "00110000", -- 3311 - 0xcef  :   48 - 0x30
    "00000000", -- 3312 - 0xcf0  :    0 - 0x0 -- Background 0xcf
    "00000000", -- 3313 - 0xcf1  :    0 - 0x0
    "00000000", -- 3314 - 0xcf2  :    0 - 0x0
    "00011110", -- 3315 - 0xcf3  :   30 - 0x1e
    "11110011", -- 3316 - 0xcf4  :  243 - 0xf3
    "00000001", -- 3317 - 0xcf5  :    1 - 0x1
    "11110011", -- 3318 - 0xcf6  :  243 - 0xf3
    "00010010", -- 3319 - 0xcf7  :   18 - 0x12
    "00000000", -- 3320 - 0xcf8  :    0 - 0x0 -- plane 1
    "00000000", -- 3321 - 0xcf9  :    0 - 0x0
    "00000000", -- 3322 - 0xcfa  :    0 - 0x0
    "00000000", -- 3323 - 0xcfb  :    0 - 0x0
    "00001100", -- 3324 - 0xcfc  :   12 - 0xc
    "11111110", -- 3325 - 0xcfd  :  254 - 0xfe
    "00001100", -- 3326 - 0xcfe  :   12 - 0xc
    "00001100", -- 3327 - 0xcff  :   12 - 0xc
    "00000000", -- 3328 - 0xd00  :    0 - 0x0 -- Background 0xd0
    "00000000", -- 3329 - 0xd01  :    0 - 0x0
    "00000000", -- 3330 - 0xd02  :    0 - 0x0
    "00000000", -- 3331 - 0xd03  :    0 - 0x0
    "00000000", -- 3332 - 0xd04  :    0 - 0x0
    "00000000", -- 3333 - 0xd05  :    0 - 0x0
    "00000000", -- 3334 - 0xd06  :    0 - 0x0
    "00000000", -- 3335 - 0xd07  :    0 - 0x0
    "00000000", -- 3336 - 0xd08  :    0 - 0x0 -- plane 1
    "00000000", -- 3337 - 0xd09  :    0 - 0x0
    "00000000", -- 3338 - 0xd0a  :    0 - 0x0
    "00000000", -- 3339 - 0xd0b  :    0 - 0x0
    "00000000", -- 3340 - 0xd0c  :    0 - 0x0
    "00000000", -- 3341 - 0xd0d  :    0 - 0x0
    "00000000", -- 3342 - 0xd0e  :    0 - 0x0
    "00000000", -- 3343 - 0xd0f  :    0 - 0x0
    "00000000", -- 3344 - 0xd10  :    0 - 0x0 -- Background 0xd1
    "00000000", -- 3345 - 0xd11  :    0 - 0x0
    "00000000", -- 3346 - 0xd12  :    0 - 0x0
    "00000000", -- 3347 - 0xd13  :    0 - 0x0
    "00000000", -- 3348 - 0xd14  :    0 - 0x0
    "00000000", -- 3349 - 0xd15  :    0 - 0x0
    "00000000", -- 3350 - 0xd16  :    0 - 0x0
    "00000000", -- 3351 - 0xd17  :    0 - 0x0
    "00000000", -- 3352 - 0xd18  :    0 - 0x0 -- plane 1
    "00000000", -- 3353 - 0xd19  :    0 - 0x0
    "00000000", -- 3354 - 0xd1a  :    0 - 0x0
    "00000000", -- 3355 - 0xd1b  :    0 - 0x0
    "00000000", -- 3356 - 0xd1c  :    0 - 0x0
    "00000000", -- 3357 - 0xd1d  :    0 - 0x0
    "00000000", -- 3358 - 0xd1e  :    0 - 0x0
    "00000000", -- 3359 - 0xd1f  :    0 - 0x0
    "00001000", -- 3360 - 0xd20  :    8 - 0x8 -- Background 0xd2
    "00001100", -- 3361 - 0xd21  :   12 - 0xc
    "00001000", -- 3362 - 0xd22  :    8 - 0x8
    "00001000", -- 3363 - 0xd23  :    8 - 0x8
    "00001010", -- 3364 - 0xd24  :   10 - 0xa
    "00001000", -- 3365 - 0xd25  :    8 - 0x8
    "00001000", -- 3366 - 0xd26  :    8 - 0x8
    "00001100", -- 3367 - 0xd27  :   12 - 0xc
    "00000111", -- 3368 - 0xd28  :    7 - 0x7 -- plane 1
    "00000111", -- 3369 - 0xd29  :    7 - 0x7
    "00000111", -- 3370 - 0xd2a  :    7 - 0x7
    "00000111", -- 3371 - 0xd2b  :    7 - 0x7
    "00000111", -- 3372 - 0xd2c  :    7 - 0x7
    "00000111", -- 3373 - 0xd2d  :    7 - 0x7
    "00000111", -- 3374 - 0xd2e  :    7 - 0x7
    "00000111", -- 3375 - 0xd2f  :    7 - 0x7
    "00010000", -- 3376 - 0xd30  :   16 - 0x10 -- Background 0xd3
    "00010000", -- 3377 - 0xd31  :   16 - 0x10
    "00110000", -- 3378 - 0xd32  :   48 - 0x30
    "00010000", -- 3379 - 0xd33  :   16 - 0x10
    "01010000", -- 3380 - 0xd34  :   80 - 0x50
    "00010000", -- 3381 - 0xd35  :   16 - 0x10
    "00110000", -- 3382 - 0xd36  :   48 - 0x30
    "00010000", -- 3383 - 0xd37  :   16 - 0x10
    "11100000", -- 3384 - 0xd38  :  224 - 0xe0 -- plane 1
    "11100000", -- 3385 - 0xd39  :  224 - 0xe0
    "11000000", -- 3386 - 0xd3a  :  192 - 0xc0
    "11100000", -- 3387 - 0xd3b  :  224 - 0xe0
    "10100000", -- 3388 - 0xd3c  :  160 - 0xa0
    "11100000", -- 3389 - 0xd3d  :  224 - 0xe0
    "11000000", -- 3390 - 0xd3e  :  192 - 0xc0
    "11100000", -- 3391 - 0xd3f  :  224 - 0xe0
    "00000000", -- 3392 - 0xd40  :    0 - 0x0 -- Background 0xd4
    "00000000", -- 3393 - 0xd41  :    0 - 0x0
    "00000000", -- 3394 - 0xd42  :    0 - 0x0
    "00000000", -- 3395 - 0xd43  :    0 - 0x0
    "00000000", -- 3396 - 0xd44  :    0 - 0x0
    "00000000", -- 3397 - 0xd45  :    0 - 0x0
    "00000000", -- 3398 - 0xd46  :    0 - 0x0
    "00000000", -- 3399 - 0xd47  :    0 - 0x0
    "00000000", -- 3400 - 0xd48  :    0 - 0x0 -- plane 1
    "00000000", -- 3401 - 0xd49  :    0 - 0x0
    "00000000", -- 3402 - 0xd4a  :    0 - 0x0
    "00000000", -- 3403 - 0xd4b  :    0 - 0x0
    "00000000", -- 3404 - 0xd4c  :    0 - 0x0
    "00000000", -- 3405 - 0xd4d  :    0 - 0x0
    "00000000", -- 3406 - 0xd4e  :    0 - 0x0
    "00000000", -- 3407 - 0xd4f  :    0 - 0x0
    "11111000", -- 3408 - 0xd50  :  248 - 0xf8 -- Background 0xd5
    "00000110", -- 3409 - 0xd51  :    6 - 0x6
    "00000001", -- 3410 - 0xd52  :    1 - 0x1
    "00000000", -- 3411 - 0xd53  :    0 - 0x0
    "00000000", -- 3412 - 0xd54  :    0 - 0x0
    "00000000", -- 3413 - 0xd55  :    0 - 0x0
    "00000000", -- 3414 - 0xd56  :    0 - 0x0
    "00000000", -- 3415 - 0xd57  :    0 - 0x0
    "00000000", -- 3416 - 0xd58  :    0 - 0x0 -- plane 1
    "11111000", -- 3417 - 0xd59  :  248 - 0xf8
    "11111110", -- 3418 - 0xd5a  :  254 - 0xfe
    "11111111", -- 3419 - 0xd5b  :  255 - 0xff
    "11111111", -- 3420 - 0xd5c  :  255 - 0xff
    "11111111", -- 3421 - 0xd5d  :  255 - 0xff
    "11111111", -- 3422 - 0xd5e  :  255 - 0xff
    "11111111", -- 3423 - 0xd5f  :  255 - 0xff
    "00000000", -- 3424 - 0xd60  :    0 - 0x0 -- Background 0xd6
    "00000000", -- 3425 - 0xd61  :    0 - 0x0
    "10000000", -- 3426 - 0xd62  :  128 - 0x80
    "01100000", -- 3427 - 0xd63  :   96 - 0x60
    "01010000", -- 3428 - 0xd64  :   80 - 0x50
    "10101000", -- 3429 - 0xd65  :  168 - 0xa8
    "01011000", -- 3430 - 0xd66  :   88 - 0x58
    "00101100", -- 3431 - 0xd67  :   44 - 0x2c
    "00000000", -- 3432 - 0xd68  :    0 - 0x0 -- plane 1
    "00000000", -- 3433 - 0xd69  :    0 - 0x0
    "00000000", -- 3434 - 0xd6a  :    0 - 0x0
    "10000000", -- 3435 - 0xd6b  :  128 - 0x80
    "10100000", -- 3436 - 0xd6c  :  160 - 0xa0
    "01010000", -- 3437 - 0xd6d  :   80 - 0x50
    "10100000", -- 3438 - 0xd6e  :  160 - 0xa0
    "11010000", -- 3439 - 0xd6f  :  208 - 0xd0
    "10100000", -- 3440 - 0xd70  :  160 - 0xa0 -- Background 0xd7
    "11000000", -- 3441 - 0xd71  :  192 - 0xc0
    "10000000", -- 3442 - 0xd72  :  128 - 0x80
    "01010000", -- 3443 - 0xd73  :   80 - 0x50
    "01100000", -- 3444 - 0xd74  :   96 - 0x60
    "00111000", -- 3445 - 0xd75  :   56 - 0x38
    "00001000", -- 3446 - 0xd76  :    8 - 0x8
    "00000111", -- 3447 - 0xd77  :    7 - 0x7
    "01111111", -- 3448 - 0xd78  :  127 - 0x7f -- plane 1
    "01111111", -- 3449 - 0xd79  :  127 - 0x7f
    "01111111", -- 3450 - 0xd7a  :  127 - 0x7f
    "00111111", -- 3451 - 0xd7b  :   63 - 0x3f
    "00111111", -- 3452 - 0xd7c  :   63 - 0x3f
    "00001111", -- 3453 - 0xd7d  :   15 - 0xf
    "00000111", -- 3454 - 0xd7e  :    7 - 0x7
    "00000000", -- 3455 - 0xd7f  :    0 - 0x0
    "00000000", -- 3456 - 0xd80  :    0 - 0x0 -- Background 0xd8
    "00000000", -- 3457 - 0xd81  :    0 - 0x0
    "00000000", -- 3458 - 0xd82  :    0 - 0x0
    "00000000", -- 3459 - 0xd83  :    0 - 0x0
    "00000000", -- 3460 - 0xd84  :    0 - 0x0
    "00000000", -- 3461 - 0xd85  :    0 - 0x0
    "00000000", -- 3462 - 0xd86  :    0 - 0x0
    "11111111", -- 3463 - 0xd87  :  255 - 0xff
    "11111111", -- 3464 - 0xd88  :  255 - 0xff -- plane 1
    "11111111", -- 3465 - 0xd89  :  255 - 0xff
    "11111111", -- 3466 - 0xd8a  :  255 - 0xff
    "11111111", -- 3467 - 0xd8b  :  255 - 0xff
    "11111111", -- 3468 - 0xd8c  :  255 - 0xff
    "11111111", -- 3469 - 0xd8d  :  255 - 0xff
    "11111111", -- 3470 - 0xd8e  :  255 - 0xff
    "00000000", -- 3471 - 0xd8f  :    0 - 0x0
    "00010101", -- 3472 - 0xd90  :   21 - 0x15 -- Background 0xd9
    "00101011", -- 3473 - 0xd91  :   43 - 0x2b
    "00010101", -- 3474 - 0xd92  :   21 - 0x15
    "00101010", -- 3475 - 0xd93  :   42 - 0x2a
    "01010110", -- 3476 - 0xd94  :   86 - 0x56
    "10101100", -- 3477 - 0xd95  :  172 - 0xac
    "01010000", -- 3478 - 0xd96  :   80 - 0x50
    "11100000", -- 3479 - 0xd97  :  224 - 0xe0
    "11101010", -- 3480 - 0xd98  :  234 - 0xea -- plane 1
    "11010100", -- 3481 - 0xd99  :  212 - 0xd4
    "11101010", -- 3482 - 0xd9a  :  234 - 0xea
    "11010100", -- 3483 - 0xd9b  :  212 - 0xd4
    "10101000", -- 3484 - 0xd9c  :  168 - 0xa8
    "01010000", -- 3485 - 0xd9d  :   80 - 0x50
    "10100000", -- 3486 - 0xd9e  :  160 - 0xa0
    "00000000", -- 3487 - 0xd9f  :    0 - 0x0
    "00000001", -- 3488 - 0xda0  :    1 - 0x1 -- Background 0xda
    "00001101", -- 3489 - 0xda1  :   13 - 0xd
    "00010011", -- 3490 - 0xda2  :   19 - 0x13
    "00001101", -- 3491 - 0xda3  :   13 - 0xd
    "00000001", -- 3492 - 0xda4  :    1 - 0x1
    "00000001", -- 3493 - 0xda5  :    1 - 0x1
    "00000001", -- 3494 - 0xda6  :    1 - 0x1
    "00000001", -- 3495 - 0xda7  :    1 - 0x1
    "00000000", -- 3496 - 0xda8  :    0 - 0x0 -- plane 1
    "00000000", -- 3497 - 0xda9  :    0 - 0x0
    "00001100", -- 3498 - 0xdaa  :   12 - 0xc
    "00000000", -- 3499 - 0xdab  :    0 - 0x0
    "00000000", -- 3500 - 0xdac  :    0 - 0x0
    "00000000", -- 3501 - 0xdad  :    0 - 0x0
    "00000000", -- 3502 - 0xdae  :    0 - 0x0
    "00000000", -- 3503 - 0xdaf  :    0 - 0x0
    "11000000", -- 3504 - 0xdb0  :  192 - 0xc0 -- Background 0xdb
    "01000000", -- 3505 - 0xdb1  :   64 - 0x40
    "01000000", -- 3506 - 0xdb2  :   64 - 0x40
    "01011000", -- 3507 - 0xdb3  :   88 - 0x58
    "01100100", -- 3508 - 0xdb4  :  100 - 0x64
    "01011000", -- 3509 - 0xdb5  :   88 - 0x58
    "01000000", -- 3510 - 0xdb6  :   64 - 0x40
    "01000000", -- 3511 - 0xdb7  :   64 - 0x40
    "00000000", -- 3512 - 0xdb8  :    0 - 0x0 -- plane 1
    "10000000", -- 3513 - 0xdb9  :  128 - 0x80
    "10000000", -- 3514 - 0xdba  :  128 - 0x80
    "10000000", -- 3515 - 0xdbb  :  128 - 0x80
    "10011000", -- 3516 - 0xdbc  :  152 - 0x98
    "10000000", -- 3517 - 0xdbd  :  128 - 0x80
    "10000000", -- 3518 - 0xdbe  :  128 - 0x80
    "10000000", -- 3519 - 0xdbf  :  128 - 0x80
    "00000000", -- 3520 - 0xdc0  :    0 - 0x0 -- Background 0xdc
    "00000000", -- 3521 - 0xdc1  :    0 - 0x0
    "00000000", -- 3522 - 0xdc2  :    0 - 0x0
    "00000110", -- 3523 - 0xdc3  :    6 - 0x6
    "00000111", -- 3524 - 0xdc4  :    7 - 0x7
    "00000111", -- 3525 - 0xdc5  :    7 - 0x7
    "00000111", -- 3526 - 0xdc6  :    7 - 0x7
    "00000011", -- 3527 - 0xdc7  :    3 - 0x3
    "00000000", -- 3528 - 0xdc8  :    0 - 0x0 -- plane 1
    "00000000", -- 3529 - 0xdc9  :    0 - 0x0
    "00000000", -- 3530 - 0xdca  :    0 - 0x0
    "00000000", -- 3531 - 0xdcb  :    0 - 0x0
    "00000010", -- 3532 - 0xdcc  :    2 - 0x2
    "00000011", -- 3533 - 0xdcd  :    3 - 0x3
    "00000011", -- 3534 - 0xdce  :    3 - 0x3
    "00000001", -- 3535 - 0xdcf  :    1 - 0x1
    "00000000", -- 3536 - 0xdd0  :    0 - 0x0 -- Background 0xdd
    "00000000", -- 3537 - 0xdd1  :    0 - 0x0
    "00000000", -- 3538 - 0xdd2  :    0 - 0x0
    "10110000", -- 3539 - 0xdd3  :  176 - 0xb0
    "11110000", -- 3540 - 0xdd4  :  240 - 0xf0
    "11110000", -- 3541 - 0xdd5  :  240 - 0xf0
    "11110000", -- 3542 - 0xdd6  :  240 - 0xf0
    "11100000", -- 3543 - 0xdd7  :  224 - 0xe0
    "00000000", -- 3544 - 0xdd8  :    0 - 0x0 -- plane 1
    "00000000", -- 3545 - 0xdd9  :    0 - 0x0
    "00000000", -- 3546 - 0xdda  :    0 - 0x0
    "00000000", -- 3547 - 0xddb  :    0 - 0x0
    "10100000", -- 3548 - 0xddc  :  160 - 0xa0
    "11100000", -- 3549 - 0xddd  :  224 - 0xe0
    "11100000", -- 3550 - 0xdde  :  224 - 0xe0
    "11000000", -- 3551 - 0xddf  :  192 - 0xc0
    "11001111", -- 3552 - 0xde0  :  207 - 0xcf -- Background 0xde
    "10000000", -- 3553 - 0xde1  :  128 - 0x80
    "11001111", -- 3554 - 0xde2  :  207 - 0xcf
    "01001000", -- 3555 - 0xde3  :   72 - 0x48
    "01001000", -- 3556 - 0xde4  :   72 - 0x48
    "01001000", -- 3557 - 0xde5  :   72 - 0x48
    "01001000", -- 3558 - 0xde6  :   72 - 0x48
    "01001000", -- 3559 - 0xde7  :   72 - 0x48
    "00110000", -- 3560 - 0xde8  :   48 - 0x30 -- plane 1
    "01111111", -- 3561 - 0xde9  :  127 - 0x7f
    "00110000", -- 3562 - 0xdea  :   48 - 0x30
    "00110000", -- 3563 - 0xdeb  :   48 - 0x30
    "00110000", -- 3564 - 0xdec  :   48 - 0x30
    "00110000", -- 3565 - 0xded  :   48 - 0x30
    "00110000", -- 3566 - 0xdee  :   48 - 0x30
    "00110000", -- 3567 - 0xdef  :   48 - 0x30
    "11110011", -- 3568 - 0xdf0  :  243 - 0xf3 -- Background 0xdf
    "00000001", -- 3569 - 0xdf1  :    1 - 0x1
    "11110011", -- 3570 - 0xdf2  :  243 - 0xf3
    "00010010", -- 3571 - 0xdf3  :   18 - 0x12
    "00010010", -- 3572 - 0xdf4  :   18 - 0x12
    "00010010", -- 3573 - 0xdf5  :   18 - 0x12
    "00010010", -- 3574 - 0xdf6  :   18 - 0x12
    "00010010", -- 3575 - 0xdf7  :   18 - 0x12
    "00001100", -- 3576 - 0xdf8  :   12 - 0xc -- plane 1
    "11111110", -- 3577 - 0xdf9  :  254 - 0xfe
    "00001100", -- 3578 - 0xdfa  :   12 - 0xc
    "00001100", -- 3579 - 0xdfb  :   12 - 0xc
    "00001100", -- 3580 - 0xdfc  :   12 - 0xc
    "00001100", -- 3581 - 0xdfd  :   12 - 0xc
    "00001100", -- 3582 - 0xdfe  :   12 - 0xc
    "00001100", -- 3583 - 0xdff  :   12 - 0xc
    "00000000", -- 3584 - 0xe00  :    0 - 0x0 -- Background 0xe0
    "00000000", -- 3585 - 0xe01  :    0 - 0x0
    "00000000", -- 3586 - 0xe02  :    0 - 0x0
    "00000000", -- 3587 - 0xe03  :    0 - 0x0
    "00000000", -- 3588 - 0xe04  :    0 - 0x0
    "00000000", -- 3589 - 0xe05  :    0 - 0x0
    "00000000", -- 3590 - 0xe06  :    0 - 0x0
    "00000000", -- 3591 - 0xe07  :    0 - 0x0
    "00000000", -- 3592 - 0xe08  :    0 - 0x0 -- plane 1
    "00000000", -- 3593 - 0xe09  :    0 - 0x0
    "00000000", -- 3594 - 0xe0a  :    0 - 0x0
    "00000000", -- 3595 - 0xe0b  :    0 - 0x0
    "00000000", -- 3596 - 0xe0c  :    0 - 0x0
    "00000000", -- 3597 - 0xe0d  :    0 - 0x0
    "00000000", -- 3598 - 0xe0e  :    0 - 0x0
    "00000000", -- 3599 - 0xe0f  :    0 - 0x0
    "00000000", -- 3600 - 0xe10  :    0 - 0x0 -- Background 0xe1
    "00000000", -- 3601 - 0xe11  :    0 - 0x0
    "00000000", -- 3602 - 0xe12  :    0 - 0x0
    "00000000", -- 3603 - 0xe13  :    0 - 0x0
    "00000000", -- 3604 - 0xe14  :    0 - 0x0
    "00000000", -- 3605 - 0xe15  :    0 - 0x0
    "00000000", -- 3606 - 0xe16  :    0 - 0x0
    "00000000", -- 3607 - 0xe17  :    0 - 0x0
    "00000000", -- 3608 - 0xe18  :    0 - 0x0 -- plane 1
    "00000000", -- 3609 - 0xe19  :    0 - 0x0
    "00000000", -- 3610 - 0xe1a  :    0 - 0x0
    "00000000", -- 3611 - 0xe1b  :    0 - 0x0
    "00000000", -- 3612 - 0xe1c  :    0 - 0x0
    "00000000", -- 3613 - 0xe1d  :    0 - 0x0
    "00000000", -- 3614 - 0xe1e  :    0 - 0x0
    "00000000", -- 3615 - 0xe1f  :    0 - 0x0
    "00000000", -- 3616 - 0xe20  :    0 - 0x0 -- Background 0xe2
    "00000000", -- 3617 - 0xe21  :    0 - 0x0
    "00000000", -- 3618 - 0xe22  :    0 - 0x0
    "00000000", -- 3619 - 0xe23  :    0 - 0x0
    "00000000", -- 3620 - 0xe24  :    0 - 0x0
    "00000000", -- 3621 - 0xe25  :    0 - 0x0
    "00000000", -- 3622 - 0xe26  :    0 - 0x0
    "00000000", -- 3623 - 0xe27  :    0 - 0x0
    "00000000", -- 3624 - 0xe28  :    0 - 0x0 -- plane 1
    "00000000", -- 3625 - 0xe29  :    0 - 0x0
    "00000000", -- 3626 - 0xe2a  :    0 - 0x0
    "00000000", -- 3627 - 0xe2b  :    0 - 0x0
    "00000000", -- 3628 - 0xe2c  :    0 - 0x0
    "00000000", -- 3629 - 0xe2d  :    0 - 0x0
    "00000000", -- 3630 - 0xe2e  :    0 - 0x0
    "00000000", -- 3631 - 0xe2f  :    0 - 0x0
    "00000000", -- 3632 - 0xe30  :    0 - 0x0 -- Background 0xe3
    "00000000", -- 3633 - 0xe31  :    0 - 0x0
    "00000000", -- 3634 - 0xe32  :    0 - 0x0
    "00000000", -- 3635 - 0xe33  :    0 - 0x0
    "00000000", -- 3636 - 0xe34  :    0 - 0x0
    "00000000", -- 3637 - 0xe35  :    0 - 0x0
    "00000000", -- 3638 - 0xe36  :    0 - 0x0
    "00000000", -- 3639 - 0xe37  :    0 - 0x0
    "00000000", -- 3640 - 0xe38  :    0 - 0x0 -- plane 1
    "00000000", -- 3641 - 0xe39  :    0 - 0x0
    "00000000", -- 3642 - 0xe3a  :    0 - 0x0
    "00000000", -- 3643 - 0xe3b  :    0 - 0x0
    "00000000", -- 3644 - 0xe3c  :    0 - 0x0
    "00000000", -- 3645 - 0xe3d  :    0 - 0x0
    "00000000", -- 3646 - 0xe3e  :    0 - 0x0
    "00000000", -- 3647 - 0xe3f  :    0 - 0x0
    "00000000", -- 3648 - 0xe40  :    0 - 0x0 -- Background 0xe4
    "00000000", -- 3649 - 0xe41  :    0 - 0x0
    "00000000", -- 3650 - 0xe42  :    0 - 0x0
    "00000000", -- 3651 - 0xe43  :    0 - 0x0
    "00000000", -- 3652 - 0xe44  :    0 - 0x0
    "00000000", -- 3653 - 0xe45  :    0 - 0x0
    "00000000", -- 3654 - 0xe46  :    0 - 0x0
    "00000000", -- 3655 - 0xe47  :    0 - 0x0
    "00000000", -- 3656 - 0xe48  :    0 - 0x0 -- plane 1
    "00000000", -- 3657 - 0xe49  :    0 - 0x0
    "00000000", -- 3658 - 0xe4a  :    0 - 0x0
    "00000000", -- 3659 - 0xe4b  :    0 - 0x0
    "00000000", -- 3660 - 0xe4c  :    0 - 0x0
    "00000000", -- 3661 - 0xe4d  :    0 - 0x0
    "00000000", -- 3662 - 0xe4e  :    0 - 0x0
    "00000000", -- 3663 - 0xe4f  :    0 - 0x0
    "00000000", -- 3664 - 0xe50  :    0 - 0x0 -- Background 0xe5
    "00000000", -- 3665 - 0xe51  :    0 - 0x0
    "00000000", -- 3666 - 0xe52  :    0 - 0x0
    "00000000", -- 3667 - 0xe53  :    0 - 0x0
    "00000000", -- 3668 - 0xe54  :    0 - 0x0
    "00000000", -- 3669 - 0xe55  :    0 - 0x0
    "00000000", -- 3670 - 0xe56  :    0 - 0x0
    "00000000", -- 3671 - 0xe57  :    0 - 0x0
    "00000000", -- 3672 - 0xe58  :    0 - 0x0 -- plane 1
    "00000000", -- 3673 - 0xe59  :    0 - 0x0
    "00000000", -- 3674 - 0xe5a  :    0 - 0x0
    "00000000", -- 3675 - 0xe5b  :    0 - 0x0
    "00000000", -- 3676 - 0xe5c  :    0 - 0x0
    "00000000", -- 3677 - 0xe5d  :    0 - 0x0
    "00000000", -- 3678 - 0xe5e  :    0 - 0x0
    "00000000", -- 3679 - 0xe5f  :    0 - 0x0
    "00000000", -- 3680 - 0xe60  :    0 - 0x0 -- Background 0xe6
    "00000000", -- 3681 - 0xe61  :    0 - 0x0
    "00000000", -- 3682 - 0xe62  :    0 - 0x0
    "00000000", -- 3683 - 0xe63  :    0 - 0x0
    "00000000", -- 3684 - 0xe64  :    0 - 0x0
    "00000000", -- 3685 - 0xe65  :    0 - 0x0
    "00000000", -- 3686 - 0xe66  :    0 - 0x0
    "00000000", -- 3687 - 0xe67  :    0 - 0x0
    "00000000", -- 3688 - 0xe68  :    0 - 0x0 -- plane 1
    "00000000", -- 3689 - 0xe69  :    0 - 0x0
    "00000000", -- 3690 - 0xe6a  :    0 - 0x0
    "00000000", -- 3691 - 0xe6b  :    0 - 0x0
    "00000000", -- 3692 - 0xe6c  :    0 - 0x0
    "00000000", -- 3693 - 0xe6d  :    0 - 0x0
    "00000000", -- 3694 - 0xe6e  :    0 - 0x0
    "00000000", -- 3695 - 0xe6f  :    0 - 0x0
    "00000000", -- 3696 - 0xe70  :    0 - 0x0 -- Background 0xe7
    "00000000", -- 3697 - 0xe71  :    0 - 0x0
    "00000000", -- 3698 - 0xe72  :    0 - 0x0
    "00000000", -- 3699 - 0xe73  :    0 - 0x0
    "00000000", -- 3700 - 0xe74  :    0 - 0x0
    "00000000", -- 3701 - 0xe75  :    0 - 0x0
    "00000000", -- 3702 - 0xe76  :    0 - 0x0
    "00000000", -- 3703 - 0xe77  :    0 - 0x0
    "00000000", -- 3704 - 0xe78  :    0 - 0x0 -- plane 1
    "00000000", -- 3705 - 0xe79  :    0 - 0x0
    "00000000", -- 3706 - 0xe7a  :    0 - 0x0
    "00000000", -- 3707 - 0xe7b  :    0 - 0x0
    "00000000", -- 3708 - 0xe7c  :    0 - 0x0
    "00000000", -- 3709 - 0xe7d  :    0 - 0x0
    "00000000", -- 3710 - 0xe7e  :    0 - 0x0
    "00000000", -- 3711 - 0xe7f  :    0 - 0x0
    "00000000", -- 3712 - 0xe80  :    0 - 0x0 -- Background 0xe8
    "00000000", -- 3713 - 0xe81  :    0 - 0x0
    "00000000", -- 3714 - 0xe82  :    0 - 0x0
    "00000000", -- 3715 - 0xe83  :    0 - 0x0
    "00000000", -- 3716 - 0xe84  :    0 - 0x0
    "00000000", -- 3717 - 0xe85  :    0 - 0x0
    "00000000", -- 3718 - 0xe86  :    0 - 0x0
    "00000000", -- 3719 - 0xe87  :    0 - 0x0
    "00000000", -- 3720 - 0xe88  :    0 - 0x0 -- plane 1
    "00000000", -- 3721 - 0xe89  :    0 - 0x0
    "00000000", -- 3722 - 0xe8a  :    0 - 0x0
    "00000000", -- 3723 - 0xe8b  :    0 - 0x0
    "00000000", -- 3724 - 0xe8c  :    0 - 0x0
    "00000000", -- 3725 - 0xe8d  :    0 - 0x0
    "00000000", -- 3726 - 0xe8e  :    0 - 0x0
    "00000000", -- 3727 - 0xe8f  :    0 - 0x0
    "00000000", -- 3728 - 0xe90  :    0 - 0x0 -- Background 0xe9
    "00000000", -- 3729 - 0xe91  :    0 - 0x0
    "00000000", -- 3730 - 0xe92  :    0 - 0x0
    "00000000", -- 3731 - 0xe93  :    0 - 0x0
    "00000000", -- 3732 - 0xe94  :    0 - 0x0
    "00000000", -- 3733 - 0xe95  :    0 - 0x0
    "00000000", -- 3734 - 0xe96  :    0 - 0x0
    "00000000", -- 3735 - 0xe97  :    0 - 0x0
    "00000000", -- 3736 - 0xe98  :    0 - 0x0 -- plane 1
    "00000000", -- 3737 - 0xe99  :    0 - 0x0
    "00000000", -- 3738 - 0xe9a  :    0 - 0x0
    "00000000", -- 3739 - 0xe9b  :    0 - 0x0
    "00000000", -- 3740 - 0xe9c  :    0 - 0x0
    "00000000", -- 3741 - 0xe9d  :    0 - 0x0
    "00000000", -- 3742 - 0xe9e  :    0 - 0x0
    "00000000", -- 3743 - 0xe9f  :    0 - 0x0
    "00000000", -- 3744 - 0xea0  :    0 - 0x0 -- Background 0xea
    "00000000", -- 3745 - 0xea1  :    0 - 0x0
    "00000000", -- 3746 - 0xea2  :    0 - 0x0
    "00000000", -- 3747 - 0xea3  :    0 - 0x0
    "00000000", -- 3748 - 0xea4  :    0 - 0x0
    "00000000", -- 3749 - 0xea5  :    0 - 0x0
    "00000000", -- 3750 - 0xea6  :    0 - 0x0
    "00000000", -- 3751 - 0xea7  :    0 - 0x0
    "00000000", -- 3752 - 0xea8  :    0 - 0x0 -- plane 1
    "00000000", -- 3753 - 0xea9  :    0 - 0x0
    "00000000", -- 3754 - 0xeaa  :    0 - 0x0
    "00000000", -- 3755 - 0xeab  :    0 - 0x0
    "00000000", -- 3756 - 0xeac  :    0 - 0x0
    "00000000", -- 3757 - 0xead  :    0 - 0x0
    "00000000", -- 3758 - 0xeae  :    0 - 0x0
    "00000000", -- 3759 - 0xeaf  :    0 - 0x0
    "00000000", -- 3760 - 0xeb0  :    0 - 0x0 -- Background 0xeb
    "00000000", -- 3761 - 0xeb1  :    0 - 0x0
    "00000000", -- 3762 - 0xeb2  :    0 - 0x0
    "00000000", -- 3763 - 0xeb3  :    0 - 0x0
    "00000000", -- 3764 - 0xeb4  :    0 - 0x0
    "00000000", -- 3765 - 0xeb5  :    0 - 0x0
    "00000000", -- 3766 - 0xeb6  :    0 - 0x0
    "00000000", -- 3767 - 0xeb7  :    0 - 0x0
    "00000000", -- 3768 - 0xeb8  :    0 - 0x0 -- plane 1
    "00000000", -- 3769 - 0xeb9  :    0 - 0x0
    "00000000", -- 3770 - 0xeba  :    0 - 0x0
    "00000000", -- 3771 - 0xebb  :    0 - 0x0
    "00000000", -- 3772 - 0xebc  :    0 - 0x0
    "00000000", -- 3773 - 0xebd  :    0 - 0x0
    "00000000", -- 3774 - 0xebe  :    0 - 0x0
    "00000000", -- 3775 - 0xebf  :    0 - 0x0
    "00000000", -- 3776 - 0xec0  :    0 - 0x0 -- Background 0xec
    "00000000", -- 3777 - 0xec1  :    0 - 0x0
    "00000000", -- 3778 - 0xec2  :    0 - 0x0
    "00000000", -- 3779 - 0xec3  :    0 - 0x0
    "00000000", -- 3780 - 0xec4  :    0 - 0x0
    "00000000", -- 3781 - 0xec5  :    0 - 0x0
    "00000000", -- 3782 - 0xec6  :    0 - 0x0
    "00000000", -- 3783 - 0xec7  :    0 - 0x0
    "00000000", -- 3784 - 0xec8  :    0 - 0x0 -- plane 1
    "00000000", -- 3785 - 0xec9  :    0 - 0x0
    "00000000", -- 3786 - 0xeca  :    0 - 0x0
    "00000000", -- 3787 - 0xecb  :    0 - 0x0
    "00000000", -- 3788 - 0xecc  :    0 - 0x0
    "00000000", -- 3789 - 0xecd  :    0 - 0x0
    "00000000", -- 3790 - 0xece  :    0 - 0x0
    "00000000", -- 3791 - 0xecf  :    0 - 0x0
    "00000000", -- 3792 - 0xed0  :    0 - 0x0 -- Background 0xed
    "00000000", -- 3793 - 0xed1  :    0 - 0x0
    "00000000", -- 3794 - 0xed2  :    0 - 0x0
    "00000000", -- 3795 - 0xed3  :    0 - 0x0
    "00000000", -- 3796 - 0xed4  :    0 - 0x0
    "00000000", -- 3797 - 0xed5  :    0 - 0x0
    "00000000", -- 3798 - 0xed6  :    0 - 0x0
    "00000000", -- 3799 - 0xed7  :    0 - 0x0
    "00000000", -- 3800 - 0xed8  :    0 - 0x0 -- plane 1
    "00000000", -- 3801 - 0xed9  :    0 - 0x0
    "00000000", -- 3802 - 0xeda  :    0 - 0x0
    "00000000", -- 3803 - 0xedb  :    0 - 0x0
    "00000000", -- 3804 - 0xedc  :    0 - 0x0
    "00000000", -- 3805 - 0xedd  :    0 - 0x0
    "00000000", -- 3806 - 0xede  :    0 - 0x0
    "00000000", -- 3807 - 0xedf  :    0 - 0x0
    "00000000", -- 3808 - 0xee0  :    0 - 0x0 -- Background 0xee
    "00000000", -- 3809 - 0xee1  :    0 - 0x0
    "00000000", -- 3810 - 0xee2  :    0 - 0x0
    "00000000", -- 3811 - 0xee3  :    0 - 0x0
    "00000000", -- 3812 - 0xee4  :    0 - 0x0
    "00000000", -- 3813 - 0xee5  :    0 - 0x0
    "00000000", -- 3814 - 0xee6  :    0 - 0x0
    "00000000", -- 3815 - 0xee7  :    0 - 0x0
    "00000000", -- 3816 - 0xee8  :    0 - 0x0 -- plane 1
    "00000000", -- 3817 - 0xee9  :    0 - 0x0
    "00000000", -- 3818 - 0xeea  :    0 - 0x0
    "00000000", -- 3819 - 0xeeb  :    0 - 0x0
    "00000000", -- 3820 - 0xeec  :    0 - 0x0
    "00000000", -- 3821 - 0xeed  :    0 - 0x0
    "00000000", -- 3822 - 0xeee  :    0 - 0x0
    "00000000", -- 3823 - 0xeef  :    0 - 0x0
    "00000000", -- 3824 - 0xef0  :    0 - 0x0 -- Background 0xef
    "00000000", -- 3825 - 0xef1  :    0 - 0x0
    "00000000", -- 3826 - 0xef2  :    0 - 0x0
    "00000000", -- 3827 - 0xef3  :    0 - 0x0
    "00000000", -- 3828 - 0xef4  :    0 - 0x0
    "00000000", -- 3829 - 0xef5  :    0 - 0x0
    "00000000", -- 3830 - 0xef6  :    0 - 0x0
    "00000000", -- 3831 - 0xef7  :    0 - 0x0
    "00000000", -- 3832 - 0xef8  :    0 - 0x0 -- plane 1
    "00000000", -- 3833 - 0xef9  :    0 - 0x0
    "00000000", -- 3834 - 0xefa  :    0 - 0x0
    "00000000", -- 3835 - 0xefb  :    0 - 0x0
    "00000000", -- 3836 - 0xefc  :    0 - 0x0
    "00000000", -- 3837 - 0xefd  :    0 - 0x0
    "00000000", -- 3838 - 0xefe  :    0 - 0x0
    "00000000", -- 3839 - 0xeff  :    0 - 0x0
    "00000000", -- 3840 - 0xf00  :    0 - 0x0 -- Background 0xf0
    "00000000", -- 3841 - 0xf01  :    0 - 0x0
    "00000000", -- 3842 - 0xf02  :    0 - 0x0
    "00000000", -- 3843 - 0xf03  :    0 - 0x0
    "00000000", -- 3844 - 0xf04  :    0 - 0x0
    "00000000", -- 3845 - 0xf05  :    0 - 0x0
    "00000000", -- 3846 - 0xf06  :    0 - 0x0
    "00000000", -- 3847 - 0xf07  :    0 - 0x0
    "00000000", -- 3848 - 0xf08  :    0 - 0x0 -- plane 1
    "00000000", -- 3849 - 0xf09  :    0 - 0x0
    "00000000", -- 3850 - 0xf0a  :    0 - 0x0
    "00000000", -- 3851 - 0xf0b  :    0 - 0x0
    "00000000", -- 3852 - 0xf0c  :    0 - 0x0
    "00000000", -- 3853 - 0xf0d  :    0 - 0x0
    "00000000", -- 3854 - 0xf0e  :    0 - 0x0
    "00000000", -- 3855 - 0xf0f  :    0 - 0x0
    "00000000", -- 3856 - 0xf10  :    0 - 0x0 -- Background 0xf1
    "00000000", -- 3857 - 0xf11  :    0 - 0x0
    "00000000", -- 3858 - 0xf12  :    0 - 0x0
    "00000000", -- 3859 - 0xf13  :    0 - 0x0
    "00000000", -- 3860 - 0xf14  :    0 - 0x0
    "00000000", -- 3861 - 0xf15  :    0 - 0x0
    "00000000", -- 3862 - 0xf16  :    0 - 0x0
    "00000000", -- 3863 - 0xf17  :    0 - 0x0
    "00000000", -- 3864 - 0xf18  :    0 - 0x0 -- plane 1
    "00000000", -- 3865 - 0xf19  :    0 - 0x0
    "00000000", -- 3866 - 0xf1a  :    0 - 0x0
    "00000000", -- 3867 - 0xf1b  :    0 - 0x0
    "00000000", -- 3868 - 0xf1c  :    0 - 0x0
    "00000000", -- 3869 - 0xf1d  :    0 - 0x0
    "00000000", -- 3870 - 0xf1e  :    0 - 0x0
    "00000000", -- 3871 - 0xf1f  :    0 - 0x0
    "00000000", -- 3872 - 0xf20  :    0 - 0x0 -- Background 0xf2
    "00000000", -- 3873 - 0xf21  :    0 - 0x0
    "00000000", -- 3874 - 0xf22  :    0 - 0x0
    "00000000", -- 3875 - 0xf23  :    0 - 0x0
    "00000000", -- 3876 - 0xf24  :    0 - 0x0
    "00000000", -- 3877 - 0xf25  :    0 - 0x0
    "00000000", -- 3878 - 0xf26  :    0 - 0x0
    "00000000", -- 3879 - 0xf27  :    0 - 0x0
    "00000000", -- 3880 - 0xf28  :    0 - 0x0 -- plane 1
    "00000000", -- 3881 - 0xf29  :    0 - 0x0
    "00000000", -- 3882 - 0xf2a  :    0 - 0x0
    "00000000", -- 3883 - 0xf2b  :    0 - 0x0
    "00000000", -- 3884 - 0xf2c  :    0 - 0x0
    "00000000", -- 3885 - 0xf2d  :    0 - 0x0
    "00000000", -- 3886 - 0xf2e  :    0 - 0x0
    "00000000", -- 3887 - 0xf2f  :    0 - 0x0
    "00000000", -- 3888 - 0xf30  :    0 - 0x0 -- Background 0xf3
    "00000000", -- 3889 - 0xf31  :    0 - 0x0
    "00000000", -- 3890 - 0xf32  :    0 - 0x0
    "00000000", -- 3891 - 0xf33  :    0 - 0x0
    "00000000", -- 3892 - 0xf34  :    0 - 0x0
    "00000000", -- 3893 - 0xf35  :    0 - 0x0
    "00000000", -- 3894 - 0xf36  :    0 - 0x0
    "00000000", -- 3895 - 0xf37  :    0 - 0x0
    "00000000", -- 3896 - 0xf38  :    0 - 0x0 -- plane 1
    "00000000", -- 3897 - 0xf39  :    0 - 0x0
    "00000000", -- 3898 - 0xf3a  :    0 - 0x0
    "00000000", -- 3899 - 0xf3b  :    0 - 0x0
    "00000000", -- 3900 - 0xf3c  :    0 - 0x0
    "00000000", -- 3901 - 0xf3d  :    0 - 0x0
    "00000000", -- 3902 - 0xf3e  :    0 - 0x0
    "00000000", -- 3903 - 0xf3f  :    0 - 0x0
    "00000000", -- 3904 - 0xf40  :    0 - 0x0 -- Background 0xf4
    "00000000", -- 3905 - 0xf41  :    0 - 0x0
    "00000000", -- 3906 - 0xf42  :    0 - 0x0
    "00000000", -- 3907 - 0xf43  :    0 - 0x0
    "00000000", -- 3908 - 0xf44  :    0 - 0x0
    "00000000", -- 3909 - 0xf45  :    0 - 0x0
    "00000000", -- 3910 - 0xf46  :    0 - 0x0
    "00000000", -- 3911 - 0xf47  :    0 - 0x0
    "00000000", -- 3912 - 0xf48  :    0 - 0x0 -- plane 1
    "00000000", -- 3913 - 0xf49  :    0 - 0x0
    "00000000", -- 3914 - 0xf4a  :    0 - 0x0
    "00000000", -- 3915 - 0xf4b  :    0 - 0x0
    "00000000", -- 3916 - 0xf4c  :    0 - 0x0
    "00000000", -- 3917 - 0xf4d  :    0 - 0x0
    "00000000", -- 3918 - 0xf4e  :    0 - 0x0
    "00000000", -- 3919 - 0xf4f  :    0 - 0x0
    "00000000", -- 3920 - 0xf50  :    0 - 0x0 -- Background 0xf5
    "00000000", -- 3921 - 0xf51  :    0 - 0x0
    "00000000", -- 3922 - 0xf52  :    0 - 0x0
    "00000000", -- 3923 - 0xf53  :    0 - 0x0
    "00000000", -- 3924 - 0xf54  :    0 - 0x0
    "00000000", -- 3925 - 0xf55  :    0 - 0x0
    "00000000", -- 3926 - 0xf56  :    0 - 0x0
    "00000000", -- 3927 - 0xf57  :    0 - 0x0
    "00000000", -- 3928 - 0xf58  :    0 - 0x0 -- plane 1
    "00000000", -- 3929 - 0xf59  :    0 - 0x0
    "00000000", -- 3930 - 0xf5a  :    0 - 0x0
    "00000000", -- 3931 - 0xf5b  :    0 - 0x0
    "00000000", -- 3932 - 0xf5c  :    0 - 0x0
    "00000000", -- 3933 - 0xf5d  :    0 - 0x0
    "00000000", -- 3934 - 0xf5e  :    0 - 0x0
    "00000000", -- 3935 - 0xf5f  :    0 - 0x0
    "00000000", -- 3936 - 0xf60  :    0 - 0x0 -- Background 0xf6
    "00000000", -- 3937 - 0xf61  :    0 - 0x0
    "00000000", -- 3938 - 0xf62  :    0 - 0x0
    "00000000", -- 3939 - 0xf63  :    0 - 0x0
    "00000000", -- 3940 - 0xf64  :    0 - 0x0
    "00000000", -- 3941 - 0xf65  :    0 - 0x0
    "00000000", -- 3942 - 0xf66  :    0 - 0x0
    "00000000", -- 3943 - 0xf67  :    0 - 0x0
    "00000000", -- 3944 - 0xf68  :    0 - 0x0 -- plane 1
    "00000000", -- 3945 - 0xf69  :    0 - 0x0
    "00000000", -- 3946 - 0xf6a  :    0 - 0x0
    "00000000", -- 3947 - 0xf6b  :    0 - 0x0
    "00000000", -- 3948 - 0xf6c  :    0 - 0x0
    "00000000", -- 3949 - 0xf6d  :    0 - 0x0
    "00000000", -- 3950 - 0xf6e  :    0 - 0x0
    "00000000", -- 3951 - 0xf6f  :    0 - 0x0
    "00000000", -- 3952 - 0xf70  :    0 - 0x0 -- Background 0xf7
    "00000000", -- 3953 - 0xf71  :    0 - 0x0
    "00000000", -- 3954 - 0xf72  :    0 - 0x0
    "00000000", -- 3955 - 0xf73  :    0 - 0x0
    "00000000", -- 3956 - 0xf74  :    0 - 0x0
    "00000000", -- 3957 - 0xf75  :    0 - 0x0
    "00000000", -- 3958 - 0xf76  :    0 - 0x0
    "00000000", -- 3959 - 0xf77  :    0 - 0x0
    "00000000", -- 3960 - 0xf78  :    0 - 0x0 -- plane 1
    "00000000", -- 3961 - 0xf79  :    0 - 0x0
    "00000000", -- 3962 - 0xf7a  :    0 - 0x0
    "00000000", -- 3963 - 0xf7b  :    0 - 0x0
    "00000000", -- 3964 - 0xf7c  :    0 - 0x0
    "00000000", -- 3965 - 0xf7d  :    0 - 0x0
    "00000000", -- 3966 - 0xf7e  :    0 - 0x0
    "00000000", -- 3967 - 0xf7f  :    0 - 0x0
    "00000000", -- 3968 - 0xf80  :    0 - 0x0 -- Background 0xf8
    "00000000", -- 3969 - 0xf81  :    0 - 0x0
    "00000000", -- 3970 - 0xf82  :    0 - 0x0
    "00000000", -- 3971 - 0xf83  :    0 - 0x0
    "00000000", -- 3972 - 0xf84  :    0 - 0x0
    "00000000", -- 3973 - 0xf85  :    0 - 0x0
    "00000000", -- 3974 - 0xf86  :    0 - 0x0
    "00000000", -- 3975 - 0xf87  :    0 - 0x0
    "00000000", -- 3976 - 0xf88  :    0 - 0x0 -- plane 1
    "00000000", -- 3977 - 0xf89  :    0 - 0x0
    "00000000", -- 3978 - 0xf8a  :    0 - 0x0
    "00000000", -- 3979 - 0xf8b  :    0 - 0x0
    "00000000", -- 3980 - 0xf8c  :    0 - 0x0
    "00000000", -- 3981 - 0xf8d  :    0 - 0x0
    "00000000", -- 3982 - 0xf8e  :    0 - 0x0
    "00000000", -- 3983 - 0xf8f  :    0 - 0x0
    "00000000", -- 3984 - 0xf90  :    0 - 0x0 -- Background 0xf9
    "00000000", -- 3985 - 0xf91  :    0 - 0x0
    "00000000", -- 3986 - 0xf92  :    0 - 0x0
    "00000000", -- 3987 - 0xf93  :    0 - 0x0
    "00000000", -- 3988 - 0xf94  :    0 - 0x0
    "00000000", -- 3989 - 0xf95  :    0 - 0x0
    "00000000", -- 3990 - 0xf96  :    0 - 0x0
    "00000000", -- 3991 - 0xf97  :    0 - 0x0
    "00000000", -- 3992 - 0xf98  :    0 - 0x0 -- plane 1
    "00000000", -- 3993 - 0xf99  :    0 - 0x0
    "00000000", -- 3994 - 0xf9a  :    0 - 0x0
    "00000000", -- 3995 - 0xf9b  :    0 - 0x0
    "00000000", -- 3996 - 0xf9c  :    0 - 0x0
    "00000000", -- 3997 - 0xf9d  :    0 - 0x0
    "00000000", -- 3998 - 0xf9e  :    0 - 0x0
    "00000000", -- 3999 - 0xf9f  :    0 - 0x0
    "00000000", -- 4000 - 0xfa0  :    0 - 0x0 -- Background 0xfa
    "00000000", -- 4001 - 0xfa1  :    0 - 0x0
    "00000000", -- 4002 - 0xfa2  :    0 - 0x0
    "00000000", -- 4003 - 0xfa3  :    0 - 0x0
    "00000000", -- 4004 - 0xfa4  :    0 - 0x0
    "00000000", -- 4005 - 0xfa5  :    0 - 0x0
    "00000000", -- 4006 - 0xfa6  :    0 - 0x0
    "00000000", -- 4007 - 0xfa7  :    0 - 0x0
    "00000000", -- 4008 - 0xfa8  :    0 - 0x0 -- plane 1
    "00000000", -- 4009 - 0xfa9  :    0 - 0x0
    "00000000", -- 4010 - 0xfaa  :    0 - 0x0
    "00000000", -- 4011 - 0xfab  :    0 - 0x0
    "00000000", -- 4012 - 0xfac  :    0 - 0x0
    "00000000", -- 4013 - 0xfad  :    0 - 0x0
    "00000000", -- 4014 - 0xfae  :    0 - 0x0
    "00000000", -- 4015 - 0xfaf  :    0 - 0x0
    "00000000", -- 4016 - 0xfb0  :    0 - 0x0 -- Background 0xfb
    "00000000", -- 4017 - 0xfb1  :    0 - 0x0
    "00000000", -- 4018 - 0xfb2  :    0 - 0x0
    "00000000", -- 4019 - 0xfb3  :    0 - 0x0
    "00000000", -- 4020 - 0xfb4  :    0 - 0x0
    "00000000", -- 4021 - 0xfb5  :    0 - 0x0
    "00000000", -- 4022 - 0xfb6  :    0 - 0x0
    "00000000", -- 4023 - 0xfb7  :    0 - 0x0
    "00000000", -- 4024 - 0xfb8  :    0 - 0x0 -- plane 1
    "00000000", -- 4025 - 0xfb9  :    0 - 0x0
    "00000000", -- 4026 - 0xfba  :    0 - 0x0
    "00000000", -- 4027 - 0xfbb  :    0 - 0x0
    "00000000", -- 4028 - 0xfbc  :    0 - 0x0
    "00000000", -- 4029 - 0xfbd  :    0 - 0x0
    "00000000", -- 4030 - 0xfbe  :    0 - 0x0
    "00000000", -- 4031 - 0xfbf  :    0 - 0x0
    "00000000", -- 4032 - 0xfc0  :    0 - 0x0 -- Background 0xfc
    "00000000", -- 4033 - 0xfc1  :    0 - 0x0
    "10001110", -- 4034 - 0xfc2  :  142 - 0x8e
    "10001010", -- 4035 - 0xfc3  :  138 - 0x8a
    "10001010", -- 4036 - 0xfc4  :  138 - 0x8a
    "10001010", -- 4037 - 0xfc5  :  138 - 0x8a
    "10001010", -- 4038 - 0xfc6  :  138 - 0x8a
    "11101110", -- 4039 - 0xfc7  :  238 - 0xee
    "00000000", -- 4040 - 0xfc8  :    0 - 0x0 -- plane 1
    "00000000", -- 4041 - 0xfc9  :    0 - 0x0
    "00000000", -- 4042 - 0xfca  :    0 - 0x0
    "00000000", -- 4043 - 0xfcb  :    0 - 0x0
    "00000000", -- 4044 - 0xfcc  :    0 - 0x0
    "00000000", -- 4045 - 0xfcd  :    0 - 0x0
    "00000000", -- 4046 - 0xfce  :    0 - 0x0
    "00000000", -- 4047 - 0xfcf  :    0 - 0x0
    "00000000", -- 4048 - 0xfd0  :    0 - 0x0 -- Background 0xfd
    "00000000", -- 4049 - 0xfd1  :    0 - 0x0
    "01001100", -- 4050 - 0xfd2  :   76 - 0x4c
    "10101010", -- 4051 - 0xfd3  :  170 - 0xaa
    "10101010", -- 4052 - 0xfd4  :  170 - 0xaa
    "11101010", -- 4053 - 0xfd5  :  234 - 0xea
    "10101010", -- 4054 - 0xfd6  :  170 - 0xaa
    "10101100", -- 4055 - 0xfd7  :  172 - 0xac
    "00000000", -- 4056 - 0xfd8  :    0 - 0x0 -- plane 1
    "00000000", -- 4057 - 0xfd9  :    0 - 0x0
    "00000000", -- 4058 - 0xfda  :    0 - 0x0
    "00000000", -- 4059 - 0xfdb  :    0 - 0x0
    "00000000", -- 4060 - 0xfdc  :    0 - 0x0
    "00000000", -- 4061 - 0xfdd  :    0 - 0x0
    "00000000", -- 4062 - 0xfde  :    0 - 0x0
    "00000000", -- 4063 - 0xfdf  :    0 - 0x0
    "00000000", -- 4064 - 0xfe0  :    0 - 0x0 -- Background 0xfe
    "00000000", -- 4065 - 0xfe1  :    0 - 0x0
    "11101100", -- 4066 - 0xfe2  :  236 - 0xec
    "01001010", -- 4067 - 0xfe3  :   74 - 0x4a
    "01001010", -- 4068 - 0xfe4  :   74 - 0x4a
    "01001010", -- 4069 - 0xfe5  :   74 - 0x4a
    "01001010", -- 4070 - 0xfe6  :   74 - 0x4a
    "11101010", -- 4071 - 0xfe7  :  234 - 0xea
    "00000000", -- 4072 - 0xfe8  :    0 - 0x0 -- plane 1
    "00000000", -- 4073 - 0xfe9  :    0 - 0x0
    "00000000", -- 4074 - 0xfea  :    0 - 0x0
    "00000000", -- 4075 - 0xfeb  :    0 - 0x0
    "00000000", -- 4076 - 0xfec  :    0 - 0x0
    "00000000", -- 4077 - 0xfed  :    0 - 0x0
    "00000000", -- 4078 - 0xfee  :    0 - 0x0
    "00000000", -- 4079 - 0xfef  :    0 - 0x0
    "00000000", -- 4080 - 0xff0  :    0 - 0x0 -- Background 0xff
    "00000000", -- 4081 - 0xff1  :    0 - 0x0
    "01100000", -- 4082 - 0xff2  :   96 - 0x60
    "10001000", -- 4083 - 0xff3  :  136 - 0x88
    "10100000", -- 4084 - 0xff4  :  160 - 0xa0
    "10100000", -- 4085 - 0xff5  :  160 - 0xa0
    "10101000", -- 4086 - 0xff6  :  168 - 0xa8
    "01000000", -- 4087 - 0xff7  :   64 - 0x40
    "00000000", -- 4088 - 0xff8  :    0 - 0x0 -- plane 1
    "00000000", -- 4089 - 0xff9  :    0 - 0x0
    "00000000", -- 4090 - 0xffa  :    0 - 0x0
    "00000000", -- 4091 - 0xffb  :    0 - 0x0
    "00000000", -- 4092 - 0xffc  :    0 - 0x0
    "00000000", -- 4093 - 0xffd  :    0 - 0x0
    "00000000", -- 4094 - 0xffe  :    0 - 0x0
    "00000000"  -- 4095 - 0xfff  :    0 - 0x0
    );
begin
  addr_int <= to_integer(unsigned(addr));
  --P_ROM: process(clk)
  --begin
  --  if clk'event and clk='1' then
      dout <= table_mem(addr_int);
  --  end if;
  --end process;
end BEHAVIORAL;
